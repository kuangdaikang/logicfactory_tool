// Benchmark "mem_ctrl" written by ABC on Fri Feb 25 15:09:03 2022

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_,
    new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_,
    new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_,
    new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_,
    new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_,
    new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_,
    new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_,
    new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_,
    new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_,
    new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_,
    new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_,
    new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_,
    new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_,
    new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_,
    new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_,
    new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_,
    new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_,
    new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_,
    new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_,
    new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_,
    new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_,
    new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_,
    new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_,
    new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_,
    new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_,
    new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_,
    new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_,
    new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_,
    new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5071_, new_n5072_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_,
    new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_,
    new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_,
    new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_,
    new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_,
    new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_,
    new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_,
    new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_,
    new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_,
    new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_,
    new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_,
    new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_,
    new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_,
    new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_,
    new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_,
    new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_,
    new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_,
    new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_,
    new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_,
    new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_,
    new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_,
    new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_,
    new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_,
    new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_,
    new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_,
    new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_,
    new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_,
    new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_,
    new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_,
    new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_,
    new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_,
    new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6275_, new_n6276_, new_n6277_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_,
    new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_,
    new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_,
    new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_,
    new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_,
    new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_,
    new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6921_,
    new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_,
    new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_,
    new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_,
    new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_,
    new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_,
    new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_,
    new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_,
    new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_,
    new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_,
    new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_,
    new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_,
    new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_,
    new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_,
    new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_,
    new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_,
    new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_,
    new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_,
    new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_,
    new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_,
    new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_,
    new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_,
    new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_,
    new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7353_, new_n7354_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7406_, new_n7407_, new_n7408_,
    new_n7409_, new_n7411_, new_n7413_, new_n7415_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_,
    new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_,
    new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_,
    new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_,
    new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_,
    new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_,
    new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_,
    new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_,
    new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_,
    new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_,
    new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_,
    new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_,
    new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_,
    new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_,
    new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_,
    new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_,
    new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_,
    new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_,
    new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_,
    new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_,
    new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_,
    new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_,
    new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_,
    new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_,
    new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_,
    new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_,
    new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_,
    new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_,
    new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_,
    new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_,
    new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_,
    new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_,
    new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_,
    new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_,
    new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_,
    new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_,
    new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_,
    new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_,
    new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_,
    new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_,
    new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_,
    new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_,
    new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_,
    new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_,
    new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_,
    new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_,
    new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_,
    new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_,
    new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_,
    new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_,
    new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_,
    new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_,
    new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_,
    new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_,
    new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_,
    new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_,
    new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_,
    new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_,
    new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_,
    new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_,
    new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_,
    new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_,
    new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_,
    new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_,
    new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_,
    new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_,
    new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_,
    new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_,
    new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_,
    new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_,
    new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_,
    new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_,
    new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_,
    new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_,
    new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_,
    new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_,
    new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_,
    new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_,
    new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_,
    new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_, new_n8444_,
    new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_,
    new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_,
    new_n8457_, new_n8458_, new_n8459_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_,
    new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_,
    new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_,
    new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_,
    new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_,
    new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_,
    new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_,
    new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_,
    new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_,
    new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_,
    new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_,
    new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_,
    new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_,
    new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8878_,
    new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_,
    new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_,
    new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_,
    new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8974_, new_n8975_, new_n8976_,
    new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_,
    new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_,
    new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_,
    new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_,
    new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_,
    new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_,
    new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_,
    new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_,
    new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_,
    new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_,
    new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_,
    new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_,
    new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_,
    new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_,
    new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_,
    new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_,
    new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_,
    new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_,
    new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_,
    new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_,
    new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_,
    new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_,
    new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_,
    new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_,
    new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_,
    new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_,
    new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_,
    new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_,
    new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_,
    new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_,
    new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_,
    new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_,
    new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_,
    new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_,
    new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_,
    new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_,
    new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_,
    new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_,
    new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_,
    new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_,
    new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_,
    new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10040_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10073_,
    new_n10074_, new_n10075_, new_n10076_, new_n10077_, new_n10078_,
    new_n10079_, new_n10080_, new_n10081_, new_n10082_, new_n10083_,
    new_n10084_, new_n10085_, new_n10086_, new_n10087_, new_n10088_,
    new_n10089_, new_n10090_, new_n10091_, new_n10092_, new_n10093_,
    new_n10094_, new_n10095_, new_n10096_, new_n10097_, new_n10098_,
    new_n10099_, new_n10100_, new_n10101_, new_n10102_, new_n10103_,
    new_n10104_, new_n10105_, new_n10106_, new_n10107_, new_n10108_,
    new_n10109_, new_n10110_, new_n10111_, new_n10112_, new_n10113_,
    new_n10114_, new_n10115_, new_n10116_, new_n10117_, new_n10118_,
    new_n10119_, new_n10120_, new_n10121_, new_n10122_, new_n10123_,
    new_n10124_, new_n10125_, new_n10126_, new_n10127_, new_n10128_,
    new_n10129_, new_n10130_, new_n10131_, new_n10132_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10200_, new_n10201_,
    new_n10202_, new_n10203_, new_n10204_, new_n10205_, new_n10206_,
    new_n10207_, new_n10208_, new_n10209_, new_n10210_, new_n10211_,
    new_n10212_, new_n10213_, new_n10214_, new_n10215_, new_n10216_,
    new_n10217_, new_n10218_, new_n10219_, new_n10220_, new_n10221_,
    new_n10222_, new_n10223_, new_n10224_, new_n10225_, new_n10226_,
    new_n10227_, new_n10228_, new_n10229_, new_n10230_, new_n10231_,
    new_n10232_, new_n10233_, new_n10234_, new_n10235_, new_n10236_,
    new_n10237_, new_n10238_, new_n10239_, new_n10240_, new_n10241_,
    new_n10242_, new_n10243_, new_n10244_, new_n10245_, new_n10246_,
    new_n10247_, new_n10248_, new_n10249_, new_n10250_, new_n10251_,
    new_n10252_, new_n10253_, new_n10254_, new_n10255_, new_n10256_,
    new_n10257_, new_n10258_, new_n10259_, new_n10260_, new_n10261_,
    new_n10262_, new_n10263_, new_n10264_, new_n10265_, new_n10266_,
    new_n10267_, new_n10268_, new_n10269_, new_n10270_, new_n10271_,
    new_n10272_, new_n10273_, new_n10274_, new_n10275_, new_n10276_,
    new_n10277_, new_n10278_, new_n10279_, new_n10281_, new_n10282_,
    new_n10283_, new_n10284_, new_n10285_, new_n10286_, new_n10287_,
    new_n10288_, new_n10289_, new_n10290_, new_n10291_, new_n10292_,
    new_n10293_, new_n10295_, new_n10296_, new_n10297_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10303_,
    new_n10304_, new_n10305_, new_n10306_, new_n10307_, new_n10308_,
    new_n10309_, new_n10310_, new_n10311_, new_n10312_, new_n10313_,
    new_n10314_, new_n10315_, new_n10316_, new_n10317_, new_n10318_,
    new_n10319_, new_n10320_, new_n10321_, new_n10322_, new_n10323_,
    new_n10324_, new_n10325_, new_n10326_, new_n10327_, new_n10328_,
    new_n10329_, new_n10330_, new_n10331_, new_n10332_, new_n10333_,
    new_n10334_, new_n10335_, new_n10336_, new_n10337_, new_n10338_,
    new_n10339_, new_n10340_, new_n10341_, new_n10342_, new_n10343_,
    new_n10344_, new_n10345_, new_n10346_, new_n10347_, new_n10348_,
    new_n10349_, new_n10350_, new_n10351_, new_n10352_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10359_, new_n10360_, new_n10361_, new_n10362_, new_n10363_,
    new_n10364_, new_n10365_, new_n10366_, new_n10367_, new_n10368_,
    new_n10369_, new_n10370_, new_n10371_, new_n10372_, new_n10373_,
    new_n10374_, new_n10375_, new_n10376_, new_n10377_, new_n10378_,
    new_n10379_, new_n10380_, new_n10381_, new_n10382_, new_n10383_,
    new_n10384_, new_n10385_, new_n10386_, new_n10387_, new_n10388_,
    new_n10389_, new_n10390_, new_n10391_, new_n10392_, new_n10393_,
    new_n10394_, new_n10395_, new_n10396_, new_n10397_, new_n10398_,
    new_n10399_, new_n10400_, new_n10401_, new_n10402_, new_n10403_,
    new_n10404_, new_n10405_, new_n10406_, new_n10407_, new_n10408_,
    new_n10409_, new_n10410_, new_n10411_, new_n10412_, new_n10413_,
    new_n10414_, new_n10415_, new_n10416_, new_n10417_, new_n10418_,
    new_n10419_, new_n10420_, new_n10421_, new_n10422_, new_n10423_,
    new_n10424_, new_n10425_, new_n10426_, new_n10427_, new_n10428_,
    new_n10429_, new_n10430_, new_n10431_, new_n10432_, new_n10433_,
    new_n10434_, new_n10435_, new_n10436_, new_n10437_, new_n10438_,
    new_n10439_, new_n10440_, new_n10441_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10448_,
    new_n10449_, new_n10450_, new_n10451_, new_n10452_, new_n10453_,
    new_n10454_, new_n10455_, new_n10456_, new_n10457_, new_n10458_,
    new_n10459_, new_n10460_, new_n10461_, new_n10462_, new_n10463_,
    new_n10464_, new_n10465_, new_n10466_, new_n10467_, new_n10468_,
    new_n10469_, new_n10470_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10478_,
    new_n10479_, new_n10480_, new_n10481_, new_n10482_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10982_,
    new_n10983_, new_n10984_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11076_, new_n11077_,
    new_n11078_, new_n11079_, new_n11080_, new_n11081_, new_n11082_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11092_,
    new_n11093_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11102_, new_n11103_,
    new_n11104_, new_n11105_, new_n11106_, new_n11107_, new_n11108_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11307_, new_n11308_,
    new_n11309_, new_n11310_, new_n11311_, new_n11312_, new_n11313_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11325_,
    new_n11326_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11343_,
    new_n11344_, new_n11345_, new_n11346_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11369_, new_n11370_, new_n11371_, new_n11373_,
    new_n11374_, new_n11375_, new_n11376_, new_n11377_, new_n11378_,
    new_n11379_, new_n11380_, new_n11381_, new_n11382_, new_n11383_,
    new_n11384_, new_n11385_, new_n11386_, new_n11387_, new_n11388_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11436_, new_n11437_, new_n11438_,
    new_n11439_, new_n11440_, new_n11441_, new_n11442_, new_n11443_,
    new_n11444_, new_n11445_, new_n11446_, new_n11447_, new_n11448_,
    new_n11449_, new_n11450_, new_n11451_, new_n11452_, new_n11453_,
    new_n11454_, new_n11455_, new_n11456_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11510_, new_n11511_, new_n11512_, new_n11513_,
    new_n11514_, new_n11515_, new_n11516_, new_n11517_, new_n11518_,
    new_n11519_, new_n11520_, new_n11521_, new_n11522_, new_n11523_,
    new_n11524_, new_n11525_, new_n11526_, new_n11527_, new_n11528_,
    new_n11529_, new_n11530_, new_n11531_, new_n11532_, new_n11533_,
    new_n11534_, new_n11535_, new_n11536_, new_n11537_, new_n11538_,
    new_n11539_, new_n11540_, new_n11541_, new_n11542_, new_n11543_,
    new_n11544_, new_n11545_, new_n11546_, new_n11547_, new_n11548_,
    new_n11549_, new_n11550_, new_n11551_, new_n11552_, new_n11553_,
    new_n11554_, new_n11555_, new_n11556_, new_n11557_, new_n11558_,
    new_n11559_, new_n11560_, new_n11561_, new_n11562_, new_n11563_,
    new_n11564_, new_n11565_, new_n11566_, new_n11567_, new_n11568_,
    new_n11569_, new_n11570_, new_n11571_, new_n11572_, new_n11573_,
    new_n11574_, new_n11575_, new_n11576_, new_n11577_, new_n11578_,
    new_n11579_, new_n11580_, new_n11581_, new_n11582_, new_n11583_,
    new_n11584_, new_n11585_, new_n11586_, new_n11587_, new_n11588_,
    new_n11589_, new_n11590_, new_n11591_, new_n11592_, new_n11593_,
    new_n11594_, new_n11595_, new_n11596_, new_n11597_, new_n11598_,
    new_n11599_, new_n11600_, new_n11601_, new_n11602_, new_n11603_,
    new_n11604_, new_n11605_, new_n11606_, new_n11607_, new_n11608_,
    new_n11609_, new_n11610_, new_n11611_, new_n11612_, new_n11613_,
    new_n11614_, new_n11615_, new_n11616_, new_n11617_, new_n11618_,
    new_n11619_, new_n11620_, new_n11621_, new_n11622_, new_n11623_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11631_, new_n11632_, new_n11633_,
    new_n11634_, new_n11635_, new_n11636_, new_n11637_, new_n11638_,
    new_n11639_, new_n11640_, new_n11641_, new_n11642_, new_n11643_,
    new_n11644_, new_n11645_, new_n11646_, new_n11647_, new_n11648_,
    new_n11649_, new_n11650_, new_n11651_, new_n11652_, new_n11653_,
    new_n11654_, new_n11655_, new_n11656_, new_n11657_, new_n11658_,
    new_n11659_, new_n11660_, new_n11661_, new_n11663_, new_n11664_,
    new_n11665_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11671_, new_n11673_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12100_, new_n12101_,
    new_n12102_, new_n12103_, new_n12104_, new_n12105_, new_n12106_,
    new_n12107_, new_n12108_, new_n12109_, new_n12110_, new_n12111_,
    new_n12112_, new_n12113_, new_n12114_, new_n12115_, new_n12116_,
    new_n12117_, new_n12118_, new_n12119_, new_n12120_, new_n12121_,
    new_n12122_, new_n12123_, new_n12124_, new_n12125_, new_n12126_,
    new_n12127_, new_n12128_, new_n12129_, new_n12130_, new_n12131_,
    new_n12132_, new_n12133_, new_n12134_, new_n12135_, new_n12136_,
    new_n12137_, new_n12138_, new_n12139_, new_n12140_, new_n12141_,
    new_n12142_, new_n12143_, new_n12144_, new_n12145_, new_n12146_,
    new_n12147_, new_n12148_, new_n12149_, new_n12150_, new_n12151_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12158_, new_n12159_, new_n12160_, new_n12161_,
    new_n12162_, new_n12163_, new_n12164_, new_n12165_, new_n12166_,
    new_n12167_, new_n12168_, new_n12169_, new_n12170_, new_n12171_,
    new_n12172_, new_n12173_, new_n12174_, new_n12175_, new_n12176_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12536_, new_n12537_,
    new_n12538_, new_n12539_, new_n12540_, new_n12541_, new_n12542_,
    new_n12543_, new_n12544_, new_n12545_, new_n12546_, new_n12547_,
    new_n12548_, new_n12549_, new_n12550_, new_n12551_, new_n12552_,
    new_n12553_, new_n12554_, new_n12555_, new_n12556_, new_n12557_,
    new_n12558_, new_n12559_, new_n12560_, new_n12561_, new_n12562_,
    new_n12563_, new_n12564_, new_n12565_, new_n12566_, new_n12567_,
    new_n12568_, new_n12569_, new_n12570_, new_n12571_, new_n12572_,
    new_n12573_, new_n12574_, new_n12575_, new_n12576_, new_n12577_,
    new_n12578_, new_n12579_, new_n12580_, new_n12581_, new_n12582_,
    new_n12583_, new_n12584_, new_n12585_, new_n12586_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12593_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12599_, new_n12600_, new_n12601_, new_n12602_,
    new_n12603_, new_n12604_, new_n12605_, new_n12606_, new_n12607_,
    new_n12608_, new_n12609_, new_n12610_, new_n12611_, new_n12612_,
    new_n12613_, new_n12614_, new_n12615_, new_n12616_, new_n12617_,
    new_n12618_, new_n12619_, new_n12620_, new_n12621_, new_n12622_,
    new_n12623_, new_n12624_, new_n12625_, new_n12626_, new_n12627_,
    new_n12628_, new_n12629_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12636_, new_n12637_,
    new_n12638_, new_n12639_, new_n12640_, new_n12641_, new_n12642_,
    new_n12643_, new_n12644_, new_n12645_, new_n12646_, new_n12647_,
    new_n12648_, new_n12649_, new_n12650_, new_n12651_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12658_, new_n12659_, new_n12660_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12791_, new_n12792_,
    new_n12793_, new_n12794_, new_n12795_, new_n12796_, new_n12797_,
    new_n12798_, new_n12799_, new_n12800_, new_n12801_, new_n12802_,
    new_n12803_, new_n12804_, new_n12805_, new_n12806_, new_n12807_,
    new_n12808_, new_n12809_, new_n12810_, new_n12811_, new_n12812_,
    new_n12813_, new_n12814_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12822_,
    new_n12823_, new_n12824_, new_n12825_, new_n12826_, new_n12827_,
    new_n12828_, new_n12829_, new_n12830_, new_n12831_, new_n12832_,
    new_n12833_, new_n12834_, new_n12835_, new_n12836_, new_n12837_,
    new_n12838_, new_n12839_, new_n12840_, new_n12841_, new_n12842_,
    new_n12843_, new_n12844_, new_n12845_, new_n12846_, new_n12847_,
    new_n12848_, new_n12849_, new_n12850_, new_n12851_, new_n12852_,
    new_n12853_, new_n12854_, new_n12855_, new_n12856_, new_n12857_,
    new_n12858_, new_n12859_, new_n12860_, new_n12861_, new_n12862_,
    new_n12863_, new_n12864_, new_n12865_, new_n12866_, new_n12867_,
    new_n12868_, new_n12869_, new_n12870_, new_n12871_, new_n12872_,
    new_n12873_, new_n12874_, new_n12875_, new_n12876_, new_n12877_,
    new_n12878_, new_n12879_, new_n12880_, new_n12881_, new_n12882_,
    new_n12883_, new_n12884_, new_n12885_, new_n12886_, new_n12887_,
    new_n12888_, new_n12889_, new_n12890_, new_n12891_, new_n12892_,
    new_n12893_, new_n12894_, new_n12895_, new_n12896_, new_n12897_,
    new_n12898_, new_n12899_, new_n12900_, new_n12901_, new_n12902_,
    new_n12903_, new_n12904_, new_n12905_, new_n12906_, new_n12907_,
    new_n12908_, new_n12909_, new_n12910_, new_n12911_, new_n12912_,
    new_n12913_, new_n12914_, new_n12915_, new_n12916_, new_n12917_,
    new_n12918_, new_n12919_, new_n12920_, new_n12921_, new_n12922_,
    new_n12923_, new_n12924_, new_n12925_, new_n12926_, new_n12927_,
    new_n12928_, new_n12929_, new_n12930_, new_n12931_, new_n12932_,
    new_n12933_, new_n12934_, new_n12935_, new_n12936_, new_n12937_,
    new_n12938_, new_n12939_, new_n12940_, new_n12941_, new_n12942_,
    new_n12943_, new_n12944_, new_n12945_, new_n12946_, new_n12947_,
    new_n12948_, new_n12949_, new_n12950_, new_n12951_, new_n12952_,
    new_n12953_, new_n12954_, new_n12955_, new_n12956_, new_n12957_,
    new_n12958_, new_n12959_, new_n12960_, new_n12961_, new_n12962_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13009_, new_n13010_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13018_, new_n13019_, new_n13020_, new_n13021_, new_n13022_,
    new_n13023_, new_n13024_, new_n13025_, new_n13026_, new_n13027_,
    new_n13029_, new_n13030_, new_n13031_, new_n13032_, new_n13033_,
    new_n13034_, new_n13035_, new_n13036_, new_n13037_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13061_,
    new_n13062_, new_n13063_, new_n13064_, new_n13065_, new_n13067_,
    new_n13068_, new_n13069_, new_n13070_, new_n13072_, new_n13073_,
    new_n13074_, new_n13076_, new_n13077_, new_n13078_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13100_, new_n13101_,
    new_n13102_, new_n13103_, new_n13104_, new_n13105_, new_n13106_,
    new_n13107_, new_n13108_, new_n13110_, new_n13111_, new_n13112_,
    new_n13113_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13120_, new_n13121_, new_n13122_, new_n13123_,
    new_n13124_, new_n13125_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13146_,
    new_n13147_, new_n13148_, new_n13149_, new_n13150_, new_n13151_,
    new_n13152_, new_n13153_, new_n13154_, new_n13155_, new_n13156_,
    new_n13157_, new_n13158_, new_n13159_, new_n13160_, new_n13161_,
    new_n13162_, new_n13164_, new_n13165_, new_n13166_, new_n13167_,
    new_n13168_, new_n13169_, new_n13170_, new_n13171_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13178_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13185_, new_n13186_, new_n13187_, new_n13188_,
    new_n13189_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13206_,
    new_n13207_, new_n13208_, new_n13209_, new_n13210_, new_n13211_,
    new_n13212_, new_n13213_, new_n13214_, new_n13215_, new_n13216_,
    new_n13217_, new_n13218_, new_n13219_, new_n13220_, new_n13221_,
    new_n13222_, new_n13223_, new_n13224_, new_n13225_, new_n13226_,
    new_n13227_, new_n13228_, new_n13229_, new_n13230_, new_n13231_,
    new_n13232_, new_n13233_, new_n13234_, new_n13235_, new_n13236_,
    new_n13237_, new_n13238_, new_n13239_, new_n13240_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13245_, new_n13246_,
    new_n13247_, new_n13248_, new_n13249_, new_n13250_, new_n13251_,
    new_n13252_, new_n13253_, new_n13254_, new_n13255_, new_n13256_,
    new_n13257_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13262_, new_n13263_, new_n13264_, new_n13265_, new_n13266_,
    new_n13267_, new_n13268_, new_n13269_, new_n13270_, new_n13271_,
    new_n13272_, new_n13273_, new_n13274_, new_n13275_, new_n13276_,
    new_n13277_, new_n13278_, new_n13279_, new_n13280_, new_n13281_,
    new_n13283_, new_n13284_, new_n13285_, new_n13286_, new_n13287_,
    new_n13288_, new_n13289_, new_n13290_, new_n13291_, new_n13292_,
    new_n13293_, new_n13294_, new_n13295_, new_n13296_, new_n13297_,
    new_n13298_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_,
    new_n13359_, new_n13360_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13367_, new_n13368_,
    new_n13369_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13376_, new_n13377_, new_n13378_,
    new_n13379_, new_n13381_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13395_, new_n13396_,
    new_n13397_, new_n13398_, new_n13399_, new_n13400_, new_n13401_,
    new_n13402_, new_n13403_, new_n13404_, new_n13405_, new_n13406_,
    new_n13407_, new_n13409_, new_n13410_, new_n13411_, new_n13412_,
    new_n13413_, new_n13414_, new_n13415_, new_n13416_, new_n13417_,
    new_n13419_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13439_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13452_,
    new_n13453_, new_n13454_, new_n13455_, new_n13456_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13597_,
    new_n13598_, new_n13599_, new_n13600_, new_n13601_, new_n13602_,
    new_n13603_, new_n13604_, new_n13605_, new_n13606_, new_n13607_,
    new_n13608_, new_n13609_, new_n13610_, new_n13611_, new_n13612_,
    new_n13613_, new_n13614_, new_n13615_, new_n13616_, new_n13617_,
    new_n13618_, new_n13619_, new_n13620_, new_n13621_, new_n13622_,
    new_n13623_, new_n13624_, new_n13625_, new_n13626_, new_n13627_,
    new_n13628_, new_n13629_, new_n13630_, new_n13631_, new_n13632_,
    new_n13633_, new_n13634_, new_n13635_, new_n13636_, new_n13637_,
    new_n13638_, new_n13639_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13648_,
    new_n13649_, new_n13650_, new_n13651_, new_n13652_, new_n13653_,
    new_n13654_, new_n13655_, new_n13656_, new_n13657_, new_n13658_,
    new_n13659_, new_n13660_, new_n13661_, new_n13662_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13695_, new_n13696_, new_n13697_, new_n13698_, new_n13699_,
    new_n13700_, new_n13701_, new_n13702_, new_n13703_, new_n13704_,
    new_n13705_, new_n13706_, new_n13707_, new_n13708_, new_n13709_,
    new_n13710_, new_n13711_, new_n13712_, new_n13713_, new_n13714_,
    new_n13715_, new_n13716_, new_n13717_, new_n13718_, new_n13719_,
    new_n13720_, new_n13721_, new_n13722_, new_n13723_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13730_, new_n13731_, new_n13732_, new_n13733_, new_n13734_,
    new_n13735_, new_n13736_, new_n13737_, new_n13738_, new_n13739_,
    new_n13740_, new_n13741_, new_n13742_, new_n13743_, new_n13744_,
    new_n13745_, new_n13746_, new_n13747_, new_n13748_, new_n13749_,
    new_n13750_, new_n13751_, new_n13752_, new_n13753_, new_n13754_,
    new_n13755_, new_n13756_, new_n13757_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13766_, new_n13767_, new_n13768_, new_n13769_,
    new_n13770_, new_n13771_, new_n13772_, new_n13773_, new_n13774_,
    new_n13775_, new_n13776_, new_n13777_, new_n13778_, new_n13779_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13806_, new_n13807_, new_n13808_, new_n13809_,
    new_n13810_, new_n13811_, new_n13812_, new_n13813_, new_n13814_,
    new_n13815_, new_n13816_, new_n13817_, new_n13818_, new_n13819_,
    new_n13820_, new_n13821_, new_n13822_, new_n13823_, new_n13824_,
    new_n13825_, new_n13826_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13853_, new_n13854_,
    new_n13855_, new_n13856_, new_n13857_, new_n13858_, new_n13859_,
    new_n13860_, new_n13861_, new_n13862_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13871_, new_n13872_, new_n13873_, new_n13874_,
    new_n13875_, new_n13876_, new_n13877_, new_n13878_, new_n13879_,
    new_n13880_, new_n13881_, new_n13882_, new_n13883_, new_n13884_,
    new_n13885_, new_n13886_, new_n13887_, new_n13888_, new_n13889_,
    new_n13890_, new_n13891_, new_n13892_, new_n13893_, new_n13894_,
    new_n13895_, new_n13896_, new_n13897_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13904_,
    new_n13905_, new_n13906_, new_n13907_, new_n13908_, new_n13909_,
    new_n13910_, new_n13911_, new_n13912_, new_n13913_, new_n13914_,
    new_n13915_, new_n13916_, new_n13917_, new_n13918_, new_n13919_,
    new_n13920_, new_n13921_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13927_, new_n13928_, new_n13929_,
    new_n13930_, new_n13931_, new_n13932_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13963_, new_n13964_,
    new_n13965_, new_n13966_, new_n13967_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14763_, new_n14764_, new_n14765_, new_n14766_, new_n14767_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14831_, new_n14832_,
    new_n14833_, new_n14834_, new_n14835_, new_n14836_, new_n14837_,
    new_n14838_, new_n14839_, new_n14840_, new_n14841_, new_n14842_,
    new_n14843_, new_n14844_, new_n14845_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15315_, new_n15316_,
    new_n15317_, new_n15318_, new_n15319_, new_n15320_, new_n15321_,
    new_n15322_, new_n15323_, new_n15324_, new_n15325_, new_n15326_,
    new_n15327_, new_n15328_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15434_, new_n15435_, new_n15436_,
    new_n15437_, new_n15438_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15470_, new_n15471_,
    new_n15472_, new_n15473_, new_n15474_, new_n15475_, new_n15476_,
    new_n15477_, new_n15478_, new_n15479_, new_n15480_, new_n15481_,
    new_n15482_, new_n15483_, new_n15484_, new_n15485_, new_n15486_,
    new_n15487_, new_n15488_, new_n15489_, new_n15490_, new_n15491_,
    new_n15492_, new_n15493_, new_n15494_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15544_, new_n15545_, new_n15546_,
    new_n15547_, new_n15548_, new_n15549_, new_n15550_, new_n15551_,
    new_n15552_, new_n15553_, new_n15554_, new_n15555_, new_n15556_,
    new_n15557_, new_n15558_, new_n15559_, new_n15560_, new_n15561_,
    new_n15562_, new_n15563_, new_n15564_, new_n15565_, new_n15566_,
    new_n15567_, new_n15568_, new_n15569_, new_n15570_, new_n15571_,
    new_n15572_, new_n15573_, new_n15574_, new_n15575_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15580_, new_n15581_,
    new_n15582_, new_n15583_, new_n15584_, new_n15585_, new_n15586_,
    new_n15587_, new_n15588_, new_n15589_, new_n15590_, new_n15591_,
    new_n15592_, new_n15593_, new_n15594_, new_n15595_, new_n15596_,
    new_n15597_, new_n15598_, new_n15599_, new_n15600_, new_n15601_,
    new_n15602_, new_n15603_, new_n15604_, new_n15605_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15611_,
    new_n15612_, new_n15613_, new_n15614_, new_n15615_, new_n15616_,
    new_n15618_, new_n15619_, new_n15620_, new_n15621_, new_n15622_,
    new_n15623_, new_n15624_, new_n15625_, new_n15626_, new_n15627_,
    new_n15628_, new_n15629_, new_n15630_, new_n15631_, new_n15632_,
    new_n15633_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15640_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15651_, new_n15652_,
    new_n15653_, new_n15654_, new_n15655_, new_n15656_, new_n15657_,
    new_n15658_, new_n15659_, new_n15660_, new_n15661_, new_n15662_,
    new_n15663_, new_n15664_, new_n15665_, new_n15666_, new_n15667_,
    new_n15668_, new_n15669_, new_n15670_, new_n15671_, new_n15672_,
    new_n15673_, new_n15674_, new_n15675_, new_n15676_, new_n15677_,
    new_n15678_, new_n15679_, new_n15680_, new_n15681_, new_n15682_,
    new_n15683_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15697_,
    new_n15698_, new_n15699_, new_n15700_, new_n15701_, new_n15702_,
    new_n15703_, new_n15704_, new_n15705_, new_n15706_, new_n15707_,
    new_n15708_, new_n15709_, new_n15710_, new_n15712_, new_n15713_,
    new_n15714_, new_n15715_, new_n15716_, new_n15717_, new_n15718_,
    new_n15719_, new_n15720_, new_n15721_, new_n15722_, new_n15723_,
    new_n15724_, new_n15725_, new_n15726_, new_n15727_, new_n15728_,
    new_n15729_, new_n15730_, new_n15731_, new_n15732_, new_n15733_,
    new_n15734_, new_n15735_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15889_, new_n15890_, new_n15891_,
    new_n15892_, new_n15893_, new_n15894_, new_n15895_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15925_, new_n15926_,
    new_n15927_, new_n15928_, new_n15929_, new_n15930_, new_n15931_,
    new_n15932_, new_n15933_, new_n15934_, new_n15935_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16011_,
    new_n16012_, new_n16013_, new_n16014_, new_n16015_, new_n16016_,
    new_n16017_, new_n16018_, new_n16019_, new_n16020_, new_n16021_,
    new_n16022_, new_n16023_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16040_, new_n16041_,
    new_n16042_, new_n16043_, new_n16044_, new_n16045_, new_n16046_,
    new_n16047_, new_n16048_, new_n16049_, new_n16050_, new_n16051_,
    new_n16052_, new_n16053_, new_n16054_, new_n16055_, new_n16056_,
    new_n16057_, new_n16058_, new_n16059_, new_n16060_, new_n16061_,
    new_n16062_, new_n16063_, new_n16064_, new_n16065_, new_n16066_,
    new_n16067_, new_n16068_, new_n16069_, new_n16070_, new_n16071_,
    new_n16072_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16082_, new_n16083_, new_n16084_, new_n16085_, new_n16086_,
    new_n16087_, new_n16088_, new_n16089_, new_n16090_, new_n16091_,
    new_n16092_, new_n16093_, new_n16094_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16100_, new_n16101_, new_n16102_,
    new_n16103_, new_n16104_, new_n16105_, new_n16106_, new_n16107_,
    new_n16108_, new_n16109_, new_n16110_, new_n16111_, new_n16112_,
    new_n16113_, new_n16114_, new_n16115_, new_n16116_, new_n16117_,
    new_n16118_, new_n16119_, new_n16120_, new_n16121_, new_n16122_,
    new_n16123_, new_n16124_, new_n16125_, new_n16126_, new_n16127_,
    new_n16128_, new_n16129_, new_n16130_, new_n16131_, new_n16132_,
    new_n16133_, new_n16134_, new_n16135_, new_n16136_, new_n16137_,
    new_n16138_, new_n16139_, new_n16140_, new_n16141_, new_n16142_,
    new_n16143_, new_n16144_, new_n16145_, new_n16146_, new_n16147_,
    new_n16148_, new_n16149_, new_n16150_, new_n16151_, new_n16152_,
    new_n16153_, new_n16154_, new_n16155_, new_n16157_, new_n16158_,
    new_n16159_, new_n16160_, new_n16161_, new_n16162_, new_n16163_,
    new_n16164_, new_n16165_, new_n16166_, new_n16167_, new_n16168_,
    new_n16169_, new_n16170_, new_n16171_, new_n16172_, new_n16173_,
    new_n16174_, new_n16175_, new_n16176_, new_n16177_, new_n16178_,
    new_n16179_, new_n16180_, new_n16181_, new_n16182_, new_n16183_,
    new_n16184_, new_n16185_, new_n16186_, new_n16187_, new_n16188_,
    new_n16189_, new_n16190_, new_n16191_, new_n16192_, new_n16193_,
    new_n16194_, new_n16195_, new_n16196_, new_n16197_, new_n16198_,
    new_n16199_, new_n16200_, new_n16201_, new_n16202_, new_n16203_,
    new_n16204_, new_n16205_, new_n16206_, new_n16207_, new_n16208_,
    new_n16209_, new_n16210_, new_n16211_, new_n16212_, new_n16213_,
    new_n16214_, new_n16215_, new_n16216_, new_n16217_, new_n16218_,
    new_n16219_, new_n16220_, new_n16221_, new_n16222_, new_n16223_,
    new_n16224_, new_n16225_, new_n16226_, new_n16227_, new_n16228_,
    new_n16229_, new_n16230_, new_n16231_, new_n16232_, new_n16233_,
    new_n16234_, new_n16235_, new_n16236_, new_n16237_, new_n16238_,
    new_n16239_, new_n16240_, new_n16241_, new_n16242_, new_n16243_,
    new_n16244_, new_n16245_, new_n16246_, new_n16247_, new_n16248_,
    new_n16249_, new_n16250_, new_n16251_, new_n16252_, new_n16253_,
    new_n16254_, new_n16255_, new_n16256_, new_n16257_, new_n16258_,
    new_n16259_, new_n16260_, new_n16261_, new_n16262_, new_n16263_,
    new_n16264_, new_n16265_, new_n16266_, new_n16267_, new_n16268_,
    new_n16269_, new_n16271_, new_n16272_, new_n16273_, new_n16274_,
    new_n16275_, new_n16276_, new_n16277_, new_n16278_, new_n16279_,
    new_n16280_, new_n16281_, new_n16282_, new_n16283_, new_n16284_,
    new_n16285_, new_n16286_, new_n16287_, new_n16288_, new_n16289_,
    new_n16290_, new_n16291_, new_n16292_, new_n16293_, new_n16294_,
    new_n16295_, new_n16296_, new_n16297_, new_n16298_, new_n16299_,
    new_n16300_, new_n16301_, new_n16302_, new_n16303_, new_n16304_,
    new_n16305_, new_n16306_, new_n16307_, new_n16308_, new_n16309_,
    new_n16310_, new_n16311_, new_n16312_, new_n16313_, new_n16314_,
    new_n16315_, new_n16316_, new_n16317_, new_n16318_, new_n16319_,
    new_n16320_, new_n16321_, new_n16322_, new_n16323_, new_n16324_,
    new_n16325_, new_n16326_, new_n16327_, new_n16328_, new_n16329_,
    new_n16330_, new_n16331_, new_n16332_, new_n16333_, new_n16334_,
    new_n16335_, new_n16336_, new_n16337_, new_n16338_, new_n16339_,
    new_n16340_, new_n16341_, new_n16342_, new_n16343_, new_n16344_,
    new_n16345_, new_n16346_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16353_, new_n16354_,
    new_n16355_, new_n16356_, new_n16357_, new_n16358_, new_n16359_,
    new_n16360_, new_n16361_, new_n16362_, new_n16363_, new_n16364_,
    new_n16365_, new_n16366_, new_n16367_, new_n16368_, new_n16369_,
    new_n16370_, new_n16371_, new_n16372_, new_n16373_, new_n16374_,
    new_n16375_, new_n16376_, new_n16377_, new_n16378_, new_n16379_,
    new_n16380_, new_n16381_, new_n16382_, new_n16383_, new_n16384_,
    new_n16385_, new_n16386_, new_n16387_, new_n16388_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16489_, new_n16490_, new_n16491_, new_n16492_,
    new_n16493_, new_n16494_, new_n16495_, new_n16496_, new_n16497_,
    new_n16498_, new_n16499_, new_n16500_, new_n16501_, new_n16502_,
    new_n16503_, new_n16504_, new_n16505_, new_n16506_, new_n16507_,
    new_n16508_, new_n16509_, new_n16510_, new_n16511_, new_n16512_,
    new_n16513_, new_n16514_, new_n16515_, new_n16516_, new_n16517_,
    new_n16518_, new_n16519_, new_n16520_, new_n16521_, new_n16522_,
    new_n16523_, new_n16524_, new_n16525_, new_n16526_, new_n16527_,
    new_n16528_, new_n16529_, new_n16530_, new_n16531_, new_n16532_,
    new_n16533_, new_n16534_, new_n16535_, new_n16536_, new_n16537_,
    new_n16538_, new_n16539_, new_n16540_, new_n16541_, new_n16542_,
    new_n16543_, new_n16544_, new_n16545_, new_n16546_, new_n16547_,
    new_n16548_, new_n16549_, new_n16550_, new_n16551_, new_n16552_,
    new_n16553_, new_n16554_, new_n16555_, new_n16556_, new_n16557_,
    new_n16558_, new_n16559_, new_n16560_, new_n16561_, new_n16562_,
    new_n16563_, new_n16564_, new_n16565_, new_n16566_, new_n16567_,
    new_n16568_, new_n16569_, new_n16570_, new_n16571_, new_n16572_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16590_, new_n16591_, new_n16592_, new_n16593_,
    new_n16594_, new_n16595_, new_n16596_, new_n16597_, new_n16598_,
    new_n16599_, new_n16600_, new_n16601_, new_n16602_, new_n16603_,
    new_n16604_, new_n16605_, new_n16606_, new_n16607_, new_n16608_,
    new_n16609_, new_n16610_, new_n16611_, new_n16612_, new_n16613_,
    new_n16614_, new_n16615_, new_n16616_, new_n16617_, new_n16618_,
    new_n16619_, new_n16620_, new_n16621_, new_n16622_, new_n16623_,
    new_n16624_, new_n16625_, new_n16626_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16862_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16868_, new_n16869_,
    new_n16870_, new_n16871_, new_n16872_, new_n16873_, new_n16874_,
    new_n16875_, new_n16876_, new_n16877_, new_n16878_, new_n16879_,
    new_n16880_, new_n16881_, new_n16882_, new_n16883_, new_n16884_,
    new_n16885_, new_n16886_, new_n16887_, new_n16888_, new_n16889_,
    new_n16890_, new_n16891_, new_n16892_, new_n16893_, new_n16894_,
    new_n16895_, new_n16896_, new_n16897_, new_n16898_, new_n16899_,
    new_n16900_, new_n16901_, new_n16902_, new_n16903_, new_n16904_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16953_, new_n16954_,
    new_n16955_, new_n16956_, new_n16957_, new_n16958_, new_n16959_,
    new_n16960_, new_n16961_, new_n16962_, new_n16963_, new_n16964_,
    new_n16965_, new_n16966_, new_n16967_, new_n16968_, new_n16969_,
    new_n16970_, new_n16971_, new_n16972_, new_n16973_, new_n16974_,
    new_n16975_, new_n16976_, new_n16977_, new_n16978_, new_n16979_,
    new_n16980_, new_n16981_, new_n16982_, new_n16983_, new_n16984_,
    new_n16985_, new_n16986_, new_n16987_, new_n16988_, new_n16989_,
    new_n16990_, new_n16991_, new_n16992_, new_n16993_, new_n16994_,
    new_n16995_, new_n16996_, new_n16997_, new_n16998_, new_n16999_,
    new_n17000_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17005_, new_n17006_, new_n17007_, new_n17008_, new_n17009_,
    new_n17010_, new_n17011_, new_n17012_, new_n17013_, new_n17014_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17024_,
    new_n17025_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17030_, new_n17031_, new_n17032_, new_n17033_, new_n17034_,
    new_n17035_, new_n17036_, new_n17037_, new_n17038_, new_n17039_,
    new_n17040_, new_n17041_, new_n17042_, new_n17043_, new_n17044_,
    new_n17045_, new_n17046_, new_n17047_, new_n17048_, new_n17049_,
    new_n17050_, new_n17051_, new_n17052_, new_n17053_, new_n17054_,
    new_n17055_, new_n17056_, new_n17057_, new_n17058_, new_n17059_,
    new_n17060_, new_n17061_, new_n17062_, new_n17063_, new_n17064_,
    new_n17065_, new_n17066_, new_n17067_, new_n17068_, new_n17069_,
    new_n17070_, new_n17071_, new_n17072_, new_n17073_, new_n17074_,
    new_n17075_, new_n17076_, new_n17077_, new_n17078_, new_n17079_,
    new_n17080_, new_n17081_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17113_, new_n17114_,
    new_n17115_, new_n17116_, new_n17117_, new_n17118_, new_n17119_,
    new_n17120_, new_n17121_, new_n17122_, new_n17123_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17130_,
    new_n17131_, new_n17132_, new_n17133_, new_n17134_, new_n17135_,
    new_n17136_, new_n17137_, new_n17138_, new_n17139_, new_n17140_,
    new_n17141_, new_n17142_, new_n17143_, new_n17144_, new_n17145_,
    new_n17146_, new_n17147_, new_n17148_, new_n17149_, new_n17150_,
    new_n17151_, new_n17152_, new_n17153_, new_n17154_, new_n17155_,
    new_n17156_, new_n17157_, new_n17158_, new_n17159_, new_n17160_,
    new_n17161_, new_n17162_, new_n17163_, new_n17164_, new_n17165_,
    new_n17166_, new_n17167_, new_n17168_, new_n17169_, new_n17170_,
    new_n17171_, new_n17172_, new_n17173_, new_n17174_, new_n17175_,
    new_n17176_, new_n17177_, new_n17178_, new_n17179_, new_n17180_,
    new_n17181_, new_n17182_, new_n17183_, new_n17184_, new_n17185_,
    new_n17186_, new_n17187_, new_n17188_, new_n17189_, new_n17190_,
    new_n17191_, new_n17192_, new_n17193_, new_n17194_, new_n17195_,
    new_n17196_, new_n17197_, new_n17198_, new_n17199_, new_n17200_,
    new_n17201_, new_n17202_, new_n17203_, new_n17204_, new_n17205_,
    new_n17206_, new_n17207_, new_n17208_, new_n17209_, new_n17210_,
    new_n17211_, new_n17212_, new_n17213_, new_n17214_, new_n17215_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17380_,
    new_n17381_, new_n17382_, new_n17383_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17389_, new_n17390_,
    new_n17391_, new_n17392_, new_n17393_, new_n17394_, new_n17395_,
    new_n17396_, new_n17397_, new_n17398_, new_n17399_, new_n17400_,
    new_n17401_, new_n17402_, new_n17403_, new_n17404_, new_n17405_,
    new_n17406_, new_n17407_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17498_, new_n17499_, new_n17500_,
    new_n17501_, new_n17502_, new_n17503_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17510_,
    new_n17511_, new_n17512_, new_n17513_, new_n17514_, new_n17515_,
    new_n17516_, new_n17517_, new_n17518_, new_n17519_, new_n17520_,
    new_n17521_, new_n17522_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17558_, new_n17559_, new_n17560_,
    new_n17561_, new_n17562_, new_n17563_, new_n17564_, new_n17565_,
    new_n17566_, new_n17567_, new_n17568_, new_n17569_, new_n17570_,
    new_n17571_, new_n17572_, new_n17573_, new_n17574_, new_n17575_,
    new_n17576_, new_n17577_, new_n17578_, new_n17579_, new_n17580_,
    new_n17581_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17586_, new_n17587_, new_n17588_, new_n17589_, new_n17590_,
    new_n17591_, new_n17592_, new_n17593_, new_n17594_, new_n17595_,
    new_n17596_, new_n17597_, new_n17598_, new_n17599_, new_n17600_,
    new_n17601_, new_n17602_, new_n17603_, new_n17604_, new_n17605_,
    new_n17606_, new_n17607_, new_n17608_, new_n17609_, new_n17610_,
    new_n17611_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17669_, new_n17670_,
    new_n17671_, new_n17672_, new_n17673_, new_n17674_, new_n17675_,
    new_n17676_, new_n17677_, new_n17678_, new_n17679_, new_n17680_,
    new_n17681_, new_n17682_, new_n17683_, new_n17684_, new_n17685_,
    new_n17686_, new_n17687_, new_n17688_, new_n17689_, new_n17690_,
    new_n17691_, new_n17692_, new_n17693_, new_n17694_, new_n17695_,
    new_n17696_, new_n17697_, new_n17698_, new_n17699_, new_n17700_,
    new_n17701_, new_n17702_, new_n17703_, new_n17704_, new_n17705_,
    new_n17706_, new_n17707_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17747_, new_n17748_, new_n17749_, new_n17750_,
    new_n17751_, new_n17752_, new_n17753_, new_n17754_, new_n17755_,
    new_n17756_, new_n17757_, new_n17758_, new_n17759_, new_n17760_,
    new_n17761_, new_n17762_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17791_, new_n17792_, new_n17793_, new_n17794_, new_n17795_,
    new_n17796_, new_n17797_, new_n17798_, new_n17799_, new_n17800_,
    new_n17801_, new_n17802_, new_n17803_, new_n17804_, new_n17805_,
    new_n17806_, new_n17807_, new_n17808_, new_n17809_, new_n17810_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17832_, new_n17833_, new_n17834_, new_n17835_,
    new_n17836_, new_n17837_, new_n17838_, new_n17839_, new_n17840_,
    new_n17841_, new_n17842_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17887_, new_n17888_, new_n17889_, new_n17890_,
    new_n17891_, new_n17892_, new_n17893_, new_n17894_, new_n17895_,
    new_n17896_, new_n17897_, new_n17898_, new_n17899_, new_n17900_,
    new_n17901_, new_n17902_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17973_, new_n17974_, new_n17975_,
    new_n17976_, new_n17977_, new_n17978_, new_n17979_, new_n17980_,
    new_n17981_, new_n17982_, new_n17983_, new_n17984_, new_n17985_,
    new_n17986_, new_n17987_, new_n17988_, new_n17989_, new_n17990_,
    new_n17991_, new_n17992_, new_n17993_, new_n17994_, new_n17995_,
    new_n17996_, new_n17997_, new_n17998_, new_n17999_, new_n18000_,
    new_n18001_, new_n18002_, new_n18003_, new_n18004_, new_n18005_,
    new_n18006_, new_n18007_, new_n18008_, new_n18009_, new_n18010_,
    new_n18011_, new_n18012_, new_n18013_, new_n18014_, new_n18015_,
    new_n18016_, new_n18017_, new_n18018_, new_n18019_, new_n18020_,
    new_n18021_, new_n18022_, new_n18023_, new_n18024_, new_n18025_,
    new_n18026_, new_n18027_, new_n18028_, new_n18029_, new_n18030_,
    new_n18031_, new_n18032_, new_n18033_, new_n18034_, new_n18035_,
    new_n18036_, new_n18037_, new_n18038_, new_n18039_, new_n18040_,
    new_n18041_, new_n18042_, new_n18043_, new_n18044_, new_n18045_,
    new_n18046_, new_n18047_, new_n18048_, new_n18049_, new_n18050_,
    new_n18051_, new_n18052_, new_n18053_, new_n18054_, new_n18055_,
    new_n18056_, new_n18057_, new_n18058_, new_n18059_, new_n18060_,
    new_n18061_, new_n18062_, new_n18063_, new_n18064_, new_n18066_,
    new_n18067_, new_n18068_, new_n18069_, new_n18070_, new_n18071_,
    new_n18072_, new_n18073_, new_n18074_, new_n18075_, new_n18076_,
    new_n18077_, new_n18078_, new_n18079_, new_n18080_, new_n18081_,
    new_n18082_, new_n18083_, new_n18084_, new_n18085_, new_n18086_,
    new_n18087_, new_n18088_, new_n18089_, new_n18090_, new_n18091_,
    new_n18092_, new_n18093_, new_n18094_, new_n18095_, new_n18096_,
    new_n18097_, new_n18098_, new_n18099_, new_n18100_, new_n18101_,
    new_n18102_, new_n18103_, new_n18104_, new_n18105_, new_n18106_,
    new_n18107_, new_n18108_, new_n18109_, new_n18110_, new_n18111_,
    new_n18112_, new_n18113_, new_n18114_, new_n18115_, new_n18116_,
    new_n18117_, new_n18118_, new_n18119_, new_n18120_, new_n18121_,
    new_n18122_, new_n18123_, new_n18124_, new_n18125_, new_n18126_,
    new_n18127_, new_n18128_, new_n18129_, new_n18130_, new_n18131_,
    new_n18132_, new_n18133_, new_n18134_, new_n18135_, new_n18136_,
    new_n18137_, new_n18138_, new_n18139_, new_n18140_, new_n18141_,
    new_n18142_, new_n18143_, new_n18144_, new_n18145_, new_n18146_,
    new_n18147_, new_n18148_, new_n18149_, new_n18150_, new_n18151_,
    new_n18152_, new_n18153_, new_n18154_, new_n18155_, new_n18156_,
    new_n18157_, new_n18158_, new_n18159_, new_n18160_, new_n18161_,
    new_n18162_, new_n18163_, new_n18164_, new_n18165_, new_n18166_,
    new_n18167_, new_n18168_, new_n18169_, new_n18170_, new_n18171_,
    new_n18172_, new_n18173_, new_n18174_, new_n18175_, new_n18176_,
    new_n18177_, new_n18178_, new_n18179_, new_n18180_, new_n18181_,
    new_n18182_, new_n18183_, new_n18184_, new_n18185_, new_n18186_,
    new_n18187_, new_n18188_, new_n18189_, new_n18190_, new_n18191_,
    new_n18192_, new_n18193_, new_n18194_, new_n18195_, new_n18196_,
    new_n18197_, new_n18198_, new_n18199_, new_n18200_, new_n18201_,
    new_n18202_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18210_, new_n18211_,
    new_n18212_, new_n18213_, new_n18214_, new_n18215_, new_n18216_,
    new_n18217_, new_n18218_, new_n18219_, new_n18220_, new_n18221_,
    new_n18222_, new_n18223_, new_n18224_, new_n18225_, new_n18226_,
    new_n18227_, new_n18228_, new_n18229_, new_n18230_, new_n18231_,
    new_n18232_, new_n18233_, new_n18234_, new_n18235_, new_n18236_,
    new_n18237_, new_n18238_, new_n18239_, new_n18240_, new_n18241_,
    new_n18242_, new_n18243_, new_n18244_, new_n18245_, new_n18246_,
    new_n18247_, new_n18248_, new_n18249_, new_n18250_, new_n18251_,
    new_n18252_, new_n18253_, new_n18254_, new_n18255_, new_n18256_,
    new_n18257_, new_n18258_, new_n18259_, new_n18260_, new_n18261_,
    new_n18262_, new_n18263_, new_n18264_, new_n18265_, new_n18266_,
    new_n18267_, new_n18268_, new_n18269_, new_n18270_, new_n18271_,
    new_n18272_, new_n18273_, new_n18274_, new_n18275_, new_n18276_,
    new_n18277_, new_n18278_, new_n18279_, new_n18280_, new_n18281_,
    new_n18282_, new_n18283_, new_n18284_, new_n18285_, new_n18286_,
    new_n18287_, new_n18288_, new_n18289_, new_n18290_, new_n18291_,
    new_n18292_, new_n18293_, new_n18294_, new_n18295_, new_n18296_,
    new_n18297_, new_n18298_, new_n18299_, new_n18300_, new_n18301_,
    new_n18302_, new_n18303_, new_n18304_, new_n18305_, new_n18306_,
    new_n18307_, new_n18308_, new_n18309_, new_n18310_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18315_, new_n18316_,
    new_n18317_, new_n18318_, new_n18319_, new_n18320_, new_n18321_,
    new_n18322_, new_n18323_, new_n18324_, new_n18325_, new_n18326_,
    new_n18327_, new_n18328_, new_n18329_, new_n18330_, new_n18331_,
    new_n18332_, new_n18333_, new_n18334_, new_n18335_, new_n18336_,
    new_n18337_, new_n18338_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18577_, new_n18578_, new_n18579_, new_n18580_, new_n18581_,
    new_n18582_, new_n18583_, new_n18584_, new_n18585_, new_n18586_,
    new_n18587_, new_n18588_, new_n18589_, new_n18591_, new_n18592_,
    new_n18593_, new_n18594_, new_n18595_, new_n18596_, new_n18597_,
    new_n18598_, new_n18599_, new_n18600_, new_n18601_, new_n18602_,
    new_n18603_, new_n18604_, new_n18605_, new_n18606_, new_n18607_,
    new_n18608_, new_n18609_, new_n18610_, new_n18611_, new_n18612_,
    new_n18613_, new_n18614_, new_n18615_, new_n18616_, new_n18617_,
    new_n18618_, new_n18619_, new_n18620_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18625_, new_n18626_, new_n18627_,
    new_n18628_, new_n18629_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18717_,
    new_n18718_, new_n18719_, new_n18720_, new_n18721_, new_n18722_,
    new_n18723_, new_n18724_, new_n18725_, new_n18726_, new_n18727_,
    new_n18728_, new_n18729_, new_n18730_, new_n18731_, new_n18732_,
    new_n18733_, new_n18734_, new_n18735_, new_n18736_, new_n18737_,
    new_n18738_, new_n18739_, new_n18740_, new_n18741_, new_n18742_,
    new_n18743_, new_n18744_, new_n18745_, new_n18746_, new_n18747_,
    new_n18748_, new_n18749_, new_n18750_, new_n18751_, new_n18752_,
    new_n18753_, new_n18754_, new_n18755_, new_n18756_, new_n18757_,
    new_n18758_, new_n18759_, new_n18760_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18765_, new_n18766_, new_n18767_,
    new_n18768_, new_n18769_, new_n18770_, new_n18771_, new_n18772_,
    new_n18773_, new_n18774_, new_n18775_, new_n18776_, new_n18777_,
    new_n18778_, new_n18779_, new_n18780_, new_n18781_, new_n18782_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18788_, new_n18789_, new_n18790_, new_n18791_, new_n18792_,
    new_n18793_, new_n18794_, new_n18795_, new_n18796_, new_n18797_,
    new_n18798_, new_n18799_, new_n18800_, new_n18801_, new_n18802_,
    new_n18803_, new_n18804_, new_n18805_, new_n18806_, new_n18807_,
    new_n18808_, new_n18809_, new_n18810_, new_n18811_, new_n18812_,
    new_n18813_, new_n18814_, new_n18815_, new_n18816_, new_n18817_,
    new_n18818_, new_n18819_, new_n18820_, new_n18821_, new_n18822_,
    new_n18823_, new_n18824_, new_n18825_, new_n18826_, new_n18827_,
    new_n18828_, new_n18829_, new_n18830_, new_n18831_, new_n18832_,
    new_n18833_, new_n18834_, new_n18835_, new_n18836_, new_n18837_,
    new_n18838_, new_n18839_, new_n18840_, new_n18841_, new_n18842_,
    new_n18843_, new_n18844_, new_n18845_, new_n18846_, new_n18847_,
    new_n18848_, new_n18849_, new_n18850_, new_n18851_, new_n18852_,
    new_n18853_, new_n18854_, new_n18855_, new_n18856_, new_n18857_,
    new_n18858_, new_n18859_, new_n18860_, new_n18861_, new_n18862_,
    new_n18863_, new_n18864_, new_n18865_, new_n18866_, new_n18867_,
    new_n18868_, new_n18869_, new_n18870_, new_n18871_, new_n18872_,
    new_n18873_, new_n18874_, new_n18875_, new_n18876_, new_n18877_,
    new_n18878_, new_n18879_, new_n18880_, new_n18881_, new_n18882_,
    new_n18883_, new_n18884_, new_n18885_, new_n18886_, new_n18887_,
    new_n18888_, new_n18889_, new_n18890_, new_n18891_, new_n18892_,
    new_n18893_, new_n18894_, new_n18895_, new_n18896_, new_n18897_,
    new_n18898_, new_n18899_, new_n18900_, new_n18901_, new_n18902_,
    new_n18903_, new_n18904_, new_n18905_, new_n18906_, new_n18907_,
    new_n18908_, new_n18909_, new_n18910_, new_n18911_, new_n18912_,
    new_n18913_, new_n18914_, new_n18915_, new_n18916_, new_n18917_,
    new_n18918_, new_n18919_, new_n18920_, new_n18921_, new_n18922_,
    new_n18923_, new_n18924_, new_n18925_, new_n18926_, new_n18927_,
    new_n18928_, new_n18929_, new_n18930_, new_n18931_, new_n18932_,
    new_n18933_, new_n18934_, new_n18935_, new_n18936_, new_n18937_,
    new_n18938_, new_n18939_, new_n18940_, new_n18941_, new_n18942_,
    new_n18943_, new_n18944_, new_n18945_, new_n18946_, new_n18947_,
    new_n18948_, new_n18949_, new_n18950_, new_n18951_, new_n18952_,
    new_n18953_, new_n18954_, new_n18955_, new_n18956_, new_n18957_,
    new_n18958_, new_n18959_, new_n18960_, new_n18961_, new_n18962_,
    new_n18963_, new_n18964_, new_n18965_, new_n18966_, new_n18967_,
    new_n18968_, new_n18969_, new_n18970_, new_n18971_, new_n18972_,
    new_n18973_, new_n18974_, new_n18975_, new_n18976_, new_n18977_,
    new_n18978_, new_n18979_, new_n18980_, new_n18981_, new_n18982_,
    new_n18983_, new_n18984_, new_n18985_, new_n18986_, new_n18987_,
    new_n18988_, new_n18989_, new_n18990_, new_n18991_, new_n18992_,
    new_n18993_, new_n18994_, new_n18995_, new_n18996_, new_n18997_,
    new_n18998_, new_n18999_, new_n19000_, new_n19001_, new_n19002_,
    new_n19003_, new_n19004_, new_n19005_, new_n19006_, new_n19007_,
    new_n19008_, new_n19009_, new_n19010_, new_n19011_, new_n19012_,
    new_n19013_, new_n19014_, new_n19015_, new_n19016_, new_n19017_,
    new_n19018_, new_n19019_, new_n19020_, new_n19021_, new_n19022_,
    new_n19023_, new_n19024_, new_n19025_, new_n19026_, new_n19027_,
    new_n19028_, new_n19029_, new_n19030_, new_n19031_, new_n19032_,
    new_n19033_, new_n19034_, new_n19035_, new_n19036_, new_n19037_,
    new_n19038_, new_n19039_, new_n19040_, new_n19041_, new_n19042_,
    new_n19043_, new_n19044_, new_n19045_, new_n19046_, new_n19047_,
    new_n19048_, new_n19049_, new_n19050_, new_n19051_, new_n19052_,
    new_n19053_, new_n19054_, new_n19055_, new_n19056_, new_n19057_,
    new_n19058_, new_n19059_, new_n19060_, new_n19061_, new_n19062_,
    new_n19063_, new_n19064_, new_n19065_, new_n19066_, new_n19067_,
    new_n19068_, new_n19069_, new_n19070_, new_n19071_, new_n19072_,
    new_n19073_, new_n19074_, new_n19075_, new_n19076_, new_n19077_,
    new_n19078_, new_n19079_, new_n19080_, new_n19081_, new_n19082_,
    new_n19083_, new_n19084_, new_n19085_, new_n19086_, new_n19087_,
    new_n19088_, new_n19089_, new_n19090_, new_n19091_, new_n19092_,
    new_n19093_, new_n19094_, new_n19095_, new_n19096_, new_n19097_,
    new_n19098_, new_n19099_, new_n19100_, new_n19101_, new_n19102_,
    new_n19103_, new_n19104_, new_n19105_, new_n19106_, new_n19107_,
    new_n19108_, new_n19109_, new_n19110_, new_n19111_, new_n19112_,
    new_n19113_, new_n19114_, new_n19115_, new_n19116_, new_n19117_,
    new_n19118_, new_n19119_, new_n19120_, new_n19121_, new_n19122_,
    new_n19123_, new_n19124_, new_n19125_, new_n19126_, new_n19127_,
    new_n19128_, new_n19129_, new_n19130_, new_n19131_, new_n19132_,
    new_n19133_, new_n19134_, new_n19135_, new_n19136_, new_n19137_,
    new_n19138_, new_n19139_, new_n19140_, new_n19141_, new_n19142_,
    new_n19143_, new_n19144_, new_n19145_, new_n19146_, new_n19147_,
    new_n19148_, new_n19149_, new_n19150_, new_n19151_, new_n19152_,
    new_n19153_, new_n19154_, new_n19155_, new_n19156_, new_n19157_,
    new_n19158_, new_n19159_, new_n19160_, new_n19161_, new_n19162_,
    new_n19163_, new_n19164_, new_n19165_, new_n19166_, new_n19167_,
    new_n19168_, new_n19169_, new_n19170_, new_n19171_, new_n19172_,
    new_n19173_, new_n19174_, new_n19175_, new_n19176_, new_n19177_,
    new_n19178_, new_n19179_, new_n19180_, new_n19181_, new_n19182_,
    new_n19183_, new_n19184_, new_n19185_, new_n19186_, new_n19187_,
    new_n19188_, new_n19189_, new_n19190_, new_n19191_, new_n19192_,
    new_n19193_, new_n19194_, new_n19195_, new_n19196_, new_n19197_,
    new_n19198_, new_n19199_, new_n19200_, new_n19201_, new_n19202_,
    new_n19203_, new_n19204_, new_n19205_, new_n19206_, new_n19207_,
    new_n19208_, new_n19209_, new_n19210_, new_n19211_, new_n19212_,
    new_n19213_, new_n19214_, new_n19215_, new_n19216_, new_n19217_,
    new_n19218_, new_n19219_, new_n19220_, new_n19221_, new_n19222_,
    new_n19223_, new_n19224_, new_n19225_, new_n19226_, new_n19227_,
    new_n19228_, new_n19229_, new_n19230_, new_n19231_, new_n19232_,
    new_n19233_, new_n19234_, new_n19235_, new_n19236_, new_n19237_,
    new_n19238_, new_n19239_, new_n19240_, new_n19241_, new_n19242_,
    new_n19243_, new_n19244_, new_n19245_, new_n19246_, new_n19247_,
    new_n19248_, new_n19249_, new_n19250_, new_n19251_, new_n19252_,
    new_n19253_, new_n19254_, new_n19255_, new_n19256_, new_n19257_,
    new_n19258_, new_n19259_, new_n19260_, new_n19261_, new_n19262_,
    new_n19263_, new_n19264_, new_n19265_, new_n19266_, new_n19267_,
    new_n19268_, new_n19269_, new_n19270_, new_n19271_, new_n19272_,
    new_n19273_, new_n19274_, new_n19275_, new_n19276_, new_n19277_,
    new_n19278_, new_n19279_, new_n19280_, new_n19281_, new_n19282_,
    new_n19283_, new_n19284_, new_n19285_, new_n19286_, new_n19287_,
    new_n19288_, new_n19289_, new_n19290_, new_n19291_, new_n19292_,
    new_n19293_, new_n19294_, new_n19295_, new_n19296_, new_n19297_,
    new_n19298_, new_n19299_, new_n19300_, new_n19301_, new_n19302_,
    new_n19303_, new_n19304_, new_n19305_, new_n19306_, new_n19307_,
    new_n19308_, new_n19309_, new_n19310_, new_n19311_, new_n19312_,
    new_n19313_, new_n19314_, new_n19315_, new_n19316_, new_n19317_,
    new_n19318_, new_n19319_, new_n19320_, new_n19321_, new_n19322_,
    new_n19323_, new_n19324_, new_n19325_, new_n19326_, new_n19327_,
    new_n19328_, new_n19329_, new_n19330_, new_n19331_, new_n19332_,
    new_n19333_, new_n19334_, new_n19335_, new_n19336_, new_n19337_,
    new_n19338_, new_n19339_, new_n19340_, new_n19341_, new_n19342_,
    new_n19343_, new_n19344_, new_n19345_, new_n19346_, new_n19347_,
    new_n19348_, new_n19349_, new_n19350_, new_n19351_, new_n19352_,
    new_n19353_, new_n19354_, new_n19355_, new_n19356_, new_n19357_,
    new_n19358_, new_n19359_, new_n19360_, new_n19361_, new_n19362_,
    new_n19363_, new_n19364_, new_n19366_, new_n19367_, new_n19368_,
    new_n19369_, new_n19370_, new_n19371_, new_n19372_, new_n19373_,
    new_n19374_, new_n19375_, new_n19376_, new_n19377_, new_n19378_,
    new_n19379_, new_n19380_, new_n19381_, new_n19382_, new_n19383_,
    new_n19384_, new_n19385_, new_n19386_, new_n19387_, new_n19388_,
    new_n19389_, new_n19390_, new_n19391_, new_n19392_, new_n19393_,
    new_n19394_, new_n19395_, new_n19396_, new_n19397_, new_n19398_,
    new_n19399_, new_n19400_, new_n19401_, new_n19402_, new_n19403_,
    new_n19404_, new_n19405_, new_n19406_, new_n19407_, new_n19408_,
    new_n19409_, new_n19410_, new_n19411_, new_n19412_, new_n19413_,
    new_n19414_, new_n19415_, new_n19416_, new_n19417_, new_n19418_,
    new_n19419_, new_n19420_, new_n19421_, new_n19422_, new_n19423_,
    new_n19424_, new_n19425_, new_n19426_, new_n19427_, new_n19428_,
    new_n19429_, new_n19430_, new_n19431_, new_n19432_, new_n19433_,
    new_n19434_, new_n19435_, new_n19436_, new_n19437_, new_n19438_,
    new_n19439_, new_n19440_, new_n19441_, new_n19442_, new_n19443_,
    new_n19444_, new_n19445_, new_n19446_, new_n19447_, new_n19448_,
    new_n19449_, new_n19450_, new_n19451_, new_n19452_, new_n19453_,
    new_n19454_, new_n19455_, new_n19456_, new_n19457_, new_n19458_,
    new_n19459_, new_n19460_, new_n19461_, new_n19462_, new_n19463_,
    new_n19464_, new_n19465_, new_n19466_, new_n19467_, new_n19468_,
    new_n19469_, new_n19470_, new_n19471_, new_n19472_, new_n19473_,
    new_n19474_, new_n19475_, new_n19476_, new_n19477_, new_n19478_,
    new_n19479_, new_n19480_, new_n19481_, new_n19482_, new_n19483_,
    new_n19484_, new_n19485_, new_n19486_, new_n19487_, new_n19488_,
    new_n19489_, new_n19490_, new_n19491_, new_n19492_, new_n19493_,
    new_n19494_, new_n19495_, new_n19496_, new_n19497_, new_n19498_,
    new_n19499_, new_n19500_, new_n19501_, new_n19502_, new_n19503_,
    new_n19504_, new_n19505_, new_n19506_, new_n19507_, new_n19508_,
    new_n19509_, new_n19510_, new_n19511_, new_n19512_, new_n19513_,
    new_n19514_, new_n19515_, new_n19516_, new_n19517_, new_n19518_,
    new_n19519_, new_n19520_, new_n19521_, new_n19522_, new_n19523_,
    new_n19524_, new_n19525_, new_n19526_, new_n19527_, new_n19528_,
    new_n19529_, new_n19530_, new_n19531_, new_n19532_, new_n19533_,
    new_n19534_, new_n19535_, new_n19536_, new_n19537_, new_n19538_,
    new_n19539_, new_n19540_, new_n19541_, new_n19542_, new_n19543_,
    new_n19544_, new_n19545_, new_n19546_, new_n19547_, new_n19548_,
    new_n19549_, new_n19550_, new_n19551_, new_n19552_, new_n19553_,
    new_n19554_, new_n19555_, new_n19556_, new_n19557_, new_n19558_,
    new_n19559_, new_n19560_, new_n19561_, new_n19562_, new_n19563_,
    new_n19564_, new_n19565_, new_n19566_, new_n19567_, new_n19568_,
    new_n19569_, new_n19570_, new_n19571_, new_n19572_, new_n19573_,
    new_n19574_, new_n19575_, new_n19576_, new_n19577_, new_n19578_,
    new_n19579_, new_n19580_, new_n19581_, new_n19582_, new_n19583_,
    new_n19584_, new_n19585_, new_n19586_, new_n19587_, new_n19588_,
    new_n19589_, new_n19590_, new_n19591_, new_n19592_, new_n19593_,
    new_n19594_, new_n19595_, new_n19596_, new_n19597_, new_n19598_,
    new_n19599_, new_n19600_, new_n19601_, new_n19602_, new_n19603_,
    new_n19604_, new_n19605_, new_n19606_, new_n19607_, new_n19608_,
    new_n19609_, new_n19610_, new_n19611_, new_n19612_, new_n19613_,
    new_n19614_, new_n19615_, new_n19616_, new_n19617_, new_n19618_,
    new_n19619_, new_n19620_, new_n19621_, new_n19622_, new_n19623_,
    new_n19624_, new_n19625_, new_n19626_, new_n19627_, new_n19628_,
    new_n19629_, new_n19630_, new_n19631_, new_n19632_, new_n19633_,
    new_n19634_, new_n19635_, new_n19636_, new_n19637_, new_n19638_,
    new_n19639_, new_n19640_, new_n19641_, new_n19642_, new_n19643_,
    new_n19644_, new_n19645_, new_n19646_, new_n19647_, new_n19648_,
    new_n19649_, new_n19650_, new_n19651_, new_n19652_, new_n19653_,
    new_n19654_, new_n19655_, new_n19656_, new_n19657_, new_n19658_,
    new_n19659_, new_n19660_, new_n19661_, new_n19662_, new_n19663_,
    new_n19664_, new_n19665_, new_n19666_, new_n19667_, new_n19668_,
    new_n19669_, new_n19670_, new_n19671_, new_n19672_, new_n19673_,
    new_n19674_, new_n19675_, new_n19676_, new_n19677_, new_n19678_,
    new_n19679_, new_n19680_, new_n19681_, new_n19682_, new_n19683_,
    new_n19684_, new_n19685_, new_n19686_, new_n19687_, new_n19688_,
    new_n19689_, new_n19690_, new_n19691_, new_n19692_, new_n19693_,
    new_n19694_, new_n19695_, new_n19696_, new_n19697_, new_n19698_,
    new_n19699_, new_n19700_, new_n19701_, new_n19702_, new_n19703_,
    new_n19704_, new_n19705_, new_n19706_, new_n19707_, new_n19708_,
    new_n19709_, new_n19710_, new_n19711_, new_n19712_, new_n19713_,
    new_n19714_, new_n19715_, new_n19716_, new_n19717_, new_n19718_,
    new_n19719_, new_n19720_, new_n19721_, new_n19722_, new_n19723_,
    new_n19724_, new_n19725_, new_n19726_, new_n19727_, new_n19728_,
    new_n19729_, new_n19730_, new_n19731_, new_n19732_, new_n19733_,
    new_n19734_, new_n19735_, new_n19736_, new_n19737_, new_n19738_,
    new_n19739_, new_n19740_, new_n19741_, new_n19742_, new_n19743_,
    new_n19744_, new_n19745_, new_n19746_, new_n19747_, new_n19748_,
    new_n19749_, new_n19750_, new_n19751_, new_n19752_, new_n19753_,
    new_n19754_, new_n19755_, new_n19756_, new_n19757_, new_n19758_,
    new_n19759_, new_n19760_, new_n19761_, new_n19762_, new_n19763_,
    new_n19764_, new_n19765_, new_n19766_, new_n19767_, new_n19768_,
    new_n19769_, new_n19770_, new_n19771_, new_n19772_, new_n19773_,
    new_n19774_, new_n19775_, new_n19776_, new_n19777_, new_n19778_,
    new_n19779_, new_n19780_, new_n19781_, new_n19782_, new_n19783_,
    new_n19784_, new_n19785_, new_n19786_, new_n19787_, new_n19788_,
    new_n19789_, new_n19790_, new_n19791_, new_n19792_, new_n19793_,
    new_n19794_, new_n19795_, new_n19796_, new_n19797_, new_n19798_,
    new_n19799_, new_n19800_, new_n19801_, new_n19802_, new_n19803_,
    new_n19804_, new_n19805_, new_n19806_, new_n19807_, new_n19808_,
    new_n19809_, new_n19810_, new_n19811_, new_n19812_, new_n19813_,
    new_n19814_, new_n19815_, new_n19816_, new_n19817_, new_n19818_,
    new_n19819_, new_n19820_, new_n19821_, new_n19822_, new_n19823_,
    new_n19824_, new_n19825_, new_n19826_, new_n19827_, new_n19828_,
    new_n19829_, new_n19830_, new_n19831_, new_n19832_, new_n19833_,
    new_n19834_, new_n19835_, new_n19836_, new_n19837_, new_n19838_,
    new_n19839_, new_n19840_, new_n19841_, new_n19842_, new_n19843_,
    new_n19844_, new_n19845_, new_n19846_, new_n19847_, new_n19848_,
    new_n19849_, new_n19850_, new_n19851_, new_n19852_, new_n19853_,
    new_n19854_, new_n19855_, new_n19856_, new_n19857_, new_n19858_,
    new_n19859_, new_n19860_, new_n19861_, new_n19862_, new_n19863_,
    new_n19864_, new_n19865_, new_n19866_, new_n19867_, new_n19868_,
    new_n19869_, new_n19870_, new_n19871_, new_n19872_, new_n19873_,
    new_n19874_, new_n19875_, new_n19876_, new_n19877_, new_n19878_,
    new_n19879_, new_n19880_, new_n19881_, new_n19882_, new_n19883_,
    new_n19884_, new_n19885_, new_n19886_, new_n19887_, new_n19888_,
    new_n19889_, new_n19890_, new_n19892_, new_n19893_, new_n19894_,
    new_n19895_, new_n19896_, new_n19897_, new_n19898_, new_n19899_,
    new_n19900_, new_n19901_, new_n19902_, new_n19903_, new_n19904_,
    new_n19905_, new_n19906_, new_n19907_, new_n19908_, new_n19909_,
    new_n19910_, new_n19911_, new_n19912_, new_n19913_, new_n19914_,
    new_n19915_, new_n19916_, new_n19917_, new_n19918_, new_n19919_,
    new_n19920_, new_n19921_, new_n19922_, new_n19923_, new_n19924_,
    new_n19925_, new_n19926_, new_n19927_, new_n19928_, new_n19929_,
    new_n19930_, new_n19931_, new_n19932_, new_n19933_, new_n19934_,
    new_n19935_, new_n19936_, new_n19937_, new_n19938_, new_n19939_,
    new_n19940_, new_n19941_, new_n19942_, new_n19943_, new_n19944_,
    new_n19945_, new_n19946_, new_n19947_, new_n19948_, new_n19949_,
    new_n19950_, new_n19951_, new_n19952_, new_n19953_, new_n19954_,
    new_n19955_, new_n19956_, new_n19957_, new_n19958_, new_n19959_,
    new_n19960_, new_n19961_, new_n19962_, new_n19963_, new_n19964_,
    new_n19965_, new_n19966_, new_n19967_, new_n19968_, new_n19969_,
    new_n19970_, new_n19971_, new_n19972_, new_n19973_, new_n19974_,
    new_n19975_, new_n19976_, new_n19977_, new_n19978_, new_n19979_,
    new_n19980_, new_n19981_, new_n19982_, new_n19983_, new_n19984_,
    new_n19985_, new_n19986_, new_n19987_, new_n19988_, new_n19989_,
    new_n19990_, new_n19991_, new_n19992_, new_n19993_, new_n19994_,
    new_n19995_, new_n19996_, new_n19997_, new_n19998_, new_n19999_,
    new_n20000_, new_n20001_, new_n20002_, new_n20003_, new_n20004_,
    new_n20005_, new_n20006_, new_n20007_, new_n20008_, new_n20009_,
    new_n20010_, new_n20011_, new_n20012_, new_n20013_, new_n20014_,
    new_n20015_, new_n20016_, new_n20017_, new_n20018_, new_n20019_,
    new_n20020_, new_n20021_, new_n20022_, new_n20023_, new_n20024_,
    new_n20025_, new_n20026_, new_n20027_, new_n20028_, new_n20029_,
    new_n20030_, new_n20031_, new_n20032_, new_n20033_, new_n20034_,
    new_n20035_, new_n20036_, new_n20037_, new_n20038_, new_n20039_,
    new_n20040_, new_n20041_, new_n20042_, new_n20043_, new_n20044_,
    new_n20045_, new_n20046_, new_n20047_, new_n20048_, new_n20049_,
    new_n20050_, new_n20051_, new_n20052_, new_n20053_, new_n20054_,
    new_n20055_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20103_, new_n20104_,
    new_n20105_, new_n20106_, new_n20107_, new_n20108_, new_n20109_,
    new_n20110_, new_n20111_, new_n20112_, new_n20113_, new_n20114_,
    new_n20115_, new_n20116_, new_n20117_, new_n20118_, new_n20119_,
    new_n20120_, new_n20121_, new_n20122_, new_n20123_, new_n20124_,
    new_n20125_, new_n20126_, new_n20127_, new_n20128_, new_n20129_,
    new_n20130_, new_n20131_, new_n20132_, new_n20133_, new_n20134_,
    new_n20135_, new_n20136_, new_n20137_, new_n20138_, new_n20139_,
    new_n20140_, new_n20141_, new_n20142_, new_n20143_, new_n20144_,
    new_n20145_, new_n20146_, new_n20147_, new_n20148_, new_n20149_,
    new_n20150_, new_n20151_, new_n20152_, new_n20153_, new_n20154_,
    new_n20155_, new_n20156_, new_n20157_, new_n20158_, new_n20159_,
    new_n20160_, new_n20161_, new_n20162_, new_n20163_, new_n20164_,
    new_n20165_, new_n20166_, new_n20167_, new_n20168_, new_n20169_,
    new_n20170_, new_n20171_, new_n20172_, new_n20173_, new_n20174_,
    new_n20175_, new_n20176_, new_n20177_, new_n20178_, new_n20179_,
    new_n20180_, new_n20181_, new_n20182_, new_n20183_, new_n20184_,
    new_n20185_, new_n20186_, new_n20187_, new_n20188_, new_n20189_,
    new_n20190_, new_n20191_, new_n20192_, new_n20193_, new_n20194_,
    new_n20195_, new_n20196_, new_n20197_, new_n20198_, new_n20199_,
    new_n20200_, new_n20201_, new_n20202_, new_n20203_, new_n20204_,
    new_n20205_, new_n20206_, new_n20207_, new_n20208_, new_n20209_,
    new_n20210_, new_n20211_, new_n20212_, new_n20213_, new_n20214_,
    new_n20215_, new_n20216_, new_n20217_, new_n20218_, new_n20219_,
    new_n20220_, new_n20221_, new_n20222_, new_n20223_, new_n20224_,
    new_n20225_, new_n20226_, new_n20227_, new_n20228_, new_n20229_,
    new_n20230_, new_n20231_, new_n20232_, new_n20233_, new_n20234_,
    new_n20235_, new_n20236_, new_n20237_, new_n20238_, new_n20239_,
    new_n20240_, new_n20241_, new_n20242_, new_n20243_, new_n20244_,
    new_n20245_, new_n20246_, new_n20247_, new_n20248_, new_n20249_,
    new_n20250_, new_n20251_, new_n20252_, new_n20253_, new_n20254_,
    new_n20255_, new_n20256_, new_n20257_, new_n20258_, new_n20259_,
    new_n20260_, new_n20261_, new_n20262_, new_n20263_, new_n20264_,
    new_n20265_, new_n20266_, new_n20267_, new_n20268_, new_n20269_,
    new_n20270_, new_n20271_, new_n20272_, new_n20273_, new_n20274_,
    new_n20275_, new_n20276_, new_n20277_, new_n20278_, new_n20279_,
    new_n20280_, new_n20281_, new_n20282_, new_n20283_, new_n20284_,
    new_n20285_, new_n20286_, new_n20287_, new_n20288_, new_n20289_,
    new_n20290_, new_n20291_, new_n20292_, new_n20293_, new_n20294_,
    new_n20295_, new_n20296_, new_n20297_, new_n20298_, new_n20299_,
    new_n20300_, new_n20301_, new_n20302_, new_n20303_, new_n20304_,
    new_n20305_, new_n20306_, new_n20307_, new_n20308_, new_n20309_,
    new_n20310_, new_n20311_, new_n20312_, new_n20313_, new_n20314_,
    new_n20315_, new_n20316_, new_n20317_, new_n20318_, new_n20319_,
    new_n20320_, new_n20321_, new_n20322_, new_n20323_, new_n20324_,
    new_n20325_, new_n20326_, new_n20327_, new_n20328_, new_n20329_,
    new_n20330_, new_n20331_, new_n20332_, new_n20333_, new_n20334_,
    new_n20335_, new_n20336_, new_n20337_, new_n20338_, new_n20339_,
    new_n20340_, new_n20341_, new_n20342_, new_n20343_, new_n20344_,
    new_n20345_, new_n20346_, new_n20347_, new_n20348_, new_n20349_,
    new_n20350_, new_n20351_, new_n20352_, new_n20353_, new_n20354_,
    new_n20355_, new_n20356_, new_n20357_, new_n20358_, new_n20359_,
    new_n20360_, new_n20361_, new_n20362_, new_n20363_, new_n20364_,
    new_n20365_, new_n20366_, new_n20367_, new_n20368_, new_n20369_,
    new_n20370_, new_n20371_, new_n20372_, new_n20373_, new_n20374_,
    new_n20375_, new_n20376_, new_n20377_, new_n20378_, new_n20379_,
    new_n20380_, new_n20381_, new_n20382_, new_n20383_, new_n20384_,
    new_n20385_, new_n20386_, new_n20387_, new_n20388_, new_n20389_,
    new_n20390_, new_n20391_, new_n20392_, new_n20393_, new_n20394_,
    new_n20395_, new_n20396_, new_n20397_, new_n20398_, new_n20399_,
    new_n20400_, new_n20401_, new_n20402_, new_n20403_, new_n20404_,
    new_n20405_, new_n20406_, new_n20407_, new_n20408_, new_n20409_,
    new_n20411_, new_n20412_, new_n20413_, new_n20414_, new_n20415_,
    new_n20416_, new_n20417_, new_n20418_, new_n20419_, new_n20420_,
    new_n20421_, new_n20422_, new_n20423_, new_n20424_, new_n20425_,
    new_n20426_, new_n20427_, new_n20428_, new_n20429_, new_n20430_,
    new_n20431_, new_n20432_, new_n20433_, new_n20434_, new_n20435_,
    new_n20436_, new_n20437_, new_n20438_, new_n20439_, new_n20440_,
    new_n20441_, new_n20442_, new_n20443_, new_n20444_, new_n20445_,
    new_n20446_, new_n20447_, new_n20448_, new_n20449_, new_n20450_,
    new_n20451_, new_n20452_, new_n20453_, new_n20454_, new_n20455_,
    new_n20456_, new_n20457_, new_n20458_, new_n20459_, new_n20460_,
    new_n20461_, new_n20462_, new_n20463_, new_n20464_, new_n20465_,
    new_n20466_, new_n20467_, new_n20468_, new_n20469_, new_n20470_,
    new_n20471_, new_n20472_, new_n20473_, new_n20474_, new_n20475_,
    new_n20476_, new_n20477_, new_n20478_, new_n20479_, new_n20480_,
    new_n20481_, new_n20482_, new_n20483_, new_n20484_, new_n20485_,
    new_n20486_, new_n20487_, new_n20488_, new_n20489_, new_n20490_,
    new_n20491_, new_n20492_, new_n20493_, new_n20494_, new_n20495_,
    new_n20496_, new_n20497_, new_n20498_, new_n20499_, new_n20500_,
    new_n20501_, new_n20502_, new_n20503_, new_n20504_, new_n20505_,
    new_n20506_, new_n20507_, new_n20508_, new_n20509_, new_n20510_,
    new_n20511_, new_n20512_, new_n20513_, new_n20514_, new_n20515_,
    new_n20516_, new_n20517_, new_n20518_, new_n20519_, new_n20520_,
    new_n20521_, new_n20522_, new_n20523_, new_n20524_, new_n20525_,
    new_n20526_, new_n20527_, new_n20528_, new_n20529_, new_n20530_,
    new_n20531_, new_n20532_, new_n20533_, new_n20534_, new_n20535_,
    new_n20536_, new_n20537_, new_n20538_, new_n20539_, new_n20540_,
    new_n20541_, new_n20542_, new_n20543_, new_n20544_, new_n20545_,
    new_n20546_, new_n20547_, new_n20548_, new_n20549_, new_n20550_,
    new_n20551_, new_n20552_, new_n20553_, new_n20554_, new_n20555_,
    new_n20556_, new_n20557_, new_n20558_, new_n20559_, new_n20560_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20569_, new_n20570_,
    new_n20571_, new_n20572_, new_n20573_, new_n20574_, new_n20575_,
    new_n20576_, new_n20577_, new_n20578_, new_n20579_, new_n20580_,
    new_n20581_, new_n20582_, new_n20583_, new_n20584_, new_n20585_,
    new_n20586_, new_n20587_, new_n20588_, new_n20589_, new_n20590_,
    new_n20591_, new_n20592_, new_n20593_, new_n20594_, new_n20595_,
    new_n20596_, new_n20597_, new_n20598_, new_n20599_, new_n20600_,
    new_n20601_, new_n20602_, new_n20603_, new_n20604_, new_n20605_,
    new_n20606_, new_n20607_, new_n20608_, new_n20609_, new_n20610_,
    new_n20611_, new_n20612_, new_n20613_, new_n20614_, new_n20615_,
    new_n20616_, new_n20617_, new_n20618_, new_n20619_, new_n20620_,
    new_n20621_, new_n20622_, new_n20623_, new_n20624_, new_n20625_,
    new_n20626_, new_n20627_, new_n20628_, new_n20629_, new_n20630_,
    new_n20631_, new_n20632_, new_n20633_, new_n20634_, new_n20635_,
    new_n20636_, new_n20637_, new_n20638_, new_n20639_, new_n20640_,
    new_n20641_, new_n20642_, new_n20643_, new_n20644_, new_n20645_,
    new_n20646_, new_n20647_, new_n20648_, new_n20649_, new_n20650_,
    new_n20651_, new_n20652_, new_n20653_, new_n20654_, new_n20655_,
    new_n20656_, new_n20657_, new_n20658_, new_n20659_, new_n20660_,
    new_n20661_, new_n20662_, new_n20663_, new_n20664_, new_n20665_,
    new_n20666_, new_n20667_, new_n20668_, new_n20669_, new_n20670_,
    new_n20671_, new_n20672_, new_n20673_, new_n20674_, new_n20675_,
    new_n20676_, new_n20677_, new_n20678_, new_n20679_, new_n20680_,
    new_n20681_, new_n20682_, new_n20683_, new_n20684_, new_n20685_,
    new_n20686_, new_n20687_, new_n20688_, new_n20689_, new_n20690_,
    new_n20691_, new_n20692_, new_n20693_, new_n20694_, new_n20695_,
    new_n20696_, new_n20697_, new_n20698_, new_n20699_, new_n20700_,
    new_n20701_, new_n20702_, new_n20703_, new_n20704_, new_n20705_,
    new_n20706_, new_n20707_, new_n20708_, new_n20709_, new_n20710_,
    new_n20711_, new_n20712_, new_n20713_, new_n20714_, new_n20715_,
    new_n20716_, new_n20717_, new_n20718_, new_n20719_, new_n20720_,
    new_n20721_, new_n20722_, new_n20723_, new_n20724_, new_n20725_,
    new_n20726_, new_n20727_, new_n20728_, new_n20729_, new_n20730_,
    new_n20731_, new_n20732_, new_n20733_, new_n20734_, new_n20735_,
    new_n20736_, new_n20737_, new_n20738_, new_n20739_, new_n20740_,
    new_n20741_, new_n20742_, new_n20743_, new_n20744_, new_n20745_,
    new_n20746_, new_n20747_, new_n20748_, new_n20749_, new_n20750_,
    new_n20751_, new_n20752_, new_n20753_, new_n20754_, new_n20755_,
    new_n20756_, new_n20757_, new_n20758_, new_n20759_, new_n20760_,
    new_n20761_, new_n20762_, new_n20763_, new_n20764_, new_n20765_,
    new_n20766_, new_n20767_, new_n20768_, new_n20769_, new_n20770_,
    new_n20771_, new_n20772_, new_n20773_, new_n20774_, new_n20775_,
    new_n20776_, new_n20777_, new_n20778_, new_n20779_, new_n20780_,
    new_n20781_, new_n20782_, new_n20783_, new_n20784_, new_n20785_,
    new_n20786_, new_n20787_, new_n20788_, new_n20789_, new_n20790_,
    new_n20791_, new_n20792_, new_n20793_, new_n20794_, new_n20795_,
    new_n20796_, new_n20797_, new_n20798_, new_n20799_, new_n20800_,
    new_n20801_, new_n20802_, new_n20803_, new_n20804_, new_n20805_,
    new_n20806_, new_n20807_, new_n20808_, new_n20809_, new_n20810_,
    new_n20811_, new_n20812_, new_n20813_, new_n20814_, new_n20815_,
    new_n20816_, new_n20817_, new_n20818_, new_n20819_, new_n20820_,
    new_n20821_, new_n20822_, new_n20823_, new_n20824_, new_n20825_,
    new_n20826_, new_n20827_, new_n20828_, new_n20829_, new_n20830_,
    new_n20831_, new_n20832_, new_n20833_, new_n20834_, new_n20835_,
    new_n20836_, new_n20837_, new_n20838_, new_n20839_, new_n20840_,
    new_n20841_, new_n20842_, new_n20843_, new_n20844_, new_n20845_,
    new_n20846_, new_n20847_, new_n20848_, new_n20849_, new_n20850_,
    new_n20851_, new_n20852_, new_n20853_, new_n20854_, new_n20855_,
    new_n20856_, new_n20857_, new_n20858_, new_n20859_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20899_, new_n20900_, new_n20901_,
    new_n20902_, new_n20903_, new_n20904_, new_n20905_, new_n20906_,
    new_n20907_, new_n20908_, new_n20909_, new_n20910_, new_n20911_,
    new_n20912_, new_n20913_, new_n20914_, new_n20915_, new_n20916_,
    new_n20917_, new_n20918_, new_n20919_, new_n20920_, new_n20921_,
    new_n20922_, new_n20923_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20969_, new_n20970_, new_n20971_,
    new_n20972_, new_n20973_, new_n20974_, new_n20975_, new_n20976_,
    new_n20977_, new_n20978_, new_n20980_, new_n20981_, new_n20982_,
    new_n20983_, new_n20984_, new_n20985_, new_n20986_, new_n20987_,
    new_n20988_, new_n20989_, new_n20990_, new_n20991_, new_n20992_,
    new_n20993_, new_n20994_, new_n20995_, new_n20996_, new_n20997_,
    new_n20998_, new_n20999_, new_n21000_, new_n21001_, new_n21002_,
    new_n21003_, new_n21004_, new_n21005_, new_n21006_, new_n21007_,
    new_n21008_, new_n21009_, new_n21010_, new_n21011_, new_n21012_,
    new_n21013_, new_n21014_, new_n21015_, new_n21016_, new_n21017_,
    new_n21018_, new_n21019_, new_n21020_, new_n21021_, new_n21022_,
    new_n21023_, new_n21024_, new_n21025_, new_n21026_, new_n21027_,
    new_n21028_, new_n21029_, new_n21030_, new_n21031_, new_n21032_,
    new_n21033_, new_n21034_, new_n21035_, new_n21036_, new_n21037_,
    new_n21038_, new_n21039_, new_n21040_, new_n21041_, new_n21042_,
    new_n21043_, new_n21044_, new_n21045_, new_n21046_, new_n21047_,
    new_n21048_, new_n21049_, new_n21050_, new_n21051_, new_n21052_,
    new_n21053_, new_n21054_, new_n21055_, new_n21056_, new_n21057_,
    new_n21058_, new_n21059_, new_n21060_, new_n21061_, new_n21062_,
    new_n21063_, new_n21064_, new_n21065_, new_n21066_, new_n21067_,
    new_n21068_, new_n21069_, new_n21070_, new_n21071_, new_n21072_,
    new_n21073_, new_n21074_, new_n21075_, new_n21076_, new_n21077_,
    new_n21078_, new_n21079_, new_n21080_, new_n21081_, new_n21082_,
    new_n21083_, new_n21084_, new_n21085_, new_n21086_, new_n21087_,
    new_n21088_, new_n21089_, new_n21090_, new_n21091_, new_n21092_,
    new_n21093_, new_n21094_, new_n21095_, new_n21096_, new_n21097_,
    new_n21098_, new_n21099_, new_n21100_, new_n21101_, new_n21102_,
    new_n21103_, new_n21104_, new_n21105_, new_n21106_, new_n21107_,
    new_n21108_, new_n21109_, new_n21110_, new_n21111_, new_n21112_,
    new_n21113_, new_n21114_, new_n21115_, new_n21116_, new_n21117_,
    new_n21118_, new_n21119_, new_n21120_, new_n21121_, new_n21122_,
    new_n21123_, new_n21124_, new_n21125_, new_n21126_, new_n21127_,
    new_n21129_, new_n21130_, new_n21131_, new_n21132_, new_n21133_,
    new_n21134_, new_n21135_, new_n21136_, new_n21137_, new_n21138_,
    new_n21139_, new_n21140_, new_n21141_, new_n21142_, new_n21143_,
    new_n21144_, new_n21145_, new_n21146_, new_n21147_, new_n21148_,
    new_n21149_, new_n21150_, new_n21151_, new_n21152_, new_n21153_,
    new_n21154_, new_n21155_, new_n21156_, new_n21157_, new_n21158_,
    new_n21159_, new_n21160_, new_n21161_, new_n21162_, new_n21163_,
    new_n21164_, new_n21165_, new_n21166_, new_n21167_, new_n21168_,
    new_n21169_, new_n21170_, new_n21171_, new_n21172_, new_n21173_,
    new_n21174_, new_n21175_, new_n21176_, new_n21177_, new_n21178_,
    new_n21179_, new_n21180_, new_n21181_, new_n21182_, new_n21183_,
    new_n21184_, new_n21185_, new_n21186_, new_n21187_, new_n21188_,
    new_n21189_, new_n21190_, new_n21191_, new_n21193_, new_n21194_,
    new_n21195_, new_n21196_, new_n21197_, new_n21198_, new_n21199_,
    new_n21200_, new_n21201_, new_n21202_, new_n21203_, new_n21204_,
    new_n21205_, new_n21206_, new_n21207_, new_n21208_, new_n21209_,
    new_n21210_, new_n21211_, new_n21212_, new_n21213_, new_n21214_,
    new_n21215_, new_n21216_, new_n21217_, new_n21218_, new_n21219_,
    new_n21220_, new_n21221_, new_n21222_, new_n21223_, new_n21224_,
    new_n21225_, new_n21226_, new_n21227_, new_n21228_, new_n21229_,
    new_n21230_, new_n21231_, new_n21232_, new_n21233_, new_n21234_,
    new_n21235_, new_n21236_, new_n21237_, new_n21238_, new_n21239_,
    new_n21240_, new_n21241_, new_n21242_, new_n21243_, new_n21244_,
    new_n21245_, new_n21246_, new_n21247_, new_n21248_, new_n21249_,
    new_n21250_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21281_, new_n21282_, new_n21283_, new_n21284_, new_n21285_,
    new_n21286_, new_n21287_, new_n21288_, new_n21289_, new_n21290_,
    new_n21291_, new_n21292_, new_n21293_, new_n21294_, new_n21295_,
    new_n21296_, new_n21297_, new_n21298_, new_n21299_, new_n21300_,
    new_n21301_, new_n21302_, new_n21303_, new_n21304_, new_n21305_,
    new_n21306_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21386_, new_n21387_,
    new_n21388_, new_n21389_, new_n21390_, new_n21391_, new_n21392_,
    new_n21393_, new_n21394_, new_n21395_, new_n21396_, new_n21397_,
    new_n21398_, new_n21399_, new_n21400_, new_n21401_, new_n21402_,
    new_n21403_, new_n21404_, new_n21405_, new_n21406_, new_n21407_,
    new_n21408_, new_n21409_, new_n21410_, new_n21411_, new_n21412_,
    new_n21413_, new_n21414_, new_n21415_, new_n21416_, new_n21417_,
    new_n21418_, new_n21419_, new_n21420_, new_n21421_, new_n21422_,
    new_n21423_, new_n21424_, new_n21425_, new_n21426_, new_n21427_,
    new_n21428_, new_n21429_, new_n21430_, new_n21431_, new_n21432_,
    new_n21433_, new_n21434_, new_n21435_, new_n21436_, new_n21437_,
    new_n21438_, new_n21439_, new_n21440_, new_n21441_, new_n21442_,
    new_n21443_, new_n21444_, new_n21445_, new_n21446_, new_n21447_,
    new_n21448_, new_n21449_, new_n21450_, new_n21451_, new_n21452_,
    new_n21453_, new_n21454_, new_n21455_, new_n21456_, new_n21457_,
    new_n21458_, new_n21459_, new_n21460_, new_n21461_, new_n21462_,
    new_n21463_, new_n21464_, new_n21465_, new_n21466_, new_n21467_,
    new_n21468_, new_n21469_, new_n21470_, new_n21471_, new_n21472_,
    new_n21473_, new_n21474_, new_n21475_, new_n21476_, new_n21477_,
    new_n21478_, new_n21479_, new_n21480_, new_n21481_, new_n21482_,
    new_n21483_, new_n21484_, new_n21485_, new_n21486_, new_n21487_,
    new_n21489_, new_n21490_, new_n21491_, new_n21492_, new_n21493_,
    new_n21494_, new_n21495_, new_n21496_, new_n21497_, new_n21498_,
    new_n21499_, new_n21500_, new_n21501_, new_n21502_, new_n21503_,
    new_n21504_, new_n21505_, new_n21506_, new_n21507_, new_n21508_,
    new_n21509_, new_n21510_, new_n21511_, new_n21512_, new_n21513_,
    new_n21514_, new_n21515_, new_n21516_, new_n21517_, new_n21518_,
    new_n21519_, new_n21520_, new_n21521_, new_n21522_, new_n21523_,
    new_n21524_, new_n21525_, new_n21526_, new_n21527_, new_n21528_,
    new_n21529_, new_n21530_, new_n21531_, new_n21532_, new_n21533_,
    new_n21534_, new_n21535_, new_n21536_, new_n21537_, new_n21538_,
    new_n21539_, new_n21540_, new_n21541_, new_n21542_, new_n21543_,
    new_n21544_, new_n21545_, new_n21546_, new_n21547_, new_n21548_,
    new_n21549_, new_n21550_, new_n21551_, new_n21552_, new_n21553_,
    new_n21554_, new_n21555_, new_n21556_, new_n21557_, new_n21558_,
    new_n21559_, new_n21560_, new_n21561_, new_n21562_, new_n21563_,
    new_n21564_, new_n21565_, new_n21566_, new_n21567_, new_n21568_,
    new_n21570_, new_n21571_, new_n21572_, new_n21573_, new_n21574_,
    new_n21575_, new_n21576_, new_n21577_, new_n21578_, new_n21579_,
    new_n21580_, new_n21581_, new_n21582_, new_n21583_, new_n21584_,
    new_n21585_, new_n21586_, new_n21587_, new_n21588_, new_n21589_,
    new_n21590_, new_n21591_, new_n21592_, new_n21593_, new_n21594_,
    new_n21595_, new_n21596_, new_n21597_, new_n21598_, new_n21599_,
    new_n21600_, new_n21601_, new_n21602_, new_n21603_, new_n21604_,
    new_n21605_, new_n21606_, new_n21607_, new_n21608_, new_n21609_,
    new_n21610_, new_n21611_, new_n21612_, new_n21613_, new_n21614_,
    new_n21615_, new_n21616_, new_n21617_, new_n21618_, new_n21619_,
    new_n21620_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21630_,
    new_n21631_, new_n21632_, new_n21633_, new_n21634_, new_n21635_,
    new_n21636_, new_n21637_, new_n21638_, new_n21639_, new_n21640_,
    new_n21641_, new_n21642_, new_n21643_, new_n21644_, new_n21645_,
    new_n21646_, new_n21647_, new_n21648_, new_n21649_, new_n21650_,
    new_n21651_, new_n21652_, new_n21653_, new_n21654_, new_n21655_,
    new_n21656_, new_n21657_, new_n21658_, new_n21659_, new_n21660_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21692_,
    new_n21693_, new_n21694_, new_n21695_, new_n21696_, new_n21697_,
    new_n21698_, new_n21699_, new_n21700_, new_n21701_, new_n21702_,
    new_n21703_, new_n21704_, new_n21705_, new_n21706_, new_n21707_,
    new_n21708_, new_n21709_, new_n21710_, new_n21711_, new_n21712_,
    new_n21713_, new_n21714_, new_n21715_, new_n21716_, new_n21717_,
    new_n21718_, new_n21719_, new_n21720_, new_n21721_, new_n21722_,
    new_n21723_, new_n21724_, new_n21725_, new_n21726_, new_n21727_,
    new_n21728_, new_n21729_, new_n21730_, new_n21731_, new_n21732_,
    new_n21733_, new_n21734_, new_n21735_, new_n21736_, new_n21737_,
    new_n21738_, new_n21739_, new_n21740_, new_n21741_, new_n21742_,
    new_n21743_, new_n21744_, new_n21745_, new_n21746_, new_n21747_,
    new_n21749_, new_n21750_, new_n21751_, new_n21752_, new_n21753_,
    new_n21754_, new_n21755_, new_n21756_, new_n21757_, new_n21758_,
    new_n21759_, new_n21760_, new_n21761_, new_n21762_, new_n21763_,
    new_n21764_, new_n21765_, new_n21766_, new_n21767_, new_n21768_,
    new_n21769_, new_n21770_, new_n21771_, new_n21772_, new_n21773_,
    new_n21774_, new_n21775_, new_n21776_, new_n21777_, new_n21778_,
    new_n21779_, new_n21780_, new_n21781_, new_n21782_, new_n21783_,
    new_n21784_, new_n21785_, new_n21786_, new_n21787_, new_n21788_,
    new_n21789_, new_n21790_, new_n21791_, new_n21792_, new_n21793_,
    new_n21794_, new_n21795_, new_n21796_, new_n21797_, new_n21798_,
    new_n21799_, new_n21800_, new_n21801_, new_n21802_, new_n21803_,
    new_n21805_, new_n21806_, new_n21807_, new_n21808_, new_n21809_,
    new_n21810_, new_n21811_, new_n21812_, new_n21813_, new_n21814_,
    new_n21815_, new_n21816_, new_n21817_, new_n21818_, new_n21819_,
    new_n21820_, new_n21821_, new_n21822_, new_n21823_, new_n21824_,
    new_n21825_, new_n21826_, new_n21827_, new_n21828_, new_n21829_,
    new_n21830_, new_n21831_, new_n21832_, new_n21833_, new_n21834_,
    new_n21835_, new_n21836_, new_n21837_, new_n21838_, new_n21839_,
    new_n21840_, new_n21841_, new_n21842_, new_n21843_, new_n21844_,
    new_n21845_, new_n21846_, new_n21847_, new_n21848_, new_n21849_,
    new_n21850_, new_n21851_, new_n21852_, new_n21853_, new_n21854_,
    new_n21855_, new_n21856_, new_n21857_, new_n21858_, new_n21859_,
    new_n21861_, new_n21862_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21880_,
    new_n21881_, new_n21882_, new_n21883_, new_n21884_, new_n21885_,
    new_n21886_, new_n21887_, new_n21888_, new_n21889_, new_n21890_,
    new_n21891_, new_n21892_, new_n21893_, new_n21894_, new_n21895_,
    new_n21896_, new_n21897_, new_n21898_, new_n21899_, new_n21900_,
    new_n21901_, new_n21902_, new_n21903_, new_n21904_, new_n21905_,
    new_n21906_, new_n21907_, new_n21908_, new_n21909_, new_n21910_,
    new_n21911_, new_n21912_, new_n21913_, new_n21914_, new_n21915_,
    new_n21916_, new_n21917_, new_n21918_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22015_, new_n22016_, new_n22017_,
    new_n22018_, new_n22019_, new_n22020_, new_n22021_, new_n22022_,
    new_n22023_, new_n22024_, new_n22025_, new_n22026_, new_n22027_,
    new_n22028_, new_n22029_, new_n22030_, new_n22031_, new_n22032_,
    new_n22033_, new_n22034_, new_n22035_, new_n22036_, new_n22037_,
    new_n22038_, new_n22039_, new_n22040_, new_n22041_, new_n22042_,
    new_n22043_, new_n22044_, new_n22045_, new_n22046_, new_n22047_,
    new_n22048_, new_n22049_, new_n22050_, new_n22051_, new_n22052_,
    new_n22053_, new_n22054_, new_n22055_, new_n22056_, new_n22057_,
    new_n22058_, new_n22059_, new_n22060_, new_n22061_, new_n22062_,
    new_n22063_, new_n22064_, new_n22065_, new_n22066_, new_n22067_,
    new_n22068_, new_n22070_, new_n22071_, new_n22072_, new_n22073_,
    new_n22074_, new_n22075_, new_n22076_, new_n22077_, new_n22078_,
    new_n22079_, new_n22080_, new_n22081_, new_n22082_, new_n22083_,
    new_n22084_, new_n22085_, new_n22086_, new_n22087_, new_n22088_,
    new_n22089_, new_n22090_, new_n22091_, new_n22092_, new_n22093_,
    new_n22094_, new_n22095_, new_n22096_, new_n22097_, new_n22098_,
    new_n22099_, new_n22100_, new_n22101_, new_n22102_, new_n22103_,
    new_n22104_, new_n22105_, new_n22106_, new_n22107_, new_n22108_,
    new_n22109_, new_n22110_, new_n22111_, new_n22112_, new_n22113_,
    new_n22114_, new_n22115_, new_n22116_, new_n22117_, new_n22118_,
    new_n22119_, new_n22120_, new_n22121_, new_n22122_, new_n22123_,
    new_n22124_, new_n22125_, new_n22126_, new_n22128_, new_n22129_,
    new_n22130_, new_n22131_, new_n22132_, new_n22133_, new_n22134_,
    new_n22135_, new_n22136_, new_n22137_, new_n22138_, new_n22139_,
    new_n22140_, new_n22141_, new_n22142_, new_n22143_, new_n22144_,
    new_n22145_, new_n22146_, new_n22147_, new_n22148_, new_n22149_,
    new_n22150_, new_n22151_, new_n22152_, new_n22153_, new_n22154_,
    new_n22155_, new_n22156_, new_n22157_, new_n22158_, new_n22159_,
    new_n22160_, new_n22161_, new_n22162_, new_n22163_, new_n22164_,
    new_n22165_, new_n22166_, new_n22168_, new_n22169_, new_n22170_,
    new_n22171_, new_n22172_, new_n22173_, new_n22174_, new_n22175_,
    new_n22176_, new_n22177_, new_n22178_, new_n22179_, new_n22180_,
    new_n22181_, new_n22182_, new_n22183_, new_n22184_, new_n22185_,
    new_n22186_, new_n22187_, new_n22188_, new_n22189_, new_n22190_,
    new_n22191_, new_n22192_, new_n22193_, new_n22194_, new_n22195_,
    new_n22196_, new_n22197_, new_n22198_, new_n22199_, new_n22200_,
    new_n22201_, new_n22202_, new_n22203_, new_n22204_, new_n22205_,
    new_n22206_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22305_, new_n22306_, new_n22307_,
    new_n22308_, new_n22309_, new_n22310_, new_n22311_, new_n22312_,
    new_n22313_, new_n22314_, new_n22315_, new_n22316_, new_n22317_,
    new_n22318_, new_n22319_, new_n22320_, new_n22321_, new_n22322_,
    new_n22323_, new_n22324_, new_n22325_, new_n22326_, new_n22327_,
    new_n22328_, new_n22329_, new_n22330_, new_n22331_, new_n22332_,
    new_n22333_, new_n22334_, new_n22335_, new_n22336_, new_n22337_,
    new_n22338_, new_n22339_, new_n22340_, new_n22341_, new_n22342_,
    new_n22343_, new_n22344_, new_n22345_, new_n22346_, new_n22348_,
    new_n22349_, new_n22350_, new_n22351_, new_n22352_, new_n22353_,
    new_n22354_, new_n22355_, new_n22356_, new_n22357_, new_n22358_,
    new_n22359_, new_n22360_, new_n22361_, new_n22362_, new_n22363_,
    new_n22364_, new_n22365_, new_n22366_, new_n22367_, new_n22368_,
    new_n22369_, new_n22370_, new_n22371_, new_n22372_, new_n22373_,
    new_n22374_, new_n22375_, new_n22376_, new_n22377_, new_n22378_,
    new_n22379_, new_n22380_, new_n22381_, new_n22382_, new_n22383_,
    new_n22384_, new_n22385_, new_n22386_, new_n22387_, new_n22388_,
    new_n22389_, new_n22390_, new_n22391_, new_n22392_, new_n22393_,
    new_n22394_, new_n22395_, new_n22396_, new_n22397_, new_n22398_,
    new_n22399_, new_n22400_, new_n22401_, new_n22402_, new_n22403_,
    new_n22404_, new_n22405_, new_n22406_, new_n22407_, new_n22408_,
    new_n22409_, new_n22410_, new_n22411_, new_n22412_, new_n22413_,
    new_n22414_, new_n22415_, new_n22416_, new_n22417_, new_n22418_,
    new_n22419_, new_n22420_, new_n22421_, new_n22422_, new_n22423_,
    new_n22424_, new_n22425_, new_n22426_, new_n22427_, new_n22429_,
    new_n22430_, new_n22431_, new_n22432_, new_n22433_, new_n22434_,
    new_n22435_, new_n22436_, new_n22437_, new_n22438_, new_n22439_,
    new_n22440_, new_n22441_, new_n22442_, new_n22443_, new_n22444_,
    new_n22445_, new_n22446_, new_n22447_, new_n22448_, new_n22449_,
    new_n22450_, new_n22451_, new_n22452_, new_n22453_, new_n22454_,
    new_n22455_, new_n22456_, new_n22457_, new_n22458_, new_n22459_,
    new_n22460_, new_n22461_, new_n22462_, new_n22463_, new_n22464_,
    new_n22465_, new_n22466_, new_n22467_, new_n22468_, new_n22469_,
    new_n22470_, new_n22471_, new_n22472_, new_n22473_, new_n22474_,
    new_n22475_, new_n22476_, new_n22477_, new_n22478_, new_n22479_,
    new_n22480_, new_n22481_, new_n22482_, new_n22483_, new_n22484_,
    new_n22485_, new_n22486_, new_n22487_, new_n22488_, new_n22489_,
    new_n22490_, new_n22491_, new_n22492_, new_n22493_, new_n22494_,
    new_n22495_, new_n22496_, new_n22497_, new_n22498_, new_n22499_,
    new_n22500_, new_n22501_, new_n22502_, new_n22503_, new_n22504_,
    new_n22505_, new_n22506_, new_n22507_, new_n22508_, new_n22510_,
    new_n22511_, new_n22512_, new_n22513_, new_n22514_, new_n22515_,
    new_n22516_, new_n22517_, new_n22518_, new_n22519_, new_n22520_,
    new_n22521_, new_n22522_, new_n22523_, new_n22524_, new_n22525_,
    new_n22526_, new_n22527_, new_n22528_, new_n22529_, new_n22530_,
    new_n22531_, new_n22532_, new_n22533_, new_n22534_, new_n22535_,
    new_n22536_, new_n22537_, new_n22538_, new_n22539_, new_n22540_,
    new_n22541_, new_n22542_, new_n22543_, new_n22544_, new_n22545_,
    new_n22546_, new_n22547_, new_n22548_, new_n22549_, new_n22550_,
    new_n22551_, new_n22552_, new_n22553_, new_n22554_, new_n22555_,
    new_n22556_, new_n22557_, new_n22558_, new_n22559_, new_n22560_,
    new_n22561_, new_n22562_, new_n22563_, new_n22564_, new_n22565_,
    new_n22566_, new_n22567_, new_n22568_, new_n22569_, new_n22570_,
    new_n22571_, new_n22572_, new_n22573_, new_n22574_, new_n22575_,
    new_n22576_, new_n22577_, new_n22578_, new_n22579_, new_n22580_,
    new_n22581_, new_n22582_, new_n22583_, new_n22584_, new_n22585_,
    new_n22586_, new_n22587_, new_n22588_, new_n22590_, new_n22591_,
    new_n22592_, new_n22593_, new_n22594_, new_n22595_, new_n22596_,
    new_n22597_, new_n22598_, new_n22599_, new_n22600_, new_n22601_,
    new_n22602_, new_n22603_, new_n22604_, new_n22605_, new_n22606_,
    new_n22607_, new_n22608_, new_n22609_, new_n22610_, new_n22611_,
    new_n22612_, new_n22613_, new_n22614_, new_n22615_, new_n22616_,
    new_n22617_, new_n22618_, new_n22619_, new_n22620_, new_n22621_,
    new_n22622_, new_n22623_, new_n22624_, new_n22625_, new_n22626_,
    new_n22627_, new_n22628_, new_n22629_, new_n22630_, new_n22631_,
    new_n22632_, new_n22633_, new_n22634_, new_n22635_, new_n22636_,
    new_n22637_, new_n22638_, new_n22639_, new_n22640_, new_n22641_,
    new_n22642_, new_n22643_, new_n22644_, new_n22645_, new_n22646_,
    new_n22647_, new_n22648_, new_n22649_, new_n22650_, new_n22651_,
    new_n22652_, new_n22653_, new_n22654_, new_n22655_, new_n22656_,
    new_n22657_, new_n22658_, new_n22659_, new_n22660_, new_n22661_,
    new_n22662_, new_n22663_, new_n22664_, new_n22665_, new_n22666_,
    new_n22667_, new_n22668_, new_n22669_, new_n22671_, new_n22672_,
    new_n22673_, new_n22674_, new_n22675_, new_n22676_, new_n22677_,
    new_n22678_, new_n22679_, new_n22680_, new_n22681_, new_n22682_,
    new_n22683_, new_n22684_, new_n22685_, new_n22686_, new_n22687_,
    new_n22688_, new_n22689_, new_n22690_, new_n22691_, new_n22692_,
    new_n22693_, new_n22694_, new_n22695_, new_n22696_, new_n22697_,
    new_n22698_, new_n22699_, new_n22700_, new_n22701_, new_n22702_,
    new_n22703_, new_n22704_, new_n22705_, new_n22706_, new_n22707_,
    new_n22708_, new_n22709_, new_n22710_, new_n22711_, new_n22712_,
    new_n22713_, new_n22714_, new_n22715_, new_n22716_, new_n22717_,
    new_n22718_, new_n22719_, new_n22720_, new_n22721_, new_n22722_,
    new_n22723_, new_n22724_, new_n22725_, new_n22726_, new_n22727_,
    new_n22728_, new_n22729_, new_n22730_, new_n22731_, new_n22732_,
    new_n22733_, new_n22734_, new_n22735_, new_n22736_, new_n22737_,
    new_n22738_, new_n22739_, new_n22740_, new_n22741_, new_n22742_,
    new_n22743_, new_n22744_, new_n22745_, new_n22746_, new_n22747_,
    new_n22748_, new_n22749_, new_n22750_, new_n22752_, new_n22753_,
    new_n22754_, new_n22755_, new_n22756_, new_n22757_, new_n22758_,
    new_n22759_, new_n22760_, new_n22761_, new_n22762_, new_n22763_,
    new_n22764_, new_n22765_, new_n22766_, new_n22767_, new_n22768_,
    new_n22769_, new_n22770_, new_n22771_, new_n22772_, new_n22773_,
    new_n22774_, new_n22775_, new_n22776_, new_n22777_, new_n22778_,
    new_n22779_, new_n22780_, new_n22781_, new_n22782_, new_n22783_,
    new_n22784_, new_n22785_, new_n22786_, new_n22787_, new_n22788_,
    new_n22789_, new_n22790_, new_n22791_, new_n22792_, new_n22793_,
    new_n22794_, new_n22795_, new_n22796_, new_n22797_, new_n22798_,
    new_n22799_, new_n22800_, new_n22801_, new_n22802_, new_n22803_,
    new_n22804_, new_n22805_, new_n22806_, new_n22807_, new_n22808_,
    new_n22809_, new_n22810_, new_n22811_, new_n22812_, new_n22813_,
    new_n22814_, new_n22815_, new_n22816_, new_n22817_, new_n22818_,
    new_n22819_, new_n22820_, new_n22821_, new_n22822_, new_n22823_,
    new_n22824_, new_n22825_, new_n22826_, new_n22827_, new_n22828_,
    new_n22829_, new_n22830_, new_n22831_, new_n22832_, new_n22833_,
    new_n22834_, new_n22835_, new_n22836_, new_n22837_, new_n22838_,
    new_n22839_, new_n22840_, new_n22841_, new_n22842_, new_n22843_,
    new_n22844_, new_n22845_, new_n22846_, new_n22847_, new_n22848_,
    new_n22849_, new_n22850_, new_n22851_, new_n22852_, new_n22853_,
    new_n22854_, new_n22855_, new_n22856_, new_n22857_, new_n22858_,
    new_n22859_, new_n22860_, new_n22861_, new_n22862_, new_n22863_,
    new_n22864_, new_n22865_, new_n22866_, new_n22867_, new_n22868_,
    new_n22869_, new_n22870_, new_n22871_, new_n22872_, new_n22873_,
    new_n22874_, new_n22875_, new_n22876_, new_n22877_, new_n22878_,
    new_n22879_, new_n22880_, new_n22881_, new_n22882_, new_n22883_,
    new_n22884_, new_n22885_, new_n22886_, new_n22887_, new_n22888_,
    new_n22889_, new_n22890_, new_n22891_, new_n22892_, new_n22893_,
    new_n22894_, new_n22895_, new_n22896_, new_n22897_, new_n22898_,
    new_n22899_, new_n22900_, new_n22901_, new_n22902_, new_n22903_,
    new_n22904_, new_n22905_, new_n22906_, new_n22907_, new_n22908_,
    new_n22909_, new_n22910_, new_n22911_, new_n22912_, new_n22913_,
    new_n22914_, new_n22915_, new_n22916_, new_n22917_, new_n22918_,
    new_n22919_, new_n22920_, new_n22921_, new_n22922_, new_n22923_,
    new_n22924_, new_n22925_, new_n22926_, new_n22927_, new_n22928_,
    new_n22929_, new_n22930_, new_n22931_, new_n22932_, new_n22933_,
    new_n22934_, new_n22935_, new_n22936_, new_n22937_, new_n22938_,
    new_n22939_, new_n22940_, new_n22941_, new_n22942_, new_n22943_,
    new_n22944_, new_n22945_, new_n22946_, new_n22947_, new_n22948_,
    new_n22949_, new_n22950_, new_n22951_, new_n22952_, new_n22953_,
    new_n22954_, new_n22955_, new_n22956_, new_n22957_, new_n22958_,
    new_n22959_, new_n22960_, new_n22961_, new_n22962_, new_n22963_,
    new_n22964_, new_n22965_, new_n22966_, new_n22967_, new_n22968_,
    new_n22969_, new_n22970_, new_n22971_, new_n22972_, new_n22973_,
    new_n22974_, new_n22975_, new_n22976_, new_n22977_, new_n22978_,
    new_n22979_, new_n22980_, new_n22981_, new_n22982_, new_n22983_,
    new_n22984_, new_n22985_, new_n22986_, new_n22987_, new_n22988_,
    new_n22989_, new_n22990_, new_n22991_, new_n22992_, new_n22993_,
    new_n22994_, new_n22995_, new_n22996_, new_n22997_, new_n22998_,
    new_n22999_, new_n23000_, new_n23001_, new_n23002_, new_n23003_,
    new_n23004_, new_n23005_, new_n23006_, new_n23007_, new_n23008_,
    new_n23009_, new_n23010_, new_n23011_, new_n23012_, new_n23013_,
    new_n23014_, new_n23015_, new_n23016_, new_n23017_, new_n23018_,
    new_n23019_, new_n23020_, new_n23021_, new_n23022_, new_n23023_,
    new_n23024_, new_n23025_, new_n23026_, new_n23027_, new_n23028_,
    new_n23029_, new_n23030_, new_n23031_, new_n23032_, new_n23033_,
    new_n23034_, new_n23035_, new_n23036_, new_n23037_, new_n23038_,
    new_n23039_, new_n23040_, new_n23041_, new_n23042_, new_n23043_,
    new_n23044_, new_n23045_, new_n23046_, new_n23047_, new_n23048_,
    new_n23049_, new_n23050_, new_n23051_, new_n23052_, new_n23053_,
    new_n23054_, new_n23055_, new_n23056_, new_n23057_, new_n23058_,
    new_n23059_, new_n23060_, new_n23061_, new_n23062_, new_n23063_,
    new_n23064_, new_n23065_, new_n23066_, new_n23067_, new_n23068_,
    new_n23069_, new_n23070_, new_n23071_, new_n23072_, new_n23073_,
    new_n23074_, new_n23075_, new_n23076_, new_n23077_, new_n23078_,
    new_n23079_, new_n23080_, new_n23081_, new_n23082_, new_n23083_,
    new_n23084_, new_n23085_, new_n23086_, new_n23087_, new_n23088_,
    new_n23089_, new_n23090_, new_n23091_, new_n23092_, new_n23093_,
    new_n23094_, new_n23095_, new_n23096_, new_n23097_, new_n23098_,
    new_n23099_, new_n23100_, new_n23101_, new_n23102_, new_n23103_,
    new_n23104_, new_n23105_, new_n23106_, new_n23107_, new_n23108_,
    new_n23109_, new_n23110_, new_n23111_, new_n23112_, new_n23113_,
    new_n23114_, new_n23115_, new_n23116_, new_n23117_, new_n23118_,
    new_n23119_, new_n23120_, new_n23121_, new_n23122_, new_n23123_,
    new_n23124_, new_n23125_, new_n23126_, new_n23127_, new_n23128_,
    new_n23129_, new_n23130_, new_n23131_, new_n23132_, new_n23133_,
    new_n23134_, new_n23135_, new_n23136_, new_n23137_, new_n23138_,
    new_n23139_, new_n23140_, new_n23141_, new_n23142_, new_n23143_,
    new_n23144_, new_n23145_, new_n23146_, new_n23147_, new_n23148_,
    new_n23149_, new_n23150_, new_n23151_, new_n23152_, new_n23153_,
    new_n23154_, new_n23155_, new_n23156_, new_n23157_, new_n23158_,
    new_n23159_, new_n23160_, new_n23161_, new_n23162_, new_n23163_,
    new_n23164_, new_n23165_, new_n23166_, new_n23167_, new_n23168_,
    new_n23169_, new_n23170_, new_n23171_, new_n23172_, new_n23173_,
    new_n23174_, new_n23175_, new_n23176_, new_n23177_, new_n23178_,
    new_n23179_, new_n23180_, new_n23181_, new_n23182_, new_n23183_,
    new_n23184_, new_n23185_, new_n23186_, new_n23187_, new_n23188_,
    new_n23189_, new_n23190_, new_n23191_, new_n23192_, new_n23193_,
    new_n23194_, new_n23195_, new_n23196_, new_n23197_, new_n23198_,
    new_n23199_, new_n23200_, new_n23201_, new_n23202_, new_n23203_,
    new_n23204_, new_n23205_, new_n23206_, new_n23207_, new_n23208_,
    new_n23209_, new_n23210_, new_n23211_, new_n23212_, new_n23213_,
    new_n23214_, new_n23215_, new_n23216_, new_n23217_, new_n23218_,
    new_n23219_, new_n23220_, new_n23221_, new_n23222_, new_n23223_,
    new_n23224_, new_n23225_, new_n23227_, new_n23228_, new_n23229_,
    new_n23230_, new_n23231_, new_n23232_, new_n23233_, new_n23234_,
    new_n23235_, new_n23236_, new_n23237_, new_n23238_, new_n23239_,
    new_n23240_, new_n23241_, new_n23242_, new_n23243_, new_n23244_,
    new_n23245_, new_n23246_, new_n23247_, new_n23248_, new_n23249_,
    new_n23250_, new_n23251_, new_n23252_, new_n23253_, new_n23254_,
    new_n23255_, new_n23256_, new_n23257_, new_n23258_, new_n23259_,
    new_n23260_, new_n23261_, new_n23262_, new_n23263_, new_n23264_,
    new_n23265_, new_n23266_, new_n23267_, new_n23268_, new_n23269_,
    new_n23270_, new_n23271_, new_n23272_, new_n23273_, new_n23274_,
    new_n23275_, new_n23276_, new_n23277_, new_n23278_, new_n23279_,
    new_n23280_, new_n23281_, new_n23282_, new_n23283_, new_n23284_,
    new_n23285_, new_n23286_, new_n23287_, new_n23288_, new_n23289_,
    new_n23290_, new_n23291_, new_n23292_, new_n23293_, new_n23294_,
    new_n23295_, new_n23296_, new_n23297_, new_n23298_, new_n23299_,
    new_n23300_, new_n23301_, new_n23302_, new_n23303_, new_n23304_,
    new_n23305_, new_n23306_, new_n23307_, new_n23308_, new_n23309_,
    new_n23310_, new_n23311_, new_n23312_, new_n23313_, new_n23314_,
    new_n23315_, new_n23316_, new_n23317_, new_n23318_, new_n23319_,
    new_n23320_, new_n23321_, new_n23322_, new_n23323_, new_n23324_,
    new_n23325_, new_n23326_, new_n23327_, new_n23328_, new_n23329_,
    new_n23330_, new_n23331_, new_n23332_, new_n23333_, new_n23334_,
    new_n23335_, new_n23336_, new_n23337_, new_n23338_, new_n23339_,
    new_n23340_, new_n23341_, new_n23342_, new_n23343_, new_n23344_,
    new_n23345_, new_n23346_, new_n23347_, new_n23348_, new_n23349_,
    new_n23350_, new_n23351_, new_n23352_, new_n23353_, new_n23354_,
    new_n23355_, new_n23356_, new_n23357_, new_n23358_, new_n23359_,
    new_n23360_, new_n23361_, new_n23362_, new_n23363_, new_n23364_,
    new_n23365_, new_n23366_, new_n23367_, new_n23368_, new_n23369_,
    new_n23370_, new_n23371_, new_n23372_, new_n23373_, new_n23374_,
    new_n23375_, new_n23376_, new_n23377_, new_n23378_, new_n23379_,
    new_n23380_, new_n23381_, new_n23382_, new_n23383_, new_n23384_,
    new_n23385_, new_n23386_, new_n23387_, new_n23388_, new_n23389_,
    new_n23390_, new_n23391_, new_n23392_, new_n23393_, new_n23394_,
    new_n23395_, new_n23396_, new_n23397_, new_n23398_, new_n23399_,
    new_n23400_, new_n23401_, new_n23402_, new_n23403_, new_n23404_,
    new_n23405_, new_n23406_, new_n23407_, new_n23408_, new_n23409_,
    new_n23410_, new_n23411_, new_n23412_, new_n23413_, new_n23414_,
    new_n23415_, new_n23416_, new_n23417_, new_n23418_, new_n23419_,
    new_n23420_, new_n23421_, new_n23422_, new_n23423_, new_n23424_,
    new_n23425_, new_n23426_, new_n23427_, new_n23428_, new_n23429_,
    new_n23430_, new_n23431_, new_n23432_, new_n23433_, new_n23434_,
    new_n23435_, new_n23436_, new_n23437_, new_n23438_, new_n23439_,
    new_n23440_, new_n23441_, new_n23442_, new_n23443_, new_n23444_,
    new_n23445_, new_n23446_, new_n23447_, new_n23448_, new_n23449_,
    new_n23450_, new_n23451_, new_n23452_, new_n23453_, new_n23454_,
    new_n23455_, new_n23456_, new_n23457_, new_n23458_, new_n23459_,
    new_n23460_, new_n23461_, new_n23462_, new_n23463_, new_n23464_,
    new_n23465_, new_n23466_, new_n23467_, new_n23468_, new_n23469_,
    new_n23470_, new_n23471_, new_n23472_, new_n23473_, new_n23474_,
    new_n23475_, new_n23476_, new_n23477_, new_n23478_, new_n23479_,
    new_n23480_, new_n23481_, new_n23482_, new_n23483_, new_n23484_,
    new_n23485_, new_n23486_, new_n23487_, new_n23488_, new_n23489_,
    new_n23490_, new_n23491_, new_n23492_, new_n23493_, new_n23494_,
    new_n23495_, new_n23496_, new_n23497_, new_n23498_, new_n23499_,
    new_n23500_, new_n23501_, new_n23502_, new_n23503_, new_n23504_,
    new_n23505_, new_n23506_, new_n23507_, new_n23508_, new_n23509_,
    new_n23510_, new_n23511_, new_n23512_, new_n23513_, new_n23514_,
    new_n23515_, new_n23516_, new_n23517_, new_n23518_, new_n23519_,
    new_n23520_, new_n23521_, new_n23522_, new_n23523_, new_n23524_,
    new_n23525_, new_n23526_, new_n23527_, new_n23528_, new_n23529_,
    new_n23530_, new_n23531_, new_n23532_, new_n23533_, new_n23534_,
    new_n23535_, new_n23536_, new_n23537_, new_n23538_, new_n23539_,
    new_n23540_, new_n23541_, new_n23542_, new_n23543_, new_n23544_,
    new_n23545_, new_n23546_, new_n23547_, new_n23548_, new_n23549_,
    new_n23550_, new_n23551_, new_n23552_, new_n23553_, new_n23554_,
    new_n23555_, new_n23556_, new_n23557_, new_n23558_, new_n23559_,
    new_n23560_, new_n23561_, new_n23562_, new_n23563_, new_n23564_,
    new_n23565_, new_n23566_, new_n23567_, new_n23568_, new_n23569_,
    new_n23570_, new_n23571_, new_n23572_, new_n23573_, new_n23574_,
    new_n23575_, new_n23576_, new_n23577_, new_n23578_, new_n23579_,
    new_n23580_, new_n23581_, new_n23582_, new_n23583_, new_n23584_,
    new_n23585_, new_n23586_, new_n23587_, new_n23588_, new_n23589_,
    new_n23590_, new_n23591_, new_n23592_, new_n23593_, new_n23594_,
    new_n23595_, new_n23596_, new_n23597_, new_n23598_, new_n23599_,
    new_n23600_, new_n23601_, new_n23602_, new_n23603_, new_n23604_,
    new_n23605_, new_n23606_, new_n23607_, new_n23608_, new_n23609_,
    new_n23610_, new_n23611_, new_n23612_, new_n23613_, new_n23614_,
    new_n23615_, new_n23616_, new_n23617_, new_n23618_, new_n23619_,
    new_n23620_, new_n23621_, new_n23622_, new_n23623_, new_n23624_,
    new_n23625_, new_n23626_, new_n23627_, new_n23628_, new_n23629_,
    new_n23630_, new_n23631_, new_n23632_, new_n23633_, new_n23634_,
    new_n23635_, new_n23636_, new_n23637_, new_n23638_, new_n23639_,
    new_n23640_, new_n23641_, new_n23642_, new_n23643_, new_n23644_,
    new_n23645_, new_n23646_, new_n23647_, new_n23648_, new_n23649_,
    new_n23650_, new_n23651_, new_n23652_, new_n23653_, new_n23654_,
    new_n23655_, new_n23656_, new_n23657_, new_n23658_, new_n23659_,
    new_n23660_, new_n23661_, new_n23662_, new_n23663_, new_n23664_,
    new_n23665_, new_n23666_, new_n23667_, new_n23668_, new_n23669_,
    new_n23670_, new_n23671_, new_n23672_, new_n23673_, new_n23674_,
    new_n23675_, new_n23676_, new_n23677_, new_n23678_, new_n23679_,
    new_n23680_, new_n23681_, new_n23682_, new_n23683_, new_n23684_,
    new_n23685_, new_n23686_, new_n23687_, new_n23688_, new_n23689_,
    new_n23690_, new_n23691_, new_n23692_, new_n23693_, new_n23694_,
    new_n23695_, new_n23696_, new_n23697_, new_n23698_, new_n23699_,
    new_n23700_, new_n23701_, new_n23702_, new_n23703_, new_n23704_,
    new_n23705_, new_n23706_, new_n23707_, new_n23708_, new_n23709_,
    new_n23711_, new_n23712_, new_n23713_, new_n23714_, new_n23715_,
    new_n23716_, new_n23717_, new_n23718_, new_n23719_, new_n23720_,
    new_n23721_, new_n23722_, new_n23723_, new_n23724_, new_n23725_,
    new_n23726_, new_n23727_, new_n23728_, new_n23729_, new_n23730_,
    new_n23731_, new_n23732_, new_n23733_, new_n23734_, new_n23735_,
    new_n23736_, new_n23737_, new_n23738_, new_n23739_, new_n23740_,
    new_n23741_, new_n23742_, new_n23743_, new_n23744_, new_n23745_,
    new_n23746_, new_n23747_, new_n23748_, new_n23749_, new_n23750_,
    new_n23751_, new_n23752_, new_n23753_, new_n23754_, new_n23755_,
    new_n23756_, new_n23757_, new_n23758_, new_n23759_, new_n23760_,
    new_n23761_, new_n23762_, new_n23763_, new_n23764_, new_n23765_,
    new_n23766_, new_n23767_, new_n23768_, new_n23769_, new_n23770_,
    new_n23771_, new_n23772_, new_n23773_, new_n23774_, new_n23775_,
    new_n23776_, new_n23777_, new_n23778_, new_n23779_, new_n23780_,
    new_n23781_, new_n23782_, new_n23783_, new_n23784_, new_n23785_,
    new_n23786_, new_n23787_, new_n23788_, new_n23789_, new_n23790_,
    new_n23791_, new_n23792_, new_n23793_, new_n23794_, new_n23795_,
    new_n23796_, new_n23797_, new_n23798_, new_n23799_, new_n23800_,
    new_n23801_, new_n23802_, new_n23803_, new_n23804_, new_n23805_,
    new_n23806_, new_n23807_, new_n23808_, new_n23809_, new_n23810_,
    new_n23811_, new_n23812_, new_n23813_, new_n23814_, new_n23815_,
    new_n23816_, new_n23817_, new_n23818_, new_n23819_, new_n23820_,
    new_n23821_, new_n23822_, new_n23823_, new_n23824_, new_n23825_,
    new_n23826_, new_n23827_, new_n23828_, new_n23829_, new_n23830_,
    new_n23831_, new_n23832_, new_n23833_, new_n23834_, new_n23835_,
    new_n23836_, new_n23837_, new_n23838_, new_n23839_, new_n23840_,
    new_n23841_, new_n23842_, new_n23843_, new_n23844_, new_n23845_,
    new_n23846_, new_n23847_, new_n23848_, new_n23849_, new_n23850_,
    new_n23851_, new_n23852_, new_n23853_, new_n23854_, new_n23855_,
    new_n23856_, new_n23857_, new_n23858_, new_n23859_, new_n23860_,
    new_n23861_, new_n23862_, new_n23863_, new_n23864_, new_n23865_,
    new_n23866_, new_n23867_, new_n23868_, new_n23869_, new_n23870_,
    new_n23871_, new_n23872_, new_n23873_, new_n23874_, new_n23875_,
    new_n23876_, new_n23877_, new_n23878_, new_n23879_, new_n23880_,
    new_n23881_, new_n23882_, new_n23883_, new_n23884_, new_n23885_,
    new_n23886_, new_n23887_, new_n23888_, new_n23889_, new_n23890_,
    new_n23891_, new_n23892_, new_n23893_, new_n23894_, new_n23895_,
    new_n23896_, new_n23897_, new_n23898_, new_n23899_, new_n23900_,
    new_n23901_, new_n23902_, new_n23903_, new_n23904_, new_n23905_,
    new_n23906_, new_n23907_, new_n23908_, new_n23909_, new_n23910_,
    new_n23911_, new_n23912_, new_n23913_, new_n23914_, new_n23915_,
    new_n23916_, new_n23917_, new_n23918_, new_n23919_, new_n23920_,
    new_n23921_, new_n23922_, new_n23923_, new_n23924_, new_n23925_,
    new_n23926_, new_n23927_, new_n23928_, new_n23929_, new_n23930_,
    new_n23931_, new_n23932_, new_n23933_, new_n23934_, new_n23935_,
    new_n23936_, new_n23937_, new_n23938_, new_n23939_, new_n23940_,
    new_n23941_, new_n23942_, new_n23943_, new_n23944_, new_n23945_,
    new_n23946_, new_n23947_, new_n23948_, new_n23949_, new_n23950_,
    new_n23951_, new_n23952_, new_n23953_, new_n23954_, new_n23955_,
    new_n23956_, new_n23957_, new_n23958_, new_n23959_, new_n23960_,
    new_n23961_, new_n23962_, new_n23963_, new_n23964_, new_n23965_,
    new_n23966_, new_n23967_, new_n23968_, new_n23969_, new_n23970_,
    new_n23971_, new_n23972_, new_n23973_, new_n23974_, new_n23975_,
    new_n23976_, new_n23977_, new_n23978_, new_n23979_, new_n23980_,
    new_n23981_, new_n23982_, new_n23983_, new_n23984_, new_n23985_,
    new_n23986_, new_n23987_, new_n23988_, new_n23989_, new_n23990_,
    new_n23991_, new_n23992_, new_n23993_, new_n23994_, new_n23995_,
    new_n23996_, new_n23997_, new_n23998_, new_n23999_, new_n24000_,
    new_n24001_, new_n24002_, new_n24003_, new_n24004_, new_n24005_,
    new_n24006_, new_n24007_, new_n24008_, new_n24009_, new_n24010_,
    new_n24011_, new_n24012_, new_n24013_, new_n24014_, new_n24015_,
    new_n24016_, new_n24017_, new_n24018_, new_n24019_, new_n24020_,
    new_n24021_, new_n24022_, new_n24023_, new_n24024_, new_n24025_,
    new_n24026_, new_n24027_, new_n24028_, new_n24029_, new_n24030_,
    new_n24031_, new_n24032_, new_n24033_, new_n24034_, new_n24035_,
    new_n24036_, new_n24037_, new_n24038_, new_n24039_, new_n24040_,
    new_n24041_, new_n24042_, new_n24043_, new_n24044_, new_n24045_,
    new_n24046_, new_n24047_, new_n24048_, new_n24049_, new_n24050_,
    new_n24051_, new_n24052_, new_n24053_, new_n24054_, new_n24055_,
    new_n24056_, new_n24057_, new_n24058_, new_n24059_, new_n24060_,
    new_n24061_, new_n24062_, new_n24063_, new_n24064_, new_n24065_,
    new_n24066_, new_n24067_, new_n24068_, new_n24069_, new_n24070_,
    new_n24071_, new_n24072_, new_n24073_, new_n24074_, new_n24075_,
    new_n24076_, new_n24077_, new_n24078_, new_n24079_, new_n24080_,
    new_n24081_, new_n24082_, new_n24083_, new_n24084_, new_n24085_,
    new_n24086_, new_n24087_, new_n24088_, new_n24089_, new_n24090_,
    new_n24091_, new_n24092_, new_n24093_, new_n24094_, new_n24095_,
    new_n24096_, new_n24097_, new_n24098_, new_n24099_, new_n24100_,
    new_n24101_, new_n24102_, new_n24103_, new_n24104_, new_n24105_,
    new_n24106_, new_n24107_, new_n24108_, new_n24109_, new_n24110_,
    new_n24111_, new_n24112_, new_n24113_, new_n24114_, new_n24115_,
    new_n24116_, new_n24117_, new_n24118_, new_n24119_, new_n24120_,
    new_n24121_, new_n24122_, new_n24123_, new_n24124_, new_n24125_,
    new_n24126_, new_n24127_, new_n24128_, new_n24129_, new_n24130_,
    new_n24131_, new_n24132_, new_n24133_, new_n24134_, new_n24135_,
    new_n24136_, new_n24137_, new_n24138_, new_n24139_, new_n24140_,
    new_n24141_, new_n24142_, new_n24143_, new_n24144_, new_n24145_,
    new_n24146_, new_n24147_, new_n24148_, new_n24149_, new_n24150_,
    new_n24151_, new_n24152_, new_n24153_, new_n24154_, new_n24155_,
    new_n24156_, new_n24157_, new_n24158_, new_n24159_, new_n24160_,
    new_n24161_, new_n24162_, new_n24163_, new_n24164_, new_n24165_,
    new_n24166_, new_n24167_, new_n24168_, new_n24169_, new_n24170_,
    new_n24171_, new_n24172_, new_n24173_, new_n24174_, new_n24175_,
    new_n24176_, new_n24177_, new_n24178_, new_n24179_, new_n24180_,
    new_n24181_, new_n24182_, new_n24183_, new_n24184_, new_n24185_,
    new_n24186_, new_n24187_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24240_, new_n24241_,
    new_n24242_, new_n24243_, new_n24244_, new_n24245_, new_n24246_,
    new_n24247_, new_n24248_, new_n24249_, new_n24250_, new_n24251_,
    new_n24252_, new_n24253_, new_n24254_, new_n24255_, new_n24256_,
    new_n24257_, new_n24258_, new_n24259_, new_n24260_, new_n24261_,
    new_n24262_, new_n24263_, new_n24264_, new_n24265_, new_n24266_,
    new_n24267_, new_n24268_, new_n24269_, new_n24270_, new_n24271_,
    new_n24272_, new_n24273_, new_n24274_, new_n24275_, new_n24276_,
    new_n24277_, new_n24278_, new_n24279_, new_n24280_, new_n24281_,
    new_n24282_, new_n24283_, new_n24284_, new_n24285_, new_n24286_,
    new_n24287_, new_n24288_, new_n24289_, new_n24290_, new_n24291_,
    new_n24292_, new_n24293_, new_n24294_, new_n24295_, new_n24296_,
    new_n24297_, new_n24298_, new_n24299_, new_n24300_, new_n24301_,
    new_n24302_, new_n24303_, new_n24304_, new_n24305_, new_n24306_,
    new_n24307_, new_n24308_, new_n24309_, new_n24310_, new_n24311_,
    new_n24312_, new_n24313_, new_n24314_, new_n24315_, new_n24316_,
    new_n24317_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24336_,
    new_n24337_, new_n24338_, new_n24339_, new_n24340_, new_n24341_,
    new_n24342_, new_n24343_, new_n24344_, new_n24345_, new_n24346_,
    new_n24347_, new_n24348_, new_n24349_, new_n24350_, new_n24351_,
    new_n24352_, new_n24353_, new_n24354_, new_n24355_, new_n24356_,
    new_n24357_, new_n24358_, new_n24359_, new_n24360_, new_n24361_,
    new_n24362_, new_n24363_, new_n24364_, new_n24365_, new_n24366_,
    new_n24367_, new_n24368_, new_n24369_, new_n24370_, new_n24371_,
    new_n24372_, new_n24373_, new_n24374_, new_n24375_, new_n24376_,
    new_n24377_, new_n24378_, new_n24379_, new_n24380_, new_n24381_,
    new_n24382_, new_n24383_, new_n24384_, new_n24385_, new_n24386_,
    new_n24387_, new_n24388_, new_n24389_, new_n24390_, new_n24391_,
    new_n24392_, new_n24393_, new_n24394_, new_n24395_, new_n24396_,
    new_n24397_, new_n24398_, new_n24399_, new_n24400_, new_n24401_,
    new_n24402_, new_n24403_, new_n24404_, new_n24405_, new_n24406_,
    new_n24407_, new_n24408_, new_n24409_, new_n24410_, new_n24411_,
    new_n24412_, new_n24413_, new_n24414_, new_n24415_, new_n24416_,
    new_n24417_, new_n24418_, new_n24419_, new_n24420_, new_n24421_,
    new_n24422_, new_n24423_, new_n24424_, new_n24425_, new_n24426_,
    new_n24427_, new_n24428_, new_n24429_, new_n24430_, new_n24431_,
    new_n24432_, new_n24433_, new_n24434_, new_n24435_, new_n24436_,
    new_n24437_, new_n24438_, new_n24439_, new_n24440_, new_n24441_,
    new_n24442_, new_n24443_, new_n24444_, new_n24445_, new_n24446_,
    new_n24447_, new_n24448_, new_n24449_, new_n24450_, new_n24451_,
    new_n24452_, new_n24453_, new_n24454_, new_n24455_, new_n24456_,
    new_n24457_, new_n24458_, new_n24459_, new_n24460_, new_n24461_,
    new_n24462_, new_n24463_, new_n24464_, new_n24465_, new_n24466_,
    new_n24467_, new_n24468_, new_n24469_, new_n24470_, new_n24471_,
    new_n24472_, new_n24473_, new_n24474_, new_n24475_, new_n24476_,
    new_n24477_, new_n24478_, new_n24479_, new_n24480_, new_n24481_,
    new_n24482_, new_n24483_, new_n24484_, new_n24485_, new_n24486_,
    new_n24487_, new_n24488_, new_n24489_, new_n24490_, new_n24491_,
    new_n24492_, new_n24493_, new_n24494_, new_n24495_, new_n24496_,
    new_n24497_, new_n24498_, new_n24499_, new_n24500_, new_n24501_,
    new_n24502_, new_n24503_, new_n24504_, new_n24505_, new_n24506_,
    new_n24507_, new_n24508_, new_n24509_, new_n24510_, new_n24511_,
    new_n24512_, new_n24513_, new_n24514_, new_n24515_, new_n24516_,
    new_n24517_, new_n24518_, new_n24519_, new_n24520_, new_n24521_,
    new_n24522_, new_n24523_, new_n24524_, new_n24525_, new_n24526_,
    new_n24527_, new_n24528_, new_n24529_, new_n24530_, new_n24531_,
    new_n24532_, new_n24533_, new_n24534_, new_n24535_, new_n24536_,
    new_n24537_, new_n24538_, new_n24539_, new_n24540_, new_n24541_,
    new_n24542_, new_n24543_, new_n24544_, new_n24545_, new_n24546_,
    new_n24547_, new_n24548_, new_n24549_, new_n24550_, new_n24551_,
    new_n24552_, new_n24553_, new_n24554_, new_n24555_, new_n24556_,
    new_n24557_, new_n24558_, new_n24559_, new_n24560_, new_n24561_,
    new_n24562_, new_n24563_, new_n24564_, new_n24565_, new_n24566_,
    new_n24567_, new_n24568_, new_n24569_, new_n24570_, new_n24571_,
    new_n24572_, new_n24573_, new_n24574_, new_n24575_, new_n24576_,
    new_n24577_, new_n24578_, new_n24579_, new_n24580_, new_n24581_,
    new_n24582_, new_n24583_, new_n24584_, new_n24585_, new_n24586_,
    new_n24587_, new_n24588_, new_n24589_, new_n24590_, new_n24591_,
    new_n24592_, new_n24593_, new_n24594_, new_n24595_, new_n24596_,
    new_n24597_, new_n24598_, new_n24599_, new_n24600_, new_n24601_,
    new_n24602_, new_n24603_, new_n24604_, new_n24605_, new_n24606_,
    new_n24607_, new_n24608_, new_n24609_, new_n24610_, new_n24611_,
    new_n24612_, new_n24613_, new_n24614_, new_n24615_, new_n24616_,
    new_n24617_, new_n24618_, new_n24619_, new_n24620_, new_n24621_,
    new_n24622_, new_n24623_, new_n24624_, new_n24625_, new_n24626_,
    new_n24627_, new_n24628_, new_n24629_, new_n24630_, new_n24631_,
    new_n24632_, new_n24633_, new_n24634_, new_n24635_, new_n24636_,
    new_n24637_, new_n24639_, new_n24640_, new_n24641_, new_n24642_,
    new_n24643_, new_n24644_, new_n24645_, new_n24646_, new_n24647_,
    new_n24648_, new_n24649_, new_n24650_, new_n24651_, new_n24652_,
    new_n24653_, new_n24654_, new_n24655_, new_n24656_, new_n24657_,
    new_n24658_, new_n24659_, new_n24660_, new_n24661_, new_n24662_,
    new_n24663_, new_n24664_, new_n24665_, new_n24666_, new_n24667_,
    new_n24668_, new_n24669_, new_n24670_, new_n24671_, new_n24672_,
    new_n24673_, new_n24674_, new_n24675_, new_n24676_, new_n24677_,
    new_n24678_, new_n24679_, new_n24680_, new_n24681_, new_n24682_,
    new_n24683_, new_n24684_, new_n24685_, new_n24686_, new_n24687_,
    new_n24688_, new_n24689_, new_n24690_, new_n24691_, new_n24692_,
    new_n24693_, new_n24694_, new_n24695_, new_n24696_, new_n24697_,
    new_n24698_, new_n24699_, new_n24700_, new_n24701_, new_n24702_,
    new_n24703_, new_n24704_, new_n24705_, new_n24706_, new_n24707_,
    new_n24708_, new_n24709_, new_n24710_, new_n24711_, new_n24712_,
    new_n24713_, new_n24714_, new_n24715_, new_n24716_, new_n24717_,
    new_n24718_, new_n24719_, new_n24720_, new_n24721_, new_n24722_,
    new_n24723_, new_n24724_, new_n24725_, new_n24726_, new_n24727_,
    new_n24728_, new_n24729_, new_n24730_, new_n24731_, new_n24732_,
    new_n24733_, new_n24734_, new_n24735_, new_n24736_, new_n24737_,
    new_n24738_, new_n24739_, new_n24740_, new_n24741_, new_n24742_,
    new_n24743_, new_n24744_, new_n24745_, new_n24746_, new_n24747_,
    new_n24748_, new_n24749_, new_n24750_, new_n24751_, new_n24752_,
    new_n24753_, new_n24754_, new_n24755_, new_n24756_, new_n24757_,
    new_n24758_, new_n24759_, new_n24760_, new_n24761_, new_n24762_,
    new_n24763_, new_n24764_, new_n24765_, new_n24766_, new_n24767_,
    new_n24768_, new_n24769_, new_n24770_, new_n24771_, new_n24772_,
    new_n24773_, new_n24774_, new_n24775_, new_n24776_, new_n24777_,
    new_n24778_, new_n24779_, new_n24780_, new_n24781_, new_n24782_,
    new_n24783_, new_n24784_, new_n24785_, new_n24786_, new_n24787_,
    new_n24788_, new_n24789_, new_n24790_, new_n24791_, new_n24792_,
    new_n24793_, new_n24794_, new_n24795_, new_n24796_, new_n24797_,
    new_n24798_, new_n24799_, new_n24800_, new_n24801_, new_n24802_,
    new_n24803_, new_n24804_, new_n24805_, new_n24806_, new_n24807_,
    new_n24808_, new_n24809_, new_n24810_, new_n24811_, new_n24812_,
    new_n24813_, new_n24814_, new_n24815_, new_n24816_, new_n24817_,
    new_n24818_, new_n24819_, new_n24820_, new_n24821_, new_n24822_,
    new_n24823_, new_n24824_, new_n24825_, new_n24826_, new_n24827_,
    new_n24828_, new_n24829_, new_n24830_, new_n24831_, new_n24832_,
    new_n24833_, new_n24834_, new_n24835_, new_n24836_, new_n24837_,
    new_n24838_, new_n24839_, new_n24840_, new_n24841_, new_n24842_,
    new_n24843_, new_n24844_, new_n24845_, new_n24846_, new_n24847_,
    new_n24848_, new_n24849_, new_n24850_, new_n24851_, new_n24852_,
    new_n24853_, new_n24854_, new_n24855_, new_n24856_, new_n24857_,
    new_n24858_, new_n24859_, new_n24860_, new_n24861_, new_n24862_,
    new_n24863_, new_n24864_, new_n24865_, new_n24866_, new_n24867_,
    new_n24868_, new_n24869_, new_n24870_, new_n24871_, new_n24872_,
    new_n24873_, new_n24874_, new_n24875_, new_n24876_, new_n24877_,
    new_n24878_, new_n24879_, new_n24880_, new_n24881_, new_n24882_,
    new_n24883_, new_n24884_, new_n24885_, new_n24886_, new_n24887_,
    new_n24888_, new_n24889_, new_n24890_, new_n24891_, new_n24892_,
    new_n24893_, new_n24894_, new_n24895_, new_n24896_, new_n24897_,
    new_n24898_, new_n24899_, new_n24900_, new_n24901_, new_n24902_,
    new_n24903_, new_n24904_, new_n24905_, new_n24906_, new_n24907_,
    new_n24908_, new_n24909_, new_n24910_, new_n24911_, new_n24912_,
    new_n24913_, new_n24914_, new_n24915_, new_n24916_, new_n24917_,
    new_n24918_, new_n24919_, new_n24920_, new_n24921_, new_n24922_,
    new_n24923_, new_n24924_, new_n24925_, new_n24926_, new_n24927_,
    new_n24928_, new_n24929_, new_n24930_, new_n24931_, new_n24932_,
    new_n24933_, new_n24934_, new_n24935_, new_n24936_, new_n24937_,
    new_n24938_, new_n24939_, new_n24940_, new_n24941_, new_n24942_,
    new_n24943_, new_n24944_, new_n24945_, new_n24946_, new_n24947_,
    new_n24948_, new_n24949_, new_n24950_, new_n24951_, new_n24952_,
    new_n24953_, new_n24954_, new_n24955_, new_n24956_, new_n24957_,
    new_n24958_, new_n24959_, new_n24960_, new_n24961_, new_n24962_,
    new_n24963_, new_n24964_, new_n24965_, new_n24966_, new_n24967_,
    new_n24968_, new_n24969_, new_n24970_, new_n24971_, new_n24972_,
    new_n24973_, new_n24974_, new_n24975_, new_n24976_, new_n24977_,
    new_n24978_, new_n24979_, new_n24980_, new_n24981_, new_n24982_,
    new_n24983_, new_n24984_, new_n24985_, new_n24986_, new_n24987_,
    new_n24988_, new_n24989_, new_n24990_, new_n24991_, new_n24992_,
    new_n24993_, new_n24994_, new_n24995_, new_n24996_, new_n24997_,
    new_n24998_, new_n24999_, new_n25000_, new_n25001_, new_n25002_,
    new_n25003_, new_n25004_, new_n25005_, new_n25006_, new_n25007_,
    new_n25008_, new_n25009_, new_n25010_, new_n25011_, new_n25012_,
    new_n25013_, new_n25014_, new_n25015_, new_n25016_, new_n25017_,
    new_n25018_, new_n25019_, new_n25020_, new_n25021_, new_n25022_,
    new_n25023_, new_n25024_, new_n25025_, new_n25026_, new_n25027_,
    new_n25028_, new_n25029_, new_n25030_, new_n25031_, new_n25032_,
    new_n25033_, new_n25034_, new_n25035_, new_n25036_, new_n25037_,
    new_n25038_, new_n25039_, new_n25040_, new_n25041_, new_n25042_,
    new_n25043_, new_n25044_, new_n25045_, new_n25046_, new_n25047_,
    new_n25048_, new_n25049_, new_n25050_, new_n25051_, new_n25052_,
    new_n25053_, new_n25054_, new_n25055_, new_n25056_, new_n25057_,
    new_n25058_, new_n25059_, new_n25060_, new_n25061_, new_n25062_,
    new_n25063_, new_n25064_, new_n25065_, new_n25066_, new_n25067_,
    new_n25068_, new_n25069_, new_n25070_, new_n25071_, new_n25072_,
    new_n25073_, new_n25074_, new_n25075_, new_n25076_, new_n25077_,
    new_n25078_, new_n25079_, new_n25080_, new_n25081_, new_n25082_,
    new_n25083_, new_n25084_, new_n25085_, new_n25086_, new_n25087_,
    new_n25088_, new_n25089_, new_n25090_, new_n25091_, new_n25092_,
    new_n25093_, new_n25094_, new_n25095_, new_n25096_, new_n25097_,
    new_n25098_, new_n25099_, new_n25100_, new_n25101_, new_n25102_,
    new_n25103_, new_n25104_, new_n25105_, new_n25106_, new_n25107_,
    new_n25108_, new_n25109_, new_n25110_, new_n25111_, new_n25112_,
    new_n25113_, new_n25114_, new_n25115_, new_n25116_, new_n25117_,
    new_n25118_, new_n25119_, new_n25120_, new_n25121_, new_n25123_,
    new_n25124_, new_n25125_, new_n25126_, new_n25127_, new_n25128_,
    new_n25129_, new_n25130_, new_n25131_, new_n25132_, new_n25133_,
    new_n25134_, new_n25135_, new_n25136_, new_n25137_, new_n25138_,
    new_n25139_, new_n25140_, new_n25141_, new_n25142_, new_n25143_,
    new_n25144_, new_n25145_, new_n25146_, new_n25147_, new_n25148_,
    new_n25149_, new_n25150_, new_n25151_, new_n25152_, new_n25153_,
    new_n25154_, new_n25155_, new_n25156_, new_n25157_, new_n25158_,
    new_n25159_, new_n25160_, new_n25161_, new_n25162_, new_n25163_,
    new_n25164_, new_n25165_, new_n25166_, new_n25167_, new_n25168_,
    new_n25169_, new_n25170_, new_n25171_, new_n25172_, new_n25173_,
    new_n25174_, new_n25175_, new_n25176_, new_n25177_, new_n25178_,
    new_n25179_, new_n25180_, new_n25181_, new_n25182_, new_n25183_,
    new_n25184_, new_n25185_, new_n25186_, new_n25187_, new_n25188_,
    new_n25189_, new_n25190_, new_n25191_, new_n25192_, new_n25193_,
    new_n25194_, new_n25195_, new_n25196_, new_n25197_, new_n25198_,
    new_n25199_, new_n25200_, new_n25201_, new_n25202_, new_n25203_,
    new_n25204_, new_n25205_, new_n25206_, new_n25207_, new_n25208_,
    new_n25209_, new_n25210_, new_n25211_, new_n25212_, new_n25213_,
    new_n25214_, new_n25215_, new_n25216_, new_n25217_, new_n25218_,
    new_n25219_, new_n25220_, new_n25221_, new_n25222_, new_n25223_,
    new_n25224_, new_n25225_, new_n25226_, new_n25227_, new_n25228_,
    new_n25229_, new_n25230_, new_n25231_, new_n25232_, new_n25233_,
    new_n25234_, new_n25235_, new_n25236_, new_n25237_, new_n25238_,
    new_n25239_, new_n25240_, new_n25241_, new_n25242_, new_n25243_,
    new_n25244_, new_n25245_, new_n25246_, new_n25247_, new_n25248_,
    new_n25249_, new_n25250_, new_n25251_, new_n25252_, new_n25253_,
    new_n25254_, new_n25255_, new_n25256_, new_n25257_, new_n25258_,
    new_n25259_, new_n25260_, new_n25261_, new_n25262_, new_n25263_,
    new_n25264_, new_n25265_, new_n25266_, new_n25267_, new_n25268_,
    new_n25269_, new_n25270_, new_n25271_, new_n25272_, new_n25273_,
    new_n25274_, new_n25275_, new_n25276_, new_n25277_, new_n25278_,
    new_n25279_, new_n25280_, new_n25281_, new_n25282_, new_n25283_,
    new_n25284_, new_n25285_, new_n25286_, new_n25287_, new_n25288_,
    new_n25289_, new_n25290_, new_n25291_, new_n25292_, new_n25293_,
    new_n25294_, new_n25295_, new_n25296_, new_n25297_, new_n25298_,
    new_n25299_, new_n25300_, new_n25301_, new_n25302_, new_n25303_,
    new_n25304_, new_n25305_, new_n25306_, new_n25307_, new_n25308_,
    new_n25309_, new_n25310_, new_n25311_, new_n25312_, new_n25313_,
    new_n25314_, new_n25315_, new_n25316_, new_n25317_, new_n25318_,
    new_n25319_, new_n25320_, new_n25321_, new_n25322_, new_n25323_,
    new_n25324_, new_n25325_, new_n25326_, new_n25327_, new_n25328_,
    new_n25329_, new_n25330_, new_n25331_, new_n25332_, new_n25333_,
    new_n25334_, new_n25335_, new_n25336_, new_n25337_, new_n25338_,
    new_n25339_, new_n25340_, new_n25341_, new_n25342_, new_n25343_,
    new_n25344_, new_n25345_, new_n25346_, new_n25347_, new_n25348_,
    new_n25349_, new_n25350_, new_n25351_, new_n25352_, new_n25353_,
    new_n25354_, new_n25355_, new_n25356_, new_n25357_, new_n25358_,
    new_n25359_, new_n25360_, new_n25361_, new_n25362_, new_n25363_,
    new_n25364_, new_n25365_, new_n25366_, new_n25367_, new_n25368_,
    new_n25369_, new_n25370_, new_n25371_, new_n25372_, new_n25373_,
    new_n25374_, new_n25375_, new_n25376_, new_n25377_, new_n25378_,
    new_n25379_, new_n25380_, new_n25381_, new_n25382_, new_n25383_,
    new_n25384_, new_n25385_, new_n25386_, new_n25387_, new_n25388_,
    new_n25389_, new_n25390_, new_n25391_, new_n25392_, new_n25393_,
    new_n25394_, new_n25395_, new_n25396_, new_n25397_, new_n25398_,
    new_n25399_, new_n25400_, new_n25401_, new_n25402_, new_n25403_,
    new_n25404_, new_n25405_, new_n25406_, new_n25407_, new_n25408_,
    new_n25409_, new_n25410_, new_n25411_, new_n25412_, new_n25413_,
    new_n25414_, new_n25415_, new_n25416_, new_n25417_, new_n25418_,
    new_n25419_, new_n25420_, new_n25421_, new_n25422_, new_n25423_,
    new_n25424_, new_n25425_, new_n25426_, new_n25427_, new_n25428_,
    new_n25429_, new_n25430_, new_n25431_, new_n25432_, new_n25433_,
    new_n25434_, new_n25435_, new_n25436_, new_n25437_, new_n25438_,
    new_n25439_, new_n25440_, new_n25441_, new_n25442_, new_n25443_,
    new_n25444_, new_n25445_, new_n25446_, new_n25447_, new_n25448_,
    new_n25449_, new_n25450_, new_n25451_, new_n25452_, new_n25453_,
    new_n25454_, new_n25455_, new_n25456_, new_n25457_, new_n25458_,
    new_n25459_, new_n25460_, new_n25461_, new_n25462_, new_n25463_,
    new_n25464_, new_n25465_, new_n25466_, new_n25467_, new_n25468_,
    new_n25469_, new_n25470_, new_n25471_, new_n25472_, new_n25473_,
    new_n25474_, new_n25475_, new_n25476_, new_n25477_, new_n25478_,
    new_n25479_, new_n25480_, new_n25481_, new_n25482_, new_n25483_,
    new_n25484_, new_n25485_, new_n25486_, new_n25487_, new_n25488_,
    new_n25489_, new_n25490_, new_n25491_, new_n25492_, new_n25493_,
    new_n25494_, new_n25495_, new_n25496_, new_n25497_, new_n25498_,
    new_n25499_, new_n25500_, new_n25501_, new_n25502_, new_n25503_,
    new_n25504_, new_n25505_, new_n25506_, new_n25507_, new_n25508_,
    new_n25509_, new_n25510_, new_n25511_, new_n25512_, new_n25513_,
    new_n25514_, new_n25515_, new_n25516_, new_n25517_, new_n25518_,
    new_n25519_, new_n25520_, new_n25521_, new_n25522_, new_n25523_,
    new_n25524_, new_n25525_, new_n25526_, new_n25527_, new_n25528_,
    new_n25529_, new_n25530_, new_n25531_, new_n25532_, new_n25533_,
    new_n25534_, new_n25535_, new_n25536_, new_n25537_, new_n25538_,
    new_n25539_, new_n25540_, new_n25541_, new_n25542_, new_n25543_,
    new_n25544_, new_n25545_, new_n25546_, new_n25547_, new_n25548_,
    new_n25549_, new_n25550_, new_n25551_, new_n25552_, new_n25553_,
    new_n25554_, new_n25555_, new_n25556_, new_n25557_, new_n25558_,
    new_n25559_, new_n25560_, new_n25561_, new_n25562_, new_n25563_,
    new_n25564_, new_n25565_, new_n25566_, new_n25567_, new_n25568_,
    new_n25569_, new_n25570_, new_n25571_, new_n25572_, new_n25573_,
    new_n25574_, new_n25575_, new_n25576_, new_n25577_, new_n25578_,
    new_n25579_, new_n25580_, new_n25581_, new_n25582_, new_n25583_,
    new_n25584_, new_n25585_, new_n25586_, new_n25587_, new_n25588_,
    new_n25589_, new_n25590_, new_n25591_, new_n25592_, new_n25594_,
    new_n25595_, new_n25596_, new_n25597_, new_n25598_, new_n25599_,
    new_n25600_, new_n25601_, new_n25602_, new_n25603_, new_n25604_,
    new_n25605_, new_n25606_, new_n25607_, new_n25608_, new_n25609_,
    new_n25610_, new_n25611_, new_n25612_, new_n25613_, new_n25614_,
    new_n25615_, new_n25616_, new_n25617_, new_n25618_, new_n25619_,
    new_n25620_, new_n25621_, new_n25622_, new_n25623_, new_n25624_,
    new_n25625_, new_n25626_, new_n25627_, new_n25628_, new_n25629_,
    new_n25630_, new_n25631_, new_n25632_, new_n25633_, new_n25634_,
    new_n25635_, new_n25636_, new_n25637_, new_n25638_, new_n25639_,
    new_n25640_, new_n25641_, new_n25642_, new_n25643_, new_n25644_,
    new_n25645_, new_n25646_, new_n25647_, new_n25648_, new_n25649_,
    new_n25650_, new_n25651_, new_n25652_, new_n25653_, new_n25654_,
    new_n25655_, new_n25656_, new_n25657_, new_n25658_, new_n25659_,
    new_n25660_, new_n25661_, new_n25662_, new_n25663_, new_n25664_,
    new_n25665_, new_n25666_, new_n25667_, new_n25668_, new_n25669_,
    new_n25670_, new_n25671_, new_n25672_, new_n25673_, new_n25674_,
    new_n25675_, new_n25676_, new_n25677_, new_n25678_, new_n25679_,
    new_n25680_, new_n25681_, new_n25682_, new_n25683_, new_n25684_,
    new_n25685_, new_n25686_, new_n25687_, new_n25688_, new_n25689_,
    new_n25690_, new_n25691_, new_n25692_, new_n25693_, new_n25694_,
    new_n25695_, new_n25696_, new_n25697_, new_n25698_, new_n25699_,
    new_n25700_, new_n25701_, new_n25702_, new_n25703_, new_n25704_,
    new_n25705_, new_n25706_, new_n25707_, new_n25708_, new_n25709_,
    new_n25710_, new_n25711_, new_n25712_, new_n25713_, new_n25714_,
    new_n25715_, new_n25716_, new_n25717_, new_n25718_, new_n25719_,
    new_n25720_, new_n25721_, new_n25722_, new_n25723_, new_n25724_,
    new_n25725_, new_n25726_, new_n25727_, new_n25728_, new_n25729_,
    new_n25730_, new_n25731_, new_n25732_, new_n25733_, new_n25734_,
    new_n25735_, new_n25736_, new_n25737_, new_n25738_, new_n25739_,
    new_n25740_, new_n25741_, new_n25742_, new_n25743_, new_n25744_,
    new_n25745_, new_n25746_, new_n25747_, new_n25748_, new_n25749_,
    new_n25750_, new_n25751_, new_n25752_, new_n25753_, new_n25754_,
    new_n25755_, new_n25756_, new_n25757_, new_n25758_, new_n25759_,
    new_n25760_, new_n25761_, new_n25762_, new_n25763_, new_n25764_,
    new_n25765_, new_n25766_, new_n25767_, new_n25768_, new_n25769_,
    new_n25770_, new_n25771_, new_n25772_, new_n25773_, new_n25774_,
    new_n25775_, new_n25776_, new_n25777_, new_n25778_, new_n25779_,
    new_n25780_, new_n25781_, new_n25782_, new_n25783_, new_n25784_,
    new_n25785_, new_n25786_, new_n25787_, new_n25788_, new_n25789_,
    new_n25790_, new_n25791_, new_n25792_, new_n25793_, new_n25794_,
    new_n25795_, new_n25796_, new_n25797_, new_n25798_, new_n25799_,
    new_n25800_, new_n25801_, new_n25802_, new_n25803_, new_n25804_,
    new_n25805_, new_n25806_, new_n25807_, new_n25808_, new_n25809_,
    new_n25810_, new_n25811_, new_n25812_, new_n25813_, new_n25814_,
    new_n25815_, new_n25816_, new_n25817_, new_n25818_, new_n25819_,
    new_n25820_, new_n25821_, new_n25822_, new_n25823_, new_n25824_,
    new_n25825_, new_n25826_, new_n25827_, new_n25828_, new_n25829_,
    new_n25830_, new_n25831_, new_n25832_, new_n25833_, new_n25834_,
    new_n25835_, new_n25836_, new_n25837_, new_n25838_, new_n25839_,
    new_n25840_, new_n25841_, new_n25842_, new_n25843_, new_n25844_,
    new_n25845_, new_n25846_, new_n25847_, new_n25848_, new_n25849_,
    new_n25850_, new_n25851_, new_n25852_, new_n25853_, new_n25854_,
    new_n25855_, new_n25856_, new_n25857_, new_n25858_, new_n25859_,
    new_n25860_, new_n25861_, new_n25862_, new_n25863_, new_n25864_,
    new_n25865_, new_n25866_, new_n25867_, new_n25868_, new_n25869_,
    new_n25870_, new_n25871_, new_n25872_, new_n25873_, new_n25874_,
    new_n25875_, new_n25876_, new_n25877_, new_n25878_, new_n25879_,
    new_n25880_, new_n25881_, new_n25882_, new_n25883_, new_n25884_,
    new_n25885_, new_n25886_, new_n25887_, new_n25888_, new_n25889_,
    new_n25890_, new_n25891_, new_n25892_, new_n25893_, new_n25894_,
    new_n25895_, new_n25896_, new_n25897_, new_n25898_, new_n25899_,
    new_n25900_, new_n25901_, new_n25902_, new_n25903_, new_n25904_,
    new_n25905_, new_n25906_, new_n25907_, new_n25908_, new_n25909_,
    new_n25910_, new_n25911_, new_n25912_, new_n25913_, new_n25914_,
    new_n25915_, new_n25916_, new_n25917_, new_n25918_, new_n25919_,
    new_n25920_, new_n25921_, new_n25922_, new_n25923_, new_n25924_,
    new_n25925_, new_n25926_, new_n25927_, new_n25928_, new_n25929_,
    new_n25930_, new_n25931_, new_n25932_, new_n25933_, new_n25934_,
    new_n25935_, new_n25936_, new_n25937_, new_n25938_, new_n25939_,
    new_n25940_, new_n25941_, new_n25942_, new_n25943_, new_n25944_,
    new_n25945_, new_n25946_, new_n25947_, new_n25948_, new_n25949_,
    new_n25950_, new_n25951_, new_n25952_, new_n25953_, new_n25954_,
    new_n25955_, new_n25956_, new_n25957_, new_n25958_, new_n25959_,
    new_n25960_, new_n25961_, new_n25962_, new_n25963_, new_n25964_,
    new_n25965_, new_n25966_, new_n25967_, new_n25968_, new_n25969_,
    new_n25970_, new_n25971_, new_n25972_, new_n25973_, new_n25974_,
    new_n25975_, new_n25976_, new_n25977_, new_n25978_, new_n25979_,
    new_n25980_, new_n25981_, new_n25982_, new_n25983_, new_n25984_,
    new_n25985_, new_n25986_, new_n25987_, new_n25988_, new_n25989_,
    new_n25990_, new_n25991_, new_n25992_, new_n25993_, new_n25994_,
    new_n25995_, new_n25996_, new_n25997_, new_n25998_, new_n25999_,
    new_n26000_, new_n26001_, new_n26002_, new_n26003_, new_n26004_,
    new_n26005_, new_n26006_, new_n26007_, new_n26008_, new_n26009_,
    new_n26010_, new_n26011_, new_n26012_, new_n26013_, new_n26014_,
    new_n26015_, new_n26016_, new_n26017_, new_n26018_, new_n26019_,
    new_n26020_, new_n26021_, new_n26022_, new_n26023_, new_n26024_,
    new_n26025_, new_n26026_, new_n26027_, new_n26028_, new_n26029_,
    new_n26030_, new_n26031_, new_n26032_, new_n26033_, new_n26034_,
    new_n26035_, new_n26036_, new_n26037_, new_n26038_, new_n26039_,
    new_n26040_, new_n26041_, new_n26042_, new_n26043_, new_n26044_,
    new_n26045_, new_n26046_, new_n26047_, new_n26048_, new_n26049_,
    new_n26050_, new_n26051_, new_n26052_, new_n26053_, new_n26054_,
    new_n26055_, new_n26056_, new_n26057_, new_n26058_, new_n26059_,
    new_n26060_, new_n26061_, new_n26062_, new_n26063_, new_n26064_,
    new_n26065_, new_n26066_, new_n26067_, new_n26068_, new_n26069_,
    new_n26070_, new_n26071_, new_n26072_, new_n26073_, new_n26074_,
    new_n26076_, new_n26077_, new_n26078_, new_n26079_, new_n26080_,
    new_n26081_, new_n26082_, new_n26083_, new_n26084_, new_n26085_,
    new_n26086_, new_n26087_, new_n26088_, new_n26089_, new_n26090_,
    new_n26091_, new_n26092_, new_n26093_, new_n26094_, new_n26095_,
    new_n26096_, new_n26097_, new_n26098_, new_n26099_, new_n26100_,
    new_n26101_, new_n26102_, new_n26103_, new_n26104_, new_n26105_,
    new_n26106_, new_n26107_, new_n26108_, new_n26109_, new_n26110_,
    new_n26111_, new_n26112_, new_n26113_, new_n26114_, new_n26115_,
    new_n26116_, new_n26117_, new_n26118_, new_n26119_, new_n26120_,
    new_n26121_, new_n26122_, new_n26123_, new_n26124_, new_n26125_,
    new_n26126_, new_n26127_, new_n26128_, new_n26129_, new_n26130_,
    new_n26131_, new_n26132_, new_n26133_, new_n26134_, new_n26135_,
    new_n26136_, new_n26137_, new_n26138_, new_n26139_, new_n26140_,
    new_n26141_, new_n26142_, new_n26143_, new_n26144_, new_n26145_,
    new_n26146_, new_n26147_, new_n26148_, new_n26149_, new_n26150_,
    new_n26151_, new_n26152_, new_n26153_, new_n26154_, new_n26155_,
    new_n26156_, new_n26157_, new_n26158_, new_n26159_, new_n26160_,
    new_n26161_, new_n26162_, new_n26163_, new_n26164_, new_n26165_,
    new_n26166_, new_n26167_, new_n26168_, new_n26169_, new_n26170_,
    new_n26171_, new_n26172_, new_n26173_, new_n26174_, new_n26175_,
    new_n26176_, new_n26177_, new_n26178_, new_n26179_, new_n26180_,
    new_n26181_, new_n26182_, new_n26183_, new_n26184_, new_n26185_,
    new_n26186_, new_n26187_, new_n26188_, new_n26189_, new_n26190_,
    new_n26191_, new_n26192_, new_n26193_, new_n26194_, new_n26195_,
    new_n26196_, new_n26197_, new_n26198_, new_n26199_, new_n26200_,
    new_n26201_, new_n26202_, new_n26203_, new_n26204_, new_n26205_,
    new_n26206_, new_n26207_, new_n26208_, new_n26209_, new_n26210_,
    new_n26211_, new_n26212_, new_n26213_, new_n26214_, new_n26215_,
    new_n26216_, new_n26217_, new_n26218_, new_n26219_, new_n26220_,
    new_n26221_, new_n26222_, new_n26223_, new_n26224_, new_n26225_,
    new_n26226_, new_n26227_, new_n26228_, new_n26229_, new_n26230_,
    new_n26231_, new_n26232_, new_n26233_, new_n26234_, new_n26235_,
    new_n26236_, new_n26237_, new_n26238_, new_n26239_, new_n26240_,
    new_n26241_, new_n26242_, new_n26243_, new_n26244_, new_n26245_,
    new_n26246_, new_n26247_, new_n26248_, new_n26249_, new_n26250_,
    new_n26251_, new_n26252_, new_n26253_, new_n26254_, new_n26255_,
    new_n26256_, new_n26257_, new_n26258_, new_n26259_, new_n26260_,
    new_n26261_, new_n26262_, new_n26263_, new_n26264_, new_n26265_,
    new_n26266_, new_n26267_, new_n26268_, new_n26269_, new_n26270_,
    new_n26271_, new_n26272_, new_n26273_, new_n26274_, new_n26275_,
    new_n26276_, new_n26277_, new_n26278_, new_n26279_, new_n26280_,
    new_n26281_, new_n26282_, new_n26283_, new_n26284_, new_n26285_,
    new_n26286_, new_n26287_, new_n26288_, new_n26289_, new_n26290_,
    new_n26291_, new_n26292_, new_n26293_, new_n26294_, new_n26295_,
    new_n26296_, new_n26297_, new_n26298_, new_n26299_, new_n26300_,
    new_n26301_, new_n26302_, new_n26303_, new_n26304_, new_n26305_,
    new_n26306_, new_n26307_, new_n26308_, new_n26309_, new_n26310_,
    new_n26311_, new_n26312_, new_n26313_, new_n26314_, new_n26315_,
    new_n26316_, new_n26317_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26326_, new_n26327_, new_n26328_, new_n26329_, new_n26330_,
    new_n26331_, new_n26332_, new_n26333_, new_n26334_, new_n26335_,
    new_n26336_, new_n26337_, new_n26338_, new_n26339_, new_n26340_,
    new_n26341_, new_n26342_, new_n26343_, new_n26344_, new_n26345_,
    new_n26346_, new_n26347_, new_n26348_, new_n26349_, new_n26350_,
    new_n26351_, new_n26352_, new_n26353_, new_n26354_, new_n26355_,
    new_n26356_, new_n26357_, new_n26358_, new_n26359_, new_n26360_,
    new_n26361_, new_n26362_, new_n26363_, new_n26364_, new_n26365_,
    new_n26366_, new_n26367_, new_n26368_, new_n26369_, new_n26370_,
    new_n26371_, new_n26372_, new_n26373_, new_n26374_, new_n26375_,
    new_n26376_, new_n26377_, new_n26378_, new_n26379_, new_n26380_,
    new_n26381_, new_n26382_, new_n26383_, new_n26384_, new_n26385_,
    new_n26386_, new_n26387_, new_n26388_, new_n26389_, new_n26390_,
    new_n26391_, new_n26392_, new_n26393_, new_n26394_, new_n26395_,
    new_n26396_, new_n26397_, new_n26398_, new_n26399_, new_n26400_,
    new_n26401_, new_n26402_, new_n26403_, new_n26404_, new_n26405_,
    new_n26406_, new_n26407_, new_n26408_, new_n26409_, new_n26410_,
    new_n26411_, new_n26412_, new_n26413_, new_n26414_, new_n26415_,
    new_n26416_, new_n26417_, new_n26418_, new_n26419_, new_n26420_,
    new_n26421_, new_n26422_, new_n26423_, new_n26424_, new_n26425_,
    new_n26426_, new_n26427_, new_n26428_, new_n26429_, new_n26430_,
    new_n26431_, new_n26432_, new_n26433_, new_n26434_, new_n26435_,
    new_n26436_, new_n26437_, new_n26438_, new_n26439_, new_n26440_,
    new_n26441_, new_n26442_, new_n26443_, new_n26444_, new_n26445_,
    new_n26446_, new_n26447_, new_n26448_, new_n26449_, new_n26450_,
    new_n26451_, new_n26452_, new_n26453_, new_n26454_, new_n26455_,
    new_n26456_, new_n26457_, new_n26458_, new_n26459_, new_n26460_,
    new_n26461_, new_n26462_, new_n26463_, new_n26464_, new_n26465_,
    new_n26466_, new_n26467_, new_n26468_, new_n26469_, new_n26470_,
    new_n26471_, new_n26472_, new_n26473_, new_n26474_, new_n26475_,
    new_n26476_, new_n26477_, new_n26478_, new_n26479_, new_n26480_,
    new_n26481_, new_n26482_, new_n26483_, new_n26484_, new_n26485_,
    new_n26486_, new_n26487_, new_n26488_, new_n26489_, new_n26490_,
    new_n26491_, new_n26492_, new_n26493_, new_n26494_, new_n26495_,
    new_n26496_, new_n26497_, new_n26498_, new_n26499_, new_n26500_,
    new_n26501_, new_n26502_, new_n26503_, new_n26504_, new_n26505_,
    new_n26506_, new_n26507_, new_n26508_, new_n26509_, new_n26510_,
    new_n26511_, new_n26512_, new_n26513_, new_n26514_, new_n26515_,
    new_n26516_, new_n26517_, new_n26518_, new_n26519_, new_n26520_,
    new_n26521_, new_n26522_, new_n26523_, new_n26524_, new_n26525_,
    new_n26526_, new_n26527_, new_n26528_, new_n26529_, new_n26530_,
    new_n26531_, new_n26532_, new_n26533_, new_n26534_, new_n26535_,
    new_n26536_, new_n26537_, new_n26538_, new_n26539_, new_n26540_,
    new_n26541_, new_n26542_, new_n26543_, new_n26544_, new_n26545_,
    new_n26546_, new_n26547_, new_n26548_, new_n26549_, new_n26550_,
    new_n26551_, new_n26553_, new_n26554_, new_n26555_, new_n26556_,
    new_n26557_, new_n26558_, new_n26559_, new_n26560_, new_n26561_,
    new_n26562_, new_n26563_, new_n26564_, new_n26565_, new_n26566_,
    new_n26567_, new_n26568_, new_n26569_, new_n26570_, new_n26571_,
    new_n26572_, new_n26573_, new_n26574_, new_n26575_, new_n26576_,
    new_n26577_, new_n26578_, new_n26579_, new_n26580_, new_n26581_,
    new_n26582_, new_n26583_, new_n26584_, new_n26585_, new_n26586_,
    new_n26587_, new_n26588_, new_n26589_, new_n26590_, new_n26591_,
    new_n26592_, new_n26593_, new_n26594_, new_n26595_, new_n26596_,
    new_n26597_, new_n26598_, new_n26599_, new_n26600_, new_n26601_,
    new_n26602_, new_n26603_, new_n26604_, new_n26605_, new_n26606_,
    new_n26607_, new_n26608_, new_n26609_, new_n26610_, new_n26611_,
    new_n26612_, new_n26613_, new_n26614_, new_n26615_, new_n26616_,
    new_n26617_, new_n26618_, new_n26619_, new_n26620_, new_n26621_,
    new_n26622_, new_n26623_, new_n26624_, new_n26625_, new_n26626_,
    new_n26627_, new_n26628_, new_n26629_, new_n26630_, new_n26631_,
    new_n26632_, new_n26633_, new_n26634_, new_n26635_, new_n26636_,
    new_n26637_, new_n26638_, new_n26639_, new_n26640_, new_n26641_,
    new_n26642_, new_n26643_, new_n26644_, new_n26645_, new_n26646_,
    new_n26647_, new_n26648_, new_n26649_, new_n26650_, new_n26651_,
    new_n26652_, new_n26653_, new_n26654_, new_n26655_, new_n26656_,
    new_n26657_, new_n26658_, new_n26659_, new_n26660_, new_n26661_,
    new_n26662_, new_n26663_, new_n26664_, new_n26665_, new_n26666_,
    new_n26667_, new_n26668_, new_n26669_, new_n26670_, new_n26671_,
    new_n26672_, new_n26673_, new_n26674_, new_n26675_, new_n26676_,
    new_n26677_, new_n26678_, new_n26679_, new_n26680_, new_n26681_,
    new_n26682_, new_n26683_, new_n26684_, new_n26685_, new_n26686_,
    new_n26687_, new_n26688_, new_n26689_, new_n26690_, new_n26691_,
    new_n26692_, new_n26693_, new_n26694_, new_n26695_, new_n26696_,
    new_n26697_, new_n26698_, new_n26699_, new_n26700_, new_n26701_,
    new_n26702_, new_n26703_, new_n26704_, new_n26705_, new_n26706_,
    new_n26707_, new_n26708_, new_n26709_, new_n26710_, new_n26711_,
    new_n26712_, new_n26713_, new_n26714_, new_n26715_, new_n26716_,
    new_n26717_, new_n26718_, new_n26719_, new_n26720_, new_n26721_,
    new_n26722_, new_n26723_, new_n26724_, new_n26725_, new_n26726_,
    new_n26727_, new_n26728_, new_n26729_, new_n26730_, new_n26731_,
    new_n26732_, new_n26733_, new_n26734_, new_n26735_, new_n26736_,
    new_n26737_, new_n26738_, new_n26739_, new_n26740_, new_n26741_,
    new_n26742_, new_n26743_, new_n26744_, new_n26745_, new_n26746_,
    new_n26747_, new_n26748_, new_n26749_, new_n26750_, new_n26751_,
    new_n26752_, new_n26753_, new_n26754_, new_n26755_, new_n26756_,
    new_n26757_, new_n26758_, new_n26759_, new_n26760_, new_n26761_,
    new_n26762_, new_n26763_, new_n26764_, new_n26765_, new_n26766_,
    new_n26767_, new_n26768_, new_n26769_, new_n26770_, new_n26771_,
    new_n26772_, new_n26773_, new_n26774_, new_n26775_, new_n26776_,
    new_n26777_, new_n26778_, new_n26779_, new_n26780_, new_n26781_,
    new_n26782_, new_n26783_, new_n26784_, new_n26785_, new_n26786_,
    new_n26787_, new_n26788_, new_n26789_, new_n26790_, new_n26791_,
    new_n26792_, new_n26793_, new_n26794_, new_n26795_, new_n26796_,
    new_n26797_, new_n26798_, new_n26799_, new_n26800_, new_n26801_,
    new_n26802_, new_n26803_, new_n26804_, new_n26805_, new_n26806_,
    new_n26807_, new_n26808_, new_n26809_, new_n26810_, new_n26811_,
    new_n26812_, new_n26813_, new_n26814_, new_n26815_, new_n26816_,
    new_n26817_, new_n26818_, new_n26819_, new_n26820_, new_n26821_,
    new_n26822_, new_n26823_, new_n26824_, new_n26825_, new_n26826_,
    new_n26827_, new_n26828_, new_n26829_, new_n26830_, new_n26831_,
    new_n26832_, new_n26833_, new_n26834_, new_n26835_, new_n26836_,
    new_n26837_, new_n26838_, new_n26839_, new_n26840_, new_n26841_,
    new_n26842_, new_n26843_, new_n26844_, new_n26845_, new_n26846_,
    new_n26847_, new_n26848_, new_n26849_, new_n26850_, new_n26851_,
    new_n26852_, new_n26853_, new_n26854_, new_n26855_, new_n26856_,
    new_n26857_, new_n26858_, new_n26859_, new_n26860_, new_n26861_,
    new_n26862_, new_n26863_, new_n26864_, new_n26865_, new_n26866_,
    new_n26867_, new_n26868_, new_n26869_, new_n26870_, new_n26871_,
    new_n26872_, new_n26873_, new_n26874_, new_n26875_, new_n26876_,
    new_n26877_, new_n26878_, new_n26879_, new_n26880_, new_n26881_,
    new_n26882_, new_n26883_, new_n26884_, new_n26885_, new_n26886_,
    new_n26887_, new_n26888_, new_n26889_, new_n26890_, new_n26891_,
    new_n26892_, new_n26893_, new_n26894_, new_n26895_, new_n26896_,
    new_n26897_, new_n26898_, new_n26899_, new_n26900_, new_n26901_,
    new_n26902_, new_n26903_, new_n26904_, new_n26905_, new_n26906_,
    new_n26907_, new_n26908_, new_n26909_, new_n26910_, new_n26911_,
    new_n26912_, new_n26913_, new_n26914_, new_n26915_, new_n26916_,
    new_n26917_, new_n26918_, new_n26919_, new_n26920_, new_n26921_,
    new_n26922_, new_n26923_, new_n26924_, new_n26925_, new_n26926_,
    new_n26927_, new_n26928_, new_n26929_, new_n26930_, new_n26931_,
    new_n26932_, new_n26933_, new_n26934_, new_n26935_, new_n26936_,
    new_n26937_, new_n26938_, new_n26939_, new_n26940_, new_n26941_,
    new_n26942_, new_n26943_, new_n26944_, new_n26945_, new_n26946_,
    new_n26947_, new_n26948_, new_n26949_, new_n26950_, new_n26951_,
    new_n26952_, new_n26953_, new_n26954_, new_n26955_, new_n26956_,
    new_n26957_, new_n26958_, new_n26959_, new_n26960_, new_n26961_,
    new_n26962_, new_n26963_, new_n26964_, new_n26965_, new_n26966_,
    new_n26967_, new_n26968_, new_n26969_, new_n26970_, new_n26971_,
    new_n26972_, new_n26973_, new_n26974_, new_n26975_, new_n26976_,
    new_n26977_, new_n26978_, new_n26979_, new_n26980_, new_n26981_,
    new_n26982_, new_n26983_, new_n26984_, new_n26985_, new_n26986_,
    new_n26987_, new_n26988_, new_n26989_, new_n26990_, new_n26991_,
    new_n26992_, new_n26993_, new_n26994_, new_n26995_, new_n26996_,
    new_n26997_, new_n26998_, new_n26999_, new_n27000_, new_n27001_,
    new_n27002_, new_n27003_, new_n27004_, new_n27005_, new_n27006_,
    new_n27007_, new_n27008_, new_n27009_, new_n27010_, new_n27011_,
    new_n27012_, new_n27013_, new_n27014_, new_n27015_, new_n27016_,
    new_n27017_, new_n27018_, new_n27019_, new_n27020_, new_n27021_,
    new_n27022_, new_n27023_, new_n27024_, new_n27025_, new_n27026_,
    new_n27027_, new_n27028_, new_n27030_, new_n27031_, new_n27032_,
    new_n27033_, new_n27034_, new_n27035_, new_n27036_, new_n27037_,
    new_n27038_, new_n27039_, new_n27040_, new_n27041_, new_n27042_,
    new_n27043_, new_n27044_, new_n27045_, new_n27046_, new_n27047_,
    new_n27048_, new_n27049_, new_n27050_, new_n27051_, new_n27052_,
    new_n27053_, new_n27054_, new_n27055_, new_n27056_, new_n27057_,
    new_n27058_, new_n27059_, new_n27060_, new_n27061_, new_n27062_,
    new_n27063_, new_n27064_, new_n27065_, new_n27066_, new_n27067_,
    new_n27068_, new_n27069_, new_n27070_, new_n27071_, new_n27072_,
    new_n27073_, new_n27074_, new_n27075_, new_n27076_, new_n27077_,
    new_n27078_, new_n27079_, new_n27080_, new_n27081_, new_n27082_,
    new_n27083_, new_n27084_, new_n27085_, new_n27086_, new_n27087_,
    new_n27088_, new_n27089_, new_n27090_, new_n27091_, new_n27092_,
    new_n27093_, new_n27094_, new_n27095_, new_n27096_, new_n27097_,
    new_n27098_, new_n27099_, new_n27100_, new_n27101_, new_n27102_,
    new_n27103_, new_n27104_, new_n27105_, new_n27106_, new_n27107_,
    new_n27108_, new_n27109_, new_n27110_, new_n27111_, new_n27112_,
    new_n27113_, new_n27114_, new_n27115_, new_n27116_, new_n27117_,
    new_n27118_, new_n27119_, new_n27120_, new_n27121_, new_n27122_,
    new_n27123_, new_n27124_, new_n27125_, new_n27126_, new_n27127_,
    new_n27128_, new_n27129_, new_n27130_, new_n27131_, new_n27132_,
    new_n27133_, new_n27134_, new_n27135_, new_n27136_, new_n27137_,
    new_n27138_, new_n27139_, new_n27140_, new_n27141_, new_n27142_,
    new_n27143_, new_n27144_, new_n27145_, new_n27146_, new_n27147_,
    new_n27148_, new_n27149_, new_n27150_, new_n27151_, new_n27152_,
    new_n27153_, new_n27154_, new_n27155_, new_n27156_, new_n27157_,
    new_n27158_, new_n27159_, new_n27160_, new_n27161_, new_n27162_,
    new_n27163_, new_n27164_, new_n27165_, new_n27166_, new_n27167_,
    new_n27168_, new_n27169_, new_n27170_, new_n27171_, new_n27172_,
    new_n27173_, new_n27174_, new_n27175_, new_n27176_, new_n27177_,
    new_n27178_, new_n27179_, new_n27180_, new_n27181_, new_n27182_,
    new_n27183_, new_n27184_, new_n27185_, new_n27186_, new_n27187_,
    new_n27188_, new_n27189_, new_n27190_, new_n27191_, new_n27192_,
    new_n27193_, new_n27194_, new_n27195_, new_n27196_, new_n27197_,
    new_n27198_, new_n27199_, new_n27200_, new_n27201_, new_n27202_,
    new_n27203_, new_n27204_, new_n27205_, new_n27206_, new_n27207_,
    new_n27208_, new_n27209_, new_n27210_, new_n27211_, new_n27212_,
    new_n27213_, new_n27214_, new_n27215_, new_n27216_, new_n27217_,
    new_n27218_, new_n27219_, new_n27220_, new_n27221_, new_n27222_,
    new_n27223_, new_n27224_, new_n27225_, new_n27226_, new_n27227_,
    new_n27228_, new_n27229_, new_n27230_, new_n27231_, new_n27232_,
    new_n27233_, new_n27234_, new_n27235_, new_n27236_, new_n27237_,
    new_n27238_, new_n27239_, new_n27240_, new_n27241_, new_n27242_,
    new_n27243_, new_n27244_, new_n27245_, new_n27246_, new_n27247_,
    new_n27248_, new_n27249_, new_n27250_, new_n27251_, new_n27252_,
    new_n27253_, new_n27254_, new_n27255_, new_n27256_, new_n27257_,
    new_n27258_, new_n27259_, new_n27260_, new_n27261_, new_n27262_,
    new_n27263_, new_n27264_, new_n27265_, new_n27266_, new_n27267_,
    new_n27268_, new_n27269_, new_n27270_, new_n27271_, new_n27272_,
    new_n27273_, new_n27274_, new_n27275_, new_n27276_, new_n27277_,
    new_n27278_, new_n27279_, new_n27280_, new_n27281_, new_n27282_,
    new_n27283_, new_n27284_, new_n27285_, new_n27286_, new_n27287_,
    new_n27288_, new_n27289_, new_n27290_, new_n27291_, new_n27292_,
    new_n27293_, new_n27294_, new_n27295_, new_n27296_, new_n27297_,
    new_n27298_, new_n27299_, new_n27300_, new_n27301_, new_n27302_,
    new_n27303_, new_n27304_, new_n27305_, new_n27306_, new_n27307_,
    new_n27308_, new_n27309_, new_n27310_, new_n27311_, new_n27312_,
    new_n27313_, new_n27314_, new_n27315_, new_n27316_, new_n27317_,
    new_n27318_, new_n27319_, new_n27320_, new_n27321_, new_n27322_,
    new_n27323_, new_n27324_, new_n27325_, new_n27326_, new_n27327_,
    new_n27328_, new_n27329_, new_n27330_, new_n27331_, new_n27332_,
    new_n27333_, new_n27334_, new_n27335_, new_n27336_, new_n27337_,
    new_n27338_, new_n27339_, new_n27340_, new_n27341_, new_n27342_,
    new_n27343_, new_n27344_, new_n27345_, new_n27346_, new_n27347_,
    new_n27348_, new_n27349_, new_n27350_, new_n27351_, new_n27352_,
    new_n27353_, new_n27354_, new_n27355_, new_n27356_, new_n27357_,
    new_n27358_, new_n27359_, new_n27360_, new_n27361_, new_n27362_,
    new_n27363_, new_n27364_, new_n27365_, new_n27366_, new_n27367_,
    new_n27368_, new_n27369_, new_n27370_, new_n27371_, new_n27372_,
    new_n27373_, new_n27374_, new_n27375_, new_n27376_, new_n27377_,
    new_n27378_, new_n27379_, new_n27380_, new_n27381_, new_n27382_,
    new_n27383_, new_n27384_, new_n27385_, new_n27386_, new_n27387_,
    new_n27388_, new_n27389_, new_n27390_, new_n27391_, new_n27392_,
    new_n27393_, new_n27394_, new_n27395_, new_n27396_, new_n27397_,
    new_n27398_, new_n27399_, new_n27400_, new_n27401_, new_n27402_,
    new_n27403_, new_n27404_, new_n27405_, new_n27406_, new_n27407_,
    new_n27408_, new_n27409_, new_n27410_, new_n27411_, new_n27412_,
    new_n27413_, new_n27414_, new_n27415_, new_n27416_, new_n27417_,
    new_n27418_, new_n27419_, new_n27420_, new_n27421_, new_n27422_,
    new_n27423_, new_n27424_, new_n27425_, new_n27426_, new_n27427_,
    new_n27428_, new_n27429_, new_n27430_, new_n27431_, new_n27432_,
    new_n27433_, new_n27434_, new_n27435_, new_n27436_, new_n27437_,
    new_n27438_, new_n27439_, new_n27440_, new_n27441_, new_n27442_,
    new_n27443_, new_n27444_, new_n27445_, new_n27446_, new_n27447_,
    new_n27448_, new_n27449_, new_n27450_, new_n27451_, new_n27452_,
    new_n27453_, new_n27454_, new_n27455_, new_n27456_, new_n27457_,
    new_n27458_, new_n27459_, new_n27460_, new_n27461_, new_n27462_,
    new_n27463_, new_n27464_, new_n27465_, new_n27466_, new_n27467_,
    new_n27468_, new_n27469_, new_n27470_, new_n27471_, new_n27472_,
    new_n27473_, new_n27474_, new_n27475_, new_n27476_, new_n27477_,
    new_n27478_, new_n27479_, new_n27480_, new_n27481_, new_n27482_,
    new_n27483_, new_n27484_, new_n27485_, new_n27486_, new_n27487_,
    new_n27488_, new_n27489_, new_n27490_, new_n27491_, new_n27492_,
    new_n27493_, new_n27494_, new_n27495_, new_n27496_, new_n27497_,
    new_n27498_, new_n27499_, new_n27501_, new_n27502_, new_n27503_,
    new_n27504_, new_n27505_, new_n27506_, new_n27507_, new_n27508_,
    new_n27509_, new_n27510_, new_n27511_, new_n27512_, new_n27513_,
    new_n27514_, new_n27515_, new_n27516_, new_n27517_, new_n27518_,
    new_n27519_, new_n27520_, new_n27521_, new_n27522_, new_n27523_,
    new_n27524_, new_n27525_, new_n27526_, new_n27527_, new_n27528_,
    new_n27529_, new_n27530_, new_n27531_, new_n27532_, new_n27533_,
    new_n27534_, new_n27535_, new_n27536_, new_n27537_, new_n27538_,
    new_n27539_, new_n27540_, new_n27541_, new_n27542_, new_n27543_,
    new_n27544_, new_n27545_, new_n27546_, new_n27547_, new_n27548_,
    new_n27549_, new_n27550_, new_n27551_, new_n27552_, new_n27553_,
    new_n27554_, new_n27555_, new_n27556_, new_n27557_, new_n27558_,
    new_n27559_, new_n27560_, new_n27561_, new_n27562_, new_n27563_,
    new_n27564_, new_n27565_, new_n27566_, new_n27567_, new_n27568_,
    new_n27569_, new_n27570_, new_n27571_, new_n27572_, new_n27573_,
    new_n27574_, new_n27575_, new_n27576_, new_n27577_, new_n27578_,
    new_n27579_, new_n27580_, new_n27581_, new_n27582_, new_n27583_,
    new_n27584_, new_n27585_, new_n27586_, new_n27587_, new_n27588_,
    new_n27589_, new_n27590_, new_n27591_, new_n27592_, new_n27593_,
    new_n27594_, new_n27595_, new_n27596_, new_n27597_, new_n27598_,
    new_n27599_, new_n27600_, new_n27601_, new_n27602_, new_n27603_,
    new_n27604_, new_n27605_, new_n27606_, new_n27607_, new_n27608_,
    new_n27609_, new_n27610_, new_n27611_, new_n27612_, new_n27613_,
    new_n27614_, new_n27615_, new_n27616_, new_n27617_, new_n27618_,
    new_n27619_, new_n27620_, new_n27621_, new_n27622_, new_n27623_,
    new_n27624_, new_n27625_, new_n27626_, new_n27627_, new_n27628_,
    new_n27629_, new_n27630_, new_n27631_, new_n27632_, new_n27633_,
    new_n27634_, new_n27635_, new_n27636_, new_n27637_, new_n27638_,
    new_n27639_, new_n27640_, new_n27641_, new_n27642_, new_n27643_,
    new_n27644_, new_n27645_, new_n27646_, new_n27647_, new_n27648_,
    new_n27649_, new_n27650_, new_n27651_, new_n27652_, new_n27653_,
    new_n27654_, new_n27655_, new_n27656_, new_n27657_, new_n27658_,
    new_n27659_, new_n27660_, new_n27661_, new_n27662_, new_n27663_,
    new_n27664_, new_n27665_, new_n27666_, new_n27667_, new_n27668_,
    new_n27669_, new_n27670_, new_n27671_, new_n27672_, new_n27673_,
    new_n27674_, new_n27675_, new_n27676_, new_n27677_, new_n27678_,
    new_n27679_, new_n27680_, new_n27681_, new_n27682_, new_n27683_,
    new_n27684_, new_n27685_, new_n27686_, new_n27687_, new_n27688_,
    new_n27689_, new_n27690_, new_n27691_, new_n27692_, new_n27693_,
    new_n27694_, new_n27695_, new_n27696_, new_n27697_, new_n27698_,
    new_n27699_, new_n27700_, new_n27701_, new_n27702_, new_n27703_,
    new_n27704_, new_n27705_, new_n27706_, new_n27707_, new_n27708_,
    new_n27709_, new_n27710_, new_n27711_, new_n27712_, new_n27713_,
    new_n27714_, new_n27715_, new_n27716_, new_n27717_, new_n27718_,
    new_n27719_, new_n27720_, new_n27721_, new_n27722_, new_n27723_,
    new_n27724_, new_n27725_, new_n27726_, new_n27727_, new_n27728_,
    new_n27729_, new_n27730_, new_n27731_, new_n27732_, new_n27733_,
    new_n27734_, new_n27735_, new_n27736_, new_n27737_, new_n27738_,
    new_n27739_, new_n27740_, new_n27741_, new_n27742_, new_n27743_,
    new_n27744_, new_n27745_, new_n27746_, new_n27747_, new_n27748_,
    new_n27749_, new_n27750_, new_n27751_, new_n27752_, new_n27753_,
    new_n27754_, new_n27755_, new_n27756_, new_n27757_, new_n27758_,
    new_n27759_, new_n27760_, new_n27761_, new_n27762_, new_n27763_,
    new_n27764_, new_n27765_, new_n27766_, new_n27767_, new_n27768_,
    new_n27769_, new_n27770_, new_n27771_, new_n27772_, new_n27773_,
    new_n27774_, new_n27775_, new_n27776_, new_n27777_, new_n27778_,
    new_n27779_, new_n27780_, new_n27781_, new_n27782_, new_n27783_,
    new_n27784_, new_n27785_, new_n27786_, new_n27787_, new_n27788_,
    new_n27789_, new_n27790_, new_n27791_, new_n27792_, new_n27793_,
    new_n27794_, new_n27795_, new_n27796_, new_n27797_, new_n27798_,
    new_n27799_, new_n27800_, new_n27801_, new_n27802_, new_n27803_,
    new_n27804_, new_n27805_, new_n27806_, new_n27807_, new_n27808_,
    new_n27809_, new_n27810_, new_n27811_, new_n27812_, new_n27813_,
    new_n27814_, new_n27815_, new_n27816_, new_n27817_, new_n27818_,
    new_n27819_, new_n27820_, new_n27821_, new_n27822_, new_n27823_,
    new_n27824_, new_n27825_, new_n27826_, new_n27827_, new_n27828_,
    new_n27829_, new_n27830_, new_n27831_, new_n27832_, new_n27833_,
    new_n27834_, new_n27835_, new_n27836_, new_n27837_, new_n27838_,
    new_n27839_, new_n27840_, new_n27841_, new_n27842_, new_n27843_,
    new_n27844_, new_n27845_, new_n27846_, new_n27847_, new_n27848_,
    new_n27849_, new_n27850_, new_n27851_, new_n27852_, new_n27853_,
    new_n27854_, new_n27855_, new_n27856_, new_n27857_, new_n27858_,
    new_n27859_, new_n27860_, new_n27861_, new_n27862_, new_n27863_,
    new_n27864_, new_n27865_, new_n27866_, new_n27867_, new_n27868_,
    new_n27869_, new_n27870_, new_n27871_, new_n27872_, new_n27873_,
    new_n27874_, new_n27875_, new_n27876_, new_n27877_, new_n27878_,
    new_n27879_, new_n27880_, new_n27881_, new_n27882_, new_n27883_,
    new_n27884_, new_n27885_, new_n27886_, new_n27887_, new_n27888_,
    new_n27889_, new_n27890_, new_n27891_, new_n27892_, new_n27893_,
    new_n27894_, new_n27895_, new_n27896_, new_n27897_, new_n27898_,
    new_n27899_, new_n27900_, new_n27901_, new_n27902_, new_n27903_,
    new_n27904_, new_n27905_, new_n27906_, new_n27907_, new_n27908_,
    new_n27909_, new_n27910_, new_n27911_, new_n27912_, new_n27913_,
    new_n27914_, new_n27915_, new_n27916_, new_n27917_, new_n27918_,
    new_n27919_, new_n27920_, new_n27921_, new_n27922_, new_n27923_,
    new_n27924_, new_n27925_, new_n27926_, new_n27927_, new_n27928_,
    new_n27929_, new_n27930_, new_n27931_, new_n27932_, new_n27933_,
    new_n27934_, new_n27935_, new_n27936_, new_n27937_, new_n27938_,
    new_n27939_, new_n27940_, new_n27941_, new_n27942_, new_n27943_,
    new_n27944_, new_n27945_, new_n27946_, new_n27947_, new_n27948_,
    new_n27949_, new_n27950_, new_n27951_, new_n27952_, new_n27953_,
    new_n27954_, new_n27955_, new_n27956_, new_n27957_, new_n27958_,
    new_n27959_, new_n27960_, new_n27961_, new_n27962_, new_n27963_,
    new_n27964_, new_n27965_, new_n27966_, new_n27967_, new_n27968_,
    new_n27969_, new_n27970_, new_n27972_, new_n27973_, new_n27974_,
    new_n27975_, new_n27976_, new_n27977_, new_n27978_, new_n27979_,
    new_n27980_, new_n27981_, new_n27982_, new_n27983_, new_n27984_,
    new_n27985_, new_n27986_, new_n27987_, new_n27988_, new_n27989_,
    new_n27990_, new_n27991_, new_n27992_, new_n27993_, new_n27994_,
    new_n27995_, new_n27996_, new_n27997_, new_n27998_, new_n27999_,
    new_n28000_, new_n28001_, new_n28002_, new_n28003_, new_n28004_,
    new_n28005_, new_n28006_, new_n28007_, new_n28008_, new_n28009_,
    new_n28010_, new_n28011_, new_n28012_, new_n28013_, new_n28014_,
    new_n28015_, new_n28016_, new_n28017_, new_n28018_, new_n28019_,
    new_n28020_, new_n28021_, new_n28022_, new_n28023_, new_n28024_,
    new_n28025_, new_n28026_, new_n28027_, new_n28028_, new_n28029_,
    new_n28030_, new_n28031_, new_n28032_, new_n28033_, new_n28034_,
    new_n28035_, new_n28036_, new_n28037_, new_n28038_, new_n28039_,
    new_n28040_, new_n28041_, new_n28042_, new_n28043_, new_n28044_,
    new_n28045_, new_n28046_, new_n28047_, new_n28048_, new_n28049_,
    new_n28050_, new_n28051_, new_n28052_, new_n28053_, new_n28054_,
    new_n28055_, new_n28056_, new_n28057_, new_n28058_, new_n28059_,
    new_n28060_, new_n28061_, new_n28062_, new_n28063_, new_n28064_,
    new_n28065_, new_n28066_, new_n28067_, new_n28068_, new_n28069_,
    new_n28070_, new_n28071_, new_n28072_, new_n28073_, new_n28074_,
    new_n28075_, new_n28076_, new_n28077_, new_n28078_, new_n28079_,
    new_n28080_, new_n28081_, new_n28082_, new_n28083_, new_n28084_,
    new_n28085_, new_n28086_, new_n28087_, new_n28088_, new_n28089_,
    new_n28090_, new_n28091_, new_n28092_, new_n28093_, new_n28094_,
    new_n28095_, new_n28096_, new_n28097_, new_n28098_, new_n28099_,
    new_n28100_, new_n28101_, new_n28102_, new_n28103_, new_n28104_,
    new_n28105_, new_n28106_, new_n28107_, new_n28108_, new_n28109_,
    new_n28110_, new_n28111_, new_n28112_, new_n28113_, new_n28114_,
    new_n28115_, new_n28116_, new_n28117_, new_n28118_, new_n28119_,
    new_n28120_, new_n28121_, new_n28122_, new_n28123_, new_n28124_,
    new_n28125_, new_n28126_, new_n28127_, new_n28128_, new_n28129_,
    new_n28130_, new_n28131_, new_n28132_, new_n28133_, new_n28134_,
    new_n28135_, new_n28136_, new_n28137_, new_n28138_, new_n28139_,
    new_n28140_, new_n28141_, new_n28142_, new_n28143_, new_n28144_,
    new_n28145_, new_n28146_, new_n28147_, new_n28148_, new_n28149_,
    new_n28150_, new_n28151_, new_n28152_, new_n28153_, new_n28154_,
    new_n28155_, new_n28156_, new_n28157_, new_n28158_, new_n28159_,
    new_n28160_, new_n28161_, new_n28162_, new_n28163_, new_n28164_,
    new_n28165_, new_n28166_, new_n28167_, new_n28168_, new_n28169_,
    new_n28170_, new_n28171_, new_n28172_, new_n28173_, new_n28174_,
    new_n28175_, new_n28176_, new_n28177_, new_n28178_, new_n28179_,
    new_n28180_, new_n28181_, new_n28182_, new_n28183_, new_n28184_,
    new_n28185_, new_n28186_, new_n28187_, new_n28188_, new_n28189_,
    new_n28190_, new_n28191_, new_n28192_, new_n28193_, new_n28194_,
    new_n28195_, new_n28196_, new_n28197_, new_n28198_, new_n28199_,
    new_n28200_, new_n28201_, new_n28202_, new_n28203_, new_n28204_,
    new_n28205_, new_n28206_, new_n28207_, new_n28208_, new_n28209_,
    new_n28210_, new_n28211_, new_n28212_, new_n28213_, new_n28214_,
    new_n28215_, new_n28216_, new_n28217_, new_n28218_, new_n28219_,
    new_n28220_, new_n28221_, new_n28222_, new_n28223_, new_n28224_,
    new_n28225_, new_n28226_, new_n28227_, new_n28228_, new_n28229_,
    new_n28230_, new_n28231_, new_n28232_, new_n28233_, new_n28234_,
    new_n28235_, new_n28236_, new_n28237_, new_n28238_, new_n28239_,
    new_n28240_, new_n28241_, new_n28242_, new_n28243_, new_n28244_,
    new_n28245_, new_n28246_, new_n28247_, new_n28248_, new_n28249_,
    new_n28250_, new_n28251_, new_n28252_, new_n28253_, new_n28254_,
    new_n28255_, new_n28256_, new_n28257_, new_n28258_, new_n28259_,
    new_n28260_, new_n28261_, new_n28262_, new_n28263_, new_n28264_,
    new_n28265_, new_n28266_, new_n28267_, new_n28268_, new_n28269_,
    new_n28270_, new_n28271_, new_n28272_, new_n28273_, new_n28274_,
    new_n28275_, new_n28276_, new_n28277_, new_n28278_, new_n28279_,
    new_n28280_, new_n28281_, new_n28282_, new_n28283_, new_n28284_,
    new_n28285_, new_n28286_, new_n28287_, new_n28288_, new_n28289_,
    new_n28290_, new_n28291_, new_n28292_, new_n28293_, new_n28294_,
    new_n28295_, new_n28296_, new_n28297_, new_n28298_, new_n28299_,
    new_n28300_, new_n28301_, new_n28302_, new_n28303_, new_n28304_,
    new_n28305_, new_n28306_, new_n28307_, new_n28308_, new_n28309_,
    new_n28310_, new_n28311_, new_n28312_, new_n28313_, new_n28314_,
    new_n28315_, new_n28316_, new_n28317_, new_n28318_, new_n28319_,
    new_n28320_, new_n28321_, new_n28322_, new_n28323_, new_n28324_,
    new_n28325_, new_n28326_, new_n28327_, new_n28328_, new_n28329_,
    new_n28330_, new_n28331_, new_n28332_, new_n28333_, new_n28334_,
    new_n28335_, new_n28336_, new_n28337_, new_n28338_, new_n28339_,
    new_n28340_, new_n28341_, new_n28342_, new_n28343_, new_n28344_,
    new_n28345_, new_n28346_, new_n28347_, new_n28348_, new_n28349_,
    new_n28350_, new_n28351_, new_n28352_, new_n28353_, new_n28354_,
    new_n28355_, new_n28356_, new_n28357_, new_n28358_, new_n28359_,
    new_n28360_, new_n28361_, new_n28362_, new_n28363_, new_n28364_,
    new_n28365_, new_n28366_, new_n28367_, new_n28368_, new_n28369_,
    new_n28370_, new_n28371_, new_n28372_, new_n28373_, new_n28374_,
    new_n28375_, new_n28376_, new_n28377_, new_n28378_, new_n28379_,
    new_n28380_, new_n28381_, new_n28382_, new_n28383_, new_n28384_,
    new_n28385_, new_n28386_, new_n28387_, new_n28388_, new_n28389_,
    new_n28390_, new_n28391_, new_n28392_, new_n28393_, new_n28394_,
    new_n28395_, new_n28396_, new_n28397_, new_n28398_, new_n28399_,
    new_n28400_, new_n28401_, new_n28402_, new_n28403_, new_n28404_,
    new_n28405_, new_n28406_, new_n28407_, new_n28408_, new_n28409_,
    new_n28410_, new_n28411_, new_n28412_, new_n28413_, new_n28414_,
    new_n28415_, new_n28416_, new_n28417_, new_n28418_, new_n28419_,
    new_n28420_, new_n28421_, new_n28422_, new_n28423_, new_n28424_,
    new_n28425_, new_n28426_, new_n28427_, new_n28428_, new_n28429_,
    new_n28430_, new_n28431_, new_n28432_, new_n28433_, new_n28434_,
    new_n28435_, new_n28436_, new_n28437_, new_n28438_, new_n28439_,
    new_n28440_, new_n28441_, new_n28443_, new_n28444_, new_n28445_,
    new_n28446_, new_n28447_, new_n28448_, new_n28449_, new_n28450_,
    new_n28451_, new_n28452_, new_n28453_, new_n28454_, new_n28455_,
    new_n28456_, new_n28457_, new_n28458_, new_n28459_, new_n28460_,
    new_n28461_, new_n28462_, new_n28463_, new_n28464_, new_n28465_,
    new_n28466_, new_n28467_, new_n28468_, new_n28469_, new_n28470_,
    new_n28471_, new_n28472_, new_n28473_, new_n28474_, new_n28475_,
    new_n28476_, new_n28477_, new_n28478_, new_n28479_, new_n28480_,
    new_n28481_, new_n28482_, new_n28483_, new_n28484_, new_n28485_,
    new_n28486_, new_n28487_, new_n28488_, new_n28489_, new_n28490_,
    new_n28491_, new_n28492_, new_n28493_, new_n28494_, new_n28495_,
    new_n28496_, new_n28497_, new_n28498_, new_n28499_, new_n28500_,
    new_n28501_, new_n28502_, new_n28503_, new_n28504_, new_n28505_,
    new_n28506_, new_n28507_, new_n28508_, new_n28509_, new_n28510_,
    new_n28511_, new_n28512_, new_n28513_, new_n28514_, new_n28515_,
    new_n28516_, new_n28517_, new_n28518_, new_n28519_, new_n28520_,
    new_n28521_, new_n28522_, new_n28523_, new_n28524_, new_n28525_,
    new_n28526_, new_n28527_, new_n28528_, new_n28529_, new_n28530_,
    new_n28531_, new_n28532_, new_n28533_, new_n28534_, new_n28535_,
    new_n28536_, new_n28537_, new_n28538_, new_n28539_, new_n28540_,
    new_n28541_, new_n28542_, new_n28543_, new_n28544_, new_n28545_,
    new_n28546_, new_n28547_, new_n28548_, new_n28549_, new_n28550_,
    new_n28551_, new_n28552_, new_n28553_, new_n28554_, new_n28555_,
    new_n28556_, new_n28557_, new_n28558_, new_n28559_, new_n28560_,
    new_n28561_, new_n28562_, new_n28563_, new_n28564_, new_n28565_,
    new_n28566_, new_n28567_, new_n28568_, new_n28569_, new_n28570_,
    new_n28571_, new_n28572_, new_n28573_, new_n28574_, new_n28575_,
    new_n28576_, new_n28577_, new_n28578_, new_n28579_, new_n28580_,
    new_n28581_, new_n28582_, new_n28583_, new_n28584_, new_n28585_,
    new_n28586_, new_n28587_, new_n28588_, new_n28589_, new_n28590_,
    new_n28591_, new_n28592_, new_n28593_, new_n28594_, new_n28595_,
    new_n28596_, new_n28597_, new_n28598_, new_n28599_, new_n28600_,
    new_n28601_, new_n28602_, new_n28603_, new_n28604_, new_n28605_,
    new_n28606_, new_n28607_, new_n28608_, new_n28609_, new_n28610_,
    new_n28611_, new_n28612_, new_n28613_, new_n28614_, new_n28615_,
    new_n28616_, new_n28617_, new_n28618_, new_n28619_, new_n28620_,
    new_n28621_, new_n28622_, new_n28623_, new_n28624_, new_n28625_,
    new_n28626_, new_n28627_, new_n28628_, new_n28629_, new_n28630_,
    new_n28631_, new_n28632_, new_n28633_, new_n28634_, new_n28635_,
    new_n28636_, new_n28637_, new_n28638_, new_n28639_, new_n28640_,
    new_n28641_, new_n28642_, new_n28643_, new_n28644_, new_n28645_,
    new_n28646_, new_n28647_, new_n28648_, new_n28649_, new_n28650_,
    new_n28651_, new_n28652_, new_n28653_, new_n28654_, new_n28655_,
    new_n28656_, new_n28657_, new_n28658_, new_n28659_, new_n28660_,
    new_n28661_, new_n28662_, new_n28663_, new_n28664_, new_n28665_,
    new_n28666_, new_n28667_, new_n28668_, new_n28669_, new_n28670_,
    new_n28671_, new_n28672_, new_n28673_, new_n28674_, new_n28675_,
    new_n28676_, new_n28677_, new_n28678_, new_n28679_, new_n28680_,
    new_n28681_, new_n28682_, new_n28683_, new_n28684_, new_n28685_,
    new_n28686_, new_n28687_, new_n28688_, new_n28689_, new_n28690_,
    new_n28691_, new_n28692_, new_n28693_, new_n28694_, new_n28695_,
    new_n28696_, new_n28697_, new_n28698_, new_n28699_, new_n28700_,
    new_n28701_, new_n28702_, new_n28703_, new_n28704_, new_n28705_,
    new_n28706_, new_n28707_, new_n28708_, new_n28709_, new_n28710_,
    new_n28711_, new_n28712_, new_n28713_, new_n28714_, new_n28715_,
    new_n28716_, new_n28717_, new_n28718_, new_n28719_, new_n28720_,
    new_n28721_, new_n28722_, new_n28723_, new_n28724_, new_n28725_,
    new_n28726_, new_n28727_, new_n28728_, new_n28729_, new_n28730_,
    new_n28731_, new_n28732_, new_n28733_, new_n28734_, new_n28735_,
    new_n28736_, new_n28737_, new_n28738_, new_n28739_, new_n28740_,
    new_n28741_, new_n28742_, new_n28743_, new_n28744_, new_n28745_,
    new_n28746_, new_n28747_, new_n28748_, new_n28749_, new_n28750_,
    new_n28751_, new_n28752_, new_n28753_, new_n28754_, new_n28755_,
    new_n28756_, new_n28757_, new_n28758_, new_n28759_, new_n28760_,
    new_n28761_, new_n28762_, new_n28763_, new_n28764_, new_n28765_,
    new_n28766_, new_n28767_, new_n28768_, new_n28769_, new_n28770_,
    new_n28771_, new_n28772_, new_n28773_, new_n28774_, new_n28775_,
    new_n28776_, new_n28777_, new_n28778_, new_n28779_, new_n28780_,
    new_n28781_, new_n28782_, new_n28783_, new_n28784_, new_n28785_,
    new_n28786_, new_n28787_, new_n28788_, new_n28789_, new_n28790_,
    new_n28791_, new_n28792_, new_n28793_, new_n28794_, new_n28795_,
    new_n28796_, new_n28797_, new_n28798_, new_n28799_, new_n28800_,
    new_n28801_, new_n28802_, new_n28803_, new_n28804_, new_n28805_,
    new_n28806_, new_n28807_, new_n28808_, new_n28809_, new_n28810_,
    new_n28811_, new_n28812_, new_n28813_, new_n28814_, new_n28815_,
    new_n28816_, new_n28817_, new_n28818_, new_n28819_, new_n28820_,
    new_n28821_, new_n28822_, new_n28823_, new_n28824_, new_n28825_,
    new_n28826_, new_n28827_, new_n28828_, new_n28829_, new_n28830_,
    new_n28831_, new_n28832_, new_n28833_, new_n28834_, new_n28835_,
    new_n28836_, new_n28837_, new_n28838_, new_n28839_, new_n28840_,
    new_n28841_, new_n28842_, new_n28843_, new_n28844_, new_n28845_,
    new_n28846_, new_n28847_, new_n28848_, new_n28849_, new_n28850_,
    new_n28851_, new_n28852_, new_n28853_, new_n28854_, new_n28855_,
    new_n28856_, new_n28857_, new_n28858_, new_n28859_, new_n28860_,
    new_n28861_, new_n28862_, new_n28863_, new_n28864_, new_n28865_,
    new_n28866_, new_n28867_, new_n28868_, new_n28869_, new_n28870_,
    new_n28871_, new_n28872_, new_n28873_, new_n28874_, new_n28875_,
    new_n28876_, new_n28877_, new_n28878_, new_n28879_, new_n28880_,
    new_n28881_, new_n28882_, new_n28883_, new_n28884_, new_n28885_,
    new_n28886_, new_n28887_, new_n28888_, new_n28889_, new_n28890_,
    new_n28891_, new_n28892_, new_n28893_, new_n28894_, new_n28895_,
    new_n28896_, new_n28897_, new_n28898_, new_n28899_, new_n28900_,
    new_n28901_, new_n28902_, new_n28903_, new_n28904_, new_n28905_,
    new_n28906_, new_n28907_, new_n28908_, new_n28909_, new_n28910_,
    new_n28911_, new_n28912_, new_n28913_, new_n28914_, new_n28915_,
    new_n28916_, new_n28917_, new_n28918_, new_n28920_, new_n28921_,
    new_n28922_, new_n28923_, new_n28924_, new_n28925_, new_n28926_,
    new_n28927_, new_n28928_, new_n28929_, new_n28930_, new_n28931_,
    new_n28932_, new_n28933_, new_n28934_, new_n28935_, new_n28936_,
    new_n28937_, new_n28938_, new_n28939_, new_n28940_, new_n28941_,
    new_n28942_, new_n28943_, new_n28944_, new_n28945_, new_n28946_,
    new_n28947_, new_n28948_, new_n28949_, new_n28950_, new_n28951_,
    new_n28952_, new_n28953_, new_n28954_, new_n28955_, new_n28956_,
    new_n28957_, new_n28958_, new_n28959_, new_n28960_, new_n28961_,
    new_n28962_, new_n28963_, new_n28964_, new_n28965_, new_n28966_,
    new_n28967_, new_n28968_, new_n28969_, new_n28970_, new_n28971_,
    new_n28972_, new_n28973_, new_n28974_, new_n28975_, new_n28976_,
    new_n28977_, new_n28978_, new_n28979_, new_n28980_, new_n28981_,
    new_n28982_, new_n28983_, new_n28984_, new_n28985_, new_n28986_,
    new_n28987_, new_n28988_, new_n28989_, new_n28990_, new_n28991_,
    new_n28992_, new_n28993_, new_n28994_, new_n28995_, new_n28996_,
    new_n28997_, new_n28998_, new_n28999_, new_n29000_, new_n29001_,
    new_n29002_, new_n29003_, new_n29004_, new_n29005_, new_n29006_,
    new_n29007_, new_n29008_, new_n29009_, new_n29010_, new_n29011_,
    new_n29012_, new_n29013_, new_n29014_, new_n29015_, new_n29016_,
    new_n29017_, new_n29018_, new_n29019_, new_n29020_, new_n29021_,
    new_n29022_, new_n29023_, new_n29024_, new_n29025_, new_n29026_,
    new_n29027_, new_n29028_, new_n29029_, new_n29030_, new_n29031_,
    new_n29032_, new_n29033_, new_n29034_, new_n29035_, new_n29036_,
    new_n29037_, new_n29038_, new_n29039_, new_n29040_, new_n29041_,
    new_n29042_, new_n29043_, new_n29044_, new_n29045_, new_n29046_,
    new_n29047_, new_n29048_, new_n29049_, new_n29050_, new_n29051_,
    new_n29052_, new_n29053_, new_n29054_, new_n29055_, new_n29056_,
    new_n29057_, new_n29058_, new_n29059_, new_n29060_, new_n29061_,
    new_n29062_, new_n29063_, new_n29064_, new_n29065_, new_n29066_,
    new_n29067_, new_n29068_, new_n29069_, new_n29070_, new_n29071_,
    new_n29072_, new_n29073_, new_n29074_, new_n29075_, new_n29076_,
    new_n29077_, new_n29078_, new_n29079_, new_n29080_, new_n29081_,
    new_n29082_, new_n29083_, new_n29084_, new_n29085_, new_n29086_,
    new_n29087_, new_n29088_, new_n29089_, new_n29090_, new_n29091_,
    new_n29092_, new_n29093_, new_n29094_, new_n29095_, new_n29096_,
    new_n29097_, new_n29098_, new_n29099_, new_n29100_, new_n29101_,
    new_n29102_, new_n29103_, new_n29104_, new_n29105_, new_n29106_,
    new_n29107_, new_n29108_, new_n29109_, new_n29110_, new_n29111_,
    new_n29112_, new_n29113_, new_n29114_, new_n29115_, new_n29116_,
    new_n29117_, new_n29118_, new_n29119_, new_n29120_, new_n29121_,
    new_n29122_, new_n29123_, new_n29124_, new_n29125_, new_n29126_,
    new_n29127_, new_n29128_, new_n29129_, new_n29130_, new_n29131_,
    new_n29132_, new_n29133_, new_n29134_, new_n29135_, new_n29136_,
    new_n29137_, new_n29138_, new_n29139_, new_n29140_, new_n29141_,
    new_n29142_, new_n29143_, new_n29144_, new_n29145_, new_n29146_,
    new_n29147_, new_n29148_, new_n29149_, new_n29150_, new_n29151_,
    new_n29152_, new_n29153_, new_n29154_, new_n29155_, new_n29156_,
    new_n29157_, new_n29158_, new_n29159_, new_n29160_, new_n29161_,
    new_n29162_, new_n29163_, new_n29164_, new_n29165_, new_n29166_,
    new_n29167_, new_n29168_, new_n29169_, new_n29170_, new_n29171_,
    new_n29172_, new_n29173_, new_n29174_, new_n29175_, new_n29176_,
    new_n29177_, new_n29178_, new_n29179_, new_n29180_, new_n29181_,
    new_n29182_, new_n29183_, new_n29184_, new_n29185_, new_n29186_,
    new_n29187_, new_n29188_, new_n29189_, new_n29190_, new_n29191_,
    new_n29192_, new_n29193_, new_n29194_, new_n29195_, new_n29196_,
    new_n29197_, new_n29198_, new_n29199_, new_n29200_, new_n29201_,
    new_n29202_, new_n29203_, new_n29204_, new_n29205_, new_n29206_,
    new_n29207_, new_n29208_, new_n29209_, new_n29210_, new_n29211_,
    new_n29212_, new_n29213_, new_n29214_, new_n29215_, new_n29216_,
    new_n29217_, new_n29218_, new_n29219_, new_n29220_, new_n29221_,
    new_n29222_, new_n29223_, new_n29224_, new_n29225_, new_n29226_,
    new_n29227_, new_n29228_, new_n29229_, new_n29230_, new_n29231_,
    new_n29232_, new_n29233_, new_n29234_, new_n29235_, new_n29236_,
    new_n29237_, new_n29238_, new_n29239_, new_n29240_, new_n29241_,
    new_n29242_, new_n29243_, new_n29244_, new_n29245_, new_n29246_,
    new_n29247_, new_n29248_, new_n29249_, new_n29250_, new_n29251_,
    new_n29252_, new_n29253_, new_n29254_, new_n29255_, new_n29256_,
    new_n29257_, new_n29258_, new_n29259_, new_n29260_, new_n29261_,
    new_n29262_, new_n29263_, new_n29264_, new_n29265_, new_n29266_,
    new_n29267_, new_n29268_, new_n29269_, new_n29270_, new_n29271_,
    new_n29272_, new_n29273_, new_n29274_, new_n29275_, new_n29276_,
    new_n29277_, new_n29278_, new_n29279_, new_n29280_, new_n29281_,
    new_n29282_, new_n29283_, new_n29284_, new_n29285_, new_n29286_,
    new_n29287_, new_n29288_, new_n29289_, new_n29290_, new_n29291_,
    new_n29292_, new_n29293_, new_n29294_, new_n29295_, new_n29296_,
    new_n29297_, new_n29298_, new_n29299_, new_n29300_, new_n29301_,
    new_n29302_, new_n29303_, new_n29304_, new_n29305_, new_n29306_,
    new_n29307_, new_n29308_, new_n29309_, new_n29310_, new_n29311_,
    new_n29312_, new_n29313_, new_n29314_, new_n29315_, new_n29316_,
    new_n29317_, new_n29318_, new_n29319_, new_n29320_, new_n29321_,
    new_n29322_, new_n29323_, new_n29324_, new_n29325_, new_n29326_,
    new_n29327_, new_n29328_, new_n29329_, new_n29330_, new_n29331_,
    new_n29332_, new_n29333_, new_n29334_, new_n29335_, new_n29336_,
    new_n29337_, new_n29338_, new_n29339_, new_n29340_, new_n29341_,
    new_n29342_, new_n29343_, new_n29344_, new_n29345_, new_n29346_,
    new_n29347_, new_n29348_, new_n29349_, new_n29350_, new_n29351_,
    new_n29352_, new_n29353_, new_n29354_, new_n29355_, new_n29356_,
    new_n29357_, new_n29358_, new_n29359_, new_n29360_, new_n29361_,
    new_n29362_, new_n29363_, new_n29364_, new_n29365_, new_n29366_,
    new_n29367_, new_n29368_, new_n29369_, new_n29370_, new_n29371_,
    new_n29372_, new_n29373_, new_n29374_, new_n29375_, new_n29376_,
    new_n29377_, new_n29378_, new_n29379_, new_n29380_, new_n29381_,
    new_n29382_, new_n29383_, new_n29384_, new_n29385_, new_n29386_,
    new_n29387_, new_n29388_, new_n29389_, new_n29390_, new_n29391_,
    new_n29392_, new_n29393_, new_n29395_, new_n29396_, new_n29397_,
    new_n29398_, new_n29399_, new_n29400_, new_n29401_, new_n29402_,
    new_n29403_, new_n29404_, new_n29405_, new_n29406_, new_n29407_,
    new_n29408_, new_n29409_, new_n29410_, new_n29411_, new_n29412_,
    new_n29413_, new_n29414_, new_n29415_, new_n29416_, new_n29417_,
    new_n29418_, new_n29419_, new_n29420_, new_n29421_, new_n29422_,
    new_n29423_, new_n29424_, new_n29425_, new_n29426_, new_n29427_,
    new_n29428_, new_n29429_, new_n29430_, new_n29431_, new_n29432_,
    new_n29433_, new_n29434_, new_n29435_, new_n29436_, new_n29437_,
    new_n29438_, new_n29439_, new_n29440_, new_n29441_, new_n29442_,
    new_n29443_, new_n29444_, new_n29445_, new_n29446_, new_n29447_,
    new_n29448_, new_n29449_, new_n29450_, new_n29451_, new_n29452_,
    new_n29453_, new_n29454_, new_n29455_, new_n29456_, new_n29457_,
    new_n29458_, new_n29459_, new_n29460_, new_n29461_, new_n29462_,
    new_n29463_, new_n29464_, new_n29465_, new_n29466_, new_n29467_,
    new_n29468_, new_n29469_, new_n29470_, new_n29471_, new_n29472_,
    new_n29473_, new_n29474_, new_n29475_, new_n29476_, new_n29477_,
    new_n29478_, new_n29479_, new_n29480_, new_n29481_, new_n29482_,
    new_n29483_, new_n29484_, new_n29485_, new_n29486_, new_n29487_,
    new_n29488_, new_n29489_, new_n29490_, new_n29491_, new_n29492_,
    new_n29493_, new_n29494_, new_n29495_, new_n29496_, new_n29497_,
    new_n29498_, new_n29499_, new_n29500_, new_n29501_, new_n29502_,
    new_n29503_, new_n29504_, new_n29505_, new_n29506_, new_n29507_,
    new_n29508_, new_n29509_, new_n29510_, new_n29511_, new_n29512_,
    new_n29513_, new_n29514_, new_n29515_, new_n29516_, new_n29517_,
    new_n29518_, new_n29519_, new_n29520_, new_n29521_, new_n29522_,
    new_n29523_, new_n29524_, new_n29525_, new_n29526_, new_n29527_,
    new_n29528_, new_n29529_, new_n29530_, new_n29531_, new_n29532_,
    new_n29533_, new_n29534_, new_n29535_, new_n29536_, new_n29537_,
    new_n29538_, new_n29539_, new_n29540_, new_n29541_, new_n29542_,
    new_n29543_, new_n29544_, new_n29545_, new_n29546_, new_n29547_,
    new_n29548_, new_n29549_, new_n29550_, new_n29551_, new_n29552_,
    new_n29553_, new_n29554_, new_n29555_, new_n29556_, new_n29557_,
    new_n29558_, new_n29559_, new_n29560_, new_n29561_, new_n29562_,
    new_n29563_, new_n29564_, new_n29565_, new_n29566_, new_n29567_,
    new_n29568_, new_n29569_, new_n29570_, new_n29571_, new_n29572_,
    new_n29573_, new_n29574_, new_n29575_, new_n29576_, new_n29577_,
    new_n29578_, new_n29579_, new_n29580_, new_n29581_, new_n29582_,
    new_n29583_, new_n29584_, new_n29585_, new_n29586_, new_n29587_,
    new_n29588_, new_n29589_, new_n29590_, new_n29591_, new_n29592_,
    new_n29593_, new_n29594_, new_n29595_, new_n29596_, new_n29597_,
    new_n29598_, new_n29599_, new_n29600_, new_n29601_, new_n29602_,
    new_n29603_, new_n29604_, new_n29605_, new_n29606_, new_n29607_,
    new_n29608_, new_n29609_, new_n29610_, new_n29611_, new_n29612_,
    new_n29613_, new_n29614_, new_n29615_, new_n29616_, new_n29617_,
    new_n29618_, new_n29619_, new_n29620_, new_n29621_, new_n29622_,
    new_n29623_, new_n29624_, new_n29625_, new_n29626_, new_n29627_,
    new_n29628_, new_n29629_, new_n29630_, new_n29631_, new_n29632_,
    new_n29633_, new_n29634_, new_n29635_, new_n29636_, new_n29637_,
    new_n29638_, new_n29639_, new_n29640_, new_n29641_, new_n29642_,
    new_n29643_, new_n29644_, new_n29645_, new_n29646_, new_n29647_,
    new_n29648_, new_n29649_, new_n29650_, new_n29651_, new_n29652_,
    new_n29653_, new_n29654_, new_n29655_, new_n29656_, new_n29657_,
    new_n29658_, new_n29659_, new_n29660_, new_n29661_, new_n29662_,
    new_n29663_, new_n29664_, new_n29665_, new_n29666_, new_n29667_,
    new_n29668_, new_n29669_, new_n29670_, new_n29671_, new_n29672_,
    new_n29673_, new_n29674_, new_n29675_, new_n29676_, new_n29677_,
    new_n29678_, new_n29679_, new_n29680_, new_n29681_, new_n29682_,
    new_n29683_, new_n29684_, new_n29685_, new_n29686_, new_n29687_,
    new_n29688_, new_n29689_, new_n29690_, new_n29691_, new_n29692_,
    new_n29693_, new_n29694_, new_n29695_, new_n29696_, new_n29697_,
    new_n29698_, new_n29699_, new_n29700_, new_n29701_, new_n29702_,
    new_n29703_, new_n29704_, new_n29705_, new_n29706_, new_n29707_,
    new_n29708_, new_n29709_, new_n29710_, new_n29711_, new_n29712_,
    new_n29713_, new_n29714_, new_n29715_, new_n29716_, new_n29717_,
    new_n29718_, new_n29719_, new_n29720_, new_n29721_, new_n29722_,
    new_n29723_, new_n29724_, new_n29725_, new_n29726_, new_n29727_,
    new_n29728_, new_n29729_, new_n29730_, new_n29731_, new_n29732_,
    new_n29733_, new_n29734_, new_n29735_, new_n29736_, new_n29737_,
    new_n29738_, new_n29739_, new_n29740_, new_n29741_, new_n29742_,
    new_n29743_, new_n29744_, new_n29745_, new_n29746_, new_n29747_,
    new_n29748_, new_n29749_, new_n29750_, new_n29751_, new_n29752_,
    new_n29753_, new_n29754_, new_n29755_, new_n29756_, new_n29757_,
    new_n29758_, new_n29759_, new_n29760_, new_n29761_, new_n29762_,
    new_n29763_, new_n29764_, new_n29765_, new_n29766_, new_n29767_,
    new_n29768_, new_n29769_, new_n29770_, new_n29771_, new_n29772_,
    new_n29773_, new_n29774_, new_n29775_, new_n29776_, new_n29777_,
    new_n29778_, new_n29779_, new_n29780_, new_n29781_, new_n29782_,
    new_n29783_, new_n29784_, new_n29785_, new_n29786_, new_n29787_,
    new_n29788_, new_n29789_, new_n29790_, new_n29791_, new_n29792_,
    new_n29793_, new_n29794_, new_n29795_, new_n29796_, new_n29797_,
    new_n29798_, new_n29799_, new_n29800_, new_n29801_, new_n29802_,
    new_n29803_, new_n29804_, new_n29805_, new_n29806_, new_n29807_,
    new_n29808_, new_n29809_, new_n29810_, new_n29811_, new_n29812_,
    new_n29813_, new_n29814_, new_n29815_, new_n29816_, new_n29817_,
    new_n29818_, new_n29819_, new_n29820_, new_n29821_, new_n29822_,
    new_n29823_, new_n29824_, new_n29825_, new_n29826_, new_n29827_,
    new_n29828_, new_n29829_, new_n29830_, new_n29831_, new_n29832_,
    new_n29833_, new_n29834_, new_n29835_, new_n29836_, new_n29837_,
    new_n29838_, new_n29839_, new_n29840_, new_n29841_, new_n29842_,
    new_n29843_, new_n29844_, new_n29845_, new_n29846_, new_n29847_,
    new_n29848_, new_n29849_, new_n29850_, new_n29851_, new_n29852_,
    new_n29853_, new_n29854_, new_n29855_, new_n29856_, new_n29857_,
    new_n29858_, new_n29859_, new_n29860_, new_n29861_, new_n29862_,
    new_n29863_, new_n29864_, new_n29865_, new_n29866_, new_n29867_,
    new_n29868_, new_n29870_, new_n29871_, new_n29872_, new_n29873_,
    new_n29874_, new_n29875_, new_n29876_, new_n29877_, new_n29878_,
    new_n29879_, new_n29880_, new_n29881_, new_n29882_, new_n29883_,
    new_n29884_, new_n29885_, new_n29886_, new_n29887_, new_n29888_,
    new_n29889_, new_n29890_, new_n29891_, new_n29892_, new_n29893_,
    new_n29894_, new_n29895_, new_n29896_, new_n29897_, new_n29898_,
    new_n29899_, new_n29900_, new_n29901_, new_n29902_, new_n29903_,
    new_n29904_, new_n29905_, new_n29906_, new_n29907_, new_n29908_,
    new_n29909_, new_n29910_, new_n29911_, new_n29912_, new_n29913_,
    new_n29914_, new_n29915_, new_n29916_, new_n29917_, new_n29918_,
    new_n29919_, new_n29920_, new_n29921_, new_n29922_, new_n29923_,
    new_n29924_, new_n29925_, new_n29926_, new_n29927_, new_n29928_,
    new_n29929_, new_n29930_, new_n29931_, new_n29932_, new_n29933_,
    new_n29934_, new_n29935_, new_n29936_, new_n29937_, new_n29938_,
    new_n29939_, new_n29940_, new_n29941_, new_n29942_, new_n29943_,
    new_n29944_, new_n29945_, new_n29946_, new_n29947_, new_n29948_,
    new_n29949_, new_n29950_, new_n29951_, new_n29952_, new_n29953_,
    new_n29954_, new_n29955_, new_n29956_, new_n29957_, new_n29958_,
    new_n29959_, new_n29960_, new_n29961_, new_n29962_, new_n29963_,
    new_n29964_, new_n29965_, new_n29966_, new_n29967_, new_n29968_,
    new_n29969_, new_n29970_, new_n29971_, new_n29972_, new_n29973_,
    new_n29974_, new_n29975_, new_n29976_, new_n29977_, new_n29978_,
    new_n29979_, new_n29980_, new_n29981_, new_n29982_, new_n29983_,
    new_n29984_, new_n29985_, new_n29986_, new_n29987_, new_n29988_,
    new_n29989_, new_n29990_, new_n29991_, new_n29992_, new_n29993_,
    new_n29994_, new_n29995_, new_n29996_, new_n29997_, new_n29998_,
    new_n29999_, new_n30000_, new_n30001_, new_n30002_, new_n30003_,
    new_n30004_, new_n30005_, new_n30006_, new_n30007_, new_n30008_,
    new_n30009_, new_n30010_, new_n30011_, new_n30012_, new_n30013_,
    new_n30014_, new_n30015_, new_n30016_, new_n30017_, new_n30018_,
    new_n30019_, new_n30020_, new_n30021_, new_n30022_, new_n30023_,
    new_n30024_, new_n30025_, new_n30026_, new_n30027_, new_n30028_,
    new_n30029_, new_n30030_, new_n30031_, new_n30032_, new_n30033_,
    new_n30034_, new_n30035_, new_n30036_, new_n30037_, new_n30038_,
    new_n30039_, new_n30040_, new_n30041_, new_n30042_, new_n30043_,
    new_n30044_, new_n30045_, new_n30046_, new_n30047_, new_n30048_,
    new_n30049_, new_n30050_, new_n30051_, new_n30052_, new_n30053_,
    new_n30054_, new_n30055_, new_n30056_, new_n30057_, new_n30058_,
    new_n30059_, new_n30060_, new_n30061_, new_n30062_, new_n30063_,
    new_n30064_, new_n30065_, new_n30066_, new_n30067_, new_n30068_,
    new_n30069_, new_n30070_, new_n30071_, new_n30072_, new_n30073_,
    new_n30074_, new_n30075_, new_n30076_, new_n30077_, new_n30078_,
    new_n30079_, new_n30080_, new_n30081_, new_n30082_, new_n30083_,
    new_n30084_, new_n30085_, new_n30086_, new_n30087_, new_n30088_,
    new_n30089_, new_n30090_, new_n30091_, new_n30092_, new_n30093_,
    new_n30094_, new_n30095_, new_n30096_, new_n30097_, new_n30098_,
    new_n30099_, new_n30100_, new_n30101_, new_n30102_, new_n30103_,
    new_n30104_, new_n30105_, new_n30106_, new_n30107_, new_n30108_,
    new_n30109_, new_n30110_, new_n30111_, new_n30112_, new_n30113_,
    new_n30114_, new_n30115_, new_n30116_, new_n30117_, new_n30118_,
    new_n30119_, new_n30120_, new_n30121_, new_n30122_, new_n30123_,
    new_n30124_, new_n30125_, new_n30126_, new_n30127_, new_n30128_,
    new_n30129_, new_n30130_, new_n30131_, new_n30132_, new_n30133_,
    new_n30134_, new_n30135_, new_n30136_, new_n30137_, new_n30138_,
    new_n30139_, new_n30140_, new_n30141_, new_n30142_, new_n30143_,
    new_n30144_, new_n30145_, new_n30146_, new_n30147_, new_n30148_,
    new_n30149_, new_n30150_, new_n30151_, new_n30152_, new_n30153_,
    new_n30154_, new_n30155_, new_n30156_, new_n30157_, new_n30158_,
    new_n30159_, new_n30160_, new_n30161_, new_n30162_, new_n30163_,
    new_n30164_, new_n30165_, new_n30166_, new_n30167_, new_n30168_,
    new_n30169_, new_n30170_, new_n30171_, new_n30172_, new_n30173_,
    new_n30174_, new_n30175_, new_n30176_, new_n30177_, new_n30178_,
    new_n30179_, new_n30180_, new_n30181_, new_n30182_, new_n30183_,
    new_n30184_, new_n30185_, new_n30186_, new_n30187_, new_n30188_,
    new_n30189_, new_n30190_, new_n30191_, new_n30192_, new_n30193_,
    new_n30194_, new_n30195_, new_n30196_, new_n30197_, new_n30198_,
    new_n30199_, new_n30200_, new_n30201_, new_n30202_, new_n30203_,
    new_n30204_, new_n30205_, new_n30206_, new_n30207_, new_n30208_,
    new_n30209_, new_n30210_, new_n30211_, new_n30212_, new_n30213_,
    new_n30214_, new_n30215_, new_n30216_, new_n30217_, new_n30218_,
    new_n30219_, new_n30220_, new_n30221_, new_n30222_, new_n30223_,
    new_n30224_, new_n30225_, new_n30226_, new_n30227_, new_n30228_,
    new_n30229_, new_n30230_, new_n30231_, new_n30232_, new_n30233_,
    new_n30234_, new_n30235_, new_n30236_, new_n30237_, new_n30238_,
    new_n30239_, new_n30240_, new_n30241_, new_n30242_, new_n30243_,
    new_n30244_, new_n30245_, new_n30246_, new_n30247_, new_n30248_,
    new_n30249_, new_n30250_, new_n30251_, new_n30252_, new_n30253_,
    new_n30254_, new_n30255_, new_n30256_, new_n30257_, new_n30258_,
    new_n30259_, new_n30260_, new_n30261_, new_n30262_, new_n30263_,
    new_n30264_, new_n30265_, new_n30266_, new_n30267_, new_n30268_,
    new_n30269_, new_n30270_, new_n30271_, new_n30272_, new_n30273_,
    new_n30274_, new_n30275_, new_n30276_, new_n30277_, new_n30278_,
    new_n30279_, new_n30280_, new_n30281_, new_n30282_, new_n30283_,
    new_n30284_, new_n30285_, new_n30286_, new_n30287_, new_n30288_,
    new_n30289_, new_n30290_, new_n30291_, new_n30292_, new_n30293_,
    new_n30294_, new_n30295_, new_n30296_, new_n30297_, new_n30298_,
    new_n30299_, new_n30300_, new_n30301_, new_n30302_, new_n30303_,
    new_n30304_, new_n30305_, new_n30306_, new_n30307_, new_n30308_,
    new_n30309_, new_n30310_, new_n30311_, new_n30312_, new_n30313_,
    new_n30314_, new_n30315_, new_n30316_, new_n30317_, new_n30318_,
    new_n30319_, new_n30320_, new_n30321_, new_n30322_, new_n30323_,
    new_n30324_, new_n30325_, new_n30326_, new_n30327_, new_n30328_,
    new_n30329_, new_n30330_, new_n30331_, new_n30332_, new_n30333_,
    new_n30334_, new_n30335_, new_n30336_, new_n30337_, new_n30338_,
    new_n30339_, new_n30340_, new_n30341_, new_n30342_, new_n30343_,
    new_n30345_, new_n30346_, new_n30347_, new_n30348_, new_n30349_,
    new_n30350_, new_n30351_, new_n30352_, new_n30353_, new_n30354_,
    new_n30355_, new_n30356_, new_n30357_, new_n30358_, new_n30359_,
    new_n30360_, new_n30361_, new_n30362_, new_n30363_, new_n30364_,
    new_n30365_, new_n30366_, new_n30367_, new_n30368_, new_n30369_,
    new_n30370_, new_n30371_, new_n30372_, new_n30373_, new_n30374_,
    new_n30375_, new_n30376_, new_n30377_, new_n30378_, new_n30379_,
    new_n30380_, new_n30381_, new_n30382_, new_n30383_, new_n30384_,
    new_n30385_, new_n30386_, new_n30387_, new_n30388_, new_n30389_,
    new_n30390_, new_n30391_, new_n30392_, new_n30393_, new_n30394_,
    new_n30395_, new_n30396_, new_n30397_, new_n30398_, new_n30399_,
    new_n30400_, new_n30401_, new_n30402_, new_n30403_, new_n30404_,
    new_n30405_, new_n30406_, new_n30407_, new_n30408_, new_n30409_,
    new_n30410_, new_n30411_, new_n30412_, new_n30413_, new_n30414_,
    new_n30415_, new_n30416_, new_n30417_, new_n30418_, new_n30419_,
    new_n30420_, new_n30421_, new_n30422_, new_n30423_, new_n30424_,
    new_n30425_, new_n30426_, new_n30427_, new_n30428_, new_n30429_,
    new_n30430_, new_n30431_, new_n30432_, new_n30433_, new_n30434_,
    new_n30435_, new_n30436_, new_n30437_, new_n30438_, new_n30439_,
    new_n30440_, new_n30441_, new_n30442_, new_n30443_, new_n30444_,
    new_n30445_, new_n30446_, new_n30447_, new_n30448_, new_n30449_,
    new_n30450_, new_n30451_, new_n30452_, new_n30453_, new_n30454_,
    new_n30455_, new_n30456_, new_n30457_, new_n30458_, new_n30459_,
    new_n30460_, new_n30461_, new_n30462_, new_n30463_, new_n30464_,
    new_n30465_, new_n30466_, new_n30467_, new_n30468_, new_n30469_,
    new_n30470_, new_n30471_, new_n30472_, new_n30473_, new_n30474_,
    new_n30475_, new_n30476_, new_n30477_, new_n30478_, new_n30479_,
    new_n30480_, new_n30481_, new_n30482_, new_n30483_, new_n30484_,
    new_n30485_, new_n30486_, new_n30487_, new_n30488_, new_n30489_,
    new_n30490_, new_n30491_, new_n30492_, new_n30493_, new_n30494_,
    new_n30495_, new_n30496_, new_n30497_, new_n30498_, new_n30499_,
    new_n30500_, new_n30501_, new_n30502_, new_n30503_, new_n30504_,
    new_n30505_, new_n30506_, new_n30507_, new_n30508_, new_n30509_,
    new_n30510_, new_n30511_, new_n30512_, new_n30513_, new_n30514_,
    new_n30515_, new_n30516_, new_n30517_, new_n30518_, new_n30519_,
    new_n30520_, new_n30521_, new_n30522_, new_n30523_, new_n30524_,
    new_n30525_, new_n30526_, new_n30527_, new_n30528_, new_n30529_,
    new_n30530_, new_n30531_, new_n30532_, new_n30533_, new_n30534_,
    new_n30535_, new_n30536_, new_n30537_, new_n30538_, new_n30539_,
    new_n30540_, new_n30541_, new_n30542_, new_n30543_, new_n30544_,
    new_n30545_, new_n30546_, new_n30547_, new_n30548_, new_n30549_,
    new_n30550_, new_n30551_, new_n30552_, new_n30553_, new_n30554_,
    new_n30555_, new_n30556_, new_n30557_, new_n30558_, new_n30559_,
    new_n30560_, new_n30561_, new_n30562_, new_n30563_, new_n30564_,
    new_n30565_, new_n30566_, new_n30567_, new_n30568_, new_n30569_,
    new_n30570_, new_n30571_, new_n30572_, new_n30573_, new_n30574_,
    new_n30575_, new_n30576_, new_n30577_, new_n30578_, new_n30579_,
    new_n30580_, new_n30581_, new_n30582_, new_n30583_, new_n30584_,
    new_n30585_, new_n30586_, new_n30587_, new_n30588_, new_n30589_,
    new_n30590_, new_n30591_, new_n30592_, new_n30593_, new_n30594_,
    new_n30595_, new_n30596_, new_n30597_, new_n30598_, new_n30599_,
    new_n30600_, new_n30601_, new_n30602_, new_n30603_, new_n30604_,
    new_n30605_, new_n30606_, new_n30607_, new_n30608_, new_n30609_,
    new_n30610_, new_n30611_, new_n30612_, new_n30613_, new_n30614_,
    new_n30615_, new_n30616_, new_n30617_, new_n30618_, new_n30619_,
    new_n30620_, new_n30621_, new_n30622_, new_n30623_, new_n30624_,
    new_n30625_, new_n30626_, new_n30627_, new_n30628_, new_n30629_,
    new_n30630_, new_n30631_, new_n30632_, new_n30633_, new_n30634_,
    new_n30635_, new_n30636_, new_n30637_, new_n30638_, new_n30639_,
    new_n30640_, new_n30641_, new_n30642_, new_n30643_, new_n30644_,
    new_n30645_, new_n30646_, new_n30647_, new_n30648_, new_n30649_,
    new_n30650_, new_n30651_, new_n30652_, new_n30653_, new_n30654_,
    new_n30655_, new_n30656_, new_n30657_, new_n30658_, new_n30659_,
    new_n30660_, new_n30661_, new_n30662_, new_n30663_, new_n30664_,
    new_n30665_, new_n30666_, new_n30667_, new_n30668_, new_n30669_,
    new_n30670_, new_n30671_, new_n30672_, new_n30673_, new_n30674_,
    new_n30675_, new_n30676_, new_n30677_, new_n30678_, new_n30679_,
    new_n30680_, new_n30681_, new_n30682_, new_n30683_, new_n30684_,
    new_n30685_, new_n30686_, new_n30687_, new_n30688_, new_n30689_,
    new_n30690_, new_n30691_, new_n30692_, new_n30693_, new_n30694_,
    new_n30695_, new_n30696_, new_n30697_, new_n30698_, new_n30699_,
    new_n30700_, new_n30701_, new_n30702_, new_n30703_, new_n30704_,
    new_n30705_, new_n30706_, new_n30707_, new_n30708_, new_n30709_,
    new_n30710_, new_n30711_, new_n30712_, new_n30713_, new_n30714_,
    new_n30715_, new_n30716_, new_n30717_, new_n30718_, new_n30719_,
    new_n30720_, new_n30721_, new_n30722_, new_n30723_, new_n30724_,
    new_n30725_, new_n30726_, new_n30727_, new_n30728_, new_n30729_,
    new_n30730_, new_n30731_, new_n30732_, new_n30733_, new_n30734_,
    new_n30735_, new_n30736_, new_n30737_, new_n30738_, new_n30739_,
    new_n30740_, new_n30741_, new_n30742_, new_n30743_, new_n30744_,
    new_n30745_, new_n30746_, new_n30747_, new_n30748_, new_n30749_,
    new_n30750_, new_n30751_, new_n30752_, new_n30753_, new_n30754_,
    new_n30755_, new_n30756_, new_n30757_, new_n30758_, new_n30759_,
    new_n30760_, new_n30761_, new_n30762_, new_n30763_, new_n30764_,
    new_n30765_, new_n30766_, new_n30767_, new_n30768_, new_n30769_,
    new_n30770_, new_n30771_, new_n30772_, new_n30773_, new_n30774_,
    new_n30775_, new_n30776_, new_n30777_, new_n30778_, new_n30779_,
    new_n30780_, new_n30781_, new_n30782_, new_n30783_, new_n30784_,
    new_n30785_, new_n30786_, new_n30787_, new_n30788_, new_n30789_,
    new_n30790_, new_n30791_, new_n30792_, new_n30793_, new_n30794_,
    new_n30795_, new_n30796_, new_n30797_, new_n30798_, new_n30799_,
    new_n30800_, new_n30801_, new_n30802_, new_n30803_, new_n30804_,
    new_n30805_, new_n30806_, new_n30807_, new_n30808_, new_n30809_,
    new_n30810_, new_n30811_, new_n30812_, new_n30813_, new_n30814_,
    new_n30815_, new_n30816_, new_n30817_, new_n30818_, new_n30819_,
    new_n30820_, new_n30821_, new_n30822_, new_n30824_, new_n30825_,
    new_n30826_, new_n30827_, new_n30828_, new_n30829_, new_n30830_,
    new_n30831_, new_n30832_, new_n30833_, new_n30834_, new_n30835_,
    new_n30836_, new_n30837_, new_n30838_, new_n30839_, new_n30840_,
    new_n30841_, new_n30842_, new_n30843_, new_n30844_, new_n30845_,
    new_n30846_, new_n30847_, new_n30848_, new_n30849_, new_n30850_,
    new_n30851_, new_n30852_, new_n30853_, new_n30854_, new_n30855_,
    new_n30856_, new_n30857_, new_n30858_, new_n30859_, new_n30860_,
    new_n30861_, new_n30862_, new_n30863_, new_n30864_, new_n30865_,
    new_n30866_, new_n30867_, new_n30868_, new_n30869_, new_n30870_,
    new_n30871_, new_n30872_, new_n30873_, new_n30874_, new_n30875_,
    new_n30876_, new_n30877_, new_n30878_, new_n30879_, new_n30880_,
    new_n30881_, new_n30882_, new_n30883_, new_n30884_, new_n30885_,
    new_n30886_, new_n30887_, new_n30888_, new_n30889_, new_n30890_,
    new_n30891_, new_n30892_, new_n30893_, new_n30894_, new_n30895_,
    new_n30896_, new_n30897_, new_n30898_, new_n30899_, new_n30900_,
    new_n30901_, new_n30902_, new_n30903_, new_n30904_, new_n30905_,
    new_n30906_, new_n30907_, new_n30908_, new_n30909_, new_n30910_,
    new_n30911_, new_n30912_, new_n30913_, new_n30914_, new_n30915_,
    new_n30916_, new_n30917_, new_n30918_, new_n30919_, new_n30920_,
    new_n30921_, new_n30922_, new_n30923_, new_n30924_, new_n30925_,
    new_n30926_, new_n30927_, new_n30928_, new_n30929_, new_n30930_,
    new_n30931_, new_n30932_, new_n30933_, new_n30934_, new_n30935_,
    new_n30936_, new_n30937_, new_n30938_, new_n30939_, new_n30940_,
    new_n30941_, new_n30942_, new_n30943_, new_n30944_, new_n30945_,
    new_n30946_, new_n30947_, new_n30948_, new_n30949_, new_n30950_,
    new_n30951_, new_n30952_, new_n30953_, new_n30954_, new_n30955_,
    new_n30956_, new_n30957_, new_n30958_, new_n30959_, new_n30960_,
    new_n30961_, new_n30962_, new_n30963_, new_n30964_, new_n30965_,
    new_n30966_, new_n30967_, new_n30968_, new_n30969_, new_n30970_,
    new_n30971_, new_n30972_, new_n30973_, new_n30974_, new_n30975_,
    new_n30976_, new_n30977_, new_n30978_, new_n30979_, new_n30980_,
    new_n30981_, new_n30982_, new_n30983_, new_n30984_, new_n30985_,
    new_n30986_, new_n30987_, new_n30988_, new_n30989_, new_n30990_,
    new_n30991_, new_n30992_, new_n30993_, new_n30994_, new_n30995_,
    new_n30996_, new_n30997_, new_n30998_, new_n30999_, new_n31000_,
    new_n31001_, new_n31002_, new_n31003_, new_n31004_, new_n31005_,
    new_n31006_, new_n31007_, new_n31008_, new_n31009_, new_n31010_,
    new_n31011_, new_n31012_, new_n31013_, new_n31014_, new_n31015_,
    new_n31016_, new_n31017_, new_n31018_, new_n31019_, new_n31020_,
    new_n31021_, new_n31022_, new_n31023_, new_n31024_, new_n31025_,
    new_n31026_, new_n31027_, new_n31028_, new_n31029_, new_n31030_,
    new_n31031_, new_n31032_, new_n31033_, new_n31034_, new_n31035_,
    new_n31036_, new_n31037_, new_n31038_, new_n31039_, new_n31040_,
    new_n31041_, new_n31042_, new_n31043_, new_n31044_, new_n31045_,
    new_n31046_, new_n31047_, new_n31048_, new_n31049_, new_n31050_,
    new_n31051_, new_n31052_, new_n31053_, new_n31054_, new_n31055_,
    new_n31056_, new_n31057_, new_n31058_, new_n31059_, new_n31060_,
    new_n31061_, new_n31062_, new_n31063_, new_n31064_, new_n31065_,
    new_n31066_, new_n31067_, new_n31068_, new_n31069_, new_n31070_,
    new_n31071_, new_n31072_, new_n31073_, new_n31074_, new_n31075_,
    new_n31076_, new_n31077_, new_n31078_, new_n31079_, new_n31080_,
    new_n31081_, new_n31082_, new_n31083_, new_n31084_, new_n31085_,
    new_n31086_, new_n31087_, new_n31088_, new_n31089_, new_n31090_,
    new_n31091_, new_n31092_, new_n31093_, new_n31094_, new_n31095_,
    new_n31096_, new_n31097_, new_n31098_, new_n31099_, new_n31100_,
    new_n31101_, new_n31102_, new_n31103_, new_n31104_, new_n31105_,
    new_n31106_, new_n31107_, new_n31108_, new_n31109_, new_n31110_,
    new_n31111_, new_n31112_, new_n31113_, new_n31114_, new_n31115_,
    new_n31116_, new_n31117_, new_n31118_, new_n31119_, new_n31120_,
    new_n31121_, new_n31122_, new_n31123_, new_n31124_, new_n31125_,
    new_n31126_, new_n31127_, new_n31128_, new_n31129_, new_n31130_,
    new_n31131_, new_n31132_, new_n31133_, new_n31134_, new_n31135_,
    new_n31136_, new_n31137_, new_n31138_, new_n31139_, new_n31140_,
    new_n31141_, new_n31142_, new_n31143_, new_n31144_, new_n31145_,
    new_n31146_, new_n31147_, new_n31148_, new_n31149_, new_n31150_,
    new_n31151_, new_n31152_, new_n31153_, new_n31154_, new_n31155_,
    new_n31156_, new_n31157_, new_n31158_, new_n31159_, new_n31160_,
    new_n31161_, new_n31162_, new_n31163_, new_n31164_, new_n31165_,
    new_n31166_, new_n31167_, new_n31168_, new_n31169_, new_n31170_,
    new_n31171_, new_n31172_, new_n31173_, new_n31174_, new_n31175_,
    new_n31176_, new_n31177_, new_n31178_, new_n31179_, new_n31180_,
    new_n31181_, new_n31182_, new_n31183_, new_n31184_, new_n31185_,
    new_n31186_, new_n31187_, new_n31188_, new_n31189_, new_n31190_,
    new_n31191_, new_n31192_, new_n31193_, new_n31194_, new_n31195_,
    new_n31196_, new_n31197_, new_n31198_, new_n31199_, new_n31200_,
    new_n31201_, new_n31202_, new_n31203_, new_n31204_, new_n31205_,
    new_n31206_, new_n31207_, new_n31208_, new_n31209_, new_n31210_,
    new_n31211_, new_n31212_, new_n31213_, new_n31214_, new_n31215_,
    new_n31216_, new_n31217_, new_n31218_, new_n31219_, new_n31220_,
    new_n31221_, new_n31222_, new_n31223_, new_n31224_, new_n31225_,
    new_n31226_, new_n31227_, new_n31228_, new_n31229_, new_n31230_,
    new_n31231_, new_n31232_, new_n31233_, new_n31234_, new_n31235_,
    new_n31236_, new_n31237_, new_n31238_, new_n31239_, new_n31240_,
    new_n31241_, new_n31242_, new_n31243_, new_n31244_, new_n31245_,
    new_n31246_, new_n31247_, new_n31248_, new_n31249_, new_n31250_,
    new_n31251_, new_n31252_, new_n31253_, new_n31254_, new_n31255_,
    new_n31256_, new_n31257_, new_n31258_, new_n31259_, new_n31260_,
    new_n31261_, new_n31262_, new_n31263_, new_n31264_, new_n31265_,
    new_n31266_, new_n31267_, new_n31268_, new_n31269_, new_n31270_,
    new_n31271_, new_n31272_, new_n31273_, new_n31274_, new_n31275_,
    new_n31276_, new_n31277_, new_n31278_, new_n31279_, new_n31280_,
    new_n31281_, new_n31282_, new_n31283_, new_n31284_, new_n31285_,
    new_n31286_, new_n31287_, new_n31288_, new_n31289_, new_n31290_,
    new_n31291_, new_n31292_, new_n31293_, new_n31294_, new_n31295_,
    new_n31296_, new_n31297_, new_n31298_, new_n31299_, new_n31301_,
    new_n31302_, new_n31303_, new_n31304_, new_n31305_, new_n31306_,
    new_n31307_, new_n31308_, new_n31309_, new_n31310_, new_n31311_,
    new_n31312_, new_n31313_, new_n31314_, new_n31315_, new_n31316_,
    new_n31317_, new_n31318_, new_n31319_, new_n31320_, new_n31321_,
    new_n31322_, new_n31323_, new_n31324_, new_n31325_, new_n31326_,
    new_n31327_, new_n31328_, new_n31329_, new_n31330_, new_n31331_,
    new_n31332_, new_n31333_, new_n31334_, new_n31335_, new_n31336_,
    new_n31337_, new_n31338_, new_n31339_, new_n31340_, new_n31341_,
    new_n31342_, new_n31343_, new_n31344_, new_n31345_, new_n31346_,
    new_n31347_, new_n31348_, new_n31349_, new_n31350_, new_n31351_,
    new_n31352_, new_n31353_, new_n31354_, new_n31355_, new_n31356_,
    new_n31357_, new_n31358_, new_n31359_, new_n31360_, new_n31361_,
    new_n31362_, new_n31363_, new_n31364_, new_n31365_, new_n31366_,
    new_n31367_, new_n31368_, new_n31369_, new_n31370_, new_n31371_,
    new_n31372_, new_n31373_, new_n31374_, new_n31375_, new_n31376_,
    new_n31377_, new_n31378_, new_n31379_, new_n31380_, new_n31381_,
    new_n31382_, new_n31383_, new_n31384_, new_n31385_, new_n31386_,
    new_n31387_, new_n31388_, new_n31389_, new_n31390_, new_n31391_,
    new_n31392_, new_n31393_, new_n31394_, new_n31395_, new_n31396_,
    new_n31397_, new_n31398_, new_n31399_, new_n31400_, new_n31401_,
    new_n31402_, new_n31403_, new_n31404_, new_n31405_, new_n31406_,
    new_n31407_, new_n31408_, new_n31409_, new_n31410_, new_n31411_,
    new_n31412_, new_n31413_, new_n31414_, new_n31415_, new_n31416_,
    new_n31417_, new_n31418_, new_n31419_, new_n31420_, new_n31421_,
    new_n31422_, new_n31423_, new_n31424_, new_n31425_, new_n31426_,
    new_n31427_, new_n31428_, new_n31429_, new_n31430_, new_n31431_,
    new_n31432_, new_n31433_, new_n31434_, new_n31435_, new_n31436_,
    new_n31437_, new_n31438_, new_n31439_, new_n31440_, new_n31441_,
    new_n31442_, new_n31443_, new_n31444_, new_n31445_, new_n31446_,
    new_n31447_, new_n31448_, new_n31449_, new_n31450_, new_n31451_,
    new_n31452_, new_n31453_, new_n31454_, new_n31455_, new_n31456_,
    new_n31457_, new_n31458_, new_n31459_, new_n31460_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31472_, new_n31473_, new_n31474_, new_n31475_, new_n31476_,
    new_n31477_, new_n31478_, new_n31479_, new_n31480_, new_n31481_,
    new_n31482_, new_n31483_, new_n31484_, new_n31485_, new_n31486_,
    new_n31487_, new_n31488_, new_n31489_, new_n31490_, new_n31491_,
    new_n31492_, new_n31493_, new_n31494_, new_n31495_, new_n31496_,
    new_n31497_, new_n31498_, new_n31499_, new_n31500_, new_n31501_,
    new_n31502_, new_n31503_, new_n31504_, new_n31505_, new_n31506_,
    new_n31507_, new_n31508_, new_n31509_, new_n31510_, new_n31511_,
    new_n31512_, new_n31513_, new_n31514_, new_n31515_, new_n31516_,
    new_n31517_, new_n31518_, new_n31519_, new_n31520_, new_n31521_,
    new_n31522_, new_n31523_, new_n31524_, new_n31525_, new_n31526_,
    new_n31527_, new_n31528_, new_n31529_, new_n31530_, new_n31531_,
    new_n31532_, new_n31533_, new_n31534_, new_n31535_, new_n31536_,
    new_n31537_, new_n31538_, new_n31539_, new_n31540_, new_n31541_,
    new_n31542_, new_n31543_, new_n31544_, new_n31545_, new_n31546_,
    new_n31547_, new_n31548_, new_n31549_, new_n31550_, new_n31551_,
    new_n31552_, new_n31553_, new_n31554_, new_n31555_, new_n31556_,
    new_n31557_, new_n31558_, new_n31559_, new_n31560_, new_n31561_,
    new_n31562_, new_n31563_, new_n31564_, new_n31565_, new_n31566_,
    new_n31567_, new_n31568_, new_n31569_, new_n31570_, new_n31571_,
    new_n31572_, new_n31573_, new_n31574_, new_n31575_, new_n31576_,
    new_n31577_, new_n31578_, new_n31579_, new_n31580_, new_n31581_,
    new_n31582_, new_n31583_, new_n31584_, new_n31585_, new_n31586_,
    new_n31587_, new_n31588_, new_n31589_, new_n31590_, new_n31591_,
    new_n31592_, new_n31593_, new_n31594_, new_n31595_, new_n31596_,
    new_n31597_, new_n31598_, new_n31599_, new_n31600_, new_n31601_,
    new_n31602_, new_n31603_, new_n31604_, new_n31605_, new_n31606_,
    new_n31607_, new_n31608_, new_n31609_, new_n31610_, new_n31611_,
    new_n31612_, new_n31613_, new_n31614_, new_n31615_, new_n31616_,
    new_n31617_, new_n31618_, new_n31619_, new_n31620_, new_n31621_,
    new_n31622_, new_n31623_, new_n31624_, new_n31625_, new_n31626_,
    new_n31627_, new_n31628_, new_n31629_, new_n31630_, new_n31631_,
    new_n31632_, new_n31633_, new_n31634_, new_n31635_, new_n31636_,
    new_n31637_, new_n31638_, new_n31639_, new_n31640_, new_n31641_,
    new_n31642_, new_n31643_, new_n31644_, new_n31645_, new_n31646_,
    new_n31647_, new_n31648_, new_n31649_, new_n31650_, new_n31651_,
    new_n31652_, new_n31653_, new_n31654_, new_n31655_, new_n31656_,
    new_n31657_, new_n31658_, new_n31659_, new_n31660_, new_n31661_,
    new_n31662_, new_n31663_, new_n31664_, new_n31665_, new_n31666_,
    new_n31667_, new_n31668_, new_n31669_, new_n31670_, new_n31671_,
    new_n31672_, new_n31673_, new_n31674_, new_n31675_, new_n31676_,
    new_n31677_, new_n31678_, new_n31679_, new_n31680_, new_n31681_,
    new_n31682_, new_n31683_, new_n31684_, new_n31685_, new_n31686_,
    new_n31687_, new_n31688_, new_n31689_, new_n31690_, new_n31691_,
    new_n31692_, new_n31693_, new_n31694_, new_n31695_, new_n31696_,
    new_n31697_, new_n31698_, new_n31699_, new_n31700_, new_n31701_,
    new_n31702_, new_n31703_, new_n31704_, new_n31705_, new_n31706_,
    new_n31707_, new_n31708_, new_n31709_, new_n31710_, new_n31711_,
    new_n31712_, new_n31713_, new_n31714_, new_n31715_, new_n31716_,
    new_n31717_, new_n31718_, new_n31719_, new_n31720_, new_n31721_,
    new_n31722_, new_n31723_, new_n31724_, new_n31725_, new_n31726_,
    new_n31727_, new_n31728_, new_n31729_, new_n31730_, new_n31731_,
    new_n31732_, new_n31733_, new_n31734_, new_n31735_, new_n31736_,
    new_n31737_, new_n31738_, new_n31739_, new_n31740_, new_n31741_,
    new_n31742_, new_n31743_, new_n31744_, new_n31745_, new_n31746_,
    new_n31747_, new_n31748_, new_n31749_, new_n31750_, new_n31751_,
    new_n31752_, new_n31753_, new_n31754_, new_n31755_, new_n31756_,
    new_n31757_, new_n31758_, new_n31759_, new_n31760_, new_n31761_,
    new_n31762_, new_n31763_, new_n31764_, new_n31765_, new_n31766_,
    new_n31767_, new_n31768_, new_n31769_, new_n31770_, new_n31771_,
    new_n31772_, new_n31773_, new_n31774_, new_n31775_, new_n31776_,
    new_n31778_, new_n31779_, new_n31780_, new_n31781_, new_n31782_,
    new_n31783_, new_n31784_, new_n31785_, new_n31786_, new_n31787_,
    new_n31788_, new_n31789_, new_n31790_, new_n31791_, new_n31792_,
    new_n31793_, new_n31794_, new_n31795_, new_n31796_, new_n31797_,
    new_n31798_, new_n31799_, new_n31800_, new_n31801_, new_n31802_,
    new_n31803_, new_n31804_, new_n31805_, new_n31806_, new_n31807_,
    new_n31808_, new_n31809_, new_n31810_, new_n31811_, new_n31812_,
    new_n31813_, new_n31814_, new_n31815_, new_n31816_, new_n31817_,
    new_n31818_, new_n31819_, new_n31820_, new_n31821_, new_n31822_,
    new_n31823_, new_n31824_, new_n31825_, new_n31826_, new_n31827_,
    new_n31828_, new_n31829_, new_n31830_, new_n31831_, new_n31832_,
    new_n31833_, new_n31834_, new_n31835_, new_n31836_, new_n31837_,
    new_n31838_, new_n31839_, new_n31840_, new_n31841_, new_n31842_,
    new_n31843_, new_n31844_, new_n31845_, new_n31846_, new_n31847_,
    new_n31848_, new_n31849_, new_n31850_, new_n31851_, new_n31852_,
    new_n31853_, new_n31854_, new_n31855_, new_n31856_, new_n31857_,
    new_n31858_, new_n31859_, new_n31860_, new_n31861_, new_n31862_,
    new_n31863_, new_n31864_, new_n31865_, new_n31866_, new_n31867_,
    new_n31868_, new_n31869_, new_n31870_, new_n31871_, new_n31872_,
    new_n31873_, new_n31874_, new_n31875_, new_n31876_, new_n31877_,
    new_n31878_, new_n31879_, new_n31880_, new_n31881_, new_n31882_,
    new_n31883_, new_n31884_, new_n31885_, new_n31886_, new_n31887_,
    new_n31888_, new_n31889_, new_n31890_, new_n31891_, new_n31892_,
    new_n31893_, new_n31894_, new_n31895_, new_n31896_, new_n31897_,
    new_n31898_, new_n31899_, new_n31900_, new_n31901_, new_n31902_,
    new_n31903_, new_n31904_, new_n31905_, new_n31906_, new_n31907_,
    new_n31908_, new_n31909_, new_n31910_, new_n31911_, new_n31912_,
    new_n31913_, new_n31914_, new_n31915_, new_n31916_, new_n31917_,
    new_n31918_, new_n31919_, new_n31920_, new_n31921_, new_n31922_,
    new_n31923_, new_n31924_, new_n31925_, new_n31926_, new_n31927_,
    new_n31928_, new_n31929_, new_n31930_, new_n31931_, new_n31932_,
    new_n31933_, new_n31934_, new_n31935_, new_n31936_, new_n31937_,
    new_n31938_, new_n31939_, new_n31940_, new_n31941_, new_n31942_,
    new_n31943_, new_n31944_, new_n31945_, new_n31946_, new_n31947_,
    new_n31948_, new_n31949_, new_n31950_, new_n31951_, new_n31952_,
    new_n31953_, new_n31954_, new_n31955_, new_n31956_, new_n31957_,
    new_n31958_, new_n31959_, new_n31960_, new_n31961_, new_n31962_,
    new_n31963_, new_n31964_, new_n31965_, new_n31966_, new_n31967_,
    new_n31968_, new_n31969_, new_n31970_, new_n31971_, new_n31972_,
    new_n31973_, new_n31974_, new_n31975_, new_n31976_, new_n31977_,
    new_n31978_, new_n31979_, new_n31980_, new_n31981_, new_n31982_,
    new_n31983_, new_n31984_, new_n31985_, new_n31986_, new_n31987_,
    new_n31988_, new_n31989_, new_n31990_, new_n31991_, new_n31992_,
    new_n31993_, new_n31994_, new_n31995_, new_n31996_, new_n31997_,
    new_n31998_, new_n31999_, new_n32000_, new_n32001_, new_n32002_,
    new_n32003_, new_n32004_, new_n32005_, new_n32006_, new_n32007_,
    new_n32008_, new_n32009_, new_n32010_, new_n32011_, new_n32012_,
    new_n32013_, new_n32014_, new_n32015_, new_n32016_, new_n32017_,
    new_n32018_, new_n32019_, new_n32020_, new_n32021_, new_n32022_,
    new_n32023_, new_n32024_, new_n32025_, new_n32026_, new_n32027_,
    new_n32028_, new_n32029_, new_n32030_, new_n32031_, new_n32032_,
    new_n32033_, new_n32034_, new_n32035_, new_n32036_, new_n32037_,
    new_n32038_, new_n32039_, new_n32040_, new_n32041_, new_n32042_,
    new_n32043_, new_n32044_, new_n32045_, new_n32046_, new_n32047_,
    new_n32048_, new_n32049_, new_n32050_, new_n32051_, new_n32052_,
    new_n32053_, new_n32054_, new_n32055_, new_n32056_, new_n32057_,
    new_n32058_, new_n32059_, new_n32060_, new_n32061_, new_n32062_,
    new_n32063_, new_n32064_, new_n32065_, new_n32066_, new_n32067_,
    new_n32068_, new_n32069_, new_n32070_, new_n32071_, new_n32072_,
    new_n32073_, new_n32074_, new_n32075_, new_n32076_, new_n32077_,
    new_n32078_, new_n32079_, new_n32080_, new_n32081_, new_n32082_,
    new_n32083_, new_n32084_, new_n32085_, new_n32086_, new_n32087_,
    new_n32088_, new_n32089_, new_n32090_, new_n32091_, new_n32092_,
    new_n32093_, new_n32094_, new_n32095_, new_n32096_, new_n32097_,
    new_n32098_, new_n32099_, new_n32100_, new_n32101_, new_n32102_,
    new_n32103_, new_n32104_, new_n32105_, new_n32106_, new_n32107_,
    new_n32108_, new_n32109_, new_n32110_, new_n32111_, new_n32112_,
    new_n32113_, new_n32114_, new_n32115_, new_n32116_, new_n32117_,
    new_n32118_, new_n32119_, new_n32120_, new_n32121_, new_n32122_,
    new_n32123_, new_n32124_, new_n32125_, new_n32126_, new_n32127_,
    new_n32128_, new_n32129_, new_n32130_, new_n32131_, new_n32132_,
    new_n32133_, new_n32134_, new_n32135_, new_n32136_, new_n32137_,
    new_n32138_, new_n32139_, new_n32140_, new_n32141_, new_n32142_,
    new_n32143_, new_n32144_, new_n32145_, new_n32146_, new_n32147_,
    new_n32148_, new_n32149_, new_n32150_, new_n32151_, new_n32152_,
    new_n32153_, new_n32154_, new_n32155_, new_n32156_, new_n32157_,
    new_n32158_, new_n32159_, new_n32160_, new_n32161_, new_n32162_,
    new_n32163_, new_n32164_, new_n32165_, new_n32166_, new_n32167_,
    new_n32168_, new_n32169_, new_n32170_, new_n32171_, new_n32172_,
    new_n32173_, new_n32174_, new_n32175_, new_n32176_, new_n32177_,
    new_n32178_, new_n32179_, new_n32180_, new_n32181_, new_n32182_,
    new_n32183_, new_n32184_, new_n32185_, new_n32186_, new_n32187_,
    new_n32188_, new_n32189_, new_n32190_, new_n32191_, new_n32192_,
    new_n32193_, new_n32194_, new_n32195_, new_n32196_, new_n32197_,
    new_n32198_, new_n32199_, new_n32200_, new_n32201_, new_n32202_,
    new_n32203_, new_n32204_, new_n32205_, new_n32206_, new_n32207_,
    new_n32208_, new_n32209_, new_n32210_, new_n32211_, new_n32212_,
    new_n32213_, new_n32214_, new_n32215_, new_n32216_, new_n32217_,
    new_n32218_, new_n32219_, new_n32220_, new_n32221_, new_n32222_,
    new_n32223_, new_n32224_, new_n32225_, new_n32226_, new_n32227_,
    new_n32228_, new_n32229_, new_n32230_, new_n32231_, new_n32232_,
    new_n32233_, new_n32234_, new_n32235_, new_n32236_, new_n32237_,
    new_n32238_, new_n32239_, new_n32240_, new_n32241_, new_n32242_,
    new_n32243_, new_n32244_, new_n32245_, new_n32246_, new_n32247_,
    new_n32248_, new_n32249_, new_n32250_, new_n32251_, new_n32252_,
    new_n32253_, new_n32255_, new_n32256_, new_n32257_, new_n32258_,
    new_n32259_, new_n32260_, new_n32261_, new_n32262_, new_n32263_,
    new_n32264_, new_n32265_, new_n32266_, new_n32267_, new_n32268_,
    new_n32269_, new_n32270_, new_n32271_, new_n32272_, new_n32273_,
    new_n32274_, new_n32275_, new_n32276_, new_n32277_, new_n32278_,
    new_n32279_, new_n32280_, new_n32281_, new_n32282_, new_n32283_,
    new_n32284_, new_n32285_, new_n32286_, new_n32287_, new_n32288_,
    new_n32289_, new_n32290_, new_n32291_, new_n32292_, new_n32293_,
    new_n32294_, new_n32295_, new_n32296_, new_n32297_, new_n32298_,
    new_n32299_, new_n32300_, new_n32301_, new_n32302_, new_n32303_,
    new_n32304_, new_n32305_, new_n32306_, new_n32307_, new_n32308_,
    new_n32309_, new_n32310_, new_n32311_, new_n32312_, new_n32313_,
    new_n32314_, new_n32315_, new_n32316_, new_n32317_, new_n32318_,
    new_n32319_, new_n32320_, new_n32321_, new_n32322_, new_n32323_,
    new_n32324_, new_n32325_, new_n32326_, new_n32327_, new_n32328_,
    new_n32329_, new_n32330_, new_n32331_, new_n32332_, new_n32333_,
    new_n32334_, new_n32335_, new_n32336_, new_n32337_, new_n32338_,
    new_n32339_, new_n32340_, new_n32341_, new_n32342_, new_n32343_,
    new_n32344_, new_n32345_, new_n32346_, new_n32347_, new_n32348_,
    new_n32349_, new_n32350_, new_n32351_, new_n32352_, new_n32353_,
    new_n32354_, new_n32355_, new_n32356_, new_n32357_, new_n32358_,
    new_n32359_, new_n32360_, new_n32361_, new_n32362_, new_n32363_,
    new_n32364_, new_n32365_, new_n32366_, new_n32367_, new_n32368_,
    new_n32369_, new_n32370_, new_n32371_, new_n32372_, new_n32373_,
    new_n32374_, new_n32375_, new_n32376_, new_n32377_, new_n32378_,
    new_n32379_, new_n32380_, new_n32381_, new_n32382_, new_n32383_,
    new_n32384_, new_n32385_, new_n32386_, new_n32387_, new_n32388_,
    new_n32389_, new_n32390_, new_n32391_, new_n32392_, new_n32393_,
    new_n32394_, new_n32395_, new_n32396_, new_n32397_, new_n32398_,
    new_n32399_, new_n32400_, new_n32401_, new_n32402_, new_n32403_,
    new_n32404_, new_n32405_, new_n32406_, new_n32407_, new_n32408_,
    new_n32409_, new_n32410_, new_n32411_, new_n32412_, new_n32413_,
    new_n32414_, new_n32415_, new_n32416_, new_n32417_, new_n32418_,
    new_n32419_, new_n32420_, new_n32421_, new_n32422_, new_n32423_,
    new_n32424_, new_n32425_, new_n32426_, new_n32427_, new_n32428_,
    new_n32429_, new_n32430_, new_n32431_, new_n32432_, new_n32433_,
    new_n32434_, new_n32435_, new_n32436_, new_n32437_, new_n32438_,
    new_n32439_, new_n32440_, new_n32441_, new_n32442_, new_n32443_,
    new_n32444_, new_n32445_, new_n32446_, new_n32447_, new_n32448_,
    new_n32449_, new_n32450_, new_n32451_, new_n32452_, new_n32453_,
    new_n32454_, new_n32455_, new_n32456_, new_n32457_, new_n32458_,
    new_n32459_, new_n32460_, new_n32461_, new_n32462_, new_n32463_,
    new_n32464_, new_n32465_, new_n32466_, new_n32467_, new_n32468_,
    new_n32469_, new_n32470_, new_n32471_, new_n32472_, new_n32473_,
    new_n32474_, new_n32475_, new_n32476_, new_n32477_, new_n32478_,
    new_n32479_, new_n32480_, new_n32481_, new_n32482_, new_n32483_,
    new_n32484_, new_n32485_, new_n32486_, new_n32487_, new_n32488_,
    new_n32489_, new_n32490_, new_n32491_, new_n32492_, new_n32493_,
    new_n32494_, new_n32495_, new_n32496_, new_n32497_, new_n32498_,
    new_n32499_, new_n32500_, new_n32501_, new_n32502_, new_n32503_,
    new_n32504_, new_n32505_, new_n32506_, new_n32507_, new_n32508_,
    new_n32509_, new_n32510_, new_n32511_, new_n32512_, new_n32513_,
    new_n32514_, new_n32515_, new_n32516_, new_n32517_, new_n32518_,
    new_n32519_, new_n32520_, new_n32521_, new_n32522_, new_n32523_,
    new_n32524_, new_n32525_, new_n32526_, new_n32527_, new_n32528_,
    new_n32529_, new_n32530_, new_n32531_, new_n32532_, new_n32533_,
    new_n32534_, new_n32535_, new_n32536_, new_n32537_, new_n32538_,
    new_n32539_, new_n32540_, new_n32541_, new_n32542_, new_n32543_,
    new_n32544_, new_n32545_, new_n32546_, new_n32547_, new_n32548_,
    new_n32549_, new_n32550_, new_n32551_, new_n32552_, new_n32553_,
    new_n32554_, new_n32555_, new_n32556_, new_n32557_, new_n32558_,
    new_n32559_, new_n32560_, new_n32561_, new_n32562_, new_n32563_,
    new_n32564_, new_n32565_, new_n32566_, new_n32567_, new_n32568_,
    new_n32569_, new_n32570_, new_n32571_, new_n32572_, new_n32573_,
    new_n32574_, new_n32575_, new_n32576_, new_n32577_, new_n32578_,
    new_n32579_, new_n32580_, new_n32581_, new_n32582_, new_n32583_,
    new_n32584_, new_n32585_, new_n32586_, new_n32587_, new_n32588_,
    new_n32589_, new_n32590_, new_n32591_, new_n32592_, new_n32593_,
    new_n32594_, new_n32595_, new_n32596_, new_n32597_, new_n32598_,
    new_n32599_, new_n32600_, new_n32601_, new_n32602_, new_n32603_,
    new_n32604_, new_n32605_, new_n32606_, new_n32607_, new_n32608_,
    new_n32609_, new_n32610_, new_n32611_, new_n32612_, new_n32613_,
    new_n32614_, new_n32615_, new_n32616_, new_n32617_, new_n32618_,
    new_n32619_, new_n32620_, new_n32621_, new_n32622_, new_n32623_,
    new_n32624_, new_n32625_, new_n32626_, new_n32627_, new_n32628_,
    new_n32629_, new_n32630_, new_n32631_, new_n32632_, new_n32633_,
    new_n32634_, new_n32635_, new_n32636_, new_n32637_, new_n32638_,
    new_n32639_, new_n32640_, new_n32641_, new_n32642_, new_n32643_,
    new_n32644_, new_n32645_, new_n32646_, new_n32647_, new_n32648_,
    new_n32649_, new_n32650_, new_n32651_, new_n32652_, new_n32653_,
    new_n32654_, new_n32655_, new_n32656_, new_n32657_, new_n32658_,
    new_n32659_, new_n32660_, new_n32661_, new_n32662_, new_n32663_,
    new_n32664_, new_n32665_, new_n32666_, new_n32667_, new_n32668_,
    new_n32669_, new_n32670_, new_n32671_, new_n32672_, new_n32673_,
    new_n32674_, new_n32675_, new_n32676_, new_n32677_, new_n32678_,
    new_n32679_, new_n32680_, new_n32681_, new_n32682_, new_n32683_,
    new_n32684_, new_n32685_, new_n32686_, new_n32687_, new_n32688_,
    new_n32689_, new_n32690_, new_n32691_, new_n32692_, new_n32693_,
    new_n32694_, new_n32695_, new_n32696_, new_n32697_, new_n32698_,
    new_n32699_, new_n32700_, new_n32701_, new_n32702_, new_n32703_,
    new_n32704_, new_n32705_, new_n32706_, new_n32707_, new_n32708_,
    new_n32709_, new_n32710_, new_n32711_, new_n32712_, new_n32713_,
    new_n32714_, new_n32715_, new_n32716_, new_n32717_, new_n32718_,
    new_n32719_, new_n32720_, new_n32721_, new_n32722_, new_n32723_,
    new_n32724_, new_n32725_, new_n32727_, new_n32728_, new_n32729_,
    new_n32730_, new_n32731_, new_n32732_, new_n32733_, new_n32734_,
    new_n32735_, new_n32736_, new_n32737_, new_n32738_, new_n32739_,
    new_n32740_, new_n32741_, new_n32742_, new_n32743_, new_n32744_,
    new_n32745_, new_n32746_, new_n32747_, new_n32748_, new_n32749_,
    new_n32750_, new_n32751_, new_n32752_, new_n32753_, new_n32754_,
    new_n32755_, new_n32756_, new_n32757_, new_n32758_, new_n32759_,
    new_n32760_, new_n32761_, new_n32762_, new_n32763_, new_n32764_,
    new_n32765_, new_n32766_, new_n32767_, new_n32768_, new_n32769_,
    new_n32770_, new_n32771_, new_n32772_, new_n32773_, new_n32774_,
    new_n32775_, new_n32776_, new_n32777_, new_n32778_, new_n32779_,
    new_n32780_, new_n32781_, new_n32782_, new_n32783_, new_n32784_,
    new_n32785_, new_n32786_, new_n32787_, new_n32788_, new_n32789_,
    new_n32790_, new_n32791_, new_n32792_, new_n32793_, new_n32794_,
    new_n32795_, new_n32796_, new_n32797_, new_n32798_, new_n32799_,
    new_n32800_, new_n32801_, new_n32802_, new_n32803_, new_n32804_,
    new_n32805_, new_n32806_, new_n32807_, new_n32808_, new_n32809_,
    new_n32810_, new_n32811_, new_n32812_, new_n32813_, new_n32814_,
    new_n32815_, new_n32816_, new_n32817_, new_n32818_, new_n32819_,
    new_n32820_, new_n32821_, new_n32822_, new_n32823_, new_n32824_,
    new_n32825_, new_n32826_, new_n32827_, new_n32828_, new_n32829_,
    new_n32830_, new_n32831_, new_n32832_, new_n32833_, new_n32834_,
    new_n32835_, new_n32836_, new_n32837_, new_n32838_, new_n32839_,
    new_n32840_, new_n32841_, new_n32842_, new_n32843_, new_n32844_,
    new_n32845_, new_n32846_, new_n32847_, new_n32848_, new_n32849_,
    new_n32850_, new_n32851_, new_n32852_, new_n32853_, new_n32854_,
    new_n32855_, new_n32856_, new_n32857_, new_n32858_, new_n32859_,
    new_n32860_, new_n32861_, new_n32862_, new_n32863_, new_n32864_,
    new_n32865_, new_n32866_, new_n32867_, new_n32868_, new_n32869_,
    new_n32870_, new_n32871_, new_n32872_, new_n32873_, new_n32874_,
    new_n32875_, new_n32876_, new_n32877_, new_n32878_, new_n32879_,
    new_n32880_, new_n32881_, new_n32882_, new_n32883_, new_n32884_,
    new_n32885_, new_n32886_, new_n32887_, new_n32888_, new_n32889_,
    new_n32890_, new_n32891_, new_n32892_, new_n32893_, new_n32894_,
    new_n32895_, new_n32896_, new_n32897_, new_n32898_, new_n32899_,
    new_n32900_, new_n32901_, new_n32902_, new_n32903_, new_n32904_,
    new_n32905_, new_n32906_, new_n32907_, new_n32908_, new_n32909_,
    new_n32910_, new_n32911_, new_n32912_, new_n32913_, new_n32914_,
    new_n32915_, new_n32916_, new_n32917_, new_n32918_, new_n32919_,
    new_n32920_, new_n32921_, new_n32922_, new_n32923_, new_n32924_,
    new_n32925_, new_n32926_, new_n32927_, new_n32928_, new_n32929_,
    new_n32930_, new_n32931_, new_n32932_, new_n32933_, new_n32934_,
    new_n32935_, new_n32936_, new_n32937_, new_n32938_, new_n32939_,
    new_n32940_, new_n32941_, new_n32942_, new_n32943_, new_n32944_,
    new_n32945_, new_n32946_, new_n32947_, new_n32948_, new_n32949_,
    new_n32950_, new_n32951_, new_n32952_, new_n32953_, new_n32954_,
    new_n32955_, new_n32956_, new_n32957_, new_n32958_, new_n32959_,
    new_n32960_, new_n32961_, new_n32962_, new_n32963_, new_n32964_,
    new_n32965_, new_n32966_, new_n32967_, new_n32968_, new_n32969_,
    new_n32970_, new_n32971_, new_n32972_, new_n32973_, new_n32974_,
    new_n32975_, new_n32976_, new_n32977_, new_n32978_, new_n32979_,
    new_n32980_, new_n32981_, new_n32982_, new_n32983_, new_n32984_,
    new_n32985_, new_n32986_, new_n32987_, new_n32988_, new_n32989_,
    new_n32990_, new_n32991_, new_n32992_, new_n32993_, new_n32994_,
    new_n32995_, new_n32996_, new_n32997_, new_n32998_, new_n32999_,
    new_n33000_, new_n33001_, new_n33002_, new_n33003_, new_n33004_,
    new_n33005_, new_n33006_, new_n33007_, new_n33008_, new_n33009_,
    new_n33010_, new_n33011_, new_n33012_, new_n33013_, new_n33014_,
    new_n33015_, new_n33016_, new_n33017_, new_n33018_, new_n33019_,
    new_n33020_, new_n33021_, new_n33022_, new_n33023_, new_n33024_,
    new_n33025_, new_n33026_, new_n33027_, new_n33028_, new_n33029_,
    new_n33030_, new_n33031_, new_n33032_, new_n33033_, new_n33034_,
    new_n33035_, new_n33036_, new_n33037_, new_n33038_, new_n33039_,
    new_n33040_, new_n33041_, new_n33042_, new_n33043_, new_n33044_,
    new_n33045_, new_n33046_, new_n33047_, new_n33048_, new_n33049_,
    new_n33050_, new_n33051_, new_n33052_, new_n33053_, new_n33054_,
    new_n33055_, new_n33056_, new_n33057_, new_n33058_, new_n33059_,
    new_n33060_, new_n33061_, new_n33062_, new_n33063_, new_n33064_,
    new_n33065_, new_n33066_, new_n33067_, new_n33068_, new_n33069_,
    new_n33070_, new_n33071_, new_n33072_, new_n33073_, new_n33074_,
    new_n33075_, new_n33076_, new_n33077_, new_n33078_, new_n33079_,
    new_n33080_, new_n33081_, new_n33082_, new_n33083_, new_n33084_,
    new_n33085_, new_n33086_, new_n33087_, new_n33088_, new_n33089_,
    new_n33090_, new_n33091_, new_n33092_, new_n33093_, new_n33094_,
    new_n33095_, new_n33096_, new_n33097_, new_n33098_, new_n33099_,
    new_n33100_, new_n33101_, new_n33102_, new_n33103_, new_n33104_,
    new_n33105_, new_n33106_, new_n33107_, new_n33108_, new_n33109_,
    new_n33110_, new_n33111_, new_n33112_, new_n33113_, new_n33114_,
    new_n33115_, new_n33116_, new_n33117_, new_n33118_, new_n33119_,
    new_n33120_, new_n33121_, new_n33122_, new_n33123_, new_n33124_,
    new_n33125_, new_n33126_, new_n33127_, new_n33128_, new_n33129_,
    new_n33130_, new_n33131_, new_n33132_, new_n33133_, new_n33134_,
    new_n33135_, new_n33136_, new_n33137_, new_n33138_, new_n33139_,
    new_n33140_, new_n33141_, new_n33142_, new_n33143_, new_n33144_,
    new_n33145_, new_n33146_, new_n33147_, new_n33148_, new_n33149_,
    new_n33150_, new_n33151_, new_n33152_, new_n33153_, new_n33154_,
    new_n33155_, new_n33156_, new_n33157_, new_n33158_, new_n33159_,
    new_n33160_, new_n33161_, new_n33162_, new_n33163_, new_n33164_,
    new_n33165_, new_n33166_, new_n33167_, new_n33168_, new_n33169_,
    new_n33170_, new_n33171_, new_n33172_, new_n33173_, new_n33174_,
    new_n33175_, new_n33176_, new_n33177_, new_n33178_, new_n33179_,
    new_n33180_, new_n33181_, new_n33182_, new_n33183_, new_n33184_,
    new_n33185_, new_n33186_, new_n33187_, new_n33188_, new_n33189_,
    new_n33190_, new_n33191_, new_n33192_, new_n33193_, new_n33195_,
    new_n33196_, new_n33197_, new_n33198_, new_n33199_, new_n33200_,
    new_n33201_, new_n33202_, new_n33203_, new_n33204_, new_n33205_,
    new_n33206_, new_n33207_, new_n33208_, new_n33209_, new_n33210_,
    new_n33211_, new_n33212_, new_n33213_, new_n33214_, new_n33215_,
    new_n33216_, new_n33217_, new_n33218_, new_n33219_, new_n33220_,
    new_n33221_, new_n33222_, new_n33223_, new_n33224_, new_n33225_,
    new_n33226_, new_n33227_, new_n33228_, new_n33229_, new_n33230_,
    new_n33231_, new_n33232_, new_n33233_, new_n33234_, new_n33235_,
    new_n33236_, new_n33237_, new_n33238_, new_n33239_, new_n33240_,
    new_n33241_, new_n33242_, new_n33243_, new_n33245_, new_n33246_,
    new_n33247_, new_n33248_, new_n33249_, new_n33250_, new_n33251_,
    new_n33252_, new_n33253_, new_n33254_, new_n33255_, new_n33256_,
    new_n33257_, new_n33258_, new_n33259_, new_n33260_, new_n33261_,
    new_n33262_, new_n33263_, new_n33264_, new_n33265_, new_n33266_,
    new_n33267_, new_n33268_, new_n33269_, new_n33270_, new_n33271_,
    new_n33272_, new_n33273_, new_n33274_, new_n33275_, new_n33276_,
    new_n33277_, new_n33278_, new_n33279_, new_n33280_, new_n33281_,
    new_n33282_, new_n33283_, new_n33284_, new_n33285_, new_n33286_,
    new_n33287_, new_n33288_, new_n33289_, new_n33290_, new_n33291_,
    new_n33292_, new_n33293_, new_n33294_, new_n33295_, new_n33296_,
    new_n33297_, new_n33298_, new_n33299_, new_n33300_, new_n33301_,
    new_n33302_, new_n33303_, new_n33304_, new_n33305_, new_n33306_,
    new_n33307_, new_n33308_, new_n33309_, new_n33310_, new_n33311_,
    new_n33312_, new_n33314_, new_n33315_, new_n33316_, new_n33317_,
    new_n33318_, new_n33319_, new_n33320_, new_n33321_, new_n33322_,
    new_n33323_, new_n33324_, new_n33325_, new_n33326_, new_n33327_,
    new_n33328_, new_n33329_, new_n33330_, new_n33331_, new_n33332_,
    new_n33333_, new_n33334_, new_n33335_, new_n33336_, new_n33337_,
    new_n33338_, new_n33339_, new_n33340_, new_n33341_, new_n33342_,
    new_n33343_, new_n33344_, new_n33345_, new_n33346_, new_n33347_,
    new_n33348_, new_n33349_, new_n33350_, new_n33351_, new_n33352_,
    new_n33353_, new_n33354_, new_n33355_, new_n33356_, new_n33357_,
    new_n33358_, new_n33359_, new_n33360_, new_n33361_, new_n33362_,
    new_n33363_, new_n33364_, new_n33365_, new_n33366_, new_n33367_,
    new_n33368_, new_n33369_, new_n33370_, new_n33371_, new_n33372_,
    new_n33373_, new_n33375_, new_n33376_, new_n33377_, new_n33378_,
    new_n33379_, new_n33380_, new_n33381_, new_n33382_, new_n33383_,
    new_n33384_, new_n33385_, new_n33386_, new_n33387_, new_n33388_,
    new_n33389_, new_n33390_, new_n33391_, new_n33392_, new_n33393_,
    new_n33394_, new_n33395_, new_n33396_, new_n33397_, new_n33398_,
    new_n33399_, new_n33400_, new_n33401_, new_n33402_, new_n33403_,
    new_n33404_, new_n33405_, new_n33406_, new_n33407_, new_n33408_,
    new_n33409_, new_n33410_, new_n33411_, new_n33412_, new_n33413_,
    new_n33414_, new_n33415_, new_n33416_, new_n33417_, new_n33418_,
    new_n33419_, new_n33420_, new_n33421_, new_n33422_, new_n33423_,
    new_n33424_, new_n33425_, new_n33426_, new_n33427_, new_n33428_,
    new_n33429_, new_n33430_, new_n33431_, new_n33432_, new_n33433_,
    new_n33434_, new_n33435_, new_n33436_, new_n33437_, new_n33438_,
    new_n33439_, new_n33440_, new_n33441_, new_n33442_, new_n33443_,
    new_n33444_, new_n33445_, new_n33446_, new_n33447_, new_n33448_,
    new_n33449_, new_n33450_, new_n33451_, new_n33452_, new_n33453_,
    new_n33454_, new_n33455_, new_n33456_, new_n33457_, new_n33458_,
    new_n33459_, new_n33460_, new_n33461_, new_n33462_, new_n33463_,
    new_n33464_, new_n33465_, new_n33466_, new_n33467_, new_n33468_,
    new_n33469_, new_n33470_, new_n33471_, new_n33472_, new_n33473_,
    new_n33474_, new_n33475_, new_n33476_, new_n33477_, new_n33478_,
    new_n33479_, new_n33480_, new_n33481_, new_n33482_, new_n33483_,
    new_n33484_, new_n33485_, new_n33486_, new_n33487_, new_n33488_,
    new_n33489_, new_n33490_, new_n33491_, new_n33492_, new_n33493_,
    new_n33494_, new_n33495_, new_n33496_, new_n33497_, new_n33498_,
    new_n33499_, new_n33500_, new_n33501_, new_n33502_, new_n33503_,
    new_n33504_, new_n33505_, new_n33506_, new_n33507_, new_n33508_,
    new_n33509_, new_n33510_, new_n33511_, new_n33512_, new_n33513_,
    new_n33514_, new_n33515_, new_n33516_, new_n33517_, new_n33518_,
    new_n33519_, new_n33520_, new_n33521_, new_n33522_, new_n33523_,
    new_n33524_, new_n33525_, new_n33526_, new_n33527_, new_n33528_,
    new_n33529_, new_n33530_, new_n33531_, new_n33532_, new_n33533_,
    new_n33534_, new_n33535_, new_n33536_, new_n33537_, new_n33538_,
    new_n33539_, new_n33540_, new_n33541_, new_n33542_, new_n33543_,
    new_n33544_, new_n33545_, new_n33546_, new_n33547_, new_n33548_,
    new_n33549_, new_n33550_, new_n33551_, new_n33552_, new_n33553_,
    new_n33554_, new_n33555_, new_n33556_, new_n33557_, new_n33558_,
    new_n33559_, new_n33560_, new_n33561_, new_n33562_, new_n33563_,
    new_n33564_, new_n33565_, new_n33566_, new_n33567_, new_n33568_,
    new_n33569_, new_n33570_, new_n33571_, new_n33572_, new_n33573_,
    new_n33574_, new_n33575_, new_n33576_, new_n33577_, new_n33578_,
    new_n33579_, new_n33580_, new_n33581_, new_n33582_, new_n33583_,
    new_n33584_, new_n33585_, new_n33586_, new_n33587_, new_n33588_,
    new_n33589_, new_n33590_, new_n33591_, new_n33592_, new_n33593_,
    new_n33594_, new_n33595_, new_n33596_, new_n33597_, new_n33598_,
    new_n33599_, new_n33600_, new_n33601_, new_n33602_, new_n33603_,
    new_n33604_, new_n33605_, new_n33606_, new_n33607_, new_n33608_,
    new_n33609_, new_n33610_, new_n33611_, new_n33612_, new_n33613_,
    new_n33614_, new_n33615_, new_n33616_, new_n33617_, new_n33618_,
    new_n33619_, new_n33620_, new_n33621_, new_n33622_, new_n33623_,
    new_n33624_, new_n33625_, new_n33626_, new_n33627_, new_n33628_,
    new_n33629_, new_n33630_, new_n33631_, new_n33632_, new_n33633_,
    new_n33634_, new_n33635_, new_n33636_, new_n33637_, new_n33638_,
    new_n33639_, new_n33640_, new_n33641_, new_n33642_, new_n33643_,
    new_n33644_, new_n33645_, new_n33646_, new_n33647_, new_n33648_,
    new_n33649_, new_n33650_, new_n33651_, new_n33652_, new_n33653_,
    new_n33654_, new_n33655_, new_n33656_, new_n33657_, new_n33658_,
    new_n33659_, new_n33660_, new_n33661_, new_n33662_, new_n33663_,
    new_n33664_, new_n33665_, new_n33666_, new_n33667_, new_n33668_,
    new_n33669_, new_n33670_, new_n33671_, new_n33672_, new_n33673_,
    new_n33674_, new_n33675_, new_n33676_, new_n33677_, new_n33678_,
    new_n33679_, new_n33680_, new_n33681_, new_n33682_, new_n33683_,
    new_n33684_, new_n33685_, new_n33686_, new_n33687_, new_n33688_,
    new_n33689_, new_n33690_, new_n33691_, new_n33692_, new_n33693_,
    new_n33694_, new_n33695_, new_n33696_, new_n33697_, new_n33698_,
    new_n33699_, new_n33700_, new_n33701_, new_n33702_, new_n33703_,
    new_n33704_, new_n33705_, new_n33706_, new_n33707_, new_n33708_,
    new_n33709_, new_n33710_, new_n33711_, new_n33712_, new_n33713_,
    new_n33714_, new_n33715_, new_n33716_, new_n33717_, new_n33718_,
    new_n33719_, new_n33720_, new_n33721_, new_n33722_, new_n33723_,
    new_n33724_, new_n33725_, new_n33726_, new_n33727_, new_n33728_,
    new_n33729_, new_n33730_, new_n33731_, new_n33732_, new_n33733_,
    new_n33734_, new_n33735_, new_n33736_, new_n33737_, new_n33738_,
    new_n33739_, new_n33740_, new_n33741_, new_n33742_, new_n33743_,
    new_n33744_, new_n33745_, new_n33746_, new_n33747_, new_n33748_,
    new_n33749_, new_n33750_, new_n33751_, new_n33752_, new_n33753_,
    new_n33754_, new_n33755_, new_n33756_, new_n33757_, new_n33758_,
    new_n33759_, new_n33760_, new_n33761_, new_n33762_, new_n33763_,
    new_n33764_, new_n33765_, new_n33766_, new_n33767_, new_n33768_,
    new_n33769_, new_n33770_, new_n33771_, new_n33772_, new_n33773_,
    new_n33774_, new_n33775_, new_n33776_, new_n33777_, new_n33778_,
    new_n33779_, new_n33780_, new_n33781_, new_n33782_, new_n33783_,
    new_n33784_, new_n33785_, new_n33786_, new_n33787_, new_n33788_,
    new_n33789_, new_n33790_, new_n33791_, new_n33792_, new_n33793_,
    new_n33794_, new_n33795_, new_n33796_, new_n33797_, new_n33798_,
    new_n33799_, new_n33800_, new_n33801_, new_n33802_, new_n33803_,
    new_n33804_, new_n33805_, new_n33806_, new_n33807_, new_n33808_,
    new_n33809_, new_n33810_, new_n33811_, new_n33812_, new_n33813_,
    new_n33814_, new_n33815_, new_n33816_, new_n33817_, new_n33818_,
    new_n33819_, new_n33820_, new_n33821_, new_n33822_, new_n33823_,
    new_n33824_, new_n33825_, new_n33826_, new_n33827_, new_n33828_,
    new_n33829_, new_n33830_, new_n33831_, new_n33832_, new_n33833_,
    new_n33834_, new_n33835_, new_n33836_, new_n33837_, new_n33838_,
    new_n33839_, new_n33840_, new_n33841_, new_n33842_, new_n33843_,
    new_n33844_, new_n33845_, new_n33846_, new_n33847_, new_n33848_,
    new_n33849_, new_n33850_, new_n33851_, new_n33852_, new_n33853_,
    new_n33854_, new_n33855_, new_n33856_, new_n33857_, new_n33858_,
    new_n33859_, new_n33860_, new_n33861_, new_n33862_, new_n33863_,
    new_n33864_, new_n33865_, new_n33866_, new_n33867_, new_n33868_,
    new_n33869_, new_n33870_, new_n33871_, new_n33872_, new_n33873_,
    new_n33874_, new_n33875_, new_n33876_, new_n33877_, new_n33878_,
    new_n33879_, new_n33880_, new_n33881_, new_n33882_, new_n33883_,
    new_n33884_, new_n33885_, new_n33886_, new_n33887_, new_n33888_,
    new_n33889_, new_n33890_, new_n33891_, new_n33892_, new_n33893_,
    new_n33894_, new_n33895_, new_n33896_, new_n33897_, new_n33898_,
    new_n33899_, new_n33900_, new_n33901_, new_n33902_, new_n33903_,
    new_n33904_, new_n33905_, new_n33906_, new_n33907_, new_n33908_,
    new_n33909_, new_n33910_, new_n33911_, new_n33912_, new_n33913_,
    new_n33914_, new_n33915_, new_n33916_, new_n33917_, new_n33918_,
    new_n33919_, new_n33920_, new_n33921_, new_n33922_, new_n33923_,
    new_n33924_, new_n33925_, new_n33926_, new_n33927_, new_n33928_,
    new_n33929_, new_n33930_, new_n33931_, new_n33932_, new_n33933_,
    new_n33934_, new_n33935_, new_n33936_, new_n33937_, new_n33938_,
    new_n33939_, new_n33940_, new_n33941_, new_n33942_, new_n33943_,
    new_n33944_, new_n33945_, new_n33946_, new_n33947_, new_n33948_,
    new_n33949_, new_n33950_, new_n33951_, new_n33952_, new_n33953_,
    new_n33954_, new_n33955_, new_n33956_, new_n33957_, new_n33958_,
    new_n33959_, new_n33960_, new_n33961_, new_n33962_, new_n33963_,
    new_n33964_, new_n33965_, new_n33966_, new_n33967_, new_n33968_,
    new_n33969_, new_n33970_, new_n33971_, new_n33972_, new_n33973_,
    new_n33974_, new_n33975_, new_n33976_, new_n33977_, new_n33978_,
    new_n33979_, new_n33980_, new_n33981_, new_n33982_, new_n33983_,
    new_n33984_, new_n33985_, new_n33986_, new_n33987_, new_n33988_,
    new_n33989_, new_n33990_, new_n33991_, new_n33992_, new_n33993_,
    new_n33994_, new_n33995_, new_n33996_, new_n33997_, new_n33998_,
    new_n33999_, new_n34000_, new_n34001_, new_n34002_, new_n34003_,
    new_n34004_, new_n34005_, new_n34006_, new_n34007_, new_n34008_,
    new_n34009_, new_n34011_, new_n34012_, new_n34013_, new_n34014_,
    new_n34015_, new_n34016_, new_n34017_, new_n34018_, new_n34019_,
    new_n34020_, new_n34021_, new_n34022_, new_n34023_, new_n34024_,
    new_n34025_, new_n34026_, new_n34027_, new_n34028_, new_n34029_,
    new_n34030_, new_n34031_, new_n34032_, new_n34033_, new_n34034_,
    new_n34035_, new_n34036_, new_n34037_, new_n34038_, new_n34039_,
    new_n34040_, new_n34041_, new_n34042_, new_n34043_, new_n34044_,
    new_n34045_, new_n34046_, new_n34047_, new_n34048_, new_n34049_,
    new_n34050_, new_n34051_, new_n34052_, new_n34053_, new_n34054_,
    new_n34055_, new_n34056_, new_n34057_, new_n34058_, new_n34059_,
    new_n34060_, new_n34061_, new_n34062_, new_n34063_, new_n34064_,
    new_n34065_, new_n34066_, new_n34067_, new_n34068_, new_n34069_,
    new_n34070_, new_n34071_, new_n34072_, new_n34073_, new_n34074_,
    new_n34075_, new_n34076_, new_n34077_, new_n34078_, new_n34079_,
    new_n34080_, new_n34081_, new_n34082_, new_n34083_, new_n34084_,
    new_n34085_, new_n34086_, new_n34087_, new_n34088_, new_n34089_,
    new_n34090_, new_n34091_, new_n34092_, new_n34093_, new_n34094_,
    new_n34095_, new_n34096_, new_n34097_, new_n34098_, new_n34099_,
    new_n34100_, new_n34101_, new_n34102_, new_n34103_, new_n34104_,
    new_n34105_, new_n34106_, new_n34107_, new_n34108_, new_n34109_,
    new_n34110_, new_n34111_, new_n34112_, new_n34113_, new_n34114_,
    new_n34115_, new_n34116_, new_n34117_, new_n34118_, new_n34119_,
    new_n34120_, new_n34121_, new_n34122_, new_n34123_, new_n34124_,
    new_n34125_, new_n34126_, new_n34127_, new_n34128_, new_n34129_,
    new_n34130_, new_n34131_, new_n34132_, new_n34133_, new_n34134_,
    new_n34135_, new_n34136_, new_n34137_, new_n34138_, new_n34139_,
    new_n34140_, new_n34141_, new_n34142_, new_n34143_, new_n34144_,
    new_n34145_, new_n34146_, new_n34147_, new_n34148_, new_n34149_,
    new_n34150_, new_n34151_, new_n34152_, new_n34153_, new_n34154_,
    new_n34155_, new_n34156_, new_n34157_, new_n34158_, new_n34159_,
    new_n34160_, new_n34161_, new_n34162_, new_n34163_, new_n34164_,
    new_n34165_, new_n34166_, new_n34167_, new_n34168_, new_n34169_,
    new_n34170_, new_n34171_, new_n34172_, new_n34173_, new_n34174_,
    new_n34175_, new_n34176_, new_n34177_, new_n34178_, new_n34179_,
    new_n34180_, new_n34181_, new_n34182_, new_n34183_, new_n34184_,
    new_n34185_, new_n34186_, new_n34187_, new_n34188_, new_n34189_,
    new_n34190_, new_n34191_, new_n34192_, new_n34193_, new_n34194_,
    new_n34195_, new_n34196_, new_n34197_, new_n34198_, new_n34199_,
    new_n34200_, new_n34201_, new_n34202_, new_n34203_, new_n34204_,
    new_n34205_, new_n34206_, new_n34207_, new_n34208_, new_n34209_,
    new_n34210_, new_n34211_, new_n34212_, new_n34213_, new_n34214_,
    new_n34215_, new_n34216_, new_n34217_, new_n34218_, new_n34219_,
    new_n34220_, new_n34221_, new_n34222_, new_n34223_, new_n34224_,
    new_n34225_, new_n34226_, new_n34227_, new_n34228_, new_n34229_,
    new_n34230_, new_n34231_, new_n34232_, new_n34233_, new_n34234_,
    new_n34235_, new_n34236_, new_n34237_, new_n34238_, new_n34239_,
    new_n34240_, new_n34241_, new_n34242_, new_n34243_, new_n34244_,
    new_n34245_, new_n34246_, new_n34247_, new_n34248_, new_n34249_,
    new_n34250_, new_n34251_, new_n34252_, new_n34253_, new_n34254_,
    new_n34255_, new_n34256_, new_n34257_, new_n34258_, new_n34259_,
    new_n34260_, new_n34261_, new_n34262_, new_n34263_, new_n34264_,
    new_n34265_, new_n34266_, new_n34267_, new_n34268_, new_n34269_,
    new_n34270_, new_n34271_, new_n34272_, new_n34273_, new_n34274_,
    new_n34275_, new_n34276_, new_n34277_, new_n34278_, new_n34279_,
    new_n34280_, new_n34281_, new_n34282_, new_n34283_, new_n34284_,
    new_n34285_, new_n34286_, new_n34287_, new_n34288_, new_n34289_,
    new_n34290_, new_n34291_, new_n34292_, new_n34293_, new_n34294_,
    new_n34295_, new_n34296_, new_n34297_, new_n34298_, new_n34299_,
    new_n34300_, new_n34302_, new_n34303_, new_n34304_, new_n34305_,
    new_n34306_, new_n34307_, new_n34308_, new_n34309_, new_n34310_,
    new_n34311_, new_n34312_, new_n34313_, new_n34314_, new_n34315_,
    new_n34316_, new_n34317_, new_n34318_, new_n34319_, new_n34320_,
    new_n34321_, new_n34322_, new_n34323_, new_n34324_, new_n34325_,
    new_n34326_, new_n34327_, new_n34328_, new_n34329_, new_n34330_,
    new_n34331_, new_n34332_, new_n34333_, new_n34334_, new_n34335_,
    new_n34336_, new_n34337_, new_n34338_, new_n34339_, new_n34340_,
    new_n34341_, new_n34342_, new_n34343_, new_n34344_, new_n34345_,
    new_n34346_, new_n34347_, new_n34348_, new_n34349_, new_n34350_,
    new_n34351_, new_n34352_, new_n34353_, new_n34354_, new_n34355_,
    new_n34356_, new_n34357_, new_n34358_, new_n34359_, new_n34360_,
    new_n34361_, new_n34362_, new_n34363_, new_n34364_, new_n34365_,
    new_n34366_, new_n34367_, new_n34368_, new_n34369_, new_n34370_,
    new_n34371_, new_n34372_, new_n34373_, new_n34374_, new_n34375_,
    new_n34376_, new_n34377_, new_n34378_, new_n34379_, new_n34380_,
    new_n34381_, new_n34382_, new_n34383_, new_n34384_, new_n34385_,
    new_n34386_, new_n34387_, new_n34388_, new_n34389_, new_n34390_,
    new_n34391_, new_n34392_, new_n34393_, new_n34394_, new_n34395_,
    new_n34396_, new_n34397_, new_n34398_, new_n34399_, new_n34400_,
    new_n34401_, new_n34402_, new_n34403_, new_n34404_, new_n34405_,
    new_n34406_, new_n34407_, new_n34408_, new_n34409_, new_n34410_,
    new_n34411_, new_n34412_, new_n34413_, new_n34414_, new_n34415_,
    new_n34416_, new_n34417_, new_n34418_, new_n34419_, new_n34420_,
    new_n34421_, new_n34422_, new_n34423_, new_n34424_, new_n34425_,
    new_n34426_, new_n34427_, new_n34428_, new_n34429_, new_n34430_,
    new_n34431_, new_n34432_, new_n34433_, new_n34434_, new_n34435_,
    new_n34436_, new_n34437_, new_n34438_, new_n34439_, new_n34440_,
    new_n34441_, new_n34442_, new_n34443_, new_n34444_, new_n34445_,
    new_n34446_, new_n34447_, new_n34448_, new_n34449_, new_n34450_,
    new_n34451_, new_n34452_, new_n34453_, new_n34454_, new_n34455_,
    new_n34456_, new_n34457_, new_n34458_, new_n34459_, new_n34460_,
    new_n34461_, new_n34462_, new_n34463_, new_n34464_, new_n34465_,
    new_n34466_, new_n34467_, new_n34468_, new_n34469_, new_n34470_,
    new_n34471_, new_n34472_, new_n34473_, new_n34474_, new_n34475_,
    new_n34476_, new_n34477_, new_n34478_, new_n34479_, new_n34480_,
    new_n34481_, new_n34482_, new_n34483_, new_n34484_, new_n34485_,
    new_n34486_, new_n34487_, new_n34488_, new_n34489_, new_n34490_,
    new_n34491_, new_n34492_, new_n34493_, new_n34494_, new_n34495_,
    new_n34496_, new_n34497_, new_n34498_, new_n34499_, new_n34500_,
    new_n34501_, new_n34502_, new_n34503_, new_n34504_, new_n34505_,
    new_n34506_, new_n34507_, new_n34508_, new_n34509_, new_n34510_,
    new_n34511_, new_n34512_, new_n34513_, new_n34514_, new_n34515_,
    new_n34516_, new_n34517_, new_n34518_, new_n34519_, new_n34520_,
    new_n34521_, new_n34522_, new_n34523_, new_n34524_, new_n34525_,
    new_n34526_, new_n34527_, new_n34528_, new_n34529_, new_n34530_,
    new_n34531_, new_n34532_, new_n34533_, new_n34534_, new_n34535_,
    new_n34536_, new_n34537_, new_n34538_, new_n34539_, new_n34540_,
    new_n34541_, new_n34542_, new_n34543_, new_n34544_, new_n34545_,
    new_n34546_, new_n34547_, new_n34548_, new_n34549_, new_n34550_,
    new_n34551_, new_n34552_, new_n34553_, new_n34554_, new_n34555_,
    new_n34556_, new_n34557_, new_n34558_, new_n34559_, new_n34560_,
    new_n34561_, new_n34562_, new_n34563_, new_n34564_, new_n34565_,
    new_n34566_, new_n34567_, new_n34568_, new_n34569_, new_n34570_,
    new_n34571_, new_n34572_, new_n34573_, new_n34574_, new_n34575_,
    new_n34576_, new_n34577_, new_n34578_, new_n34579_, new_n34580_,
    new_n34581_, new_n34583_, new_n34584_, new_n34585_, new_n34586_,
    new_n34587_, new_n34588_, new_n34589_, new_n34590_, new_n34591_,
    new_n34592_, new_n34593_, new_n34594_, new_n34595_, new_n34596_,
    new_n34597_, new_n34598_, new_n34599_, new_n34600_, new_n34601_,
    new_n34602_, new_n34603_, new_n34604_, new_n34605_, new_n34606_,
    new_n34607_, new_n34608_, new_n34609_, new_n34610_, new_n34611_,
    new_n34612_, new_n34613_, new_n34614_, new_n34615_, new_n34616_,
    new_n34617_, new_n34618_, new_n34619_, new_n34620_, new_n34621_,
    new_n34622_, new_n34623_, new_n34624_, new_n34625_, new_n34626_,
    new_n34627_, new_n34628_, new_n34629_, new_n34630_, new_n34631_,
    new_n34632_, new_n34633_, new_n34634_, new_n34635_, new_n34636_,
    new_n34637_, new_n34638_, new_n34639_, new_n34640_, new_n34641_,
    new_n34642_, new_n34643_, new_n34644_, new_n34645_, new_n34646_,
    new_n34647_, new_n34648_, new_n34649_, new_n34650_, new_n34651_,
    new_n34652_, new_n34653_, new_n34654_, new_n34655_, new_n34656_,
    new_n34657_, new_n34658_, new_n34659_, new_n34660_, new_n34661_,
    new_n34662_, new_n34663_, new_n34664_, new_n34665_, new_n34666_,
    new_n34667_, new_n34668_, new_n34669_, new_n34670_, new_n34671_,
    new_n34672_, new_n34673_, new_n34674_, new_n34675_, new_n34676_,
    new_n34677_, new_n34678_, new_n34679_, new_n34680_, new_n34681_,
    new_n34682_, new_n34683_, new_n34684_, new_n34685_, new_n34686_,
    new_n34687_, new_n34688_, new_n34689_, new_n34690_, new_n34691_,
    new_n34692_, new_n34693_, new_n34694_, new_n34695_, new_n34696_,
    new_n34697_, new_n34698_, new_n34699_, new_n34700_, new_n34701_,
    new_n34702_, new_n34703_, new_n34704_, new_n34705_, new_n34706_,
    new_n34707_, new_n34708_, new_n34709_, new_n34710_, new_n34711_,
    new_n34712_, new_n34713_, new_n34714_, new_n34715_, new_n34716_,
    new_n34717_, new_n34718_, new_n34719_, new_n34720_, new_n34721_,
    new_n34722_, new_n34723_, new_n34724_, new_n34725_, new_n34726_,
    new_n34727_, new_n34728_, new_n34729_, new_n34730_, new_n34731_,
    new_n34732_, new_n34733_, new_n34734_, new_n34735_, new_n34736_,
    new_n34737_, new_n34738_, new_n34739_, new_n34740_, new_n34741_,
    new_n34742_, new_n34743_, new_n34744_, new_n34745_, new_n34746_,
    new_n34747_, new_n34748_, new_n34749_, new_n34750_, new_n34751_,
    new_n34752_, new_n34753_, new_n34754_, new_n34755_, new_n34756_,
    new_n34757_, new_n34758_, new_n34759_, new_n34760_, new_n34761_,
    new_n34762_, new_n34763_, new_n34764_, new_n34765_, new_n34766_,
    new_n34767_, new_n34768_, new_n34769_, new_n34770_, new_n34771_,
    new_n34772_, new_n34773_, new_n34774_, new_n34775_, new_n34776_,
    new_n34778_, new_n34779_, new_n34780_, new_n34781_, new_n34782_,
    new_n34783_, new_n34784_, new_n34786_, new_n34787_, new_n34788_,
    new_n34789_, new_n34790_, new_n34791_, new_n34792_, new_n34794_,
    new_n34795_, new_n34796_, new_n34797_, new_n34798_, new_n34799_,
    new_n34800_, new_n34801_, new_n34802_, new_n34803_, new_n34804_,
    new_n34805_, new_n34806_, new_n34807_, new_n34808_, new_n34809_,
    new_n34810_, new_n34811_, new_n34812_, new_n34813_, new_n34814_,
    new_n34815_, new_n34816_, new_n34817_, new_n34818_, new_n34819_,
    new_n34820_, new_n34821_, new_n34822_, new_n34823_, new_n34824_,
    new_n34825_, new_n34826_, new_n34827_, new_n34828_, new_n34829_,
    new_n34830_, new_n34831_, new_n34832_, new_n34833_, new_n34834_,
    new_n34835_, new_n34836_, new_n34837_, new_n34838_, new_n34839_,
    new_n34840_, new_n34841_, new_n34842_, new_n34843_, new_n34844_,
    new_n34845_, new_n34846_, new_n34847_, new_n34848_, new_n34849_,
    new_n34850_, new_n34851_, new_n34852_, new_n34853_, new_n34854_,
    new_n34855_, new_n34856_, new_n34857_, new_n34858_, new_n34859_,
    new_n34860_, new_n34861_, new_n34862_, new_n34863_, new_n34864_,
    new_n34865_, new_n34866_, new_n34867_, new_n34868_, new_n34869_,
    new_n34870_, new_n34871_, new_n34872_, new_n34873_, new_n34874_,
    new_n34875_, new_n34876_, new_n34877_, new_n34878_, new_n34879_,
    new_n34880_, new_n34881_, new_n34882_, new_n34883_, new_n34884_,
    new_n34885_, new_n34886_, new_n34887_, new_n34888_, new_n34889_,
    new_n34890_, new_n34891_, new_n34892_, new_n34893_, new_n34894_,
    new_n34895_, new_n34896_, new_n34897_, new_n34898_, new_n34899_,
    new_n34900_, new_n34901_, new_n34903_, new_n34904_, new_n34905_,
    new_n34906_, new_n34907_, new_n34908_, new_n34910_, new_n34911_,
    new_n34912_, new_n34913_, new_n34914_, new_n34915_, new_n34916_,
    new_n34918_, new_n34919_, new_n34920_, new_n34921_, new_n34922_,
    new_n34923_, new_n34924_, new_n34925_, new_n34926_, new_n34927_,
    new_n34928_, new_n34929_, new_n34930_, new_n34931_, new_n34932_,
    new_n34933_, new_n34934_, new_n34935_, new_n34936_, new_n34937_,
    new_n34938_, new_n34939_, new_n34940_, new_n34941_, new_n34942_,
    new_n34943_, new_n34944_, new_n34945_, new_n34946_, new_n34947_,
    new_n34948_, new_n34949_, new_n34950_, new_n34951_, new_n34952_,
    new_n34953_, new_n34954_, new_n34955_, new_n34956_, new_n34957_,
    new_n34958_, new_n34959_, new_n34960_, new_n34961_, new_n34962_,
    new_n34963_, new_n34964_, new_n34965_, new_n34966_, new_n34967_,
    new_n34968_, new_n34969_, new_n34970_, new_n34971_, new_n34972_,
    new_n34973_, new_n34974_, new_n34975_, new_n34976_, new_n34977_,
    new_n34978_, new_n34979_, new_n34980_, new_n34981_, new_n34982_,
    new_n34983_, new_n34984_, new_n34985_, new_n34986_, new_n34987_,
    new_n34988_, new_n34989_, new_n34990_, new_n34991_, new_n34992_,
    new_n34993_, new_n34994_, new_n34995_, new_n34996_, new_n34997_,
    new_n34998_, new_n34999_, new_n35000_, new_n35001_, new_n35002_,
    new_n35003_, new_n35004_, new_n35005_, new_n35006_, new_n35007_,
    new_n35008_, new_n35009_, new_n35010_, new_n35011_, new_n35012_,
    new_n35013_, new_n35014_, new_n35015_, new_n35016_, new_n35017_,
    new_n35018_, new_n35019_, new_n35020_, new_n35021_, new_n35022_,
    new_n35023_, new_n35024_, new_n35025_, new_n35026_, new_n35027_,
    new_n35028_, new_n35029_, new_n35030_, new_n35031_, new_n35032_,
    new_n35033_, new_n35034_, new_n35035_, new_n35036_, new_n35037_,
    new_n35038_, new_n35039_, new_n35040_, new_n35041_, new_n35042_,
    new_n35043_, new_n35044_, new_n35045_, new_n35046_, new_n35047_,
    new_n35048_, new_n35049_, new_n35050_, new_n35051_, new_n35052_,
    new_n35053_, new_n35054_, new_n35055_, new_n35056_, new_n35057_,
    new_n35058_, new_n35059_, new_n35060_, new_n35061_, new_n35062_,
    new_n35063_, new_n35064_, new_n35065_, new_n35066_, new_n35067_,
    new_n35068_, new_n35069_, new_n35070_, new_n35071_, new_n35072_,
    new_n35073_, new_n35074_, new_n35075_, new_n35076_, new_n35077_,
    new_n35078_, new_n35079_, new_n35080_, new_n35081_, new_n35082_,
    new_n35083_, new_n35084_, new_n35085_, new_n35086_, new_n35087_,
    new_n35088_, new_n35089_, new_n35090_, new_n35091_, new_n35092_,
    new_n35093_, new_n35094_, new_n35095_, new_n35096_, new_n35097_,
    new_n35098_, new_n35099_, new_n35100_, new_n35101_, new_n35102_,
    new_n35103_, new_n35104_, new_n35105_, new_n35106_, new_n35107_,
    new_n35108_, new_n35109_, new_n35110_, new_n35111_, new_n35112_,
    new_n35113_, new_n35114_, new_n35115_, new_n35116_, new_n35117_,
    new_n35118_, new_n35119_, new_n35120_, new_n35121_, new_n35122_,
    new_n35123_, new_n35124_, new_n35125_, new_n35126_, new_n35127_,
    new_n35128_, new_n35129_, new_n35130_, new_n35131_, new_n35132_,
    new_n35133_, new_n35134_, new_n35135_, new_n35136_, new_n35137_,
    new_n35138_, new_n35139_, new_n35140_, new_n35141_, new_n35142_,
    new_n35143_, new_n35144_, new_n35145_, new_n35146_, new_n35147_,
    new_n35148_, new_n35149_, new_n35150_, new_n35151_, new_n35152_,
    new_n35153_, new_n35154_, new_n35155_, new_n35156_, new_n35157_,
    new_n35158_, new_n35159_, new_n35160_, new_n35161_, new_n35162_,
    new_n35163_, new_n35164_, new_n35165_, new_n35166_, new_n35167_,
    new_n35168_, new_n35169_, new_n35170_, new_n35171_, new_n35172_,
    new_n35173_, new_n35174_, new_n35175_, new_n35176_, new_n35177_,
    new_n35178_, new_n35179_, new_n35180_, new_n35181_, new_n35182_,
    new_n35183_, new_n35184_, new_n35185_, new_n35186_, new_n35187_,
    new_n35188_, new_n35189_, new_n35190_, new_n35191_, new_n35192_,
    new_n35193_, new_n35194_, new_n35195_, new_n35196_, new_n35197_,
    new_n35198_, new_n35199_, new_n35200_, new_n35201_, new_n35202_,
    new_n35203_, new_n35204_, new_n35205_, new_n35206_, new_n35207_,
    new_n35208_, new_n35209_, new_n35210_, new_n35211_, new_n35212_,
    new_n35213_, new_n35214_, new_n35215_, new_n35216_, new_n35217_,
    new_n35218_, new_n35219_, new_n35220_, new_n35221_, new_n35222_,
    new_n35223_, new_n35224_, new_n35225_, new_n35226_, new_n35227_,
    new_n35228_, new_n35229_, new_n35230_, new_n35231_, new_n35232_,
    new_n35233_, new_n35234_, new_n35235_, new_n35236_, new_n35237_,
    new_n35238_, new_n35239_, new_n35240_, new_n35241_, new_n35242_,
    new_n35243_, new_n35244_, new_n35245_, new_n35246_, new_n35247_,
    new_n35248_, new_n35249_, new_n35250_, new_n35251_, new_n35252_,
    new_n35253_, new_n35254_, new_n35255_, new_n35256_, new_n35257_,
    new_n35258_, new_n35259_, new_n35260_, new_n35261_, new_n35262_,
    new_n35263_, new_n35264_, new_n35265_, new_n35266_, new_n35267_,
    new_n35268_, new_n35269_, new_n35270_, new_n35271_, new_n35272_,
    new_n35273_, new_n35274_, new_n35275_, new_n35276_, new_n35277_,
    new_n35278_, new_n35279_, new_n35280_, new_n35281_, new_n35282_,
    new_n35283_, new_n35284_, new_n35285_, new_n35286_, new_n35287_,
    new_n35288_, new_n35289_, new_n35290_, new_n35291_, new_n35292_,
    new_n35293_, new_n35294_, new_n35295_, new_n35296_, new_n35297_,
    new_n35298_, new_n35299_, new_n35300_, new_n35301_, new_n35302_,
    new_n35303_, new_n35304_, new_n35305_, new_n35306_, new_n35307_,
    new_n35308_, new_n35309_, new_n35310_, new_n35311_, new_n35312_,
    new_n35313_, new_n35314_, new_n35315_, new_n35316_, new_n35317_,
    new_n35318_, new_n35319_, new_n35320_, new_n35321_, new_n35322_,
    new_n35323_, new_n35324_, new_n35325_, new_n35326_, new_n35327_,
    new_n35328_, new_n35329_, new_n35330_, new_n35331_, new_n35332_,
    new_n35333_, new_n35334_, new_n35335_, new_n35336_, new_n35337_,
    new_n35338_, new_n35339_, new_n35340_, new_n35341_, new_n35342_,
    new_n35343_, new_n35344_, new_n35345_, new_n35346_, new_n35347_,
    new_n35348_, new_n35349_, new_n35350_, new_n35351_, new_n35352_,
    new_n35353_, new_n35354_, new_n35355_, new_n35356_, new_n35357_,
    new_n35358_, new_n35359_, new_n35360_, new_n35361_, new_n35362_,
    new_n35363_, new_n35364_, new_n35365_, new_n35366_, new_n35367_,
    new_n35368_, new_n35369_, new_n35370_, new_n35371_, new_n35372_,
    new_n35373_, new_n35374_, new_n35375_, new_n35376_, new_n35377_,
    new_n35378_, new_n35379_, new_n35380_, new_n35381_, new_n35382_,
    new_n35383_, new_n35384_, new_n35385_, new_n35386_, new_n35387_,
    new_n35388_, new_n35389_, new_n35390_, new_n35391_, new_n35392_,
    new_n35393_, new_n35394_, new_n35395_, new_n35396_, new_n35397_,
    new_n35398_, new_n35399_, new_n35400_, new_n35401_, new_n35402_,
    new_n35403_, new_n35404_, new_n35405_, new_n35406_, new_n35407_,
    new_n35408_, new_n35410_, new_n35411_, new_n35412_, new_n35413_,
    new_n35414_, new_n35415_, new_n35416_, new_n35417_, new_n35418_,
    new_n35419_, new_n35420_, new_n35421_, new_n35422_, new_n35423_,
    new_n35424_, new_n35425_, new_n35426_, new_n35427_, new_n35428_,
    new_n35429_, new_n35430_, new_n35431_, new_n35432_, new_n35433_,
    new_n35434_, new_n35435_, new_n35436_, new_n35437_, new_n35438_,
    new_n35439_, new_n35440_, new_n35441_, new_n35442_, new_n35443_,
    new_n35444_, new_n35445_, new_n35446_, new_n35447_, new_n35448_,
    new_n35449_, new_n35450_, new_n35451_, new_n35452_, new_n35453_,
    new_n35454_, new_n35455_, new_n35456_, new_n35457_, new_n35458_,
    new_n35459_, new_n35460_, new_n35461_, new_n35462_, new_n35463_,
    new_n35464_, new_n35465_, new_n35466_, new_n35467_, new_n35468_,
    new_n35469_, new_n35470_, new_n35471_, new_n35472_, new_n35473_,
    new_n35474_, new_n35475_, new_n35476_, new_n35477_, new_n35478_,
    new_n35479_, new_n35480_, new_n35481_, new_n35482_, new_n35483_,
    new_n35485_, new_n35486_, new_n35487_, new_n35488_, new_n35489_,
    new_n35490_, new_n35491_, new_n35492_, new_n35493_, new_n35494_,
    new_n35495_, new_n35496_, new_n35497_, new_n35498_, new_n35499_,
    new_n35500_, new_n35501_, new_n35502_, new_n35503_, new_n35504_,
    new_n35505_, new_n35506_, new_n35507_, new_n35508_, new_n35509_,
    new_n35510_, new_n35511_, new_n35512_, new_n35513_, new_n35514_,
    new_n35515_, new_n35516_, new_n35517_, new_n35518_, new_n35519_,
    new_n35520_, new_n35521_, new_n35522_, new_n35523_, new_n35524_,
    new_n35525_, new_n35526_, new_n35527_, new_n35528_, new_n35529_,
    new_n35530_, new_n35531_, new_n35532_, new_n35533_, new_n35534_,
    new_n35535_, new_n35536_, new_n35537_, new_n35538_, new_n35539_,
    new_n35540_, new_n35541_, new_n35542_, new_n35543_, new_n35544_,
    new_n35545_, new_n35546_, new_n35547_, new_n35548_, new_n35549_,
    new_n35550_, new_n35551_, new_n35552_, new_n35553_, new_n35554_,
    new_n35555_, new_n35556_, new_n35557_, new_n35558_, new_n35559_,
    new_n35560_, new_n35561_, new_n35562_, new_n35563_, new_n35564_,
    new_n35565_, new_n35566_, new_n35567_, new_n35568_, new_n35569_,
    new_n35570_, new_n35571_, new_n35572_, new_n35573_, new_n35574_,
    new_n35575_, new_n35576_, new_n35577_, new_n35578_, new_n35579_,
    new_n35580_, new_n35581_, new_n35582_, new_n35583_, new_n35584_,
    new_n35585_, new_n35586_, new_n35587_, new_n35588_, new_n35589_,
    new_n35590_, new_n35591_, new_n35592_, new_n35593_, new_n35594_,
    new_n35595_, new_n35596_, new_n35597_, new_n35598_, new_n35599_,
    new_n35600_, new_n35601_, new_n35602_, new_n35603_, new_n35604_,
    new_n35605_, new_n35606_, new_n35607_, new_n35608_, new_n35609_,
    new_n35610_, new_n35611_, new_n35612_, new_n35613_, new_n35614_,
    new_n35615_, new_n35616_, new_n35617_, new_n35618_, new_n35619_,
    new_n35620_, new_n35621_, new_n35622_, new_n35623_, new_n35624_,
    new_n35625_, new_n35626_, new_n35627_, new_n35628_, new_n35629_,
    new_n35630_, new_n35631_, new_n35632_, new_n35633_, new_n35634_,
    new_n35635_, new_n35636_, new_n35637_, new_n35638_, new_n35639_,
    new_n35640_, new_n35641_, new_n35642_, new_n35643_, new_n35645_,
    new_n35646_, new_n35647_, new_n35648_, new_n35649_, new_n35650_,
    new_n35651_, new_n35652_, new_n35653_, new_n35654_, new_n35655_,
    new_n35656_, new_n35657_, new_n35658_, new_n35659_, new_n35660_,
    new_n35661_, new_n35662_, new_n35663_, new_n35664_, new_n35665_,
    new_n35666_, new_n35667_, new_n35668_, new_n35669_, new_n35670_,
    new_n35671_, new_n35672_, new_n35673_, new_n35674_, new_n35675_,
    new_n35676_, new_n35677_, new_n35678_, new_n35679_, new_n35680_,
    new_n35681_, new_n35682_, new_n35683_, new_n35684_, new_n35685_,
    new_n35686_, new_n35687_, new_n35688_, new_n35689_, new_n35690_,
    new_n35691_, new_n35692_, new_n35693_, new_n35694_, new_n35695_,
    new_n35696_, new_n35697_, new_n35698_, new_n35699_, new_n35700_,
    new_n35701_, new_n35702_, new_n35703_, new_n35704_, new_n35705_,
    new_n35706_, new_n35707_, new_n35708_, new_n35709_, new_n35710_,
    new_n35711_, new_n35712_, new_n35713_, new_n35714_, new_n35715_,
    new_n35716_, new_n35717_, new_n35718_, new_n35719_, new_n35720_,
    new_n35721_, new_n35722_, new_n35723_, new_n35724_, new_n35725_,
    new_n35726_, new_n35727_, new_n35728_, new_n35729_, new_n35730_,
    new_n35731_, new_n35732_, new_n35733_, new_n35734_, new_n35735_,
    new_n35736_, new_n35737_, new_n35738_, new_n35739_, new_n35740_,
    new_n35741_, new_n35742_, new_n35743_, new_n35744_, new_n35745_,
    new_n35746_, new_n35747_, new_n35748_, new_n35749_, new_n35750_,
    new_n35751_, new_n35752_, new_n35753_, new_n35754_, new_n35755_,
    new_n35756_, new_n35757_, new_n35758_, new_n35759_, new_n35760_,
    new_n35761_, new_n35762_, new_n35763_, new_n35764_, new_n35765_,
    new_n35766_, new_n35767_, new_n35768_, new_n35769_, new_n35771_,
    new_n35772_, new_n35773_, new_n35774_, new_n35775_, new_n35776_,
    new_n35777_, new_n35778_, new_n35779_, new_n35780_, new_n35781_,
    new_n35782_, new_n35783_, new_n35784_, new_n35785_, new_n35786_,
    new_n35787_, new_n35788_, new_n35789_, new_n35790_, new_n35791_,
    new_n35792_, new_n35793_, new_n35794_, new_n35795_, new_n35796_,
    new_n35798_, new_n35799_, new_n35800_, new_n35801_, new_n35802_,
    new_n35803_, new_n35804_, new_n35805_, new_n35806_, new_n35807_,
    new_n35808_, new_n35809_, new_n35810_, new_n35811_, new_n35812_,
    new_n35813_, new_n35814_, new_n35815_, new_n35816_, new_n35817_,
    new_n35819_, new_n35820_, new_n35821_, new_n35822_, new_n35823_,
    new_n35824_, new_n35825_, new_n35826_, new_n35827_, new_n35828_,
    new_n35829_, new_n35830_, new_n35831_, new_n35832_, new_n35833_,
    new_n35834_, new_n35835_, new_n35836_, new_n35837_, new_n35838_,
    new_n35840_, new_n35841_, new_n35842_, new_n35843_, new_n35844_,
    new_n35845_, new_n35846_, new_n35847_, new_n35848_, new_n35849_,
    new_n35850_, new_n35851_, new_n35852_, new_n35853_, new_n35854_,
    new_n35855_, new_n35856_, new_n35857_, new_n35858_, new_n35859_,
    new_n35861_, new_n35862_, new_n35863_, new_n35864_, new_n35865_,
    new_n35866_, new_n35867_, new_n35868_, new_n35869_, new_n35870_,
    new_n35871_, new_n35872_, new_n35873_, new_n35874_, new_n35875_,
    new_n35876_, new_n35877_, new_n35878_, new_n35879_, new_n35880_,
    new_n35881_, new_n35882_, new_n35883_, new_n35884_, new_n35885_,
    new_n35886_, new_n35887_, new_n35888_, new_n35889_, new_n35890_,
    new_n35891_, new_n35892_, new_n35893_, new_n35894_, new_n35895_,
    new_n35896_, new_n35897_, new_n35898_, new_n35899_, new_n35900_,
    new_n35901_, new_n35902_, new_n35903_, new_n35904_, new_n35905_,
    new_n35906_, new_n35907_, new_n35908_, new_n35909_, new_n35910_,
    new_n35911_, new_n35912_, new_n35913_, new_n35914_, new_n35915_,
    new_n35916_, new_n35917_, new_n35918_, new_n35919_, new_n35920_,
    new_n35921_, new_n35922_, new_n35923_, new_n35924_, new_n35925_,
    new_n35926_, new_n35927_, new_n35928_, new_n35929_, new_n35930_,
    new_n35931_, new_n35932_, new_n35933_, new_n35934_, new_n35935_,
    new_n35936_, new_n35937_, new_n35938_, new_n35939_, new_n35940_,
    new_n35941_, new_n35942_, new_n35943_, new_n35944_, new_n35945_,
    new_n35946_, new_n35947_, new_n35948_, new_n35949_, new_n35950_,
    new_n35951_, new_n35952_, new_n35953_, new_n35954_, new_n35955_,
    new_n35956_, new_n35957_, new_n35958_, new_n35959_, new_n35960_,
    new_n35961_, new_n35962_, new_n35963_, new_n35964_, new_n35965_,
    new_n35966_, new_n35967_, new_n35968_, new_n35969_, new_n35970_,
    new_n35971_, new_n35972_, new_n35973_, new_n35974_, new_n35975_,
    new_n35977_, new_n35978_, new_n35979_, new_n35980_, new_n35981_,
    new_n35982_, new_n35983_, new_n35984_, new_n35985_, new_n35986_,
    new_n35987_, new_n35988_, new_n35989_, new_n35990_, new_n35991_,
    new_n35992_, new_n35993_, new_n35994_, new_n35995_, new_n35996_,
    new_n35997_, new_n35998_, new_n35999_, new_n36000_, new_n36001_,
    new_n36002_, new_n36003_, new_n36004_, new_n36005_, new_n36006_,
    new_n36007_, new_n36008_, new_n36009_, new_n36010_, new_n36011_,
    new_n36012_, new_n36013_, new_n36014_, new_n36015_, new_n36016_,
    new_n36017_, new_n36018_, new_n36019_, new_n36020_, new_n36021_,
    new_n36022_, new_n36023_, new_n36024_, new_n36025_, new_n36026_,
    new_n36027_, new_n36028_, new_n36029_, new_n36030_, new_n36031_,
    new_n36032_, new_n36033_, new_n36034_, new_n36035_, new_n36036_,
    new_n36037_, new_n36038_, new_n36039_, new_n36040_, new_n36041_,
    new_n36042_, new_n36043_, new_n36044_, new_n36045_, new_n36046_,
    new_n36047_, new_n36048_, new_n36049_, new_n36050_, new_n36051_,
    new_n36052_, new_n36053_, new_n36054_, new_n36055_, new_n36056_,
    new_n36057_, new_n36058_, new_n36059_, new_n36060_, new_n36061_,
    new_n36062_, new_n36063_, new_n36064_, new_n36065_, new_n36066_,
    new_n36067_, new_n36068_, new_n36069_, new_n36070_, new_n36071_,
    new_n36072_, new_n36073_, new_n36074_, new_n36075_, new_n36076_,
    new_n36077_, new_n36078_, new_n36079_, new_n36080_, new_n36081_,
    new_n36082_, new_n36083_, new_n36084_, new_n36085_, new_n36086_,
    new_n36088_, new_n36089_, new_n36090_, new_n36091_, new_n36092_,
    new_n36093_, new_n36094_, new_n36095_, new_n36096_, new_n36097_,
    new_n36098_, new_n36099_, new_n36100_, new_n36101_, new_n36102_,
    new_n36103_, new_n36104_, new_n36105_, new_n36107_, new_n36108_,
    new_n36109_, new_n36110_, new_n36111_, new_n36112_, new_n36114_,
    new_n36115_, new_n36116_, new_n36117_, new_n36118_, new_n36119_,
    new_n36120_, new_n36121_, new_n36122_, new_n36123_, new_n36124_,
    new_n36125_, new_n36126_, new_n36127_, new_n36128_, new_n36129_,
    new_n36130_, new_n36131_, new_n36132_, new_n36133_, new_n36135_,
    new_n36136_, new_n36137_, new_n36138_, new_n36139_, new_n36140_,
    new_n36142_, new_n36143_, new_n36144_, new_n36145_, new_n36146_,
    new_n36147_, new_n36148_, new_n36149_, new_n36150_, new_n36151_,
    new_n36152_, new_n36153_, new_n36154_, new_n36155_, new_n36156_,
    new_n36157_, new_n36158_, new_n36159_, new_n36160_, new_n36161_,
    new_n36162_, new_n36163_, new_n36164_, new_n36165_, new_n36166_,
    new_n36167_, new_n36168_, new_n36169_, new_n36170_, new_n36171_,
    new_n36172_, new_n36173_, new_n36174_, new_n36175_, new_n36176_,
    new_n36177_, new_n36178_, new_n36179_, new_n36180_, new_n36181_,
    new_n36182_, new_n36183_, new_n36184_, new_n36185_, new_n36186_,
    new_n36187_, new_n36188_, new_n36189_, new_n36190_, new_n36191_,
    new_n36192_, new_n36193_, new_n36194_, new_n36195_, new_n36196_,
    new_n36197_, new_n36198_, new_n36199_, new_n36200_, new_n36201_,
    new_n36202_, new_n36203_, new_n36204_, new_n36205_, new_n36206_,
    new_n36207_, new_n36208_, new_n36209_, new_n36210_, new_n36211_,
    new_n36212_, new_n36213_, new_n36214_, new_n36215_, new_n36216_,
    new_n36217_, new_n36218_, new_n36219_, new_n36220_, new_n36221_,
    new_n36222_, new_n36223_, new_n36224_, new_n36225_, new_n36226_,
    new_n36227_, new_n36228_, new_n36229_, new_n36230_, new_n36231_,
    new_n36232_, new_n36233_, new_n36234_, new_n36235_, new_n36236_,
    new_n36237_, new_n36238_, new_n36239_, new_n36240_, new_n36241_,
    new_n36242_, new_n36243_, new_n36244_, new_n36245_, new_n36246_,
    new_n36247_, new_n36248_, new_n36249_, new_n36251_, new_n36252_,
    new_n36253_, new_n36254_, new_n36255_, new_n36256_, new_n36257_,
    new_n36258_, new_n36259_, new_n36260_, new_n36261_, new_n36262_,
    new_n36263_, new_n36264_, new_n36265_, new_n36266_, new_n36267_,
    new_n36268_, new_n36269_, new_n36270_, new_n36271_, new_n36272_,
    new_n36273_, new_n36274_, new_n36275_, new_n36276_, new_n36277_,
    new_n36278_, new_n36279_, new_n36280_, new_n36281_, new_n36282_,
    new_n36283_, new_n36284_, new_n36285_, new_n36286_, new_n36287_,
    new_n36288_, new_n36289_, new_n36290_, new_n36291_, new_n36292_,
    new_n36293_, new_n36294_, new_n36295_, new_n36296_, new_n36297_,
    new_n36298_, new_n36299_, new_n36300_, new_n36301_, new_n36302_,
    new_n36303_, new_n36304_, new_n36305_, new_n36306_, new_n36307_,
    new_n36308_, new_n36309_, new_n36310_, new_n36311_, new_n36312_,
    new_n36313_, new_n36314_, new_n36315_, new_n36316_, new_n36317_,
    new_n36318_, new_n36319_, new_n36320_, new_n36321_, new_n36322_,
    new_n36323_, new_n36324_, new_n36325_, new_n36326_, new_n36327_,
    new_n36328_, new_n36329_, new_n36330_, new_n36331_, new_n36332_,
    new_n36333_, new_n36334_, new_n36335_, new_n36336_, new_n36337_,
    new_n36338_, new_n36339_, new_n36340_, new_n36341_, new_n36342_,
    new_n36343_, new_n36344_, new_n36345_, new_n36346_, new_n36347_,
    new_n36348_, new_n36349_, new_n36350_, new_n36351_, new_n36352_,
    new_n36353_, new_n36354_, new_n36355_, new_n36356_, new_n36357_,
    new_n36358_, new_n36359_, new_n36360_, new_n36361_, new_n36362_,
    new_n36363_, new_n36364_, new_n36365_, new_n36366_, new_n36367_,
    new_n36368_, new_n36369_, new_n36370_, new_n36371_, new_n36372_,
    new_n36373_, new_n36374_, new_n36375_, new_n36376_, new_n36377_,
    new_n36378_, new_n36379_, new_n36380_, new_n36381_, new_n36382_,
    new_n36383_, new_n36384_, new_n36385_, new_n36386_, new_n36387_,
    new_n36388_, new_n36389_, new_n36390_, new_n36391_, new_n36392_,
    new_n36393_, new_n36394_, new_n36395_, new_n36396_, new_n36397_,
    new_n36398_, new_n36399_, new_n36400_, new_n36401_, new_n36402_,
    new_n36403_, new_n36404_, new_n36405_, new_n36406_, new_n36407_,
    new_n36408_, new_n36409_, new_n36410_, new_n36411_, new_n36412_,
    new_n36413_, new_n36414_, new_n36415_, new_n36416_, new_n36417_,
    new_n36418_, new_n36419_, new_n36420_, new_n36421_, new_n36422_,
    new_n36423_, new_n36424_, new_n36425_, new_n36426_, new_n36427_,
    new_n36428_, new_n36429_, new_n36430_, new_n36431_, new_n36432_,
    new_n36433_, new_n36434_, new_n36435_, new_n36436_, new_n36437_,
    new_n36438_, new_n36439_, new_n36440_, new_n36441_, new_n36442_,
    new_n36443_, new_n36444_, new_n36445_, new_n36446_, new_n36447_,
    new_n36448_, new_n36449_, new_n36450_, new_n36451_, new_n36452_,
    new_n36453_, new_n36454_, new_n36455_, new_n36456_, new_n36457_,
    new_n36458_, new_n36459_, new_n36460_, new_n36461_, new_n36462_,
    new_n36463_, new_n36464_, new_n36465_, new_n36466_, new_n36467_,
    new_n36468_, new_n36469_, new_n36470_, new_n36471_, new_n36472_,
    new_n36473_, new_n36474_, new_n36475_, new_n36476_, new_n36477_,
    new_n36478_, new_n36479_, new_n36480_, new_n36481_, new_n36482_,
    new_n36483_, new_n36484_, new_n36485_, new_n36486_, new_n36487_,
    new_n36488_, new_n36489_, new_n36490_, new_n36491_, new_n36492_,
    new_n36493_, new_n36494_, new_n36495_, new_n36496_, new_n36497_,
    new_n36498_, new_n36499_, new_n36500_, new_n36501_, new_n36502_,
    new_n36503_, new_n36504_, new_n36505_, new_n36506_, new_n36507_,
    new_n36508_, new_n36509_, new_n36510_, new_n36511_, new_n36512_,
    new_n36513_, new_n36514_, new_n36515_, new_n36516_, new_n36517_,
    new_n36518_, new_n36519_, new_n36520_, new_n36521_, new_n36522_,
    new_n36523_, new_n36524_, new_n36525_, new_n36526_, new_n36527_,
    new_n36528_, new_n36529_, new_n36530_, new_n36531_, new_n36532_,
    new_n36533_, new_n36534_, new_n36535_, new_n36536_, new_n36537_,
    new_n36538_, new_n36539_, new_n36540_, new_n36541_, new_n36542_,
    new_n36543_, new_n36544_, new_n36545_, new_n36546_, new_n36547_,
    new_n36548_, new_n36549_, new_n36550_, new_n36551_, new_n36552_,
    new_n36553_, new_n36554_, new_n36555_, new_n36556_, new_n36557_,
    new_n36558_, new_n36559_, new_n36560_, new_n36561_, new_n36562_,
    new_n36563_, new_n36564_, new_n36565_, new_n36566_, new_n36567_,
    new_n36568_, new_n36569_, new_n36570_, new_n36571_, new_n36572_,
    new_n36573_, new_n36574_, new_n36575_, new_n36576_, new_n36577_,
    new_n36578_, new_n36579_, new_n36580_, new_n36581_, new_n36582_,
    new_n36583_, new_n36584_, new_n36585_, new_n36586_, new_n36587_,
    new_n36588_, new_n36589_, new_n36590_, new_n36591_, new_n36592_,
    new_n36593_, new_n36594_, new_n36595_, new_n36596_, new_n36597_,
    new_n36598_, new_n36599_, new_n36600_, new_n36601_, new_n36602_,
    new_n36603_, new_n36604_, new_n36605_, new_n36606_, new_n36607_,
    new_n36608_, new_n36609_, new_n36610_, new_n36611_, new_n36612_,
    new_n36613_, new_n36614_, new_n36615_, new_n36616_, new_n36617_,
    new_n36618_, new_n36619_, new_n36620_, new_n36621_, new_n36622_,
    new_n36623_, new_n36624_, new_n36625_, new_n36626_, new_n36627_,
    new_n36628_, new_n36629_, new_n36630_, new_n36631_, new_n36632_,
    new_n36633_, new_n36634_, new_n36635_, new_n36636_, new_n36637_,
    new_n36638_, new_n36639_, new_n36640_, new_n36641_, new_n36642_,
    new_n36643_, new_n36644_, new_n36645_, new_n36646_, new_n36647_,
    new_n36648_, new_n36649_, new_n36650_, new_n36651_, new_n36652_,
    new_n36653_, new_n36654_, new_n36655_, new_n36656_, new_n36657_,
    new_n36658_, new_n36659_, new_n36660_, new_n36661_, new_n36662_,
    new_n36663_, new_n36664_, new_n36665_, new_n36666_, new_n36667_,
    new_n36668_, new_n36669_, new_n36670_, new_n36671_, new_n36672_,
    new_n36673_, new_n36674_, new_n36675_, new_n36676_, new_n36677_,
    new_n36678_, new_n36679_, new_n36680_, new_n36681_, new_n36682_,
    new_n36683_, new_n36684_, new_n36685_, new_n36686_, new_n36687_,
    new_n36688_, new_n36689_, new_n36690_, new_n36691_, new_n36692_,
    new_n36693_, new_n36694_, new_n36695_, new_n36696_, new_n36697_,
    new_n36698_, new_n36699_, new_n36700_, new_n36701_, new_n36702_,
    new_n36703_, new_n36704_, new_n36705_, new_n36706_, new_n36707_,
    new_n36708_, new_n36709_, new_n36710_, new_n36711_, new_n36712_,
    new_n36713_, new_n36714_, new_n36715_, new_n36716_, new_n36717_,
    new_n36718_, new_n36719_, new_n36720_, new_n36721_, new_n36722_,
    new_n36723_, new_n36724_, new_n36725_, new_n36726_, new_n36727_,
    new_n36728_, new_n36729_, new_n36730_, new_n36731_, new_n36732_,
    new_n36733_, new_n36734_, new_n36735_, new_n36736_, new_n36737_,
    new_n36738_, new_n36739_, new_n36740_, new_n36741_, new_n36742_,
    new_n36743_, new_n36744_, new_n36745_, new_n36746_, new_n36747_,
    new_n36748_, new_n36749_, new_n36750_, new_n36751_, new_n36752_,
    new_n36753_, new_n36754_, new_n36755_, new_n36756_, new_n36757_,
    new_n36758_, new_n36759_, new_n36760_, new_n36761_, new_n36762_,
    new_n36763_, new_n36764_, new_n36765_, new_n36766_, new_n36767_,
    new_n36768_, new_n36769_, new_n36770_, new_n36771_, new_n36772_,
    new_n36773_, new_n36774_, new_n36775_, new_n36776_, new_n36777_,
    new_n36778_, new_n36779_, new_n36780_, new_n36781_, new_n36782_,
    new_n36783_, new_n36784_, new_n36785_, new_n36786_, new_n36787_,
    new_n36788_, new_n36789_, new_n36790_, new_n36791_, new_n36792_,
    new_n36793_, new_n36794_, new_n36795_, new_n36796_, new_n36797_,
    new_n36798_, new_n36799_, new_n36800_, new_n36801_, new_n36802_,
    new_n36803_, new_n36804_, new_n36805_, new_n36806_, new_n36807_,
    new_n36808_, new_n36809_, new_n36810_, new_n36811_, new_n36812_,
    new_n36813_, new_n36814_, new_n36815_, new_n36816_, new_n36817_,
    new_n36818_, new_n36819_, new_n36820_, new_n36821_, new_n36822_,
    new_n36823_, new_n36824_, new_n36825_, new_n36826_, new_n36827_,
    new_n36828_, new_n36829_, new_n36830_, new_n36831_, new_n36832_,
    new_n36833_, new_n36834_, new_n36835_, new_n36836_, new_n36837_,
    new_n36838_, new_n36839_, new_n36840_, new_n36841_, new_n36842_,
    new_n36843_, new_n36844_, new_n36845_, new_n36846_, new_n36847_,
    new_n36848_, new_n36849_, new_n36850_, new_n36851_, new_n36852_,
    new_n36853_, new_n36854_, new_n36855_, new_n36856_, new_n36857_,
    new_n36858_, new_n36859_, new_n36860_, new_n36861_, new_n36862_,
    new_n36863_, new_n36864_, new_n36865_, new_n36866_, new_n36867_,
    new_n36868_, new_n36869_, new_n36870_, new_n36871_, new_n36872_,
    new_n36873_, new_n36874_, new_n36875_, new_n36877_, new_n36878_,
    new_n36879_, new_n36880_, new_n36881_, new_n36882_, new_n36883_,
    new_n36884_, new_n36885_, new_n36886_, new_n36887_, new_n36888_,
    new_n36889_, new_n36890_, new_n36891_, new_n36892_, new_n36893_,
    new_n36894_, new_n36895_, new_n36896_, new_n36897_, new_n36898_,
    new_n36899_, new_n36900_, new_n36901_, new_n36902_, new_n36903_,
    new_n36904_, new_n36905_, new_n36906_, new_n36907_, new_n36908_,
    new_n36909_, new_n36910_, new_n36911_, new_n36912_, new_n36913_,
    new_n36914_, new_n36915_, new_n36916_, new_n36917_, new_n36918_,
    new_n36919_, new_n36920_, new_n36921_, new_n36922_, new_n36923_,
    new_n36924_, new_n36925_, new_n36926_, new_n36927_, new_n36928_,
    new_n36929_, new_n36930_, new_n36931_, new_n36932_, new_n36933_,
    new_n36934_, new_n36935_, new_n36936_, new_n36937_, new_n36938_,
    new_n36939_, new_n36940_, new_n36941_, new_n36942_, new_n36943_,
    new_n36944_, new_n36945_, new_n36946_, new_n36947_, new_n36948_,
    new_n36949_, new_n36950_, new_n36951_, new_n36952_, new_n36953_,
    new_n36954_, new_n36955_, new_n36956_, new_n36957_, new_n36958_,
    new_n36959_, new_n36960_, new_n36961_, new_n36962_, new_n36963_,
    new_n36964_, new_n36965_, new_n36966_, new_n36967_, new_n36968_,
    new_n36969_, new_n36970_, new_n36971_, new_n36972_, new_n36973_,
    new_n36974_, new_n36975_, new_n36976_, new_n36977_, new_n36978_,
    new_n36979_, new_n36980_, new_n36981_, new_n36982_, new_n36983_,
    new_n36984_, new_n36985_, new_n36986_, new_n36987_, new_n36988_,
    new_n36989_, new_n36990_, new_n36991_, new_n36992_, new_n36993_,
    new_n36994_, new_n36995_, new_n36996_, new_n36997_, new_n36998_,
    new_n36999_, new_n37000_, new_n37001_, new_n37002_, new_n37003_,
    new_n37004_, new_n37005_, new_n37006_, new_n37007_, new_n37008_,
    new_n37009_, new_n37010_, new_n37011_, new_n37012_, new_n37013_,
    new_n37014_, new_n37015_, new_n37016_, new_n37017_, new_n37018_,
    new_n37019_, new_n37020_, new_n37021_, new_n37022_, new_n37023_,
    new_n37024_, new_n37025_, new_n37026_, new_n37027_, new_n37028_,
    new_n37029_, new_n37030_, new_n37031_, new_n37032_, new_n37033_,
    new_n37034_, new_n37035_, new_n37036_, new_n37037_, new_n37038_,
    new_n37039_, new_n37040_, new_n37041_, new_n37042_, new_n37043_,
    new_n37044_, new_n37045_, new_n37046_, new_n37047_, new_n37048_,
    new_n37049_, new_n37050_, new_n37051_, new_n37052_, new_n37053_,
    new_n37054_, new_n37055_, new_n37056_, new_n37057_, new_n37058_,
    new_n37059_, new_n37060_, new_n37061_, new_n37062_, new_n37063_,
    new_n37064_, new_n37065_, new_n37066_, new_n37067_, new_n37068_,
    new_n37069_, new_n37070_, new_n37071_, new_n37072_, new_n37073_,
    new_n37074_, new_n37075_, new_n37076_, new_n37077_, new_n37078_,
    new_n37079_, new_n37080_, new_n37081_, new_n37082_, new_n37083_,
    new_n37084_, new_n37085_, new_n37086_, new_n37087_, new_n37088_,
    new_n37089_, new_n37090_, new_n37091_, new_n37092_, new_n37093_,
    new_n37094_, new_n37095_, new_n37096_, new_n37097_, new_n37098_,
    new_n37099_, new_n37100_, new_n37101_, new_n37102_, new_n37103_,
    new_n37104_, new_n37105_, new_n37106_, new_n37107_, new_n37108_,
    new_n37109_, new_n37110_, new_n37111_, new_n37112_, new_n37113_,
    new_n37114_, new_n37115_, new_n37116_, new_n37117_, new_n37118_,
    new_n37119_, new_n37120_, new_n37121_, new_n37122_, new_n37123_,
    new_n37124_, new_n37125_, new_n37126_, new_n37127_, new_n37128_,
    new_n37129_, new_n37130_, new_n37131_, new_n37132_, new_n37133_,
    new_n37134_, new_n37135_, new_n37136_, new_n37137_, new_n37138_,
    new_n37139_, new_n37140_, new_n37141_, new_n37142_, new_n37143_,
    new_n37144_, new_n37145_, new_n37146_, new_n37147_, new_n37148_,
    new_n37149_, new_n37150_, new_n37151_, new_n37152_, new_n37153_,
    new_n37154_, new_n37155_, new_n37156_, new_n37157_, new_n37158_,
    new_n37159_, new_n37160_, new_n37161_, new_n37162_, new_n37163_,
    new_n37164_, new_n37165_, new_n37166_, new_n37167_, new_n37168_,
    new_n37169_, new_n37170_, new_n37171_, new_n37172_, new_n37173_,
    new_n37174_, new_n37175_, new_n37176_, new_n37177_, new_n37178_,
    new_n37179_, new_n37180_, new_n37181_, new_n37182_, new_n37183_,
    new_n37184_, new_n37185_, new_n37186_, new_n37187_, new_n37188_,
    new_n37189_, new_n37190_, new_n37191_, new_n37192_, new_n37193_,
    new_n37194_, new_n37195_, new_n37196_, new_n37197_, new_n37198_,
    new_n37199_, new_n37200_, new_n37201_, new_n37202_, new_n37203_,
    new_n37204_, new_n37205_, new_n37206_, new_n37207_, new_n37208_,
    new_n37209_, new_n37210_, new_n37211_, new_n37212_, new_n37213_,
    new_n37214_, new_n37215_, new_n37216_, new_n37217_, new_n37218_,
    new_n37219_, new_n37220_, new_n37221_, new_n37222_, new_n37223_,
    new_n37224_, new_n37225_, new_n37226_, new_n37227_, new_n37228_,
    new_n37229_, new_n37230_, new_n37231_, new_n37232_, new_n37233_,
    new_n37234_, new_n37235_, new_n37236_, new_n37237_, new_n37238_,
    new_n37239_, new_n37240_, new_n37241_, new_n37242_, new_n37243_,
    new_n37244_, new_n37245_, new_n37246_, new_n37247_, new_n37248_,
    new_n37249_, new_n37250_, new_n37251_, new_n37252_, new_n37253_,
    new_n37254_, new_n37255_, new_n37256_, new_n37257_, new_n37258_,
    new_n37259_, new_n37260_, new_n37261_, new_n37262_, new_n37263_,
    new_n37264_, new_n37265_, new_n37266_, new_n37267_, new_n37268_,
    new_n37269_, new_n37270_, new_n37271_, new_n37272_, new_n37273_,
    new_n37274_, new_n37275_, new_n37276_, new_n37277_, new_n37278_,
    new_n37279_, new_n37280_, new_n37281_, new_n37282_, new_n37283_,
    new_n37284_, new_n37285_, new_n37286_, new_n37287_, new_n37288_,
    new_n37289_, new_n37290_, new_n37291_, new_n37292_, new_n37293_,
    new_n37294_, new_n37295_, new_n37296_, new_n37297_, new_n37298_,
    new_n37299_, new_n37300_, new_n37301_, new_n37302_, new_n37303_,
    new_n37304_, new_n37305_, new_n37306_, new_n37307_, new_n37308_,
    new_n37309_, new_n37310_, new_n37311_, new_n37312_, new_n37313_,
    new_n37314_, new_n37315_, new_n37316_, new_n37317_, new_n37318_,
    new_n37319_, new_n37320_, new_n37321_, new_n37322_, new_n37323_,
    new_n37324_, new_n37325_, new_n37326_, new_n37327_, new_n37328_,
    new_n37329_, new_n37330_, new_n37331_, new_n37332_, new_n37333_,
    new_n37334_, new_n37335_, new_n37336_, new_n37337_, new_n37338_,
    new_n37339_, new_n37340_, new_n37341_, new_n37342_, new_n37343_,
    new_n37344_, new_n37345_, new_n37346_, new_n37347_, new_n37348_,
    new_n37349_, new_n37350_, new_n37351_, new_n37352_, new_n37353_,
    new_n37354_, new_n37355_, new_n37356_, new_n37357_, new_n37358_,
    new_n37359_, new_n37360_, new_n37361_, new_n37362_, new_n37363_,
    new_n37364_, new_n37365_, new_n37366_, new_n37367_, new_n37368_,
    new_n37369_, new_n37370_, new_n37371_, new_n37372_, new_n37373_,
    new_n37374_, new_n37375_, new_n37376_, new_n37377_, new_n37378_,
    new_n37379_, new_n37380_, new_n37381_, new_n37382_, new_n37383_,
    new_n37384_, new_n37385_, new_n37386_, new_n37387_, new_n37388_,
    new_n37389_, new_n37390_, new_n37391_, new_n37392_, new_n37393_,
    new_n37394_, new_n37395_, new_n37396_, new_n37397_, new_n37398_,
    new_n37399_, new_n37400_, new_n37401_, new_n37402_, new_n37403_,
    new_n37404_, new_n37405_, new_n37406_, new_n37407_, new_n37408_,
    new_n37409_, new_n37410_, new_n37411_, new_n37412_, new_n37413_,
    new_n37414_, new_n37415_, new_n37416_, new_n37417_, new_n37418_,
    new_n37419_, new_n37420_, new_n37421_, new_n37422_, new_n37423_,
    new_n37424_, new_n37425_, new_n37426_, new_n37427_, new_n37428_,
    new_n37429_, new_n37430_, new_n37431_, new_n37432_, new_n37433_,
    new_n37434_, new_n37435_, new_n37436_, new_n37437_, new_n37438_,
    new_n37439_, new_n37440_, new_n37441_, new_n37442_, new_n37443_,
    new_n37444_, new_n37445_, new_n37446_, new_n37447_, new_n37448_,
    new_n37449_, new_n37450_, new_n37451_, new_n37452_, new_n37453_,
    new_n37454_, new_n37455_, new_n37456_, new_n37457_, new_n37459_,
    new_n37460_, new_n37461_, new_n37462_, new_n37463_, new_n37464_,
    new_n37465_, new_n37466_, new_n37467_, new_n37468_, new_n37469_,
    new_n37470_, new_n37471_, new_n37472_, new_n37473_, new_n37474_,
    new_n37475_, new_n37476_, new_n37477_, new_n37478_, new_n37479_,
    new_n37480_, new_n37481_, new_n37482_, new_n37483_, new_n37484_,
    new_n37485_, new_n37486_, new_n37487_, new_n37488_, new_n37489_,
    new_n37490_, new_n37491_, new_n37492_, new_n37493_, new_n37494_,
    new_n37495_, new_n37496_, new_n37497_, new_n37498_, new_n37499_,
    new_n37500_, new_n37501_, new_n37502_, new_n37503_, new_n37504_,
    new_n37505_, new_n37506_, new_n37507_, new_n37508_, new_n37509_,
    new_n37510_, new_n37511_, new_n37512_, new_n37513_, new_n37514_,
    new_n37515_, new_n37516_, new_n37517_, new_n37518_, new_n37519_,
    new_n37520_, new_n37521_, new_n37522_, new_n37523_, new_n37524_,
    new_n37525_, new_n37526_, new_n37527_, new_n37528_, new_n37529_,
    new_n37530_, new_n37531_, new_n37532_, new_n37533_, new_n37534_,
    new_n37535_, new_n37536_, new_n37537_, new_n37538_, new_n37539_,
    new_n37540_, new_n37541_, new_n37542_, new_n37543_, new_n37544_,
    new_n37545_, new_n37546_, new_n37547_, new_n37548_, new_n37549_,
    new_n37550_, new_n37551_, new_n37552_, new_n37553_, new_n37554_,
    new_n37555_, new_n37556_, new_n37557_, new_n37558_, new_n37559_,
    new_n37560_, new_n37561_, new_n37562_, new_n37563_, new_n37564_,
    new_n37565_, new_n37566_, new_n37567_, new_n37568_, new_n37569_,
    new_n37570_, new_n37571_, new_n37572_, new_n37573_, new_n37574_,
    new_n37575_, new_n37576_, new_n37577_, new_n37578_, new_n37579_,
    new_n37580_, new_n37581_, new_n37582_, new_n37583_, new_n37584_,
    new_n37585_, new_n37586_, new_n37587_, new_n37588_, new_n37589_,
    new_n37590_, new_n37591_, new_n37592_, new_n37593_, new_n37594_,
    new_n37595_, new_n37596_, new_n37597_, new_n37598_, new_n37599_,
    new_n37600_, new_n37601_, new_n37602_, new_n37603_, new_n37604_,
    new_n37605_, new_n37606_, new_n37607_, new_n37608_, new_n37609_,
    new_n37610_, new_n37611_, new_n37612_, new_n37613_, new_n37614_,
    new_n37615_, new_n37616_, new_n37617_, new_n37618_, new_n37619_,
    new_n37620_, new_n37621_, new_n37622_, new_n37623_, new_n37624_,
    new_n37625_, new_n37626_, new_n37627_, new_n37628_, new_n37629_,
    new_n37630_, new_n37631_, new_n37632_, new_n37633_, new_n37634_,
    new_n37635_, new_n37636_, new_n37637_, new_n37638_, new_n37639_,
    new_n37640_, new_n37641_, new_n37642_, new_n37643_, new_n37644_,
    new_n37645_, new_n37646_, new_n37647_, new_n37648_, new_n37649_,
    new_n37650_, new_n37651_, new_n37652_, new_n37653_, new_n37654_,
    new_n37655_, new_n37656_, new_n37657_, new_n37658_, new_n37659_,
    new_n37660_, new_n37661_, new_n37662_, new_n37663_, new_n37664_,
    new_n37665_, new_n37666_, new_n37667_, new_n37668_, new_n37669_,
    new_n37670_, new_n37671_, new_n37672_, new_n37673_, new_n37674_,
    new_n37675_, new_n37676_, new_n37677_, new_n37678_, new_n37679_,
    new_n37680_, new_n37681_, new_n37682_, new_n37683_, new_n37684_,
    new_n37685_, new_n37686_, new_n37687_, new_n37688_, new_n37689_,
    new_n37690_, new_n37691_, new_n37692_, new_n37693_, new_n37694_,
    new_n37695_, new_n37696_, new_n37697_, new_n37698_, new_n37699_,
    new_n37700_, new_n37701_, new_n37702_, new_n37703_, new_n37704_,
    new_n37705_, new_n37706_, new_n37707_, new_n37708_, new_n37709_,
    new_n37710_, new_n37711_, new_n37712_, new_n37713_, new_n37714_,
    new_n37715_, new_n37716_, new_n37717_, new_n37718_, new_n37719_,
    new_n37720_, new_n37721_, new_n37722_, new_n37723_, new_n37724_,
    new_n37725_, new_n37726_, new_n37727_, new_n37728_, new_n37729_,
    new_n37730_, new_n37731_, new_n37732_, new_n37733_, new_n37734_,
    new_n37735_, new_n37736_, new_n37737_, new_n37738_, new_n37739_,
    new_n37740_, new_n37741_, new_n37742_, new_n37743_, new_n37744_,
    new_n37745_, new_n37746_, new_n37747_, new_n37748_, new_n37749_,
    new_n37750_, new_n37751_, new_n37752_, new_n37753_, new_n37754_,
    new_n37755_, new_n37756_, new_n37757_, new_n37758_, new_n37759_,
    new_n37760_, new_n37761_, new_n37762_, new_n37763_, new_n37764_,
    new_n37765_, new_n37766_, new_n37767_, new_n37768_, new_n37769_,
    new_n37770_, new_n37771_, new_n37772_, new_n37773_, new_n37774_,
    new_n37775_, new_n37776_, new_n37777_, new_n37778_, new_n37779_,
    new_n37780_, new_n37781_, new_n37782_, new_n37783_, new_n37784_,
    new_n37785_, new_n37786_, new_n37787_, new_n37788_, new_n37789_,
    new_n37790_, new_n37791_, new_n37792_, new_n37793_, new_n37794_,
    new_n37795_, new_n37796_, new_n37797_, new_n37798_, new_n37799_,
    new_n37800_, new_n37801_, new_n37802_, new_n37803_, new_n37804_,
    new_n37805_, new_n37806_, new_n37807_, new_n37808_, new_n37809_,
    new_n37810_, new_n37811_, new_n37812_, new_n37813_, new_n37814_,
    new_n37815_, new_n37816_, new_n37817_, new_n37818_, new_n37819_,
    new_n37820_, new_n37821_, new_n37822_, new_n37823_, new_n37824_,
    new_n37825_, new_n37826_, new_n37827_, new_n37828_, new_n37829_,
    new_n37830_, new_n37831_, new_n37832_, new_n37833_, new_n37834_,
    new_n37835_, new_n37836_, new_n37837_, new_n37838_, new_n37839_,
    new_n37840_, new_n37841_, new_n37842_, new_n37843_, new_n37844_,
    new_n37845_, new_n37846_, new_n37847_, new_n37848_, new_n37849_,
    new_n37850_, new_n37851_, new_n37852_, new_n37853_, new_n37854_,
    new_n37855_, new_n37856_, new_n37857_, new_n37858_, new_n37859_,
    new_n37860_, new_n37861_, new_n37862_, new_n37863_, new_n37864_,
    new_n37865_, new_n37866_, new_n37867_, new_n37868_, new_n37869_,
    new_n37870_, new_n37871_, new_n37872_, new_n37873_, new_n37874_,
    new_n37875_, new_n37876_, new_n37877_, new_n37878_, new_n37879_,
    new_n37880_, new_n37881_, new_n37882_, new_n37883_, new_n37884_,
    new_n37885_, new_n37886_, new_n37887_, new_n37888_, new_n37889_,
    new_n37890_, new_n37891_, new_n37892_, new_n37893_, new_n37894_,
    new_n37895_, new_n37896_, new_n37897_, new_n37898_, new_n37899_,
    new_n37900_, new_n37901_, new_n37902_, new_n37903_, new_n37904_,
    new_n37905_, new_n37906_, new_n37907_, new_n37908_, new_n37909_,
    new_n37910_, new_n37911_, new_n37912_, new_n37913_, new_n37914_,
    new_n37915_, new_n37916_, new_n37917_, new_n37918_, new_n37919_,
    new_n37920_, new_n37921_, new_n37922_, new_n37923_, new_n37924_,
    new_n37925_, new_n37926_, new_n37927_, new_n37928_, new_n37929_,
    new_n37930_, new_n37931_, new_n37932_, new_n37933_, new_n37934_,
    new_n37935_, new_n37936_, new_n37937_, new_n37938_, new_n37939_,
    new_n37940_, new_n37941_, new_n37942_, new_n37943_, new_n37944_,
    new_n37945_, new_n37946_, new_n37947_, new_n37948_, new_n37949_,
    new_n37950_, new_n37951_, new_n37952_, new_n37953_, new_n37954_,
    new_n37955_, new_n37956_, new_n37957_, new_n37958_, new_n37959_,
    new_n37960_, new_n37961_, new_n37962_, new_n37963_, new_n37964_,
    new_n37965_, new_n37966_, new_n37967_, new_n37968_, new_n37969_,
    new_n37970_, new_n37971_, new_n37972_, new_n37973_, new_n37974_,
    new_n37975_, new_n37976_, new_n37977_, new_n37978_, new_n37979_,
    new_n37980_, new_n37981_, new_n37982_, new_n37983_, new_n37984_,
    new_n37985_, new_n37986_, new_n37987_, new_n37988_, new_n37989_,
    new_n37990_, new_n37991_, new_n37992_, new_n37993_, new_n37994_,
    new_n37995_, new_n37996_, new_n37997_, new_n37998_, new_n37999_,
    new_n38000_, new_n38001_, new_n38002_, new_n38003_, new_n38004_,
    new_n38005_, new_n38006_, new_n38007_, new_n38008_, new_n38009_,
    new_n38010_, new_n38011_, new_n38012_, new_n38013_, new_n38014_,
    new_n38015_, new_n38016_, new_n38017_, new_n38018_, new_n38019_,
    new_n38020_, new_n38021_, new_n38022_, new_n38023_, new_n38024_,
    new_n38025_, new_n38026_, new_n38027_, new_n38028_, new_n38029_,
    new_n38030_, new_n38031_, new_n38032_, new_n38033_, new_n38034_,
    new_n38035_, new_n38036_, new_n38037_, new_n38038_, new_n38039_,
    new_n38040_, new_n38041_, new_n38042_, new_n38043_, new_n38044_,
    new_n38045_, new_n38046_, new_n38048_, new_n38049_, new_n38050_,
    new_n38051_, new_n38052_, new_n38053_, new_n38054_, new_n38055_,
    new_n38056_, new_n38057_, new_n38058_, new_n38059_, new_n38060_,
    new_n38061_, new_n38062_, new_n38063_, new_n38064_, new_n38065_,
    new_n38066_, new_n38067_, new_n38068_, new_n38069_, new_n38070_,
    new_n38071_, new_n38072_, new_n38073_, new_n38074_, new_n38075_,
    new_n38076_, new_n38077_, new_n38078_, new_n38079_, new_n38080_,
    new_n38081_, new_n38082_, new_n38083_, new_n38084_, new_n38085_,
    new_n38086_, new_n38087_, new_n38088_, new_n38089_, new_n38090_,
    new_n38091_, new_n38092_, new_n38093_, new_n38094_, new_n38095_,
    new_n38096_, new_n38097_, new_n38098_, new_n38099_, new_n38100_,
    new_n38101_, new_n38102_, new_n38103_, new_n38104_, new_n38105_,
    new_n38106_, new_n38107_, new_n38108_, new_n38109_, new_n38110_,
    new_n38111_, new_n38112_, new_n38113_, new_n38114_, new_n38115_,
    new_n38116_, new_n38117_, new_n38118_, new_n38119_, new_n38120_,
    new_n38121_, new_n38122_, new_n38123_, new_n38124_, new_n38125_,
    new_n38126_, new_n38127_, new_n38128_, new_n38129_, new_n38130_,
    new_n38131_, new_n38132_, new_n38133_, new_n38134_, new_n38135_,
    new_n38136_, new_n38137_, new_n38138_, new_n38139_, new_n38140_,
    new_n38141_, new_n38142_, new_n38143_, new_n38144_, new_n38145_,
    new_n38146_, new_n38147_, new_n38148_, new_n38149_, new_n38150_,
    new_n38151_, new_n38152_, new_n38153_, new_n38154_, new_n38155_,
    new_n38156_, new_n38157_, new_n38158_, new_n38159_, new_n38160_,
    new_n38161_, new_n38162_, new_n38163_, new_n38164_, new_n38165_,
    new_n38166_, new_n38167_, new_n38168_, new_n38169_, new_n38170_,
    new_n38171_, new_n38173_, new_n38174_, new_n38175_, new_n38176_,
    new_n38177_, new_n38178_, new_n38179_, new_n38180_, new_n38181_,
    new_n38182_, new_n38183_, new_n38184_, new_n38185_, new_n38186_,
    new_n38187_, new_n38188_, new_n38189_, new_n38190_, new_n38191_,
    new_n38192_, new_n38193_, new_n38194_, new_n38195_, new_n38196_,
    new_n38197_, new_n38198_, new_n38199_, new_n38200_, new_n38201_,
    new_n38202_, new_n38203_, new_n38204_, new_n38205_, new_n38206_,
    new_n38207_, new_n38208_, new_n38209_, new_n38210_, new_n38211_,
    new_n38212_, new_n38213_, new_n38214_, new_n38215_, new_n38216_,
    new_n38217_, new_n38218_, new_n38219_, new_n38220_, new_n38221_,
    new_n38222_, new_n38223_, new_n38224_, new_n38226_, new_n38227_,
    new_n38228_, new_n38229_, new_n38230_, new_n38231_, new_n38232_,
    new_n38233_, new_n38234_, new_n38235_, new_n38236_, new_n38237_,
    new_n38238_, new_n38239_, new_n38240_, new_n38241_, new_n38242_,
    new_n38243_, new_n38244_, new_n38245_, new_n38246_, new_n38247_,
    new_n38248_, new_n38249_, new_n38250_, new_n38251_, new_n38252_,
    new_n38253_, new_n38254_, new_n38255_, new_n38257_, new_n38258_,
    new_n38259_, new_n38260_, new_n38261_, new_n38262_, new_n38263_,
    new_n38264_, new_n38265_, new_n38266_, new_n38267_, new_n38269_,
    new_n38270_, new_n38271_, new_n38272_, new_n38273_, new_n38274_,
    new_n38275_, new_n38276_, new_n38277_, new_n38278_, new_n38279_,
    new_n38280_, new_n38281_, new_n38282_, new_n38283_, new_n38284_,
    new_n38285_, new_n38286_, new_n38287_, new_n38288_, new_n38289_,
    new_n38290_, new_n38291_, new_n38292_, new_n38293_, new_n38294_,
    new_n38295_, new_n38296_, new_n38297_, new_n38298_, new_n38299_,
    new_n38300_, new_n38301_, new_n38302_, new_n38303_, new_n38304_,
    new_n38305_, new_n38306_, new_n38307_, new_n38308_, new_n38309_,
    new_n38310_, new_n38311_, new_n38312_, new_n38313_, new_n38314_,
    new_n38315_, new_n38316_, new_n38317_, new_n38318_, new_n38319_,
    new_n38320_, new_n38321_, new_n38322_, new_n38323_, new_n38324_,
    new_n38325_, new_n38326_, new_n38327_, new_n38328_, new_n38329_,
    new_n38330_, new_n38331_, new_n38332_, new_n38333_, new_n38334_,
    new_n38335_, new_n38336_, new_n38337_, new_n38338_, new_n38339_,
    new_n38340_, new_n38341_, new_n38342_, new_n38343_, new_n38344_,
    new_n38345_, new_n38346_, new_n38347_, new_n38348_, new_n38349_,
    new_n38350_, new_n38352_, new_n38353_, new_n38354_, new_n38355_,
    new_n38356_, new_n38357_, new_n38358_, new_n38359_, new_n38360_,
    new_n38361_, new_n38362_, new_n38363_, new_n38364_, new_n38365_,
    new_n38366_, new_n38367_, new_n38368_, new_n38369_, new_n38370_,
    new_n38371_, new_n38372_, new_n38373_, new_n38374_, new_n38375_,
    new_n38376_, new_n38377_, new_n38378_, new_n38379_, new_n38380_,
    new_n38381_, new_n38382_, new_n38383_, new_n38384_, new_n38385_,
    new_n38386_, new_n38387_, new_n38389_, new_n38390_, new_n38391_,
    new_n38392_, new_n38393_, new_n38394_, new_n38395_, new_n38396_,
    new_n38397_, new_n38398_, new_n38399_, new_n38400_, new_n38401_,
    new_n38402_, new_n38403_, new_n38404_, new_n38405_, new_n38406_,
    new_n38407_, new_n38408_, new_n38409_, new_n38410_, new_n38412_,
    new_n38413_, new_n38414_, new_n38415_, new_n38416_, new_n38417_,
    new_n38418_, new_n38419_, new_n38420_, new_n38421_, new_n38422_,
    new_n38423_, new_n38424_, new_n38425_, new_n38426_, new_n38427_,
    new_n38428_, new_n38429_, new_n38430_, new_n38431_, new_n38432_,
    new_n38433_, new_n38434_, new_n38435_, new_n38436_, new_n38437_,
    new_n38438_, new_n38439_, new_n38440_, new_n38441_, new_n38442_,
    new_n38443_, new_n38444_, new_n38445_, new_n38446_, new_n38447_,
    new_n38448_, new_n38449_, new_n38450_, new_n38451_, new_n38452_,
    new_n38453_, new_n38454_, new_n38455_, new_n38456_, new_n38457_,
    new_n38458_, new_n38459_, new_n38460_, new_n38461_, new_n38462_,
    new_n38463_, new_n38464_, new_n38465_, new_n38466_, new_n38467_,
    new_n38468_, new_n38469_, new_n38470_, new_n38471_, new_n38472_,
    new_n38473_, new_n38474_, new_n38475_, new_n38476_, new_n38477_,
    new_n38478_, new_n38479_, new_n38480_, new_n38481_, new_n38482_,
    new_n38483_, new_n38484_, new_n38485_, new_n38486_, new_n38487_,
    new_n38488_, new_n38489_, new_n38490_, new_n38491_, new_n38492_,
    new_n38493_, new_n38494_, new_n38495_, new_n38496_, new_n38497_,
    new_n38498_, new_n38499_, new_n38500_, new_n38501_, new_n38502_,
    new_n38503_, new_n38504_, new_n38505_, new_n38506_, new_n38507_,
    new_n38508_, new_n38509_, new_n38510_, new_n38511_, new_n38512_,
    new_n38513_, new_n38514_, new_n38515_, new_n38516_, new_n38517_,
    new_n38518_, new_n38519_, new_n38520_, new_n38521_, new_n38522_,
    new_n38523_, new_n38524_, new_n38525_, new_n38526_, new_n38527_,
    new_n38528_, new_n38529_, new_n38530_, new_n38531_, new_n38532_,
    new_n38533_, new_n38534_, new_n38535_, new_n38536_, new_n38537_,
    new_n38538_, new_n38539_, new_n38540_, new_n38541_, new_n38542_,
    new_n38543_, new_n38544_, new_n38545_, new_n38546_, new_n38547_,
    new_n38548_, new_n38549_, new_n38550_, new_n38551_, new_n38552_,
    new_n38553_, new_n38554_, new_n38555_, new_n38556_, new_n38557_,
    new_n38558_, new_n38559_, new_n38560_, new_n38561_, new_n38562_,
    new_n38563_, new_n38564_, new_n38565_, new_n38566_, new_n38567_,
    new_n38568_, new_n38569_, new_n38570_, new_n38571_, new_n38572_,
    new_n38573_, new_n38574_, new_n38575_, new_n38576_, new_n38577_,
    new_n38578_, new_n38579_, new_n38580_, new_n38581_, new_n38582_,
    new_n38583_, new_n38584_, new_n38585_, new_n38586_, new_n38587_,
    new_n38588_, new_n38589_, new_n38590_, new_n38591_, new_n38592_,
    new_n38593_, new_n38594_, new_n38595_, new_n38596_, new_n38597_,
    new_n38598_, new_n38599_, new_n38600_, new_n38601_, new_n38602_,
    new_n38603_, new_n38604_, new_n38605_, new_n38606_, new_n38607_,
    new_n38608_, new_n38609_, new_n38610_, new_n38611_, new_n38612_,
    new_n38613_, new_n38614_, new_n38615_, new_n38616_, new_n38617_,
    new_n38618_, new_n38619_, new_n38620_, new_n38621_, new_n38622_,
    new_n38623_, new_n38624_, new_n38625_, new_n38626_, new_n38627_,
    new_n38628_, new_n38629_, new_n38630_, new_n38631_, new_n38632_,
    new_n38633_, new_n38634_, new_n38635_, new_n38636_, new_n38637_,
    new_n38638_, new_n38639_, new_n38640_, new_n38641_, new_n38642_,
    new_n38643_, new_n38644_, new_n38645_, new_n38646_, new_n38647_,
    new_n38648_, new_n38649_, new_n38650_, new_n38651_, new_n38652_,
    new_n38653_, new_n38654_, new_n38655_, new_n38656_, new_n38657_,
    new_n38658_, new_n38659_, new_n38660_, new_n38661_, new_n38662_,
    new_n38663_, new_n38664_, new_n38665_, new_n38666_, new_n38667_,
    new_n38668_, new_n38669_, new_n38670_, new_n38671_, new_n38672_,
    new_n38673_, new_n38674_, new_n38675_, new_n38676_, new_n38677_,
    new_n38678_, new_n38679_, new_n38680_, new_n38681_, new_n38682_,
    new_n38683_, new_n38684_, new_n38685_, new_n38686_, new_n38687_,
    new_n38688_, new_n38689_, new_n38690_, new_n38691_, new_n38692_,
    new_n38693_, new_n38694_, new_n38695_, new_n38696_, new_n38697_,
    new_n38698_, new_n38699_, new_n38700_, new_n38701_, new_n38702_,
    new_n38703_, new_n38704_, new_n38705_, new_n38706_, new_n38707_,
    new_n38708_, new_n38709_, new_n38710_, new_n38711_, new_n38712_,
    new_n38713_, new_n38714_, new_n38715_, new_n38716_, new_n38717_,
    new_n38718_, new_n38719_, new_n38720_, new_n38721_, new_n38722_,
    new_n38723_, new_n38724_, new_n38725_, new_n38726_, new_n38727_,
    new_n38728_, new_n38729_, new_n38730_, new_n38731_, new_n38732_,
    new_n38733_, new_n38734_, new_n38735_, new_n38736_, new_n38737_,
    new_n38738_, new_n38739_, new_n38740_, new_n38741_, new_n38742_,
    new_n38743_, new_n38744_, new_n38745_, new_n38746_, new_n38747_,
    new_n38748_, new_n38749_, new_n38750_, new_n38751_, new_n38752_,
    new_n38753_, new_n38754_, new_n38755_, new_n38756_, new_n38757_,
    new_n38758_, new_n38759_, new_n38760_, new_n38761_, new_n38762_,
    new_n38763_, new_n38764_, new_n38765_, new_n38766_, new_n38767_,
    new_n38768_, new_n38769_, new_n38770_, new_n38771_, new_n38772_,
    new_n38773_, new_n38774_, new_n38775_, new_n38776_, new_n38777_,
    new_n38778_, new_n38779_, new_n38780_, new_n38781_, new_n38782_,
    new_n38783_, new_n38784_, new_n38785_, new_n38786_, new_n38787_,
    new_n38788_, new_n38789_, new_n38790_, new_n38791_, new_n38792_,
    new_n38793_, new_n38794_, new_n38795_, new_n38796_, new_n38797_,
    new_n38798_, new_n38799_, new_n38800_, new_n38801_, new_n38802_,
    new_n38803_, new_n38804_, new_n38805_, new_n38806_, new_n38807_,
    new_n38808_, new_n38809_, new_n38810_, new_n38811_, new_n38812_,
    new_n38813_, new_n38814_, new_n38815_, new_n38816_, new_n38817_,
    new_n38818_, new_n38819_, new_n38820_, new_n38821_, new_n38822_,
    new_n38824_, new_n38825_, new_n38826_, new_n38827_, new_n38828_,
    new_n38829_, new_n38830_, new_n38831_, new_n38832_, new_n38833_,
    new_n38834_, new_n38835_, new_n38836_, new_n38837_, new_n38838_,
    new_n38839_, new_n38840_, new_n38841_, new_n38842_, new_n38843_,
    new_n38844_, new_n38845_, new_n38846_, new_n38847_, new_n38848_,
    new_n38849_, new_n38850_, new_n38851_, new_n38852_, new_n38853_,
    new_n38854_, new_n38855_, new_n38856_, new_n38857_, new_n38858_,
    new_n38859_, new_n38860_, new_n38861_, new_n38862_, new_n38863_,
    new_n38864_, new_n38865_, new_n38866_, new_n38867_, new_n38868_,
    new_n38869_, new_n38870_, new_n38871_, new_n38872_, new_n38873_,
    new_n38874_, new_n38875_, new_n38876_, new_n38877_, new_n38878_,
    new_n38879_, new_n38880_, new_n38881_, new_n38882_, new_n38883_,
    new_n38884_, new_n38885_, new_n38886_, new_n38887_, new_n38888_,
    new_n38889_, new_n38890_, new_n38891_, new_n38892_, new_n38893_,
    new_n38894_, new_n38895_, new_n38896_, new_n38897_, new_n38898_,
    new_n38899_, new_n38900_, new_n38901_, new_n38902_, new_n38903_,
    new_n38904_, new_n38905_, new_n38906_, new_n38907_, new_n38908_,
    new_n38909_, new_n38910_, new_n38911_, new_n38912_, new_n38913_,
    new_n38914_, new_n38915_, new_n38916_, new_n38917_, new_n38918_,
    new_n38919_, new_n38920_, new_n38921_, new_n38922_, new_n38923_,
    new_n38924_, new_n38925_, new_n38926_, new_n38927_, new_n38928_,
    new_n38929_, new_n38930_, new_n38931_, new_n38932_, new_n38933_,
    new_n38934_, new_n38935_, new_n38936_, new_n38937_, new_n38938_,
    new_n38939_, new_n38940_, new_n38941_, new_n38942_, new_n38943_,
    new_n38944_, new_n38945_, new_n38946_, new_n38947_, new_n38948_,
    new_n38949_, new_n38950_, new_n38951_, new_n38952_, new_n38953_,
    new_n38954_, new_n38955_, new_n38956_, new_n38957_, new_n38958_,
    new_n38959_, new_n38960_, new_n38961_, new_n38962_, new_n38963_,
    new_n38964_, new_n38965_, new_n38966_, new_n38967_, new_n38968_,
    new_n38969_, new_n38970_, new_n38971_, new_n38972_, new_n38973_,
    new_n38974_, new_n38975_, new_n38976_, new_n38977_, new_n38978_,
    new_n38979_, new_n38980_, new_n38981_, new_n38982_, new_n38983_,
    new_n38984_, new_n38985_, new_n38986_, new_n38987_, new_n38988_,
    new_n38989_, new_n38990_, new_n38991_, new_n38992_, new_n38993_,
    new_n38994_, new_n38995_, new_n38996_, new_n38997_, new_n38998_,
    new_n38999_, new_n39000_, new_n39001_, new_n39002_, new_n39003_,
    new_n39004_, new_n39005_, new_n39006_, new_n39007_, new_n39008_,
    new_n39009_, new_n39010_, new_n39011_, new_n39012_, new_n39013_,
    new_n39014_, new_n39015_, new_n39016_, new_n39017_, new_n39018_,
    new_n39019_, new_n39020_, new_n39021_, new_n39022_, new_n39023_,
    new_n39024_, new_n39025_, new_n39026_, new_n39027_, new_n39028_,
    new_n39029_, new_n39030_, new_n39031_, new_n39032_, new_n39033_,
    new_n39034_, new_n39035_, new_n39036_, new_n39037_, new_n39038_,
    new_n39039_, new_n39040_, new_n39041_, new_n39042_, new_n39043_,
    new_n39044_, new_n39045_, new_n39046_, new_n39047_, new_n39048_,
    new_n39049_, new_n39050_, new_n39051_, new_n39052_, new_n39053_,
    new_n39054_, new_n39055_, new_n39056_, new_n39057_, new_n39058_,
    new_n39059_, new_n39060_, new_n39061_, new_n39062_, new_n39063_,
    new_n39064_, new_n39065_, new_n39066_, new_n39067_, new_n39068_,
    new_n39069_, new_n39070_, new_n39071_, new_n39072_, new_n39073_,
    new_n39074_, new_n39075_, new_n39076_, new_n39077_, new_n39078_,
    new_n39079_, new_n39080_, new_n39081_, new_n39082_, new_n39083_,
    new_n39084_, new_n39085_, new_n39086_, new_n39087_, new_n39088_,
    new_n39089_, new_n39090_, new_n39091_, new_n39092_, new_n39093_,
    new_n39094_, new_n39095_, new_n39096_, new_n39097_, new_n39098_,
    new_n39099_, new_n39100_, new_n39101_, new_n39102_, new_n39103_,
    new_n39104_, new_n39105_, new_n39106_, new_n39107_, new_n39108_,
    new_n39109_, new_n39110_, new_n39111_, new_n39112_, new_n39113_,
    new_n39114_, new_n39115_, new_n39116_, new_n39117_, new_n39118_,
    new_n39119_, new_n39120_, new_n39121_, new_n39122_, new_n39123_,
    new_n39124_, new_n39125_, new_n39126_, new_n39127_, new_n39128_,
    new_n39129_, new_n39130_, new_n39131_, new_n39132_, new_n39133_,
    new_n39134_, new_n39135_, new_n39136_, new_n39137_, new_n39138_,
    new_n39139_, new_n39140_, new_n39141_, new_n39142_, new_n39143_,
    new_n39144_, new_n39145_, new_n39146_, new_n39147_, new_n39148_,
    new_n39149_, new_n39150_, new_n39151_, new_n39152_, new_n39153_,
    new_n39154_, new_n39155_, new_n39156_, new_n39158_, new_n39159_,
    new_n39160_, new_n39161_, new_n39162_, new_n39163_, new_n39164_,
    new_n39165_, new_n39166_, new_n39167_, new_n39168_, new_n39169_,
    new_n39170_, new_n39171_, new_n39172_, new_n39173_, new_n39174_,
    new_n39175_, new_n39176_, new_n39177_, new_n39178_, new_n39179_,
    new_n39180_, new_n39181_, new_n39182_, new_n39183_, new_n39184_,
    new_n39185_, new_n39186_, new_n39187_, new_n39188_, new_n39189_,
    new_n39190_, new_n39191_, new_n39192_, new_n39193_, new_n39194_,
    new_n39195_, new_n39196_, new_n39197_, new_n39198_, new_n39199_,
    new_n39200_, new_n39201_, new_n39202_, new_n39203_, new_n39204_,
    new_n39205_, new_n39206_, new_n39207_, new_n39208_, new_n39209_,
    new_n39210_, new_n39211_, new_n39212_, new_n39213_, new_n39214_,
    new_n39215_, new_n39216_, new_n39217_, new_n39218_, new_n39219_,
    new_n39220_, new_n39221_, new_n39222_, new_n39223_, new_n39224_,
    new_n39225_, new_n39226_, new_n39227_, new_n39228_, new_n39229_,
    new_n39230_, new_n39231_, new_n39232_, new_n39233_, new_n39234_,
    new_n39235_, new_n39236_, new_n39237_, new_n39238_, new_n39239_,
    new_n39240_, new_n39241_, new_n39242_, new_n39243_, new_n39244_,
    new_n39245_, new_n39246_, new_n39247_, new_n39248_, new_n39249_,
    new_n39250_, new_n39251_, new_n39252_, new_n39253_, new_n39254_,
    new_n39255_, new_n39256_, new_n39257_, new_n39258_, new_n39259_,
    new_n39260_, new_n39261_, new_n39262_, new_n39263_, new_n39264_,
    new_n39265_, new_n39266_, new_n39267_, new_n39268_, new_n39269_,
    new_n39270_, new_n39271_, new_n39272_, new_n39273_, new_n39274_,
    new_n39275_, new_n39276_, new_n39277_, new_n39278_, new_n39279_,
    new_n39280_, new_n39281_, new_n39282_, new_n39283_, new_n39284_,
    new_n39285_, new_n39286_, new_n39287_, new_n39288_, new_n39289_,
    new_n39290_, new_n39291_, new_n39292_, new_n39293_, new_n39294_,
    new_n39295_, new_n39296_, new_n39297_, new_n39298_, new_n39299_,
    new_n39300_, new_n39301_, new_n39302_, new_n39303_, new_n39304_,
    new_n39305_, new_n39306_, new_n39307_, new_n39308_, new_n39309_,
    new_n39310_, new_n39311_, new_n39312_, new_n39313_, new_n39314_,
    new_n39315_, new_n39316_, new_n39317_, new_n39318_, new_n39319_,
    new_n39320_, new_n39321_, new_n39322_, new_n39323_, new_n39324_,
    new_n39325_, new_n39326_, new_n39327_, new_n39328_, new_n39329_,
    new_n39330_, new_n39331_, new_n39332_, new_n39333_, new_n39334_,
    new_n39335_, new_n39336_, new_n39337_, new_n39338_, new_n39339_,
    new_n39340_, new_n39341_, new_n39342_, new_n39343_, new_n39344_,
    new_n39345_, new_n39346_, new_n39347_, new_n39348_, new_n39349_,
    new_n39350_, new_n39351_, new_n39352_, new_n39353_, new_n39354_,
    new_n39356_, new_n39357_, new_n39358_, new_n39359_, new_n39360_,
    new_n39361_, new_n39362_, new_n39363_, new_n39364_, new_n39365_,
    new_n39366_, new_n39367_, new_n39369_, new_n39370_, new_n39371_,
    new_n39372_, new_n39373_, new_n39374_, new_n39375_, new_n39376_,
    new_n39377_, new_n39378_, new_n39379_, new_n39380_, new_n39381_,
    new_n39382_, new_n39383_, new_n39384_, new_n39385_, new_n39386_,
    new_n39387_, new_n39388_, new_n39389_, new_n39390_, new_n39391_,
    new_n39392_, new_n39393_, new_n39394_, new_n39395_, new_n39396_,
    new_n39397_, new_n39398_, new_n39399_, new_n39400_, new_n39401_,
    new_n39402_, new_n39403_, new_n39404_, new_n39405_, new_n39406_,
    new_n39407_, new_n39408_, new_n39409_, new_n39410_, new_n39411_,
    new_n39412_, new_n39413_, new_n39414_, new_n39415_, new_n39416_,
    new_n39417_, new_n39418_, new_n39419_, new_n39420_, new_n39421_,
    new_n39422_, new_n39423_, new_n39424_, new_n39425_, new_n39426_,
    new_n39427_, new_n39428_, new_n39429_, new_n39430_, new_n39431_,
    new_n39432_, new_n39433_, new_n39434_, new_n39435_, new_n39436_,
    new_n39437_, new_n39438_, new_n39439_, new_n39440_, new_n39441_,
    new_n39442_, new_n39443_, new_n39444_, new_n39445_, new_n39446_,
    new_n39447_, new_n39448_, new_n39449_, new_n39450_, new_n39451_,
    new_n39452_, new_n39453_, new_n39454_, new_n39455_, new_n39456_,
    new_n39457_, new_n39458_, new_n39459_, new_n39460_, new_n39461_,
    new_n39462_, new_n39463_, new_n39464_, new_n39465_, new_n39466_,
    new_n39467_, new_n39468_, new_n39469_, new_n39470_, new_n39471_,
    new_n39472_, new_n39473_, new_n39474_, new_n39475_, new_n39476_,
    new_n39477_, new_n39478_, new_n39479_, new_n39480_, new_n39481_,
    new_n39482_, new_n39483_, new_n39484_, new_n39485_, new_n39486_,
    new_n39487_, new_n39488_, new_n39489_, new_n39490_, new_n39491_,
    new_n39492_, new_n39493_, new_n39494_, new_n39495_, new_n39496_,
    new_n39497_, new_n39498_, new_n39499_, new_n39500_, new_n39501_,
    new_n39502_, new_n39503_, new_n39504_, new_n39505_, new_n39506_,
    new_n39507_, new_n39508_, new_n39509_, new_n39510_, new_n39511_,
    new_n39512_, new_n39513_, new_n39514_, new_n39515_, new_n39516_,
    new_n39517_, new_n39518_, new_n39519_, new_n39520_, new_n39521_,
    new_n39522_, new_n39523_, new_n39524_, new_n39525_, new_n39526_,
    new_n39527_, new_n39528_, new_n39529_, new_n39530_, new_n39531_,
    new_n39532_, new_n39533_, new_n39534_, new_n39535_, new_n39536_,
    new_n39537_, new_n39538_, new_n39539_, new_n39540_, new_n39541_,
    new_n39542_, new_n39543_, new_n39544_, new_n39545_, new_n39546_,
    new_n39547_, new_n39548_, new_n39549_, new_n39550_, new_n39551_,
    new_n39552_, new_n39553_, new_n39554_, new_n39555_, new_n39556_,
    new_n39557_, new_n39558_, new_n39559_, new_n39560_, new_n39561_,
    new_n39562_, new_n39563_, new_n39564_, new_n39565_, new_n39566_,
    new_n39567_, new_n39568_, new_n39569_, new_n39570_, new_n39571_,
    new_n39572_, new_n39573_, new_n39574_, new_n39575_, new_n39576_,
    new_n39577_, new_n39578_, new_n39579_, new_n39580_, new_n39581_,
    new_n39582_, new_n39583_, new_n39584_, new_n39585_, new_n39586_,
    new_n39587_, new_n39588_, new_n39589_, new_n39590_, new_n39591_,
    new_n39592_, new_n39593_, new_n39594_, new_n39595_, new_n39596_,
    new_n39597_, new_n39598_, new_n39599_, new_n39600_, new_n39601_,
    new_n39602_, new_n39603_, new_n39604_, new_n39605_, new_n39606_,
    new_n39607_, new_n39608_, new_n39609_, new_n39610_, new_n39611_,
    new_n39612_, new_n39613_, new_n39614_, new_n39615_, new_n39616_,
    new_n39617_, new_n39618_, new_n39619_, new_n39620_, new_n39621_,
    new_n39622_, new_n39623_, new_n39624_, new_n39625_, new_n39626_,
    new_n39627_, new_n39628_, new_n39629_, new_n39631_, new_n39632_,
    new_n39633_, new_n39634_, new_n39635_, new_n39636_, new_n39637_,
    new_n39638_, new_n39639_, new_n39640_, new_n39641_, new_n39642_,
    new_n39643_, new_n39644_, new_n39645_, new_n39646_, new_n39647_,
    new_n39648_, new_n39649_, new_n39650_, new_n39651_, new_n39652_,
    new_n39653_, new_n39654_, new_n39655_, new_n39656_, new_n39657_,
    new_n39658_, new_n39659_, new_n39660_, new_n39661_, new_n39662_,
    new_n39663_, new_n39664_, new_n39665_, new_n39666_, new_n39667_,
    new_n39668_, new_n39669_, new_n39670_, new_n39671_, new_n39672_,
    new_n39673_, new_n39674_, new_n39675_, new_n39676_, new_n39677_,
    new_n39678_, new_n39679_, new_n39680_, new_n39681_, new_n39682_,
    new_n39683_, new_n39684_, new_n39685_, new_n39686_, new_n39687_,
    new_n39688_, new_n39689_, new_n39690_, new_n39691_, new_n39692_,
    new_n39693_, new_n39694_, new_n39695_, new_n39696_, new_n39697_,
    new_n39698_, new_n39699_, new_n39700_, new_n39701_, new_n39702_,
    new_n39703_, new_n39704_, new_n39705_, new_n39706_, new_n39707_,
    new_n39708_, new_n39709_, new_n39710_, new_n39711_, new_n39712_,
    new_n39713_, new_n39714_, new_n39715_, new_n39716_, new_n39717_,
    new_n39718_, new_n39719_, new_n39720_, new_n39721_, new_n39722_,
    new_n39723_, new_n39724_, new_n39725_, new_n39726_, new_n39727_,
    new_n39728_, new_n39729_, new_n39730_, new_n39731_, new_n39732_,
    new_n39733_, new_n39734_, new_n39735_, new_n39736_, new_n39737_,
    new_n39738_, new_n39739_, new_n39740_, new_n39741_, new_n39742_,
    new_n39743_, new_n39744_, new_n39745_, new_n39746_, new_n39747_,
    new_n39748_, new_n39749_, new_n39750_, new_n39751_, new_n39752_,
    new_n39753_, new_n39754_, new_n39755_, new_n39756_, new_n39757_,
    new_n39758_, new_n39759_, new_n39760_, new_n39761_, new_n39762_,
    new_n39763_, new_n39764_, new_n39765_, new_n39766_, new_n39767_,
    new_n39768_, new_n39769_, new_n39770_, new_n39771_, new_n39772_,
    new_n39773_, new_n39774_, new_n39775_, new_n39776_, new_n39777_,
    new_n39778_, new_n39779_, new_n39780_, new_n39781_, new_n39782_,
    new_n39783_, new_n39784_, new_n39785_, new_n39786_, new_n39787_,
    new_n39788_, new_n39789_, new_n39790_, new_n39791_, new_n39792_,
    new_n39793_, new_n39794_, new_n39795_, new_n39796_, new_n39797_,
    new_n39798_, new_n39799_, new_n39800_, new_n39801_, new_n39802_,
    new_n39803_, new_n39804_, new_n39805_, new_n39806_, new_n39807_,
    new_n39808_, new_n39809_, new_n39810_, new_n39811_, new_n39812_,
    new_n39813_, new_n39814_, new_n39815_, new_n39816_, new_n39817_,
    new_n39818_, new_n39819_, new_n39820_, new_n39821_, new_n39822_,
    new_n39823_, new_n39824_, new_n39825_, new_n39826_, new_n39827_,
    new_n39828_, new_n39829_, new_n39830_, new_n39831_, new_n39832_,
    new_n39833_, new_n39834_, new_n39835_, new_n39836_, new_n39837_,
    new_n39838_, new_n39839_, new_n39840_, new_n39841_, new_n39842_,
    new_n39843_, new_n39844_, new_n39845_, new_n39846_, new_n39847_,
    new_n39848_, new_n39849_, new_n39850_, new_n39851_, new_n39852_,
    new_n39853_, new_n39854_, new_n39855_, new_n39856_, new_n39857_,
    new_n39858_, new_n39859_, new_n39860_, new_n39861_, new_n39862_,
    new_n39863_, new_n39864_, new_n39865_, new_n39866_, new_n39867_,
    new_n39868_, new_n39869_, new_n39870_, new_n39871_, new_n39872_,
    new_n39873_, new_n39874_, new_n39875_, new_n39876_, new_n39877_,
    new_n39878_, new_n39879_, new_n39880_, new_n39881_, new_n39882_,
    new_n39883_, new_n39884_, new_n39885_, new_n39886_, new_n39887_,
    new_n39888_, new_n39889_, new_n39890_, new_n39891_, new_n39892_,
    new_n39893_, new_n39894_, new_n39895_, new_n39896_, new_n39897_,
    new_n39898_, new_n39899_, new_n39900_, new_n39901_, new_n39902_,
    new_n39903_, new_n39904_, new_n39905_, new_n39906_, new_n39907_,
    new_n39908_, new_n39909_, new_n39910_, new_n39911_, new_n39912_,
    new_n39913_, new_n39914_, new_n39915_, new_n39916_, new_n39917_,
    new_n39918_, new_n39919_, new_n39920_, new_n39921_, new_n39922_,
    new_n39923_, new_n39924_, new_n39925_, new_n39926_, new_n39927_,
    new_n39928_, new_n39929_, new_n39930_, new_n39931_, new_n39932_,
    new_n39933_, new_n39934_, new_n39935_, new_n39936_, new_n39937_,
    new_n39938_, new_n39939_, new_n39940_, new_n39941_, new_n39942_,
    new_n39943_, new_n39944_, new_n39945_, new_n39946_, new_n39947_,
    new_n39948_, new_n39949_, new_n39950_, new_n39951_, new_n39952_,
    new_n39953_, new_n39954_, new_n39955_, new_n39956_, new_n39957_,
    new_n39958_, new_n39959_, new_n39960_, new_n39961_, new_n39962_,
    new_n39963_, new_n39964_, new_n39965_, new_n39966_, new_n39967_,
    new_n39969_, new_n39970_, new_n39971_, new_n39972_, new_n39973_,
    new_n39974_, new_n39975_, new_n39976_, new_n39977_, new_n39978_,
    new_n39979_, new_n39980_, new_n39981_, new_n39982_, new_n39983_,
    new_n39984_, new_n39985_, new_n39986_, new_n39987_, new_n39988_,
    new_n39989_, new_n39990_, new_n39991_, new_n39992_, new_n39993_,
    new_n39994_, new_n39995_, new_n39996_, new_n39997_, new_n39998_,
    new_n39999_, new_n40000_, new_n40001_, new_n40002_, new_n40003_,
    new_n40004_, new_n40005_, new_n40006_, new_n40007_, new_n40008_,
    new_n40009_, new_n40010_, new_n40011_, new_n40012_, new_n40013_,
    new_n40014_, new_n40015_, new_n40016_, new_n40017_, new_n40018_,
    new_n40019_, new_n40020_, new_n40021_, new_n40022_, new_n40023_,
    new_n40024_, new_n40025_, new_n40026_, new_n40027_, new_n40028_,
    new_n40029_, new_n40030_, new_n40031_, new_n40032_, new_n40033_,
    new_n40034_, new_n40035_, new_n40036_, new_n40037_, new_n40038_,
    new_n40039_, new_n40040_, new_n40041_, new_n40042_, new_n40043_,
    new_n40044_, new_n40045_, new_n40046_, new_n40047_, new_n40048_,
    new_n40049_, new_n40050_, new_n40051_, new_n40052_, new_n40053_,
    new_n40054_, new_n40055_, new_n40056_, new_n40057_, new_n40058_,
    new_n40060_, new_n40061_, new_n40062_, new_n40063_, new_n40064_,
    new_n40065_, new_n40066_, new_n40067_, new_n40068_, new_n40069_,
    new_n40070_, new_n40071_, new_n40072_, new_n40073_, new_n40074_,
    new_n40075_, new_n40076_, new_n40077_, new_n40078_, new_n40079_,
    new_n40080_, new_n40081_, new_n40082_, new_n40083_, new_n40084_,
    new_n40085_, new_n40086_, new_n40087_, new_n40088_, new_n40089_,
    new_n40090_, new_n40091_, new_n40092_, new_n40093_, new_n40094_,
    new_n40095_, new_n40096_, new_n40097_, new_n40098_, new_n40099_,
    new_n40100_, new_n40101_, new_n40102_, new_n40103_, new_n40104_,
    new_n40105_, new_n40106_, new_n40107_, new_n40108_, new_n40109_,
    new_n40110_, new_n40111_, new_n40112_, new_n40113_, new_n40114_,
    new_n40115_, new_n40116_, new_n40117_, new_n40118_, new_n40119_,
    new_n40120_, new_n40121_, new_n40122_, new_n40123_, new_n40124_,
    new_n40125_, new_n40126_, new_n40127_, new_n40128_, new_n40129_,
    new_n40130_, new_n40131_, new_n40132_, new_n40133_, new_n40134_,
    new_n40135_, new_n40136_, new_n40137_, new_n40138_, new_n40139_,
    new_n40140_, new_n40141_, new_n40142_, new_n40143_, new_n40144_,
    new_n40145_, new_n40146_, new_n40147_, new_n40148_, new_n40149_,
    new_n40150_, new_n40151_, new_n40152_, new_n40153_, new_n40154_,
    new_n40155_, new_n40156_, new_n40157_, new_n40158_, new_n40159_,
    new_n40160_, new_n40161_, new_n40162_, new_n40163_, new_n40164_,
    new_n40165_, new_n40166_, new_n40167_, new_n40168_, new_n40169_,
    new_n40170_, new_n40171_, new_n40172_, new_n40173_, new_n40174_,
    new_n40175_, new_n40176_, new_n40177_, new_n40178_, new_n40179_,
    new_n40180_, new_n40181_, new_n40182_, new_n40183_, new_n40184_,
    new_n40185_, new_n40186_, new_n40187_, new_n40188_, new_n40189_,
    new_n40190_, new_n40191_, new_n40192_, new_n40193_, new_n40194_,
    new_n40195_, new_n40196_, new_n40197_, new_n40198_, new_n40199_,
    new_n40200_, new_n40201_, new_n40202_, new_n40203_, new_n40204_,
    new_n40205_, new_n40206_, new_n40207_, new_n40208_, new_n40209_,
    new_n40210_, new_n40211_, new_n40212_, new_n40213_, new_n40214_,
    new_n40215_, new_n40216_, new_n40217_, new_n40218_, new_n40219_,
    new_n40220_, new_n40221_, new_n40222_, new_n40223_, new_n40224_,
    new_n40225_, new_n40226_, new_n40227_, new_n40228_, new_n40229_,
    new_n40230_, new_n40231_, new_n40232_, new_n40233_, new_n40234_,
    new_n40235_, new_n40236_, new_n40237_, new_n40238_, new_n40239_,
    new_n40240_, new_n40241_, new_n40242_, new_n40243_, new_n40244_,
    new_n40245_, new_n40246_, new_n40247_, new_n40248_, new_n40249_,
    new_n40250_, new_n40251_, new_n40252_, new_n40253_, new_n40254_,
    new_n40255_, new_n40256_, new_n40257_, new_n40258_, new_n40259_,
    new_n40260_, new_n40261_, new_n40262_, new_n40263_, new_n40264_,
    new_n40265_, new_n40266_, new_n40267_, new_n40268_, new_n40269_,
    new_n40270_, new_n40271_, new_n40272_, new_n40273_, new_n40274_,
    new_n40275_, new_n40276_, new_n40277_, new_n40278_, new_n40279_,
    new_n40280_, new_n40281_, new_n40282_, new_n40283_, new_n40284_,
    new_n40285_, new_n40286_, new_n40287_, new_n40288_, new_n40289_,
    new_n40290_, new_n40291_, new_n40292_, new_n40293_, new_n40294_,
    new_n40295_, new_n40296_, new_n40297_, new_n40298_, new_n40299_,
    new_n40300_, new_n40301_, new_n40302_, new_n40303_, new_n40304_,
    new_n40305_, new_n40306_, new_n40307_, new_n40308_, new_n40309_,
    new_n40310_, new_n40311_, new_n40312_, new_n40313_, new_n40314_,
    new_n40315_, new_n40316_, new_n40317_, new_n40318_, new_n40319_,
    new_n40320_, new_n40321_, new_n40322_, new_n40323_, new_n40324_,
    new_n40325_, new_n40326_, new_n40327_, new_n40328_, new_n40329_,
    new_n40330_, new_n40331_, new_n40332_, new_n40333_, new_n40334_,
    new_n40335_, new_n40336_, new_n40337_, new_n40338_, new_n40339_,
    new_n40340_, new_n40341_, new_n40342_, new_n40343_, new_n40344_,
    new_n40345_, new_n40346_, new_n40347_, new_n40348_, new_n40349_,
    new_n40350_, new_n40351_, new_n40352_, new_n40353_, new_n40354_,
    new_n40355_, new_n40356_, new_n40357_, new_n40358_, new_n40359_,
    new_n40360_, new_n40361_, new_n40362_, new_n40363_, new_n40364_,
    new_n40365_, new_n40366_, new_n40367_, new_n40368_, new_n40369_,
    new_n40370_, new_n40371_, new_n40372_, new_n40373_, new_n40374_,
    new_n40375_, new_n40376_, new_n40377_, new_n40378_, new_n40379_,
    new_n40380_, new_n40381_, new_n40382_, new_n40383_, new_n40384_,
    new_n40385_, new_n40386_, new_n40387_, new_n40388_, new_n40389_,
    new_n40390_, new_n40391_, new_n40392_, new_n40393_, new_n40394_,
    new_n40395_, new_n40396_, new_n40397_, new_n40398_, new_n40399_,
    new_n40400_, new_n40401_, new_n40402_, new_n40403_, new_n40404_,
    new_n40405_, new_n40406_, new_n40407_, new_n40408_, new_n40409_,
    new_n40410_, new_n40411_, new_n40412_, new_n40413_, new_n40414_,
    new_n40415_, new_n40416_, new_n40417_, new_n40418_, new_n40419_,
    new_n40420_, new_n40421_, new_n40422_, new_n40423_, new_n40424_,
    new_n40425_, new_n40426_, new_n40427_, new_n40428_, new_n40429_,
    new_n40430_, new_n40431_, new_n40432_, new_n40433_, new_n40434_,
    new_n40435_, new_n40436_, new_n40437_, new_n40438_, new_n40439_,
    new_n40440_, new_n40441_, new_n40442_, new_n40443_, new_n40444_,
    new_n40445_, new_n40446_, new_n40447_, new_n40448_, new_n40449_,
    new_n40450_, new_n40451_, new_n40452_, new_n40453_, new_n40454_,
    new_n40455_, new_n40456_, new_n40457_, new_n40458_, new_n40459_,
    new_n40460_, new_n40461_, new_n40462_, new_n40463_, new_n40464_,
    new_n40465_, new_n40466_, new_n40467_, new_n40468_, new_n40469_,
    new_n40470_, new_n40471_, new_n40472_, new_n40473_, new_n40474_,
    new_n40475_, new_n40476_, new_n40477_, new_n40478_, new_n40479_,
    new_n40481_, new_n40482_, new_n40483_, new_n40484_, new_n40485_,
    new_n40486_, new_n40487_, new_n40488_, new_n40489_, new_n40490_,
    new_n40491_, new_n40492_, new_n40493_, new_n40494_, new_n40495_,
    new_n40496_, new_n40497_, new_n40498_, new_n40499_, new_n40500_,
    new_n40501_, new_n40502_, new_n40503_, new_n40504_, new_n40505_,
    new_n40506_, new_n40507_, new_n40508_, new_n40509_, new_n40510_,
    new_n40511_, new_n40512_, new_n40513_, new_n40514_, new_n40515_,
    new_n40516_, new_n40517_, new_n40518_, new_n40519_, new_n40520_,
    new_n40521_, new_n40522_, new_n40523_, new_n40524_, new_n40525_,
    new_n40526_, new_n40527_, new_n40528_, new_n40529_, new_n40530_,
    new_n40531_, new_n40532_, new_n40533_, new_n40534_, new_n40535_,
    new_n40536_, new_n40537_, new_n40538_, new_n40539_, new_n40540_,
    new_n40541_, new_n40542_, new_n40543_, new_n40544_, new_n40545_,
    new_n40546_, new_n40547_, new_n40548_, new_n40549_, new_n40550_,
    new_n40551_, new_n40552_, new_n40553_, new_n40554_, new_n40555_,
    new_n40556_, new_n40557_, new_n40558_, new_n40559_, new_n40560_,
    new_n40561_, new_n40562_, new_n40563_, new_n40564_, new_n40565_,
    new_n40566_, new_n40567_, new_n40568_, new_n40569_, new_n40570_,
    new_n40571_, new_n40572_, new_n40573_, new_n40574_, new_n40575_,
    new_n40576_, new_n40577_, new_n40578_, new_n40579_, new_n40580_,
    new_n40581_, new_n40582_, new_n40583_, new_n40584_, new_n40585_,
    new_n40586_, new_n40587_, new_n40588_, new_n40589_, new_n40590_,
    new_n40591_, new_n40592_, new_n40593_, new_n40594_, new_n40595_,
    new_n40596_, new_n40597_, new_n40598_, new_n40599_, new_n40600_,
    new_n40601_, new_n40602_, new_n40603_, new_n40604_, new_n40605_,
    new_n40606_, new_n40607_, new_n40608_, new_n40609_, new_n40610_,
    new_n40611_, new_n40612_, new_n40613_, new_n40614_, new_n40615_,
    new_n40616_, new_n40617_, new_n40618_, new_n40619_, new_n40620_,
    new_n40621_, new_n40622_, new_n40623_, new_n40624_, new_n40625_,
    new_n40626_, new_n40627_, new_n40628_, new_n40629_, new_n40630_,
    new_n40631_, new_n40632_, new_n40633_, new_n40634_, new_n40635_,
    new_n40636_, new_n40637_, new_n40638_, new_n40639_, new_n40640_,
    new_n40641_, new_n40642_, new_n40643_, new_n40644_, new_n40645_,
    new_n40646_, new_n40647_, new_n40648_, new_n40649_, new_n40650_,
    new_n40651_, new_n40652_, new_n40653_, new_n40654_, new_n40655_,
    new_n40656_, new_n40657_, new_n40658_, new_n40659_, new_n40660_,
    new_n40661_, new_n40662_, new_n40663_, new_n40664_, new_n40665_,
    new_n40666_, new_n40667_, new_n40668_, new_n40669_, new_n40670_,
    new_n40671_, new_n40672_, new_n40673_, new_n40674_, new_n40675_,
    new_n40676_, new_n40677_, new_n40678_, new_n40679_, new_n40680_,
    new_n40681_, new_n40682_, new_n40683_, new_n40684_, new_n40685_,
    new_n40686_, new_n40687_, new_n40688_, new_n40689_, new_n40690_,
    new_n40691_, new_n40692_, new_n40693_, new_n40694_, new_n40695_,
    new_n40696_, new_n40697_, new_n40698_, new_n40699_, new_n40700_,
    new_n40701_, new_n40702_, new_n40703_, new_n40704_, new_n40705_,
    new_n40706_, new_n40707_, new_n40708_, new_n40709_, new_n40710_,
    new_n40711_, new_n40712_, new_n40713_, new_n40714_, new_n40715_,
    new_n40716_, new_n40717_, new_n40718_, new_n40719_, new_n40720_,
    new_n40721_, new_n40722_, new_n40723_, new_n40724_, new_n40725_,
    new_n40726_, new_n40727_, new_n40728_, new_n40729_, new_n40730_,
    new_n40731_, new_n40732_, new_n40733_, new_n40734_, new_n40735_,
    new_n40736_, new_n40737_, new_n40738_, new_n40739_, new_n40740_,
    new_n40741_, new_n40742_, new_n40743_, new_n40744_, new_n40745_,
    new_n40746_, new_n40747_, new_n40748_, new_n40749_, new_n40750_,
    new_n40751_, new_n40752_, new_n40753_, new_n40754_, new_n40755_,
    new_n40756_, new_n40757_, new_n40758_, new_n40759_, new_n40760_,
    new_n40761_, new_n40762_, new_n40763_, new_n40764_, new_n40765_,
    new_n40766_, new_n40767_, new_n40768_, new_n40770_, new_n40771_,
    new_n40772_, new_n40773_, new_n40774_, new_n40775_, new_n40776_,
    new_n40777_, new_n40778_, new_n40779_, new_n40780_, new_n40781_,
    new_n40782_, new_n40783_, new_n40784_, new_n40785_, new_n40786_,
    new_n40787_, new_n40788_, new_n40789_, new_n40790_, new_n40791_,
    new_n40792_, new_n40793_, new_n40794_, new_n40795_, new_n40796_,
    new_n40797_, new_n40798_, new_n40799_, new_n40800_, new_n40801_,
    new_n40802_, new_n40803_, new_n40804_, new_n40805_, new_n40806_,
    new_n40807_, new_n40808_, new_n40809_, new_n40810_, new_n40811_,
    new_n40812_, new_n40813_, new_n40814_, new_n40815_, new_n40816_,
    new_n40817_, new_n40818_, new_n40819_, new_n40820_, new_n40821_,
    new_n40822_, new_n40823_, new_n40824_, new_n40825_, new_n40826_,
    new_n40827_, new_n40828_, new_n40829_, new_n40830_, new_n40831_,
    new_n40832_, new_n40833_, new_n40834_, new_n40835_, new_n40836_,
    new_n40837_, new_n40838_, new_n40839_, new_n40840_, new_n40841_,
    new_n40842_, new_n40843_, new_n40844_, new_n40845_, new_n40846_,
    new_n40847_, new_n40848_, new_n40849_, new_n40850_, new_n40851_,
    new_n40852_, new_n40853_, new_n40854_, new_n40855_, new_n40856_,
    new_n40857_, new_n40859_, new_n40860_, new_n40861_, new_n40862_,
    new_n40863_, new_n40864_, new_n40865_, new_n40866_, new_n40867_,
    new_n40868_, new_n40869_, new_n40870_, new_n40871_, new_n40872_,
    new_n40873_, new_n40874_, new_n40875_, new_n40876_, new_n40877_,
    new_n40878_, new_n40879_, new_n40880_, new_n40881_, new_n40882_,
    new_n40883_, new_n40884_, new_n40885_, new_n40886_, new_n40887_,
    new_n40888_, new_n40889_, new_n40890_, new_n40891_, new_n40892_,
    new_n40893_, new_n40894_, new_n40895_, new_n40896_, new_n40897_,
    new_n40898_, new_n40899_, new_n40900_, new_n40901_, new_n40902_,
    new_n40903_, new_n40904_, new_n40905_, new_n40906_, new_n40907_,
    new_n40908_, new_n40909_, new_n40910_, new_n40911_, new_n40912_,
    new_n40913_, new_n40914_, new_n40915_, new_n40916_, new_n40917_,
    new_n40918_, new_n40919_, new_n40920_, new_n40921_, new_n40922_,
    new_n40923_, new_n40924_, new_n40925_, new_n40926_, new_n40927_,
    new_n40928_, new_n40929_, new_n40930_, new_n40931_, new_n40932_,
    new_n40933_, new_n40934_, new_n40935_, new_n40936_, new_n40937_,
    new_n40938_, new_n40939_, new_n40940_, new_n40941_, new_n40942_,
    new_n40943_, new_n40944_, new_n40945_, new_n40946_, new_n40947_,
    new_n40948_, new_n40949_, new_n40950_, new_n40951_, new_n40952_,
    new_n40953_, new_n40954_, new_n40955_, new_n40956_, new_n40957_,
    new_n40958_, new_n40959_, new_n40960_, new_n40961_, new_n40962_,
    new_n40963_, new_n40964_, new_n40965_, new_n40966_, new_n40967_,
    new_n40968_, new_n40969_, new_n40970_, new_n40971_, new_n40972_,
    new_n40973_, new_n40974_, new_n40975_, new_n40976_, new_n40977_,
    new_n40978_, new_n40979_, new_n40980_, new_n40981_, new_n40982_,
    new_n40983_, new_n40984_, new_n40985_, new_n40986_, new_n40987_,
    new_n40988_, new_n40989_, new_n40990_, new_n40991_, new_n40992_,
    new_n40993_, new_n40994_, new_n40995_, new_n40996_, new_n40997_,
    new_n40998_, new_n40999_, new_n41000_, new_n41001_, new_n41002_,
    new_n41003_, new_n41004_, new_n41005_, new_n41006_, new_n41007_,
    new_n41008_, new_n41009_, new_n41010_, new_n41011_, new_n41012_,
    new_n41013_, new_n41014_, new_n41015_, new_n41016_, new_n41017_,
    new_n41018_, new_n41019_, new_n41020_, new_n41021_, new_n41022_,
    new_n41023_, new_n41024_, new_n41025_, new_n41026_, new_n41027_,
    new_n41028_, new_n41029_, new_n41030_, new_n41031_, new_n41032_,
    new_n41033_, new_n41034_, new_n41035_, new_n41036_, new_n41037_,
    new_n41038_, new_n41039_, new_n41040_, new_n41041_, new_n41042_,
    new_n41043_, new_n41044_, new_n41045_, new_n41046_, new_n41047_,
    new_n41048_, new_n41049_, new_n41050_, new_n41051_, new_n41052_,
    new_n41053_, new_n41054_, new_n41055_, new_n41056_, new_n41057_,
    new_n41058_, new_n41059_, new_n41060_, new_n41061_, new_n41062_,
    new_n41063_, new_n41064_, new_n41065_, new_n41066_, new_n41067_,
    new_n41068_, new_n41069_, new_n41070_, new_n41071_, new_n41072_,
    new_n41073_, new_n41074_, new_n41075_, new_n41076_, new_n41077_,
    new_n41078_, new_n41079_, new_n41080_, new_n41081_, new_n41082_,
    new_n41083_, new_n41084_, new_n41085_, new_n41086_, new_n41087_,
    new_n41088_, new_n41089_, new_n41090_, new_n41091_, new_n41092_,
    new_n41093_, new_n41094_, new_n41095_, new_n41096_, new_n41097_,
    new_n41098_, new_n41099_, new_n41100_, new_n41101_, new_n41102_,
    new_n41103_, new_n41104_, new_n41105_, new_n41106_, new_n41107_,
    new_n41108_, new_n41109_, new_n41110_, new_n41111_, new_n41112_,
    new_n41113_, new_n41114_, new_n41115_, new_n41116_, new_n41117_,
    new_n41118_, new_n41119_, new_n41120_, new_n41121_, new_n41122_,
    new_n41123_, new_n41124_, new_n41125_, new_n41126_, new_n41127_,
    new_n41128_, new_n41129_, new_n41130_, new_n41131_, new_n41132_,
    new_n41133_, new_n41134_, new_n41135_, new_n41136_, new_n41137_,
    new_n41138_, new_n41139_, new_n41140_, new_n41141_, new_n41142_,
    new_n41143_, new_n41144_, new_n41145_, new_n41146_, new_n41147_,
    new_n41148_, new_n41149_, new_n41150_, new_n41151_, new_n41152_,
    new_n41153_, new_n41154_, new_n41155_, new_n41156_, new_n41157_,
    new_n41158_, new_n41159_, new_n41160_, new_n41161_, new_n41162_,
    new_n41163_, new_n41164_, new_n41165_, new_n41166_, new_n41167_,
    new_n41168_, new_n41170_, new_n41171_, new_n41172_, new_n41173_,
    new_n41174_, new_n41175_, new_n41176_, new_n41177_, new_n41178_,
    new_n41179_, new_n41180_, new_n41181_, new_n41182_, new_n41183_,
    new_n41184_, new_n41185_, new_n41186_, new_n41187_, new_n41188_,
    new_n41189_, new_n41190_, new_n41191_, new_n41192_, new_n41193_,
    new_n41194_, new_n41195_, new_n41196_, new_n41197_, new_n41198_,
    new_n41199_, new_n41200_, new_n41201_, new_n41202_, new_n41203_,
    new_n41204_, new_n41205_, new_n41206_, new_n41207_, new_n41208_,
    new_n41209_, new_n41210_, new_n41211_, new_n41212_, new_n41213_,
    new_n41214_, new_n41215_, new_n41216_, new_n41217_, new_n41218_,
    new_n41219_, new_n41220_, new_n41221_, new_n41223_, new_n41224_,
    new_n41225_, new_n41226_, new_n41227_, new_n41228_, new_n41229_,
    new_n41230_, new_n41231_, new_n41232_, new_n41233_, new_n41234_,
    new_n41235_, new_n41236_, new_n41237_, new_n41238_, new_n41239_,
    new_n41240_, new_n41241_, new_n41242_, new_n41243_, new_n41244_,
    new_n41245_, new_n41246_, new_n41247_, new_n41248_, new_n41249_,
    new_n41250_, new_n41251_, new_n41252_, new_n41253_, new_n41254_,
    new_n41255_, new_n41256_, new_n41257_, new_n41258_, new_n41259_,
    new_n41260_, new_n41261_, new_n41262_, new_n41263_, new_n41264_,
    new_n41265_, new_n41266_, new_n41267_, new_n41268_, new_n41269_,
    new_n41270_, new_n41271_, new_n41272_, new_n41273_, new_n41274_,
    new_n41275_, new_n41276_, new_n41277_, new_n41278_, new_n41279_,
    new_n41280_, new_n41281_, new_n41282_, new_n41283_, new_n41284_,
    new_n41285_, new_n41286_, new_n41287_, new_n41288_, new_n41289_,
    new_n41290_, new_n41291_, new_n41292_, new_n41293_, new_n41294_,
    new_n41295_, new_n41296_, new_n41297_, new_n41298_, new_n41299_,
    new_n41300_, new_n41301_, new_n41302_, new_n41303_, new_n41304_,
    new_n41305_, new_n41306_, new_n41307_, new_n41308_, new_n41309_,
    new_n41310_, new_n41311_, new_n41312_, new_n41313_, new_n41314_,
    new_n41315_, new_n41316_, new_n41317_, new_n41318_, new_n41319_,
    new_n41320_, new_n41321_, new_n41322_, new_n41323_, new_n41324_,
    new_n41325_, new_n41326_, new_n41327_, new_n41328_, new_n41329_,
    new_n41330_, new_n41331_, new_n41332_, new_n41333_, new_n41334_,
    new_n41335_, new_n41336_, new_n41337_, new_n41338_, new_n41339_,
    new_n41340_, new_n41341_, new_n41342_, new_n41343_, new_n41344_,
    new_n41345_, new_n41346_, new_n41347_, new_n41348_, new_n41349_,
    new_n41350_, new_n41351_, new_n41352_, new_n41353_, new_n41354_,
    new_n41355_, new_n41356_, new_n41357_, new_n41358_, new_n41359_,
    new_n41360_, new_n41361_, new_n41362_, new_n41363_, new_n41364_,
    new_n41365_, new_n41366_, new_n41367_, new_n41368_, new_n41369_,
    new_n41370_, new_n41371_, new_n41372_, new_n41373_, new_n41374_,
    new_n41375_, new_n41376_, new_n41377_, new_n41378_, new_n41379_,
    new_n41380_, new_n41381_, new_n41382_, new_n41383_, new_n41384_,
    new_n41385_, new_n41386_, new_n41387_, new_n41388_, new_n41389_,
    new_n41390_, new_n41391_, new_n41392_, new_n41393_, new_n41394_,
    new_n41395_, new_n41396_, new_n41397_, new_n41398_, new_n41399_,
    new_n41400_, new_n41401_, new_n41402_, new_n41403_, new_n41404_,
    new_n41405_, new_n41406_, new_n41407_, new_n41408_, new_n41409_,
    new_n41410_, new_n41411_, new_n41412_, new_n41413_, new_n41414_,
    new_n41415_, new_n41416_, new_n41417_, new_n41418_, new_n41419_,
    new_n41420_, new_n41421_, new_n41422_, new_n41423_, new_n41424_,
    new_n41425_, new_n41426_, new_n41427_, new_n41428_, new_n41429_,
    new_n41430_, new_n41431_, new_n41432_, new_n41433_, new_n41434_,
    new_n41435_, new_n41436_, new_n41437_, new_n41438_, new_n41439_,
    new_n41440_, new_n41441_, new_n41442_, new_n41443_, new_n41444_,
    new_n41445_, new_n41446_, new_n41447_, new_n41448_, new_n41449_,
    new_n41450_, new_n41451_, new_n41452_, new_n41453_, new_n41454_,
    new_n41455_, new_n41456_, new_n41457_, new_n41458_, new_n41459_,
    new_n41460_, new_n41461_, new_n41462_, new_n41463_, new_n41464_,
    new_n41465_, new_n41466_, new_n41467_, new_n41468_, new_n41470_,
    new_n41471_, new_n41472_, new_n41473_, new_n41474_, new_n41475_,
    new_n41476_, new_n41477_, new_n41478_, new_n41479_, new_n41480_,
    new_n41481_, new_n41482_, new_n41483_, new_n41484_, new_n41485_,
    new_n41486_, new_n41487_, new_n41488_, new_n41489_, new_n41490_,
    new_n41491_, new_n41492_, new_n41493_, new_n41494_, new_n41495_,
    new_n41496_, new_n41497_, new_n41498_, new_n41499_, new_n41500_,
    new_n41501_, new_n41502_, new_n41503_, new_n41504_, new_n41505_,
    new_n41506_, new_n41507_, new_n41508_, new_n41509_, new_n41510_,
    new_n41511_, new_n41512_, new_n41513_, new_n41514_, new_n41515_,
    new_n41516_, new_n41517_, new_n41518_, new_n41519_, new_n41520_,
    new_n41521_, new_n41522_, new_n41523_, new_n41524_, new_n41525_,
    new_n41526_, new_n41527_, new_n41528_, new_n41529_, new_n41530_,
    new_n41531_, new_n41532_, new_n41533_, new_n41534_, new_n41535_,
    new_n41536_, new_n41537_, new_n41538_, new_n41539_, new_n41540_,
    new_n41541_, new_n41542_, new_n41543_, new_n41544_, new_n41545_,
    new_n41546_, new_n41547_, new_n41548_, new_n41549_, new_n41550_,
    new_n41551_, new_n41552_, new_n41553_, new_n41554_, new_n41555_,
    new_n41556_, new_n41557_, new_n41558_, new_n41559_, new_n41560_,
    new_n41561_, new_n41562_, new_n41563_, new_n41564_, new_n41565_,
    new_n41566_, new_n41567_, new_n41568_, new_n41569_, new_n41570_,
    new_n41571_, new_n41572_, new_n41573_, new_n41574_, new_n41575_,
    new_n41576_, new_n41577_, new_n41578_, new_n41579_, new_n41580_,
    new_n41581_, new_n41582_, new_n41583_, new_n41584_, new_n41585_,
    new_n41586_, new_n41587_, new_n41588_, new_n41589_, new_n41590_,
    new_n41591_, new_n41592_, new_n41593_, new_n41594_, new_n41595_,
    new_n41596_, new_n41597_, new_n41598_, new_n41599_, new_n41600_,
    new_n41601_, new_n41602_, new_n41603_, new_n41604_, new_n41605_,
    new_n41606_, new_n41607_, new_n41608_, new_n41609_, new_n41610_,
    new_n41611_, new_n41612_, new_n41613_, new_n41614_, new_n41615_,
    new_n41616_, new_n41617_, new_n41618_, new_n41619_, new_n41620_,
    new_n41621_, new_n41622_, new_n41623_, new_n41624_, new_n41625_,
    new_n41626_, new_n41627_, new_n41628_, new_n41629_, new_n41630_,
    new_n41631_, new_n41632_, new_n41633_, new_n41634_, new_n41635_,
    new_n41636_, new_n41637_, new_n41638_, new_n41639_, new_n41640_,
    new_n41641_, new_n41642_, new_n41643_, new_n41644_, new_n41645_,
    new_n41646_, new_n41647_, new_n41648_, new_n41649_, new_n41650_,
    new_n41651_, new_n41652_, new_n41653_, new_n41654_, new_n41655_,
    new_n41656_, new_n41657_, new_n41658_, new_n41659_, new_n41660_,
    new_n41661_, new_n41662_, new_n41663_, new_n41664_, new_n41665_,
    new_n41666_, new_n41667_, new_n41668_, new_n41669_, new_n41670_,
    new_n41671_, new_n41672_, new_n41673_, new_n41674_, new_n41675_,
    new_n41676_, new_n41677_, new_n41678_, new_n41679_, new_n41680_,
    new_n41681_, new_n41682_, new_n41683_, new_n41684_, new_n41685_,
    new_n41686_, new_n41687_, new_n41688_, new_n41689_, new_n41690_,
    new_n41691_, new_n41692_, new_n41693_, new_n41694_, new_n41695_,
    new_n41696_, new_n41697_, new_n41698_, new_n41699_, new_n41700_,
    new_n41701_, new_n41702_, new_n41703_, new_n41704_, new_n41705_,
    new_n41706_, new_n41707_, new_n41708_, new_n41709_, new_n41710_,
    new_n41711_, new_n41712_, new_n41713_, new_n41714_, new_n41715_,
    new_n41716_, new_n41717_, new_n41718_, new_n41719_, new_n41720_,
    new_n41721_, new_n41722_, new_n41723_, new_n41724_, new_n41725_,
    new_n41726_, new_n41727_, new_n41728_, new_n41729_, new_n41730_,
    new_n41731_, new_n41732_, new_n41733_, new_n41734_, new_n41735_,
    new_n41736_, new_n41737_, new_n41738_, new_n41739_, new_n41740_,
    new_n41741_, new_n41742_, new_n41744_, new_n41745_, new_n41746_,
    new_n41747_, new_n41748_, new_n41749_, new_n41750_, new_n41751_,
    new_n41752_, new_n41753_, new_n41754_, new_n41755_, new_n41756_,
    new_n41757_, new_n41758_, new_n41759_, new_n41760_, new_n41761_,
    new_n41762_, new_n41763_, new_n41764_, new_n41765_, new_n41766_,
    new_n41767_, new_n41768_, new_n41769_, new_n41770_, new_n41771_,
    new_n41772_, new_n41773_, new_n41774_, new_n41775_, new_n41776_,
    new_n41777_, new_n41778_, new_n41779_, new_n41780_, new_n41781_,
    new_n41782_, new_n41783_, new_n41784_, new_n41785_, new_n41786_,
    new_n41787_, new_n41788_, new_n41789_, new_n41790_, new_n41791_,
    new_n41792_, new_n41793_, new_n41794_, new_n41795_, new_n41796_,
    new_n41797_, new_n41798_, new_n41799_, new_n41800_, new_n41801_,
    new_n41802_, new_n41803_, new_n41804_, new_n41805_, new_n41806_,
    new_n41807_, new_n41808_, new_n41809_, new_n41810_, new_n41811_,
    new_n41812_, new_n41813_, new_n41814_, new_n41815_, new_n41816_,
    new_n41817_, new_n41818_, new_n41819_, new_n41820_, new_n41821_,
    new_n41822_, new_n41823_, new_n41824_, new_n41825_, new_n41826_,
    new_n41827_, new_n41828_, new_n41829_, new_n41830_, new_n41831_,
    new_n41832_, new_n41833_, new_n41834_, new_n41835_, new_n41836_,
    new_n41837_, new_n41838_, new_n41839_, new_n41840_, new_n41841_,
    new_n41842_, new_n41843_, new_n41844_, new_n41845_, new_n41846_,
    new_n41847_, new_n41848_, new_n41849_, new_n41850_, new_n41851_,
    new_n41852_, new_n41853_, new_n41854_, new_n41855_, new_n41856_,
    new_n41857_, new_n41858_, new_n41859_, new_n41860_, new_n41861_,
    new_n41862_, new_n41863_, new_n41864_, new_n41865_, new_n41866_,
    new_n41867_, new_n41868_, new_n41869_, new_n41870_, new_n41871_,
    new_n41872_, new_n41873_, new_n41874_, new_n41875_, new_n41876_,
    new_n41877_, new_n41878_, new_n41879_, new_n41880_, new_n41881_,
    new_n41882_, new_n41883_, new_n41884_, new_n41885_, new_n41886_,
    new_n41887_, new_n41888_, new_n41889_, new_n41890_, new_n41891_,
    new_n41892_, new_n41893_, new_n41894_, new_n41895_, new_n41896_,
    new_n41897_, new_n41898_, new_n41899_, new_n41900_, new_n41901_,
    new_n41902_, new_n41903_, new_n41904_, new_n41905_, new_n41906_,
    new_n41907_, new_n41908_, new_n41909_, new_n41910_, new_n41911_,
    new_n41912_, new_n41913_, new_n41914_, new_n41915_, new_n41916_,
    new_n41917_, new_n41918_, new_n41919_, new_n41920_, new_n41921_,
    new_n41922_, new_n41923_, new_n41924_, new_n41925_, new_n41926_,
    new_n41927_, new_n41928_, new_n41929_, new_n41930_, new_n41931_,
    new_n41932_, new_n41933_, new_n41934_, new_n41935_, new_n41936_,
    new_n41937_, new_n41938_, new_n41939_, new_n41940_, new_n41941_,
    new_n41942_, new_n41943_, new_n41944_, new_n41945_, new_n41946_,
    new_n41947_, new_n41948_, new_n41949_, new_n41950_, new_n41951_,
    new_n41952_, new_n41953_, new_n41954_, new_n41955_, new_n41956_,
    new_n41957_, new_n41958_, new_n41959_, new_n41960_, new_n41961_,
    new_n41962_, new_n41963_, new_n41964_, new_n41965_, new_n41966_,
    new_n41967_, new_n41968_, new_n41969_, new_n41970_, new_n41971_,
    new_n41972_, new_n41974_, new_n41975_, new_n41976_, new_n41977_,
    new_n41978_, new_n41979_, new_n41980_, new_n41981_, new_n41982_,
    new_n41983_, new_n41984_, new_n41985_, new_n41986_, new_n41987_,
    new_n41988_, new_n41989_, new_n41990_, new_n41991_, new_n41992_,
    new_n41993_, new_n41994_, new_n41995_, new_n41996_, new_n41997_,
    new_n41998_, new_n41999_, new_n42000_, new_n42001_, new_n42002_,
    new_n42003_, new_n42004_, new_n42005_, new_n42006_, new_n42007_,
    new_n42008_, new_n42009_, new_n42010_, new_n42011_, new_n42012_,
    new_n42013_, new_n42014_, new_n42015_, new_n42016_, new_n42017_,
    new_n42018_, new_n42019_, new_n42020_, new_n42021_, new_n42022_,
    new_n42023_, new_n42024_, new_n42025_, new_n42026_, new_n42027_,
    new_n42028_, new_n42029_, new_n42030_, new_n42031_, new_n42032_,
    new_n42033_, new_n42034_, new_n42035_, new_n42036_, new_n42037_,
    new_n42038_, new_n42039_, new_n42040_, new_n42041_, new_n42042_,
    new_n42043_, new_n42044_, new_n42045_, new_n42046_, new_n42047_,
    new_n42048_, new_n42049_, new_n42050_, new_n42051_, new_n42052_,
    new_n42053_, new_n42054_, new_n42055_, new_n42056_, new_n42057_,
    new_n42058_, new_n42059_, new_n42060_, new_n42061_, new_n42062_,
    new_n42063_, new_n42064_, new_n42065_, new_n42066_, new_n42067_,
    new_n42068_, new_n42069_, new_n42070_, new_n42071_, new_n42072_,
    new_n42073_, new_n42074_, new_n42075_, new_n42076_, new_n42077_,
    new_n42078_, new_n42079_, new_n42080_, new_n42081_, new_n42082_,
    new_n42083_, new_n42084_, new_n42085_, new_n42086_, new_n42087_,
    new_n42088_, new_n42089_, new_n42090_, new_n42091_, new_n42092_,
    new_n42093_, new_n42094_, new_n42095_, new_n42096_, new_n42097_,
    new_n42098_, new_n42099_, new_n42100_, new_n42101_, new_n42102_,
    new_n42103_, new_n42104_, new_n42105_, new_n42106_, new_n42107_,
    new_n42108_, new_n42109_, new_n42110_, new_n42111_, new_n42112_,
    new_n42113_, new_n42114_, new_n42115_, new_n42116_, new_n42117_,
    new_n42118_, new_n42119_, new_n42120_, new_n42121_, new_n42122_,
    new_n42123_, new_n42124_, new_n42125_, new_n42126_, new_n42127_,
    new_n42128_, new_n42129_, new_n42130_, new_n42131_, new_n42132_,
    new_n42133_, new_n42134_, new_n42135_, new_n42137_, new_n42138_,
    new_n42139_, new_n42140_, new_n42141_, new_n42142_, new_n42143_,
    new_n42144_, new_n42145_, new_n42146_, new_n42147_, new_n42148_,
    new_n42149_, new_n42150_, new_n42151_, new_n42152_, new_n42153_,
    new_n42154_, new_n42155_, new_n42156_, new_n42157_, new_n42158_,
    new_n42159_, new_n42160_, new_n42161_, new_n42162_, new_n42163_,
    new_n42164_, new_n42165_, new_n42166_, new_n42167_, new_n42168_,
    new_n42169_, new_n42170_, new_n42171_, new_n42172_, new_n42173_,
    new_n42174_, new_n42175_, new_n42176_, new_n42177_, new_n42178_,
    new_n42179_, new_n42180_, new_n42181_, new_n42182_, new_n42183_,
    new_n42184_, new_n42185_, new_n42186_, new_n42187_, new_n42188_,
    new_n42189_, new_n42190_, new_n42191_, new_n42192_, new_n42193_,
    new_n42194_, new_n42195_, new_n42196_, new_n42197_, new_n42198_,
    new_n42199_, new_n42200_, new_n42201_, new_n42202_, new_n42203_,
    new_n42204_, new_n42205_, new_n42206_, new_n42207_, new_n42208_,
    new_n42209_, new_n42210_, new_n42211_, new_n42212_, new_n42213_,
    new_n42214_, new_n42215_, new_n42216_, new_n42217_, new_n42218_,
    new_n42219_, new_n42220_, new_n42221_, new_n42222_, new_n42223_,
    new_n42224_, new_n42225_, new_n42226_, new_n42227_, new_n42228_,
    new_n42229_, new_n42230_, new_n42231_, new_n42232_, new_n42233_,
    new_n42234_, new_n42235_, new_n42236_, new_n42237_, new_n42238_,
    new_n42239_, new_n42240_, new_n42241_, new_n42242_, new_n42243_,
    new_n42244_, new_n42245_, new_n42246_, new_n42247_, new_n42248_,
    new_n42249_, new_n42250_, new_n42251_, new_n42252_, new_n42253_,
    new_n42254_, new_n42255_, new_n42256_, new_n42257_, new_n42258_,
    new_n42259_, new_n42260_, new_n42261_, new_n42262_, new_n42263_,
    new_n42264_, new_n42265_, new_n42266_, new_n42267_, new_n42268_,
    new_n42269_, new_n42270_, new_n42271_, new_n42272_, new_n42273_,
    new_n42274_, new_n42275_, new_n42276_, new_n42277_, new_n42278_,
    new_n42279_, new_n42280_, new_n42281_, new_n42282_, new_n42283_,
    new_n42284_, new_n42285_, new_n42286_, new_n42287_, new_n42288_,
    new_n42289_, new_n42290_, new_n42291_, new_n42292_, new_n42293_,
    new_n42294_, new_n42295_, new_n42296_, new_n42297_, new_n42298_,
    new_n42299_, new_n42300_, new_n42301_, new_n42302_, new_n42303_,
    new_n42304_, new_n42305_, new_n42306_, new_n42307_, new_n42308_,
    new_n42309_, new_n42310_, new_n42311_, new_n42312_, new_n42313_,
    new_n42314_, new_n42315_, new_n42316_, new_n42317_, new_n42318_,
    new_n42319_, new_n42320_, new_n42321_, new_n42322_, new_n42323_,
    new_n42325_, new_n42326_, new_n42327_, new_n42328_, new_n42329_,
    new_n42330_, new_n42331_, new_n42333_, new_n42334_, new_n42335_,
    new_n42336_, new_n42337_, new_n42338_, new_n42339_, new_n42340_,
    new_n42341_, new_n42343_, new_n42344_, new_n42345_, new_n42346_,
    new_n42347_, new_n42348_, new_n42349_, new_n42350_, new_n42351_,
    new_n42352_, new_n42353_, new_n42354_, new_n42355_, new_n42356_,
    new_n42357_, new_n42358_, new_n42359_, new_n42360_, new_n42361_,
    new_n42362_, new_n42363_, new_n42364_, new_n42365_, new_n42366_,
    new_n42367_, new_n42368_, new_n42369_, new_n42370_, new_n42371_,
    new_n42372_, new_n42373_, new_n42374_, new_n42375_, new_n42376_,
    new_n42377_, new_n42378_, new_n42379_, new_n42380_, new_n42381_,
    new_n42382_, new_n42383_, new_n42385_, new_n42386_, new_n42387_,
    new_n42388_, new_n42389_, new_n42390_, new_n42391_, new_n42392_,
    new_n42393_, new_n42394_, new_n42395_, new_n42396_, new_n42397_,
    new_n42398_, new_n42399_, new_n42400_, new_n42401_, new_n42402_,
    new_n42403_, new_n42404_, new_n42405_, new_n42406_, new_n42407_,
    new_n42408_, new_n42409_, new_n42410_, new_n42411_, new_n42412_,
    new_n42413_, new_n42414_, new_n42415_, new_n42416_, new_n42417_,
    new_n42418_, new_n42419_, new_n42420_, new_n42421_, new_n42422_,
    new_n42423_, new_n42424_, new_n42425_, new_n42426_, new_n42427_,
    new_n42428_, new_n42429_, new_n42430_, new_n42431_, new_n42432_,
    new_n42433_, new_n42434_, new_n42435_, new_n42436_, new_n42437_,
    new_n42438_, new_n42439_, new_n42440_, new_n42441_, new_n42442_,
    new_n42443_, new_n42444_, new_n42445_, new_n42446_, new_n42447_,
    new_n42448_, new_n42449_, new_n42450_, new_n42451_, new_n42452_,
    new_n42453_, new_n42454_, new_n42455_, new_n42456_, new_n42457_,
    new_n42458_, new_n42459_, new_n42460_, new_n42461_, new_n42462_,
    new_n42463_, new_n42464_, new_n42465_, new_n42466_, new_n42467_,
    new_n42468_, new_n42469_, new_n42470_, new_n42471_, new_n42472_,
    new_n42473_, new_n42474_, new_n42475_, new_n42476_, new_n42477_,
    new_n42478_, new_n42479_, new_n42480_, new_n42481_, new_n42482_,
    new_n42483_, new_n42484_, new_n42485_, new_n42486_, new_n42487_,
    new_n42488_, new_n42489_, new_n42490_, new_n42491_, new_n42492_,
    new_n42493_, new_n42494_, new_n42495_, new_n42496_, new_n42497_,
    new_n42498_, new_n42499_, new_n42500_, new_n42501_, new_n42502_,
    new_n42503_, new_n42504_, new_n42505_, new_n42506_, new_n42507_,
    new_n42508_, new_n42509_, new_n42510_, new_n42511_, new_n42512_,
    new_n42513_, new_n42514_, new_n42515_, new_n42516_, new_n42517_,
    new_n42518_, new_n42519_, new_n42520_, new_n42521_, new_n42522_,
    new_n42523_, new_n42524_, new_n42525_, new_n42526_, new_n42527_,
    new_n42528_, new_n42529_, new_n42530_, new_n42531_, new_n42532_,
    new_n42533_, new_n42534_, new_n42535_, new_n42536_, new_n42537_,
    new_n42538_, new_n42539_, new_n42540_, new_n42541_, new_n42542_,
    new_n42543_, new_n42544_, new_n42545_, new_n42546_, new_n42547_,
    new_n42548_, new_n42549_, new_n42550_, new_n42551_, new_n42552_,
    new_n42553_, new_n42554_, new_n42555_, new_n42556_, new_n42557_,
    new_n42558_, new_n42559_, new_n42560_, new_n42561_, new_n42562_,
    new_n42563_, new_n42564_, new_n42565_, new_n42566_, new_n42567_,
    new_n42568_, new_n42569_, new_n42570_, new_n42571_, new_n42572_,
    new_n42573_, new_n42574_, new_n42575_, new_n42576_, new_n42577_,
    new_n42578_, new_n42579_, new_n42580_, new_n42581_, new_n42582_,
    new_n42583_, new_n42584_, new_n42585_, new_n42586_, new_n42587_,
    new_n42588_, new_n42589_, new_n42590_, new_n42591_, new_n42592_,
    new_n42593_, new_n42594_, new_n42595_, new_n42596_, new_n42597_,
    new_n42598_, new_n42599_, new_n42600_, new_n42601_, new_n42602_,
    new_n42603_, new_n42604_, new_n42605_, new_n42606_, new_n42607_,
    new_n42608_, new_n42609_, new_n42610_, new_n42611_, new_n42612_,
    new_n42613_, new_n42614_, new_n42615_, new_n42616_, new_n42617_,
    new_n42618_, new_n42619_, new_n42621_, new_n42622_, new_n42623_,
    new_n42624_, new_n42625_, new_n42626_, new_n42627_, new_n42628_,
    new_n42629_, new_n42630_, new_n42631_, new_n42632_, new_n42633_,
    new_n42634_, new_n42635_, new_n42636_, new_n42637_, new_n42638_,
    new_n42639_, new_n42640_, new_n42641_, new_n42642_, new_n42643_,
    new_n42644_, new_n42645_, new_n42646_, new_n42647_, new_n42648_,
    new_n42649_, new_n42650_, new_n42651_, new_n42652_, new_n42653_,
    new_n42654_, new_n42655_, new_n42656_, new_n42657_, new_n42658_,
    new_n42659_, new_n42660_, new_n42661_, new_n42662_, new_n42663_,
    new_n42664_, new_n42665_, new_n42666_, new_n42667_, new_n42668_,
    new_n42669_, new_n42670_, new_n42671_, new_n42672_, new_n42673_,
    new_n42674_, new_n42675_, new_n42676_, new_n42677_, new_n42678_,
    new_n42679_, new_n42680_, new_n42681_, new_n42682_, new_n42683_,
    new_n42684_, new_n42685_, new_n42686_, new_n42687_, new_n42688_,
    new_n42689_, new_n42690_, new_n42691_, new_n42692_, new_n42693_,
    new_n42694_, new_n42695_, new_n42696_, new_n42697_, new_n42698_,
    new_n42699_, new_n42700_, new_n42701_, new_n42702_, new_n42703_,
    new_n42704_, new_n42705_, new_n42706_, new_n42707_, new_n42708_,
    new_n42709_, new_n42710_, new_n42711_, new_n42712_, new_n42713_,
    new_n42714_, new_n42715_, new_n42716_, new_n42717_, new_n42718_,
    new_n42719_, new_n42720_, new_n42721_, new_n42722_, new_n42723_,
    new_n42724_, new_n42725_, new_n42726_, new_n42727_, new_n42728_,
    new_n42729_, new_n42730_, new_n42731_, new_n42732_, new_n42733_,
    new_n42734_, new_n42735_, new_n42736_, new_n42737_, new_n42738_,
    new_n42739_, new_n42740_, new_n42741_, new_n42742_, new_n42743_,
    new_n42744_, new_n42745_, new_n42746_, new_n42747_, new_n42748_,
    new_n42749_, new_n42750_, new_n42751_, new_n42752_, new_n42753_,
    new_n42754_, new_n42755_, new_n42756_, new_n42757_, new_n42758_,
    new_n42759_, new_n42760_, new_n42761_, new_n42762_, new_n42763_,
    new_n42764_, new_n42765_, new_n42766_, new_n42767_, new_n42768_,
    new_n42769_, new_n42770_, new_n42771_, new_n42772_, new_n42773_,
    new_n42774_, new_n42775_, new_n42776_, new_n42777_, new_n42778_,
    new_n42779_, new_n42780_, new_n42781_, new_n42782_, new_n42783_,
    new_n42784_, new_n42785_, new_n42786_, new_n42787_, new_n42788_,
    new_n42789_, new_n42790_, new_n42791_, new_n42792_, new_n42793_,
    new_n42794_, new_n42795_, new_n42796_, new_n42797_, new_n42798_,
    new_n42799_, new_n42800_, new_n42801_, new_n42802_, new_n42803_,
    new_n42804_, new_n42805_, new_n42806_, new_n42807_, new_n42808_,
    new_n42809_, new_n42810_, new_n42811_, new_n42812_, new_n42813_,
    new_n42814_, new_n42815_, new_n42816_, new_n42817_, new_n42818_,
    new_n42819_, new_n42820_, new_n42821_, new_n42822_, new_n42823_,
    new_n42824_, new_n42825_, new_n42826_, new_n42827_, new_n42828_,
    new_n42829_, new_n42830_, new_n42831_, new_n42832_, new_n42833_,
    new_n42834_, new_n42835_, new_n42836_, new_n42837_, new_n42838_,
    new_n42839_, new_n42840_, new_n42841_, new_n42842_, new_n42843_,
    new_n42844_, new_n42845_, new_n42847_, new_n42848_, new_n42849_,
    new_n42850_, new_n42851_, new_n42853_, new_n42854_, new_n42855_,
    new_n42856_, new_n42857_, new_n42859_, new_n42860_, new_n42861_,
    new_n42862_, new_n42863_, new_n42865_, new_n42866_, new_n42867_,
    new_n42868_, new_n42869_, new_n42871_, new_n42872_, new_n42873_,
    new_n42874_, new_n42875_, new_n42877_, new_n42878_, new_n42879_,
    new_n42880_, new_n42881_, new_n42882_, new_n42884_, new_n42885_,
    new_n42886_, new_n42887_, new_n42888_, new_n42889_, new_n42891_,
    new_n42892_, new_n42893_, new_n42894_, new_n42895_, new_n42896_,
    new_n42897_, new_n42898_, new_n42899_, new_n42900_, new_n42901_,
    new_n42902_, new_n42903_, new_n42904_, new_n42905_, new_n42906_,
    new_n42907_, new_n42908_, new_n42909_, new_n42910_, new_n42911_,
    new_n42912_, new_n42913_, new_n42914_, new_n42915_, new_n42916_,
    new_n42917_, new_n42918_, new_n42919_, new_n42920_, new_n42921_,
    new_n42922_, new_n42923_, new_n42925_, new_n42926_, new_n42927_,
    new_n42928_, new_n42929_, new_n42930_, new_n42931_, new_n42932_,
    new_n42933_, new_n42934_, new_n42935_, new_n42936_, new_n42937_,
    new_n42938_, new_n42939_, new_n42940_, new_n42941_, new_n42942_,
    new_n42943_, new_n42944_, new_n42945_, new_n42946_, new_n42947_,
    new_n42948_, new_n42949_, new_n42950_, new_n42951_, new_n42952_,
    new_n42953_, new_n42954_, new_n42955_, new_n42956_, new_n42957_,
    new_n42958_, new_n42959_, new_n42960_, new_n42961_, new_n42962_,
    new_n42963_, new_n42964_, new_n42965_, new_n42966_, new_n42967_,
    new_n42968_, new_n42969_, new_n42970_, new_n42971_, new_n42972_,
    new_n42973_, new_n42974_, new_n42975_, new_n42976_, new_n42977_,
    new_n42978_, new_n42979_, new_n42980_, new_n42981_, new_n42982_,
    new_n42983_, new_n42984_, new_n42985_, new_n42986_, new_n42987_,
    new_n42988_, new_n42989_, new_n42990_, new_n42991_, new_n42992_,
    new_n42993_, new_n42994_, new_n42995_, new_n42996_, new_n42997_,
    new_n42998_, new_n42999_, new_n43000_, new_n43001_, new_n43002_,
    new_n43003_, new_n43004_, new_n43005_, new_n43006_, new_n43007_,
    new_n43008_, new_n43009_, new_n43010_, new_n43011_, new_n43012_,
    new_n43013_, new_n43014_, new_n43015_, new_n43016_, new_n43017_,
    new_n43018_, new_n43019_, new_n43020_, new_n43021_, new_n43022_,
    new_n43023_, new_n43024_, new_n43025_, new_n43026_, new_n43027_,
    new_n43028_, new_n43029_, new_n43030_, new_n43031_, new_n43032_,
    new_n43033_, new_n43034_, new_n43035_, new_n43036_, new_n43037_,
    new_n43038_, new_n43039_, new_n43040_, new_n43041_, new_n43042_,
    new_n43043_, new_n43044_, new_n43045_, new_n43046_, new_n43047_,
    new_n43048_, new_n43049_, new_n43050_, new_n43051_, new_n43052_,
    new_n43053_, new_n43054_, new_n43055_, new_n43056_, new_n43057_,
    new_n43058_, new_n43059_, new_n43060_, new_n43061_, new_n43062_,
    new_n43063_, new_n43064_, new_n43065_, new_n43066_, new_n43067_,
    new_n43068_, new_n43069_, new_n43070_, new_n43071_, new_n43072_,
    new_n43073_, new_n43074_, new_n43075_, new_n43076_, new_n43077_,
    new_n43078_, new_n43079_, new_n43080_, new_n43081_, new_n43082_,
    new_n43083_, new_n43084_, new_n43085_, new_n43086_, new_n43087_,
    new_n43088_, new_n43089_, new_n43090_, new_n43091_, new_n43092_,
    new_n43093_, new_n43094_, new_n43095_, new_n43096_, new_n43097_,
    new_n43098_, new_n43099_, new_n43100_, new_n43101_, new_n43102_,
    new_n43103_, new_n43104_, new_n43105_, new_n43106_, new_n43107_,
    new_n43108_, new_n43109_, new_n43110_, new_n43111_, new_n43112_,
    new_n43113_, new_n43114_, new_n43115_, new_n43116_, new_n43117_,
    new_n43118_, new_n43119_, new_n43120_, new_n43121_, new_n43122_,
    new_n43123_, new_n43124_, new_n43125_, new_n43126_, new_n43127_,
    new_n43128_, new_n43129_, new_n43130_, new_n43131_, new_n43132_,
    new_n43133_, new_n43135_, new_n43136_, new_n43137_, new_n43138_,
    new_n43139_, new_n43140_, new_n43141_, new_n43142_, new_n43143_,
    new_n43144_, new_n43145_, new_n43146_, new_n43147_, new_n43148_,
    new_n43149_, new_n43150_, new_n43151_, new_n43152_, new_n43153_,
    new_n43154_, new_n43155_, new_n43156_, new_n43157_, new_n43158_,
    new_n43159_, new_n43160_, new_n43161_, new_n43162_, new_n43163_,
    new_n43164_, new_n43165_, new_n43166_, new_n43167_, new_n43168_,
    new_n43169_, new_n43170_, new_n43171_, new_n43172_, new_n43173_,
    new_n43174_, new_n43175_, new_n43176_, new_n43177_, new_n43178_,
    new_n43180_, new_n43181_, new_n43182_, new_n43183_, new_n43184_,
    new_n43185_, new_n43186_, new_n43187_, new_n43188_, new_n43189_,
    new_n43190_, new_n43191_, new_n43192_, new_n43193_, new_n43194_,
    new_n43195_, new_n43196_, new_n43197_, new_n43198_, new_n43199_,
    new_n43200_, new_n43201_, new_n43202_, new_n43203_, new_n43204_,
    new_n43205_, new_n43206_, new_n43207_, new_n43208_, new_n43209_,
    new_n43210_, new_n43211_, new_n43212_, new_n43213_, new_n43214_,
    new_n43215_, new_n43216_, new_n43217_, new_n43218_, new_n43219_,
    new_n43221_, new_n43222_, new_n43223_, new_n43224_, new_n43225_,
    new_n43226_, new_n43227_, new_n43228_, new_n43229_, new_n43230_,
    new_n43231_, new_n43232_, new_n43233_, new_n43234_, new_n43235_,
    new_n43236_, new_n43237_, new_n43238_, new_n43239_, new_n43240_,
    new_n43241_, new_n43242_, new_n43243_, new_n43244_, new_n43245_,
    new_n43246_, new_n43247_, new_n43248_, new_n43249_, new_n43250_,
    new_n43251_, new_n43252_, new_n43253_, new_n43254_, new_n43255_,
    new_n43256_, new_n43257_, new_n43258_, new_n43259_, new_n43260_,
    new_n43261_, new_n43262_, new_n43263_, new_n43264_, new_n43265_,
    new_n43266_, new_n43267_, new_n43268_, new_n43269_, new_n43270_,
    new_n43271_, new_n43272_, new_n43273_, new_n43274_, new_n43275_,
    new_n43276_, new_n43277_, new_n43278_, new_n43279_, new_n43280_,
    new_n43281_, new_n43282_, new_n43283_, new_n43284_, new_n43285_,
    new_n43286_, new_n43288_, new_n43289_, new_n43290_, new_n43291_,
    new_n43292_, new_n43293_, new_n43294_, new_n43295_, new_n43296_,
    new_n43297_, new_n43298_, new_n43299_, new_n43300_, new_n43301_,
    new_n43302_, new_n43303_, new_n43304_, new_n43305_, new_n43306_,
    new_n43307_, new_n43308_, new_n43309_, new_n43310_, new_n43311_,
    new_n43312_, new_n43313_, new_n43314_, new_n43315_, new_n43316_,
    new_n43317_, new_n43318_, new_n43319_, new_n43320_, new_n43321_,
    new_n43322_, new_n43323_, new_n43324_, new_n43325_, new_n43326_,
    new_n43327_, new_n43328_, new_n43329_, new_n43330_, new_n43331_,
    new_n43332_, new_n43333_, new_n43334_, new_n43335_, new_n43336_,
    new_n43337_, new_n43338_, new_n43339_, new_n43340_, new_n43341_,
    new_n43342_, new_n43343_, new_n43344_, new_n43345_, new_n43346_,
    new_n43347_, new_n43348_, new_n43349_, new_n43350_, new_n43351_,
    new_n43352_, new_n43353_, new_n43354_, new_n43355_, new_n43356_,
    new_n43357_, new_n43358_, new_n43359_, new_n43360_, new_n43361_,
    new_n43362_, new_n43363_, new_n43364_, new_n43365_, new_n43366_,
    new_n43367_, new_n43368_, new_n43369_, new_n43370_, new_n43371_,
    new_n43372_, new_n43373_, new_n43374_, new_n43375_, new_n43376_,
    new_n43377_, new_n43378_, new_n43379_, new_n43380_, new_n43381_,
    new_n43382_, new_n43383_, new_n43384_, new_n43385_, new_n43386_,
    new_n43387_, new_n43388_, new_n43389_, new_n43390_, new_n43391_,
    new_n43392_, new_n43393_, new_n43394_, new_n43395_, new_n43396_,
    new_n43397_, new_n43398_, new_n43399_, new_n43400_, new_n43401_,
    new_n43402_, new_n43403_, new_n43404_, new_n43405_, new_n43406_,
    new_n43407_, new_n43408_, new_n43409_, new_n43410_, new_n43411_,
    new_n43412_, new_n43413_, new_n43414_, new_n43415_, new_n43416_,
    new_n43417_, new_n43418_, new_n43419_, new_n43420_, new_n43421_,
    new_n43422_, new_n43423_, new_n43424_, new_n43425_, new_n43426_,
    new_n43427_, new_n43428_, new_n43429_, new_n43430_, new_n43431_,
    new_n43432_, new_n43433_, new_n43434_, new_n43435_, new_n43436_,
    new_n43437_, new_n43438_, new_n43439_, new_n43440_, new_n43441_,
    new_n43442_, new_n43443_, new_n43444_, new_n43445_, new_n43446_,
    new_n43447_, new_n43448_, new_n43449_, new_n43450_, new_n43451_,
    new_n43452_, new_n43453_, new_n43454_, new_n43455_, new_n43456_,
    new_n43457_, new_n43458_, new_n43459_, new_n43460_, new_n43461_,
    new_n43462_, new_n43463_, new_n43464_, new_n43465_, new_n43466_,
    new_n43467_, new_n43468_, new_n43469_, new_n43470_, new_n43471_,
    new_n43472_, new_n43473_, new_n43474_, new_n43475_, new_n43476_,
    new_n43477_, new_n43478_, new_n43479_, new_n43480_, new_n43481_,
    new_n43482_, new_n43483_, new_n43484_, new_n43485_, new_n43486_,
    new_n43487_, new_n43488_, new_n43489_, new_n43490_, new_n43491_,
    new_n43492_, new_n43493_, new_n43495_, new_n43496_, new_n43497_,
    new_n43498_, new_n43499_, new_n43500_, new_n43501_, new_n43502_,
    new_n43503_, new_n43504_, new_n43505_, new_n43506_, new_n43507_,
    new_n43508_, new_n43509_, new_n43510_, new_n43511_, new_n43512_,
    new_n43513_, new_n43514_, new_n43515_, new_n43516_, new_n43517_,
    new_n43518_, new_n43519_, new_n43520_, new_n43521_, new_n43522_,
    new_n43523_, new_n43524_, new_n43525_, new_n43526_, new_n43527_,
    new_n43528_, new_n43529_, new_n43530_, new_n43531_, new_n43532_,
    new_n43533_, new_n43534_, new_n43535_, new_n43536_, new_n43537_,
    new_n43538_, new_n43539_, new_n43540_, new_n43541_, new_n43542_,
    new_n43543_, new_n43544_, new_n43545_, new_n43546_, new_n43547_,
    new_n43548_, new_n43549_, new_n43550_, new_n43551_, new_n43552_,
    new_n43553_, new_n43554_, new_n43555_, new_n43556_, new_n43557_,
    new_n43558_, new_n43559_, new_n43560_, new_n43561_, new_n43562_,
    new_n43563_, new_n43564_, new_n43565_, new_n43566_, new_n43567_,
    new_n43568_, new_n43569_, new_n43570_, new_n43571_, new_n43572_,
    new_n43573_, new_n43574_, new_n43575_, new_n43576_, new_n43577_,
    new_n43578_, new_n43579_, new_n43580_, new_n43581_, new_n43582_,
    new_n43583_, new_n43584_, new_n43585_, new_n43586_, new_n43587_,
    new_n43588_, new_n43589_, new_n43590_, new_n43591_, new_n43592_,
    new_n43593_, new_n43594_, new_n43595_, new_n43596_, new_n43597_,
    new_n43598_, new_n43599_, new_n43600_, new_n43601_, new_n43602_,
    new_n43603_, new_n43604_, new_n43605_, new_n43606_, new_n43607_,
    new_n43608_, new_n43609_, new_n43610_, new_n43611_, new_n43612_,
    new_n43613_, new_n43614_, new_n43615_, new_n43616_, new_n43617_,
    new_n43618_, new_n43619_, new_n43620_, new_n43621_, new_n43622_,
    new_n43623_, new_n43624_, new_n43625_, new_n43626_, new_n43627_,
    new_n43628_, new_n43629_, new_n43630_, new_n43631_, new_n43632_,
    new_n43633_, new_n43634_, new_n43635_, new_n43636_, new_n43637_,
    new_n43638_, new_n43639_, new_n43640_, new_n43641_, new_n43642_,
    new_n43643_, new_n43644_, new_n43645_, new_n43646_, new_n43647_,
    new_n43648_, new_n43649_, new_n43650_, new_n43652_, new_n43653_,
    new_n43654_, new_n43655_, new_n43656_, new_n43657_, new_n43658_,
    new_n43659_, new_n43660_, new_n43661_, new_n43662_, new_n43663_,
    new_n43664_, new_n43665_, new_n43666_, new_n43667_, new_n43668_,
    new_n43669_, new_n43670_, new_n43671_, new_n43672_, new_n43673_,
    new_n43674_, new_n43675_, new_n43676_, new_n43677_, new_n43678_,
    new_n43679_, new_n43680_, new_n43681_, new_n43682_, new_n43683_,
    new_n43684_, new_n43685_, new_n43686_, new_n43687_, new_n43688_,
    new_n43689_, new_n43690_, new_n43691_, new_n43692_, new_n43693_,
    new_n43694_, new_n43695_, new_n43697_, new_n43698_, new_n43699_,
    new_n43700_, new_n43701_, new_n43702_, new_n43703_, new_n43704_,
    new_n43705_, new_n43706_, new_n43707_, new_n43708_, new_n43709_,
    new_n43710_, new_n43711_, new_n43712_, new_n43713_, new_n43714_,
    new_n43715_, new_n43716_, new_n43717_, new_n43718_, new_n43719_,
    new_n43720_, new_n43721_, new_n43722_, new_n43723_, new_n43724_,
    new_n43725_, new_n43726_, new_n43727_, new_n43728_, new_n43729_,
    new_n43730_, new_n43731_, new_n43732_, new_n43733_, new_n43734_,
    new_n43735_, new_n43736_, new_n43737_, new_n43738_, new_n43739_,
    new_n43741_, new_n43742_, new_n43743_, new_n43744_, new_n43745_,
    new_n43746_, new_n43747_, new_n43748_, new_n43749_, new_n43750_,
    new_n43751_, new_n43752_, new_n43753_, new_n43754_, new_n43755_,
    new_n43756_, new_n43757_, new_n43758_, new_n43759_, new_n43760_,
    new_n43761_, new_n43762_, new_n43763_, new_n43764_, new_n43765_,
    new_n43766_, new_n43767_, new_n43768_, new_n43769_, new_n43770_,
    new_n43771_, new_n43772_, new_n43773_, new_n43774_, new_n43775_,
    new_n43776_, new_n43777_, new_n43778_, new_n43779_, new_n43780_,
    new_n43781_, new_n43782_, new_n43783_, new_n43784_, new_n43785_,
    new_n43786_, new_n43787_, new_n43788_, new_n43790_, new_n43791_,
    new_n43792_, new_n43793_, new_n43794_, new_n43795_, new_n43796_,
    new_n43797_, new_n43798_, new_n43799_, new_n43800_, new_n43801_,
    new_n43802_, new_n43803_, new_n43804_, new_n43805_, new_n43806_,
    new_n43807_, new_n43808_, new_n43809_, new_n43810_, new_n43811_,
    new_n43812_, new_n43813_, new_n43814_, new_n43815_, new_n43816_,
    new_n43817_, new_n43818_, new_n43819_, new_n43820_, new_n43821_,
    new_n43822_, new_n43823_, new_n43824_, new_n43825_, new_n43826_,
    new_n43827_, new_n43828_, new_n43829_, new_n43830_, new_n43831_,
    new_n43832_, new_n43833_, new_n43834_, new_n43835_, new_n43836_,
    new_n43837_, new_n43838_, new_n43839_, new_n43840_, new_n43841_,
    new_n43842_, new_n43843_, new_n43844_, new_n43845_, new_n43846_,
    new_n43847_, new_n43848_, new_n43849_, new_n43850_, new_n43851_,
    new_n43852_, new_n43853_, new_n43854_, new_n43855_, new_n43856_,
    new_n43857_, new_n43858_, new_n43859_, new_n43860_, new_n43861_,
    new_n43862_, new_n43863_, new_n43864_, new_n43865_, new_n43866_,
    new_n43867_, new_n43868_, new_n43869_, new_n43870_, new_n43871_,
    new_n43872_, new_n43873_, new_n43874_, new_n43875_, new_n43876_,
    new_n43877_, new_n43878_, new_n43879_, new_n43880_, new_n43881_,
    new_n43882_, new_n43883_, new_n43884_, new_n43885_, new_n43886_,
    new_n43887_, new_n43888_, new_n43889_, new_n43891_, new_n43892_,
    new_n43893_, new_n43894_, new_n43895_, new_n43896_, new_n43897_,
    new_n43898_, new_n43899_, new_n43900_, new_n43901_, new_n43902_,
    new_n43903_, new_n43904_, new_n43905_, new_n43906_, new_n43907_,
    new_n43908_, new_n43909_, new_n43910_, new_n43911_, new_n43912_,
    new_n43913_, new_n43914_, new_n43915_, new_n43916_, new_n43917_,
    new_n43918_, new_n43919_, new_n43920_, new_n43921_, new_n43922_,
    new_n43923_, new_n43924_, new_n43925_, new_n43926_, new_n43927_,
    new_n43928_, new_n43929_, new_n43930_, new_n43931_, new_n43932_,
    new_n43933_, new_n43934_, new_n43935_, new_n43936_, new_n43937_,
    new_n43938_, new_n43939_, new_n43940_, new_n43941_, new_n43942_,
    new_n43943_, new_n43944_, new_n43945_, new_n43946_, new_n43947_,
    new_n43948_, new_n43949_, new_n43950_, new_n43951_, new_n43952_,
    new_n43954_, new_n43955_, new_n43956_, new_n43957_, new_n43958_,
    new_n43959_, new_n43960_, new_n43961_, new_n43962_, new_n43963_,
    new_n43964_, new_n43965_, new_n43966_, new_n43967_, new_n43968_,
    new_n43969_, new_n43970_, new_n43971_, new_n43972_, new_n43973_,
    new_n43974_, new_n43975_, new_n43976_, new_n43977_, new_n43978_,
    new_n43979_, new_n43980_, new_n43981_, new_n43982_, new_n43983_,
    new_n43984_, new_n43985_, new_n43986_, new_n43987_, new_n43988_,
    new_n43989_, new_n43990_, new_n43991_, new_n43992_, new_n43993_,
    new_n43995_, new_n43996_, new_n43997_, new_n43998_, new_n43999_,
    new_n44000_, new_n44001_, new_n44002_, new_n44003_, new_n44004_,
    new_n44005_, new_n44006_, new_n44007_, new_n44008_, new_n44009_,
    new_n44010_, new_n44011_, new_n44012_, new_n44013_, new_n44014_,
    new_n44015_, new_n44016_, new_n44017_, new_n44018_, new_n44019_,
    new_n44020_, new_n44021_, new_n44022_, new_n44023_, new_n44024_,
    new_n44025_, new_n44026_, new_n44027_, new_n44028_, new_n44029_,
    new_n44030_, new_n44031_, new_n44032_, new_n44033_, new_n44034_,
    new_n44035_, new_n44036_, new_n44037_, new_n44038_, new_n44039_,
    new_n44040_, new_n44041_, new_n44042_, new_n44043_, new_n44044_,
    new_n44045_, new_n44046_, new_n44047_, new_n44048_, new_n44049_,
    new_n44050_, new_n44051_, new_n44052_, new_n44053_, new_n44054_,
    new_n44055_, new_n44056_, new_n44057_, new_n44058_, new_n44059_,
    new_n44060_, new_n44061_, new_n44062_, new_n44063_, new_n44064_,
    new_n44065_, new_n44066_, new_n44067_, new_n44069_, new_n44070_,
    new_n44071_, new_n44072_, new_n44073_, new_n44074_, new_n44075_,
    new_n44076_, new_n44077_, new_n44078_, new_n44079_, new_n44080_,
    new_n44081_, new_n44082_, new_n44083_, new_n44084_, new_n44085_,
    new_n44086_, new_n44087_, new_n44088_, new_n44089_, new_n44090_,
    new_n44091_, new_n44092_, new_n44093_, new_n44094_, new_n44095_,
    new_n44096_, new_n44098_, new_n44099_, new_n44100_, new_n44101_,
    new_n44102_, new_n44103_, new_n44104_, new_n44105_, new_n44106_,
    new_n44107_, new_n44108_, new_n44109_, new_n44110_, new_n44111_,
    new_n44112_, new_n44113_, new_n44114_, new_n44115_, new_n44116_,
    new_n44117_, new_n44118_, new_n44119_, new_n44120_, new_n44121_,
    new_n44122_, new_n44123_, new_n44124_, new_n44125_, new_n44126_,
    new_n44127_, new_n44128_, new_n44129_, new_n44130_, new_n44131_,
    new_n44132_, new_n44133_, new_n44134_, new_n44135_, new_n44136_,
    new_n44137_, new_n44138_, new_n44139_, new_n44141_, new_n44142_,
    new_n44143_, new_n44144_, new_n44145_, new_n44146_, new_n44147_,
    new_n44148_, new_n44149_, new_n44150_, new_n44151_, new_n44152_,
    new_n44153_, new_n44154_, new_n44155_, new_n44156_, new_n44157_,
    new_n44158_, new_n44159_, new_n44160_, new_n44161_, new_n44162_,
    new_n44163_, new_n44164_, new_n44165_, new_n44166_, new_n44167_,
    new_n44168_, new_n44169_, new_n44170_, new_n44171_, new_n44172_,
    new_n44173_, new_n44174_, new_n44175_, new_n44176_, new_n44177_,
    new_n44178_, new_n44179_, new_n44180_, new_n44181_, new_n44182_,
    new_n44183_, new_n44184_, new_n44185_, new_n44186_, new_n44187_,
    new_n44188_, new_n44189_, new_n44190_, new_n44191_, new_n44192_,
    new_n44193_, new_n44194_, new_n44195_, new_n44196_, new_n44197_,
    new_n44198_, new_n44199_, new_n44200_, new_n44201_, new_n44202_,
    new_n44203_, new_n44204_, new_n44205_, new_n44206_, new_n44207_,
    new_n44208_, new_n44210_, new_n44211_, new_n44212_, new_n44213_,
    new_n44214_, new_n44215_, new_n44216_, new_n44217_, new_n44218_,
    new_n44219_, new_n44220_, new_n44221_, new_n44222_, new_n44223_,
    new_n44224_, new_n44225_, new_n44226_, new_n44227_, new_n44228_,
    new_n44229_, new_n44230_, new_n44231_, new_n44232_, new_n44233_,
    new_n44234_, new_n44235_, new_n44236_, new_n44237_, new_n44238_,
    new_n44239_, new_n44240_, new_n44241_, new_n44242_, new_n44243_,
    new_n44244_, new_n44245_, new_n44246_, new_n44247_, new_n44248_,
    new_n44249_, new_n44250_, new_n44251_, new_n44252_, new_n44253_,
    new_n44254_, new_n44255_, new_n44256_, new_n44257_, new_n44258_,
    new_n44259_, new_n44260_, new_n44261_, new_n44262_, new_n44263_,
    new_n44264_, new_n44265_, new_n44266_, new_n44267_, new_n44269_,
    new_n44270_, new_n44271_, new_n44272_, new_n44273_, new_n44274_,
    new_n44275_, new_n44276_, new_n44277_, new_n44278_, new_n44279_,
    new_n44280_, new_n44281_, new_n44282_, new_n44283_, new_n44284_,
    new_n44285_, new_n44286_, new_n44287_, new_n44288_, new_n44289_,
    new_n44290_, new_n44291_, new_n44292_, new_n44293_, new_n44294_,
    new_n44295_, new_n44296_, new_n44297_, new_n44298_, new_n44299_,
    new_n44300_, new_n44301_, new_n44302_, new_n44303_, new_n44304_,
    new_n44305_, new_n44306_, new_n44307_, new_n44308_, new_n44309_,
    new_n44310_, new_n44311_, new_n44313_, new_n44314_, new_n44315_,
    new_n44316_, new_n44317_, new_n44318_, new_n44319_, new_n44320_,
    new_n44321_, new_n44322_, new_n44323_, new_n44324_, new_n44325_,
    new_n44326_, new_n44327_, new_n44328_, new_n44329_, new_n44330_,
    new_n44331_, new_n44332_, new_n44333_, new_n44334_, new_n44335_,
    new_n44336_, new_n44337_, new_n44338_, new_n44339_, new_n44340_,
    new_n44341_, new_n44342_, new_n44343_, new_n44344_, new_n44345_,
    new_n44346_, new_n44347_, new_n44348_, new_n44349_, new_n44350_,
    new_n44352_, new_n44353_, new_n44354_, new_n44355_, new_n44356_,
    new_n44357_, new_n44358_, new_n44359_, new_n44360_, new_n44361_,
    new_n44362_, new_n44363_, new_n44364_, new_n44365_, new_n44366_,
    new_n44367_, new_n44368_, new_n44369_, new_n44370_, new_n44371_,
    new_n44372_, new_n44373_, new_n44374_, new_n44375_, new_n44376_,
    new_n44377_, new_n44378_, new_n44379_, new_n44380_, new_n44381_,
    new_n44382_, new_n44383_, new_n44384_, new_n44385_, new_n44386_,
    new_n44387_, new_n44388_, new_n44389_, new_n44391_, new_n44392_,
    new_n44393_, new_n44394_, new_n44395_, new_n44396_, new_n44397_,
    new_n44398_, new_n44399_, new_n44400_, new_n44401_, new_n44402_,
    new_n44403_, new_n44404_, new_n44405_, new_n44406_, new_n44407_,
    new_n44408_, new_n44409_, new_n44410_, new_n44411_, new_n44412_,
    new_n44413_, new_n44414_, new_n44415_, new_n44416_, new_n44417_,
    new_n44418_, new_n44419_, new_n44420_, new_n44421_, new_n44422_,
    new_n44423_, new_n44424_, new_n44425_, new_n44426_, new_n44427_,
    new_n44428_, new_n44429_, new_n44430_, new_n44431_, new_n44432_,
    new_n44433_, new_n44434_, new_n44435_, new_n44436_, new_n44437_,
    new_n44438_, new_n44439_, new_n44440_, new_n44441_, new_n44442_,
    new_n44443_, new_n44444_, new_n44445_, new_n44446_, new_n44447_,
    new_n44448_, new_n44450_, new_n44451_, new_n44452_, new_n44454_,
    new_n44455_, new_n44456_, new_n44457_, new_n44458_, new_n44459_,
    new_n44460_, new_n44461_, new_n44462_, new_n44463_, new_n44464_,
    new_n44465_, new_n44466_, new_n44467_, new_n44468_, new_n44469_,
    new_n44470_, new_n44472_, new_n44473_, new_n44474_, new_n44475_,
    new_n44476_, new_n44477_, new_n44478_, new_n44479_, new_n44480_,
    new_n44481_, new_n44482_, new_n44483_, new_n44484_, new_n44485_,
    new_n44486_, new_n44487_, new_n44488_, new_n44490_, new_n44492_,
    new_n44493_, new_n44495_, new_n44496_, new_n44497_, new_n44499_,
    new_n44500_, new_n44501_, new_n44502_, new_n44503_, new_n44504_,
    new_n44505_, new_n44506_, new_n44507_, new_n44508_, new_n44509_,
    new_n44510_, new_n44511_, new_n44512_, new_n44514_, new_n44515_,
    new_n44517_, new_n44518_, new_n44520_, new_n44521_, new_n44523_,
    new_n44524_, new_n44526_, new_n44527_, new_n44529_, new_n44530_,
    new_n44532_, new_n44533_, new_n44535_, new_n44536_, new_n44538_,
    new_n44539_, new_n44541_, new_n44542_, new_n44543_, new_n44544_,
    new_n44545_, new_n44546_, new_n44547_, new_n44549_, new_n44550_,
    new_n44551_, new_n44552_, new_n44553_, new_n44554_, new_n44556_,
    new_n44557_, new_n44558_, new_n44560_, new_n44561_, new_n44562_,
    new_n44563_, new_n44564_, new_n44565_, new_n44566_, new_n44567_,
    new_n44568_, new_n44569_, new_n44570_, new_n44571_, new_n44572_,
    new_n44573_, new_n44574_, new_n44575_, new_n44576_, new_n44577_,
    new_n44578_, new_n44579_, new_n44580_, new_n44582_, new_n44583_,
    new_n44585_, new_n44586_, new_n44588_, new_n44589_, new_n44591_,
    new_n44592_, new_n44594_, new_n44595_, new_n44597_, new_n44598_,
    new_n44600_, new_n44601_, new_n44603_, new_n44604_, new_n44605_,
    new_n44606_, new_n44607_, new_n44608_, new_n44609_, new_n44610_,
    new_n44611_, new_n44612_, new_n44613_, new_n44614_, new_n44615_,
    new_n44616_, new_n44617_, new_n44618_, new_n44619_, new_n44620_,
    new_n44621_, new_n44622_, new_n44623_, new_n44624_, new_n44625_,
    new_n44626_, new_n44627_, new_n44628_, new_n44630_, new_n44631_,
    new_n44632_, new_n44634_, new_n44635_, new_n44637_, new_n44638_,
    new_n44639_, new_n44641_, new_n44642_, new_n44644_, new_n44645_,
    new_n44646_, new_n44647_, new_n44648_, new_n44649_, new_n44650_,
    new_n44651_, new_n44652_, new_n44653_, new_n44654_, new_n44656_,
    new_n44657_, new_n44658_, new_n44659_, new_n44661_, new_n44662_,
    new_n44664_, new_n44665_, new_n44666_, new_n44668_, new_n44669_,
    new_n44670_, new_n44671_, new_n44673_, new_n44674_, new_n44676_,
    new_n44677_, new_n44679_, new_n44680_, new_n44682_, new_n44683_,
    new_n44685_, new_n44686_, new_n44688_, new_n44689_, new_n44691_,
    new_n44692_, new_n44694_, new_n44695_, new_n44697_, new_n44698_,
    new_n44700_, new_n44701_, new_n44703_, new_n44704_, new_n44706_,
    new_n44707_, new_n44708_, new_n44709_, new_n44710_, new_n44711_,
    new_n44712_, new_n44714_, new_n44715_, new_n44716_, new_n44717_,
    new_n44719_, new_n44720_, new_n44721_, new_n44722_, new_n44723_,
    new_n44724_, new_n44725_, new_n44726_, new_n44727_, new_n44728_,
    new_n44729_, new_n44731_, new_n44732_, new_n44734_, new_n44735_,
    new_n44737_, new_n44738_, new_n44740_, new_n44741_, new_n44743_,
    new_n44744_, new_n44746_, new_n44747_, new_n44749_, new_n44750_,
    new_n44752_, new_n44753_, new_n44754_, new_n44755_, new_n44756_,
    new_n44758_, new_n44759_, new_n44761_, new_n44762_, new_n44764_,
    new_n44765_, new_n44767_, new_n44768_, new_n44770_, new_n44771_,
    new_n44773_, new_n44774_, new_n44776_, new_n44777_, new_n44779_,
    new_n44780_, new_n44782_, new_n44783_, new_n44785_, new_n44786_,
    new_n44788_, new_n44789_, new_n44791_, new_n44792_, new_n44794_,
    new_n44795_, new_n44797_, new_n44798_, new_n44800_, new_n44801_,
    new_n44803_, new_n44804_, new_n44806_, new_n44807_, new_n44809_,
    new_n44810_, new_n44812_, new_n44813_, new_n44815_, new_n44816_,
    new_n44818_, new_n44819_, new_n44821_, new_n44822_, new_n44824_,
    new_n44825_, new_n44827_, new_n44828_, new_n44830_, new_n44831_,
    new_n44833_, new_n44834_, new_n44836_, new_n44837_, new_n44839_,
    new_n44840_, new_n44842_, new_n44843_, new_n44845_, new_n44846_,
    new_n44848_, new_n44849_, new_n44851_, new_n44852_, new_n44854_,
    new_n44855_, new_n44857_, new_n44858_, new_n44860_, new_n44861_,
    new_n44863_, new_n44864_, new_n44866_, new_n44867_, new_n44869_,
    new_n44870_, new_n44872_, new_n44873_, new_n44875_, new_n44876_,
    new_n44878_, new_n44879_, new_n44881_, new_n44882_, new_n44884_,
    new_n44885_, new_n44887_, new_n44888_, new_n44890_, new_n44891_,
    new_n44893_, new_n44894_, new_n44896_, new_n44897_, new_n44899_,
    new_n44900_, new_n44902_, new_n44903_, new_n44905_, new_n44906_,
    new_n44908_, new_n44909_, new_n44911_, new_n44912_, new_n44914_,
    new_n44915_, new_n44917_, new_n44918_, new_n44920_, new_n44921_,
    new_n44923_, new_n44924_, new_n44926_, new_n44927_, new_n44929_,
    new_n44930_, new_n44932_, new_n44933_, new_n44935_, new_n44936_,
    new_n44938_, new_n44939_, new_n44941_, new_n44942_, new_n44944_,
    new_n44945_, new_n44947_, new_n44948_, new_n44950_, new_n44951_,
    new_n44953_, new_n44954_, new_n44956_, new_n44957_, new_n44959_,
    new_n44960_, new_n44962_, new_n44963_, new_n44965_, new_n44966_,
    new_n44968_, new_n44969_, new_n44971_, new_n44972_, new_n44974_,
    new_n44975_, new_n44977_, new_n44978_, new_n44979_, new_n44981_,
    new_n44982_, new_n44984_, new_n44985_, new_n44987_, new_n44988_,
    new_n44990_, new_n44991_, new_n44993_, new_n44994_, new_n44996_,
    new_n44997_, new_n44999_, new_n45000_, new_n45002_, new_n45003_,
    new_n45005_, new_n45006_, new_n45008_, new_n45009_, new_n45011_,
    new_n45012_, new_n45014_, new_n45015_, new_n45017_, new_n45018_,
    new_n45020_, new_n45021_, new_n45023_, new_n45024_, new_n45026_,
    new_n45027_, new_n45029_, new_n45030_, new_n45032_, new_n45033_,
    new_n45035_, new_n45036_, new_n45038_, new_n45039_, new_n45041_,
    new_n45042_, new_n45044_, new_n45045_, new_n45047_, new_n45048_,
    new_n45050_, new_n45051_, new_n45053_, new_n45054_, new_n45056_,
    new_n45057_, new_n45059_, new_n45060_, new_n45062_, new_n45063_,
    new_n45065_, new_n45066_, new_n45068_, new_n45069_, new_n45071_,
    new_n45072_, new_n45074_, new_n45075_, new_n45077_, new_n45078_,
    new_n45080_, new_n45081_, new_n45083_, new_n45084_, new_n45086_,
    new_n45087_, new_n45089_, new_n45090_, new_n45092_, new_n45093_,
    new_n45095_, new_n45096_, new_n45098_, new_n45099_, new_n45101_,
    new_n45102_, new_n45104_, new_n45105_, new_n45107_, new_n45108_,
    new_n45109_, new_n45110_, new_n45111_, new_n45112_, new_n45113_,
    new_n45114_, new_n45115_, new_n45116_, new_n45117_, new_n45118_,
    new_n45119_, new_n45120_, new_n45121_, new_n45122_, new_n45123_,
    new_n45124_, new_n45125_, new_n45126_, new_n45127_, new_n45128_,
    new_n45129_, new_n45131_, new_n45132_, new_n45134_, new_n45135_,
    new_n45137_, new_n45138_, new_n45140_, new_n45141_, new_n45143_,
    new_n45144_, new_n45146_, new_n45147_, new_n45149_, new_n45150_,
    new_n45152_, new_n45153_, new_n45154_, new_n45155_, new_n45156_,
    new_n45157_, new_n45158_, new_n45159_, new_n45160_, new_n45161_,
    new_n45162_, new_n45163_, new_n45164_, new_n45165_, new_n45166_,
    new_n45167_, new_n45168_, new_n45169_, new_n45170_, new_n45171_,
    new_n45172_, new_n45173_, new_n45174_, new_n45175_, new_n45177_,
    new_n45178_, new_n45179_, new_n45180_, new_n45181_, new_n45182_,
    new_n45183_, new_n45184_, new_n45185_, new_n45186_, new_n45187_,
    new_n45188_, new_n45189_, new_n45190_, new_n45191_, new_n45192_,
    new_n45193_, new_n45195_, new_n45196_, new_n45197_, new_n45198_,
    new_n45199_, new_n45200_, new_n45201_, new_n45202_, new_n45203_,
    new_n45204_, new_n45205_, new_n45206_, new_n45207_, new_n45208_,
    new_n45209_, new_n45210_, new_n45211_, new_n45212_, new_n45213_,
    new_n45214_, new_n45215_, new_n45216_, new_n45217_, new_n45218_,
    new_n45219_, new_n45220_, new_n45221_, new_n45222_, new_n45223_,
    new_n45225_, new_n45226_, new_n45227_, new_n45228_, new_n45229_,
    new_n45231_, new_n45232_, new_n45233_, new_n45234_, new_n45235_,
    new_n45236_, new_n45237_, new_n45238_, new_n45239_, new_n45240_,
    new_n45241_, new_n45242_, new_n45243_, new_n45244_, new_n45245_,
    new_n45246_, new_n45247_, new_n45248_, new_n45249_, new_n45251_,
    new_n45252_, new_n45253_, new_n45254_, new_n45255_, new_n45256_,
    new_n45257_, new_n45258_, new_n45259_, new_n45260_, new_n45261_,
    new_n45262_, new_n45263_, new_n45264_, new_n45265_, new_n45266_,
    new_n45267_, new_n45268_, new_n45269_, new_n45271_, new_n45272_,
    new_n45273_, new_n45274_, new_n45275_, new_n45276_, new_n45277_,
    new_n45278_, new_n45279_, new_n45280_, new_n45281_, new_n45282_,
    new_n45283_, new_n45284_, new_n45285_, new_n45286_, new_n45287_,
    new_n45288_, new_n45289_, new_n45291_, new_n45292_, new_n45293_,
    new_n45294_, new_n45295_, new_n45296_, new_n45297_, new_n45298_,
    new_n45299_, new_n45300_, new_n45301_, new_n45302_, new_n45303_,
    new_n45304_, new_n45305_, new_n45306_, new_n45307_, new_n45308_,
    new_n45309_, new_n45311_, new_n45312_, new_n45313_, new_n45314_,
    new_n45315_, new_n45316_, new_n45317_, new_n45318_, new_n45319_,
    new_n45320_, new_n45322_, new_n45323_, new_n45324_, new_n45325_,
    new_n45326_, new_n45327_, new_n45328_, new_n45329_, new_n45330_,
    new_n45331_, new_n45333_, new_n45334_, new_n45335_, new_n45336_,
    new_n45337_, new_n45338_, new_n45339_, new_n45340_, new_n45341_,
    new_n45342_, new_n45344_, new_n45345_, new_n45346_, new_n45347_,
    new_n45348_, new_n45349_, new_n45350_, new_n45351_, new_n45352_,
    new_n45353_, new_n45354_, new_n45357_, new_n45358_, new_n45360_,
    new_n45361_, new_n45363_, new_n45364_, new_n45366_, new_n45367_,
    new_n45369_, new_n45370_, new_n45372_, new_n45373_, new_n45375_,
    new_n45376_, new_n45378_, new_n45379_, new_n45381_, new_n45382_,
    new_n45384_, new_n45385_, new_n45387_, new_n45388_, new_n45390_,
    new_n45391_, new_n45393_, new_n45394_, new_n45396_, new_n45397_,
    new_n45399_, new_n45400_, new_n45402_, new_n45403_, new_n45405_,
    new_n45406_, new_n45408_, new_n45409_, new_n45411_, new_n45412_,
    new_n45414_, new_n45415_, new_n45417_, new_n45418_, new_n45420_,
    new_n45421_, new_n45423_, new_n45424_, new_n45426_, new_n45427_,
    new_n45429_, new_n45430_, new_n45431_, new_n45432_, new_n45433_,
    new_n45434_, new_n45435_, new_n45436_, new_n45438_, new_n45439_,
    new_n45441_, new_n45442_, new_n45444_, new_n45445_, new_n45447_,
    new_n45448_, new_n45450_, new_n45451_, new_n45453_, new_n45454_,
    new_n45455_, new_n45456_, new_n45457_, new_n45459_, new_n45460_,
    new_n45462_, new_n45463_, new_n45465_, new_n45466_, new_n45468_,
    new_n45469_, new_n45471_, new_n45472_, new_n45474_, new_n45475_,
    new_n45477_, new_n45478_, new_n45479_, new_n45480_, new_n45481_,
    new_n45483_, new_n45484_, new_n45486_, new_n45487_, new_n45489_,
    new_n45490_, new_n45492_, new_n45493_, new_n45495_, new_n45496_,
    new_n45497_, new_n45498_, new_n45500_, new_n45501_, new_n45503_,
    new_n45504_, new_n45506_, new_n45507_, new_n45509_, new_n45510_,
    new_n45512_, new_n45513_, new_n45515_, new_n45516_, new_n45518_,
    new_n45519_, new_n45521_, new_n45522_, new_n45524_, new_n45525_,
    new_n45527_, new_n45528_, new_n45530_, new_n45531_, new_n45533_,
    new_n45534_, new_n45536_, new_n45537_, new_n45539_, new_n45540_,
    new_n45542_, new_n45543_, new_n45545_, new_n45546_, new_n45548_,
    new_n45549_, new_n45551_, new_n45552_, new_n45554_, new_n45555_,
    new_n45557_, new_n45558_, new_n45560_, new_n45561_, new_n45562_,
    new_n45563_, new_n45565_, new_n45566_, new_n45568_, new_n45569_,
    new_n45571_, new_n45572_, new_n45574_, new_n45575_, new_n45577_,
    new_n45578_, new_n45580_, new_n45581_, new_n45583_, new_n45584_,
    new_n45586_, new_n45587_, new_n45589_, new_n45590_, new_n45592_,
    new_n45593_, new_n45595_, new_n45596_, new_n45598_, new_n45599_,
    new_n45601_, new_n45602_, new_n45603_, new_n45604_, new_n45606_,
    new_n45607_, new_n45609_, new_n45610_, new_n45612_, new_n45613_,
    new_n45615_, new_n45616_, new_n45618_, new_n45619_, new_n45621_,
    new_n45622_, new_n45624_, new_n45625_, new_n45627_, new_n45628_,
    new_n45630_, new_n45631_, new_n45633_, new_n45634_, new_n45635_,
    new_n45636_, new_n45637_, new_n45638_, new_n45639_, new_n45640_,
    new_n45641_, new_n45642_, new_n45643_, new_n45644_, new_n45645_,
    new_n45646_, new_n45647_, new_n45648_, new_n45649_, new_n45650_,
    new_n45651_, new_n45652_, new_n45653_, new_n45654_, new_n45655_,
    new_n45656_, new_n45657_, new_n45658_, new_n45659_, new_n45660_,
    new_n45661_, new_n45662_, new_n45663_, new_n45664_, new_n45665_,
    new_n45666_, new_n45667_, new_n45668_, new_n45669_, new_n45670_,
    new_n45671_, new_n45672_, new_n45673_, new_n45674_, new_n45675_,
    new_n45676_, new_n45677_, new_n45678_, new_n45679_, new_n45680_,
    new_n45681_, new_n45682_, new_n45683_, new_n45684_, new_n45685_,
    new_n45686_, new_n45687_, new_n45688_, new_n45689_, new_n45690_,
    new_n45691_, new_n45692_, new_n45693_, new_n45694_, new_n45695_,
    new_n45696_, new_n45697_, new_n45698_, new_n45699_, new_n45700_,
    new_n45701_, new_n45702_, new_n45703_, new_n45704_, new_n45705_,
    new_n45706_, new_n45707_, new_n45708_, new_n45709_, new_n45710_,
    new_n45711_, new_n45712_, new_n45713_, new_n45714_, new_n45715_,
    new_n45716_, new_n45717_, new_n45718_, new_n45719_, new_n45720_,
    new_n45721_, new_n45722_, new_n45723_, new_n45724_, new_n45725_,
    new_n45726_, new_n45727_, new_n45728_, new_n45729_, new_n45730_,
    new_n45731_, new_n45732_, new_n45733_, new_n45734_, new_n45735_,
    new_n45736_, new_n45737_, new_n45738_, new_n45739_, new_n45740_,
    new_n45741_, new_n45742_, new_n45744_, new_n45745_, new_n45747_,
    new_n45748_, new_n45750_, new_n45751_, new_n45752_, new_n45753_,
    new_n45755_, new_n45756_, new_n45758_, new_n45759_, new_n45761_,
    new_n45762_, new_n45764_, new_n45765_, new_n45767_, new_n45768_,
    new_n45770_, new_n45771_, new_n45773_, new_n45774_, new_n45776_,
    new_n45777_, new_n45779_, new_n45780_, new_n45782_, new_n45783_,
    new_n45785_, new_n45786_, new_n45788_, new_n45789_, new_n45791_,
    new_n45792_, new_n45794_, new_n45795_, new_n45797_, new_n45798_,
    new_n45800_, new_n45801_, new_n45802_, new_n45803_, new_n45804_,
    new_n45805_, new_n45807_, new_n45808_, new_n45809_, new_n45810_,
    new_n45812_, new_n45813_, new_n45814_, new_n45815_, new_n45816_,
    new_n45817_, new_n45818_, new_n45819_, new_n45820_, new_n45821_,
    new_n45822_, new_n45823_, new_n45824_, new_n45825_, new_n45826_,
    new_n45827_, new_n45828_, new_n45829_, new_n45830_, new_n45831_,
    new_n45833_, new_n45834_, new_n45835_, new_n45837_, new_n45838_,
    new_n45839_, new_n45841_, new_n45842_, new_n45843_, new_n45845_,
    new_n45846_, new_n45847_, new_n45848_, new_n45849_, new_n45850_,
    new_n45851_, new_n45852_, new_n45853_, new_n45854_, new_n45855_,
    new_n45856_, new_n45857_, new_n45858_, new_n45859_, new_n45860_,
    new_n45861_, new_n45862_, new_n45863_, new_n45864_, new_n45865_,
    new_n45866_, new_n45867_, new_n45868_, new_n45869_, new_n45870_,
    new_n45871_, new_n45872_, new_n45873_, new_n45874_, new_n45875_,
    new_n45876_, new_n45877_, new_n45878_, new_n45879_, new_n45880_,
    new_n45881_, new_n45882_, new_n45883_, new_n45884_, new_n45885_,
    new_n45886_, new_n45887_, new_n45888_, new_n45889_, new_n45890_,
    new_n45891_, new_n45892_, new_n45893_, new_n45894_, new_n45895_,
    new_n45896_, new_n45897_, new_n45898_, new_n45899_, new_n45900_,
    new_n45901_, new_n45902_, new_n45903_, new_n45904_, new_n45905_,
    new_n45906_, new_n45907_, new_n45908_, new_n45909_, new_n45910_,
    new_n45911_, new_n45912_, new_n45913_, new_n45914_, new_n45915_,
    new_n45916_, new_n45917_, new_n45918_, new_n45919_, new_n45920_,
    new_n45921_, new_n45922_, new_n45923_, new_n45924_, new_n45925_,
    new_n45926_, new_n45927_, new_n45928_, new_n45929_, new_n45930_,
    new_n45931_, new_n45932_, new_n45933_, new_n45934_, new_n45935_,
    new_n45936_, new_n45937_, new_n45938_, new_n45939_, new_n45940_,
    new_n45941_, new_n45942_, new_n45943_, new_n45944_, new_n45945_,
    new_n45946_, new_n45947_, new_n45948_, new_n45949_, new_n45950_,
    new_n45951_, new_n45952_, new_n45953_, new_n45954_, new_n45955_,
    new_n45956_, new_n45957_, new_n45958_, new_n45959_, new_n45960_,
    new_n45961_, new_n45962_, new_n45963_, new_n45964_, new_n45965_,
    new_n45966_, new_n45967_, new_n45968_, new_n45969_, new_n45970_,
    new_n45971_, new_n45972_, new_n45973_, new_n45974_, new_n45975_,
    new_n45976_, new_n45977_, new_n45978_, new_n45979_, new_n45980_,
    new_n45981_, new_n45982_, new_n45983_, new_n45984_, new_n45985_,
    new_n45986_, new_n45987_, new_n45988_, new_n45989_, new_n45990_,
    new_n45991_, new_n45992_, new_n45993_, new_n45994_, new_n45995_,
    new_n45996_, new_n45997_, new_n45998_, new_n45999_, new_n46000_,
    new_n46001_, new_n46002_, new_n46003_, new_n46004_, new_n46005_,
    new_n46006_, new_n46007_, new_n46008_, new_n46009_, new_n46010_,
    new_n46011_, new_n46012_, new_n46013_, new_n46014_, new_n46015_,
    new_n46016_, new_n46017_, new_n46018_, new_n46019_, new_n46020_,
    new_n46021_, new_n46022_, new_n46023_, new_n46024_, new_n46025_,
    new_n46026_, new_n46027_, new_n46028_, new_n46029_, new_n46030_,
    new_n46031_, new_n46032_, new_n46033_, new_n46034_, new_n46035_,
    new_n46036_, new_n46037_, new_n46038_, new_n46039_, new_n46040_,
    new_n46041_, new_n46042_, new_n46043_, new_n46044_, new_n46045_,
    new_n46046_, new_n46047_, new_n46048_, new_n46049_, new_n46050_,
    new_n46051_, new_n46052_, new_n46053_, new_n46054_, new_n46055_,
    new_n46056_, new_n46057_, new_n46058_, new_n46059_, new_n46060_,
    new_n46061_, new_n46062_, new_n46063_, new_n46064_, new_n46065_,
    new_n46066_, new_n46067_, new_n46068_, new_n46069_, new_n46070_,
    new_n46071_, new_n46072_, new_n46073_, new_n46074_, new_n46075_,
    new_n46076_, new_n46077_, new_n46078_, new_n46079_, new_n46080_,
    new_n46081_, new_n46082_, new_n46083_, new_n46084_, new_n46085_,
    new_n46086_, new_n46087_, new_n46088_, new_n46089_, new_n46090_,
    new_n46091_, new_n46092_, new_n46093_, new_n46094_, new_n46095_,
    new_n46096_, new_n46097_, new_n46098_, new_n46099_, new_n46100_,
    new_n46101_, new_n46102_, new_n46103_, new_n46104_, new_n46105_,
    new_n46106_, new_n46107_, new_n46108_, new_n46109_, new_n46110_,
    new_n46111_, new_n46112_, new_n46113_, new_n46114_, new_n46115_,
    new_n46116_, new_n46117_, new_n46118_, new_n46119_, new_n46120_,
    new_n46121_, new_n46122_, new_n46123_, new_n46124_, new_n46125_,
    new_n46126_, new_n46127_, new_n46128_, new_n46129_, new_n46130_,
    new_n46131_, new_n46132_, new_n46133_, new_n46134_, new_n46135_,
    new_n46136_, new_n46137_, new_n46138_, new_n46139_, new_n46140_,
    new_n46141_, new_n46142_, new_n46143_, new_n46144_, new_n46145_,
    new_n46146_, new_n46147_, new_n46148_, new_n46149_, new_n46150_,
    new_n46151_, new_n46152_, new_n46153_, new_n46154_, new_n46155_,
    new_n46156_, new_n46157_, new_n46158_, new_n46159_, new_n46160_,
    new_n46161_, new_n46162_, new_n46163_, new_n46164_, new_n46165_,
    new_n46166_, new_n46167_, new_n46168_, new_n46169_, new_n46170_,
    new_n46171_, new_n46172_, new_n46173_, new_n46174_, new_n46175_,
    new_n46176_, new_n46177_, new_n46178_, new_n46179_, new_n46180_,
    new_n46181_, new_n46182_, new_n46183_, new_n46184_, new_n46185_,
    new_n46186_, new_n46187_, new_n46188_, new_n46189_, new_n46190_,
    new_n46191_, new_n46192_, new_n46193_, new_n46194_, new_n46195_,
    new_n46196_, new_n46197_, new_n46198_, new_n46199_, new_n46200_,
    new_n46201_, new_n46202_, new_n46203_, new_n46204_, new_n46205_,
    new_n46206_, new_n46207_, new_n46208_, new_n46209_, new_n46210_,
    new_n46211_, new_n46212_, new_n46213_, new_n46214_, new_n46215_,
    new_n46216_, new_n46217_, new_n46218_, new_n46219_, new_n46220_,
    new_n46221_, new_n46222_, new_n46223_, new_n46224_, new_n46225_,
    new_n46226_, new_n46227_, new_n46228_, new_n46229_, new_n46230_,
    new_n46231_, new_n46232_, new_n46233_, new_n46234_, new_n46235_,
    new_n46236_, new_n46237_, new_n46238_, new_n46239_, new_n46240_,
    new_n46241_, new_n46242_, new_n46243_, new_n46244_, new_n46245_,
    new_n46246_, new_n46247_, new_n46248_, new_n46249_, new_n46250_,
    new_n46251_, new_n46252_, new_n46253_, new_n46254_, new_n46255_,
    new_n46256_, new_n46257_, new_n46258_, new_n46259_, new_n46260_,
    new_n46261_, new_n46262_, new_n46263_, new_n46264_, new_n46265_,
    new_n46266_, new_n46267_, new_n46268_, new_n46269_, new_n46270_,
    new_n46271_, new_n46272_, new_n46273_, new_n46274_, new_n46275_,
    new_n46276_, new_n46277_, new_n46278_, new_n46279_, new_n46280_,
    new_n46281_, new_n46282_, new_n46283_, new_n46284_, new_n46285_,
    new_n46286_, new_n46287_, new_n46288_, new_n46289_, new_n46290_,
    new_n46291_, new_n46292_, new_n46293_, new_n46294_, new_n46295_,
    new_n46296_, new_n46297_, new_n46298_, new_n46299_, new_n46300_,
    new_n46301_, new_n46302_, new_n46303_, new_n46304_, new_n46305_,
    new_n46306_, new_n46307_, new_n46308_, new_n46309_, new_n46310_,
    new_n46311_, new_n46312_, new_n46313_, new_n46314_, new_n46315_,
    new_n46316_, new_n46317_, new_n46318_, new_n46319_, new_n46320_,
    new_n46321_, new_n46322_, new_n46323_, new_n46324_, new_n46325_,
    new_n46326_, new_n46327_, new_n46328_, new_n46329_, new_n46330_,
    new_n46331_, new_n46332_, new_n46333_, new_n46334_, new_n46335_,
    new_n46336_, new_n46337_, new_n46338_, new_n46339_, new_n46340_,
    new_n46341_, new_n46342_, new_n46343_, new_n46344_, new_n46345_,
    new_n46346_, new_n46347_, new_n46348_, new_n46349_, new_n46350_,
    new_n46351_, new_n46352_, new_n46353_, new_n46354_, new_n46355_,
    new_n46356_, new_n46357_, new_n46358_, new_n46359_, new_n46360_,
    new_n46361_, new_n46362_, new_n46363_, new_n46364_, new_n46365_,
    new_n46366_, new_n46367_, new_n46368_, new_n46369_, new_n46370_,
    new_n46371_, new_n46372_, new_n46373_, new_n46374_, new_n46375_,
    new_n46376_, new_n46377_, new_n46378_, new_n46379_, new_n46380_,
    new_n46381_, new_n46382_, new_n46383_, new_n46384_, new_n46385_,
    new_n46386_, new_n46387_, new_n46388_, new_n46389_, new_n46390_,
    new_n46391_, new_n46392_, new_n46393_, new_n46394_, new_n46395_,
    new_n46396_, new_n46397_, new_n46398_, new_n46399_, new_n46400_,
    new_n46401_, new_n46402_, new_n46403_, new_n46404_, new_n46405_,
    new_n46406_, new_n46407_, new_n46408_, new_n46409_, new_n46410_,
    new_n46411_, new_n46412_, new_n46413_, new_n46414_, new_n46415_,
    new_n46416_, new_n46417_, new_n46418_, new_n46419_, new_n46420_,
    new_n46421_, new_n46422_, new_n46423_, new_n46424_, new_n46425_,
    new_n46426_, new_n46427_, new_n46428_, new_n46429_, new_n46430_,
    new_n46431_, new_n46432_, new_n46433_, new_n46434_, new_n46435_,
    new_n46436_, new_n46437_, new_n46438_, new_n46439_, new_n46440_,
    new_n46441_, new_n46442_, new_n46443_, new_n46444_, new_n46445_,
    new_n46446_, new_n46447_, new_n46448_, new_n46449_, new_n46450_,
    new_n46451_, new_n46452_, new_n46453_, new_n46454_, new_n46455_,
    new_n46456_, new_n46457_, new_n46458_, new_n46459_, new_n46460_,
    new_n46461_, new_n46462_, new_n46463_, new_n46464_, new_n46465_,
    new_n46466_, new_n46467_, new_n46468_, new_n46469_, new_n46470_,
    new_n46471_, new_n46472_, new_n46473_, new_n46474_, new_n46475_,
    new_n46476_, new_n46477_, new_n46478_, new_n46479_, new_n46480_,
    new_n46481_, new_n46482_, new_n46483_, new_n46484_, new_n46485_,
    new_n46486_, new_n46487_, new_n46488_, new_n46489_, new_n46490_,
    new_n46491_, new_n46492_, new_n46493_, new_n46494_, new_n46495_,
    new_n46496_, new_n46497_, new_n46498_, new_n46499_, new_n46500_,
    new_n46501_, new_n46502_, new_n46503_, new_n46504_, new_n46505_,
    new_n46506_, new_n46507_, new_n46508_, new_n46509_, new_n46510_,
    new_n46511_, new_n46512_, new_n46513_, new_n46514_, new_n46515_,
    new_n46516_, new_n46517_, new_n46518_, new_n46519_, new_n46520_,
    new_n46521_, new_n46522_, new_n46523_, new_n46524_, new_n46525_,
    new_n46526_, new_n46527_, new_n46528_, new_n46529_, new_n46530_,
    new_n46531_, new_n46532_, new_n46533_, new_n46534_, new_n46535_,
    new_n46536_, new_n46537_, new_n46538_, new_n46539_, new_n46540_,
    new_n46541_, new_n46542_, new_n46543_, new_n46544_, new_n46545_,
    new_n46546_, new_n46547_, new_n46548_, new_n46549_, new_n46550_,
    new_n46551_, new_n46552_, new_n46553_, new_n46554_, new_n46555_,
    new_n46556_, new_n46557_, new_n46558_, new_n46559_, new_n46560_,
    new_n46561_, new_n46562_, new_n46563_, new_n46564_, new_n46565_,
    new_n46566_, new_n46567_, new_n46568_, new_n46569_, new_n46570_,
    new_n46571_, new_n46572_, new_n46573_, new_n46574_, new_n46575_,
    new_n46576_, new_n46577_, new_n46578_, new_n46579_, new_n46580_,
    new_n46581_, new_n46582_, new_n46583_, new_n46584_, new_n46585_,
    new_n46586_, new_n46587_, new_n46588_, new_n46589_, new_n46590_,
    new_n46591_, new_n46592_, new_n46593_, new_n46594_, new_n46595_,
    new_n46596_, new_n46597_, new_n46598_, new_n46599_, new_n46600_,
    new_n46601_, new_n46602_, new_n46603_, new_n46604_, new_n46605_,
    new_n46606_, new_n46607_, new_n46608_, new_n46609_, new_n46610_,
    new_n46611_, new_n46612_, new_n46613_, new_n46614_, new_n46615_,
    new_n46616_, new_n46617_, new_n46618_, new_n46619_, new_n46620_,
    new_n46621_, new_n46622_, new_n46623_, new_n46624_, new_n46625_,
    new_n46626_, new_n46627_, new_n46628_, new_n46629_, new_n46630_,
    new_n46631_, new_n46632_, new_n46633_, new_n46634_, new_n46635_,
    new_n46636_, new_n46637_, new_n46638_, new_n46639_, new_n46640_,
    new_n46641_, new_n46642_, new_n46643_, new_n46644_, new_n46645_,
    new_n46646_, new_n46647_, new_n46648_, new_n46649_, new_n46650_,
    new_n46651_, new_n46652_, new_n46653_, new_n46654_, new_n46655_,
    new_n46656_, new_n46657_, new_n46658_, new_n46659_, new_n46660_,
    new_n46661_, new_n46662_, new_n46663_, new_n46664_, new_n46665_,
    new_n46666_, new_n46667_, new_n46668_, new_n46669_, new_n46670_,
    new_n46671_, new_n46672_, new_n46673_, new_n46674_, new_n46675_,
    new_n46676_, new_n46677_, new_n46678_, new_n46679_, new_n46680_,
    new_n46681_, new_n46682_, new_n46683_, new_n46684_, new_n46685_,
    new_n46686_, new_n46687_, new_n46688_, new_n46689_, new_n46690_,
    new_n46691_, new_n46692_, new_n46693_, new_n46694_, new_n46695_,
    new_n46696_, new_n46697_, new_n46698_, new_n46699_, new_n46700_,
    new_n46701_, new_n46702_, new_n46703_, new_n46704_, new_n46705_,
    new_n46706_, new_n46707_, new_n46708_, new_n46709_, new_n46710_,
    new_n46711_, new_n46712_, new_n46713_, new_n46714_, new_n46715_,
    new_n46716_, new_n46717_, new_n46718_, new_n46719_, new_n46720_,
    new_n46721_, new_n46722_, new_n46724_, new_n46725_, new_n46726_,
    new_n46727_, new_n46728_, new_n46729_, new_n46731_, new_n46732_,
    new_n46733_, new_n46734_, new_n46735_, new_n46737_, new_n46738_,
    new_n46739_, new_n46740_, new_n46741_, new_n46743_, new_n46744_,
    new_n46745_, new_n46747_, new_n46748_, new_n46749_, new_n46750_,
    new_n46751_, new_n46753_, new_n46754_, new_n46755_, new_n46757_,
    new_n46758_, new_n46760_, new_n46761_, new_n46762_, new_n46764_,
    new_n46765_, new_n46766_, new_n46767_, new_n46768_, new_n46769_,
    new_n46770_, new_n46771_, new_n46772_, new_n46773_, new_n46774_,
    new_n46776_, new_n46777_, new_n46778_, new_n46779_, new_n46781_,
    new_n46782_, new_n46783_, new_n46784_, new_n46785_, new_n46786_,
    new_n46787_, new_n46788_, new_n46790_, new_n46791_, new_n46792_,
    new_n46793_, new_n46794_, new_n46795_, new_n46797_, new_n46798_,
    new_n46800_, new_n46801_, new_n46802_, new_n46803_, new_n46804_,
    new_n46806_, new_n46807_, new_n46808_, new_n46810_, new_n46811_,
    new_n46812_, new_n46814_, new_n46815_, new_n46816_, new_n46818_,
    new_n46819_, new_n46820_, new_n46822_, new_n46823_, new_n46824_,
    new_n46826_, new_n46827_, new_n46828_, new_n46830_, new_n46831_,
    new_n46832_, new_n46834_, new_n46835_, new_n46836_, new_n46837_,
    new_n46839_, new_n46840_, new_n46841_, new_n46842_, new_n46844_,
    new_n46845_, new_n46846_, new_n46847_, new_n46849_, new_n46850_,
    new_n46851_, new_n46852_, new_n46853_, new_n46855_, new_n46856_,
    new_n46857_, new_n46859_, new_n46860_, new_n46861_, new_n46863_,
    new_n46864_, new_n46865_, new_n46867_, new_n46868_, new_n46869_,
    new_n46871_, new_n46872_, new_n46873_, new_n46875_, new_n46876_,
    new_n46877_, new_n46879_, new_n46880_, new_n46881_, new_n46882_,
    new_n46883_, new_n46885_, new_n46886_, new_n46887_, new_n46888_,
    new_n46890_, new_n46891_, new_n46892_, new_n46894_, new_n46895_,
    new_n46896_, new_n46898_, new_n46899_, new_n46900_, new_n46902_,
    new_n46903_, new_n46904_, new_n46906_, new_n46907_, new_n46908_,
    new_n46910_, new_n46911_, new_n46912_, new_n46914_, new_n46915_,
    new_n46916_, new_n46918_, new_n46919_, new_n46920_, new_n46922_,
    new_n46923_, new_n46924_, new_n46926_, new_n46927_, new_n46928_,
    new_n46930_, new_n46931_, new_n46932_, new_n46934_, new_n46935_,
    new_n46936_, new_n46938_, new_n46939_, new_n46940_, new_n46942_,
    new_n46943_, new_n46944_, new_n46946_, new_n46947_, new_n46948_,
    new_n46950_, new_n46951_, new_n46952_, new_n46954_, new_n46955_,
    new_n46956_, new_n46958_, new_n46959_, new_n46960_, new_n46962_,
    new_n46963_, new_n46964_, new_n46966_, new_n46967_, new_n46968_,
    new_n46970_, new_n46971_, new_n46972_, new_n46974_, new_n46975_,
    new_n46976_, new_n46978_, new_n46979_, new_n46980_, new_n46982_,
    new_n46983_, new_n46984_, new_n46986_, new_n46987_, new_n46988_,
    new_n46990_, new_n46991_, new_n46992_, new_n46994_, new_n46995_,
    new_n46996_, new_n46998_, new_n46999_, new_n47000_, new_n47002_,
    new_n47003_, new_n47004_, new_n47006_, new_n47007_, new_n47008_,
    new_n47010_, new_n47011_, new_n47012_, new_n47014_, new_n47015_,
    new_n47016_, new_n47018_, new_n47019_, new_n47020_, new_n47022_,
    new_n47023_, new_n47024_, new_n47026_, new_n47027_, new_n47028_,
    new_n47029_, new_n47030_, new_n47031_, new_n47032_, new_n47033_,
    new_n47034_, new_n47036_, new_n47038_, new_n47039_, new_n47040_,
    new_n47042_, new_n47043_, new_n47044_, new_n47046_, new_n47047_,
    new_n47048_, new_n47050_, new_n47051_, new_n47052_, new_n47053_,
    new_n47054_, new_n47055_, new_n47056_, new_n47057_, new_n47058_,
    new_n47059_, new_n47060_, new_n47061_, new_n47062_, new_n47063_,
    new_n47064_, new_n47065_, new_n47066_, new_n47067_, new_n47068_,
    new_n47069_, new_n47070_, new_n47071_, new_n47072_, new_n47073_,
    new_n47074_, new_n47075_, new_n47076_, new_n47077_, new_n47078_,
    new_n47079_, new_n47080_, new_n47081_, new_n47082_, new_n47083_,
    new_n47084_, new_n47085_, new_n47086_, new_n47087_, new_n47088_,
    new_n47089_, new_n47090_, new_n47091_, new_n47092_, new_n47093_,
    new_n47094_, new_n47095_, new_n47096_, new_n47097_, new_n47099_,
    new_n47100_, new_n47101_, new_n47102_, new_n47103_, new_n47104_,
    new_n47105_, new_n47106_, new_n47107_, new_n47108_, new_n47109_,
    new_n47110_, new_n47111_, new_n47112_, new_n47113_, new_n47114_,
    new_n47115_, new_n47116_, new_n47117_, new_n47118_, new_n47119_,
    new_n47120_, new_n47121_, new_n47122_, new_n47123_, new_n47124_,
    new_n47125_, new_n47126_, new_n47127_, new_n47128_, new_n47129_,
    new_n47130_, new_n47131_, new_n47132_, new_n47133_, new_n47134_,
    new_n47135_, new_n47136_, new_n47137_, new_n47138_, new_n47139_,
    new_n47141_, new_n47142_, new_n47143_, new_n47145_, new_n47146_,
    new_n47147_, new_n47148_, new_n47149_, new_n47150_, new_n47151_,
    new_n47152_, new_n47153_, new_n47154_, new_n47155_, new_n47156_,
    new_n47157_, new_n47158_, new_n47159_, new_n47160_, new_n47161_,
    new_n47162_, new_n47163_, new_n47164_, new_n47165_, new_n47166_,
    new_n47167_, new_n47168_, new_n47169_, new_n47170_, new_n47171_,
    new_n47172_, new_n47173_, new_n47174_, new_n47175_, new_n47176_,
    new_n47177_, new_n47178_, new_n47179_, new_n47181_, new_n47182_,
    new_n47183_, new_n47184_, new_n47185_, new_n47186_, new_n47187_,
    new_n47188_, new_n47189_, new_n47190_, new_n47191_, new_n47192_,
    new_n47193_, new_n47194_, new_n47195_, new_n47196_, new_n47197_,
    new_n47198_, new_n47199_, new_n47200_, new_n47201_, new_n47202_,
    new_n47203_, new_n47204_, new_n47205_, new_n47206_, new_n47207_,
    new_n47208_, new_n47209_, new_n47210_, new_n47211_, new_n47212_,
    new_n47213_, new_n47214_, new_n47215_, new_n47216_, new_n47218_,
    new_n47219_, new_n47220_, new_n47221_, new_n47222_, new_n47223_,
    new_n47224_, new_n47225_, new_n47226_, new_n47227_, new_n47228_,
    new_n47229_, new_n47230_, new_n47231_, new_n47232_, new_n47233_,
    new_n47234_, new_n47235_, new_n47236_, new_n47237_, new_n47238_,
    new_n47239_, new_n47240_, new_n47241_, new_n47242_, new_n47243_,
    new_n47244_, new_n47245_, new_n47246_, new_n47247_, new_n47248_,
    new_n47249_, new_n47250_, new_n47251_, new_n47252_, new_n47254_,
    new_n47255_, new_n47256_, new_n47258_, new_n47259_, new_n47260_,
    new_n47261_, new_n47262_, new_n47263_, new_n47264_, new_n47265_,
    new_n47266_, new_n47267_, new_n47268_, new_n47269_, new_n47270_,
    new_n47271_, new_n47272_, new_n47273_, new_n47274_, new_n47275_,
    new_n47276_, new_n47277_, new_n47278_, new_n47279_, new_n47280_,
    new_n47281_, new_n47282_, new_n47283_, new_n47284_, new_n47285_,
    new_n47286_, new_n47287_, new_n47288_, new_n47289_, new_n47291_,
    new_n47292_, new_n47293_, new_n47294_, new_n47295_, new_n47296_,
    new_n47297_, new_n47298_, new_n47299_, new_n47300_, new_n47301_,
    new_n47302_, new_n47303_, new_n47304_, new_n47305_, new_n47306_,
    new_n47307_, new_n47308_, new_n47309_, new_n47310_, new_n47311_,
    new_n47312_, new_n47313_, new_n47314_, new_n47315_, new_n47316_,
    new_n47317_, new_n47318_, new_n47319_, new_n47320_, new_n47321_,
    new_n47323_, new_n47324_, new_n47325_, new_n47326_, new_n47327_,
    new_n47328_, new_n47329_, new_n47330_, new_n47331_, new_n47332_,
    new_n47333_, new_n47334_, new_n47335_, new_n47336_, new_n47337_,
    new_n47338_, new_n47339_, new_n47340_, new_n47341_, new_n47342_,
    new_n47343_, new_n47344_, new_n47345_, new_n47346_, new_n47347_,
    new_n47348_, new_n47349_, new_n47350_, new_n47351_, new_n47352_,
    new_n47353_, new_n47354_, new_n47355_, new_n47356_, new_n47357_,
    new_n47359_, new_n47360_, new_n47361_, new_n47362_, new_n47363_,
    new_n47364_, new_n47365_, new_n47366_, new_n47367_, new_n47368_,
    new_n47369_, new_n47370_, new_n47371_, new_n47372_, new_n47373_,
    new_n47374_, new_n47375_, new_n47376_, new_n47377_, new_n47378_,
    new_n47379_, new_n47380_, new_n47381_, new_n47382_, new_n47383_,
    new_n47384_, new_n47385_, new_n47386_, new_n47387_, new_n47388_,
    new_n47389_, new_n47390_, new_n47391_, new_n47392_, new_n47393_,
    new_n47395_, new_n47396_, new_n47397_, new_n47398_, new_n47399_,
    new_n47400_, new_n47401_, new_n47402_, new_n47403_, new_n47404_,
    new_n47405_, new_n47406_, new_n47407_, new_n47408_, new_n47409_,
    new_n47410_, new_n47411_, new_n47412_, new_n47413_, new_n47414_,
    new_n47415_, new_n47416_, new_n47417_, new_n47418_, new_n47419_,
    new_n47420_, new_n47421_, new_n47422_, new_n47423_, new_n47424_,
    new_n47425_, new_n47426_, new_n47427_, new_n47428_, new_n47429_,
    new_n47430_, new_n47431_, new_n47433_, new_n47434_, new_n47435_,
    new_n47436_, new_n47437_, new_n47438_, new_n47439_, new_n47440_,
    new_n47441_, new_n47442_, new_n47443_, new_n47444_, new_n47445_,
    new_n47446_, new_n47447_, new_n47448_, new_n47449_, new_n47450_,
    new_n47451_, new_n47452_, new_n47453_, new_n47454_, new_n47455_,
    new_n47456_, new_n47457_, new_n47458_, new_n47459_, new_n47460_,
    new_n47461_, new_n47462_, new_n47463_, new_n47464_, new_n47465_,
    new_n47466_, new_n47467_, new_n47469_, new_n47470_, new_n47471_,
    new_n47472_, new_n47473_, new_n47474_, new_n47475_, new_n47476_,
    new_n47477_, new_n47478_, new_n47479_, new_n47480_, new_n47481_,
    new_n47482_, new_n47483_, new_n47484_, new_n47485_, new_n47486_,
    new_n47487_, new_n47488_, new_n47489_, new_n47490_, new_n47491_,
    new_n47492_, new_n47493_, new_n47494_, new_n47495_, new_n47496_,
    new_n47497_, new_n47498_, new_n47499_, new_n47500_, new_n47501_,
    new_n47502_, new_n47503_, new_n47505_, new_n47506_, new_n47507_,
    new_n47508_, new_n47509_, new_n47510_, new_n47511_, new_n47512_,
    new_n47513_, new_n47514_, new_n47515_, new_n47516_, new_n47517_,
    new_n47518_, new_n47519_, new_n47520_, new_n47521_, new_n47522_,
    new_n47523_, new_n47524_, new_n47525_, new_n47526_, new_n47527_,
    new_n47528_, new_n47529_, new_n47530_, new_n47531_, new_n47532_,
    new_n47533_, new_n47534_, new_n47535_, new_n47537_, new_n47538_,
    new_n47539_, new_n47540_, new_n47541_, new_n47542_, new_n47543_,
    new_n47544_, new_n47545_, new_n47546_, new_n47547_, new_n47548_,
    new_n47549_, new_n47550_, new_n47551_, new_n47552_, new_n47553_,
    new_n47554_, new_n47555_, new_n47556_, new_n47557_, new_n47558_,
    new_n47559_, new_n47560_, new_n47561_, new_n47562_, new_n47563_,
    new_n47564_, new_n47565_, new_n47566_, new_n47567_, new_n47569_,
    new_n47570_, new_n47571_, new_n47572_, new_n47573_, new_n47574_,
    new_n47575_, new_n47576_, new_n47577_, new_n47578_, new_n47579_,
    new_n47580_, new_n47581_, new_n47582_, new_n47583_, new_n47584_,
    new_n47585_, new_n47586_, new_n47587_, new_n47588_, new_n47589_,
    new_n47590_, new_n47591_, new_n47592_, new_n47593_, new_n47594_,
    new_n47595_, new_n47596_, new_n47597_, new_n47598_, new_n47599_,
    new_n47600_, new_n47601_, new_n47602_, new_n47603_, new_n47604_,
    new_n47606_, new_n47607_, new_n47608_, new_n47610_, new_n47611_,
    new_n47612_, new_n47614_, new_n47615_, new_n47616_, new_n47617_,
    new_n47618_, new_n47619_, new_n47620_, new_n47621_, new_n47622_,
    new_n47623_, new_n47624_, new_n47625_, new_n47626_, new_n47627_,
    new_n47628_, new_n47629_, new_n47630_, new_n47631_, new_n47632_,
    new_n47633_, new_n47634_, new_n47635_, new_n47636_, new_n47637_,
    new_n47638_, new_n47639_, new_n47640_, new_n47641_, new_n47642_,
    new_n47643_, new_n47644_, new_n47647_, new_n47648_, new_n47649_,
    new_n47651_, new_n47652_, new_n47653_, new_n47654_, new_n47655_,
    new_n47656_, new_n47657_, new_n47658_, new_n47659_, new_n47660_,
    new_n47661_, new_n47662_, new_n47663_, new_n47664_, new_n47665_,
    new_n47666_, new_n47667_, new_n47668_, new_n47669_, new_n47670_,
    new_n47671_, new_n47672_, new_n47673_, new_n47674_, new_n47675_,
    new_n47676_, new_n47677_, new_n47678_, new_n47679_, new_n47680_,
    new_n47681_, new_n47682_, new_n47683_, new_n47684_, new_n47685_,
    new_n47686_, new_n47687_, new_n47688_, new_n47689_, new_n47691_,
    new_n47692_, new_n47693_, new_n47695_, new_n47696_, new_n47697_,
    new_n47699_, new_n47700_, new_n47701_, new_n47703_, new_n47704_,
    new_n47705_, new_n47706_, new_n47707_, new_n47708_, new_n47709_,
    new_n47710_, new_n47711_, new_n47712_, new_n47713_, new_n47714_,
    new_n47715_, new_n47716_, new_n47717_, new_n47718_, new_n47719_,
    new_n47720_, new_n47721_, new_n47722_, new_n47723_, new_n47724_,
    new_n47725_, new_n47726_, new_n47727_, new_n47728_, new_n47729_,
    new_n47730_, new_n47731_, new_n47732_, new_n47733_, new_n47734_,
    new_n47735_, new_n47737_, new_n47738_, new_n47739_, new_n47741_,
    new_n47742_, new_n47743_, new_n47745_, new_n47746_, new_n47747_,
    new_n47748_, new_n47749_, new_n47750_, new_n47751_, new_n47752_,
    new_n47753_, new_n47754_, new_n47755_, new_n47756_, new_n47757_,
    new_n47758_, new_n47759_, new_n47760_, new_n47761_, new_n47762_,
    new_n47763_, new_n47764_, new_n47765_, new_n47766_, new_n47767_,
    new_n47768_, new_n47769_, new_n47770_, new_n47771_, new_n47772_,
    new_n47773_, new_n47774_, new_n47775_, new_n47776_, new_n47777_,
    new_n47778_, new_n47780_, new_n47781_, new_n47782_, new_n47784_,
    new_n47785_, new_n47786_, new_n47788_, new_n47789_, new_n47790_,
    new_n47792_, new_n47793_, new_n47794_, new_n47796_, new_n47797_,
    new_n47798_, new_n47800_, new_n47801_, new_n47802_, new_n47804_,
    new_n47805_, new_n47806_, new_n47808_, new_n47809_, new_n47810_,
    new_n47812_, new_n47813_, new_n47814_, new_n47816_, new_n47817_,
    new_n47818_, new_n47820_, new_n47821_, new_n47822_, new_n47824_,
    new_n47825_, new_n47826_, new_n47828_, new_n47829_, new_n47830_,
    new_n47832_, new_n47833_, new_n47834_, new_n47836_, new_n47837_,
    new_n47838_, new_n47839_, new_n47840_, new_n47841_, new_n47842_,
    new_n47843_, new_n47844_, new_n47845_, new_n47846_, new_n47847_,
    new_n47848_, new_n47849_, new_n47850_, new_n47851_, new_n47852_,
    new_n47853_, new_n47854_, new_n47855_, new_n47856_, new_n47857_,
    new_n47858_, new_n47859_, new_n47860_, new_n47861_, new_n47862_,
    new_n47863_, new_n47864_, new_n47865_, new_n47866_, new_n47867_,
    new_n47868_, new_n47869_, new_n47870_, new_n47872_, new_n47873_,
    new_n47874_, new_n47875_, new_n47876_, new_n47877_, new_n47878_,
    new_n47879_, new_n47880_, new_n47881_, new_n47882_, new_n47883_,
    new_n47884_, new_n47885_, new_n47886_, new_n47887_, new_n47888_,
    new_n47889_, new_n47890_, new_n47891_, new_n47892_, new_n47893_,
    new_n47894_, new_n47895_, new_n47896_, new_n47897_, new_n47898_,
    new_n47899_, new_n47900_, new_n47901_, new_n47902_, new_n47903_,
    new_n47904_, new_n47905_, new_n47906_, new_n47907_, new_n47908_,
    new_n47909_, new_n47910_, new_n47912_, new_n47913_, new_n47914_,
    new_n47916_, new_n47917_, new_n47918_, new_n47920_, new_n47921_,
    new_n47922_, new_n47923_, new_n47924_, new_n47925_, new_n47926_,
    new_n47927_, new_n47928_, new_n47929_, new_n47930_, new_n47931_,
    new_n47932_, new_n47933_, new_n47934_, new_n47935_, new_n47936_,
    new_n47937_, new_n47938_, new_n47939_, new_n47940_, new_n47941_,
    new_n47942_, new_n47943_, new_n47944_, new_n47945_, new_n47946_,
    new_n47947_, new_n47948_, new_n47949_, new_n47950_, new_n47951_,
    new_n47952_, new_n47954_, new_n47955_, new_n47956_, new_n47957_,
    new_n47958_, new_n47959_, new_n47960_, new_n47961_, new_n47962_,
    new_n47963_, new_n47964_, new_n47965_, new_n47966_, new_n47967_,
    new_n47968_, new_n47969_, new_n47970_, new_n47971_, new_n47972_,
    new_n47973_, new_n47974_, new_n47975_, new_n47976_, new_n47977_,
    new_n47978_, new_n47979_, new_n47980_, new_n47981_, new_n47982_,
    new_n47983_, new_n47984_, new_n47985_, new_n47986_, new_n47987_,
    new_n47989_, new_n47990_, new_n47991_, new_n47992_, new_n47993_,
    new_n47994_, new_n47995_, new_n47996_, new_n47997_, new_n47998_,
    new_n47999_, new_n48000_, new_n48001_, new_n48002_, new_n48003_,
    new_n48004_, new_n48005_, new_n48006_, new_n48007_, new_n48008_,
    new_n48009_, new_n48010_, new_n48011_, new_n48012_, new_n48013_,
    new_n48014_, new_n48015_, new_n48016_, new_n48017_, new_n48018_,
    new_n48019_, new_n48020_, new_n48021_, new_n48023_, new_n48024_,
    new_n48025_, new_n48026_, new_n48027_, new_n48028_, new_n48029_,
    new_n48030_, new_n48031_, new_n48032_, new_n48033_, new_n48034_,
    new_n48035_, new_n48036_, new_n48037_, new_n48038_, new_n48039_,
    new_n48040_, new_n48041_, new_n48042_, new_n48043_, new_n48044_,
    new_n48045_, new_n48046_, new_n48047_, new_n48048_, new_n48049_,
    new_n48050_, new_n48051_, new_n48052_, new_n48053_, new_n48054_,
    new_n48055_, new_n48056_, new_n48058_, new_n48059_, new_n48060_,
    new_n48062_, new_n48063_, new_n48064_, new_n48065_, new_n48066_,
    new_n48067_, new_n48068_, new_n48069_, new_n48070_, new_n48071_,
    new_n48072_, new_n48073_, new_n48074_, new_n48075_, new_n48076_,
    new_n48077_, new_n48078_, new_n48079_, new_n48080_, new_n48081_,
    new_n48082_, new_n48083_, new_n48084_, new_n48085_, new_n48086_,
    new_n48087_, new_n48088_, new_n48089_, new_n48090_, new_n48091_,
    new_n48092_, new_n48093_, new_n48094_, new_n48095_, new_n48096_,
    new_n48098_, new_n48099_, new_n48100_, new_n48101_, new_n48102_,
    new_n48103_, new_n48104_, new_n48105_, new_n48106_, new_n48107_,
    new_n48108_, new_n48109_, new_n48110_, new_n48111_, new_n48112_,
    new_n48113_, new_n48114_, new_n48115_, new_n48116_, new_n48117_,
    new_n48118_, new_n48119_, new_n48120_, new_n48121_, new_n48122_,
    new_n48123_, new_n48124_, new_n48125_, new_n48126_, new_n48127_,
    new_n48128_, new_n48129_, new_n48130_, new_n48132_, new_n48133_,
    new_n48134_, new_n48135_, new_n48136_, new_n48137_, new_n48138_,
    new_n48139_, new_n48140_, new_n48141_, new_n48142_, new_n48143_,
    new_n48144_, new_n48145_, new_n48146_, new_n48147_, new_n48148_,
    new_n48149_, new_n48150_, new_n48151_, new_n48152_, new_n48153_,
    new_n48154_, new_n48155_, new_n48156_, new_n48157_, new_n48158_,
    new_n48159_, new_n48160_, new_n48161_, new_n48162_, new_n48163_,
    new_n48164_, new_n48165_, new_n48166_, new_n48168_, new_n48169_,
    new_n48170_, new_n48171_, new_n48172_, new_n48173_, new_n48174_,
    new_n48175_, new_n48176_, new_n48177_, new_n48178_, new_n48179_,
    new_n48180_, new_n48181_, new_n48182_, new_n48183_, new_n48184_,
    new_n48185_, new_n48186_, new_n48187_, new_n48188_, new_n48189_,
    new_n48190_, new_n48191_, new_n48192_, new_n48193_, new_n48194_,
    new_n48195_, new_n48196_, new_n48197_, new_n48198_, new_n48199_,
    new_n48200_, new_n48202_, new_n48203_, new_n48204_, new_n48205_,
    new_n48206_, new_n48207_, new_n48208_, new_n48209_, new_n48210_,
    new_n48211_, new_n48212_, new_n48213_, new_n48214_, new_n48215_,
    new_n48216_, new_n48217_, new_n48218_, new_n48219_, new_n48220_,
    new_n48221_, new_n48222_, new_n48223_, new_n48224_, new_n48225_,
    new_n48226_, new_n48227_, new_n48228_, new_n48229_, new_n48230_,
    new_n48231_, new_n48232_, new_n48233_, new_n48234_, new_n48235_,
    new_n48237_, new_n48238_, new_n48239_, new_n48240_, new_n48241_,
    new_n48242_, new_n48243_, new_n48244_, new_n48245_, new_n48246_,
    new_n48247_, new_n48248_, new_n48249_, new_n48250_, new_n48251_,
    new_n48252_, new_n48253_, new_n48254_, new_n48255_, new_n48256_,
    new_n48257_, new_n48258_, new_n48259_, new_n48260_, new_n48261_,
    new_n48262_, new_n48263_, new_n48264_, new_n48265_, new_n48266_,
    new_n48267_, new_n48268_, new_n48269_, new_n48270_, new_n48271_,
    new_n48272_, new_n48273_, new_n48274_, new_n48275_, new_n48276_,
    new_n48277_, new_n48278_, new_n48279_, new_n48280_, new_n48281_,
    new_n48282_, new_n48283_, new_n48284_, new_n48285_, new_n48286_,
    new_n48287_, new_n48288_, new_n48289_, new_n48290_, new_n48291_,
    new_n48293_, new_n48294_, new_n48295_, new_n48296_, new_n48297_,
    new_n48298_, new_n48299_, new_n48300_, new_n48301_, new_n48302_,
    new_n48303_, new_n48304_, new_n48305_, new_n48306_, new_n48307_,
    new_n48308_, new_n48309_, new_n48310_, new_n48311_, new_n48312_,
    new_n48313_, new_n48314_, new_n48315_, new_n48316_, new_n48317_,
    new_n48318_, new_n48319_, new_n48320_, new_n48321_, new_n48322_,
    new_n48323_, new_n48324_, new_n48325_, new_n48326_, new_n48328_,
    new_n48329_, new_n48330_, new_n48332_, new_n48333_, new_n48334_,
    new_n48336_, new_n48337_, new_n48338_, new_n48340_, new_n48341_,
    new_n48342_, new_n48344_, new_n48345_, new_n48346_, new_n48348_,
    new_n48349_, new_n48350_, new_n48352_, new_n48353_, new_n48354_,
    new_n48356_, new_n48357_, new_n48358_, new_n48360_, new_n48361_,
    new_n48362_, new_n48363_, new_n48364_, new_n48365_, new_n48366_,
    new_n48367_, new_n48368_, new_n48369_, new_n48370_, new_n48371_,
    new_n48372_, new_n48373_, new_n48374_, new_n48375_, new_n48377_,
    new_n48378_, new_n48379_, new_n48381_, new_n48382_, new_n48383_,
    new_n48384_, new_n48385_, new_n48386_, new_n48387_, new_n48388_,
    new_n48389_, new_n48390_, new_n48391_, new_n48392_, new_n48393_,
    new_n48394_, new_n48395_, new_n48396_, new_n48397_, new_n48398_,
    new_n48399_, new_n48400_, new_n48401_, new_n48402_, new_n48403_,
    new_n48404_, new_n48405_, new_n48406_, new_n48407_, new_n48408_,
    new_n48409_, new_n48410_, new_n48411_, new_n48412_, new_n48413_,
    new_n48414_, new_n48415_, new_n48417_, new_n48418_, new_n48419_,
    new_n48421_, new_n48422_, new_n48423_, new_n48425_, new_n48426_,
    new_n48427_, new_n48429_, new_n48430_, new_n48431_, new_n48433_,
    new_n48434_, new_n48435_, new_n48437_, new_n48438_, new_n48440_,
    new_n48441_, new_n48442_, new_n48444_, new_n48445_, new_n48446_,
    new_n48448_, new_n48449_, new_n48450_, new_n48452_, new_n48453_,
    new_n48454_, new_n48456_, new_n48457_, new_n48458_, new_n48460_,
    new_n48461_, new_n48462_, new_n48464_, new_n48465_, new_n48466_,
    new_n48468_, new_n48469_, new_n48470_, new_n48471_, new_n48472_,
    new_n48473_, new_n48474_, new_n48475_, new_n48476_, new_n48477_,
    new_n48478_, new_n48479_, new_n48481_, new_n48482_, new_n48483_,
    new_n48485_, new_n48486_, new_n48487_, new_n48489_, new_n48490_,
    new_n48491_, new_n48493_, new_n48494_, new_n48495_, new_n48497_,
    new_n48498_, new_n48499_, new_n48501_, new_n48502_, new_n48503_,
    new_n48505_, new_n48506_, new_n48507_, new_n48509_, new_n48510_,
    new_n48511_, new_n48513_, new_n48514_, new_n48515_, new_n48517_,
    new_n48518_, new_n48519_, new_n48521_, new_n48522_, new_n48523_,
    new_n48525_, new_n48526_, new_n48527_, new_n48529_, new_n48530_,
    new_n48531_, new_n48533_, new_n48534_, new_n48535_, new_n48537_,
    new_n48538_, new_n48539_, new_n48541_, new_n48542_, new_n48543_,
    new_n48545_, new_n48546_, new_n48547_, new_n48550_, new_n48551_,
    new_n48552_, new_n48553_, new_n48554_, new_n48555_, new_n48556_,
    new_n48557_, new_n48558_, new_n48559_, new_n48560_, new_n48561_,
    new_n48562_, new_n48563_, new_n48564_, new_n48565_, new_n48566_,
    new_n48567_, new_n48568_, new_n48569_, new_n48570_, new_n48571_,
    new_n48573_, new_n48574_, new_n48575_, new_n48577_, new_n48578_,
    new_n48579_, new_n48581_, new_n48582_, new_n48583_, new_n48585_,
    new_n48586_, new_n48587_, new_n48588_, new_n48589_, new_n48590_,
    new_n48591_, new_n48592_, new_n48593_, new_n48594_, new_n48595_,
    new_n48596_, new_n48597_, new_n48598_, new_n48599_, new_n48600_,
    new_n48602_, new_n48603_, new_n48604_, new_n48606_, new_n48607_,
    new_n48608_, new_n48609_, new_n48611_, new_n48612_, new_n48613_,
    new_n48614_, new_n48616_, new_n48617_, new_n48618_, new_n48620_,
    new_n48621_, new_n48622_, new_n48623_, new_n48624_, new_n48625_,
    new_n48626_, new_n48628_, new_n48629_, new_n48630_, new_n48632_,
    new_n48633_, new_n48634_, new_n48635_, new_n48636_, new_n48637_,
    new_n48638_, new_n48639_, new_n48640_, new_n48641_, new_n48642_,
    new_n48643_, new_n48644_, new_n48645_, new_n48646_, new_n48647_,
    new_n48649_, new_n48650_, new_n48651_, new_n48653_, new_n48654_,
    new_n48655_, new_n48657_, new_n48658_, new_n48659_, new_n48660_,
    new_n48661_, new_n48662_, new_n48663_, new_n48667_, new_n48668_,
    new_n48670_, new_n48672_, new_n48673_, new_n48675_, new_n48676_,
    new_n48678_, new_n48679_, new_n48681_, new_n48682_, new_n48684_,
    new_n48685_, new_n48687_, new_n48688_, new_n48690_, new_n48691_,
    new_n48693_, new_n48694_, new_n48696_, new_n48697_, new_n48699_,
    new_n48700_, new_n48702_, new_n48703_, new_n48704_, new_n48706_,
    new_n48707_, new_n48709_, new_n48710_, new_n48711_, new_n48712_,
    new_n48713_, new_n48714_, new_n48715_, new_n48716_, new_n48718_,
    new_n48719_, new_n48721_, new_n48722_, new_n48724_, new_n48725_,
    new_n48727_, new_n48728_, new_n48730_, new_n48731_, new_n48733_,
    new_n48734_, new_n48736_, new_n48737_, new_n48738_, new_n48740_,
    new_n48741_, new_n48743_, new_n48744_, new_n48746_, new_n48747_,
    new_n48749_, new_n48750_, new_n48752_, new_n48753_, new_n48755_,
    new_n48756_, new_n48758_, new_n48759_, new_n48761_, new_n48762_,
    new_n48764_, new_n48765_, new_n48767_, new_n48768_, new_n48770_,
    new_n48772_, new_n48774_, new_n48776_, new_n48779_, new_n48780_,
    new_n48781_, new_n48783_, new_n48784_, new_n48785_, new_n48786_,
    new_n48787_, new_n48788_, new_n48789_, new_n48790_, new_n48791_,
    new_n48792_, new_n48793_, new_n48794_, new_n48795_, new_n48796_,
    new_n48797_, new_n48798_, new_n48799_, new_n48800_, new_n48801_,
    new_n48802_, new_n48803_, new_n48804_, new_n48805_, new_n48806_,
    new_n48807_, new_n48808_, new_n48809_, new_n48810_, new_n48812_,
    new_n48813_, new_n48814_, new_n48815_, new_n48816_, new_n48817_,
    new_n48818_, new_n48819_, new_n48820_, new_n48821_, new_n48822_,
    new_n48823_, new_n48824_, new_n48825_, new_n48826_, new_n48827_,
    new_n48828_, new_n48829_, new_n48830_, new_n48831_, new_n48832_,
    new_n48833_, new_n48834_, new_n48835_, new_n48836_, new_n48837_,
    new_n48838_, new_n48840_, new_n48841_, new_n48842_, new_n48843_,
    new_n48844_, new_n48845_, new_n48846_, new_n48847_, new_n48848_,
    new_n48849_, new_n48850_, new_n48851_, new_n48852_, new_n48853_,
    new_n48854_, new_n48855_, new_n48856_, new_n48857_, new_n48858_,
    new_n48859_, new_n48860_, new_n48861_, new_n48862_, new_n48863_,
    new_n48864_, new_n48865_, new_n48866_, new_n48868_, new_n48869_,
    new_n48870_, new_n48871_, new_n48872_, new_n48873_, new_n48874_,
    new_n48875_, new_n48876_, new_n48877_, new_n48878_, new_n48879_,
    new_n48880_, new_n48881_, new_n48882_, new_n48883_, new_n48884_,
    new_n48885_, new_n48886_, new_n48887_, new_n48888_, new_n48889_,
    new_n48890_, new_n48891_, new_n48892_, new_n48893_, new_n48894_,
    new_n48896_, new_n48897_, new_n48899_, new_n48901_, new_n48902_,
    new_n48904_, new_n48907_, new_n48909_, new_n48910_, new_n48912_,
    new_n48913_, new_n48915_, new_n48916_, new_n48918_, new_n48919_,
    new_n48922_, new_n48923_, new_n48925_, new_n48926_, new_n48928_,
    new_n48929_, new_n48931_, new_n48932_, new_n48934_, new_n48935_,
    new_n48937_, new_n48938_, new_n48940_, new_n48941_, new_n48943_,
    new_n48944_, new_n48946_, new_n48947_, new_n48949_, new_n48950_,
    new_n48952_, new_n48953_, new_n48955_, new_n48956_, new_n48958_,
    new_n48959_, new_n48961_, new_n48962_, new_n48964_, new_n48965_,
    new_n48967_, new_n48968_, new_n48970_, new_n48971_, new_n48973_,
    new_n48974_, new_n48976_, new_n48977_, new_n48979_, new_n48980_,
    new_n48981_, new_n48982_, new_n48983_, new_n48984_, new_n48985_,
    new_n48986_, new_n48988_, new_n48989_, new_n48991_, new_n48992_,
    new_n48994_, new_n48995_, new_n48997_, new_n48998_, new_n49000_,
    new_n49001_, new_n49003_, new_n49004_, new_n49006_, new_n49007_,
    new_n49009_, new_n49010_, new_n49011_, new_n49012_, new_n49013_,
    new_n49014_, new_n49015_, new_n49016_, new_n49018_, new_n49019_,
    new_n49021_, new_n49022_, new_n49024_, new_n49025_, new_n49027_,
    new_n49028_, new_n49030_, new_n49031_, new_n49033_, new_n49034_,
    new_n49035_, new_n49036_, new_n49037_, new_n49038_, new_n49039_,
    new_n49040_, new_n49042_, new_n49043_, new_n49045_, new_n49046_,
    new_n49047_, new_n49048_, new_n49049_, new_n49050_, new_n49051_,
    new_n49052_, new_n49054_, new_n49055_, new_n49056_, new_n49057_,
    new_n49058_, new_n49059_, new_n49060_, new_n49061_, new_n49063_,
    new_n49064_, new_n49065_, new_n49066_, new_n49067_, new_n49068_,
    new_n49069_, new_n49070_, new_n49072_, new_n49073_, new_n49075_,
    new_n49076_, new_n49078_, new_n49080_, new_n49081_, new_n49083_,
    new_n49084_, new_n49086_, new_n49087_, new_n49089_, new_n49091_,
    new_n49092_, new_n49094_, new_n49095_, new_n49097_, new_n49098_,
    new_n49100_, new_n49101_, new_n49103_, new_n49104_, new_n49106_,
    new_n49107_, new_n49109_, new_n49110_, new_n49112_, new_n49113_,
    new_n49115_, new_n49116_, new_n49118_, new_n49120_, new_n49121_,
    new_n49123_, new_n49124_, new_n49126_, new_n49127_, new_n49129_,
    new_n49131_, new_n49133_, new_n49134_, new_n49136_, new_n49137_,
    new_n49138_, new_n49139_, new_n49140_, new_n49141_, new_n49142_,
    new_n49143_, new_n49144_, new_n49145_, new_n49147_, new_n49149_,
    new_n49150_, new_n49152_, new_n49153_, new_n49155_, new_n49156_,
    new_n49158_, new_n49160_, new_n49161_, new_n49163_, new_n49165_,
    new_n49166_, new_n49168_, new_n49170_, new_n49171_, new_n49173_,
    new_n49174_, new_n49176_, new_n49177_, new_n49179_, new_n49180_,
    new_n49182_, new_n49184_, new_n49185_, new_n49187_, new_n49188_,
    new_n49190_, new_n49191_, new_n49193_, new_n49194_, new_n49196_,
    new_n49197_, new_n49199_, new_n49200_, new_n49202_, new_n49204_,
    new_n49205_, new_n49207_, new_n49208_, new_n49210_, new_n49211_,
    new_n49213_, new_n49215_, new_n49217_, new_n49218_, new_n49220_,
    new_n49222_, new_n49223_, new_n49225_, new_n49226_, new_n49228_,
    new_n49230_, new_n49231_, new_n49233_, new_n49235_, new_n49236_,
    new_n49238_, new_n49239_, new_n49241_, new_n49242_, new_n49244_,
    new_n49245_, new_n49248_, new_n49250_, new_n49252_, new_n49253_,
    new_n49256_;
  assign new_n2437_ = ~pi0216 & pi0833;
  assign new_n2438_ = pi0929 & new_n2437_;
  assign new_n2439_ = pi1144 & ~new_n2437_;
  assign new_n2440_ = ~pi0332 & ~new_n2439_;
  assign new_n2441_ = ~new_n2438_ & new_n2440_;
  assign new_n2442_ = pi0221 & ~new_n2441_;
  assign new_n2443_ = pi0265 & ~pi0332;
  assign new_n2444_ = pi0216 & ~new_n2443_;
  assign new_n2445_ = pi0153 & ~pi0332;
  assign new_n2446_ = ~pi0105 & ~new_n2445_;
  assign new_n2447_ = ~pi0152 & ~pi0161;
  assign new_n2448_ = ~pi0166 & new_n2447_;
  assign new_n2449_ = pi0095 & ~pi0479;
  assign new_n2450_ = ~pi0040 & ~pi0072;
  assign new_n2451_ = ~pi0088 & ~pi0098;
  assign new_n2452_ = ~pi0077 & new_n2451_;
  assign new_n2453_ = ~pi0050 & new_n2452_;
  assign new_n2454_ = ~pi0102 & new_n2453_;
  assign new_n2455_ = ~pi0065 & ~pi0071;
  assign new_n2456_ = ~pi0083 & ~pi0103;
  assign new_n2457_ = ~pi0067 & ~pi0069;
  assign new_n2458_ = ~pi0066 & ~pi0073;
  assign new_n2459_ = ~pi0061 & ~pi0076;
  assign new_n2460_ = ~pi0085 & ~pi0106;
  assign new_n2461_ = new_n2459_ & new_n2460_;
  assign new_n2462_ = ~pi0048 & new_n2461_;
  assign new_n2463_ = ~pi0089 & new_n2462_;
  assign new_n2464_ = ~pi0049 & new_n2463_;
  assign new_n2465_ = ~pi0104 & new_n2464_;
  assign new_n2466_ = ~pi0045 & new_n2465_;
  assign new_n2467_ = ~pi0068 & ~pi0084;
  assign new_n2468_ = ~pi0082 & ~pi0111;
  assign new_n2469_ = ~pi0036 & new_n2468_;
  assign new_n2470_ = new_n2467_ & new_n2469_;
  assign new_n2471_ = new_n2466_ & new_n2470_;
  assign new_n2472_ = new_n2458_ & new_n2471_;
  assign new_n2473_ = new_n2457_ & new_n2472_;
  assign new_n2474_ = new_n2456_ & new_n2473_;
  assign new_n2475_ = new_n2455_ & new_n2474_;
  assign new_n2476_ = ~pi0063 & ~pi0107;
  assign new_n2477_ = new_n2475_ & new_n2476_;
  assign new_n2478_ = ~pi0064 & new_n2477_;
  assign new_n2479_ = ~pi0081 & new_n2478_;
  assign new_n2480_ = new_n2454_ & new_n2479_;
  assign new_n2481_ = ~pi0097 & ~pi0108;
  assign new_n2482_ = ~pi0094 & new_n2481_;
  assign new_n2483_ = ~pi0053 & ~pi0060;
  assign new_n2484_ = ~pi0086 & new_n2483_;
  assign new_n2485_ = ~pi0046 & new_n2484_;
  assign new_n2486_ = new_n2482_ & new_n2485_;
  assign new_n2487_ = new_n2480_ & new_n2486_;
  assign new_n2488_ = ~pi0109 & ~pi0110;
  assign new_n2489_ = ~pi0058 & ~pi0091;
  assign new_n2490_ = ~pi0047 & new_n2489_;
  assign new_n2491_ = new_n2488_ & new_n2490_;
  assign new_n2492_ = new_n2487_ & new_n2491_;
  assign new_n2493_ = ~pi0090 & ~pi0093;
  assign new_n2494_ = ~pi0070 & ~pi0096;
  assign new_n2495_ = ~pi0035 & ~pi0051;
  assign new_n2496_ = new_n2494_ & new_n2495_;
  assign new_n2497_ = new_n2493_ & new_n2496_;
  assign new_n2498_ = new_n2492_ & new_n2497_;
  assign new_n2499_ = new_n2450_ & new_n2498_;
  assign new_n2500_ = pi0225 & new_n2499_;
  assign new_n2501_ = pi0032 & ~new_n2500_;
  assign new_n2502_ = ~pi0095 & ~new_n2501_;
  assign new_n2503_ = pi0060 & new_n2480_;
  assign new_n2504_ = ~pi0053 & ~new_n2503_;
  assign new_n2505_ = ~pi0086 & ~pi0094;
  assign new_n2506_ = ~pi0060 & new_n2480_;
  assign new_n2507_ = pi0053 & ~new_n2506_;
  assign new_n2508_ = new_n2505_ & ~new_n2507_;
  assign new_n2509_ = ~new_n2504_ & new_n2508_;
  assign new_n2510_ = ~pi0046 & new_n2488_;
  assign new_n2511_ = ~pi0047 & ~pi0091;
  assign new_n2512_ = new_n2481_ & new_n2511_;
  assign new_n2513_ = new_n2510_ & new_n2512_;
  assign new_n2514_ = ~pi0058 & new_n2513_;
  assign new_n2515_ = new_n2493_ & new_n2514_;
  assign new_n2516_ = new_n2509_ & new_n2515_;
  assign new_n2517_ = ~pi0035 & ~new_n2516_;
  assign new_n2518_ = ~pi0058 & ~pi0090;
  assign new_n2519_ = new_n2486_ & new_n2488_;
  assign new_n2520_ = new_n2511_ & new_n2519_;
  assign new_n2521_ = new_n2480_ & new_n2520_;
  assign new_n2522_ = new_n2518_ & new_n2521_;
  assign new_n2523_ = ~pi0093 & new_n2522_;
  assign new_n2524_ = pi0035 & ~new_n2523_;
  assign new_n2525_ = pi0035 & new_n2523_;
  assign new_n2526_ = ~pi0225 & new_n2525_;
  assign new_n2527_ = ~pi0070 & ~new_n2526_;
  assign new_n2528_ = ~pi0051 & new_n2527_;
  assign new_n2529_ = ~new_n2524_ & new_n2528_;
  assign new_n2530_ = ~new_n2517_ & new_n2529_;
  assign new_n2531_ = ~pi0096 & ~new_n2530_;
  assign new_n2532_ = ~pi0047 & new_n2519_;
  assign new_n2533_ = new_n2480_ & new_n2532_;
  assign new_n2534_ = ~pi0035 & ~pi0070;
  assign new_n2535_ = ~pi0051 & new_n2534_;
  assign new_n2536_ = ~pi0093 & new_n2518_;
  assign new_n2537_ = ~pi0091 & new_n2536_;
  assign new_n2538_ = new_n2535_ & new_n2537_;
  assign new_n2539_ = new_n2533_ & new_n2538_;
  assign new_n2540_ = pi0096 & ~new_n2539_;
  assign new_n2541_ = new_n2450_ & ~new_n2540_;
  assign new_n2542_ = ~new_n2531_ & new_n2541_;
  assign new_n2543_ = ~pi0032 & ~new_n2542_;
  assign new_n2544_ = new_n2502_ & ~new_n2543_;
  assign new_n2545_ = ~new_n2449_ & ~new_n2544_;
  assign new_n2546_ = ~pi0137 & new_n2545_;
  assign new_n2547_ = ~pi0035 & ~pi0093;
  assign new_n2548_ = new_n2522_ & new_n2547_;
  assign new_n2549_ = ~pi0072 & ~pi0096;
  assign new_n2550_ = ~pi0051 & ~pi0070;
  assign new_n2551_ = new_n2549_ & new_n2550_;
  assign new_n2552_ = new_n2548_ & new_n2551_;
  assign new_n2553_ = pi0040 & new_n2552_;
  assign new_n2554_ = ~pi0032 & ~new_n2553_;
  assign new_n2555_ = pi0072 & ~new_n2498_;
  assign new_n2556_ = ~pi0040 & ~new_n2555_;
  assign new_n2557_ = ~pi0070 & new_n2548_;
  assign new_n2558_ = pi0051 & ~new_n2557_;
  assign new_n2559_ = ~pi0096 & ~new_n2558_;
  assign new_n2560_ = ~pi0051 & pi0070;
  assign new_n2561_ = new_n2559_ & ~new_n2560_;
  assign new_n2562_ = ~new_n2524_ & ~new_n2526_;
  assign new_n2563_ = pi0093 & new_n2522_;
  assign new_n2564_ = ~pi0035 & ~new_n2563_;
  assign new_n2565_ = pi0091 & new_n2533_;
  assign new_n2566_ = new_n2518_ & ~new_n2565_;
  assign new_n2567_ = ~pi0109 & new_n2487_;
  assign new_n2568_ = pi0110 & ~new_n2567_;
  assign new_n2569_ = pi0047 & new_n2480_;
  assign new_n2570_ = new_n2519_ & new_n2569_;
  assign new_n2571_ = pi0047 & ~new_n2570_;
  assign new_n2572_ = ~pi0091 & ~new_n2571_;
  assign new_n2573_ = ~new_n2568_ & new_n2572_;
  assign new_n2574_ = ~pi0047 & ~pi0110;
  assign new_n2575_ = pi0109 & ~new_n2487_;
  assign new_n2576_ = ~pi0102 & new_n2479_;
  assign new_n2577_ = new_n2451_ & new_n2576_;
  assign new_n2578_ = ~pi0050 & new_n2483_;
  assign new_n2579_ = ~pi0077 & new_n2578_;
  assign new_n2580_ = new_n2505_ & new_n2579_;
  assign new_n2581_ = new_n2577_ & new_n2580_;
  assign new_n2582_ = ~pi0097 & new_n2581_;
  assign new_n2583_ = pi0108 & ~new_n2582_;
  assign new_n2584_ = ~pi0046 & ~new_n2583_;
  assign new_n2585_ = pi0097 & ~new_n2581_;
  assign new_n2586_ = new_n2452_ & new_n2576_;
  assign new_n2587_ = new_n2578_ & new_n2586_;
  assign new_n2588_ = ~pi0086 & pi0094;
  assign new_n2589_ = new_n2587_ & new_n2588_;
  assign new_n2590_ = ~pi0097 & ~new_n2589_;
  assign new_n2591_ = pi0086 & ~new_n2587_;
  assign new_n2592_ = ~pi0094 & ~new_n2591_;
  assign new_n2593_ = pi0077 & new_n2577_;
  assign new_n2594_ = ~pi0050 & ~new_n2593_;
  assign new_n2595_ = pi0081 & ~new_n2478_;
  assign new_n2596_ = pi0102 & ~new_n2479_;
  assign new_n2597_ = ~new_n2595_ & ~new_n2596_;
  assign new_n2598_ = pi0064 & ~new_n2477_;
  assign new_n2599_ = pi0071 & ~new_n2474_;
  assign new_n2600_ = ~pi0065 & ~new_n2599_;
  assign new_n2601_ = ~pi0067 & new_n2472_;
  assign new_n2602_ = pi0069 & ~new_n2601_;
  assign new_n2603_ = pi0083 & ~new_n2473_;
  assign new_n2604_ = ~pi0103 & ~new_n2603_;
  assign new_n2605_ = ~new_n2602_ & new_n2604_;
  assign new_n2606_ = ~pi0069 & ~pi0083;
  assign new_n2607_ = ~pi0068 & ~pi0111;
  assign new_n2608_ = new_n2458_ & new_n2466_;
  assign new_n2609_ = pi0084 & ~new_n2608_;
  assign new_n2610_ = pi0085 & pi0106;
  assign new_n2611_ = new_n2459_ & ~new_n2610_;
  assign new_n2612_ = pi0061 & pi0076;
  assign new_n2613_ = new_n2460_ & ~new_n2612_;
  assign new_n2614_ = ~new_n2611_ & ~new_n2613_;
  assign new_n2615_ = ~pi0048 & ~new_n2614_;
  assign new_n2616_ = ~new_n2461_ & ~new_n2615_;
  assign new_n2617_ = pi0089 & ~new_n2462_;
  assign new_n2618_ = ~pi0049 & ~new_n2617_;
  assign new_n2619_ = ~new_n2616_ & new_n2618_;
  assign new_n2620_ = ~new_n2463_ & ~new_n2619_;
  assign new_n2621_ = pi0104 & ~new_n2464_;
  assign new_n2622_ = ~pi0045 & ~new_n2621_;
  assign new_n2623_ = ~new_n2620_ & new_n2622_;
  assign new_n2624_ = ~new_n2465_ & ~new_n2623_;
  assign new_n2625_ = ~new_n2466_ & ~new_n2624_;
  assign new_n2626_ = new_n2458_ & ~new_n2625_;
  assign new_n2627_ = pi0066 & pi0073;
  assign new_n2628_ = ~new_n2458_ & ~new_n2466_;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = ~new_n2626_ & new_n2629_;
  assign new_n2631_ = ~pi0084 & ~new_n2630_;
  assign new_n2632_ = ~new_n2609_ & ~new_n2631_;
  assign new_n2633_ = new_n2607_ & ~new_n2632_;
  assign new_n2634_ = ~pi0084 & new_n2608_;
  assign new_n2635_ = ~pi0068 & new_n2634_;
  assign new_n2636_ = pi0111 & ~new_n2635_;
  assign new_n2637_ = ~pi0082 & ~new_n2636_;
  assign new_n2638_ = pi0068 & ~new_n2634_;
  assign new_n2639_ = new_n2637_ & ~new_n2638_;
  assign new_n2640_ = ~new_n2633_ & new_n2639_;
  assign new_n2641_ = ~pi0036 & ~pi0067;
  assign new_n2642_ = pi0082 & new_n2607_;
  assign new_n2643_ = new_n2634_ & new_n2642_;
  assign new_n2644_ = new_n2641_ & ~new_n2643_;
  assign new_n2645_ = ~new_n2640_ & new_n2644_;
  assign new_n2646_ = pi0067 & ~new_n2472_;
  assign new_n2647_ = new_n2468_ & new_n2635_;
  assign new_n2648_ = pi0036 & ~new_n2647_;
  assign new_n2649_ = ~new_n2646_ & ~new_n2648_;
  assign new_n2650_ = ~new_n2645_ & new_n2649_;
  assign new_n2651_ = new_n2606_ & ~new_n2650_;
  assign new_n2652_ = new_n2605_ & ~new_n2651_;
  assign new_n2653_ = pi0103 & new_n2606_;
  assign new_n2654_ = new_n2601_ & new_n2653_;
  assign new_n2655_ = ~pi0071 & ~new_n2654_;
  assign new_n2656_ = ~new_n2652_ & new_n2655_;
  assign new_n2657_ = new_n2600_ & ~new_n2656_;
  assign new_n2658_ = ~pi0107 & ~new_n2657_;
  assign new_n2659_ = pi0065 & ~pi0071;
  assign new_n2660_ = new_n2474_ & new_n2659_;
  assign new_n2661_ = new_n2658_ & ~new_n2660_;
  assign new_n2662_ = pi0107 & ~new_n2475_;
  assign new_n2663_ = ~pi0063 & ~new_n2662_;
  assign new_n2664_ = ~new_n2661_ & new_n2663_;
  assign new_n2665_ = ~pi0064 & ~new_n2664_;
  assign new_n2666_ = ~new_n2598_ & ~new_n2665_;
  assign new_n2667_ = ~pi0081 & ~pi0102;
  assign new_n2668_ = ~new_n2666_ & new_n2667_;
  assign new_n2669_ = ~new_n2658_ & new_n2663_;
  assign new_n2670_ = pi0063 & ~pi0107;
  assign new_n2671_ = new_n2475_ & new_n2670_;
  assign new_n2672_ = ~pi0064 & ~new_n2671_;
  assign new_n2673_ = ~new_n2669_ & new_n2672_;
  assign new_n2674_ = ~new_n2598_ & ~new_n2673_;
  assign new_n2675_ = new_n2668_ & ~new_n2674_;
  assign new_n2676_ = new_n2597_ & ~new_n2675_;
  assign new_n2677_ = new_n2451_ & ~new_n2676_;
  assign new_n2678_ = ~pi0098 & new_n2576_;
  assign new_n2679_ = pi0088 & ~new_n2678_;
  assign new_n2680_ = pi0098 & ~new_n2576_;
  assign new_n2681_ = ~pi0077 & ~new_n2680_;
  assign new_n2682_ = ~new_n2679_ & new_n2681_;
  assign new_n2683_ = ~new_n2677_ & new_n2682_;
  assign new_n2684_ = new_n2594_ & ~new_n2683_;
  assign new_n2685_ = pi0050 & ~new_n2586_;
  assign new_n2686_ = ~pi0060 & ~new_n2685_;
  assign new_n2687_ = ~new_n2684_ & new_n2686_;
  assign new_n2688_ = new_n2504_ & ~new_n2687_;
  assign new_n2689_ = ~new_n2507_ & ~new_n2688_;
  assign new_n2690_ = ~pi0086 & ~new_n2689_;
  assign new_n2691_ = new_n2592_ & ~new_n2690_;
  assign new_n2692_ = new_n2590_ & ~new_n2691_;
  assign new_n2693_ = ~new_n2585_ & ~new_n2692_;
  assign new_n2694_ = ~pi0108 & ~new_n2693_;
  assign new_n2695_ = new_n2584_ & ~new_n2694_;
  assign new_n2696_ = pi0046 & new_n2481_;
  assign new_n2697_ = new_n2581_ & new_n2696_;
  assign new_n2698_ = ~pi0109 & ~new_n2697_;
  assign new_n2699_ = ~new_n2695_ & new_n2698_;
  assign new_n2700_ = ~new_n2575_ & ~new_n2699_;
  assign new_n2701_ = new_n2574_ & ~new_n2700_;
  assign new_n2702_ = new_n2573_ & ~new_n2701_;
  assign new_n2703_ = new_n2566_ & ~new_n2702_;
  assign new_n2704_ = pi0058 & ~new_n2521_;
  assign new_n2705_ = pi0090 & ~new_n2492_;
  assign new_n2706_ = ~pi0093 & ~new_n2705_;
  assign new_n2707_ = ~new_n2704_ & new_n2706_;
  assign new_n2708_ = ~new_n2703_ & new_n2707_;
  assign new_n2709_ = new_n2564_ & ~new_n2708_;
  assign new_n2710_ = new_n2562_ & ~new_n2709_;
  assign new_n2711_ = ~pi0051 & ~new_n2710_;
  assign new_n2712_ = new_n2561_ & ~new_n2711_;
  assign new_n2713_ = ~pi0072 & ~new_n2712_;
  assign new_n2714_ = new_n2556_ & ~new_n2713_;
  assign new_n2715_ = new_n2554_ & ~new_n2714_;
  assign new_n2716_ = pi0096 & new_n2539_;
  assign new_n2717_ = ~pi0051 & ~pi0072;
  assign new_n2718_ = ~pi0040 & new_n2717_;
  assign new_n2719_ = new_n2548_ & new_n2718_;
  assign new_n2720_ = new_n2716_ & new_n2719_;
  assign new_n2721_ = new_n2715_ & ~new_n2720_;
  assign new_n2722_ = ~new_n2501_ & ~new_n2721_;
  assign new_n2723_ = ~pi0095 & ~new_n2722_;
  assign new_n2724_ = ~pi0032 & ~pi0040;
  assign new_n2725_ = new_n2552_ & new_n2724_;
  assign new_n2726_ = pi0095 & ~new_n2725_;
  assign new_n2727_ = pi0479 & new_n2726_;
  assign new_n2728_ = ~new_n2723_ & ~new_n2727_;
  assign new_n2729_ = pi0137 & ~new_n2728_;
  assign new_n2730_ = ~new_n2546_ & ~new_n2729_;
  assign new_n2731_ = pi0210 & ~new_n2730_;
  assign new_n2732_ = ~pi0833 & pi0957;
  assign new_n2733_ = pi1091 & ~new_n2732_;
  assign new_n2734_ = pi0841 & new_n2522_;
  assign new_n2735_ = ~pi0093 & new_n2734_;
  assign new_n2736_ = new_n2717_ & new_n2735_;
  assign new_n2737_ = ~pi0035 & ~pi0040;
  assign new_n2738_ = pi0225 & new_n2737_;
  assign new_n2739_ = new_n2494_ & new_n2738_;
  assign new_n2740_ = new_n2736_ & new_n2739_;
  assign new_n2741_ = pi0032 & ~new_n2740_;
  assign new_n2742_ = ~new_n2721_ & ~new_n2741_;
  assign new_n2743_ = ~pi0095 & ~new_n2742_;
  assign new_n2744_ = ~new_n2727_ & ~new_n2743_;
  assign new_n2745_ = pi0137 & ~new_n2744_;
  assign new_n2746_ = pi0095 & pi0479;
  assign new_n2747_ = ~new_n2543_ & ~new_n2741_;
  assign new_n2748_ = ~pi0095 & ~new_n2747_;
  assign new_n2749_ = ~new_n2746_ & ~new_n2748_;
  assign new_n2750_ = ~pi0137 & ~new_n2749_;
  assign new_n2751_ = ~new_n2745_ & ~new_n2750_;
  assign new_n2752_ = ~new_n2733_ & new_n2751_;
  assign new_n2753_ = pi0829 & pi0950;
  assign new_n2754_ = pi1092 & pi1093;
  assign new_n2755_ = new_n2753_ & new_n2754_;
  assign new_n2756_ = new_n2749_ & ~new_n2755_;
  assign new_n2757_ = ~pi0097 & ~new_n2509_;
  assign new_n2758_ = ~pi0108 & ~new_n2585_;
  assign new_n2759_ = ~pi0110 & new_n2758_;
  assign new_n2760_ = ~pi0046 & ~pi0109;
  assign new_n2761_ = new_n2511_ & new_n2760_;
  assign new_n2762_ = new_n2536_ & new_n2761_;
  assign new_n2763_ = new_n2759_ & new_n2762_;
  assign new_n2764_ = ~new_n2757_ & new_n2763_;
  assign new_n2765_ = ~pi0035 & ~new_n2764_;
  assign new_n2766_ = new_n2529_ & ~new_n2765_;
  assign new_n2767_ = ~pi0096 & ~new_n2766_;
  assign new_n2768_ = new_n2541_ & ~new_n2767_;
  assign new_n2769_ = ~pi0032 & ~new_n2768_;
  assign new_n2770_ = ~new_n2741_ & ~new_n2769_;
  assign new_n2771_ = ~pi0095 & ~new_n2770_;
  assign new_n2772_ = ~new_n2746_ & new_n2755_;
  assign new_n2773_ = ~new_n2771_ & new_n2772_;
  assign new_n2774_ = ~pi0137 & ~new_n2773_;
  assign new_n2775_ = ~new_n2756_ & new_n2774_;
  assign new_n2776_ = new_n2733_ & ~new_n2775_;
  assign new_n2777_ = ~new_n2745_ & new_n2776_;
  assign new_n2778_ = ~new_n2752_ & ~new_n2777_;
  assign new_n2779_ = ~pi0210 & new_n2778_;
  assign new_n2780_ = ~new_n2731_ & ~new_n2779_;
  assign new_n2781_ = pi0234 & new_n2780_;
  assign new_n2782_ = ~pi0040 & new_n2549_;
  assign new_n2783_ = new_n2530_ & new_n2782_;
  assign new_n2784_ = ~pi0032 & ~new_n2783_;
  assign new_n2785_ = new_n2502_ & ~new_n2784_;
  assign new_n2786_ = ~pi0137 & ~new_n2785_;
  assign new_n2787_ = ~new_n2449_ & ~new_n2726_;
  assign new_n2788_ = ~new_n2501_ & ~new_n2715_;
  assign new_n2789_ = ~pi0095 & ~new_n2788_;
  assign new_n2790_ = new_n2787_ & ~new_n2789_;
  assign new_n2791_ = pi0137 & ~new_n2790_;
  assign new_n2792_ = ~new_n2786_ & ~new_n2791_;
  assign new_n2793_ = pi0210 & ~new_n2792_;
  assign new_n2794_ = ~pi0095 & ~new_n2741_;
  assign new_n2795_ = new_n2733_ & new_n2755_;
  assign new_n2796_ = ~new_n2517_ & ~new_n2795_;
  assign new_n2797_ = pi1091 & pi1093;
  assign new_n2798_ = ~new_n2732_ & new_n2797_;
  assign new_n2799_ = pi0950 & pi1092;
  assign new_n2800_ = pi0829 & new_n2799_;
  assign new_n2801_ = new_n2798_ & new_n2800_;
  assign new_n2802_ = ~new_n2765_ & new_n2801_;
  assign new_n2803_ = ~new_n2796_ & ~new_n2802_;
  assign new_n2804_ = new_n2529_ & new_n2782_;
  assign new_n2805_ = ~new_n2803_ & new_n2804_;
  assign new_n2806_ = ~pi0032 & ~new_n2805_;
  assign new_n2807_ = new_n2794_ & ~new_n2806_;
  assign new_n2808_ = ~pi0137 & ~new_n2807_;
  assign new_n2809_ = ~new_n2715_ & ~new_n2741_;
  assign new_n2810_ = ~pi0095 & ~new_n2809_;
  assign new_n2811_ = new_n2787_ & ~new_n2810_;
  assign new_n2812_ = pi0137 & ~new_n2811_;
  assign new_n2813_ = ~new_n2808_ & ~new_n2812_;
  assign new_n2814_ = ~pi0210 & ~new_n2813_;
  assign new_n2815_ = ~new_n2793_ & ~new_n2814_;
  assign new_n2816_ = ~pi0234 & new_n2815_;
  assign new_n2817_ = ~pi0332 & ~new_n2816_;
  assign new_n2818_ = ~new_n2781_ & new_n2817_;
  assign new_n2819_ = new_n2448_ & ~new_n2818_;
  assign new_n2820_ = pi0146 & new_n2780_;
  assign new_n2821_ = pi0234 & ~pi0332;
  assign new_n2822_ = ~pi0210 & ~new_n2751_;
  assign new_n2823_ = ~pi0146 & ~new_n2731_;
  assign new_n2824_ = ~new_n2822_ & new_n2823_;
  assign new_n2825_ = new_n2821_ & ~new_n2824_;
  assign new_n2826_ = ~new_n2820_ & new_n2825_;
  assign new_n2827_ = ~new_n2784_ & new_n2794_;
  assign new_n2828_ = ~pi0137 & ~new_n2827_;
  assign new_n2829_ = ~new_n2812_ & ~new_n2828_;
  assign new_n2830_ = ~pi0210 & ~new_n2829_;
  assign new_n2831_ = ~pi0146 & ~new_n2793_;
  assign new_n2832_ = ~new_n2830_ & new_n2831_;
  assign new_n2833_ = ~pi0234 & ~pi0332;
  assign new_n2834_ = pi0146 & new_n2815_;
  assign new_n2835_ = new_n2833_ & ~new_n2834_;
  assign new_n2836_ = ~new_n2832_ & new_n2835_;
  assign new_n2837_ = ~new_n2448_ & ~new_n2836_;
  assign new_n2838_ = ~new_n2826_ & new_n2837_;
  assign new_n2839_ = ~new_n2819_ & ~new_n2838_;
  assign new_n2840_ = pi0105 & ~new_n2839_;
  assign new_n2841_ = ~new_n2446_ & ~new_n2840_;
  assign new_n2842_ = pi0228 & ~new_n2841_;
  assign new_n2843_ = pi0225 & pi0841;
  assign new_n2844_ = new_n2499_ & ~new_n2843_;
  assign new_n2845_ = pi0032 & ~new_n2844_;
  assign new_n2846_ = ~pi0095 & ~new_n2845_;
  assign new_n2847_ = ~pi0051 & ~pi0096;
  assign new_n2848_ = pi0070 & ~new_n2548_;
  assign new_n2849_ = new_n2847_ & ~new_n2848_;
  assign new_n2850_ = new_n2450_ & new_n2849_;
  assign new_n2851_ = ~new_n2527_ & new_n2850_;
  assign new_n2852_ = ~pi0032 & ~new_n2851_;
  assign new_n2853_ = new_n2846_ & ~new_n2852_;
  assign new_n2854_ = pi0137 & ~new_n2853_;
  assign new_n2855_ = pi0093 & ~new_n2522_;
  assign new_n2856_ = ~pi0035 & ~new_n2855_;
  assign new_n2857_ = ~new_n2704_ & ~new_n2705_;
  assign new_n2858_ = ~pi0053 & new_n2687_;
  assign new_n2859_ = ~pi0086 & ~new_n2858_;
  assign new_n2860_ = new_n2592_ & ~new_n2859_;
  assign new_n2861_ = new_n2590_ & ~new_n2860_;
  assign new_n2862_ = ~new_n2585_ & ~new_n2861_;
  assign new_n2863_ = ~pi0108 & ~new_n2862_;
  assign new_n2864_ = new_n2584_ & ~new_n2863_;
  assign new_n2865_ = ~pi0109 & ~new_n2864_;
  assign new_n2866_ = ~new_n2575_ & ~new_n2865_;
  assign new_n2867_ = new_n2574_ & ~new_n2866_;
  assign new_n2868_ = new_n2573_ & ~new_n2867_;
  assign new_n2869_ = new_n2566_ & ~new_n2868_;
  assign new_n2870_ = new_n2857_ & ~new_n2869_;
  assign new_n2871_ = ~pi0093 & ~new_n2870_;
  assign new_n2872_ = new_n2856_ & ~new_n2871_;
  assign new_n2873_ = new_n2528_ & ~new_n2872_;
  assign new_n2874_ = new_n2559_ & ~new_n2848_;
  assign new_n2875_ = ~new_n2873_ & new_n2874_;
  assign new_n2876_ = ~pi0072 & ~new_n2875_;
  assign new_n2877_ = new_n2556_ & ~new_n2876_;
  assign new_n2878_ = new_n2554_ & ~new_n2877_;
  assign new_n2879_ = ~new_n2795_ & new_n2878_;
  assign new_n2880_ = new_n2554_ & new_n2795_;
  assign new_n2881_ = ~pi0097 & ~new_n2861_;
  assign new_n2882_ = ~pi0108 & ~new_n2881_;
  assign new_n2883_ = new_n2584_ & ~new_n2882_;
  assign new_n2884_ = ~pi0109 & ~new_n2883_;
  assign new_n2885_ = ~new_n2575_ & ~new_n2884_;
  assign new_n2886_ = new_n2574_ & ~new_n2885_;
  assign new_n2887_ = new_n2573_ & ~new_n2886_;
  assign new_n2888_ = new_n2566_ & ~new_n2887_;
  assign new_n2889_ = new_n2857_ & ~new_n2888_;
  assign new_n2890_ = ~pi0093 & ~new_n2889_;
  assign new_n2891_ = new_n2856_ & ~new_n2890_;
  assign new_n2892_ = new_n2528_ & ~new_n2891_;
  assign new_n2893_ = new_n2874_ & ~new_n2892_;
  assign new_n2894_ = ~pi0072 & ~new_n2893_;
  assign new_n2895_ = new_n2556_ & ~new_n2894_;
  assign new_n2896_ = new_n2880_ & ~new_n2895_;
  assign new_n2897_ = ~new_n2845_ & ~new_n2896_;
  assign new_n2898_ = ~new_n2879_ & new_n2897_;
  assign new_n2899_ = ~pi0095 & ~new_n2898_;
  assign new_n2900_ = new_n2787_ & ~new_n2899_;
  assign new_n2901_ = ~pi0137 & ~new_n2900_;
  assign new_n2902_ = ~new_n2854_ & ~new_n2901_;
  assign new_n2903_ = ~pi0210 & ~new_n2902_;
  assign new_n2904_ = pi0146 & new_n2903_;
  assign new_n2905_ = ~pi0225 & new_n2499_;
  assign new_n2906_ = pi0032 & ~new_n2905_;
  assign new_n2907_ = ~new_n2878_ & ~new_n2906_;
  assign new_n2908_ = ~pi0095 & ~new_n2907_;
  assign new_n2909_ = ~pi0137 & new_n2787_;
  assign new_n2910_ = ~new_n2908_ & new_n2909_;
  assign new_n2911_ = ~pi0095 & ~new_n2906_;
  assign new_n2912_ = pi0137 & new_n2911_;
  assign new_n2913_ = ~new_n2852_ & new_n2912_;
  assign new_n2914_ = pi0210 & ~new_n2913_;
  assign new_n2915_ = ~new_n2910_ & new_n2914_;
  assign new_n2916_ = new_n2821_ & ~new_n2915_;
  assign new_n2917_ = ~pi0146 & ~pi0210;
  assign new_n2918_ = ~new_n2845_ & ~new_n2878_;
  assign new_n2919_ = ~pi0095 & ~new_n2918_;
  assign new_n2920_ = new_n2787_ & ~new_n2919_;
  assign new_n2921_ = ~pi0137 & ~new_n2920_;
  assign new_n2922_ = ~new_n2854_ & ~new_n2921_;
  assign new_n2923_ = new_n2917_ & ~new_n2922_;
  assign new_n2924_ = new_n2916_ & ~new_n2923_;
  assign new_n2925_ = ~new_n2904_ & new_n2924_;
  assign new_n2926_ = ~pi0072 & ~new_n2716_;
  assign new_n2927_ = ~new_n2875_ & new_n2926_;
  assign new_n2928_ = new_n2556_ & ~new_n2927_;
  assign new_n2929_ = new_n2554_ & ~new_n2928_;
  assign new_n2930_ = ~new_n2795_ & new_n2929_;
  assign new_n2931_ = ~new_n2893_ & new_n2926_;
  assign new_n2932_ = new_n2556_ & ~new_n2931_;
  assign new_n2933_ = new_n2880_ & ~new_n2932_;
  assign new_n2934_ = ~new_n2845_ & ~new_n2933_;
  assign new_n2935_ = ~new_n2930_ & new_n2934_;
  assign new_n2936_ = ~pi0095 & ~new_n2935_;
  assign new_n2937_ = ~new_n2726_ & ~new_n2936_;
  assign new_n2938_ = ~pi0137 & ~new_n2937_;
  assign new_n2939_ = ~pi0072 & new_n2724_;
  assign new_n2940_ = new_n2716_ & new_n2939_;
  assign new_n2941_ = new_n2852_ & ~new_n2940_;
  assign new_n2942_ = new_n2846_ & ~new_n2941_;
  assign new_n2943_ = new_n2449_ & new_n2725_;
  assign new_n2944_ = pi0137 & ~new_n2943_;
  assign new_n2945_ = ~new_n2942_ & new_n2944_;
  assign new_n2946_ = ~new_n2938_ & ~new_n2945_;
  assign new_n2947_ = ~pi0210 & ~new_n2946_;
  assign new_n2948_ = pi0146 & new_n2947_;
  assign new_n2949_ = ~pi0137 & ~new_n2726_;
  assign new_n2950_ = ~new_n2906_ & ~new_n2929_;
  assign new_n2951_ = ~pi0095 & ~new_n2950_;
  assign new_n2952_ = new_n2949_ & ~new_n2951_;
  assign new_n2953_ = new_n2911_ & ~new_n2941_;
  assign new_n2954_ = ~new_n2943_ & ~new_n2953_;
  assign new_n2955_ = pi0137 & ~new_n2954_;
  assign new_n2956_ = pi0210 & ~new_n2955_;
  assign new_n2957_ = ~new_n2952_ & new_n2956_;
  assign new_n2958_ = new_n2833_ & ~new_n2957_;
  assign new_n2959_ = ~new_n2845_ & ~new_n2929_;
  assign new_n2960_ = ~pi0095 & ~new_n2959_;
  assign new_n2961_ = ~new_n2726_ & ~new_n2960_;
  assign new_n2962_ = ~pi0137 & ~new_n2961_;
  assign new_n2963_ = ~new_n2945_ & ~new_n2962_;
  assign new_n2964_ = new_n2917_ & ~new_n2963_;
  assign new_n2965_ = new_n2958_ & ~new_n2964_;
  assign new_n2966_ = ~new_n2948_ & new_n2965_;
  assign new_n2967_ = ~new_n2448_ & ~new_n2966_;
  assign new_n2968_ = ~new_n2925_ & new_n2967_;
  assign new_n2969_ = ~new_n2947_ & new_n2958_;
  assign new_n2970_ = ~new_n2903_ & new_n2916_;
  assign new_n2971_ = new_n2448_ & ~new_n2970_;
  assign new_n2972_ = ~new_n2969_ & new_n2971_;
  assign new_n2973_ = ~pi0153 & ~new_n2972_;
  assign new_n2974_ = ~new_n2968_ & new_n2973_;
  assign new_n2975_ = ~pi0109 & ~new_n2695_;
  assign new_n2976_ = ~new_n2575_ & ~new_n2975_;
  assign new_n2977_ = new_n2574_ & ~new_n2976_;
  assign new_n2978_ = new_n2573_ & ~new_n2977_;
  assign new_n2979_ = new_n2566_ & ~new_n2978_;
  assign new_n2980_ = new_n2707_ & ~new_n2979_;
  assign new_n2981_ = new_n2564_ & ~new_n2980_;
  assign new_n2982_ = new_n2562_ & ~new_n2981_;
  assign new_n2983_ = ~pi0051 & ~new_n2982_;
  assign new_n2984_ = new_n2561_ & ~new_n2983_;
  assign new_n2985_ = ~pi0072 & ~new_n2984_;
  assign new_n2986_ = new_n2556_ & ~new_n2985_;
  assign new_n2987_ = new_n2554_ & ~new_n2986_;
  assign new_n2988_ = ~new_n2720_ & new_n2987_;
  assign new_n2989_ = ~new_n2741_ & ~new_n2988_;
  assign new_n2990_ = ~pi0095 & ~new_n2989_;
  assign new_n2991_ = ~new_n2726_ & ~new_n2990_;
  assign new_n2992_ = pi0137 & ~new_n2991_;
  assign new_n2993_ = ~pi0146 & ~new_n2448_;
  assign new_n2994_ = new_n2733_ & ~new_n2993_;
  assign new_n2995_ = ~new_n2756_ & new_n2994_;
  assign new_n2996_ = ~new_n2726_ & new_n2749_;
  assign new_n2997_ = ~new_n2995_ & new_n2996_;
  assign new_n2998_ = ~new_n2726_ & new_n2994_;
  assign new_n2999_ = new_n2773_ & new_n2998_;
  assign new_n3000_ = ~pi0137 & ~new_n2999_;
  assign new_n3001_ = ~new_n2997_ & new_n3000_;
  assign new_n3002_ = ~new_n2992_ & ~new_n3001_;
  assign new_n3003_ = ~pi0210 & ~new_n3002_;
  assign new_n3004_ = pi0234 & ~new_n3003_;
  assign new_n3005_ = ~new_n2741_ & ~new_n2987_;
  assign new_n3006_ = ~pi0095 & ~new_n3005_;
  assign new_n3007_ = new_n2787_ & ~new_n3006_;
  assign new_n3008_ = pi0137 & ~new_n3007_;
  assign new_n3009_ = new_n2808_ & ~new_n2993_;
  assign new_n3010_ = new_n2828_ & new_n2993_;
  assign new_n3011_ = ~pi0210 & ~pi0234;
  assign new_n3012_ = ~new_n3010_ & new_n3011_;
  assign new_n3013_ = ~new_n3009_ & new_n3012_;
  assign new_n3014_ = ~new_n3008_ & new_n3013_;
  assign new_n3015_ = ~new_n2501_ & ~new_n2987_;
  assign new_n3016_ = ~pi0095 & ~new_n3015_;
  assign new_n3017_ = new_n2787_ & ~new_n3016_;
  assign new_n3018_ = pi0137 & ~new_n3017_;
  assign new_n3019_ = pi0210 & ~new_n2786_;
  assign new_n3020_ = ~new_n3018_ & new_n3019_;
  assign new_n3021_ = ~new_n3014_ & ~new_n3020_;
  assign new_n3022_ = ~new_n3004_ & new_n3021_;
  assign new_n3023_ = ~new_n2501_ & ~new_n2988_;
  assign new_n3024_ = ~pi0095 & ~new_n3023_;
  assign new_n3025_ = pi0137 & ~new_n2726_;
  assign new_n3026_ = ~new_n3024_ & new_n3025_;
  assign new_n3027_ = ~new_n2545_ & new_n2949_;
  assign new_n3028_ = pi0210 & pi0234;
  assign new_n3029_ = ~new_n3027_ & new_n3028_;
  assign new_n3030_ = ~new_n3026_ & new_n3029_;
  assign new_n3031_ = ~new_n3022_ & ~new_n3030_;
  assign new_n3032_ = new_n2445_ & ~new_n3031_;
  assign new_n3033_ = ~pi0228 & ~new_n3032_;
  assign new_n3034_ = ~new_n2974_ & new_n3033_;
  assign new_n3035_ = ~new_n2842_ & ~new_n3034_;
  assign new_n3036_ = ~pi0216 & ~new_n3035_;
  assign new_n3037_ = ~new_n2444_ & ~new_n3036_;
  assign new_n3038_ = ~pi0221 & ~new_n3037_;
  assign new_n3039_ = ~new_n2442_ & ~new_n3038_;
  assign new_n3040_ = ~pi0215 & ~new_n3039_;
  assign new_n3041_ = ~pi0332 & ~pi1144;
  assign new_n3042_ = pi0215 & ~new_n3041_;
  assign new_n3043_ = pi0299 & ~new_n3042_;
  assign new_n3044_ = ~new_n3040_ & new_n3043_;
  assign new_n3045_ = ~pi0224 & pi0833;
  assign new_n3046_ = pi0222 & ~new_n3045_;
  assign new_n3047_ = ~pi0223 & ~new_n3046_;
  assign new_n3048_ = new_n3041_ & ~new_n3047_;
  assign new_n3049_ = pi0224 & ~new_n2443_;
  assign new_n3050_ = ~pi0222 & ~new_n3049_;
  assign new_n3051_ = ~pi0332 & ~pi0929;
  assign new_n3052_ = new_n3045_ & new_n3051_;
  assign new_n3053_ = ~new_n3050_ & ~new_n3052_;
  assign new_n3054_ = ~pi0223 & ~new_n3053_;
  assign new_n3055_ = ~new_n3048_ & ~new_n3054_;
  assign new_n3056_ = ~pi0299 & ~new_n3055_;
  assign new_n3057_ = ~pi0222 & ~pi0224;
  assign new_n3058_ = pi0198 & ~new_n2730_;
  assign new_n3059_ = ~pi0198 & new_n2778_;
  assign new_n3060_ = ~new_n3058_ & ~new_n3059_;
  assign new_n3061_ = pi0142 & new_n3060_;
  assign new_n3062_ = ~pi0198 & ~new_n2751_;
  assign new_n3063_ = ~pi0142 & ~new_n3058_;
  assign new_n3064_ = ~new_n3062_ & new_n3063_;
  assign new_n3065_ = new_n2821_ & ~new_n3064_;
  assign new_n3066_ = ~new_n3061_ & new_n3065_;
  assign new_n3067_ = ~pi0144 & ~pi0174;
  assign new_n3068_ = ~pi0189 & new_n3067_;
  assign new_n3069_ = ~pi0223 & ~new_n3068_;
  assign new_n3070_ = ~pi0198 & ~new_n2829_;
  assign new_n3071_ = pi0198 & ~new_n2792_;
  assign new_n3072_ = ~pi0142 & ~new_n3071_;
  assign new_n3073_ = ~new_n3070_ & new_n3072_;
  assign new_n3074_ = ~pi0198 & ~new_n2813_;
  assign new_n3075_ = ~new_n3071_ & ~new_n3074_;
  assign new_n3076_ = pi0142 & new_n3075_;
  assign new_n3077_ = new_n2833_ & ~new_n3076_;
  assign new_n3078_ = ~new_n3073_ & new_n3077_;
  assign new_n3079_ = new_n3069_ & ~new_n3078_;
  assign new_n3080_ = ~new_n3066_ & new_n3079_;
  assign new_n3081_ = ~pi0223 & new_n3068_;
  assign new_n3082_ = pi0234 & new_n3060_;
  assign new_n3083_ = ~pi0234 & new_n3075_;
  assign new_n3084_ = ~pi0332 & ~new_n3083_;
  assign new_n3085_ = ~new_n3082_ & new_n3084_;
  assign new_n3086_ = new_n3081_ & ~new_n3085_;
  assign new_n3087_ = ~new_n3080_ & ~new_n3086_;
  assign new_n3088_ = new_n3057_ & ~new_n3087_;
  assign new_n3089_ = new_n3056_ & ~new_n3088_;
  assign new_n3090_ = ~pi0039 & ~new_n3089_;
  assign new_n3091_ = ~new_n3044_ & new_n3090_;
  assign new_n3092_ = pi0234 & new_n2449_;
  assign new_n3093_ = ~pi0332 & ~new_n3092_;
  assign new_n3094_ = ~pi0095 & new_n2725_;
  assign new_n3095_ = ~new_n2449_ & ~new_n3094_;
  assign new_n3096_ = pi0234 & ~new_n3095_;
  assign new_n3097_ = ~pi0032 & ~pi0095;
  assign new_n3098_ = new_n2450_ & new_n3097_;
  assign new_n3099_ = new_n2847_ & new_n3098_;
  assign new_n3100_ = new_n2557_ & new_n3099_;
  assign new_n3101_ = ~pi0234 & new_n3100_;
  assign new_n3102_ = ~new_n3096_ & ~new_n3101_;
  assign new_n3103_ = pi0137 & ~new_n3102_;
  assign new_n3104_ = new_n3093_ & ~new_n3103_;
  assign new_n3105_ = ~pi0223 & new_n3057_;
  assign new_n3106_ = ~new_n3104_ & new_n3105_;
  assign new_n3107_ = ~new_n3055_ & ~new_n3106_;
  assign new_n3108_ = ~pi0299 & ~new_n3107_;
  assign new_n3109_ = pi0105 & ~new_n3104_;
  assign new_n3110_ = ~new_n2446_ & ~new_n3109_;
  assign new_n3111_ = pi0228 & ~new_n3110_;
  assign new_n3112_ = ~pi0332 & new_n3094_;
  assign new_n3113_ = ~pi0137 & ~pi0153;
  assign new_n3114_ = new_n3112_ & new_n3113_;
  assign new_n3115_ = pi0137 & new_n3100_;
  assign new_n3116_ = new_n2445_ & ~new_n3115_;
  assign new_n3117_ = ~pi0228 & ~new_n3116_;
  assign new_n3118_ = ~new_n3114_ & new_n3117_;
  assign new_n3119_ = ~new_n3111_ & ~new_n3118_;
  assign new_n3120_ = ~pi0216 & ~new_n3119_;
  assign new_n3121_ = ~new_n2444_ & ~new_n3120_;
  assign new_n3122_ = ~pi0221 & ~new_n3121_;
  assign new_n3123_ = ~new_n2442_ & ~new_n3122_;
  assign new_n3124_ = ~pi0215 & ~new_n3123_;
  assign new_n3125_ = ~new_n3042_ & ~new_n3124_;
  assign new_n3126_ = pi0299 & ~new_n3125_;
  assign new_n3127_ = ~new_n3108_ & ~new_n3126_;
  assign new_n3128_ = pi0039 & ~new_n3127_;
  assign new_n3129_ = ~pi0038 & ~new_n3128_;
  assign new_n3130_ = ~new_n3091_ & new_n3129_;
  assign new_n3131_ = pi0105 & pi0228;
  assign new_n3132_ = new_n3093_ & new_n3131_;
  assign new_n3133_ = new_n2445_ & ~new_n3131_;
  assign new_n3134_ = ~pi0216 & ~new_n3133_;
  assign new_n3135_ = ~new_n3132_ & new_n3134_;
  assign new_n3136_ = ~new_n2444_ & ~new_n3135_;
  assign new_n3137_ = ~pi0221 & ~new_n3136_;
  assign new_n3138_ = ~new_n2442_ & ~new_n3137_;
  assign new_n3139_ = ~pi0215 & ~new_n3138_;
  assign new_n3140_ = ~new_n3042_ & ~new_n3139_;
  assign new_n3141_ = ~pi0215 & ~pi0221;
  assign new_n3142_ = new_n3134_ & new_n3141_;
  assign new_n3143_ = ~new_n3104_ & new_n3142_;
  assign new_n3144_ = new_n3140_ & ~new_n3143_;
  assign new_n3145_ = pi0299 & ~new_n3144_;
  assign new_n3146_ = ~new_n3108_ & ~new_n3145_;
  assign new_n3147_ = ~pi0039 & ~new_n3146_;
  assign new_n3148_ = pi0299 & new_n3140_;
  assign new_n3149_ = ~new_n3093_ & new_n3105_;
  assign new_n3150_ = new_n3056_ & ~new_n3149_;
  assign new_n3151_ = ~new_n3148_ & ~new_n3150_;
  assign new_n3152_ = pi0039 & new_n3151_;
  assign new_n3153_ = pi0038 & ~new_n3152_;
  assign new_n3154_ = ~new_n3147_ & new_n3153_;
  assign new_n3155_ = ~pi0100 & ~new_n3154_;
  assign new_n3156_ = ~new_n3130_ & new_n3155_;
  assign new_n3157_ = pi0228 & ~new_n2446_;
  assign new_n3158_ = ~pi0210 & ~new_n2993_;
  assign new_n3159_ = pi0095 & pi0234;
  assign new_n3160_ = ~pi0137 & ~new_n3159_;
  assign new_n3161_ = ~new_n3158_ & new_n3160_;
  assign new_n3162_ = ~new_n3102_ & ~new_n3161_;
  assign new_n3163_ = ~pi0332 & ~new_n3162_;
  assign new_n3164_ = pi0105 & ~new_n3163_;
  assign new_n3165_ = new_n3157_ & ~new_n3164_;
  assign new_n3166_ = ~pi0137 & pi0210;
  assign new_n3167_ = ~pi0252 & ~new_n3166_;
  assign new_n3168_ = ~new_n2993_ & new_n3167_;
  assign new_n3169_ = new_n3112_ & new_n3168_;
  assign new_n3170_ = new_n2993_ & new_n3115_;
  assign new_n3171_ = new_n2445_ & ~new_n3170_;
  assign new_n3172_ = ~new_n3169_ & new_n3171_;
  assign new_n3173_ = pi0252 & ~new_n2993_;
  assign new_n3174_ = ~new_n3158_ & ~new_n3173_;
  assign new_n3175_ = new_n3114_ & new_n3174_;
  assign new_n3176_ = ~new_n3172_ & ~new_n3175_;
  assign new_n3177_ = ~pi0228 & ~new_n3176_;
  assign new_n3178_ = ~pi0216 & ~new_n3177_;
  assign new_n3179_ = ~new_n3165_ & new_n3178_;
  assign new_n3180_ = ~new_n2444_ & ~new_n3179_;
  assign new_n3181_ = ~pi0221 & ~new_n3180_;
  assign new_n3182_ = ~new_n2442_ & ~new_n3181_;
  assign new_n3183_ = ~pi0215 & ~new_n3182_;
  assign new_n3184_ = ~new_n3042_ & ~new_n3183_;
  assign new_n3185_ = pi0299 & ~new_n3184_;
  assign new_n3186_ = ~pi0038 & ~pi0039;
  assign new_n3187_ = pi0142 & ~pi0198;
  assign new_n3188_ = ~pi0137 & ~new_n3187_;
  assign new_n3189_ = ~new_n3102_ & ~new_n3188_;
  assign new_n3190_ = new_n3093_ & ~new_n3189_;
  assign new_n3191_ = new_n3069_ & ~new_n3190_;
  assign new_n3192_ = ~pi0137 & pi0198;
  assign new_n3193_ = ~pi0095 & new_n3192_;
  assign new_n3194_ = ~new_n3095_ & ~new_n3193_;
  assign new_n3195_ = new_n2821_ & ~new_n3194_;
  assign new_n3196_ = new_n3100_ & ~new_n3192_;
  assign new_n3197_ = new_n2833_ & ~new_n3196_;
  assign new_n3198_ = new_n3081_ & ~new_n3197_;
  assign new_n3199_ = ~new_n3195_ & new_n3198_;
  assign new_n3200_ = ~new_n3191_ & ~new_n3199_;
  assign new_n3201_ = new_n3057_ & ~new_n3200_;
  assign new_n3202_ = ~new_n3055_ & ~new_n3201_;
  assign new_n3203_ = ~pi0299 & ~new_n3202_;
  assign new_n3204_ = new_n3186_ & ~new_n3203_;
  assign new_n3205_ = ~new_n3185_ & new_n3204_;
  assign new_n3206_ = ~new_n3151_ & ~new_n3186_;
  assign new_n3207_ = pi0100 & ~new_n3206_;
  assign new_n3208_ = ~new_n3205_ & new_n3207_;
  assign new_n3209_ = ~pi0087 & ~new_n3208_;
  assign new_n3210_ = ~new_n3156_ & new_n3209_;
  assign new_n3211_ = ~pi0038 & ~pi0100;
  assign new_n3212_ = ~pi0039 & new_n3211_;
  assign new_n3213_ = ~new_n3151_ & ~new_n3212_;
  assign new_n3214_ = new_n3127_ & new_n3212_;
  assign new_n3215_ = ~new_n3213_ & ~new_n3214_;
  assign new_n3216_ = pi0087 & ~new_n3215_;
  assign new_n3217_ = ~pi0075 & ~new_n3216_;
  assign new_n3218_ = ~new_n3210_ & new_n3217_;
  assign new_n3219_ = new_n3134_ & ~new_n3165_;
  assign new_n3220_ = ~new_n2444_ & ~new_n3219_;
  assign new_n3221_ = ~pi0221 & ~new_n3220_;
  assign new_n3222_ = ~new_n2442_ & ~new_n3221_;
  assign new_n3223_ = ~pi0215 & ~new_n3222_;
  assign new_n3224_ = ~new_n3042_ & ~new_n3223_;
  assign new_n3225_ = pi0299 & ~new_n3224_;
  assign new_n3226_ = ~pi0039 & ~pi0087;
  assign new_n3227_ = new_n3211_ & new_n3226_;
  assign new_n3228_ = ~new_n3203_ & new_n3227_;
  assign new_n3229_ = ~new_n3225_ & new_n3228_;
  assign new_n3230_ = ~new_n3151_ & ~new_n3227_;
  assign new_n3231_ = pi0075 & ~new_n3230_;
  assign new_n3232_ = ~new_n3229_ & new_n3231_;
  assign new_n3233_ = ~new_n3218_ & ~new_n3232_;
  assign new_n3234_ = ~pi0092 & ~new_n3233_;
  assign new_n3235_ = ~pi0075 & ~pi0087;
  assign new_n3236_ = ~new_n3215_ & new_n3235_;
  assign new_n3237_ = ~new_n3151_ & ~new_n3235_;
  assign new_n3238_ = pi0092 & ~new_n3237_;
  assign new_n3239_ = ~new_n3236_ & new_n3238_;
  assign new_n3240_ = ~pi0054 & ~new_n3239_;
  assign new_n3241_ = ~new_n3234_ & new_n3240_;
  assign new_n3242_ = ~pi0075 & ~pi0092;
  assign new_n3243_ = new_n3227_ & new_n3242_;
  assign new_n3244_ = new_n3151_ & ~new_n3243_;
  assign new_n3245_ = ~pi0087 & ~pi0100;
  assign new_n3246_ = ~pi0038 & new_n3245_;
  assign new_n3247_ = new_n3242_ & new_n3246_;
  assign new_n3248_ = new_n3147_ & new_n3247_;
  assign new_n3249_ = ~new_n3244_ & ~new_n3248_;
  assign new_n3250_ = pi0054 & new_n3249_;
  assign new_n3251_ = ~pi0074 & ~new_n3250_;
  assign new_n3252_ = ~new_n3241_ & new_n3251_;
  assign new_n3253_ = ~pi0054 & new_n3249_;
  assign new_n3254_ = pi0054 & ~new_n3151_;
  assign new_n3255_ = pi0074 & ~new_n3254_;
  assign new_n3256_ = ~new_n3253_ & new_n3255_;
  assign new_n3257_ = ~new_n3252_ & ~new_n3256_;
  assign new_n3258_ = ~pi0055 & ~new_n3257_;
  assign new_n3259_ = ~pi0332 & new_n3102_;
  assign new_n3260_ = pi0105 & ~new_n3259_;
  assign new_n3261_ = new_n3157_ & ~new_n3260_;
  assign new_n3262_ = ~pi0228 & new_n2445_;
  assign new_n3263_ = ~new_n3100_ & new_n3262_;
  assign new_n3264_ = ~pi0216 & ~new_n3263_;
  assign new_n3265_ = ~new_n3261_ & new_n3264_;
  assign new_n3266_ = ~new_n2444_ & ~new_n3265_;
  assign new_n3267_ = ~pi0221 & ~new_n3266_;
  assign new_n3268_ = ~new_n2442_ & ~new_n3267_;
  assign new_n3269_ = ~pi0215 & ~new_n3268_;
  assign new_n3270_ = ~pi0054 & ~pi0074;
  assign new_n3271_ = new_n3242_ & new_n3270_;
  assign new_n3272_ = new_n3245_ & new_n3271_;
  assign new_n3273_ = new_n3186_ & new_n3272_;
  assign new_n3274_ = ~new_n3042_ & new_n3273_;
  assign new_n3275_ = ~new_n3269_ & new_n3274_;
  assign new_n3276_ = new_n3140_ & ~new_n3273_;
  assign new_n3277_ = pi0055 & ~new_n3276_;
  assign new_n3278_ = ~new_n3275_ & new_n3277_;
  assign new_n3279_ = ~pi0056 & ~new_n3278_;
  assign new_n3280_ = ~new_n3258_ & new_n3279_;
  assign new_n3281_ = ~pi0100 & new_n3186_;
  assign new_n3282_ = ~pi0092 & new_n3235_;
  assign new_n3283_ = new_n3270_ & new_n3282_;
  assign new_n3284_ = ~pi0055 & new_n3283_;
  assign new_n3285_ = new_n3281_ & new_n3284_;
  assign new_n3286_ = new_n3140_ & ~new_n3285_;
  assign new_n3287_ = new_n3125_ & new_n3285_;
  assign new_n3288_ = ~new_n3286_ & ~new_n3287_;
  assign new_n3289_ = pi0056 & ~new_n3288_;
  assign new_n3290_ = ~pi0062 & ~new_n3289_;
  assign new_n3291_ = ~new_n3280_ & new_n3290_;
  assign new_n3292_ = ~pi0056 & ~new_n3288_;
  assign new_n3293_ = pi0056 & new_n3140_;
  assign new_n3294_ = pi0062 & ~new_n3293_;
  assign new_n3295_ = ~new_n3292_ & new_n3294_;
  assign new_n3296_ = ~pi0059 & ~new_n3295_;
  assign new_n3297_ = ~new_n3291_ & new_n3296_;
  assign new_n3298_ = ~pi0056 & ~pi0062;
  assign new_n3299_ = new_n3285_ & new_n3298_;
  assign new_n3300_ = new_n3143_ & new_n3299_;
  assign new_n3301_ = pi0059 & new_n3140_;
  assign new_n3302_ = ~new_n3300_ & new_n3301_;
  assign new_n3303_ = ~pi0057 & ~new_n3302_;
  assign new_n3304_ = ~new_n3297_ & new_n3303_;
  assign new_n3305_ = ~pi0059 & new_n3300_;
  assign new_n3306_ = new_n3140_ & ~new_n3305_;
  assign new_n3307_ = pi0057 & ~new_n3306_;
  assign po0153 = new_n3304_ | new_n3307_;
  assign new_n3309_ = ~pi0939 & new_n3045_;
  assign new_n3310_ = ~pi1146 & ~new_n3045_;
  assign new_n3311_ = pi0222 & ~new_n3310_;
  assign new_n3312_ = ~new_n3309_ & new_n3311_;
  assign new_n3313_ = ~pi0222 & pi0224;
  assign new_n3314_ = pi0276 & new_n3313_;
  assign new_n3315_ = ~pi0223 & ~new_n3314_;
  assign new_n3316_ = ~new_n3312_ & new_n3315_;
  assign new_n3317_ = pi0223 & ~pi1146;
  assign new_n3318_ = ~pi0299 & ~new_n3317_;
  assign new_n3319_ = ~new_n3316_ & new_n3318_;
  assign new_n3320_ = pi0215 & pi1146;
  assign new_n3321_ = ~pi0939 & new_n2437_;
  assign new_n3322_ = ~pi1146 & ~new_n2437_;
  assign new_n3323_ = pi0221 & ~new_n3322_;
  assign new_n3324_ = ~new_n3321_ & new_n3323_;
  assign new_n3325_ = ~new_n3320_ & ~new_n3324_;
  assign new_n3326_ = ~pi0228 & new_n3100_;
  assign new_n3327_ = ~pi0216 & new_n3326_;
  assign new_n3328_ = new_n3325_ & new_n3327_;
  assign new_n3329_ = pi0216 & ~pi0221;
  assign new_n3330_ = pi0276 & new_n3329_;
  assign new_n3331_ = ~pi0216 & ~new_n3131_;
  assign new_n3332_ = ~new_n3330_ & ~new_n3331_;
  assign new_n3333_ = ~pi0221 & ~new_n3332_;
  assign new_n3334_ = ~new_n3324_ & ~new_n3333_;
  assign new_n3335_ = ~pi0215 & ~new_n3334_;
  assign new_n3336_ = ~new_n3320_ & ~new_n3335_;
  assign new_n3337_ = pi0299 & ~new_n3336_;
  assign new_n3338_ = ~new_n3328_ & new_n3337_;
  assign new_n3339_ = ~new_n3319_ & ~new_n3338_;
  assign new_n3340_ = ~pi0154 & ~new_n3339_;
  assign new_n3341_ = ~new_n3324_ & ~new_n3330_;
  assign new_n3342_ = ~pi0215 & ~new_n3341_;
  assign new_n3343_ = ~new_n3320_ & ~new_n3342_;
  assign new_n3344_ = pi0299 & ~new_n3343_;
  assign new_n3345_ = ~new_n3319_ & ~new_n3344_;
  assign new_n3346_ = pi0154 & ~new_n3345_;
  assign new_n3347_ = new_n3212_ & ~new_n3346_;
  assign new_n3348_ = ~new_n3340_ & new_n3347_;
  assign new_n3349_ = pi0154 & ~new_n3343_;
  assign new_n3350_ = ~pi0154 & ~new_n3336_;
  assign new_n3351_ = ~new_n3349_ & ~new_n3350_;
  assign new_n3352_ = pi0299 & ~new_n3351_;
  assign new_n3353_ = ~new_n3319_ & ~new_n3352_;
  assign new_n3354_ = ~new_n3212_ & new_n3353_;
  assign new_n3355_ = ~new_n3348_ & ~new_n3354_;
  assign new_n3356_ = pi0087 & ~new_n3355_;
  assign new_n3357_ = pi0039 & ~new_n3100_;
  assign new_n3358_ = ~pi0070 & new_n2981_;
  assign new_n3359_ = ~new_n2524_ & ~new_n2848_;
  assign new_n3360_ = ~new_n3358_ & new_n3359_;
  assign new_n3361_ = ~pi0051 & ~new_n3360_;
  assign new_n3362_ = new_n2559_ & ~new_n3361_;
  assign new_n3363_ = new_n2926_ & ~new_n3362_;
  assign new_n3364_ = ~new_n2555_ & ~new_n3363_;
  assign new_n3365_ = new_n2724_ & ~new_n3364_;
  assign new_n3366_ = pi0040 & ~new_n2552_;
  assign new_n3367_ = pi0032 & ~new_n2499_;
  assign new_n3368_ = ~new_n3366_ & ~new_n3367_;
  assign new_n3369_ = ~new_n3365_ & new_n3368_;
  assign new_n3370_ = ~pi0095 & ~new_n3369_;
  assign new_n3371_ = ~new_n2726_ & ~new_n3370_;
  assign new_n3372_ = ~pi0039 & ~new_n3371_;
  assign new_n3373_ = ~new_n3357_ & ~new_n3372_;
  assign new_n3374_ = ~pi0216 & ~pi0228;
  assign new_n3375_ = new_n3325_ & new_n3374_;
  assign new_n3376_ = new_n3373_ & new_n3375_;
  assign new_n3377_ = new_n3337_ & ~new_n3376_;
  assign new_n3378_ = ~new_n3319_ & ~new_n3377_;
  assign new_n3379_ = ~pi0154 & ~new_n3378_;
  assign new_n3380_ = ~pi0038 & ~new_n3346_;
  assign new_n3381_ = ~new_n3379_ & new_n3380_;
  assign new_n3382_ = pi0038 & new_n3353_;
  assign new_n3383_ = ~pi0100 & ~new_n3382_;
  assign new_n3384_ = ~new_n3381_ & new_n3383_;
  assign new_n3385_ = ~pi0146 & ~new_n3100_;
  assign new_n3386_ = ~pi0252 & new_n3100_;
  assign new_n3387_ = pi0146 & ~new_n3386_;
  assign new_n3388_ = ~new_n3385_ & ~new_n3387_;
  assign new_n3389_ = pi0152 & ~new_n3388_;
  assign new_n3390_ = ~pi0161 & ~pi0166;
  assign new_n3391_ = new_n3388_ & ~new_n3390_;
  assign new_n3392_ = new_n3386_ & new_n3390_;
  assign new_n3393_ = ~pi0152 & ~new_n3392_;
  assign new_n3394_ = ~new_n3391_ & new_n3393_;
  assign new_n3395_ = ~new_n3389_ & ~new_n3394_;
  assign new_n3396_ = ~pi0038 & ~pi0216;
  assign new_n3397_ = ~pi0228 & new_n3396_;
  assign new_n3398_ = ~pi0154 & pi0299;
  assign new_n3399_ = ~pi0039 & new_n3398_;
  assign new_n3400_ = new_n3397_ & new_n3399_;
  assign new_n3401_ = new_n3325_ & new_n3400_;
  assign new_n3402_ = new_n3395_ & new_n3401_;
  assign new_n3403_ = pi0100 & ~new_n3353_;
  assign new_n3404_ = ~new_n3402_ & new_n3403_;
  assign new_n3405_ = ~pi0087 & ~new_n3404_;
  assign new_n3406_ = ~new_n3384_ & new_n3405_;
  assign new_n3407_ = ~new_n3356_ & ~new_n3406_;
  assign new_n3408_ = ~pi0075 & ~new_n3407_;
  assign new_n3409_ = pi0075 & new_n3353_;
  assign new_n3410_ = ~pi0092 & ~new_n3409_;
  assign new_n3411_ = ~new_n3408_ & new_n3410_;
  assign new_n3412_ = new_n3235_ & new_n3348_;
  assign new_n3413_ = new_n3235_ & new_n3281_;
  assign new_n3414_ = new_n3353_ & ~new_n3413_;
  assign new_n3415_ = pi0092 & ~new_n3414_;
  assign new_n3416_ = ~new_n3412_ & new_n3415_;
  assign new_n3417_ = new_n3270_ & ~new_n3416_;
  assign new_n3418_ = ~new_n3411_ & new_n3417_;
  assign new_n3419_ = ~new_n3270_ & new_n3353_;
  assign new_n3420_ = ~pi0055 & ~new_n3419_;
  assign new_n3421_ = ~new_n3418_ & new_n3420_;
  assign new_n3422_ = new_n3328_ & ~new_n3349_;
  assign new_n3423_ = new_n3273_ & new_n3422_;
  assign new_n3424_ = pi0055 & ~new_n3351_;
  assign new_n3425_ = ~new_n3423_ & new_n3424_;
  assign new_n3426_ = ~pi0056 & ~new_n3425_;
  assign new_n3427_ = ~new_n3421_ & new_n3426_;
  assign new_n3428_ = ~pi0055 & new_n3273_;
  assign new_n3429_ = ~new_n3351_ & new_n3428_;
  assign new_n3430_ = ~new_n3422_ & new_n3429_;
  assign new_n3431_ = ~new_n3285_ & ~new_n3351_;
  assign new_n3432_ = pi0056 & ~new_n3431_;
  assign new_n3433_ = ~new_n3430_ & new_n3432_;
  assign new_n3434_ = ~pi0062 & ~new_n3433_;
  assign new_n3435_ = ~new_n3427_ & new_n3434_;
  assign new_n3436_ = ~pi0057 & ~pi0059;
  assign new_n3437_ = ~pi0056 & new_n3284_;
  assign new_n3438_ = new_n3281_ & new_n3437_;
  assign new_n3439_ = ~new_n3351_ & ~new_n3438_;
  assign new_n3440_ = ~new_n3430_ & ~new_n3439_;
  assign new_n3441_ = pi0062 & ~new_n3440_;
  assign new_n3442_ = new_n3436_ & ~new_n3441_;
  assign new_n3443_ = ~new_n3435_ & new_n3442_;
  assign new_n3444_ = new_n3351_ & ~new_n3436_;
  assign new_n3445_ = ~pi0239 & ~new_n3444_;
  assign new_n3446_ = ~new_n3443_ & new_n3445_;
  assign new_n3447_ = new_n2716_ & new_n3098_;
  assign new_n3448_ = ~new_n2449_ & ~new_n3447_;
  assign new_n3449_ = ~pi0224 & new_n3448_;
  assign new_n3450_ = pi0224 & ~pi0276;
  assign new_n3451_ = ~pi0222 & ~new_n3450_;
  assign new_n3452_ = ~new_n3449_ & new_n3451_;
  assign new_n3453_ = ~pi0223 & ~new_n3312_;
  assign new_n3454_ = ~new_n3452_ & new_n3453_;
  assign new_n3455_ = ~new_n3317_ & ~new_n3454_;
  assign new_n3456_ = ~pi0299 & ~new_n3455_;
  assign new_n3457_ = ~pi0072 & ~new_n3362_;
  assign new_n3458_ = ~new_n2555_ & ~new_n3457_;
  assign new_n3459_ = new_n2724_ & ~new_n3458_;
  assign new_n3460_ = new_n3368_ & ~new_n3459_;
  assign new_n3461_ = ~pi0095 & ~new_n3460_;
  assign new_n3462_ = new_n2787_ & ~new_n3461_;
  assign new_n3463_ = ~pi0228 & new_n3462_;
  assign new_n3464_ = new_n3131_ & new_n3448_;
  assign new_n3465_ = ~new_n3463_ & ~new_n3464_;
  assign new_n3466_ = ~pi0154 & ~new_n3465_;
  assign new_n3467_ = ~pi0216 & ~pi0221;
  assign new_n3468_ = ~pi0215 & new_n3467_;
  assign new_n3469_ = pi0105 & ~new_n3448_;
  assign new_n3470_ = pi0228 & ~new_n3469_;
  assign new_n3471_ = ~new_n2726_ & ~new_n3448_;
  assign new_n3472_ = ~pi0228 & ~new_n3471_;
  assign new_n3473_ = ~new_n3470_ & ~new_n3472_;
  assign new_n3474_ = pi0154 & ~new_n3473_;
  assign new_n3475_ = new_n3468_ & ~new_n3474_;
  assign new_n3476_ = ~new_n3466_ & new_n3475_;
  assign new_n3477_ = pi0299 & new_n3343_;
  assign new_n3478_ = ~new_n3476_ & new_n3477_;
  assign new_n3479_ = ~new_n3456_ & ~new_n3478_;
  assign new_n3480_ = ~pi0039 & ~new_n3479_;
  assign new_n3481_ = new_n2449_ & new_n3131_;
  assign new_n3482_ = new_n3468_ & new_n3481_;
  assign new_n3483_ = new_n3343_ & ~new_n3482_;
  assign new_n3484_ = pi0154 & ~new_n3483_;
  assign new_n3485_ = ~pi0215 & ~new_n3483_;
  assign new_n3486_ = ~new_n3350_ & ~new_n3485_;
  assign new_n3487_ = ~new_n3484_ & new_n3486_;
  assign new_n3488_ = pi0299 & ~new_n3487_;
  assign new_n3489_ = ~pi0223 & ~pi0299;
  assign new_n3490_ = new_n3057_ & new_n3489_;
  assign new_n3491_ = new_n2449_ & new_n3490_;
  assign new_n3492_ = ~new_n3319_ & ~new_n3491_;
  assign new_n3493_ = ~new_n3488_ & new_n3492_;
  assign new_n3494_ = new_n3328_ & ~new_n3484_;
  assign new_n3495_ = ~new_n3487_ & ~new_n3494_;
  assign new_n3496_ = pi0299 & ~new_n3495_;
  assign new_n3497_ = ~new_n3493_ & ~new_n3496_;
  assign new_n3498_ = pi0039 & ~new_n3497_;
  assign new_n3499_ = new_n3211_ & ~new_n3498_;
  assign new_n3500_ = ~new_n3480_ & new_n3499_;
  assign new_n3501_ = pi0100 & new_n3402_;
  assign new_n3502_ = ~new_n3211_ & ~new_n3493_;
  assign new_n3503_ = ~new_n3501_ & new_n3502_;
  assign new_n3504_ = ~new_n3500_ & ~new_n3503_;
  assign new_n3505_ = ~pi0087 & ~new_n3504_;
  assign new_n3506_ = new_n3212_ & new_n3496_;
  assign new_n3507_ = pi0087 & ~new_n3493_;
  assign new_n3508_ = ~new_n3506_ & new_n3507_;
  assign new_n3509_ = ~pi0075 & ~new_n3508_;
  assign new_n3510_ = ~new_n3505_ & new_n3509_;
  assign new_n3511_ = pi0075 & new_n3493_;
  assign new_n3512_ = ~pi0092 & ~new_n3511_;
  assign new_n3513_ = ~new_n3510_ & new_n3512_;
  assign new_n3514_ = new_n3413_ & new_n3496_;
  assign new_n3515_ = pi0092 & ~new_n3493_;
  assign new_n3516_ = ~new_n3514_ & new_n3515_;
  assign new_n3517_ = new_n3270_ & ~new_n3516_;
  assign new_n3518_ = ~new_n3513_ & new_n3517_;
  assign new_n3519_ = ~new_n3270_ & new_n3493_;
  assign new_n3520_ = ~pi0055 & ~new_n3519_;
  assign new_n3521_ = ~new_n3518_ & new_n3520_;
  assign new_n3522_ = new_n3273_ & new_n3494_;
  assign new_n3523_ = pi0055 & ~new_n3487_;
  assign new_n3524_ = ~new_n3522_ & new_n3523_;
  assign new_n3525_ = ~pi0056 & ~new_n3524_;
  assign new_n3526_ = ~new_n3521_ & new_n3525_;
  assign new_n3527_ = new_n3428_ & new_n3495_;
  assign new_n3528_ = ~new_n3285_ & ~new_n3487_;
  assign new_n3529_ = pi0056 & ~new_n3528_;
  assign new_n3530_ = ~new_n3527_ & new_n3529_;
  assign new_n3531_ = ~pi0062 & ~new_n3530_;
  assign new_n3532_ = ~new_n3526_ & new_n3531_;
  assign new_n3533_ = ~new_n3438_ & ~new_n3487_;
  assign new_n3534_ = ~pi0056 & new_n3527_;
  assign new_n3535_ = ~new_n3533_ & ~new_n3534_;
  assign new_n3536_ = pi0062 & ~new_n3535_;
  assign new_n3537_ = new_n3436_ & ~new_n3536_;
  assign new_n3538_ = ~new_n3532_ & new_n3537_;
  assign new_n3539_ = ~new_n3436_ & new_n3487_;
  assign new_n3540_ = pi0239 & ~new_n3539_;
  assign new_n3541_ = ~new_n3538_ & new_n3540_;
  assign po0154 = new_n3446_ | new_n3541_;
  assign new_n3543_ = ~pi0927 & new_n2437_;
  assign new_n3544_ = ~pi1145 & ~new_n2437_;
  assign new_n3545_ = pi0221 & ~new_n3544_;
  assign new_n3546_ = ~new_n3543_ & new_n3545_;
  assign new_n3547_ = pi0216 & pi0274;
  assign new_n3548_ = ~pi0221 & ~new_n3547_;
  assign new_n3549_ = ~pi0151 & new_n3465_;
  assign new_n3550_ = pi0151 & new_n3473_;
  assign new_n3551_ = ~pi0216 & ~new_n3550_;
  assign new_n3552_ = ~new_n3549_ & new_n3551_;
  assign new_n3553_ = new_n3548_ & ~new_n3552_;
  assign new_n3554_ = ~new_n3546_ & ~new_n3553_;
  assign new_n3555_ = ~pi0215 & ~new_n3554_;
  assign new_n3556_ = pi0215 & pi1145;
  assign new_n3557_ = pi0299 & ~new_n3556_;
  assign new_n3558_ = ~new_n3555_ & new_n3557_;
  assign new_n3559_ = ~pi0927 & new_n3045_;
  assign new_n3560_ = ~pi1145 & ~new_n3045_;
  assign new_n3561_ = pi0222 & ~new_n3560_;
  assign new_n3562_ = ~new_n3559_ & new_n3561_;
  assign new_n3563_ = pi0224 & pi0274;
  assign new_n3564_ = ~pi0222 & ~new_n3563_;
  assign new_n3565_ = ~new_n3449_ & new_n3564_;
  assign new_n3566_ = ~new_n3562_ & ~new_n3565_;
  assign new_n3567_ = ~pi0223 & ~new_n3566_;
  assign new_n3568_ = pi0223 & pi1145;
  assign new_n3569_ = ~pi0299 & ~new_n3568_;
  assign new_n3570_ = ~new_n3567_ & new_n3569_;
  assign new_n3571_ = ~pi0039 & ~new_n3570_;
  assign new_n3572_ = ~new_n3558_ & new_n3571_;
  assign new_n3573_ = new_n3313_ & ~new_n3563_;
  assign new_n3574_ = ~new_n3562_ & ~new_n3573_;
  assign new_n3575_ = ~pi0223 & ~new_n3574_;
  assign new_n3576_ = ~new_n3568_ & ~new_n3575_;
  assign new_n3577_ = ~pi0299 & ~new_n3576_;
  assign new_n3578_ = ~new_n3491_ & ~new_n3577_;
  assign new_n3579_ = ~pi0151 & ~new_n3131_;
  assign new_n3580_ = ~new_n3481_ & ~new_n3579_;
  assign new_n3581_ = ~pi0151 & new_n3326_;
  assign new_n3582_ = ~new_n3580_ & ~new_n3581_;
  assign new_n3583_ = ~pi0216 & ~new_n3582_;
  assign new_n3584_ = new_n3548_ & ~new_n3583_;
  assign new_n3585_ = ~new_n3546_ & ~new_n3584_;
  assign new_n3586_ = ~pi0215 & ~new_n3585_;
  assign new_n3587_ = ~new_n3556_ & ~new_n3586_;
  assign new_n3588_ = pi0299 & ~new_n3587_;
  assign new_n3589_ = new_n3578_ & ~new_n3588_;
  assign new_n3590_ = pi0039 & ~new_n3589_;
  assign new_n3591_ = ~pi0038 & ~new_n3590_;
  assign new_n3592_ = ~new_n3572_ & new_n3591_;
  assign new_n3593_ = ~pi0216 & ~new_n3579_;
  assign new_n3594_ = new_n3548_ & ~new_n3593_;
  assign new_n3595_ = ~new_n3546_ & ~new_n3594_;
  assign new_n3596_ = ~pi0215 & ~new_n3595_;
  assign new_n3597_ = ~new_n3556_ & ~new_n3596_;
  assign new_n3598_ = new_n3141_ & new_n3481_;
  assign new_n3599_ = ~new_n3547_ & new_n3598_;
  assign new_n3600_ = new_n3597_ & ~new_n3599_;
  assign new_n3601_ = pi0299 & ~new_n3600_;
  assign new_n3602_ = new_n3578_ & ~new_n3601_;
  assign new_n3603_ = pi0038 & new_n3602_;
  assign new_n3604_ = ~pi0100 & ~new_n3603_;
  assign new_n3605_ = ~new_n3592_ & new_n3604_;
  assign new_n3606_ = ~pi0228 & new_n3395_;
  assign new_n3607_ = ~new_n2449_ & new_n3131_;
  assign new_n3608_ = ~new_n3606_ & ~new_n3607_;
  assign new_n3609_ = ~pi0151 & new_n3608_;
  assign new_n3610_ = new_n3583_ & ~new_n3609_;
  assign new_n3611_ = new_n3548_ & ~new_n3610_;
  assign new_n3612_ = ~new_n3546_ & ~new_n3611_;
  assign new_n3613_ = ~pi0215 & ~new_n3612_;
  assign new_n3614_ = ~new_n3556_ & ~new_n3613_;
  assign new_n3615_ = pi0299 & ~new_n3614_;
  assign new_n3616_ = new_n3186_ & new_n3578_;
  assign new_n3617_ = ~new_n3615_ & new_n3616_;
  assign new_n3618_ = ~new_n3186_ & new_n3602_;
  assign new_n3619_ = pi0100 & ~new_n3618_;
  assign new_n3620_ = ~new_n3617_ & new_n3619_;
  assign new_n3621_ = ~new_n3605_ & ~new_n3620_;
  assign new_n3622_ = ~pi0087 & ~new_n3621_;
  assign new_n3623_ = ~new_n3212_ & new_n3602_;
  assign new_n3624_ = new_n3212_ & new_n3589_;
  assign new_n3625_ = ~new_n3623_ & ~new_n3624_;
  assign new_n3626_ = pi0087 & new_n3625_;
  assign new_n3627_ = ~pi0075 & ~new_n3626_;
  assign new_n3628_ = ~new_n3622_ & new_n3627_;
  assign new_n3629_ = pi0075 & new_n3602_;
  assign new_n3630_ = ~pi0092 & ~new_n3629_;
  assign new_n3631_ = ~new_n3628_ & new_n3630_;
  assign new_n3632_ = new_n3235_ & ~new_n3625_;
  assign new_n3633_ = ~new_n3235_ & new_n3602_;
  assign new_n3634_ = pi0092 & ~new_n3633_;
  assign new_n3635_ = ~new_n3632_ & new_n3634_;
  assign new_n3636_ = new_n3270_ & ~new_n3635_;
  assign new_n3637_ = ~new_n3631_ & new_n3636_;
  assign new_n3638_ = ~new_n3270_ & new_n3602_;
  assign new_n3639_ = ~pi0055 & ~new_n3638_;
  assign new_n3640_ = ~new_n3637_ & new_n3639_;
  assign new_n3641_ = new_n3273_ & new_n3587_;
  assign new_n3642_ = ~new_n3273_ & new_n3600_;
  assign new_n3643_ = pi0055 & ~new_n3642_;
  assign new_n3644_ = ~new_n3641_ & new_n3643_;
  assign new_n3645_ = ~pi0056 & ~new_n3644_;
  assign new_n3646_ = ~new_n3640_ & new_n3645_;
  assign new_n3647_ = new_n3285_ & ~new_n3587_;
  assign new_n3648_ = ~new_n3285_ & ~new_n3600_;
  assign new_n3649_ = pi0056 & ~new_n3648_;
  assign new_n3650_ = ~new_n3647_ & new_n3649_;
  assign new_n3651_ = ~pi0062 & ~new_n3650_;
  assign new_n3652_ = ~new_n3646_ & new_n3651_;
  assign new_n3653_ = new_n3438_ & new_n3587_;
  assign new_n3654_ = ~new_n3438_ & new_n3600_;
  assign new_n3655_ = pi0062 & ~new_n3654_;
  assign new_n3656_ = ~new_n3653_ & new_n3655_;
  assign new_n3657_ = pi0235 & new_n3436_;
  assign new_n3658_ = ~new_n3656_ & new_n3657_;
  assign new_n3659_ = ~new_n3652_ & new_n3658_;
  assign new_n3660_ = ~new_n3546_ & ~new_n3556_;
  assign new_n3661_ = new_n3327_ & new_n3660_;
  assign new_n3662_ = pi0299 & ~new_n3597_;
  assign new_n3663_ = ~new_n3661_ & new_n3662_;
  assign new_n3664_ = new_n3281_ & ~new_n3577_;
  assign new_n3665_ = ~new_n3663_ & new_n3664_;
  assign new_n3666_ = ~new_n3577_ & ~new_n3662_;
  assign new_n3667_ = ~new_n3212_ & new_n3666_;
  assign new_n3668_ = ~new_n3665_ & ~new_n3667_;
  assign new_n3669_ = pi0087 & ~new_n3668_;
  assign new_n3670_ = ~pi0100 & new_n3373_;
  assign new_n3671_ = ~pi0039 & pi0100;
  assign new_n3672_ = new_n3395_ & new_n3671_;
  assign new_n3673_ = ~new_n3670_ & ~new_n3672_;
  assign new_n3674_ = new_n3397_ & new_n3660_;
  assign new_n3675_ = ~new_n3673_ & new_n3674_;
  assign new_n3676_ = new_n3662_ & ~new_n3675_;
  assign new_n3677_ = ~pi0087 & ~new_n3577_;
  assign new_n3678_ = ~new_n3676_ & new_n3677_;
  assign new_n3679_ = ~new_n3669_ & ~new_n3678_;
  assign new_n3680_ = ~pi0075 & ~new_n3679_;
  assign new_n3681_ = pi0075 & new_n3666_;
  assign new_n3682_ = ~pi0092 & ~new_n3681_;
  assign new_n3683_ = ~new_n3680_ & new_n3682_;
  assign new_n3684_ = new_n3235_ & new_n3665_;
  assign new_n3685_ = ~new_n3413_ & new_n3666_;
  assign new_n3686_ = pi0092 & ~new_n3685_;
  assign new_n3687_ = ~new_n3684_ & new_n3686_;
  assign new_n3688_ = new_n3270_ & ~new_n3687_;
  assign new_n3689_ = ~new_n3683_ & new_n3688_;
  assign new_n3690_ = ~new_n3270_ & new_n3666_;
  assign new_n3691_ = ~pi0055 & ~new_n3690_;
  assign new_n3692_ = ~new_n3689_ & new_n3691_;
  assign new_n3693_ = new_n3273_ & new_n3661_;
  assign new_n3694_ = pi0055 & ~new_n3597_;
  assign new_n3695_ = ~new_n3693_ & new_n3694_;
  assign new_n3696_ = ~pi0056 & ~new_n3695_;
  assign new_n3697_ = ~new_n3692_ & new_n3696_;
  assign new_n3698_ = new_n3285_ & new_n3661_;
  assign new_n3699_ = ~new_n3597_ & ~new_n3698_;
  assign new_n3700_ = pi0056 & ~new_n3699_;
  assign new_n3701_ = ~pi0062 & ~new_n3700_;
  assign new_n3702_ = ~new_n3697_ & new_n3701_;
  assign new_n3703_ = ~pi0056 & new_n3698_;
  assign new_n3704_ = pi0062 & ~new_n3597_;
  assign new_n3705_ = ~new_n3703_ & new_n3704_;
  assign new_n3706_ = ~pi0235 & new_n3436_;
  assign new_n3707_ = ~new_n3705_ & new_n3706_;
  assign new_n3708_ = ~new_n3702_ & new_n3707_;
  assign new_n3709_ = pi0235 & new_n3599_;
  assign new_n3710_ = ~new_n3436_ & ~new_n3709_;
  assign new_n3711_ = new_n3597_ & new_n3710_;
  assign new_n3712_ = ~new_n3708_ & ~new_n3711_;
  assign po0155 = ~new_n3659_ & new_n3712_;
  assign new_n3714_ = pi0223 & pi1143;
  assign new_n3715_ = ~pi0299 & ~new_n3714_;
  assign new_n3716_ = ~pi0944 & new_n3045_;
  assign new_n3717_ = ~pi1143 & ~new_n3045_;
  assign new_n3718_ = pi0222 & ~new_n3717_;
  assign new_n3719_ = ~new_n3716_ & new_n3718_;
  assign new_n3720_ = pi0224 & pi0264;
  assign new_n3721_ = ~pi0222 & ~new_n3720_;
  assign new_n3722_ = ~pi0284 & new_n3448_;
  assign new_n3723_ = ~pi0224 & ~new_n3722_;
  assign new_n3724_ = new_n3721_ & ~new_n3723_;
  assign new_n3725_ = ~new_n3719_ & ~new_n3724_;
  assign new_n3726_ = ~new_n3448_ & new_n3721_;
  assign new_n3727_ = new_n3725_ & ~new_n3726_;
  assign new_n3728_ = ~pi0223 & ~new_n3727_;
  assign new_n3729_ = new_n3715_ & ~new_n3728_;
  assign new_n3730_ = ~pi0039 & ~new_n3729_;
  assign new_n3731_ = pi0215 & pi1143;
  assign new_n3732_ = pi0299 & ~new_n3731_;
  assign new_n3733_ = ~pi0944 & new_n2437_;
  assign new_n3734_ = ~pi1143 & ~new_n2437_;
  assign new_n3735_ = pi0221 & ~new_n3734_;
  assign new_n3736_ = ~new_n3733_ & new_n3735_;
  assign new_n3737_ = pi0216 & pi0264;
  assign new_n3738_ = ~pi0221 & ~new_n3737_;
  assign new_n3739_ = pi0284 & ~new_n2449_;
  assign new_n3740_ = pi0105 & ~new_n3739_;
  assign new_n3741_ = ~pi0105 & pi0146;
  assign new_n3742_ = pi0228 & ~new_n3741_;
  assign new_n3743_ = ~new_n3740_ & new_n3742_;
  assign new_n3744_ = ~new_n3469_ & new_n3743_;
  assign new_n3745_ = pi0146 & ~new_n3462_;
  assign new_n3746_ = ~pi0146 & new_n3471_;
  assign new_n3747_ = pi0284 & ~new_n3746_;
  assign new_n3748_ = ~new_n3745_ & new_n3747_;
  assign new_n3749_ = ~pi0146 & ~pi0284;
  assign new_n3750_ = ~new_n3371_ & new_n3749_;
  assign new_n3751_ = ~new_n3748_ & ~new_n3750_;
  assign new_n3752_ = ~pi0228 & ~new_n3751_;
  assign new_n3753_ = ~new_n3744_ & ~new_n3752_;
  assign new_n3754_ = ~pi0216 & ~new_n3753_;
  assign new_n3755_ = new_n3738_ & ~new_n3754_;
  assign new_n3756_ = ~new_n3736_ & ~new_n3755_;
  assign new_n3757_ = ~pi0215 & ~new_n3756_;
  assign new_n3758_ = new_n3732_ & ~new_n3757_;
  assign new_n3759_ = new_n3730_ & ~new_n3758_;
  assign new_n3760_ = ~pi0224 & new_n3739_;
  assign new_n3761_ = new_n3721_ & ~new_n3760_;
  assign new_n3762_ = ~new_n3719_ & ~new_n3761_;
  assign new_n3763_ = ~pi0223 & ~new_n3762_;
  assign new_n3764_ = ~new_n3714_ & ~new_n3763_;
  assign new_n3765_ = ~pi0299 & ~new_n3764_;
  assign new_n3766_ = pi0284 & new_n3100_;
  assign new_n3767_ = ~new_n3385_ & ~new_n3766_;
  assign new_n3768_ = ~pi0228 & ~new_n3767_;
  assign new_n3769_ = ~new_n3743_ & ~new_n3768_;
  assign new_n3770_ = ~pi0216 & ~new_n3769_;
  assign new_n3771_ = new_n3738_ & ~new_n3770_;
  assign new_n3772_ = ~new_n3736_ & ~new_n3771_;
  assign new_n3773_ = ~pi0215 & ~new_n3772_;
  assign new_n3774_ = ~new_n3731_ & ~new_n3773_;
  assign new_n3775_ = pi0299 & ~new_n3774_;
  assign new_n3776_ = ~new_n3765_ & ~new_n3775_;
  assign new_n3777_ = pi0039 & ~new_n3776_;
  assign new_n3778_ = ~pi0038 & ~new_n3777_;
  assign new_n3779_ = ~new_n3759_ & new_n3778_;
  assign new_n3780_ = ~new_n3481_ & ~new_n3743_;
  assign new_n3781_ = ~pi0146 & ~pi0228;
  assign new_n3782_ = new_n3780_ & ~new_n3781_;
  assign new_n3783_ = ~pi0216 & ~new_n3782_;
  assign new_n3784_ = new_n3738_ & ~new_n3783_;
  assign new_n3785_ = ~new_n3736_ & ~new_n3784_;
  assign new_n3786_ = ~pi0215 & ~new_n3785_;
  assign new_n3787_ = ~new_n3731_ & ~new_n3786_;
  assign new_n3788_ = new_n3598_ & ~new_n3737_;
  assign new_n3789_ = new_n3787_ & ~new_n3788_;
  assign new_n3790_ = pi0299 & ~new_n3789_;
  assign new_n3791_ = ~new_n3765_ & ~new_n3790_;
  assign new_n3792_ = pi0038 & new_n3791_;
  assign new_n3793_ = ~pi0100 & ~new_n3792_;
  assign new_n3794_ = ~new_n3779_ & new_n3793_;
  assign new_n3795_ = pi0252 & new_n2448_;
  assign new_n3796_ = ~pi0284 & ~new_n3795_;
  assign new_n3797_ = new_n3100_ & new_n3796_;
  assign new_n3798_ = ~pi0228 & ~new_n3797_;
  assign new_n3799_ = ~new_n3387_ & new_n3798_;
  assign new_n3800_ = ~new_n3743_ & ~new_n3799_;
  assign new_n3801_ = ~pi0216 & ~new_n3800_;
  assign new_n3802_ = new_n3738_ & ~new_n3801_;
  assign new_n3803_ = ~new_n3736_ & ~new_n3802_;
  assign new_n3804_ = ~pi0215 & ~new_n3803_;
  assign new_n3805_ = ~new_n3731_ & ~new_n3804_;
  assign new_n3806_ = pi0299 & ~new_n3805_;
  assign new_n3807_ = new_n3186_ & ~new_n3765_;
  assign new_n3808_ = ~new_n3806_ & new_n3807_;
  assign new_n3809_ = ~new_n3186_ & new_n3791_;
  assign new_n3810_ = pi0100 & ~new_n3809_;
  assign new_n3811_ = ~new_n3808_ & new_n3810_;
  assign new_n3812_ = ~new_n3794_ & ~new_n3811_;
  assign new_n3813_ = ~pi0087 & ~new_n3812_;
  assign new_n3814_ = ~new_n3212_ & new_n3791_;
  assign new_n3815_ = new_n3212_ & new_n3776_;
  assign new_n3816_ = ~new_n3814_ & ~new_n3815_;
  assign new_n3817_ = pi0087 & new_n3816_;
  assign new_n3818_ = ~pi0075 & ~new_n3817_;
  assign new_n3819_ = ~new_n3813_ & new_n3818_;
  assign new_n3820_ = pi0075 & new_n3791_;
  assign new_n3821_ = ~pi0092 & ~new_n3820_;
  assign new_n3822_ = ~new_n3819_ & new_n3821_;
  assign new_n3823_ = new_n3235_ & ~new_n3816_;
  assign new_n3824_ = ~new_n3235_ & new_n3791_;
  assign new_n3825_ = pi0092 & ~new_n3824_;
  assign new_n3826_ = ~new_n3823_ & new_n3825_;
  assign new_n3827_ = new_n3270_ & ~new_n3826_;
  assign new_n3828_ = ~new_n3822_ & new_n3827_;
  assign new_n3829_ = ~new_n3270_ & new_n3791_;
  assign new_n3830_ = ~pi0055 & ~new_n3829_;
  assign new_n3831_ = ~new_n3828_ & new_n3830_;
  assign new_n3832_ = new_n3273_ & new_n3774_;
  assign new_n3833_ = ~new_n3273_ & new_n3789_;
  assign new_n3834_ = pi0055 & ~new_n3833_;
  assign new_n3835_ = ~new_n3832_ & new_n3834_;
  assign new_n3836_ = ~pi0056 & ~new_n3835_;
  assign new_n3837_ = ~new_n3831_ & new_n3836_;
  assign new_n3838_ = new_n3285_ & ~new_n3774_;
  assign new_n3839_ = ~new_n3285_ & ~new_n3789_;
  assign new_n3840_ = pi0056 & ~new_n3839_;
  assign new_n3841_ = ~new_n3838_ & new_n3840_;
  assign new_n3842_ = ~pi0062 & ~new_n3841_;
  assign new_n3843_ = ~new_n3837_ & new_n3842_;
  assign new_n3844_ = new_n3438_ & new_n3774_;
  assign new_n3845_ = ~new_n3438_ & new_n3789_;
  assign new_n3846_ = pi0062 & ~new_n3845_;
  assign new_n3847_ = ~new_n3844_ & new_n3846_;
  assign new_n3848_ = pi0238 & new_n3436_;
  assign new_n3849_ = ~new_n3847_ & new_n3848_;
  assign new_n3850_ = ~new_n3843_ & new_n3849_;
  assign new_n3851_ = ~pi0146 & ~new_n3462_;
  assign new_n3852_ = pi0146 & new_n3471_;
  assign new_n3853_ = ~pi0284 & ~new_n3852_;
  assign new_n3854_ = pi0146 & pi0284;
  assign new_n3855_ = ~new_n3371_ & new_n3854_;
  assign new_n3856_ = ~new_n3853_ & ~new_n3855_;
  assign new_n3857_ = ~new_n3851_ & ~new_n3856_;
  assign new_n3858_ = ~pi0228 & ~new_n3857_;
  assign new_n3859_ = new_n3131_ & ~new_n3448_;
  assign new_n3860_ = ~new_n3743_ & ~new_n3859_;
  assign new_n3861_ = ~new_n3858_ & new_n3860_;
  assign new_n3862_ = ~pi0216 & ~new_n3861_;
  assign new_n3863_ = new_n3738_ & ~new_n3862_;
  assign new_n3864_ = ~new_n3736_ & ~new_n3863_;
  assign new_n3865_ = ~pi0215 & ~new_n3864_;
  assign new_n3866_ = new_n3732_ & ~new_n3865_;
  assign new_n3867_ = new_n3715_ & new_n3725_;
  assign new_n3868_ = new_n3730_ & ~new_n3867_;
  assign new_n3869_ = ~new_n3866_ & new_n3868_;
  assign new_n3870_ = new_n2449_ & new_n3105_;
  assign new_n3871_ = new_n3765_ & ~new_n3870_;
  assign new_n3872_ = ~new_n3768_ & new_n3780_;
  assign new_n3873_ = ~pi0216 & ~new_n3872_;
  assign new_n3874_ = new_n3738_ & ~new_n3873_;
  assign new_n3875_ = ~new_n3736_ & ~new_n3874_;
  assign new_n3876_ = ~pi0215 & ~new_n3875_;
  assign new_n3877_ = ~new_n3731_ & ~new_n3876_;
  assign new_n3878_ = pi0299 & ~new_n3877_;
  assign new_n3879_ = ~new_n3871_ & ~new_n3878_;
  assign new_n3880_ = pi0039 & ~new_n3879_;
  assign new_n3881_ = ~pi0038 & ~new_n3880_;
  assign new_n3882_ = ~new_n3869_ & new_n3881_;
  assign new_n3883_ = pi0299 & ~new_n3787_;
  assign new_n3884_ = ~new_n3871_ & ~new_n3883_;
  assign new_n3885_ = pi0038 & new_n3884_;
  assign new_n3886_ = ~pi0100 & ~new_n3885_;
  assign new_n3887_ = ~new_n3882_ & new_n3886_;
  assign new_n3888_ = new_n3780_ & ~new_n3799_;
  assign new_n3889_ = ~pi0216 & ~new_n3888_;
  assign new_n3890_ = new_n3738_ & ~new_n3889_;
  assign new_n3891_ = ~new_n3736_ & ~new_n3890_;
  assign new_n3892_ = ~pi0215 & ~new_n3891_;
  assign new_n3893_ = ~new_n3731_ & ~new_n3892_;
  assign new_n3894_ = pi0299 & ~new_n3893_;
  assign new_n3895_ = new_n3186_ & ~new_n3871_;
  assign new_n3896_ = ~new_n3894_ & new_n3895_;
  assign new_n3897_ = ~new_n3186_ & new_n3884_;
  assign new_n3898_ = pi0100 & ~new_n3897_;
  assign new_n3899_ = ~new_n3896_ & new_n3898_;
  assign new_n3900_ = ~new_n3887_ & ~new_n3899_;
  assign new_n3901_ = ~pi0087 & ~new_n3900_;
  assign new_n3902_ = ~new_n3212_ & new_n3884_;
  assign new_n3903_ = new_n3212_ & new_n3879_;
  assign new_n3904_ = ~new_n3902_ & ~new_n3903_;
  assign new_n3905_ = pi0087 & new_n3904_;
  assign new_n3906_ = ~pi0075 & ~new_n3905_;
  assign new_n3907_ = ~new_n3901_ & new_n3906_;
  assign new_n3908_ = pi0075 & new_n3884_;
  assign new_n3909_ = ~pi0092 & ~new_n3908_;
  assign new_n3910_ = ~new_n3907_ & new_n3909_;
  assign new_n3911_ = new_n3235_ & ~new_n3904_;
  assign new_n3912_ = ~new_n3235_ & new_n3884_;
  assign new_n3913_ = pi0092 & ~new_n3912_;
  assign new_n3914_ = ~new_n3911_ & new_n3913_;
  assign new_n3915_ = new_n3270_ & ~new_n3914_;
  assign new_n3916_ = ~new_n3910_ & new_n3915_;
  assign new_n3917_ = ~new_n3270_ & new_n3884_;
  assign new_n3918_ = ~pi0055 & ~new_n3917_;
  assign new_n3919_ = ~new_n3916_ & new_n3918_;
  assign new_n3920_ = new_n3273_ & new_n3877_;
  assign new_n3921_ = ~new_n3273_ & new_n3787_;
  assign new_n3922_ = pi0055 & ~new_n3921_;
  assign new_n3923_ = ~new_n3920_ & new_n3922_;
  assign new_n3924_ = ~pi0056 & ~new_n3923_;
  assign new_n3925_ = ~new_n3919_ & new_n3924_;
  assign new_n3926_ = new_n3285_ & ~new_n3877_;
  assign new_n3927_ = ~new_n3285_ & ~new_n3787_;
  assign new_n3928_ = pi0056 & ~new_n3927_;
  assign new_n3929_ = ~new_n3926_ & new_n3928_;
  assign new_n3930_ = ~pi0062 & ~new_n3929_;
  assign new_n3931_ = ~new_n3925_ & new_n3930_;
  assign new_n3932_ = new_n3438_ & new_n3877_;
  assign new_n3933_ = ~new_n3438_ & new_n3787_;
  assign new_n3934_ = pi0062 & ~new_n3933_;
  assign new_n3935_ = ~new_n3932_ & new_n3934_;
  assign new_n3936_ = ~pi0238 & new_n3436_;
  assign new_n3937_ = ~new_n3935_ & new_n3936_;
  assign new_n3938_ = ~new_n3931_ & new_n3937_;
  assign new_n3939_ = pi0238 & new_n3788_;
  assign new_n3940_ = ~new_n3436_ & ~new_n3939_;
  assign new_n3941_ = new_n3787_ & new_n3940_;
  assign new_n3942_ = ~new_n3938_ & ~new_n3941_;
  assign po0156 = ~new_n3850_ & new_n3942_;
  assign new_n3944_ = pi0215 & pi1142;
  assign new_n3945_ = pi0299 & ~new_n3944_;
  assign new_n3946_ = ~pi0932 & new_n2437_;
  assign new_n3947_ = ~pi1142 & ~new_n2437_;
  assign new_n3948_ = pi0221 & ~new_n3947_;
  assign new_n3949_ = ~new_n3946_ & new_n3948_;
  assign new_n3950_ = pi0216 & pi0277;
  assign new_n3951_ = ~pi0221 & ~new_n3950_;
  assign new_n3952_ = ~pi0262 & new_n3471_;
  assign new_n3953_ = ~pi0172 & ~new_n3952_;
  assign new_n3954_ = pi0172 & ~pi0262;
  assign new_n3955_ = new_n3462_ & new_n3954_;
  assign new_n3956_ = ~new_n3953_ & ~new_n3955_;
  assign new_n3957_ = pi0262 & new_n3371_;
  assign new_n3958_ = ~pi0228 & ~new_n3957_;
  assign new_n3959_ = ~new_n3956_ & new_n3958_;
  assign new_n3960_ = pi0262 & ~new_n2449_;
  assign new_n3961_ = pi0105 & new_n3960_;
  assign new_n3962_ = ~new_n3447_ & new_n3961_;
  assign new_n3963_ = ~pi0105 & pi0172;
  assign new_n3964_ = pi0228 & ~new_n3963_;
  assign new_n3965_ = ~new_n3962_ & new_n3964_;
  assign new_n3966_ = ~new_n3469_ & new_n3965_;
  assign new_n3967_ = ~pi0216 & ~new_n3966_;
  assign new_n3968_ = ~new_n3959_ & new_n3967_;
  assign new_n3969_ = new_n3951_ & ~new_n3968_;
  assign new_n3970_ = ~new_n3949_ & ~new_n3969_;
  assign new_n3971_ = ~pi0215 & ~new_n3970_;
  assign new_n3972_ = new_n3945_ & ~new_n3971_;
  assign new_n3973_ = pi0223 & pi1142;
  assign new_n3974_ = ~pi0299 & ~new_n3973_;
  assign new_n3975_ = ~pi0932 & new_n3045_;
  assign new_n3976_ = ~pi1142 & ~new_n3045_;
  assign new_n3977_ = pi0222 & ~new_n3976_;
  assign new_n3978_ = ~new_n3975_ & new_n3977_;
  assign new_n3979_ = pi0224 & pi0277;
  assign new_n3980_ = ~pi0222 & ~new_n3979_;
  assign new_n3981_ = ~pi0262 & new_n3448_;
  assign new_n3982_ = ~pi0224 & ~new_n3981_;
  assign new_n3983_ = new_n3980_ & ~new_n3982_;
  assign new_n3984_ = ~new_n3978_ & ~new_n3983_;
  assign new_n3985_ = new_n3974_ & new_n3984_;
  assign new_n3986_ = ~new_n3448_ & new_n3980_;
  assign new_n3987_ = new_n3984_ & ~new_n3986_;
  assign new_n3988_ = ~pi0223 & ~new_n3987_;
  assign new_n3989_ = new_n3974_ & ~new_n3988_;
  assign new_n3990_ = ~pi0039 & ~new_n3989_;
  assign new_n3991_ = ~new_n3985_ & new_n3990_;
  assign new_n3992_ = ~new_n3972_ & new_n3991_;
  assign new_n3993_ = ~pi0224 & new_n3960_;
  assign new_n3994_ = new_n3980_ & ~new_n3993_;
  assign new_n3995_ = ~new_n3978_ & ~new_n3994_;
  assign new_n3996_ = ~pi0223 & ~new_n3995_;
  assign new_n3997_ = ~new_n3973_ & ~new_n3996_;
  assign new_n3998_ = ~pi0299 & ~new_n3997_;
  assign new_n3999_ = ~new_n3870_ & new_n3998_;
  assign new_n4000_ = ~pi0262 & new_n3100_;
  assign new_n4001_ = pi0172 & ~pi0228;
  assign new_n4002_ = ~new_n3326_ & ~new_n4001_;
  assign new_n4003_ = ~new_n4000_ & ~new_n4002_;
  assign new_n4004_ = ~new_n3961_ & ~new_n3963_;
  assign new_n4005_ = pi0228 & ~new_n4004_;
  assign new_n4006_ = ~new_n3481_ & ~new_n4005_;
  assign new_n4007_ = ~new_n4003_ & new_n4006_;
  assign new_n4008_ = ~pi0216 & ~new_n4007_;
  assign new_n4009_ = new_n3951_ & ~new_n4008_;
  assign new_n4010_ = ~new_n3949_ & ~new_n4009_;
  assign new_n4011_ = ~pi0215 & ~new_n4010_;
  assign new_n4012_ = ~new_n3944_ & ~new_n4011_;
  assign new_n4013_ = pi0299 & ~new_n4012_;
  assign new_n4014_ = ~new_n3999_ & ~new_n4013_;
  assign new_n4015_ = pi0039 & ~new_n4014_;
  assign new_n4016_ = ~pi0038 & ~new_n4015_;
  assign new_n4017_ = ~new_n3992_ & new_n4016_;
  assign new_n4018_ = ~new_n4001_ & ~new_n4005_;
  assign new_n4019_ = ~pi0216 & ~new_n4018_;
  assign new_n4020_ = new_n3951_ & ~new_n4019_;
  assign new_n4021_ = ~new_n3949_ & ~new_n4020_;
  assign new_n4022_ = ~pi0215 & ~new_n4021_;
  assign new_n4023_ = ~new_n3944_ & ~new_n4022_;
  assign new_n4024_ = ~new_n3482_ & ~new_n4023_;
  assign new_n4025_ = pi0299 & new_n4024_;
  assign new_n4026_ = ~new_n3999_ & ~new_n4025_;
  assign new_n4027_ = pi0038 & new_n4026_;
  assign new_n4028_ = ~pi0100 & ~new_n4027_;
  assign new_n4029_ = ~new_n4017_ & new_n4028_;
  assign new_n4030_ = ~pi0262 & new_n3395_;
  assign new_n4031_ = ~new_n3606_ & ~new_n4001_;
  assign new_n4032_ = ~new_n4030_ & ~new_n4031_;
  assign new_n4033_ = new_n4006_ & ~new_n4032_;
  assign new_n4034_ = ~pi0216 & ~new_n4033_;
  assign new_n4035_ = new_n3951_ & ~new_n4034_;
  assign new_n4036_ = ~new_n3949_ & ~new_n4035_;
  assign new_n4037_ = ~pi0215 & ~new_n4036_;
  assign new_n4038_ = ~new_n3944_ & ~new_n4037_;
  assign new_n4039_ = pi0299 & ~new_n4038_;
  assign new_n4040_ = new_n3186_ & ~new_n3999_;
  assign new_n4041_ = ~new_n4039_ & new_n4040_;
  assign new_n4042_ = ~new_n3186_ & new_n4026_;
  assign new_n4043_ = pi0100 & ~new_n4042_;
  assign new_n4044_ = ~new_n4041_ & new_n4043_;
  assign new_n4045_ = ~new_n4029_ & ~new_n4044_;
  assign new_n4046_ = ~pi0087 & ~new_n4045_;
  assign new_n4047_ = ~new_n3212_ & new_n4026_;
  assign new_n4048_ = new_n3212_ & new_n4014_;
  assign new_n4049_ = ~new_n4047_ & ~new_n4048_;
  assign new_n4050_ = pi0087 & new_n4049_;
  assign new_n4051_ = ~pi0075 & ~new_n4050_;
  assign new_n4052_ = ~new_n4046_ & new_n4051_;
  assign new_n4053_ = pi0075 & new_n4026_;
  assign new_n4054_ = ~pi0092 & ~new_n4053_;
  assign new_n4055_ = ~new_n4052_ & new_n4054_;
  assign new_n4056_ = new_n3235_ & ~new_n4049_;
  assign new_n4057_ = ~new_n3235_ & new_n4026_;
  assign new_n4058_ = pi0092 & ~new_n4057_;
  assign new_n4059_ = ~new_n4056_ & new_n4058_;
  assign new_n4060_ = new_n3270_ & ~new_n4059_;
  assign new_n4061_ = ~new_n4055_ & new_n4060_;
  assign new_n4062_ = ~new_n3270_ & new_n4026_;
  assign new_n4063_ = ~pi0055 & ~new_n4062_;
  assign new_n4064_ = ~new_n4061_ & new_n4063_;
  assign new_n4065_ = new_n3273_ & new_n4012_;
  assign new_n4066_ = ~new_n3273_ & ~new_n4024_;
  assign new_n4067_ = pi0055 & ~new_n4066_;
  assign new_n4068_ = ~new_n4065_ & new_n4067_;
  assign new_n4069_ = ~pi0056 & ~new_n4068_;
  assign new_n4070_ = ~new_n4064_ & new_n4069_;
  assign new_n4071_ = new_n3285_ & ~new_n4012_;
  assign new_n4072_ = ~new_n3285_ & new_n4024_;
  assign new_n4073_ = pi0056 & ~new_n4072_;
  assign new_n4074_ = ~new_n4071_ & new_n4073_;
  assign new_n4075_ = ~pi0062 & ~new_n4074_;
  assign new_n4076_ = ~new_n4070_ & new_n4075_;
  assign new_n4077_ = new_n3438_ & new_n4012_;
  assign new_n4078_ = ~new_n3438_ & ~new_n4024_;
  assign new_n4079_ = pi0062 & ~new_n4078_;
  assign new_n4080_ = ~new_n4077_ & new_n4079_;
  assign new_n4081_ = new_n3436_ & ~new_n4080_;
  assign new_n4082_ = ~new_n4076_ & new_n4081_;
  assign new_n4083_ = ~new_n3436_ & ~new_n4024_;
  assign new_n4084_ = ~pi0249 & ~new_n4083_;
  assign new_n4085_ = ~new_n4082_ & new_n4084_;
  assign new_n4086_ = pi0262 & new_n3462_;
  assign new_n4087_ = ~pi0172 & ~new_n4086_;
  assign new_n4088_ = ~pi0262 & ~new_n3371_;
  assign new_n4089_ = pi0262 & ~new_n3471_;
  assign new_n4090_ = pi0172 & ~new_n4089_;
  assign new_n4091_ = ~new_n4088_ & new_n4090_;
  assign new_n4092_ = ~new_n4087_ & ~new_n4091_;
  assign new_n4093_ = ~pi0228 & ~new_n4092_;
  assign new_n4094_ = ~pi0216 & ~new_n3965_;
  assign new_n4095_ = ~new_n4093_ & new_n4094_;
  assign new_n4096_ = new_n3951_ & ~new_n4095_;
  assign new_n4097_ = ~new_n3949_ & ~new_n4096_;
  assign new_n4098_ = ~pi0215 & ~new_n4097_;
  assign new_n4099_ = new_n3945_ & ~new_n4098_;
  assign new_n4100_ = new_n3990_ & ~new_n4099_;
  assign new_n4101_ = ~new_n4003_ & ~new_n4005_;
  assign new_n4102_ = ~pi0216 & ~new_n4101_;
  assign new_n4103_ = new_n3951_ & ~new_n4102_;
  assign new_n4104_ = ~new_n3949_ & ~new_n4103_;
  assign new_n4105_ = ~pi0215 & ~new_n4104_;
  assign new_n4106_ = ~new_n3944_ & ~new_n4105_;
  assign new_n4107_ = pi0299 & ~new_n4106_;
  assign new_n4108_ = ~new_n3998_ & ~new_n4107_;
  assign new_n4109_ = pi0039 & ~new_n4108_;
  assign new_n4110_ = ~pi0038 & ~new_n4109_;
  assign new_n4111_ = ~new_n4100_ & new_n4110_;
  assign new_n4112_ = pi0299 & ~new_n4023_;
  assign new_n4113_ = ~new_n3998_ & ~new_n4112_;
  assign new_n4114_ = pi0038 & new_n4113_;
  assign new_n4115_ = ~pi0100 & ~new_n4114_;
  assign new_n4116_ = ~new_n4111_ & new_n4115_;
  assign new_n4117_ = ~new_n4005_ & ~new_n4032_;
  assign new_n4118_ = ~pi0216 & ~new_n4117_;
  assign new_n4119_ = new_n3951_ & ~new_n4118_;
  assign new_n4120_ = ~new_n3949_ & ~new_n4119_;
  assign new_n4121_ = ~pi0215 & ~new_n4120_;
  assign new_n4122_ = ~new_n3944_ & ~new_n4121_;
  assign new_n4123_ = pi0299 & ~new_n4122_;
  assign new_n4124_ = new_n3186_ & ~new_n3998_;
  assign new_n4125_ = ~new_n4123_ & new_n4124_;
  assign new_n4126_ = ~new_n3186_ & new_n4113_;
  assign new_n4127_ = pi0100 & ~new_n4126_;
  assign new_n4128_ = ~new_n4125_ & new_n4127_;
  assign new_n4129_ = ~new_n4116_ & ~new_n4128_;
  assign new_n4130_ = ~pi0087 & ~new_n4129_;
  assign new_n4131_ = ~new_n3212_ & new_n4113_;
  assign new_n4132_ = new_n3212_ & new_n4108_;
  assign new_n4133_ = ~new_n4131_ & ~new_n4132_;
  assign new_n4134_ = pi0087 & new_n4133_;
  assign new_n4135_ = ~pi0075 & ~new_n4134_;
  assign new_n4136_ = ~new_n4130_ & new_n4135_;
  assign new_n4137_ = pi0075 & new_n4113_;
  assign new_n4138_ = ~pi0092 & ~new_n4137_;
  assign new_n4139_ = ~new_n4136_ & new_n4138_;
  assign new_n4140_ = new_n3235_ & ~new_n4133_;
  assign new_n4141_ = ~new_n3235_ & new_n4113_;
  assign new_n4142_ = pi0092 & ~new_n4141_;
  assign new_n4143_ = ~new_n4140_ & new_n4142_;
  assign new_n4144_ = new_n3270_ & ~new_n4143_;
  assign new_n4145_ = ~new_n4139_ & new_n4144_;
  assign new_n4146_ = ~new_n3270_ & new_n4113_;
  assign new_n4147_ = ~pi0055 & ~new_n4146_;
  assign new_n4148_ = ~new_n4145_ & new_n4147_;
  assign new_n4149_ = new_n3273_ & new_n4106_;
  assign new_n4150_ = ~new_n3273_ & new_n4023_;
  assign new_n4151_ = pi0055 & ~new_n4150_;
  assign new_n4152_ = ~new_n4149_ & new_n4151_;
  assign new_n4153_ = ~pi0056 & ~new_n4152_;
  assign new_n4154_ = ~new_n4148_ & new_n4153_;
  assign new_n4155_ = new_n3285_ & ~new_n4106_;
  assign new_n4156_ = ~new_n3285_ & ~new_n4023_;
  assign new_n4157_ = pi0056 & ~new_n4156_;
  assign new_n4158_ = ~new_n4155_ & new_n4157_;
  assign new_n4159_ = ~pi0062 & ~new_n4158_;
  assign new_n4160_ = ~new_n4154_ & new_n4159_;
  assign new_n4161_ = new_n3438_ & new_n4106_;
  assign new_n4162_ = ~new_n3438_ & new_n4023_;
  assign new_n4163_ = pi0062 & ~new_n4162_;
  assign new_n4164_ = ~new_n4161_ & new_n4163_;
  assign new_n4165_ = new_n3436_ & ~new_n4164_;
  assign new_n4166_ = ~new_n4160_ & new_n4165_;
  assign new_n4167_ = ~new_n3436_ & new_n4023_;
  assign new_n4168_ = pi0249 & ~new_n4167_;
  assign new_n4169_ = ~new_n4166_ & new_n4168_;
  assign po0157 = new_n4085_ | new_n4169_;
  assign new_n4171_ = pi0215 & pi1141;
  assign new_n4172_ = pi0299 & ~new_n4171_;
  assign new_n4173_ = ~pi0935 & new_n2437_;
  assign new_n4174_ = ~pi1141 & ~new_n2437_;
  assign new_n4175_ = pi0221 & ~new_n4174_;
  assign new_n4176_ = ~new_n4173_ & new_n4175_;
  assign new_n4177_ = pi0216 & pi0270;
  assign new_n4178_ = ~pi0221 & ~new_n4177_;
  assign new_n4179_ = pi0861 & new_n3471_;
  assign new_n4180_ = ~pi0171 & ~new_n4179_;
  assign new_n4181_ = pi0171 & new_n3462_;
  assign new_n4182_ = ~new_n4180_ & ~new_n4181_;
  assign new_n4183_ = pi0861 & ~new_n4182_;
  assign new_n4184_ = ~new_n3371_ & new_n4180_;
  assign new_n4185_ = ~new_n4183_ & ~new_n4184_;
  assign new_n4186_ = ~pi0228 & ~new_n4185_;
  assign new_n4187_ = pi0861 & ~new_n2449_;
  assign new_n4188_ = pi0105 & ~new_n4187_;
  assign new_n4189_ = ~pi0105 & pi0171;
  assign new_n4190_ = pi0228 & ~new_n4189_;
  assign new_n4191_ = ~new_n4188_ & new_n4190_;
  assign new_n4192_ = ~new_n3469_ & new_n4191_;
  assign new_n4193_ = ~pi0216 & ~new_n4192_;
  assign new_n4194_ = ~new_n4186_ & new_n4193_;
  assign new_n4195_ = new_n4178_ & ~new_n4194_;
  assign new_n4196_ = ~new_n4176_ & ~new_n4195_;
  assign new_n4197_ = ~pi0215 & ~new_n4196_;
  assign new_n4198_ = new_n4172_ & ~new_n4197_;
  assign new_n4199_ = pi0223 & pi1141;
  assign new_n4200_ = ~pi0299 & ~new_n4199_;
  assign new_n4201_ = ~pi0935 & new_n3045_;
  assign new_n4202_ = ~pi1141 & ~new_n3045_;
  assign new_n4203_ = pi0222 & ~new_n4202_;
  assign new_n4204_ = ~new_n4201_ & new_n4203_;
  assign new_n4205_ = pi0224 & pi0270;
  assign new_n4206_ = ~pi0222 & ~new_n4205_;
  assign new_n4207_ = pi0861 & new_n3448_;
  assign new_n4208_ = ~pi0224 & ~new_n4207_;
  assign new_n4209_ = new_n4206_ & ~new_n4208_;
  assign new_n4210_ = ~new_n4204_ & ~new_n4209_;
  assign new_n4211_ = new_n4200_ & new_n4210_;
  assign new_n4212_ = ~new_n3448_ & new_n4206_;
  assign new_n4213_ = new_n4210_ & ~new_n4212_;
  assign new_n4214_ = ~pi0223 & ~new_n4213_;
  assign new_n4215_ = new_n4200_ & ~new_n4214_;
  assign new_n4216_ = ~pi0039 & ~new_n4215_;
  assign new_n4217_ = ~new_n4211_ & new_n4216_;
  assign new_n4218_ = ~new_n4198_ & new_n4217_;
  assign new_n4219_ = ~pi0224 & ~new_n4187_;
  assign new_n4220_ = new_n4206_ & ~new_n4219_;
  assign new_n4221_ = ~new_n4204_ & ~new_n4220_;
  assign new_n4222_ = ~pi0223 & ~new_n4221_;
  assign new_n4223_ = ~new_n4199_ & ~new_n4222_;
  assign new_n4224_ = ~pi0299 & ~new_n4223_;
  assign new_n4225_ = ~pi0216 & ~new_n4191_;
  assign new_n4226_ = pi0171 & ~new_n3100_;
  assign new_n4227_ = ~pi0861 & new_n3100_;
  assign new_n4228_ = ~pi0228 & ~new_n4227_;
  assign new_n4229_ = ~new_n4226_ & new_n4228_;
  assign new_n4230_ = new_n4225_ & ~new_n4229_;
  assign new_n4231_ = new_n4178_ & ~new_n4230_;
  assign new_n4232_ = ~new_n4176_ & ~new_n4231_;
  assign new_n4233_ = ~pi0215 & ~new_n4232_;
  assign new_n4234_ = ~new_n4171_ & ~new_n4233_;
  assign new_n4235_ = pi0299 & ~new_n4234_;
  assign new_n4236_ = ~new_n4224_ & ~new_n4235_;
  assign new_n4237_ = pi0039 & ~new_n4236_;
  assign new_n4238_ = ~pi0038 & ~new_n4237_;
  assign new_n4239_ = ~new_n4218_ & new_n4238_;
  assign new_n4240_ = ~pi0171 & ~pi0228;
  assign new_n4241_ = new_n4225_ & ~new_n4240_;
  assign new_n4242_ = new_n4178_ & ~new_n4241_;
  assign new_n4243_ = ~new_n4176_ & ~new_n4242_;
  assign new_n4244_ = ~pi0215 & ~new_n4243_;
  assign new_n4245_ = ~new_n4171_ & ~new_n4244_;
  assign new_n4246_ = pi0299 & ~new_n4245_;
  assign new_n4247_ = ~new_n4224_ & ~new_n4246_;
  assign new_n4248_ = pi0038 & new_n4247_;
  assign new_n4249_ = ~pi0100 & ~new_n4248_;
  assign new_n4250_ = ~new_n4239_ & new_n4249_;
  assign new_n4251_ = pi0171 & ~new_n3395_;
  assign new_n4252_ = ~pi0861 & new_n3395_;
  assign new_n4253_ = ~pi0228 & ~new_n4252_;
  assign new_n4254_ = ~new_n4251_ & new_n4253_;
  assign new_n4255_ = new_n4225_ & ~new_n4254_;
  assign new_n4256_ = new_n4178_ & ~new_n4255_;
  assign new_n4257_ = ~new_n4176_ & ~new_n4256_;
  assign new_n4258_ = ~pi0215 & ~new_n4257_;
  assign new_n4259_ = ~new_n4171_ & ~new_n4258_;
  assign new_n4260_ = pi0299 & ~new_n4259_;
  assign new_n4261_ = new_n3186_ & ~new_n4224_;
  assign new_n4262_ = ~new_n4260_ & new_n4261_;
  assign new_n4263_ = ~new_n3186_ & new_n4247_;
  assign new_n4264_ = pi0100 & ~new_n4263_;
  assign new_n4265_ = ~new_n4262_ & new_n4264_;
  assign new_n4266_ = ~new_n4250_ & ~new_n4265_;
  assign new_n4267_ = ~pi0087 & ~new_n4266_;
  assign new_n4268_ = ~new_n3212_ & new_n4247_;
  assign new_n4269_ = new_n3212_ & new_n4236_;
  assign new_n4270_ = ~new_n4268_ & ~new_n4269_;
  assign new_n4271_ = pi0087 & new_n4270_;
  assign new_n4272_ = ~pi0075 & ~new_n4271_;
  assign new_n4273_ = ~new_n4267_ & new_n4272_;
  assign new_n4274_ = pi0075 & new_n4247_;
  assign new_n4275_ = ~pi0092 & ~new_n4274_;
  assign new_n4276_ = ~new_n4273_ & new_n4275_;
  assign new_n4277_ = new_n3235_ & ~new_n4270_;
  assign new_n4278_ = ~new_n3235_ & new_n4247_;
  assign new_n4279_ = pi0092 & ~new_n4278_;
  assign new_n4280_ = ~new_n4277_ & new_n4279_;
  assign new_n4281_ = new_n3270_ & ~new_n4280_;
  assign new_n4282_ = ~new_n4276_ & new_n4281_;
  assign new_n4283_ = ~new_n3270_ & new_n4247_;
  assign new_n4284_ = ~pi0055 & ~new_n4283_;
  assign new_n4285_ = ~new_n4282_ & new_n4284_;
  assign new_n4286_ = new_n3273_ & new_n4234_;
  assign new_n4287_ = ~new_n3273_ & new_n4245_;
  assign new_n4288_ = pi0055 & ~new_n4287_;
  assign new_n4289_ = ~new_n4286_ & new_n4288_;
  assign new_n4290_ = ~pi0056 & ~new_n4289_;
  assign new_n4291_ = ~new_n4285_ & new_n4290_;
  assign new_n4292_ = new_n3285_ & ~new_n4234_;
  assign new_n4293_ = ~new_n3285_ & ~new_n4245_;
  assign new_n4294_ = pi0056 & ~new_n4293_;
  assign new_n4295_ = ~new_n4292_ & new_n4294_;
  assign new_n4296_ = ~pi0062 & ~new_n4295_;
  assign new_n4297_ = ~new_n4291_ & new_n4296_;
  assign new_n4298_ = new_n3438_ & new_n4234_;
  assign new_n4299_ = ~new_n3438_ & new_n4245_;
  assign new_n4300_ = pi0062 & ~new_n4299_;
  assign new_n4301_ = ~new_n4298_ & new_n4300_;
  assign new_n4302_ = ~pi0241 & new_n3436_;
  assign new_n4303_ = ~new_n4301_ & new_n4302_;
  assign new_n4304_ = ~new_n4297_ & new_n4303_;
  assign new_n4305_ = ~pi0861 & new_n3462_;
  assign new_n4306_ = ~pi0171 & ~new_n4305_;
  assign new_n4307_ = pi0861 & ~new_n3371_;
  assign new_n4308_ = ~pi0861 & ~new_n3471_;
  assign new_n4309_ = pi0171 & ~new_n4308_;
  assign new_n4310_ = ~new_n4307_ & new_n4309_;
  assign new_n4311_ = ~new_n4306_ & ~new_n4310_;
  assign new_n4312_ = ~pi0228 & ~new_n4311_;
  assign new_n4313_ = ~new_n3859_ & new_n4225_;
  assign new_n4314_ = ~new_n4312_ & new_n4313_;
  assign new_n4315_ = new_n4178_ & ~new_n4314_;
  assign new_n4316_ = ~new_n4176_ & ~new_n4315_;
  assign new_n4317_ = ~pi0215 & ~new_n4316_;
  assign new_n4318_ = new_n4172_ & ~new_n4317_;
  assign new_n4319_ = new_n4216_ & ~new_n4318_;
  assign new_n4320_ = ~new_n3491_ & ~new_n4224_;
  assign new_n4321_ = ~new_n3481_ & new_n4225_;
  assign new_n4322_ = ~new_n4229_ & new_n4321_;
  assign new_n4323_ = new_n4178_ & ~new_n4322_;
  assign new_n4324_ = ~new_n4176_ & ~new_n4323_;
  assign new_n4325_ = ~pi0215 & ~new_n4324_;
  assign new_n4326_ = ~new_n4171_ & ~new_n4325_;
  assign new_n4327_ = pi0299 & ~new_n4326_;
  assign new_n4328_ = new_n4320_ & ~new_n4327_;
  assign new_n4329_ = pi0039 & ~new_n4328_;
  assign new_n4330_ = ~pi0038 & ~new_n4329_;
  assign new_n4331_ = ~new_n4319_ & new_n4330_;
  assign new_n4332_ = new_n3598_ & ~new_n4177_;
  assign new_n4333_ = new_n4245_ & ~new_n4332_;
  assign new_n4334_ = pi0299 & ~new_n4333_;
  assign new_n4335_ = new_n4320_ & ~new_n4334_;
  assign new_n4336_ = pi0038 & new_n4335_;
  assign new_n4337_ = ~pi0100 & ~new_n4336_;
  assign new_n4338_ = ~new_n4331_ & new_n4337_;
  assign new_n4339_ = ~new_n4254_ & new_n4321_;
  assign new_n4340_ = new_n4178_ & ~new_n4339_;
  assign new_n4341_ = ~new_n4176_ & ~new_n4340_;
  assign new_n4342_ = ~pi0215 & ~new_n4341_;
  assign new_n4343_ = ~new_n4171_ & ~new_n4342_;
  assign new_n4344_ = pi0299 & ~new_n4343_;
  assign new_n4345_ = new_n3186_ & new_n4320_;
  assign new_n4346_ = ~new_n4344_ & new_n4345_;
  assign new_n4347_ = ~new_n3186_ & new_n4335_;
  assign new_n4348_ = pi0100 & ~new_n4347_;
  assign new_n4349_ = ~new_n4346_ & new_n4348_;
  assign new_n4350_ = ~new_n4338_ & ~new_n4349_;
  assign new_n4351_ = ~pi0087 & ~new_n4350_;
  assign new_n4352_ = ~new_n3212_ & new_n4335_;
  assign new_n4353_ = new_n3212_ & new_n4328_;
  assign new_n4354_ = ~new_n4352_ & ~new_n4353_;
  assign new_n4355_ = pi0087 & new_n4354_;
  assign new_n4356_ = ~pi0075 & ~new_n4355_;
  assign new_n4357_ = ~new_n4351_ & new_n4356_;
  assign new_n4358_ = pi0075 & new_n4335_;
  assign new_n4359_ = ~pi0092 & ~new_n4358_;
  assign new_n4360_ = ~new_n4357_ & new_n4359_;
  assign new_n4361_ = new_n3235_ & ~new_n4354_;
  assign new_n4362_ = ~new_n3235_ & new_n4335_;
  assign new_n4363_ = pi0092 & ~new_n4362_;
  assign new_n4364_ = ~new_n4361_ & new_n4363_;
  assign new_n4365_ = new_n3270_ & ~new_n4364_;
  assign new_n4366_ = ~new_n4360_ & new_n4365_;
  assign new_n4367_ = ~new_n3270_ & new_n4335_;
  assign new_n4368_ = ~pi0055 & ~new_n4367_;
  assign new_n4369_ = ~new_n4366_ & new_n4368_;
  assign new_n4370_ = new_n3273_ & new_n4326_;
  assign new_n4371_ = ~new_n3273_ & new_n4333_;
  assign new_n4372_ = pi0055 & ~new_n4371_;
  assign new_n4373_ = ~new_n4370_ & new_n4372_;
  assign new_n4374_ = ~pi0056 & ~new_n4373_;
  assign new_n4375_ = ~new_n4369_ & new_n4374_;
  assign new_n4376_ = new_n3285_ & ~new_n4326_;
  assign new_n4377_ = ~new_n3285_ & ~new_n4333_;
  assign new_n4378_ = pi0056 & ~new_n4377_;
  assign new_n4379_ = ~new_n4376_ & new_n4378_;
  assign new_n4380_ = ~pi0062 & ~new_n4379_;
  assign new_n4381_ = ~new_n4375_ & new_n4380_;
  assign new_n4382_ = new_n3438_ & new_n4326_;
  assign new_n4383_ = ~new_n3438_ & new_n4333_;
  assign new_n4384_ = pi0062 & ~new_n4383_;
  assign new_n4385_ = ~new_n4382_ & new_n4384_;
  assign new_n4386_ = pi0241 & new_n3436_;
  assign new_n4387_ = ~new_n4385_ & new_n4386_;
  assign new_n4388_ = ~new_n4381_ & new_n4387_;
  assign new_n4389_ = pi0241 & new_n4332_;
  assign new_n4390_ = ~new_n3436_ & ~new_n4389_;
  assign new_n4391_ = new_n4245_ & new_n4390_;
  assign new_n4392_ = ~new_n4388_ & ~new_n4391_;
  assign po0158 = ~new_n4304_ & new_n4392_;
  assign new_n4394_ = pi0215 & pi1140;
  assign new_n4395_ = pi0299 & ~new_n4394_;
  assign new_n4396_ = ~pi0921 & new_n2437_;
  assign new_n4397_ = ~pi1140 & ~new_n2437_;
  assign new_n4398_ = pi0221 & ~new_n4397_;
  assign new_n4399_ = ~new_n4396_ & new_n4398_;
  assign new_n4400_ = pi0216 & pi0282;
  assign new_n4401_ = ~pi0221 & ~new_n4400_;
  assign new_n4402_ = pi0869 & new_n3471_;
  assign new_n4403_ = ~pi0170 & ~new_n4402_;
  assign new_n4404_ = pi0170 & new_n3462_;
  assign new_n4405_ = ~new_n4403_ & ~new_n4404_;
  assign new_n4406_ = pi0869 & ~new_n4405_;
  assign new_n4407_ = ~new_n3371_ & new_n4403_;
  assign new_n4408_ = ~new_n4406_ & ~new_n4407_;
  assign new_n4409_ = ~pi0228 & ~new_n4408_;
  assign new_n4410_ = pi0869 & ~new_n2449_;
  assign new_n4411_ = pi0105 & ~new_n4410_;
  assign new_n4412_ = ~pi0105 & pi0170;
  assign new_n4413_ = pi0228 & ~new_n4412_;
  assign new_n4414_ = ~new_n4411_ & new_n4413_;
  assign new_n4415_ = ~new_n3469_ & new_n4414_;
  assign new_n4416_ = ~pi0216 & ~new_n4415_;
  assign new_n4417_ = ~new_n4409_ & new_n4416_;
  assign new_n4418_ = new_n4401_ & ~new_n4417_;
  assign new_n4419_ = ~new_n4399_ & ~new_n4418_;
  assign new_n4420_ = ~pi0215 & ~new_n4419_;
  assign new_n4421_ = new_n4395_ & ~new_n4420_;
  assign new_n4422_ = pi0223 & pi1140;
  assign new_n4423_ = ~pi0299 & ~new_n4422_;
  assign new_n4424_ = ~pi0921 & new_n3045_;
  assign new_n4425_ = ~pi1140 & ~new_n3045_;
  assign new_n4426_ = pi0222 & ~new_n4425_;
  assign new_n4427_ = ~new_n4424_ & new_n4426_;
  assign new_n4428_ = pi0224 & pi0282;
  assign new_n4429_ = ~pi0222 & ~new_n4428_;
  assign new_n4430_ = pi0869 & new_n3448_;
  assign new_n4431_ = ~pi0224 & ~new_n4430_;
  assign new_n4432_ = new_n4429_ & ~new_n4431_;
  assign new_n4433_ = ~new_n4427_ & ~new_n4432_;
  assign new_n4434_ = new_n4423_ & new_n4433_;
  assign new_n4435_ = ~new_n3448_ & new_n4429_;
  assign new_n4436_ = new_n4433_ & ~new_n4435_;
  assign new_n4437_ = ~pi0223 & ~new_n4436_;
  assign new_n4438_ = new_n4423_ & ~new_n4437_;
  assign new_n4439_ = ~pi0039 & ~new_n4438_;
  assign new_n4440_ = ~new_n4434_ & new_n4439_;
  assign new_n4441_ = ~new_n4421_ & new_n4440_;
  assign new_n4442_ = ~pi0224 & ~new_n4410_;
  assign new_n4443_ = new_n4429_ & ~new_n4442_;
  assign new_n4444_ = ~new_n4427_ & ~new_n4443_;
  assign new_n4445_ = ~pi0223 & ~new_n4444_;
  assign new_n4446_ = ~new_n4422_ & ~new_n4445_;
  assign new_n4447_ = ~pi0299 & ~new_n4446_;
  assign new_n4448_ = ~pi0216 & ~new_n4414_;
  assign new_n4449_ = pi0170 & ~new_n3100_;
  assign new_n4450_ = ~pi0869 & new_n3100_;
  assign new_n4451_ = ~pi0228 & ~new_n4450_;
  assign new_n4452_ = ~new_n4449_ & new_n4451_;
  assign new_n4453_ = new_n4448_ & ~new_n4452_;
  assign new_n4454_ = new_n4401_ & ~new_n4453_;
  assign new_n4455_ = ~new_n4399_ & ~new_n4454_;
  assign new_n4456_ = ~pi0215 & ~new_n4455_;
  assign new_n4457_ = ~new_n4394_ & ~new_n4456_;
  assign new_n4458_ = pi0299 & ~new_n4457_;
  assign new_n4459_ = ~new_n4447_ & ~new_n4458_;
  assign new_n4460_ = pi0039 & ~new_n4459_;
  assign new_n4461_ = ~pi0038 & ~new_n4460_;
  assign new_n4462_ = ~new_n4441_ & new_n4461_;
  assign new_n4463_ = ~pi0170 & ~pi0228;
  assign new_n4464_ = new_n4448_ & ~new_n4463_;
  assign new_n4465_ = new_n4401_ & ~new_n4464_;
  assign new_n4466_ = ~new_n4399_ & ~new_n4465_;
  assign new_n4467_ = ~pi0215 & ~new_n4466_;
  assign new_n4468_ = ~new_n4394_ & ~new_n4467_;
  assign new_n4469_ = pi0299 & ~new_n4468_;
  assign new_n4470_ = ~new_n4447_ & ~new_n4469_;
  assign new_n4471_ = pi0038 & new_n4470_;
  assign new_n4472_ = ~pi0100 & ~new_n4471_;
  assign new_n4473_ = ~new_n4462_ & new_n4472_;
  assign new_n4474_ = pi0170 & ~new_n3395_;
  assign new_n4475_ = ~pi0869 & new_n3395_;
  assign new_n4476_ = ~pi0228 & ~new_n4475_;
  assign new_n4477_ = ~new_n4474_ & new_n4476_;
  assign new_n4478_ = new_n4448_ & ~new_n4477_;
  assign new_n4479_ = new_n4401_ & ~new_n4478_;
  assign new_n4480_ = ~new_n4399_ & ~new_n4479_;
  assign new_n4481_ = ~pi0215 & ~new_n4480_;
  assign new_n4482_ = ~new_n4394_ & ~new_n4481_;
  assign new_n4483_ = pi0299 & ~new_n4482_;
  assign new_n4484_ = new_n3186_ & ~new_n4447_;
  assign new_n4485_ = ~new_n4483_ & new_n4484_;
  assign new_n4486_ = ~new_n3186_ & new_n4470_;
  assign new_n4487_ = pi0100 & ~new_n4486_;
  assign new_n4488_ = ~new_n4485_ & new_n4487_;
  assign new_n4489_ = ~new_n4473_ & ~new_n4488_;
  assign new_n4490_ = ~pi0087 & ~new_n4489_;
  assign new_n4491_ = ~new_n3212_ & new_n4470_;
  assign new_n4492_ = new_n3212_ & new_n4459_;
  assign new_n4493_ = ~new_n4491_ & ~new_n4492_;
  assign new_n4494_ = pi0087 & new_n4493_;
  assign new_n4495_ = ~pi0075 & ~new_n4494_;
  assign new_n4496_ = ~new_n4490_ & new_n4495_;
  assign new_n4497_ = pi0075 & new_n4470_;
  assign new_n4498_ = ~pi0092 & ~new_n4497_;
  assign new_n4499_ = ~new_n4496_ & new_n4498_;
  assign new_n4500_ = new_n3235_ & ~new_n4493_;
  assign new_n4501_ = ~new_n3235_ & new_n4470_;
  assign new_n4502_ = pi0092 & ~new_n4501_;
  assign new_n4503_ = ~new_n4500_ & new_n4502_;
  assign new_n4504_ = new_n3270_ & ~new_n4503_;
  assign new_n4505_ = ~new_n4499_ & new_n4504_;
  assign new_n4506_ = ~new_n3270_ & new_n4470_;
  assign new_n4507_ = ~pi0055 & ~new_n4506_;
  assign new_n4508_ = ~new_n4505_ & new_n4507_;
  assign new_n4509_ = new_n3273_ & new_n4457_;
  assign new_n4510_ = ~new_n3273_ & new_n4468_;
  assign new_n4511_ = pi0055 & ~new_n4510_;
  assign new_n4512_ = ~new_n4509_ & new_n4511_;
  assign new_n4513_ = ~pi0056 & ~new_n4512_;
  assign new_n4514_ = ~new_n4508_ & new_n4513_;
  assign new_n4515_ = new_n3285_ & ~new_n4457_;
  assign new_n4516_ = ~new_n3285_ & ~new_n4468_;
  assign new_n4517_ = pi0056 & ~new_n4516_;
  assign new_n4518_ = ~new_n4515_ & new_n4517_;
  assign new_n4519_ = ~pi0062 & ~new_n4518_;
  assign new_n4520_ = ~new_n4514_ & new_n4519_;
  assign new_n4521_ = new_n3438_ & new_n4457_;
  assign new_n4522_ = ~new_n3438_ & new_n4468_;
  assign new_n4523_ = pi0062 & ~new_n4522_;
  assign new_n4524_ = ~new_n4521_ & new_n4523_;
  assign new_n4525_ = ~pi0248 & new_n3436_;
  assign new_n4526_ = ~new_n4524_ & new_n4525_;
  assign new_n4527_ = ~new_n4520_ & new_n4526_;
  assign new_n4528_ = ~pi0869 & new_n3462_;
  assign new_n4529_ = ~pi0170 & ~new_n4528_;
  assign new_n4530_ = pi0869 & ~new_n3371_;
  assign new_n4531_ = ~pi0869 & ~new_n3471_;
  assign new_n4532_ = pi0170 & ~new_n4531_;
  assign new_n4533_ = ~new_n4530_ & new_n4532_;
  assign new_n4534_ = ~new_n4529_ & ~new_n4533_;
  assign new_n4535_ = ~pi0228 & ~new_n4534_;
  assign new_n4536_ = ~new_n3859_ & new_n4448_;
  assign new_n4537_ = ~new_n4535_ & new_n4536_;
  assign new_n4538_ = new_n4401_ & ~new_n4537_;
  assign new_n4539_ = ~new_n4399_ & ~new_n4538_;
  assign new_n4540_ = ~pi0215 & ~new_n4539_;
  assign new_n4541_ = new_n4395_ & ~new_n4540_;
  assign new_n4542_ = new_n4439_ & ~new_n4541_;
  assign new_n4543_ = ~new_n3491_ & ~new_n4447_;
  assign new_n4544_ = ~new_n3481_ & new_n4448_;
  assign new_n4545_ = ~new_n4452_ & new_n4544_;
  assign new_n4546_ = new_n4401_ & ~new_n4545_;
  assign new_n4547_ = ~new_n4399_ & ~new_n4546_;
  assign new_n4548_ = ~pi0215 & ~new_n4547_;
  assign new_n4549_ = ~new_n4394_ & ~new_n4548_;
  assign new_n4550_ = pi0299 & ~new_n4549_;
  assign new_n4551_ = new_n4543_ & ~new_n4550_;
  assign new_n4552_ = pi0039 & ~new_n4551_;
  assign new_n4553_ = ~pi0038 & ~new_n4552_;
  assign new_n4554_ = ~new_n4542_ & new_n4553_;
  assign new_n4555_ = new_n3598_ & ~new_n4400_;
  assign new_n4556_ = new_n4468_ & ~new_n4555_;
  assign new_n4557_ = pi0299 & ~new_n4556_;
  assign new_n4558_ = new_n4543_ & ~new_n4557_;
  assign new_n4559_ = pi0038 & new_n4558_;
  assign new_n4560_ = ~pi0100 & ~new_n4559_;
  assign new_n4561_ = ~new_n4554_ & new_n4560_;
  assign new_n4562_ = ~new_n4477_ & new_n4544_;
  assign new_n4563_ = new_n4401_ & ~new_n4562_;
  assign new_n4564_ = ~new_n4399_ & ~new_n4563_;
  assign new_n4565_ = ~pi0215 & ~new_n4564_;
  assign new_n4566_ = ~new_n4394_ & ~new_n4565_;
  assign new_n4567_ = pi0299 & ~new_n4566_;
  assign new_n4568_ = new_n3186_ & new_n4543_;
  assign new_n4569_ = ~new_n4567_ & new_n4568_;
  assign new_n4570_ = ~new_n3186_ & new_n4558_;
  assign new_n4571_ = pi0100 & ~new_n4570_;
  assign new_n4572_ = ~new_n4569_ & new_n4571_;
  assign new_n4573_ = ~new_n4561_ & ~new_n4572_;
  assign new_n4574_ = ~pi0087 & ~new_n4573_;
  assign new_n4575_ = ~new_n3212_ & new_n4558_;
  assign new_n4576_ = new_n3212_ & new_n4551_;
  assign new_n4577_ = ~new_n4575_ & ~new_n4576_;
  assign new_n4578_ = pi0087 & new_n4577_;
  assign new_n4579_ = ~pi0075 & ~new_n4578_;
  assign new_n4580_ = ~new_n4574_ & new_n4579_;
  assign new_n4581_ = pi0075 & new_n4558_;
  assign new_n4582_ = ~pi0092 & ~new_n4581_;
  assign new_n4583_ = ~new_n4580_ & new_n4582_;
  assign new_n4584_ = new_n3235_ & ~new_n4577_;
  assign new_n4585_ = ~new_n3235_ & new_n4558_;
  assign new_n4586_ = pi0092 & ~new_n4585_;
  assign new_n4587_ = ~new_n4584_ & new_n4586_;
  assign new_n4588_ = new_n3270_ & ~new_n4587_;
  assign new_n4589_ = ~new_n4583_ & new_n4588_;
  assign new_n4590_ = ~new_n3270_ & new_n4558_;
  assign new_n4591_ = ~pi0055 & ~new_n4590_;
  assign new_n4592_ = ~new_n4589_ & new_n4591_;
  assign new_n4593_ = new_n3273_ & new_n4549_;
  assign new_n4594_ = ~new_n3273_ & new_n4556_;
  assign new_n4595_ = pi0055 & ~new_n4594_;
  assign new_n4596_ = ~new_n4593_ & new_n4595_;
  assign new_n4597_ = ~pi0056 & ~new_n4596_;
  assign new_n4598_ = ~new_n4592_ & new_n4597_;
  assign new_n4599_ = new_n3285_ & ~new_n4549_;
  assign new_n4600_ = ~new_n3285_ & ~new_n4556_;
  assign new_n4601_ = pi0056 & ~new_n4600_;
  assign new_n4602_ = ~new_n4599_ & new_n4601_;
  assign new_n4603_ = ~pi0062 & ~new_n4602_;
  assign new_n4604_ = ~new_n4598_ & new_n4603_;
  assign new_n4605_ = new_n3438_ & new_n4549_;
  assign new_n4606_ = ~new_n3438_ & new_n4556_;
  assign new_n4607_ = pi0062 & ~new_n4606_;
  assign new_n4608_ = ~new_n4605_ & new_n4607_;
  assign new_n4609_ = pi0248 & new_n3436_;
  assign new_n4610_ = ~new_n4608_ & new_n4609_;
  assign new_n4611_ = ~new_n4604_ & new_n4610_;
  assign new_n4612_ = pi0248 & new_n4555_;
  assign new_n4613_ = ~new_n3436_ & ~new_n4612_;
  assign new_n4614_ = new_n4468_ & new_n4613_;
  assign new_n4615_ = ~new_n4611_ & ~new_n4614_;
  assign po0159 = ~new_n4527_ & new_n4615_;
  assign new_n4617_ = pi0216 & ~pi1139;
  assign new_n4618_ = ~pi0833 & pi1139;
  assign new_n4619_ = pi0833 & pi0920;
  assign new_n4620_ = ~pi0216 & ~new_n4619_;
  assign new_n4621_ = ~new_n4618_ & new_n4620_;
  assign new_n4622_ = pi0221 & ~new_n4621_;
  assign new_n4623_ = ~new_n4617_ & new_n4622_;
  assign new_n4624_ = pi0216 & pi0281;
  assign new_n4625_ = ~pi0221 & ~new_n4624_;
  assign new_n4626_ = ~pi0216 & ~pi0862;
  assign new_n4627_ = ~new_n3326_ & ~new_n3607_;
  assign new_n4628_ = new_n4626_ & ~new_n4627_;
  assign new_n4629_ = new_n4625_ & ~new_n4628_;
  assign new_n4630_ = ~new_n4623_ & ~new_n4629_;
  assign new_n4631_ = new_n3608_ & new_n4625_;
  assign new_n4632_ = new_n4630_ & ~new_n4631_;
  assign new_n4633_ = pi0148 & ~pi0215;
  assign new_n4634_ = ~pi0216 & ~new_n4622_;
  assign new_n4635_ = new_n3608_ & new_n4634_;
  assign new_n4636_ = new_n4633_ & ~new_n4635_;
  assign new_n4637_ = ~new_n4632_ & new_n4636_;
  assign new_n4638_ = pi0215 & pi1139;
  assign new_n4639_ = ~pi0148 & ~pi0215;
  assign new_n4640_ = ~new_n3131_ & ~new_n3326_;
  assign new_n4641_ = pi0862 & ~new_n3481_;
  assign new_n4642_ = ~pi0216 & ~new_n4641_;
  assign new_n4643_ = ~new_n4640_ & new_n4642_;
  assign new_n4644_ = new_n4625_ & ~new_n4643_;
  assign new_n4645_ = ~new_n4623_ & ~new_n4644_;
  assign new_n4646_ = ~new_n3131_ & ~new_n3606_;
  assign new_n4647_ = new_n4625_ & new_n4646_;
  assign new_n4648_ = new_n4645_ & ~new_n4647_;
  assign new_n4649_ = new_n4639_ & ~new_n4648_;
  assign new_n4650_ = ~new_n4638_ & ~new_n4649_;
  assign new_n4651_ = ~new_n4637_ & new_n4650_;
  assign new_n4652_ = pi0299 & ~new_n4651_;
  assign new_n4653_ = ~pi0920 & new_n3045_;
  assign new_n4654_ = ~pi1139 & ~new_n3045_;
  assign new_n4655_ = pi0222 & ~new_n4654_;
  assign new_n4656_ = ~new_n4653_ & new_n4655_;
  assign new_n4657_ = pi0223 & pi1139;
  assign new_n4658_ = ~pi0224 & ~new_n4657_;
  assign new_n4659_ = ~new_n4656_ & new_n4658_;
  assign new_n4660_ = new_n2449_ & new_n4659_;
  assign new_n4661_ = ~pi0862 & new_n4659_;
  assign new_n4662_ = pi0224 & pi0281;
  assign new_n4663_ = ~pi0222 & ~new_n4662_;
  assign new_n4664_ = ~new_n4656_ & ~new_n4663_;
  assign new_n4665_ = ~pi0223 & ~new_n4664_;
  assign new_n4666_ = ~new_n4657_ & ~new_n4665_;
  assign new_n4667_ = ~pi0299 & ~new_n4666_;
  assign new_n4668_ = ~new_n4661_ & new_n4667_;
  assign new_n4669_ = ~new_n4660_ & new_n4668_;
  assign new_n4670_ = new_n3186_ & ~new_n4669_;
  assign new_n4671_ = ~new_n4652_ & new_n4670_;
  assign new_n4672_ = new_n3607_ & new_n4626_;
  assign new_n4673_ = new_n4625_ & ~new_n4672_;
  assign new_n4674_ = ~new_n4623_ & ~new_n4673_;
  assign new_n4675_ = pi0148 & ~new_n3131_;
  assign new_n4676_ = new_n4634_ & new_n4675_;
  assign new_n4677_ = ~pi0215 & ~new_n4676_;
  assign new_n4678_ = ~new_n4674_ & new_n4677_;
  assign new_n4679_ = ~new_n4638_ & ~new_n4678_;
  assign new_n4680_ = ~new_n3482_ & ~new_n4679_;
  assign new_n4681_ = pi0299 & new_n4680_;
  assign new_n4682_ = ~new_n4669_ & ~new_n4681_;
  assign new_n4683_ = ~new_n3186_ & new_n4682_;
  assign new_n4684_ = pi0100 & ~new_n4683_;
  assign new_n4685_ = ~new_n4671_ & new_n4684_;
  assign new_n4686_ = ~pi0228 & new_n3371_;
  assign new_n4687_ = ~new_n3131_ & ~new_n4686_;
  assign new_n4688_ = ~pi0862 & new_n4687_;
  assign new_n4689_ = pi0862 & ~new_n3473_;
  assign new_n4690_ = ~pi0216 & ~new_n4689_;
  assign new_n4691_ = ~new_n4688_ & new_n4690_;
  assign new_n4692_ = new_n4625_ & ~new_n4691_;
  assign new_n4693_ = ~new_n4623_ & ~new_n4692_;
  assign new_n4694_ = new_n4639_ & ~new_n4693_;
  assign new_n4695_ = ~new_n3465_ & new_n4626_;
  assign new_n4696_ = new_n4625_ & ~new_n4695_;
  assign new_n4697_ = ~new_n4623_ & ~new_n4696_;
  assign new_n4698_ = new_n3465_ & new_n4634_;
  assign new_n4699_ = new_n4633_ & ~new_n4698_;
  assign new_n4700_ = ~new_n4697_ & new_n4699_;
  assign new_n4701_ = pi0299 & ~new_n4638_;
  assign new_n4702_ = ~new_n4700_ & new_n4701_;
  assign new_n4703_ = ~new_n4694_ & new_n4702_;
  assign new_n4704_ = ~new_n3448_ & new_n4659_;
  assign new_n4705_ = ~new_n4661_ & ~new_n4666_;
  assign new_n4706_ = ~new_n4704_ & new_n4705_;
  assign new_n4707_ = ~pi0299 & ~new_n4706_;
  assign new_n4708_ = ~pi0039 & ~new_n4707_;
  assign new_n4709_ = ~new_n4703_ & new_n4708_;
  assign new_n4710_ = new_n4639_ & ~new_n4645_;
  assign new_n4711_ = new_n4627_ & new_n4634_;
  assign new_n4712_ = new_n4633_ & ~new_n4711_;
  assign new_n4713_ = ~new_n4630_ & new_n4712_;
  assign new_n4714_ = ~new_n4638_ & ~new_n4713_;
  assign new_n4715_ = ~new_n4710_ & new_n4714_;
  assign new_n4716_ = pi0299 & ~new_n4715_;
  assign new_n4717_ = ~new_n4669_ & ~new_n4716_;
  assign new_n4718_ = pi0039 & ~new_n4717_;
  assign new_n4719_ = ~pi0038 & ~new_n4718_;
  assign new_n4720_ = ~new_n4709_ & new_n4719_;
  assign new_n4721_ = pi0038 & new_n4682_;
  assign new_n4722_ = ~pi0100 & ~new_n4721_;
  assign new_n4723_ = ~new_n4720_ & new_n4722_;
  assign new_n4724_ = ~new_n4685_ & ~new_n4723_;
  assign new_n4725_ = ~pi0087 & ~new_n4724_;
  assign new_n4726_ = ~new_n3212_ & new_n4682_;
  assign new_n4727_ = new_n3212_ & new_n4717_;
  assign new_n4728_ = ~new_n4726_ & ~new_n4727_;
  assign new_n4729_ = pi0087 & new_n4728_;
  assign new_n4730_ = ~pi0075 & ~new_n4729_;
  assign new_n4731_ = ~new_n4725_ & new_n4730_;
  assign new_n4732_ = pi0075 & new_n4682_;
  assign new_n4733_ = ~pi0092 & ~new_n4732_;
  assign new_n4734_ = ~new_n4731_ & new_n4733_;
  assign new_n4735_ = new_n3235_ & ~new_n4728_;
  assign new_n4736_ = ~new_n3235_ & new_n4682_;
  assign new_n4737_ = pi0092 & ~new_n4736_;
  assign new_n4738_ = ~new_n4735_ & new_n4737_;
  assign new_n4739_ = new_n3270_ & ~new_n4738_;
  assign new_n4740_ = ~new_n4734_ & new_n4739_;
  assign new_n4741_ = ~new_n3270_ & new_n4682_;
  assign new_n4742_ = ~pi0055 & ~new_n4741_;
  assign new_n4743_ = ~new_n4740_ & new_n4742_;
  assign new_n4744_ = new_n3273_ & new_n4715_;
  assign new_n4745_ = ~new_n3273_ & ~new_n4680_;
  assign new_n4746_ = pi0055 & ~new_n4745_;
  assign new_n4747_ = ~new_n4744_ & new_n4746_;
  assign new_n4748_ = ~pi0056 & ~new_n4747_;
  assign new_n4749_ = ~new_n4743_ & new_n4748_;
  assign new_n4750_ = new_n3285_ & ~new_n4715_;
  assign new_n4751_ = ~new_n3285_ & new_n4680_;
  assign new_n4752_ = pi0056 & ~new_n4751_;
  assign new_n4753_ = ~new_n4750_ & new_n4752_;
  assign new_n4754_ = ~pi0062 & ~new_n4753_;
  assign new_n4755_ = ~new_n4749_ & new_n4754_;
  assign new_n4756_ = new_n3438_ & new_n4715_;
  assign new_n4757_ = ~new_n3438_ & ~new_n4680_;
  assign new_n4758_ = pi0062 & ~new_n4757_;
  assign new_n4759_ = ~new_n4756_ & new_n4758_;
  assign new_n4760_ = new_n3436_ & ~new_n4759_;
  assign new_n4761_ = ~new_n4755_ & new_n4760_;
  assign new_n4762_ = ~new_n3436_ & ~new_n4680_;
  assign new_n4763_ = ~pi0247 & ~new_n4762_;
  assign new_n4764_ = ~new_n4761_ & new_n4763_;
  assign new_n4765_ = ~new_n4632_ & new_n4639_;
  assign new_n4766_ = ~pi0216 & ~new_n4623_;
  assign new_n4767_ = new_n4646_ & new_n4766_;
  assign new_n4768_ = ~new_n4630_ & new_n4633_;
  assign new_n4769_ = ~new_n4767_ & new_n4768_;
  assign new_n4770_ = ~new_n4638_ & ~new_n4769_;
  assign new_n4771_ = ~new_n4765_ & new_n4770_;
  assign new_n4772_ = pi0299 & ~new_n4771_;
  assign new_n4773_ = ~new_n3491_ & ~new_n4668_;
  assign new_n4774_ = new_n3186_ & new_n4773_;
  assign new_n4775_ = ~new_n4772_ & new_n4774_;
  assign new_n4776_ = pi0299 & ~new_n4679_;
  assign new_n4777_ = new_n4773_ & ~new_n4776_;
  assign new_n4778_ = ~new_n3186_ & new_n4777_;
  assign new_n4779_ = pi0100 & ~new_n4778_;
  assign new_n4780_ = ~new_n4775_ & new_n4779_;
  assign new_n4781_ = new_n3448_ & new_n4661_;
  assign new_n4782_ = new_n4667_ & ~new_n4781_;
  assign new_n4783_ = pi0862 & ~new_n4687_;
  assign new_n4784_ = ~pi0862 & new_n3473_;
  assign new_n4785_ = ~pi0216 & ~new_n4784_;
  assign new_n4786_ = ~new_n4783_ & new_n4785_;
  assign new_n4787_ = new_n4625_ & ~new_n4786_;
  assign new_n4788_ = ~new_n4623_ & ~new_n4787_;
  assign new_n4789_ = new_n4633_ & ~new_n4788_;
  assign new_n4790_ = new_n4639_ & ~new_n4697_;
  assign new_n4791_ = ~new_n4638_ & ~new_n4790_;
  assign new_n4792_ = ~new_n4789_ & new_n4791_;
  assign new_n4793_ = pi0299 & ~new_n4792_;
  assign new_n4794_ = ~new_n4782_ & ~new_n4793_;
  assign new_n4795_ = ~pi0039 & ~new_n4794_;
  assign new_n4796_ = ~new_n4630_ & new_n4677_;
  assign new_n4797_ = new_n4714_ & ~new_n4796_;
  assign new_n4798_ = pi0299 & ~new_n4797_;
  assign new_n4799_ = new_n4773_ & ~new_n4798_;
  assign new_n4800_ = pi0039 & ~new_n4799_;
  assign new_n4801_ = ~pi0038 & ~new_n4800_;
  assign new_n4802_ = ~new_n4795_ & new_n4801_;
  assign new_n4803_ = pi0038 & new_n4777_;
  assign new_n4804_ = ~pi0100 & ~new_n4803_;
  assign new_n4805_ = ~new_n4802_ & new_n4804_;
  assign new_n4806_ = ~new_n4780_ & ~new_n4805_;
  assign new_n4807_ = ~pi0087 & ~new_n4806_;
  assign new_n4808_ = ~new_n3212_ & new_n4777_;
  assign new_n4809_ = new_n3212_ & new_n4799_;
  assign new_n4810_ = ~new_n4808_ & ~new_n4809_;
  assign new_n4811_ = pi0087 & new_n4810_;
  assign new_n4812_ = ~pi0075 & ~new_n4811_;
  assign new_n4813_ = ~new_n4807_ & new_n4812_;
  assign new_n4814_ = pi0075 & new_n4777_;
  assign new_n4815_ = ~pi0092 & ~new_n4814_;
  assign new_n4816_ = ~new_n4813_ & new_n4815_;
  assign new_n4817_ = new_n3235_ & ~new_n4810_;
  assign new_n4818_ = ~new_n3235_ & new_n4777_;
  assign new_n4819_ = pi0092 & ~new_n4818_;
  assign new_n4820_ = ~new_n4817_ & new_n4819_;
  assign new_n4821_ = new_n3270_ & ~new_n4820_;
  assign new_n4822_ = ~new_n4816_ & new_n4821_;
  assign new_n4823_ = ~new_n3270_ & new_n4777_;
  assign new_n4824_ = ~pi0055 & ~new_n4823_;
  assign new_n4825_ = ~new_n4822_ & new_n4824_;
  assign new_n4826_ = new_n3273_ & new_n4797_;
  assign new_n4827_ = ~new_n3273_ & new_n4679_;
  assign new_n4828_ = pi0055 & ~new_n4827_;
  assign new_n4829_ = ~new_n4826_ & new_n4828_;
  assign new_n4830_ = ~pi0056 & ~new_n4829_;
  assign new_n4831_ = ~new_n4825_ & new_n4830_;
  assign new_n4832_ = new_n3285_ & ~new_n4797_;
  assign new_n4833_ = ~new_n3285_ & ~new_n4679_;
  assign new_n4834_ = pi0056 & ~new_n4833_;
  assign new_n4835_ = ~new_n4832_ & new_n4834_;
  assign new_n4836_ = ~pi0062 & ~new_n4835_;
  assign new_n4837_ = ~new_n4831_ & new_n4836_;
  assign new_n4838_ = new_n3438_ & new_n4797_;
  assign new_n4839_ = ~new_n3438_ & new_n4679_;
  assign new_n4840_ = pi0062 & ~new_n4839_;
  assign new_n4841_ = ~new_n4838_ & new_n4840_;
  assign new_n4842_ = new_n3436_ & ~new_n4841_;
  assign new_n4843_ = ~new_n4837_ & new_n4842_;
  assign new_n4844_ = ~new_n3436_ & new_n4679_;
  assign new_n4845_ = pi0247 & ~new_n4844_;
  assign new_n4846_ = ~new_n4843_ & new_n4845_;
  assign po0160 = new_n4764_ | new_n4846_;
  assign new_n4848_ = pi0215 & pi1138;
  assign new_n4849_ = pi0299 & ~new_n4848_;
  assign new_n4850_ = ~pi0940 & new_n2437_;
  assign new_n4851_ = ~pi1138 & ~new_n2437_;
  assign new_n4852_ = pi0221 & ~new_n4851_;
  assign new_n4853_ = ~new_n4850_ & new_n4852_;
  assign new_n4854_ = pi0216 & pi0269;
  assign new_n4855_ = ~pi0221 & ~new_n4854_;
  assign new_n4856_ = pi0877 & new_n3471_;
  assign new_n4857_ = ~pi0169 & ~new_n4856_;
  assign new_n4858_ = pi0169 & new_n3462_;
  assign new_n4859_ = ~new_n4857_ & ~new_n4858_;
  assign new_n4860_ = pi0877 & ~new_n4859_;
  assign new_n4861_ = ~new_n3371_ & new_n4857_;
  assign new_n4862_ = ~new_n4860_ & ~new_n4861_;
  assign new_n4863_ = ~pi0228 & ~new_n4862_;
  assign new_n4864_ = pi0877 & ~new_n2449_;
  assign new_n4865_ = pi0105 & ~new_n4864_;
  assign new_n4866_ = ~pi0105 & pi0169;
  assign new_n4867_ = pi0228 & ~new_n4866_;
  assign new_n4868_ = ~new_n4865_ & new_n4867_;
  assign new_n4869_ = ~new_n3469_ & new_n4868_;
  assign new_n4870_ = ~pi0216 & ~new_n4869_;
  assign new_n4871_ = ~new_n4863_ & new_n4870_;
  assign new_n4872_ = new_n4855_ & ~new_n4871_;
  assign new_n4873_ = ~new_n4853_ & ~new_n4872_;
  assign new_n4874_ = ~pi0215 & ~new_n4873_;
  assign new_n4875_ = new_n4849_ & ~new_n4874_;
  assign new_n4876_ = pi0223 & pi1138;
  assign new_n4877_ = ~pi0299 & ~new_n4876_;
  assign new_n4878_ = ~pi0940 & new_n3045_;
  assign new_n4879_ = ~pi1138 & ~new_n3045_;
  assign new_n4880_ = pi0222 & ~new_n4879_;
  assign new_n4881_ = ~new_n4878_ & new_n4880_;
  assign new_n4882_ = pi0224 & pi0269;
  assign new_n4883_ = ~pi0222 & ~new_n4882_;
  assign new_n4884_ = pi0877 & new_n3448_;
  assign new_n4885_ = ~pi0224 & ~new_n4884_;
  assign new_n4886_ = new_n4883_ & ~new_n4885_;
  assign new_n4887_ = ~new_n4881_ & ~new_n4886_;
  assign new_n4888_ = new_n4877_ & new_n4887_;
  assign new_n4889_ = ~new_n3448_ & new_n4883_;
  assign new_n4890_ = new_n4887_ & ~new_n4889_;
  assign new_n4891_ = ~pi0223 & ~new_n4890_;
  assign new_n4892_ = new_n4877_ & ~new_n4891_;
  assign new_n4893_ = ~pi0039 & ~new_n4892_;
  assign new_n4894_ = ~new_n4888_ & new_n4893_;
  assign new_n4895_ = ~new_n4875_ & new_n4894_;
  assign new_n4896_ = ~pi0224 & ~new_n4864_;
  assign new_n4897_ = new_n4883_ & ~new_n4896_;
  assign new_n4898_ = ~new_n4881_ & ~new_n4897_;
  assign new_n4899_ = ~pi0223 & ~new_n4898_;
  assign new_n4900_ = ~new_n4876_ & ~new_n4899_;
  assign new_n4901_ = ~pi0299 & ~new_n4900_;
  assign new_n4902_ = ~pi0216 & ~new_n4868_;
  assign new_n4903_ = pi0169 & ~new_n3100_;
  assign new_n4904_ = ~pi0877 & new_n3100_;
  assign new_n4905_ = ~pi0228 & ~new_n4904_;
  assign new_n4906_ = ~new_n4903_ & new_n4905_;
  assign new_n4907_ = new_n4902_ & ~new_n4906_;
  assign new_n4908_ = new_n4855_ & ~new_n4907_;
  assign new_n4909_ = ~new_n4853_ & ~new_n4908_;
  assign new_n4910_ = ~pi0215 & ~new_n4909_;
  assign new_n4911_ = ~new_n4848_ & ~new_n4910_;
  assign new_n4912_ = pi0299 & ~new_n4911_;
  assign new_n4913_ = ~new_n4901_ & ~new_n4912_;
  assign new_n4914_ = pi0039 & ~new_n4913_;
  assign new_n4915_ = ~pi0038 & ~new_n4914_;
  assign new_n4916_ = ~new_n4895_ & new_n4915_;
  assign new_n4917_ = ~pi0169 & ~pi0228;
  assign new_n4918_ = new_n4902_ & ~new_n4917_;
  assign new_n4919_ = new_n4855_ & ~new_n4918_;
  assign new_n4920_ = ~new_n4853_ & ~new_n4919_;
  assign new_n4921_ = ~pi0215 & ~new_n4920_;
  assign new_n4922_ = ~new_n4848_ & ~new_n4921_;
  assign new_n4923_ = pi0299 & ~new_n4922_;
  assign new_n4924_ = ~new_n4901_ & ~new_n4923_;
  assign new_n4925_ = pi0038 & new_n4924_;
  assign new_n4926_ = ~pi0100 & ~new_n4925_;
  assign new_n4927_ = ~new_n4916_ & new_n4926_;
  assign new_n4928_ = pi0169 & ~new_n3395_;
  assign new_n4929_ = ~pi0877 & new_n3395_;
  assign new_n4930_ = ~pi0228 & ~new_n4929_;
  assign new_n4931_ = ~new_n4928_ & new_n4930_;
  assign new_n4932_ = new_n4902_ & ~new_n4931_;
  assign new_n4933_ = new_n4855_ & ~new_n4932_;
  assign new_n4934_ = ~new_n4853_ & ~new_n4933_;
  assign new_n4935_ = ~pi0215 & ~new_n4934_;
  assign new_n4936_ = ~new_n4848_ & ~new_n4935_;
  assign new_n4937_ = pi0299 & ~new_n4936_;
  assign new_n4938_ = new_n3186_ & ~new_n4901_;
  assign new_n4939_ = ~new_n4937_ & new_n4938_;
  assign new_n4940_ = ~new_n3186_ & new_n4924_;
  assign new_n4941_ = pi0100 & ~new_n4940_;
  assign new_n4942_ = ~new_n4939_ & new_n4941_;
  assign new_n4943_ = ~new_n4927_ & ~new_n4942_;
  assign new_n4944_ = ~pi0087 & ~new_n4943_;
  assign new_n4945_ = ~new_n3212_ & new_n4924_;
  assign new_n4946_ = new_n3212_ & new_n4913_;
  assign new_n4947_ = ~new_n4945_ & ~new_n4946_;
  assign new_n4948_ = pi0087 & new_n4947_;
  assign new_n4949_ = ~pi0075 & ~new_n4948_;
  assign new_n4950_ = ~new_n4944_ & new_n4949_;
  assign new_n4951_ = pi0075 & new_n4924_;
  assign new_n4952_ = ~pi0092 & ~new_n4951_;
  assign new_n4953_ = ~new_n4950_ & new_n4952_;
  assign new_n4954_ = new_n3235_ & ~new_n4947_;
  assign new_n4955_ = ~new_n3235_ & new_n4924_;
  assign new_n4956_ = pi0092 & ~new_n4955_;
  assign new_n4957_ = ~new_n4954_ & new_n4956_;
  assign new_n4958_ = new_n3270_ & ~new_n4957_;
  assign new_n4959_ = ~new_n4953_ & new_n4958_;
  assign new_n4960_ = ~new_n3270_ & new_n4924_;
  assign new_n4961_ = ~pi0055 & ~new_n4960_;
  assign new_n4962_ = ~new_n4959_ & new_n4961_;
  assign new_n4963_ = new_n3273_ & new_n4911_;
  assign new_n4964_ = ~new_n3273_ & new_n4922_;
  assign new_n4965_ = pi0055 & ~new_n4964_;
  assign new_n4966_ = ~new_n4963_ & new_n4965_;
  assign new_n4967_ = ~pi0056 & ~new_n4966_;
  assign new_n4968_ = ~new_n4962_ & new_n4967_;
  assign new_n4969_ = new_n3285_ & ~new_n4911_;
  assign new_n4970_ = ~new_n3285_ & ~new_n4922_;
  assign new_n4971_ = pi0056 & ~new_n4970_;
  assign new_n4972_ = ~new_n4969_ & new_n4971_;
  assign new_n4973_ = ~pi0062 & ~new_n4972_;
  assign new_n4974_ = ~new_n4968_ & new_n4973_;
  assign new_n4975_ = new_n3438_ & new_n4911_;
  assign new_n4976_ = ~new_n3438_ & new_n4922_;
  assign new_n4977_ = pi0062 & ~new_n4976_;
  assign new_n4978_ = ~new_n4975_ & new_n4977_;
  assign new_n4979_ = ~pi0246 & new_n3436_;
  assign new_n4980_ = ~new_n4978_ & new_n4979_;
  assign new_n4981_ = ~new_n4974_ & new_n4980_;
  assign new_n4982_ = ~pi0877 & new_n3462_;
  assign new_n4983_ = ~pi0169 & ~new_n4982_;
  assign new_n4984_ = pi0877 & ~new_n3371_;
  assign new_n4985_ = ~pi0877 & ~new_n3471_;
  assign new_n4986_ = pi0169 & ~new_n4985_;
  assign new_n4987_ = ~new_n4984_ & new_n4986_;
  assign new_n4988_ = ~new_n4983_ & ~new_n4987_;
  assign new_n4989_ = ~pi0228 & ~new_n4988_;
  assign new_n4990_ = ~new_n3859_ & new_n4902_;
  assign new_n4991_ = ~new_n4989_ & new_n4990_;
  assign new_n4992_ = new_n4855_ & ~new_n4991_;
  assign new_n4993_ = ~new_n4853_ & ~new_n4992_;
  assign new_n4994_ = ~pi0215 & ~new_n4993_;
  assign new_n4995_ = new_n4849_ & ~new_n4994_;
  assign new_n4996_ = new_n4893_ & ~new_n4995_;
  assign new_n4997_ = ~new_n3491_ & ~new_n4901_;
  assign new_n4998_ = ~new_n3481_ & new_n4902_;
  assign new_n4999_ = ~new_n4906_ & new_n4998_;
  assign new_n5000_ = new_n4855_ & ~new_n4999_;
  assign new_n5001_ = ~new_n4853_ & ~new_n5000_;
  assign new_n5002_ = ~pi0215 & ~new_n5001_;
  assign new_n5003_ = ~new_n4848_ & ~new_n5002_;
  assign new_n5004_ = pi0299 & ~new_n5003_;
  assign new_n5005_ = new_n4997_ & ~new_n5004_;
  assign new_n5006_ = pi0039 & ~new_n5005_;
  assign new_n5007_ = ~pi0038 & ~new_n5006_;
  assign new_n5008_ = ~new_n4996_ & new_n5007_;
  assign new_n5009_ = new_n3598_ & ~new_n4854_;
  assign new_n5010_ = new_n4922_ & ~new_n5009_;
  assign new_n5011_ = pi0299 & ~new_n5010_;
  assign new_n5012_ = new_n4997_ & ~new_n5011_;
  assign new_n5013_ = pi0038 & new_n5012_;
  assign new_n5014_ = ~pi0100 & ~new_n5013_;
  assign new_n5015_ = ~new_n5008_ & new_n5014_;
  assign new_n5016_ = ~new_n4931_ & new_n4998_;
  assign new_n5017_ = new_n4855_ & ~new_n5016_;
  assign new_n5018_ = ~new_n4853_ & ~new_n5017_;
  assign new_n5019_ = ~pi0215 & ~new_n5018_;
  assign new_n5020_ = ~new_n4848_ & ~new_n5019_;
  assign new_n5021_ = pi0299 & ~new_n5020_;
  assign new_n5022_ = new_n3186_ & new_n4997_;
  assign new_n5023_ = ~new_n5021_ & new_n5022_;
  assign new_n5024_ = ~new_n3186_ & new_n5012_;
  assign new_n5025_ = pi0100 & ~new_n5024_;
  assign new_n5026_ = ~new_n5023_ & new_n5025_;
  assign new_n5027_ = ~new_n5015_ & ~new_n5026_;
  assign new_n5028_ = ~pi0087 & ~new_n5027_;
  assign new_n5029_ = ~new_n3212_ & new_n5012_;
  assign new_n5030_ = new_n3212_ & new_n5005_;
  assign new_n5031_ = ~new_n5029_ & ~new_n5030_;
  assign new_n5032_ = pi0087 & new_n5031_;
  assign new_n5033_ = ~pi0075 & ~new_n5032_;
  assign new_n5034_ = ~new_n5028_ & new_n5033_;
  assign new_n5035_ = pi0075 & new_n5012_;
  assign new_n5036_ = ~pi0092 & ~new_n5035_;
  assign new_n5037_ = ~new_n5034_ & new_n5036_;
  assign new_n5038_ = new_n3235_ & ~new_n5031_;
  assign new_n5039_ = ~new_n3235_ & new_n5012_;
  assign new_n5040_ = pi0092 & ~new_n5039_;
  assign new_n5041_ = ~new_n5038_ & new_n5040_;
  assign new_n5042_ = new_n3270_ & ~new_n5041_;
  assign new_n5043_ = ~new_n5037_ & new_n5042_;
  assign new_n5044_ = ~new_n3270_ & new_n5012_;
  assign new_n5045_ = ~pi0055 & ~new_n5044_;
  assign new_n5046_ = ~new_n5043_ & new_n5045_;
  assign new_n5047_ = new_n3273_ & new_n5003_;
  assign new_n5048_ = ~new_n3273_ & new_n5010_;
  assign new_n5049_ = pi0055 & ~new_n5048_;
  assign new_n5050_ = ~new_n5047_ & new_n5049_;
  assign new_n5051_ = ~pi0056 & ~new_n5050_;
  assign new_n5052_ = ~new_n5046_ & new_n5051_;
  assign new_n5053_ = new_n3285_ & ~new_n5003_;
  assign new_n5054_ = ~new_n3285_ & ~new_n5010_;
  assign new_n5055_ = pi0056 & ~new_n5054_;
  assign new_n5056_ = ~new_n5053_ & new_n5055_;
  assign new_n5057_ = ~pi0062 & ~new_n5056_;
  assign new_n5058_ = ~new_n5052_ & new_n5057_;
  assign new_n5059_ = new_n3438_ & new_n5003_;
  assign new_n5060_ = ~new_n3438_ & new_n5010_;
  assign new_n5061_ = pi0062 & ~new_n5060_;
  assign new_n5062_ = ~new_n5059_ & new_n5061_;
  assign new_n5063_ = pi0246 & new_n3436_;
  assign new_n5064_ = ~new_n5062_ & new_n5063_;
  assign new_n5065_ = ~new_n5058_ & new_n5064_;
  assign new_n5066_ = pi0246 & new_n5009_;
  assign new_n5067_ = ~new_n3436_ & ~new_n5066_;
  assign new_n5068_ = new_n4922_ & new_n5067_;
  assign new_n5069_ = ~new_n5065_ & ~new_n5068_;
  assign po0161 = ~new_n4981_ & new_n5069_;
  assign new_n5071_ = pi0215 & pi1137;
  assign new_n5072_ = pi0299 & ~new_n5071_;
  assign new_n5073_ = ~pi0933 & new_n2437_;
  assign new_n5074_ = ~pi1137 & ~new_n2437_;
  assign new_n5075_ = pi0221 & ~new_n5074_;
  assign new_n5076_ = ~new_n5073_ & new_n5075_;
  assign new_n5077_ = pi0216 & pi0280;
  assign new_n5078_ = ~pi0221 & ~new_n5077_;
  assign new_n5079_ = pi0878 & new_n3471_;
  assign new_n5080_ = ~pi0168 & ~new_n5079_;
  assign new_n5081_ = pi0168 & new_n3462_;
  assign new_n5082_ = ~new_n5080_ & ~new_n5081_;
  assign new_n5083_ = pi0878 & ~new_n5082_;
  assign new_n5084_ = ~new_n3371_ & new_n5080_;
  assign new_n5085_ = ~new_n5083_ & ~new_n5084_;
  assign new_n5086_ = ~pi0228 & ~new_n5085_;
  assign new_n5087_ = pi0878 & ~new_n2449_;
  assign new_n5088_ = pi0105 & ~new_n5087_;
  assign new_n5089_ = ~pi0105 & pi0168;
  assign new_n5090_ = pi0228 & ~new_n5089_;
  assign new_n5091_ = ~new_n5088_ & new_n5090_;
  assign new_n5092_ = ~new_n3469_ & new_n5091_;
  assign new_n5093_ = ~pi0216 & ~new_n5092_;
  assign new_n5094_ = ~new_n5086_ & new_n5093_;
  assign new_n5095_ = new_n5078_ & ~new_n5094_;
  assign new_n5096_ = ~new_n5076_ & ~new_n5095_;
  assign new_n5097_ = ~pi0215 & ~new_n5096_;
  assign new_n5098_ = new_n5072_ & ~new_n5097_;
  assign new_n5099_ = pi0223 & pi1137;
  assign new_n5100_ = ~pi0299 & ~new_n5099_;
  assign new_n5101_ = ~pi0933 & new_n3045_;
  assign new_n5102_ = ~pi1137 & ~new_n3045_;
  assign new_n5103_ = pi0222 & ~new_n5102_;
  assign new_n5104_ = ~new_n5101_ & new_n5103_;
  assign new_n5105_ = pi0224 & pi0280;
  assign new_n5106_ = ~pi0222 & ~new_n5105_;
  assign new_n5107_ = pi0878 & new_n3448_;
  assign new_n5108_ = ~pi0224 & ~new_n5107_;
  assign new_n5109_ = new_n5106_ & ~new_n5108_;
  assign new_n5110_ = ~new_n5104_ & ~new_n5109_;
  assign new_n5111_ = new_n5100_ & new_n5110_;
  assign new_n5112_ = ~new_n3448_ & new_n5106_;
  assign new_n5113_ = new_n5110_ & ~new_n5112_;
  assign new_n5114_ = ~pi0223 & ~new_n5113_;
  assign new_n5115_ = new_n5100_ & ~new_n5114_;
  assign new_n5116_ = ~pi0039 & ~new_n5115_;
  assign new_n5117_ = ~new_n5111_ & new_n5116_;
  assign new_n5118_ = ~new_n5098_ & new_n5117_;
  assign new_n5119_ = ~pi0224 & ~new_n5087_;
  assign new_n5120_ = new_n5106_ & ~new_n5119_;
  assign new_n5121_ = ~new_n5104_ & ~new_n5120_;
  assign new_n5122_ = ~pi0223 & ~new_n5121_;
  assign new_n5123_ = ~new_n5099_ & ~new_n5122_;
  assign new_n5124_ = ~pi0299 & ~new_n5123_;
  assign new_n5125_ = ~pi0216 & ~new_n5091_;
  assign new_n5126_ = pi0168 & ~new_n3100_;
  assign new_n5127_ = ~pi0878 & new_n3100_;
  assign new_n5128_ = ~pi0228 & ~new_n5127_;
  assign new_n5129_ = ~new_n5126_ & new_n5128_;
  assign new_n5130_ = new_n5125_ & ~new_n5129_;
  assign new_n5131_ = new_n5078_ & ~new_n5130_;
  assign new_n5132_ = ~new_n5076_ & ~new_n5131_;
  assign new_n5133_ = ~pi0215 & ~new_n5132_;
  assign new_n5134_ = ~new_n5071_ & ~new_n5133_;
  assign new_n5135_ = pi0299 & ~new_n5134_;
  assign new_n5136_ = ~new_n5124_ & ~new_n5135_;
  assign new_n5137_ = pi0039 & ~new_n5136_;
  assign new_n5138_ = ~pi0038 & ~new_n5137_;
  assign new_n5139_ = ~new_n5118_ & new_n5138_;
  assign new_n5140_ = ~pi0168 & ~pi0228;
  assign new_n5141_ = new_n5125_ & ~new_n5140_;
  assign new_n5142_ = new_n5078_ & ~new_n5141_;
  assign new_n5143_ = ~new_n5076_ & ~new_n5142_;
  assign new_n5144_ = ~pi0215 & ~new_n5143_;
  assign new_n5145_ = ~new_n5071_ & ~new_n5144_;
  assign new_n5146_ = pi0299 & ~new_n5145_;
  assign new_n5147_ = ~new_n5124_ & ~new_n5146_;
  assign new_n5148_ = pi0038 & new_n5147_;
  assign new_n5149_ = ~pi0100 & ~new_n5148_;
  assign new_n5150_ = ~new_n5139_ & new_n5149_;
  assign new_n5151_ = pi0168 & ~new_n3395_;
  assign new_n5152_ = ~pi0878 & new_n3395_;
  assign new_n5153_ = ~pi0228 & ~new_n5152_;
  assign new_n5154_ = ~new_n5151_ & new_n5153_;
  assign new_n5155_ = new_n5125_ & ~new_n5154_;
  assign new_n5156_ = new_n5078_ & ~new_n5155_;
  assign new_n5157_ = ~new_n5076_ & ~new_n5156_;
  assign new_n5158_ = ~pi0215 & ~new_n5157_;
  assign new_n5159_ = ~new_n5071_ & ~new_n5158_;
  assign new_n5160_ = pi0299 & ~new_n5159_;
  assign new_n5161_ = new_n3186_ & ~new_n5124_;
  assign new_n5162_ = ~new_n5160_ & new_n5161_;
  assign new_n5163_ = ~new_n3186_ & new_n5147_;
  assign new_n5164_ = pi0100 & ~new_n5163_;
  assign new_n5165_ = ~new_n5162_ & new_n5164_;
  assign new_n5166_ = ~new_n5150_ & ~new_n5165_;
  assign new_n5167_ = ~pi0087 & ~new_n5166_;
  assign new_n5168_ = ~new_n3212_ & new_n5147_;
  assign new_n5169_ = new_n3212_ & new_n5136_;
  assign new_n5170_ = ~new_n5168_ & ~new_n5169_;
  assign new_n5171_ = pi0087 & new_n5170_;
  assign new_n5172_ = ~pi0075 & ~new_n5171_;
  assign new_n5173_ = ~new_n5167_ & new_n5172_;
  assign new_n5174_ = pi0075 & new_n5147_;
  assign new_n5175_ = ~pi0092 & ~new_n5174_;
  assign new_n5176_ = ~new_n5173_ & new_n5175_;
  assign new_n5177_ = new_n3235_ & ~new_n5170_;
  assign new_n5178_ = ~new_n3235_ & new_n5147_;
  assign new_n5179_ = pi0092 & ~new_n5178_;
  assign new_n5180_ = ~new_n5177_ & new_n5179_;
  assign new_n5181_ = new_n3270_ & ~new_n5180_;
  assign new_n5182_ = ~new_n5176_ & new_n5181_;
  assign new_n5183_ = ~new_n3270_ & new_n5147_;
  assign new_n5184_ = ~pi0055 & ~new_n5183_;
  assign new_n5185_ = ~new_n5182_ & new_n5184_;
  assign new_n5186_ = new_n3273_ & new_n5134_;
  assign new_n5187_ = ~new_n3273_ & new_n5145_;
  assign new_n5188_ = pi0055 & ~new_n5187_;
  assign new_n5189_ = ~new_n5186_ & new_n5188_;
  assign new_n5190_ = ~pi0056 & ~new_n5189_;
  assign new_n5191_ = ~new_n5185_ & new_n5190_;
  assign new_n5192_ = new_n3285_ & ~new_n5134_;
  assign new_n5193_ = ~new_n3285_ & ~new_n5145_;
  assign new_n5194_ = pi0056 & ~new_n5193_;
  assign new_n5195_ = ~new_n5192_ & new_n5194_;
  assign new_n5196_ = ~pi0062 & ~new_n5195_;
  assign new_n5197_ = ~new_n5191_ & new_n5196_;
  assign new_n5198_ = new_n3438_ & new_n5134_;
  assign new_n5199_ = ~new_n3438_ & new_n5145_;
  assign new_n5200_ = pi0062 & ~new_n5199_;
  assign new_n5201_ = ~new_n5198_ & new_n5200_;
  assign new_n5202_ = ~pi0240 & new_n3436_;
  assign new_n5203_ = ~new_n5201_ & new_n5202_;
  assign new_n5204_ = ~new_n5197_ & new_n5203_;
  assign new_n5205_ = ~pi0878 & new_n3462_;
  assign new_n5206_ = ~pi0168 & ~new_n5205_;
  assign new_n5207_ = pi0878 & ~new_n3371_;
  assign new_n5208_ = ~pi0878 & ~new_n3471_;
  assign new_n5209_ = pi0168 & ~new_n5208_;
  assign new_n5210_ = ~new_n5207_ & new_n5209_;
  assign new_n5211_ = ~new_n5206_ & ~new_n5210_;
  assign new_n5212_ = ~pi0228 & ~new_n5211_;
  assign new_n5213_ = ~new_n3859_ & new_n5125_;
  assign new_n5214_ = ~new_n5212_ & new_n5213_;
  assign new_n5215_ = new_n5078_ & ~new_n5214_;
  assign new_n5216_ = ~new_n5076_ & ~new_n5215_;
  assign new_n5217_ = ~pi0215 & ~new_n5216_;
  assign new_n5218_ = new_n5072_ & ~new_n5217_;
  assign new_n5219_ = new_n5116_ & ~new_n5218_;
  assign new_n5220_ = ~new_n3491_ & ~new_n5124_;
  assign new_n5221_ = ~new_n3481_ & new_n5125_;
  assign new_n5222_ = ~new_n5129_ & new_n5221_;
  assign new_n5223_ = new_n5078_ & ~new_n5222_;
  assign new_n5224_ = ~new_n5076_ & ~new_n5223_;
  assign new_n5225_ = ~pi0215 & ~new_n5224_;
  assign new_n5226_ = ~new_n5071_ & ~new_n5225_;
  assign new_n5227_ = pi0299 & ~new_n5226_;
  assign new_n5228_ = new_n5220_ & ~new_n5227_;
  assign new_n5229_ = pi0039 & ~new_n5228_;
  assign new_n5230_ = ~pi0038 & ~new_n5229_;
  assign new_n5231_ = ~new_n5219_ & new_n5230_;
  assign new_n5232_ = new_n3598_ & ~new_n5077_;
  assign new_n5233_ = new_n5145_ & ~new_n5232_;
  assign new_n5234_ = pi0299 & ~new_n5233_;
  assign new_n5235_ = new_n5220_ & ~new_n5234_;
  assign new_n5236_ = pi0038 & new_n5235_;
  assign new_n5237_ = ~pi0100 & ~new_n5236_;
  assign new_n5238_ = ~new_n5231_ & new_n5237_;
  assign new_n5239_ = ~new_n5154_ & new_n5221_;
  assign new_n5240_ = new_n5078_ & ~new_n5239_;
  assign new_n5241_ = ~new_n5076_ & ~new_n5240_;
  assign new_n5242_ = ~pi0215 & ~new_n5241_;
  assign new_n5243_ = ~new_n5071_ & ~new_n5242_;
  assign new_n5244_ = pi0299 & ~new_n5243_;
  assign new_n5245_ = new_n3186_ & new_n5220_;
  assign new_n5246_ = ~new_n5244_ & new_n5245_;
  assign new_n5247_ = ~new_n3186_ & new_n5235_;
  assign new_n5248_ = pi0100 & ~new_n5247_;
  assign new_n5249_ = ~new_n5246_ & new_n5248_;
  assign new_n5250_ = ~new_n5238_ & ~new_n5249_;
  assign new_n5251_ = ~pi0087 & ~new_n5250_;
  assign new_n5252_ = ~new_n3212_ & new_n5235_;
  assign new_n5253_ = new_n3212_ & new_n5228_;
  assign new_n5254_ = ~new_n5252_ & ~new_n5253_;
  assign new_n5255_ = pi0087 & new_n5254_;
  assign new_n5256_ = ~pi0075 & ~new_n5255_;
  assign new_n5257_ = ~new_n5251_ & new_n5256_;
  assign new_n5258_ = pi0075 & new_n5235_;
  assign new_n5259_ = ~pi0092 & ~new_n5258_;
  assign new_n5260_ = ~new_n5257_ & new_n5259_;
  assign new_n5261_ = new_n3235_ & ~new_n5254_;
  assign new_n5262_ = ~new_n3235_ & new_n5235_;
  assign new_n5263_ = pi0092 & ~new_n5262_;
  assign new_n5264_ = ~new_n5261_ & new_n5263_;
  assign new_n5265_ = new_n3270_ & ~new_n5264_;
  assign new_n5266_ = ~new_n5260_ & new_n5265_;
  assign new_n5267_ = ~new_n3270_ & new_n5235_;
  assign new_n5268_ = ~pi0055 & ~new_n5267_;
  assign new_n5269_ = ~new_n5266_ & new_n5268_;
  assign new_n5270_ = new_n3273_ & new_n5226_;
  assign new_n5271_ = ~new_n3273_ & new_n5233_;
  assign new_n5272_ = pi0055 & ~new_n5271_;
  assign new_n5273_ = ~new_n5270_ & new_n5272_;
  assign new_n5274_ = ~pi0056 & ~new_n5273_;
  assign new_n5275_ = ~new_n5269_ & new_n5274_;
  assign new_n5276_ = new_n3285_ & ~new_n5226_;
  assign new_n5277_ = ~new_n3285_ & ~new_n5233_;
  assign new_n5278_ = pi0056 & ~new_n5277_;
  assign new_n5279_ = ~new_n5276_ & new_n5278_;
  assign new_n5280_ = ~pi0062 & ~new_n5279_;
  assign new_n5281_ = ~new_n5275_ & new_n5280_;
  assign new_n5282_ = new_n3438_ & new_n5226_;
  assign new_n5283_ = ~new_n3438_ & new_n5233_;
  assign new_n5284_ = pi0062 & ~new_n5283_;
  assign new_n5285_ = ~new_n5282_ & new_n5284_;
  assign new_n5286_ = pi0240 & new_n3436_;
  assign new_n5287_ = ~new_n5285_ & new_n5286_;
  assign new_n5288_ = ~new_n5281_ & new_n5287_;
  assign new_n5289_ = pi0240 & new_n5232_;
  assign new_n5290_ = ~new_n3436_ & ~new_n5289_;
  assign new_n5291_ = new_n5145_ & new_n5290_;
  assign new_n5292_ = ~new_n5288_ & ~new_n5291_;
  assign po0162 = ~new_n5204_ & new_n5292_;
  assign new_n5294_ = ~pi0928 & new_n2437_;
  assign new_n5295_ = ~pi1136 & ~new_n2437_;
  assign new_n5296_ = pi0221 & ~new_n5295_;
  assign new_n5297_ = ~new_n5294_ & new_n5296_;
  assign new_n5298_ = pi0216 & pi0266;
  assign new_n5299_ = pi0875 & ~new_n2449_;
  assign new_n5300_ = pi0105 & ~new_n5299_;
  assign new_n5301_ = ~pi0105 & ~pi0166;
  assign new_n5302_ = ~new_n5300_ & ~new_n5301_;
  assign new_n5303_ = new_n3470_ & ~new_n5302_;
  assign new_n5304_ = ~pi0216 & ~new_n5303_;
  assign new_n5305_ = ~pi0166 & ~new_n3462_;
  assign new_n5306_ = pi0166 & new_n3471_;
  assign new_n5307_ = pi0875 & ~new_n5306_;
  assign new_n5308_ = ~new_n5305_ & new_n5307_;
  assign new_n5309_ = pi0166 & ~pi0875;
  assign new_n5310_ = ~new_n3371_ & new_n5309_;
  assign new_n5311_ = ~new_n5308_ & ~new_n5310_;
  assign new_n5312_ = ~pi0228 & ~new_n5311_;
  assign new_n5313_ = ~new_n3470_ & ~new_n5312_;
  assign new_n5314_ = new_n5304_ & ~new_n5313_;
  assign new_n5315_ = ~new_n5298_ & ~new_n5314_;
  assign new_n5316_ = ~pi0221 & ~new_n5315_;
  assign new_n5317_ = ~new_n5297_ & ~new_n5316_;
  assign new_n5318_ = ~pi0215 & ~new_n5317_;
  assign new_n5319_ = pi0215 & pi1136;
  assign new_n5320_ = pi0299 & ~new_n5319_;
  assign new_n5321_ = ~new_n5318_ & new_n5320_;
  assign new_n5322_ = ~pi0224 & ~pi0875;
  assign new_n5323_ = ~new_n2449_ & new_n5322_;
  assign new_n5324_ = pi0224 & ~pi0266;
  assign new_n5325_ = ~pi0222 & ~new_n5324_;
  assign new_n5326_ = ~new_n5323_ & new_n5325_;
  assign new_n5327_ = new_n3057_ & ~new_n3448_;
  assign new_n5328_ = new_n5326_ & ~new_n5327_;
  assign new_n5329_ = ~pi0928 & new_n3045_;
  assign new_n5330_ = ~pi1136 & ~new_n3045_;
  assign new_n5331_ = pi0222 & ~new_n5330_;
  assign new_n5332_ = ~new_n5329_ & new_n5331_;
  assign new_n5333_ = pi0223 & pi1136;
  assign new_n5334_ = ~pi0299 & ~new_n5333_;
  assign new_n5335_ = ~new_n5332_ & new_n5334_;
  assign new_n5336_ = ~new_n5328_ & new_n5335_;
  assign new_n5337_ = ~new_n5326_ & ~new_n5332_;
  assign new_n5338_ = ~new_n5327_ & new_n5337_;
  assign new_n5339_ = ~pi0223 & ~new_n5338_;
  assign new_n5340_ = new_n5334_ & ~new_n5339_;
  assign new_n5341_ = ~pi0039 & ~new_n5340_;
  assign new_n5342_ = ~new_n5336_ & new_n5341_;
  assign new_n5343_ = ~new_n5321_ & new_n5342_;
  assign new_n5344_ = ~pi0223 & ~new_n5337_;
  assign new_n5345_ = ~new_n5333_ & ~new_n5344_;
  assign new_n5346_ = ~pi0299 & ~new_n5345_;
  assign new_n5347_ = new_n3105_ & ~new_n5299_;
  assign new_n5348_ = new_n5346_ & ~new_n5347_;
  assign new_n5349_ = pi0228 & new_n5302_;
  assign new_n5350_ = ~pi0875 & new_n3100_;
  assign new_n5351_ = ~pi0166 & ~new_n3100_;
  assign new_n5352_ = ~pi0228 & ~new_n5351_;
  assign new_n5353_ = ~new_n5350_ & new_n5352_;
  assign new_n5354_ = ~new_n5349_ & ~new_n5353_;
  assign new_n5355_ = ~pi0216 & ~new_n5354_;
  assign new_n5356_ = ~new_n5298_ & ~new_n5355_;
  assign new_n5357_ = ~pi0221 & ~new_n5356_;
  assign new_n5358_ = ~new_n5297_ & ~new_n5357_;
  assign new_n5359_ = ~pi0215 & ~new_n5358_;
  assign new_n5360_ = ~new_n5319_ & ~new_n5359_;
  assign new_n5361_ = pi0299 & ~new_n5360_;
  assign new_n5362_ = ~new_n5348_ & ~new_n5361_;
  assign new_n5363_ = pi0039 & ~new_n5362_;
  assign new_n5364_ = ~pi0038 & ~new_n5363_;
  assign new_n5365_ = ~new_n5343_ & new_n5364_;
  assign new_n5366_ = pi0166 & ~pi0228;
  assign new_n5367_ = ~new_n5349_ & ~new_n5366_;
  assign new_n5368_ = ~pi0216 & ~new_n5367_;
  assign new_n5369_ = ~new_n5298_ & ~new_n5368_;
  assign new_n5370_ = ~pi0221 & ~new_n5369_;
  assign new_n5371_ = ~new_n5297_ & ~new_n5370_;
  assign new_n5372_ = ~pi0215 & ~new_n5371_;
  assign new_n5373_ = ~new_n5319_ & ~new_n5372_;
  assign new_n5374_ = pi0299 & ~new_n5373_;
  assign new_n5375_ = ~new_n5348_ & ~new_n5374_;
  assign new_n5376_ = pi0038 & new_n5375_;
  assign new_n5377_ = ~pi0100 & ~new_n5376_;
  assign new_n5378_ = ~new_n5365_ & new_n5377_;
  assign new_n5379_ = ~pi0875 & new_n3388_;
  assign new_n5380_ = pi0166 & ~new_n5379_;
  assign new_n5381_ = ~new_n2447_ & ~new_n3388_;
  assign new_n5382_ = new_n2447_ & ~new_n3386_;
  assign new_n5383_ = pi0875 & ~new_n5382_;
  assign new_n5384_ = ~new_n5381_ & new_n5383_;
  assign new_n5385_ = ~new_n5380_ & ~new_n5384_;
  assign new_n5386_ = ~pi0228 & ~new_n5385_;
  assign new_n5387_ = ~new_n5349_ & ~new_n5386_;
  assign new_n5388_ = ~pi0216 & ~new_n5387_;
  assign new_n5389_ = ~new_n5298_ & ~new_n5388_;
  assign new_n5390_ = ~pi0221 & ~new_n5389_;
  assign new_n5391_ = ~new_n5297_ & ~new_n5390_;
  assign new_n5392_ = ~pi0215 & ~new_n5391_;
  assign new_n5393_ = ~new_n5319_ & ~new_n5392_;
  assign new_n5394_ = pi0299 & ~new_n5393_;
  assign new_n5395_ = new_n3186_ & ~new_n5348_;
  assign new_n5396_ = ~new_n5394_ & new_n5395_;
  assign new_n5397_ = ~new_n3186_ & new_n5375_;
  assign new_n5398_ = pi0100 & ~new_n5397_;
  assign new_n5399_ = ~new_n5396_ & new_n5398_;
  assign new_n5400_ = ~new_n5378_ & ~new_n5399_;
  assign new_n5401_ = ~pi0087 & ~new_n5400_;
  assign new_n5402_ = ~new_n3212_ & new_n5375_;
  assign new_n5403_ = new_n3212_ & new_n5362_;
  assign new_n5404_ = ~new_n5402_ & ~new_n5403_;
  assign new_n5405_ = pi0087 & new_n5404_;
  assign new_n5406_ = ~pi0075 & ~new_n5405_;
  assign new_n5407_ = ~new_n5401_ & new_n5406_;
  assign new_n5408_ = pi0075 & new_n5375_;
  assign new_n5409_ = ~pi0092 & ~new_n5408_;
  assign new_n5410_ = ~new_n5407_ & new_n5409_;
  assign new_n5411_ = new_n3235_ & ~new_n5404_;
  assign new_n5412_ = ~new_n3235_ & new_n5375_;
  assign new_n5413_ = pi0092 & ~new_n5412_;
  assign new_n5414_ = ~new_n5411_ & new_n5413_;
  assign new_n5415_ = new_n3270_ & ~new_n5414_;
  assign new_n5416_ = ~new_n5410_ & new_n5415_;
  assign new_n5417_ = ~new_n3270_ & new_n5375_;
  assign new_n5418_ = ~pi0055 & ~new_n5417_;
  assign new_n5419_ = ~new_n5416_ & new_n5418_;
  assign new_n5420_ = new_n3273_ & new_n5360_;
  assign new_n5421_ = ~new_n3273_ & new_n5373_;
  assign new_n5422_ = pi0055 & ~new_n5421_;
  assign new_n5423_ = ~new_n5420_ & new_n5422_;
  assign new_n5424_ = ~pi0056 & ~new_n5423_;
  assign new_n5425_ = ~new_n5419_ & new_n5424_;
  assign new_n5426_ = new_n3285_ & ~new_n5360_;
  assign new_n5427_ = ~new_n3285_ & ~new_n5373_;
  assign new_n5428_ = pi0056 & ~new_n5427_;
  assign new_n5429_ = ~new_n5426_ & new_n5428_;
  assign new_n5430_ = ~pi0062 & ~new_n5429_;
  assign new_n5431_ = ~new_n5425_ & new_n5430_;
  assign new_n5432_ = new_n3438_ & new_n5360_;
  assign new_n5433_ = ~new_n3438_ & new_n5373_;
  assign new_n5434_ = pi0062 & ~new_n5433_;
  assign new_n5435_ = ~new_n5432_ & new_n5434_;
  assign new_n5436_ = new_n3436_ & ~new_n5435_;
  assign new_n5437_ = ~new_n5431_ & new_n5436_;
  assign new_n5438_ = ~new_n3436_ & new_n5373_;
  assign new_n5439_ = ~pi0245 & ~new_n5438_;
  assign new_n5440_ = ~new_n5437_ & new_n5439_;
  assign new_n5441_ = ~pi0166 & ~new_n3371_;
  assign new_n5442_ = pi0875 & ~new_n5441_;
  assign new_n5443_ = pi0166 & new_n3462_;
  assign new_n5444_ = ~pi0166 & ~new_n3471_;
  assign new_n5445_ = ~pi0875 & ~new_n5444_;
  assign new_n5446_ = ~new_n5443_ & new_n5445_;
  assign new_n5447_ = ~pi0228 & ~new_n5446_;
  assign new_n5448_ = ~new_n5442_ & new_n5447_;
  assign new_n5449_ = new_n5304_ & ~new_n5448_;
  assign new_n5450_ = ~new_n5298_ & ~new_n5449_;
  assign new_n5451_ = ~pi0221 & ~new_n5450_;
  assign new_n5452_ = ~new_n5297_ & ~new_n5451_;
  assign new_n5453_ = ~pi0215 & ~new_n5452_;
  assign new_n5454_ = new_n5320_ & ~new_n5453_;
  assign new_n5455_ = new_n5341_ & ~new_n5454_;
  assign new_n5456_ = ~new_n3481_ & ~new_n5349_;
  assign new_n5457_ = ~new_n5353_ & new_n5456_;
  assign new_n5458_ = ~pi0216 & ~new_n5457_;
  assign new_n5459_ = ~new_n5298_ & ~new_n5458_;
  assign new_n5460_ = ~pi0221 & ~new_n5459_;
  assign new_n5461_ = ~new_n5297_ & ~new_n5460_;
  assign new_n5462_ = ~pi0215 & ~new_n5461_;
  assign new_n5463_ = ~new_n5319_ & ~new_n5462_;
  assign new_n5464_ = pi0299 & ~new_n5463_;
  assign new_n5465_ = ~new_n5346_ & ~new_n5464_;
  assign new_n5466_ = pi0039 & ~new_n5465_;
  assign new_n5467_ = ~pi0038 & ~new_n5466_;
  assign new_n5468_ = ~new_n5455_ & new_n5467_;
  assign new_n5469_ = ~new_n3482_ & new_n5373_;
  assign new_n5470_ = pi0299 & ~new_n5469_;
  assign new_n5471_ = ~new_n5346_ & ~new_n5470_;
  assign new_n5472_ = pi0038 & new_n5471_;
  assign new_n5473_ = ~pi0100 & ~new_n5472_;
  assign new_n5474_ = ~new_n5468_ & new_n5473_;
  assign new_n5475_ = ~new_n5386_ & new_n5456_;
  assign new_n5476_ = ~pi0216 & ~new_n5475_;
  assign new_n5477_ = ~new_n5298_ & ~new_n5476_;
  assign new_n5478_ = ~pi0221 & ~new_n5477_;
  assign new_n5479_ = ~new_n5297_ & ~new_n5478_;
  assign new_n5480_ = ~pi0215 & ~new_n5479_;
  assign new_n5481_ = ~new_n5319_ & ~new_n5480_;
  assign new_n5482_ = pi0299 & ~new_n5481_;
  assign new_n5483_ = new_n3186_ & ~new_n5346_;
  assign new_n5484_ = ~new_n5482_ & new_n5483_;
  assign new_n5485_ = ~new_n3186_ & new_n5471_;
  assign new_n5486_ = pi0100 & ~new_n5485_;
  assign new_n5487_ = ~new_n5484_ & new_n5486_;
  assign new_n5488_ = ~new_n5474_ & ~new_n5487_;
  assign new_n5489_ = ~pi0087 & ~new_n5488_;
  assign new_n5490_ = ~new_n3212_ & new_n5471_;
  assign new_n5491_ = new_n3212_ & new_n5465_;
  assign new_n5492_ = ~new_n5490_ & ~new_n5491_;
  assign new_n5493_ = pi0087 & new_n5492_;
  assign new_n5494_ = ~pi0075 & ~new_n5493_;
  assign new_n5495_ = ~new_n5489_ & new_n5494_;
  assign new_n5496_ = pi0075 & new_n5471_;
  assign new_n5497_ = ~pi0092 & ~new_n5496_;
  assign new_n5498_ = ~new_n5495_ & new_n5497_;
  assign new_n5499_ = new_n3235_ & ~new_n5492_;
  assign new_n5500_ = ~new_n3235_ & new_n5471_;
  assign new_n5501_ = pi0092 & ~new_n5500_;
  assign new_n5502_ = ~new_n5499_ & new_n5501_;
  assign new_n5503_ = new_n3270_ & ~new_n5502_;
  assign new_n5504_ = ~new_n5498_ & new_n5503_;
  assign new_n5505_ = ~new_n3270_ & new_n5471_;
  assign new_n5506_ = ~pi0055 & ~new_n5505_;
  assign new_n5507_ = ~new_n5504_ & new_n5506_;
  assign new_n5508_ = new_n3273_ & new_n5463_;
  assign new_n5509_ = ~new_n3273_ & new_n5469_;
  assign new_n5510_ = pi0055 & ~new_n5509_;
  assign new_n5511_ = ~new_n5508_ & new_n5510_;
  assign new_n5512_ = ~pi0056 & ~new_n5511_;
  assign new_n5513_ = ~new_n5507_ & new_n5512_;
  assign new_n5514_ = new_n3285_ & ~new_n5463_;
  assign new_n5515_ = ~new_n3285_ & ~new_n5469_;
  assign new_n5516_ = pi0056 & ~new_n5515_;
  assign new_n5517_ = ~new_n5514_ & new_n5516_;
  assign new_n5518_ = ~pi0062 & ~new_n5517_;
  assign new_n5519_ = ~new_n5513_ & new_n5518_;
  assign new_n5520_ = new_n3438_ & new_n5463_;
  assign new_n5521_ = ~new_n3438_ & new_n5469_;
  assign new_n5522_ = pi0062 & ~new_n5521_;
  assign new_n5523_ = ~new_n5520_ & new_n5522_;
  assign new_n5524_ = new_n3436_ & ~new_n5523_;
  assign new_n5525_ = ~new_n5519_ & new_n5524_;
  assign new_n5526_ = ~new_n3436_ & new_n5469_;
  assign new_n5527_ = pi0245 & ~new_n5526_;
  assign new_n5528_ = ~new_n5525_ & new_n5527_;
  assign po0163 = new_n5440_ | new_n5528_;
  assign new_n5530_ = ~pi0938 & new_n2437_;
  assign new_n5531_ = ~pi1135 & ~new_n2437_;
  assign new_n5532_ = pi0221 & ~new_n5531_;
  assign new_n5533_ = ~new_n5530_ & new_n5532_;
  assign new_n5534_ = pi0216 & pi0279;
  assign new_n5535_ = pi0879 & ~new_n2449_;
  assign new_n5536_ = pi0105 & ~new_n5535_;
  assign new_n5537_ = ~pi0105 & ~pi0161;
  assign new_n5538_ = ~new_n5536_ & ~new_n5537_;
  assign new_n5539_ = new_n3470_ & ~new_n5538_;
  assign new_n5540_ = ~pi0216 & ~new_n5539_;
  assign new_n5541_ = ~pi0161 & ~new_n3462_;
  assign new_n5542_ = pi0161 & new_n3471_;
  assign new_n5543_ = pi0879 & ~new_n5542_;
  assign new_n5544_ = ~new_n5541_ & new_n5543_;
  assign new_n5545_ = pi0161 & ~pi0879;
  assign new_n5546_ = ~new_n3371_ & new_n5545_;
  assign new_n5547_ = ~new_n5544_ & ~new_n5546_;
  assign new_n5548_ = ~pi0228 & ~new_n5547_;
  assign new_n5549_ = ~new_n3470_ & ~new_n5548_;
  assign new_n5550_ = new_n5540_ & ~new_n5549_;
  assign new_n5551_ = ~new_n5534_ & ~new_n5550_;
  assign new_n5552_ = ~pi0221 & ~new_n5551_;
  assign new_n5553_ = ~new_n5533_ & ~new_n5552_;
  assign new_n5554_ = ~pi0215 & ~new_n5553_;
  assign new_n5555_ = pi0215 & pi1135;
  assign new_n5556_ = pi0299 & ~new_n5555_;
  assign new_n5557_ = ~new_n5554_ & new_n5556_;
  assign new_n5558_ = pi0223 & pi1135;
  assign new_n5559_ = ~pi0299 & ~new_n5558_;
  assign new_n5560_ = ~pi0938 & new_n3045_;
  assign new_n5561_ = ~pi1135 & ~new_n3045_;
  assign new_n5562_ = pi0222 & ~new_n5561_;
  assign new_n5563_ = ~new_n5560_ & new_n5562_;
  assign new_n5564_ = ~pi0224 & ~pi0879;
  assign new_n5565_ = ~new_n2449_ & new_n5564_;
  assign new_n5566_ = pi0224 & ~pi0279;
  assign new_n5567_ = ~pi0222 & ~new_n5566_;
  assign new_n5568_ = ~new_n5565_ & new_n5567_;
  assign new_n5569_ = ~new_n5563_ & ~new_n5568_;
  assign new_n5570_ = ~pi0223 & ~new_n5569_;
  assign new_n5571_ = new_n5327_ & ~new_n5563_;
  assign new_n5572_ = new_n5570_ & ~new_n5571_;
  assign new_n5573_ = new_n5559_ & ~new_n5572_;
  assign new_n5574_ = ~pi0039 & ~new_n5573_;
  assign new_n5575_ = ~new_n5557_ & new_n5574_;
  assign new_n5576_ = ~new_n5558_ & ~new_n5570_;
  assign new_n5577_ = ~pi0299 & ~new_n5576_;
  assign new_n5578_ = new_n3105_ & ~new_n5535_;
  assign new_n5579_ = new_n5577_ & ~new_n5578_;
  assign new_n5580_ = pi0228 & new_n5538_;
  assign new_n5581_ = ~pi0879 & new_n3100_;
  assign new_n5582_ = pi0161 & ~pi0228;
  assign new_n5583_ = ~new_n3326_ & ~new_n5582_;
  assign new_n5584_ = ~new_n5581_ & ~new_n5583_;
  assign new_n5585_ = ~new_n5580_ & ~new_n5584_;
  assign new_n5586_ = ~pi0216 & ~new_n5585_;
  assign new_n5587_ = ~new_n5534_ & ~new_n5586_;
  assign new_n5588_ = ~pi0221 & ~new_n5587_;
  assign new_n5589_ = ~new_n5533_ & ~new_n5588_;
  assign new_n5590_ = ~pi0215 & ~new_n5589_;
  assign new_n5591_ = ~new_n5555_ & ~new_n5590_;
  assign new_n5592_ = pi0299 & ~new_n5591_;
  assign new_n5593_ = ~new_n5579_ & ~new_n5592_;
  assign new_n5594_ = pi0039 & ~new_n5593_;
  assign new_n5595_ = ~pi0038 & ~new_n5594_;
  assign new_n5596_ = ~new_n5575_ & new_n5595_;
  assign new_n5597_ = ~new_n5580_ & ~new_n5582_;
  assign new_n5598_ = ~pi0216 & ~new_n5597_;
  assign new_n5599_ = ~new_n5534_ & ~new_n5598_;
  assign new_n5600_ = ~pi0221 & ~new_n5599_;
  assign new_n5601_ = ~new_n5533_ & ~new_n5600_;
  assign new_n5602_ = ~pi0215 & ~new_n5601_;
  assign new_n5603_ = ~new_n5555_ & ~new_n5602_;
  assign new_n5604_ = pi0299 & ~new_n5603_;
  assign new_n5605_ = ~new_n5579_ & ~new_n5604_;
  assign new_n5606_ = pi0038 & new_n5605_;
  assign new_n5607_ = ~pi0100 & ~new_n5606_;
  assign new_n5608_ = ~new_n5596_ & new_n5607_;
  assign new_n5609_ = ~pi0879 & new_n3388_;
  assign new_n5610_ = pi0161 & ~new_n5609_;
  assign new_n5611_ = ~pi0152 & ~pi0166;
  assign new_n5612_ = ~new_n3388_ & ~new_n5611_;
  assign new_n5613_ = ~new_n3386_ & new_n5611_;
  assign new_n5614_ = pi0879 & ~new_n5613_;
  assign new_n5615_ = ~new_n5612_ & new_n5614_;
  assign new_n5616_ = ~new_n5610_ & ~new_n5615_;
  assign new_n5617_ = ~pi0228 & ~new_n5616_;
  assign new_n5618_ = ~new_n5580_ & ~new_n5617_;
  assign new_n5619_ = ~pi0216 & ~new_n5618_;
  assign new_n5620_ = ~new_n5534_ & ~new_n5619_;
  assign new_n5621_ = ~pi0221 & ~new_n5620_;
  assign new_n5622_ = ~new_n5533_ & ~new_n5621_;
  assign new_n5623_ = ~pi0215 & ~new_n5622_;
  assign new_n5624_ = ~new_n5555_ & ~new_n5623_;
  assign new_n5625_ = pi0299 & ~new_n5624_;
  assign new_n5626_ = new_n3186_ & ~new_n5579_;
  assign new_n5627_ = ~new_n5625_ & new_n5626_;
  assign new_n5628_ = ~new_n3186_ & new_n5605_;
  assign new_n5629_ = pi0100 & ~new_n5628_;
  assign new_n5630_ = ~new_n5627_ & new_n5629_;
  assign new_n5631_ = ~new_n5608_ & ~new_n5630_;
  assign new_n5632_ = ~pi0087 & ~new_n5631_;
  assign new_n5633_ = ~new_n3212_ & new_n5605_;
  assign new_n5634_ = new_n3212_ & new_n5593_;
  assign new_n5635_ = ~new_n5633_ & ~new_n5634_;
  assign new_n5636_ = pi0087 & new_n5635_;
  assign new_n5637_ = ~pi0075 & ~new_n5636_;
  assign new_n5638_ = ~new_n5632_ & new_n5637_;
  assign new_n5639_ = pi0075 & new_n5605_;
  assign new_n5640_ = ~pi0092 & ~new_n5639_;
  assign new_n5641_ = ~new_n5638_ & new_n5640_;
  assign new_n5642_ = new_n3235_ & ~new_n5635_;
  assign new_n5643_ = ~new_n3235_ & new_n5605_;
  assign new_n5644_ = pi0092 & ~new_n5643_;
  assign new_n5645_ = ~new_n5642_ & new_n5644_;
  assign new_n5646_ = new_n3270_ & ~new_n5645_;
  assign new_n5647_ = ~new_n5641_ & new_n5646_;
  assign new_n5648_ = ~new_n3270_ & new_n5605_;
  assign new_n5649_ = ~pi0055 & ~new_n5648_;
  assign new_n5650_ = ~new_n5647_ & new_n5649_;
  assign new_n5651_ = new_n3273_ & new_n5591_;
  assign new_n5652_ = ~new_n3273_ & new_n5603_;
  assign new_n5653_ = pi0055 & ~new_n5652_;
  assign new_n5654_ = ~new_n5651_ & new_n5653_;
  assign new_n5655_ = ~pi0056 & ~new_n5654_;
  assign new_n5656_ = ~new_n5650_ & new_n5655_;
  assign new_n5657_ = new_n3285_ & ~new_n5591_;
  assign new_n5658_ = ~new_n3285_ & ~new_n5603_;
  assign new_n5659_ = pi0056 & ~new_n5658_;
  assign new_n5660_ = ~new_n5657_ & new_n5659_;
  assign new_n5661_ = ~pi0062 & ~new_n5660_;
  assign new_n5662_ = ~new_n5656_ & new_n5661_;
  assign new_n5663_ = new_n3438_ & new_n5591_;
  assign new_n5664_ = ~new_n3438_ & new_n5603_;
  assign new_n5665_ = pi0062 & ~new_n5664_;
  assign new_n5666_ = ~new_n5663_ & new_n5665_;
  assign new_n5667_ = new_n3436_ & ~new_n5666_;
  assign new_n5668_ = ~new_n5662_ & new_n5667_;
  assign new_n5669_ = ~new_n3436_ & new_n5603_;
  assign new_n5670_ = ~pi0244 & ~new_n5669_;
  assign new_n5671_ = ~new_n5668_ & new_n5670_;
  assign new_n5672_ = ~pi0161 & ~new_n3371_;
  assign new_n5673_ = pi0879 & ~new_n5672_;
  assign new_n5674_ = pi0161 & new_n3462_;
  assign new_n5675_ = ~pi0161 & ~new_n3471_;
  assign new_n5676_ = ~pi0879 & ~new_n5675_;
  assign new_n5677_ = ~new_n5674_ & new_n5676_;
  assign new_n5678_ = ~pi0228 & ~new_n5677_;
  assign new_n5679_ = ~new_n5673_ & new_n5678_;
  assign new_n5680_ = new_n5540_ & ~new_n5679_;
  assign new_n5681_ = ~new_n5534_ & ~new_n5680_;
  assign new_n5682_ = ~pi0221 & ~new_n5681_;
  assign new_n5683_ = ~new_n5533_ & ~new_n5682_;
  assign new_n5684_ = ~pi0215 & ~new_n5683_;
  assign new_n5685_ = new_n5556_ & ~new_n5684_;
  assign new_n5686_ = ~new_n5327_ & new_n5569_;
  assign new_n5687_ = ~pi0223 & ~new_n5686_;
  assign new_n5688_ = new_n5559_ & ~new_n5687_;
  assign new_n5689_ = ~pi0039 & ~new_n5688_;
  assign new_n5690_ = ~new_n5685_ & new_n5689_;
  assign new_n5691_ = ~new_n3481_ & ~new_n5580_;
  assign new_n5692_ = ~new_n5584_ & new_n5691_;
  assign new_n5693_ = ~pi0216 & ~new_n5692_;
  assign new_n5694_ = ~new_n5534_ & ~new_n5693_;
  assign new_n5695_ = ~pi0221 & ~new_n5694_;
  assign new_n5696_ = ~new_n5533_ & ~new_n5695_;
  assign new_n5697_ = ~pi0215 & ~new_n5696_;
  assign new_n5698_ = ~new_n5555_ & ~new_n5697_;
  assign new_n5699_ = pi0299 & ~new_n5698_;
  assign new_n5700_ = ~new_n5577_ & ~new_n5699_;
  assign new_n5701_ = pi0039 & ~new_n5700_;
  assign new_n5702_ = ~pi0038 & ~new_n5701_;
  assign new_n5703_ = ~new_n5690_ & new_n5702_;
  assign new_n5704_ = ~new_n3482_ & new_n5603_;
  assign new_n5705_ = pi0299 & ~new_n5704_;
  assign new_n5706_ = ~new_n5577_ & ~new_n5705_;
  assign new_n5707_ = pi0038 & new_n5706_;
  assign new_n5708_ = ~pi0100 & ~new_n5707_;
  assign new_n5709_ = ~new_n5703_ & new_n5708_;
  assign new_n5710_ = ~new_n5617_ & new_n5691_;
  assign new_n5711_ = ~pi0216 & ~new_n5710_;
  assign new_n5712_ = ~new_n5534_ & ~new_n5711_;
  assign new_n5713_ = ~pi0221 & ~new_n5712_;
  assign new_n5714_ = ~new_n5533_ & ~new_n5713_;
  assign new_n5715_ = ~pi0215 & ~new_n5714_;
  assign new_n5716_ = ~new_n5555_ & ~new_n5715_;
  assign new_n5717_ = pi0299 & ~new_n5716_;
  assign new_n5718_ = new_n3186_ & ~new_n5577_;
  assign new_n5719_ = ~new_n5717_ & new_n5718_;
  assign new_n5720_ = ~new_n3186_ & new_n5706_;
  assign new_n5721_ = pi0100 & ~new_n5720_;
  assign new_n5722_ = ~new_n5719_ & new_n5721_;
  assign new_n5723_ = ~new_n5709_ & ~new_n5722_;
  assign new_n5724_ = ~pi0087 & ~new_n5723_;
  assign new_n5725_ = ~new_n3212_ & new_n5706_;
  assign new_n5726_ = new_n3212_ & new_n5700_;
  assign new_n5727_ = ~new_n5725_ & ~new_n5726_;
  assign new_n5728_ = pi0087 & new_n5727_;
  assign new_n5729_ = ~pi0075 & ~new_n5728_;
  assign new_n5730_ = ~new_n5724_ & new_n5729_;
  assign new_n5731_ = pi0075 & new_n5706_;
  assign new_n5732_ = ~pi0092 & ~new_n5731_;
  assign new_n5733_ = ~new_n5730_ & new_n5732_;
  assign new_n5734_ = new_n3235_ & ~new_n5727_;
  assign new_n5735_ = ~new_n3235_ & new_n5706_;
  assign new_n5736_ = pi0092 & ~new_n5735_;
  assign new_n5737_ = ~new_n5734_ & new_n5736_;
  assign new_n5738_ = new_n3270_ & ~new_n5737_;
  assign new_n5739_ = ~new_n5733_ & new_n5738_;
  assign new_n5740_ = ~new_n3270_ & new_n5706_;
  assign new_n5741_ = ~pi0055 & ~new_n5740_;
  assign new_n5742_ = ~new_n5739_ & new_n5741_;
  assign new_n5743_ = new_n3273_ & new_n5698_;
  assign new_n5744_ = ~new_n3273_ & new_n5704_;
  assign new_n5745_ = pi0055 & ~new_n5744_;
  assign new_n5746_ = ~new_n5743_ & new_n5745_;
  assign new_n5747_ = ~pi0056 & ~new_n5746_;
  assign new_n5748_ = ~new_n5742_ & new_n5747_;
  assign new_n5749_ = new_n3285_ & ~new_n5698_;
  assign new_n5750_ = ~new_n3285_ & ~new_n5704_;
  assign new_n5751_ = pi0056 & ~new_n5750_;
  assign new_n5752_ = ~new_n5749_ & new_n5751_;
  assign new_n5753_ = ~pi0062 & ~new_n5752_;
  assign new_n5754_ = ~new_n5748_ & new_n5753_;
  assign new_n5755_ = new_n3438_ & new_n5698_;
  assign new_n5756_ = ~new_n3438_ & new_n5704_;
  assign new_n5757_ = pi0062 & ~new_n5756_;
  assign new_n5758_ = ~new_n5755_ & new_n5757_;
  assign new_n5759_ = new_n3436_ & ~new_n5758_;
  assign new_n5760_ = ~new_n5754_ & new_n5759_;
  assign new_n5761_ = ~new_n3436_ & new_n5704_;
  assign new_n5762_ = pi0244 & ~new_n5761_;
  assign new_n5763_ = ~new_n5760_ & new_n5762_;
  assign po0164 = new_n5671_ | new_n5763_;
  assign new_n5765_ = pi0833 & ~pi0930;
  assign new_n5766_ = ~pi0216 & pi0221;
  assign new_n5767_ = new_n5765_ & new_n5766_;
  assign new_n5768_ = pi0216 & pi0278;
  assign new_n5769_ = ~pi0221 & ~new_n5768_;
  assign new_n5770_ = ~pi0105 & pi0152;
  assign new_n5771_ = pi0228 & ~new_n5770_;
  assign new_n5772_ = ~pi0846 & new_n3448_;
  assign new_n5773_ = pi0105 & ~new_n5772_;
  assign new_n5774_ = new_n5771_ & ~new_n5773_;
  assign new_n5775_ = ~pi0216 & ~new_n5774_;
  assign new_n5776_ = pi0152 & ~new_n3462_;
  assign new_n5777_ = ~pi0152 & new_n3471_;
  assign new_n5778_ = ~pi0846 & ~new_n5777_;
  assign new_n5779_ = ~new_n5776_ & new_n5778_;
  assign new_n5780_ = ~pi0152 & pi0846;
  assign new_n5781_ = ~new_n3371_ & new_n5780_;
  assign new_n5782_ = ~new_n5779_ & ~new_n5781_;
  assign new_n5783_ = ~pi0228 & ~new_n5782_;
  assign new_n5784_ = new_n5775_ & ~new_n5783_;
  assign new_n5785_ = new_n5769_ & ~new_n5784_;
  assign new_n5786_ = ~new_n5767_ & ~new_n5785_;
  assign new_n5787_ = pi0221 & ~new_n2437_;
  assign new_n5788_ = ~pi0215 & pi0299;
  assign new_n5789_ = ~new_n5787_ & new_n5788_;
  assign new_n5790_ = new_n5786_ & new_n5789_;
  assign new_n5791_ = pi0222 & ~pi0224;
  assign new_n5792_ = new_n5765_ & new_n5791_;
  assign new_n5793_ = pi0224 & pi0278;
  assign new_n5794_ = ~pi0222 & ~new_n5793_;
  assign new_n5795_ = ~pi0224 & ~new_n5772_;
  assign new_n5796_ = new_n5794_ & ~new_n5795_;
  assign new_n5797_ = ~new_n5792_ & ~new_n5796_;
  assign new_n5798_ = ~new_n3046_ & new_n3489_;
  assign new_n5799_ = new_n5797_ & new_n5798_;
  assign new_n5800_ = ~pi0039 & ~new_n5799_;
  assign new_n5801_ = ~new_n5790_ & new_n5800_;
  assign new_n5802_ = pi0846 & ~new_n2449_;
  assign new_n5803_ = ~pi0224 & new_n5802_;
  assign new_n5804_ = new_n5794_ & ~new_n5803_;
  assign new_n5805_ = new_n3047_ & ~new_n5792_;
  assign new_n5806_ = ~new_n5804_ & new_n5805_;
  assign new_n5807_ = ~pi0299 & ~new_n5806_;
  assign new_n5808_ = ~new_n3870_ & new_n5807_;
  assign new_n5809_ = ~pi0215 & ~new_n5787_;
  assign new_n5810_ = ~new_n5767_ & new_n5809_;
  assign new_n5811_ = pi0105 & new_n5802_;
  assign new_n5812_ = ~new_n5770_ & ~new_n5811_;
  assign new_n5813_ = pi0228 & ~new_n5812_;
  assign new_n5814_ = ~new_n3481_ & ~new_n5813_;
  assign new_n5815_ = ~pi0846 & new_n3100_;
  assign new_n5816_ = ~pi0152 & ~new_n3100_;
  assign new_n5817_ = ~pi0228 & ~new_n5816_;
  assign new_n5818_ = ~new_n5815_ & new_n5817_;
  assign new_n5819_ = new_n5814_ & ~new_n5818_;
  assign new_n5820_ = ~pi0216 & ~new_n5819_;
  assign new_n5821_ = new_n5769_ & ~new_n5820_;
  assign new_n5822_ = new_n5810_ & ~new_n5821_;
  assign new_n5823_ = pi0299 & ~new_n5822_;
  assign new_n5824_ = ~new_n5808_ & ~new_n5823_;
  assign new_n5825_ = pi0039 & ~new_n5824_;
  assign new_n5826_ = ~pi0038 & ~new_n5825_;
  assign new_n5827_ = ~new_n5801_ & new_n5826_;
  assign new_n5828_ = pi0152 & ~pi0228;
  assign new_n5829_ = ~new_n5813_ & ~new_n5828_;
  assign new_n5830_ = ~pi0216 & ~new_n5829_;
  assign new_n5831_ = new_n5769_ & ~new_n5830_;
  assign new_n5832_ = new_n5810_ & ~new_n5831_;
  assign new_n5833_ = ~new_n3482_ & ~new_n5832_;
  assign new_n5834_ = pi0299 & new_n5833_;
  assign new_n5835_ = ~new_n5808_ & ~new_n5834_;
  assign new_n5836_ = pi0038 & new_n5835_;
  assign new_n5837_ = ~pi0100 & ~new_n5836_;
  assign new_n5838_ = ~new_n5827_ & new_n5837_;
  assign new_n5839_ = pi0846 & ~new_n3394_;
  assign new_n5840_ = ~new_n3389_ & ~new_n5839_;
  assign new_n5841_ = ~pi0228 & ~new_n5840_;
  assign new_n5842_ = new_n5814_ & ~new_n5841_;
  assign new_n5843_ = ~pi0216 & ~new_n5842_;
  assign new_n5844_ = new_n5769_ & ~new_n5843_;
  assign new_n5845_ = new_n5810_ & ~new_n5844_;
  assign new_n5846_ = pi0299 & ~new_n5845_;
  assign new_n5847_ = new_n3186_ & ~new_n5808_;
  assign new_n5848_ = ~new_n5846_ & new_n5847_;
  assign new_n5849_ = ~new_n3186_ & new_n5835_;
  assign new_n5850_ = pi0100 & ~new_n5849_;
  assign new_n5851_ = ~new_n5848_ & new_n5850_;
  assign new_n5852_ = ~new_n5838_ & ~new_n5851_;
  assign new_n5853_ = ~pi0087 & ~new_n5852_;
  assign new_n5854_ = ~new_n3212_ & new_n5835_;
  assign new_n5855_ = new_n3212_ & new_n5824_;
  assign new_n5856_ = ~new_n5854_ & ~new_n5855_;
  assign new_n5857_ = pi0087 & new_n5856_;
  assign new_n5858_ = ~pi0075 & ~new_n5857_;
  assign new_n5859_ = ~new_n5853_ & new_n5858_;
  assign new_n5860_ = pi0075 & new_n5835_;
  assign new_n5861_ = ~pi0092 & ~new_n5860_;
  assign new_n5862_ = ~new_n5859_ & new_n5861_;
  assign new_n5863_ = new_n3235_ & ~new_n5856_;
  assign new_n5864_ = ~new_n3235_ & new_n5835_;
  assign new_n5865_ = pi0092 & ~new_n5864_;
  assign new_n5866_ = ~new_n5863_ & new_n5865_;
  assign new_n5867_ = new_n3270_ & ~new_n5866_;
  assign new_n5868_ = ~new_n5862_ & new_n5867_;
  assign new_n5869_ = ~new_n3270_ & new_n5835_;
  assign new_n5870_ = ~pi0055 & ~new_n5869_;
  assign new_n5871_ = ~new_n5868_ & new_n5870_;
  assign new_n5872_ = new_n3273_ & new_n5822_;
  assign new_n5873_ = ~new_n3273_ & ~new_n5833_;
  assign new_n5874_ = pi0055 & ~new_n5873_;
  assign new_n5875_ = ~new_n5872_ & new_n5874_;
  assign new_n5876_ = ~pi0056 & ~new_n5875_;
  assign new_n5877_ = ~new_n5871_ & new_n5876_;
  assign new_n5878_ = new_n3285_ & ~new_n5822_;
  assign new_n5879_ = ~new_n3285_ & new_n5833_;
  assign new_n5880_ = pi0056 & ~new_n5879_;
  assign new_n5881_ = ~new_n5878_ & new_n5880_;
  assign new_n5882_ = ~pi0062 & ~new_n5881_;
  assign new_n5883_ = ~new_n5877_ & new_n5882_;
  assign new_n5884_ = new_n3438_ & new_n5822_;
  assign new_n5885_ = ~new_n3438_ & ~new_n5833_;
  assign new_n5886_ = pi0062 & ~new_n5885_;
  assign new_n5887_ = ~new_n5884_ & new_n5886_;
  assign new_n5888_ = new_n3436_ & ~new_n5887_;
  assign new_n5889_ = ~new_n5883_ & new_n5888_;
  assign new_n5890_ = ~new_n3436_ & ~new_n5833_;
  assign new_n5891_ = pi0242 & ~new_n5890_;
  assign new_n5892_ = ~new_n5889_ & new_n5891_;
  assign new_n5893_ = ~pi0152 & ~new_n3462_;
  assign new_n5894_ = pi0152 & new_n3471_;
  assign new_n5895_ = pi0846 & ~new_n5894_;
  assign new_n5896_ = ~new_n5893_ & new_n5895_;
  assign new_n5897_ = pi0152 & ~pi0846;
  assign new_n5898_ = ~new_n3371_ & new_n5897_;
  assign new_n5899_ = ~pi0228 & ~new_n5898_;
  assign new_n5900_ = ~new_n5896_ & new_n5899_;
  assign new_n5901_ = ~new_n3448_ & new_n5771_;
  assign new_n5902_ = new_n5775_ & ~new_n5901_;
  assign new_n5903_ = ~new_n5900_ & new_n5902_;
  assign new_n5904_ = new_n5769_ & ~new_n5903_;
  assign new_n5905_ = ~new_n5767_ & ~new_n5904_;
  assign new_n5906_ = new_n5789_ & new_n5905_;
  assign new_n5907_ = ~new_n3447_ & new_n5803_;
  assign new_n5908_ = new_n5794_ & ~new_n5907_;
  assign new_n5909_ = ~new_n5792_ & new_n5798_;
  assign new_n5910_ = ~new_n5908_ & new_n5909_;
  assign new_n5911_ = ~pi0039 & ~new_n5910_;
  assign new_n5912_ = ~new_n5906_ & new_n5911_;
  assign new_n5913_ = ~new_n5813_ & ~new_n5818_;
  assign new_n5914_ = ~pi0216 & ~new_n5913_;
  assign new_n5915_ = new_n5769_ & ~new_n5914_;
  assign new_n5916_ = new_n5810_ & ~new_n5915_;
  assign new_n5917_ = pi0299 & ~new_n5916_;
  assign new_n5918_ = ~new_n5807_ & ~new_n5917_;
  assign new_n5919_ = pi0039 & ~new_n5918_;
  assign new_n5920_ = ~pi0038 & ~new_n5919_;
  assign new_n5921_ = ~new_n5912_ & new_n5920_;
  assign new_n5922_ = pi0299 & ~new_n5832_;
  assign new_n5923_ = ~new_n5807_ & ~new_n5922_;
  assign new_n5924_ = pi0038 & new_n5923_;
  assign new_n5925_ = ~pi0100 & ~new_n5924_;
  assign new_n5926_ = ~new_n5921_ & new_n5925_;
  assign new_n5927_ = ~new_n5813_ & ~new_n5841_;
  assign new_n5928_ = ~pi0216 & ~new_n5927_;
  assign new_n5929_ = new_n5769_ & ~new_n5928_;
  assign new_n5930_ = new_n5810_ & ~new_n5929_;
  assign new_n5931_ = pi0299 & ~new_n5930_;
  assign new_n5932_ = new_n3186_ & ~new_n5807_;
  assign new_n5933_ = ~new_n5931_ & new_n5932_;
  assign new_n5934_ = ~new_n3186_ & new_n5923_;
  assign new_n5935_ = pi0100 & ~new_n5934_;
  assign new_n5936_ = ~new_n5933_ & new_n5935_;
  assign new_n5937_ = ~new_n5926_ & ~new_n5936_;
  assign new_n5938_ = ~pi0087 & ~new_n5937_;
  assign new_n5939_ = ~new_n3212_ & new_n5923_;
  assign new_n5940_ = new_n3212_ & new_n5918_;
  assign new_n5941_ = ~new_n5939_ & ~new_n5940_;
  assign new_n5942_ = pi0087 & new_n5941_;
  assign new_n5943_ = ~pi0075 & ~new_n5942_;
  assign new_n5944_ = ~new_n5938_ & new_n5943_;
  assign new_n5945_ = pi0075 & new_n5923_;
  assign new_n5946_ = ~pi0092 & ~new_n5945_;
  assign new_n5947_ = ~new_n5944_ & new_n5946_;
  assign new_n5948_ = new_n3235_ & ~new_n5941_;
  assign new_n5949_ = ~new_n3235_ & new_n5923_;
  assign new_n5950_ = pi0092 & ~new_n5949_;
  assign new_n5951_ = ~new_n5948_ & new_n5950_;
  assign new_n5952_ = new_n3270_ & ~new_n5951_;
  assign new_n5953_ = ~new_n5947_ & new_n5952_;
  assign new_n5954_ = ~new_n3270_ & new_n5923_;
  assign new_n5955_ = ~pi0055 & ~new_n5954_;
  assign new_n5956_ = ~new_n5953_ & new_n5955_;
  assign new_n5957_ = new_n3273_ & new_n5916_;
  assign new_n5958_ = ~new_n3273_ & new_n5832_;
  assign new_n5959_ = pi0055 & ~new_n5958_;
  assign new_n5960_ = ~new_n5957_ & new_n5959_;
  assign new_n5961_ = ~pi0056 & ~new_n5960_;
  assign new_n5962_ = ~new_n5956_ & new_n5961_;
  assign new_n5963_ = new_n3285_ & ~new_n5916_;
  assign new_n5964_ = ~new_n3285_ & ~new_n5832_;
  assign new_n5965_ = pi0056 & ~new_n5964_;
  assign new_n5966_ = ~new_n5963_ & new_n5965_;
  assign new_n5967_ = ~pi0062 & ~new_n5966_;
  assign new_n5968_ = ~new_n5962_ & new_n5967_;
  assign new_n5969_ = new_n3438_ & new_n5916_;
  assign new_n5970_ = ~new_n3438_ & new_n5832_;
  assign new_n5971_ = pi0062 & ~new_n5970_;
  assign new_n5972_ = ~new_n5969_ & new_n5971_;
  assign new_n5973_ = new_n3436_ & ~new_n5972_;
  assign new_n5974_ = ~new_n5968_ & new_n5973_;
  assign new_n5975_ = ~new_n3436_ & new_n5832_;
  assign new_n5976_ = ~pi0242 & ~new_n5975_;
  assign new_n5977_ = ~new_n5974_ & new_n5976_;
  assign new_n5978_ = ~new_n5892_ & ~new_n5977_;
  assign new_n5979_ = ~pi1134 & ~new_n5978_;
  assign new_n5980_ = new_n3489_ & ~new_n5797_;
  assign new_n5981_ = ~pi0039 & ~new_n5980_;
  assign new_n5982_ = ~new_n5786_ & new_n5788_;
  assign new_n5983_ = new_n5981_ & ~new_n5982_;
  assign new_n5984_ = new_n3047_ & new_n5808_;
  assign new_n5985_ = ~pi0299 & ~new_n5984_;
  assign new_n5986_ = ~new_n5767_ & ~new_n5821_;
  assign new_n5987_ = ~pi0215 & ~new_n5986_;
  assign new_n5988_ = pi0299 & ~new_n5987_;
  assign new_n5989_ = ~new_n5985_ & ~new_n5988_;
  assign new_n5990_ = pi0039 & ~new_n5989_;
  assign new_n5991_ = ~pi0038 & ~new_n5990_;
  assign new_n5992_ = ~new_n5983_ & new_n5991_;
  assign new_n5993_ = ~new_n5767_ & ~new_n5831_;
  assign new_n5994_ = ~pi0215 & ~new_n5993_;
  assign new_n5995_ = ~new_n3482_ & new_n5994_;
  assign new_n5996_ = pi0299 & ~new_n5995_;
  assign new_n5997_ = ~new_n5985_ & ~new_n5996_;
  assign new_n5998_ = pi0038 & new_n5997_;
  assign new_n5999_ = ~pi0100 & ~new_n5998_;
  assign new_n6000_ = ~new_n5992_ & new_n5999_;
  assign new_n6001_ = ~new_n5767_ & ~new_n5844_;
  assign new_n6002_ = ~pi0215 & ~new_n6001_;
  assign new_n6003_ = pi0299 & ~new_n6002_;
  assign new_n6004_ = new_n3186_ & ~new_n5985_;
  assign new_n6005_ = ~new_n6003_ & new_n6004_;
  assign new_n6006_ = ~new_n3186_ & new_n5997_;
  assign new_n6007_ = pi0100 & ~new_n6006_;
  assign new_n6008_ = ~new_n6005_ & new_n6007_;
  assign new_n6009_ = ~new_n6000_ & ~new_n6008_;
  assign new_n6010_ = ~pi0087 & ~new_n6009_;
  assign new_n6011_ = ~new_n3212_ & new_n5997_;
  assign new_n6012_ = new_n3212_ & new_n5989_;
  assign new_n6013_ = ~new_n6011_ & ~new_n6012_;
  assign new_n6014_ = pi0087 & new_n6013_;
  assign new_n6015_ = ~pi0075 & ~new_n6014_;
  assign new_n6016_ = ~new_n6010_ & new_n6015_;
  assign new_n6017_ = pi0075 & new_n5997_;
  assign new_n6018_ = ~pi0092 & ~new_n6017_;
  assign new_n6019_ = ~new_n6016_ & new_n6018_;
  assign new_n6020_ = new_n3235_ & ~new_n6013_;
  assign new_n6021_ = ~new_n3235_ & new_n5997_;
  assign new_n6022_ = pi0092 & ~new_n6021_;
  assign new_n6023_ = ~new_n6020_ & new_n6022_;
  assign new_n6024_ = new_n3270_ & ~new_n6023_;
  assign new_n6025_ = ~new_n6019_ & new_n6024_;
  assign new_n6026_ = ~new_n3270_ & new_n5997_;
  assign new_n6027_ = ~pi0055 & ~new_n6026_;
  assign new_n6028_ = ~new_n6025_ & new_n6027_;
  assign new_n6029_ = new_n3273_ & new_n5987_;
  assign new_n6030_ = ~new_n3273_ & new_n5995_;
  assign new_n6031_ = pi0055 & ~new_n6030_;
  assign new_n6032_ = ~new_n6029_ & new_n6031_;
  assign new_n6033_ = ~pi0056 & ~new_n6032_;
  assign new_n6034_ = ~new_n6028_ & new_n6033_;
  assign new_n6035_ = new_n3285_ & ~new_n5987_;
  assign new_n6036_ = ~new_n3285_ & ~new_n5995_;
  assign new_n6037_ = pi0056 & ~new_n6036_;
  assign new_n6038_ = ~new_n6035_ & new_n6037_;
  assign new_n6039_ = ~pi0062 & ~new_n6038_;
  assign new_n6040_ = ~new_n6034_ & new_n6039_;
  assign new_n6041_ = new_n3438_ & new_n5987_;
  assign new_n6042_ = ~new_n3438_ & new_n5995_;
  assign new_n6043_ = pi0062 & ~new_n6042_;
  assign new_n6044_ = ~new_n6041_ & new_n6043_;
  assign new_n6045_ = new_n3436_ & ~new_n6044_;
  assign new_n6046_ = ~new_n6040_ & new_n6045_;
  assign new_n6047_ = ~new_n3436_ & new_n5995_;
  assign new_n6048_ = pi0242 & ~new_n6047_;
  assign new_n6049_ = ~new_n6046_ & new_n6048_;
  assign new_n6050_ = new_n5788_ & ~new_n5905_;
  assign new_n6051_ = new_n3489_ & new_n5908_;
  assign new_n6052_ = new_n5981_ & ~new_n6051_;
  assign new_n6053_ = ~new_n6050_ & new_n6052_;
  assign new_n6054_ = ~pi0223 & new_n5804_;
  assign new_n6055_ = new_n5985_ & ~new_n6054_;
  assign new_n6056_ = ~new_n5767_ & ~new_n5915_;
  assign new_n6057_ = ~pi0215 & ~new_n6056_;
  assign new_n6058_ = pi0299 & ~new_n6057_;
  assign new_n6059_ = ~new_n6055_ & ~new_n6058_;
  assign new_n6060_ = pi0039 & ~new_n6059_;
  assign new_n6061_ = ~pi0038 & ~new_n6060_;
  assign new_n6062_ = ~new_n6053_ & new_n6061_;
  assign new_n6063_ = pi0299 & ~new_n5994_;
  assign new_n6064_ = ~new_n6055_ & ~new_n6063_;
  assign new_n6065_ = pi0038 & new_n6064_;
  assign new_n6066_ = ~pi0100 & ~new_n6065_;
  assign new_n6067_ = ~new_n6062_ & new_n6066_;
  assign new_n6068_ = ~new_n5767_ & ~new_n5929_;
  assign new_n6069_ = ~pi0215 & ~new_n6068_;
  assign new_n6070_ = pi0299 & ~new_n6069_;
  assign new_n6071_ = new_n3186_ & ~new_n6055_;
  assign new_n6072_ = ~new_n6070_ & new_n6071_;
  assign new_n6073_ = ~new_n3186_ & new_n6064_;
  assign new_n6074_ = pi0100 & ~new_n6073_;
  assign new_n6075_ = ~new_n6072_ & new_n6074_;
  assign new_n6076_ = ~new_n6067_ & ~new_n6075_;
  assign new_n6077_ = ~pi0087 & ~new_n6076_;
  assign new_n6078_ = ~new_n3212_ & new_n6064_;
  assign new_n6079_ = new_n3212_ & new_n6059_;
  assign new_n6080_ = ~new_n6078_ & ~new_n6079_;
  assign new_n6081_ = pi0087 & new_n6080_;
  assign new_n6082_ = ~pi0075 & ~new_n6081_;
  assign new_n6083_ = ~new_n6077_ & new_n6082_;
  assign new_n6084_ = pi0075 & new_n6064_;
  assign new_n6085_ = ~pi0092 & ~new_n6084_;
  assign new_n6086_ = ~new_n6083_ & new_n6085_;
  assign new_n6087_ = new_n3235_ & ~new_n6080_;
  assign new_n6088_ = ~new_n3235_ & new_n6064_;
  assign new_n6089_ = pi0092 & ~new_n6088_;
  assign new_n6090_ = ~new_n6087_ & new_n6089_;
  assign new_n6091_ = new_n3270_ & ~new_n6090_;
  assign new_n6092_ = ~new_n6086_ & new_n6091_;
  assign new_n6093_ = ~new_n3270_ & new_n6064_;
  assign new_n6094_ = ~pi0055 & ~new_n6093_;
  assign new_n6095_ = ~new_n6092_ & new_n6094_;
  assign new_n6096_ = new_n3273_ & new_n6057_;
  assign new_n6097_ = ~new_n3273_ & new_n5994_;
  assign new_n6098_ = pi0055 & ~new_n6097_;
  assign new_n6099_ = ~new_n6096_ & new_n6098_;
  assign new_n6100_ = ~pi0056 & ~new_n6099_;
  assign new_n6101_ = ~new_n6095_ & new_n6100_;
  assign new_n6102_ = new_n3285_ & ~new_n6057_;
  assign new_n6103_ = ~new_n3285_ & ~new_n5994_;
  assign new_n6104_ = pi0056 & ~new_n6103_;
  assign new_n6105_ = ~new_n6102_ & new_n6104_;
  assign new_n6106_ = ~pi0062 & ~new_n6105_;
  assign new_n6107_ = ~new_n6101_ & new_n6106_;
  assign new_n6108_ = new_n3438_ & new_n6057_;
  assign new_n6109_ = ~new_n3438_ & new_n5994_;
  assign new_n6110_ = pi0062 & ~new_n6109_;
  assign new_n6111_ = ~new_n6108_ & new_n6110_;
  assign new_n6112_ = new_n3436_ & ~new_n6111_;
  assign new_n6113_ = ~new_n6107_ & new_n6112_;
  assign new_n6114_ = ~new_n3436_ & new_n5994_;
  assign new_n6115_ = ~pi0242 & ~new_n6114_;
  assign new_n6116_ = ~new_n6113_ & new_n6115_;
  assign new_n6117_ = pi1134 & ~new_n6116_;
  assign new_n6118_ = ~new_n6049_ & new_n6117_;
  assign po0165 = ~new_n5979_ & ~new_n6118_;
  assign new_n6120_ = pi0057 & pi0059;
  assign new_n6121_ = new_n3100_ & new_n3299_;
  assign new_n6122_ = ~new_n3436_ & ~new_n6121_;
  assign new_n6123_ = ~new_n6120_ & ~new_n6122_;
  assign new_n6124_ = pi0057 & ~new_n6123_;
  assign new_n6125_ = new_n3094_ & new_n3212_;
  assign new_n6126_ = new_n3284_ & new_n6125_;
  assign new_n6127_ = pi0056 & ~new_n6126_;
  assign new_n6128_ = ~pi0054 & new_n3282_;
  assign new_n6129_ = new_n6125_ & new_n6128_;
  assign new_n6130_ = pi0074 & ~new_n6129_;
  assign new_n6131_ = ~pi0055 & ~new_n6130_;
  assign new_n6132_ = ~pi0039 & new_n3094_;
  assign new_n6133_ = pi0038 & ~new_n6132_;
  assign new_n6134_ = ~pi0100 & ~new_n6133_;
  assign new_n6135_ = pi0058 & new_n2521_;
  assign new_n6136_ = ~pi0090 & ~new_n6135_;
  assign new_n6137_ = new_n2505_ & new_n2578_;
  assign new_n6138_ = new_n2683_ & new_n6137_;
  assign new_n6139_ = new_n2590_ & ~new_n6138_;
  assign new_n6140_ = ~new_n2585_ & ~new_n6139_;
  assign new_n6141_ = ~pi0108 & ~new_n6140_;
  assign new_n6142_ = new_n2584_ & ~new_n6141_;
  assign new_n6143_ = ~pi0110 & new_n2698_;
  assign new_n6144_ = ~new_n6142_ & new_n6143_;
  assign new_n6145_ = ~new_n2568_ & ~new_n2575_;
  assign new_n6146_ = ~new_n6144_ & new_n6145_;
  assign new_n6147_ = ~pi0047 & ~new_n6146_;
  assign new_n6148_ = new_n2489_ & ~new_n2571_;
  assign new_n6149_ = ~new_n6147_ & new_n6148_;
  assign new_n6150_ = new_n6136_ & ~new_n6149_;
  assign new_n6151_ = ~new_n2705_ & ~new_n6150_;
  assign new_n6152_ = ~pi0093 & ~new_n6151_;
  assign new_n6153_ = ~pi0841 & new_n2522_;
  assign new_n6154_ = pi0093 & ~new_n6153_;
  assign new_n6155_ = ~new_n6152_ & ~new_n6154_;
  assign new_n6156_ = ~pi0035 & ~new_n6155_;
  assign new_n6157_ = ~pi0070 & ~new_n2524_;
  assign new_n6158_ = ~new_n6156_ & new_n6157_;
  assign new_n6159_ = ~pi0051 & ~new_n6158_;
  assign new_n6160_ = new_n2559_ & ~new_n6159_;
  assign new_n6161_ = new_n2926_ & ~new_n6160_;
  assign new_n6162_ = new_n2556_ & ~new_n6161_;
  assign new_n6163_ = new_n2554_ & ~new_n6162_;
  assign new_n6164_ = ~pi0198 & ~pi0299;
  assign new_n6165_ = ~pi0210 & pi0299;
  assign new_n6166_ = ~new_n6164_ & ~new_n6165_;
  assign new_n6167_ = ~pi0035 & new_n2551_;
  assign new_n6168_ = ~pi0040 & new_n6167_;
  assign new_n6169_ = new_n2735_ & new_n6168_;
  assign new_n6170_ = pi0032 & ~new_n6169_;
  assign new_n6171_ = ~new_n6166_ & ~new_n6170_;
  assign new_n6172_ = ~new_n3367_ & new_n6166_;
  assign new_n6173_ = ~new_n6171_ & ~new_n6172_;
  assign new_n6174_ = ~new_n6163_ & ~new_n6173_;
  assign new_n6175_ = ~pi0095 & ~new_n6174_;
  assign new_n6176_ = ~new_n2726_ & ~new_n6175_;
  assign new_n6177_ = ~pi0039 & ~new_n6176_;
  assign new_n6178_ = pi0603 & ~pi0642;
  assign new_n6179_ = ~pi0614 & ~pi0616;
  assign new_n6180_ = new_n6178_ & new_n6179_;
  assign new_n6181_ = ~pi0662 & pi0680;
  assign new_n6182_ = ~pi0661 & new_n6181_;
  assign new_n6183_ = ~pi0681 & new_n6182_;
  assign po1101 = new_n6180_ | new_n6183_;
  assign new_n6185_ = ~pi0332 & ~pi0468;
  assign new_n6186_ = pi0835 & pi0984;
  assign new_n6187_ = ~pi0252 & ~pi1001;
  assign new_n6188_ = ~pi0979 & ~new_n6187_;
  assign new_n6189_ = ~new_n6186_ & new_n6188_;
  assign new_n6190_ = ~pi0287 & new_n6189_;
  assign new_n6191_ = pi0835 & pi0950;
  assign new_n6192_ = new_n6190_ & new_n6191_;
  assign new_n6193_ = pi1092 & new_n6192_;
  assign new_n6194_ = ~pi0824 & ~pi0829;
  assign new_n6195_ = pi0824 & ~pi1091;
  assign new_n6196_ = pi1093 & ~new_n2733_;
  assign new_n6197_ = ~new_n6195_ & new_n6196_;
  assign new_n6198_ = ~new_n6194_ & ~new_n6197_;
  assign new_n6199_ = new_n6193_ & new_n6198_;
  assign new_n6200_ = ~new_n6185_ & ~new_n6199_;
  assign new_n6201_ = po1101 & ~new_n6200_;
  assign new_n6202_ = new_n3100_ & ~new_n6201_;
  assign new_n6203_ = new_n3094_ & new_n6185_;
  assign new_n6204_ = po1101 & new_n6203_;
  assign new_n6205_ = ~new_n6202_ & ~new_n6204_;
  assign new_n6206_ = ~pi0907 & ~pi0947;
  assign new_n6207_ = ~pi0960 & ~pi0963;
  assign new_n6208_ = ~pi0970 & ~pi0972;
  assign new_n6209_ = ~pi0975 & ~pi0978;
  assign new_n6210_ = new_n6208_ & new_n6209_;
  assign new_n6211_ = new_n6207_ & new_n6210_;
  assign new_n6212_ = new_n6206_ & new_n6211_;
  assign new_n6213_ = ~new_n6205_ & new_n6212_;
  assign new_n6214_ = ~new_n6180_ & ~new_n6185_;
  assign new_n6215_ = ~new_n6183_ & new_n6214_;
  assign new_n6216_ = new_n6199_ & ~new_n6215_;
  assign new_n6217_ = new_n3100_ & ~new_n6216_;
  assign new_n6218_ = ~new_n6212_ & new_n6217_;
  assign new_n6219_ = pi0215 & ~new_n6218_;
  assign new_n6220_ = ~new_n6213_ & new_n6219_;
  assign new_n6221_ = po1101 & ~new_n6185_;
  assign new_n6222_ = new_n6185_ & ~new_n6212_;
  assign new_n6223_ = ~new_n6221_ & ~new_n6222_;
  assign new_n6224_ = new_n2795_ & new_n6192_;
  assign new_n6225_ = pi0216 & pi0221;
  assign new_n6226_ = new_n6224_ & new_n6225_;
  assign new_n6227_ = ~new_n6223_ & new_n6226_;
  assign new_n6228_ = new_n3100_ & ~new_n6227_;
  assign new_n6229_ = ~pi0215 & ~new_n6228_;
  assign new_n6230_ = pi0299 & ~new_n6229_;
  assign new_n6231_ = ~new_n6220_ & new_n6230_;
  assign new_n6232_ = ~pi0969 & ~pi0971;
  assign new_n6233_ = ~pi0974 & ~pi0977;
  assign new_n6234_ = new_n6232_ & new_n6233_;
  assign new_n6235_ = ~pi0587 & ~pi0602;
  assign new_n6236_ = ~pi0961 & ~pi0967;
  assign new_n6237_ = new_n6235_ & new_n6236_;
  assign new_n6238_ = new_n6234_ & new_n6237_;
  assign new_n6239_ = ~new_n6205_ & new_n6238_;
  assign new_n6240_ = new_n6217_ & ~new_n6238_;
  assign new_n6241_ = pi0223 & ~new_n6240_;
  assign new_n6242_ = ~new_n6239_ & new_n6241_;
  assign new_n6243_ = new_n6185_ & ~new_n6238_;
  assign new_n6244_ = ~new_n6221_ & ~new_n6243_;
  assign new_n6245_ = pi0222 & pi0224;
  assign new_n6246_ = new_n6224_ & new_n6245_;
  assign new_n6247_ = ~new_n6244_ & new_n6246_;
  assign new_n6248_ = new_n3100_ & ~new_n6247_;
  assign new_n6249_ = ~pi0223 & ~new_n6248_;
  assign new_n6250_ = ~pi0299 & ~new_n6249_;
  assign new_n6251_ = ~new_n6242_ & new_n6250_;
  assign new_n6252_ = pi0039 & ~new_n6251_;
  assign new_n6253_ = ~new_n6231_ & new_n6252_;
  assign new_n6254_ = ~new_n6177_ & ~new_n6253_;
  assign new_n6255_ = ~pi0038 & ~new_n6254_;
  assign new_n6256_ = new_n6134_ & ~new_n6255_;
  assign new_n6257_ = ~pi0039 & new_n3100_;
  assign new_n6258_ = ~pi0038 & pi0100;
  assign new_n6259_ = new_n6257_ & new_n6258_;
  assign new_n6260_ = ~pi0142 & ~new_n3068_;
  assign new_n6261_ = ~pi0299 & new_n6260_;
  assign new_n6262_ = pi0299 & new_n2993_;
  assign new_n6263_ = ~new_n6261_ & ~new_n6262_;
  assign new_n6264_ = ~new_n3386_ & new_n6263_;
  assign new_n6265_ = ~pi0041 & ~pi0099;
  assign new_n6266_ = ~pi0101 & new_n6265_;
  assign new_n6267_ = ~pi0042 & ~pi0043;
  assign new_n6268_ = ~pi0052 & new_n6267_;
  assign new_n6269_ = ~pi0113 & ~pi0116;
  assign new_n6270_ = ~pi0114 & ~pi0115;
  assign new_n6271_ = new_n6269_ & new_n6270_;
  assign new_n6272_ = new_n6268_ & new_n6271_;
  assign new_n6273_ = new_n6266_ & new_n6272_;
  assign po1057 = pi0044 | ~new_n6273_;
  assign new_n6275_ = ~pi0683 & po1057;
  assign new_n6276_ = pi0129 & pi0250;
  assign new_n6277_ = new_n2799_ & ~new_n6194_;
  assign po0740 = ~pi1093 & new_n6277_;
  assign new_n6279_ = ~pi0250 & ~po0740;
  assign new_n6280_ = ~new_n6276_ & ~new_n6279_;
  assign new_n6281_ = ~new_n6275_ & ~new_n6280_;
  assign new_n6282_ = ~new_n6263_ & po1057;
  assign new_n6283_ = new_n6281_ & new_n6282_;
  assign new_n6284_ = ~new_n6264_ & ~new_n6283_;
  assign new_n6285_ = new_n6259_ & new_n6284_;
  assign new_n6286_ = ~pi0087 & ~new_n6285_;
  assign new_n6287_ = ~new_n6256_ & new_n6286_;
  assign new_n6288_ = pi0087 & ~new_n6125_;
  assign new_n6289_ = ~pi0075 & ~new_n6288_;
  assign new_n6290_ = ~pi0054 & ~pi0092;
  assign new_n6291_ = new_n6289_ & new_n6290_;
  assign new_n6292_ = ~new_n6287_ & new_n6291_;
  assign new_n6293_ = ~pi0074 & ~new_n6292_;
  assign new_n6294_ = new_n6131_ & ~new_n6293_;
  assign new_n6295_ = ~pi0056 & ~new_n6294_;
  assign new_n6296_ = ~new_n6127_ & ~new_n6295_;
  assign new_n6297_ = ~pi0062 & ~new_n6296_;
  assign new_n6298_ = new_n3437_ & new_n6125_;
  assign new_n6299_ = pi0062 & ~new_n6298_;
  assign new_n6300_ = ~pi0059 & ~new_n6299_;
  assign new_n6301_ = ~new_n6297_ & new_n6300_;
  assign new_n6302_ = ~pi0057 & ~new_n6301_;
  assign po0167 = ~new_n6124_ & ~new_n6302_;
  assign new_n6304_ = ~pi0055 & new_n3298_;
  assign new_n6305_ = ~pi0059 & new_n6304_;
  assign new_n6306_ = ~pi0228 & ~new_n6305_;
  assign new_n6307_ = pi0057 & ~new_n6306_;
  assign new_n6308_ = ~new_n6183_ & ~new_n6185_;
  assign new_n6309_ = ~pi0907 & new_n6185_;
  assign new_n6310_ = ~new_n6308_ & ~new_n6309_;
  assign new_n6311_ = ~pi0228 & ~new_n3273_;
  assign new_n6312_ = pi0030 & pi0228;
  assign new_n6313_ = ~new_n3326_ & ~new_n6312_;
  assign new_n6314_ = ~new_n6311_ & ~new_n6313_;
  assign new_n6315_ = new_n6310_ & new_n6314_;
  assign new_n6316_ = new_n6307_ & new_n6315_;
  assign new_n6317_ = ~pi0602 & new_n6185_;
  assign new_n6318_ = ~new_n6308_ & ~new_n6317_;
  assign new_n6319_ = ~pi0091 & ~pi0314;
  assign new_n6320_ = new_n2574_ & ~new_n2575_;
  assign new_n6321_ = pi0085 & new_n2625_;
  assign new_n6322_ = new_n2458_ & ~new_n6321_;
  assign new_n6323_ = new_n2629_ & ~new_n6322_;
  assign new_n6324_ = new_n2467_ & ~new_n6323_;
  assign new_n6325_ = ~new_n2609_ & ~new_n2638_;
  assign new_n6326_ = ~new_n6324_ & new_n6325_;
  assign new_n6327_ = new_n2468_ & new_n6326_;
  assign new_n6328_ = ~new_n2643_ & ~new_n6327_;
  assign new_n6329_ = new_n2641_ & ~new_n6328_;
  assign new_n6330_ = pi0067 & new_n2472_;
  assign new_n6331_ = new_n2606_ & ~new_n6330_;
  assign new_n6332_ = ~new_n6329_ & new_n6331_;
  assign new_n6333_ = new_n2605_ & ~new_n6332_;
  assign new_n6334_ = ~pi0071 & ~new_n6333_;
  assign po1049 = pi0064 | ~new_n2476_;
  assign new_n6336_ = new_n2600_ & ~po1049;
  assign new_n6337_ = ~new_n6334_ & new_n6336_;
  assign new_n6338_ = ~pi0081 & ~new_n6337_;
  assign new_n6339_ = new_n2654_ & new_n6336_;
  assign new_n6340_ = new_n6338_ & ~new_n6339_;
  assign new_n6341_ = ~pi0102 & ~new_n2595_;
  assign new_n6342_ = new_n2452_ & new_n6341_;
  assign new_n6343_ = ~new_n6340_ & new_n6342_;
  assign new_n6344_ = new_n2594_ & ~new_n6343_;
  assign new_n6345_ = new_n2686_ & ~new_n6344_;
  assign new_n6346_ = new_n2504_ & ~new_n6345_;
  assign new_n6347_ = ~new_n2507_ & ~new_n6346_;
  assign new_n6348_ = ~pi0086 & ~new_n6347_;
  assign new_n6349_ = ~pi0046 & new_n2481_;
  assign new_n6350_ = new_n2592_ & new_n6349_;
  assign new_n6351_ = ~new_n6348_ & new_n6350_;
  assign new_n6352_ = new_n2698_ & ~new_n6351_;
  assign new_n6353_ = new_n6320_ & ~new_n6352_;
  assign new_n6354_ = new_n6319_ & ~new_n6353_;
  assign new_n6355_ = pi0091 & ~new_n2533_;
  assign new_n6356_ = ~pi0058 & ~new_n6355_;
  assign new_n6357_ = ~pi0091 & pi0314;
  assign new_n6358_ = ~new_n6338_ & new_n6342_;
  assign new_n6359_ = new_n2594_ & ~new_n6358_;
  assign new_n6360_ = new_n2686_ & ~new_n6359_;
  assign new_n6361_ = new_n2504_ & ~new_n6360_;
  assign new_n6362_ = ~new_n2507_ & ~new_n6361_;
  assign new_n6363_ = ~pi0086 & ~new_n6362_;
  assign new_n6364_ = new_n6350_ & ~new_n6363_;
  assign new_n6365_ = new_n2698_ & ~new_n6364_;
  assign new_n6366_ = new_n6320_ & ~new_n6365_;
  assign new_n6367_ = new_n6357_ & ~new_n6366_;
  assign new_n6368_ = new_n6356_ & ~new_n6367_;
  assign new_n6369_ = ~new_n6354_ & new_n6368_;
  assign new_n6370_ = ~pi0090 & ~new_n6369_;
  assign new_n6371_ = ~new_n2705_ & ~new_n6370_;
  assign new_n6372_ = ~pi0093 & ~new_n6371_;
  assign new_n6373_ = pi0093 & ~new_n2734_;
  assign new_n6374_ = ~pi0035 & ~new_n6373_;
  assign new_n6375_ = ~new_n6372_ & new_n6374_;
  assign new_n6376_ = ~pi0070 & ~new_n6375_;
  assign new_n6377_ = new_n2849_ & ~new_n6376_;
  assign new_n6378_ = ~pi0072 & ~new_n6377_;
  assign new_n6379_ = ~pi0095 & new_n2724_;
  assign new_n6380_ = ~new_n2555_ & new_n6379_;
  assign new_n6381_ = ~new_n6378_ & new_n6380_;
  assign new_n6382_ = ~new_n2943_ & ~new_n6381_;
  assign new_n6383_ = ~pi0841 & new_n2523_;
  assign new_n6384_ = new_n2535_ & new_n6383_;
  assign new_n6385_ = new_n2782_ & new_n6384_;
  assign new_n6386_ = pi0032 & new_n6385_;
  assign new_n6387_ = ~pi0095 & new_n6386_;
  assign new_n6388_ = ~pi0198 & new_n6387_;
  assign new_n6389_ = new_n6382_ & ~new_n6388_;
  assign new_n6390_ = ~pi0228 & ~new_n6389_;
  assign new_n6391_ = ~new_n6312_ & ~new_n6390_;
  assign new_n6392_ = new_n6318_ & ~new_n6391_;
  assign new_n6393_ = ~pi0299 & ~new_n6392_;
  assign new_n6394_ = pi0145 & pi0180;
  assign new_n6395_ = pi0181 & pi0182;
  assign new_n6396_ = new_n6394_ & new_n6395_;
  assign new_n6397_ = ~pi0299 & new_n6396_;
  assign new_n6398_ = ~new_n6393_ & ~new_n6397_;
  assign new_n6399_ = new_n6312_ & new_n6318_;
  assign new_n6400_ = ~new_n6185_ & ~new_n6389_;
  assign new_n6401_ = ~pi0047 & new_n2488_;
  assign new_n6402_ = ~new_n2697_ & ~new_n6351_;
  assign new_n6403_ = new_n6401_ & ~new_n6402_;
  assign new_n6404_ = new_n6319_ & ~new_n6403_;
  assign new_n6405_ = ~new_n2697_ & ~new_n6364_;
  assign new_n6406_ = new_n6401_ & ~new_n6405_;
  assign new_n6407_ = new_n6357_ & ~new_n6406_;
  assign new_n6408_ = new_n6356_ & ~new_n6407_;
  assign new_n6409_ = ~new_n6404_ & new_n6408_;
  assign new_n6410_ = ~pi0090 & ~new_n6409_;
  assign new_n6411_ = ~new_n2705_ & ~new_n6410_;
  assign new_n6412_ = ~pi0093 & ~new_n6411_;
  assign new_n6413_ = new_n6374_ & ~new_n6412_;
  assign new_n6414_ = ~pi0070 & ~new_n6413_;
  assign new_n6415_ = new_n2849_ & ~new_n6414_;
  assign new_n6416_ = ~pi0072 & ~new_n6415_;
  assign new_n6417_ = new_n6380_ & ~new_n6416_;
  assign new_n6418_ = ~new_n2943_ & ~new_n6417_;
  assign new_n6419_ = ~new_n6388_ & new_n6418_;
  assign new_n6420_ = new_n6185_ & ~new_n6419_;
  assign new_n6421_ = ~new_n6400_ & ~new_n6420_;
  assign new_n6422_ = ~pi0228 & new_n6318_;
  assign new_n6423_ = ~new_n6421_ & new_n6422_;
  assign new_n6424_ = ~new_n6399_ & ~new_n6423_;
  assign new_n6425_ = new_n6396_ & ~new_n6424_;
  assign new_n6426_ = ~new_n6398_ & ~new_n6425_;
  assign new_n6427_ = new_n6310_ & new_n6312_;
  assign new_n6428_ = pi0299 & ~new_n6427_;
  assign new_n6429_ = pi0158 & pi0159;
  assign new_n6430_ = pi0160 & pi0197;
  assign new_n6431_ = new_n6429_ & new_n6430_;
  assign new_n6432_ = ~pi0210 & new_n6387_;
  assign new_n6433_ = new_n6382_ & ~new_n6432_;
  assign new_n6434_ = ~new_n6185_ & ~new_n6433_;
  assign new_n6435_ = new_n6418_ & ~new_n6432_;
  assign new_n6436_ = new_n6185_ & ~new_n6435_;
  assign new_n6437_ = ~new_n6434_ & ~new_n6436_;
  assign new_n6438_ = new_n6310_ & ~new_n6437_;
  assign new_n6439_ = new_n6431_ & ~new_n6438_;
  assign new_n6440_ = new_n6310_ & ~new_n6433_;
  assign new_n6441_ = ~new_n6431_ & ~new_n6440_;
  assign new_n6442_ = ~pi0228 & ~new_n6441_;
  assign new_n6443_ = ~new_n6439_ & new_n6442_;
  assign new_n6444_ = new_n6428_ & ~new_n6443_;
  assign new_n6445_ = pi0232 & ~new_n6444_;
  assign new_n6446_ = ~new_n6426_ & new_n6445_;
  assign new_n6447_ = ~pi0228 & new_n6440_;
  assign new_n6448_ = new_n6428_ & ~new_n6447_;
  assign new_n6449_ = ~pi0232 & ~new_n6448_;
  assign new_n6450_ = ~new_n6393_ & new_n6449_;
  assign new_n6451_ = ~new_n6446_ & ~new_n6450_;
  assign new_n6452_ = ~pi0039 & ~new_n6451_;
  assign new_n6453_ = ~pi0215 & pi0221;
  assign new_n6454_ = ~pi0287 & new_n3100_;
  assign new_n6455_ = pi0835 & new_n6189_;
  assign new_n6456_ = new_n6454_ & new_n6455_;
  assign new_n6457_ = pi0824 & pi1093;
  assign new_n6458_ = new_n2799_ & new_n6457_;
  assign new_n6459_ = new_n6456_ & new_n6458_;
  assign new_n6460_ = ~pi1091 & new_n6459_;
  assign new_n6461_ = pi1091 & new_n2732_;
  assign new_n6462_ = new_n6458_ & ~new_n6461_;
  assign new_n6463_ = ~new_n2795_ & ~new_n6462_;
  assign new_n6464_ = pi1091 & ~new_n6463_;
  assign new_n6465_ = new_n6456_ & new_n6464_;
  assign new_n6466_ = ~new_n6460_ & ~new_n6465_;
  assign new_n6467_ = pi0216 & ~new_n6466_;
  assign new_n6468_ = ~pi0829 & ~new_n2732_;
  assign new_n6469_ = pi1091 & ~new_n6468_;
  assign new_n6470_ = new_n6459_ & ~new_n6469_;
  assign new_n6471_ = ~pi0216 & new_n6470_;
  assign new_n6472_ = ~new_n6467_ & ~new_n6471_;
  assign new_n6473_ = ~pi0228 & ~new_n6472_;
  assign new_n6474_ = ~new_n6312_ & ~new_n6473_;
  assign new_n6475_ = new_n6453_ & ~new_n6474_;
  assign new_n6476_ = ~new_n6312_ & ~new_n6475_;
  assign new_n6477_ = new_n6310_ & ~new_n6476_;
  assign new_n6478_ = pi0299 & ~new_n6477_;
  assign new_n6479_ = pi0224 & new_n6466_;
  assign new_n6480_ = pi0222 & ~pi0223;
  assign new_n6481_ = ~pi0224 & ~new_n6470_;
  assign new_n6482_ = new_n6480_ & ~new_n6481_;
  assign new_n6483_ = ~new_n6479_ & new_n6482_;
  assign new_n6484_ = ~pi0228 & new_n6483_;
  assign new_n6485_ = ~new_n6312_ & ~new_n6484_;
  assign new_n6486_ = new_n6318_ & ~new_n6485_;
  assign new_n6487_ = ~pi0299 & ~new_n6486_;
  assign new_n6488_ = pi0039 & ~new_n6487_;
  assign new_n6489_ = ~new_n6478_ & new_n6488_;
  assign new_n6490_ = ~pi0038 & ~new_n6489_;
  assign new_n6491_ = ~new_n6452_ & new_n6490_;
  assign new_n6492_ = pi0299 & new_n6310_;
  assign new_n6493_ = ~pi0299 & new_n6318_;
  assign new_n6494_ = ~new_n6492_ & ~new_n6493_;
  assign new_n6495_ = ~pi0039 & ~new_n6313_;
  assign new_n6496_ = ~new_n6494_ & new_n6495_;
  assign new_n6497_ = new_n6312_ & ~new_n6494_;
  assign new_n6498_ = pi0038 & ~new_n6497_;
  assign new_n6499_ = ~new_n6496_ & new_n6498_;
  assign new_n6500_ = ~new_n6491_ & ~new_n6499_;
  assign new_n6501_ = ~pi0100 & ~new_n6500_;
  assign new_n6502_ = new_n3100_ & ~new_n6280_;
  assign new_n6503_ = pi0683 & po1057;
  assign new_n6504_ = new_n6502_ & new_n6503_;
  assign new_n6505_ = ~new_n6308_ & new_n6504_;
  assign new_n6506_ = new_n6260_ & new_n6505_;
  assign new_n6507_ = pi0252 & ~new_n6260_;
  assign new_n6508_ = pi0252 & new_n6203_;
  assign new_n6509_ = ~new_n6183_ & new_n6508_;
  assign new_n6510_ = pi0252 & new_n3100_;
  assign new_n6511_ = new_n6183_ & new_n6510_;
  assign new_n6512_ = ~new_n6509_ & ~new_n6511_;
  assign new_n6513_ = new_n6507_ & ~new_n6512_;
  assign new_n6514_ = ~new_n6506_ & ~new_n6513_;
  assign new_n6515_ = ~pi0228 & ~new_n6317_;
  assign new_n6516_ = ~new_n6514_ & new_n6515_;
  assign new_n6517_ = ~pi0299 & ~new_n6399_;
  assign new_n6518_ = ~new_n6516_ & new_n6517_;
  assign new_n6519_ = ~new_n2993_ & new_n6512_;
  assign new_n6520_ = new_n2993_ & ~new_n6505_;
  assign new_n6521_ = ~pi0228 & ~new_n6309_;
  assign new_n6522_ = ~new_n6520_ & new_n6521_;
  assign new_n6523_ = ~new_n6519_ & new_n6522_;
  assign new_n6524_ = new_n6428_ & ~new_n6523_;
  assign new_n6525_ = new_n3186_ & ~new_n6524_;
  assign new_n6526_ = ~new_n6518_ & new_n6525_;
  assign new_n6527_ = ~new_n3186_ & new_n6497_;
  assign new_n6528_ = pi0100 & ~new_n6527_;
  assign new_n6529_ = ~new_n6526_ & new_n6528_;
  assign new_n6530_ = ~pi0087 & ~new_n6529_;
  assign new_n6531_ = ~new_n6501_ & new_n6530_;
  assign new_n6532_ = pi0087 & new_n6497_;
  assign new_n6533_ = ~pi0075 & ~new_n6532_;
  assign new_n6534_ = ~new_n6531_ & new_n6533_;
  assign new_n6535_ = ~new_n3227_ & new_n6497_;
  assign new_n6536_ = new_n3246_ & new_n6496_;
  assign new_n6537_ = ~new_n6535_ & ~new_n6536_;
  assign new_n6538_ = pi0075 & new_n6537_;
  assign new_n6539_ = ~pi0092 & ~new_n6538_;
  assign new_n6540_ = ~new_n6534_ & new_n6539_;
  assign new_n6541_ = ~pi0075 & new_n6537_;
  assign new_n6542_ = pi0075 & ~new_n6497_;
  assign new_n6543_ = pi0092 & ~new_n6542_;
  assign new_n6544_ = ~new_n6541_ & new_n6543_;
  assign new_n6545_ = ~pi0054 & ~new_n6544_;
  assign new_n6546_ = ~new_n6540_ & new_n6545_;
  assign new_n6547_ = new_n3242_ & new_n6537_;
  assign new_n6548_ = ~new_n3242_ & ~new_n6497_;
  assign new_n6549_ = ~new_n6547_ & ~new_n6548_;
  assign new_n6550_ = pi0054 & ~new_n6549_;
  assign new_n6551_ = ~pi0074 & ~new_n6550_;
  assign new_n6552_ = ~new_n6546_ & new_n6551_;
  assign new_n6553_ = ~pi0054 & new_n6547_;
  assign new_n6554_ = ~pi0054 & new_n3242_;
  assign new_n6555_ = ~new_n6497_ & ~new_n6554_;
  assign new_n6556_ = pi0074 & ~new_n6555_;
  assign new_n6557_ = ~new_n6553_ & new_n6556_;
  assign new_n6558_ = ~pi0055 & ~new_n6557_;
  assign new_n6559_ = ~new_n6552_ & new_n6558_;
  assign new_n6560_ = pi0055 & ~new_n6315_;
  assign new_n6561_ = new_n3298_ & ~new_n6560_;
  assign new_n6562_ = ~new_n6559_ & new_n6561_;
  assign new_n6563_ = ~new_n3298_ & new_n6427_;
  assign new_n6564_ = ~pi0059 & ~new_n6563_;
  assign new_n6565_ = ~new_n6562_ & new_n6564_;
  assign new_n6566_ = ~pi0228 & ~new_n6304_;
  assign new_n6567_ = new_n6315_ & ~new_n6566_;
  assign new_n6568_ = pi0059 & ~new_n6567_;
  assign new_n6569_ = ~pi0057 & ~new_n6568_;
  assign new_n6570_ = ~new_n6565_ & new_n6569_;
  assign po0171 = ~new_n6316_ & ~new_n6570_;
  assign new_n6572_ = ~pi0947 & new_n6185_;
  assign new_n6573_ = ~new_n6214_ & ~new_n6572_;
  assign new_n6574_ = new_n6314_ & new_n6573_;
  assign new_n6575_ = new_n6307_ & new_n6574_;
  assign new_n6576_ = ~pi0587 & new_n6185_;
  assign new_n6577_ = ~new_n6214_ & ~new_n6576_;
  assign new_n6578_ = new_n6312_ & new_n6577_;
  assign new_n6579_ = ~pi0228 & new_n6577_;
  assign new_n6580_ = ~new_n6421_ & new_n6579_;
  assign new_n6581_ = ~new_n6578_ & ~new_n6580_;
  assign new_n6582_ = new_n6396_ & ~new_n6581_;
  assign new_n6583_ = ~new_n6391_ & new_n6577_;
  assign new_n6584_ = ~new_n6396_ & new_n6583_;
  assign new_n6585_ = ~pi0299 & ~new_n6584_;
  assign new_n6586_ = ~new_n6582_ & new_n6585_;
  assign new_n6587_ = new_n6312_ & new_n6573_;
  assign new_n6588_ = pi0299 & ~new_n6587_;
  assign new_n6589_ = ~new_n6437_ & new_n6573_;
  assign new_n6590_ = new_n6431_ & ~new_n6589_;
  assign new_n6591_ = ~new_n6433_ & new_n6573_;
  assign new_n6592_ = ~new_n6431_ & ~new_n6591_;
  assign new_n6593_ = ~pi0228 & ~new_n6592_;
  assign new_n6594_ = ~new_n6590_ & new_n6593_;
  assign new_n6595_ = new_n6588_ & ~new_n6594_;
  assign new_n6596_ = pi0232 & ~new_n6595_;
  assign new_n6597_ = ~new_n6586_ & new_n6596_;
  assign new_n6598_ = ~pi0299 & ~new_n6583_;
  assign new_n6599_ = ~pi0228 & new_n6591_;
  assign new_n6600_ = new_n6588_ & ~new_n6599_;
  assign new_n6601_ = ~pi0232 & ~new_n6600_;
  assign new_n6602_ = ~new_n6598_ & new_n6601_;
  assign new_n6603_ = ~new_n6597_ & ~new_n6602_;
  assign new_n6604_ = ~pi0039 & ~new_n6603_;
  assign new_n6605_ = pi0299 & new_n6453_;
  assign new_n6606_ = ~new_n6588_ & ~new_n6605_;
  assign new_n6607_ = new_n6475_ & new_n6573_;
  assign new_n6608_ = ~new_n6606_ & ~new_n6607_;
  assign new_n6609_ = ~new_n6485_ & new_n6577_;
  assign new_n6610_ = ~pi0299 & ~new_n6609_;
  assign new_n6611_ = pi0039 & ~new_n6610_;
  assign new_n6612_ = ~new_n6608_ & new_n6611_;
  assign new_n6613_ = ~pi0038 & ~new_n6612_;
  assign new_n6614_ = ~new_n6604_ & new_n6613_;
  assign new_n6615_ = pi0299 & ~new_n6573_;
  assign new_n6616_ = ~pi0299 & ~new_n6577_;
  assign new_n6617_ = ~new_n6615_ & ~new_n6616_;
  assign new_n6618_ = new_n6495_ & new_n6617_;
  assign new_n6619_ = new_n6312_ & new_n6617_;
  assign new_n6620_ = pi0038 & ~new_n6619_;
  assign new_n6621_ = ~new_n6618_ & new_n6620_;
  assign new_n6622_ = ~new_n6614_ & ~new_n6621_;
  assign new_n6623_ = ~pi0100 & ~new_n6622_;
  assign new_n6624_ = ~pi0228 & new_n3068_;
  assign new_n6625_ = ~new_n6180_ & ~new_n6508_;
  assign new_n6626_ = new_n6180_ & ~new_n6510_;
  assign new_n6627_ = ~new_n6625_ & ~new_n6626_;
  assign new_n6628_ = ~new_n6576_ & new_n6627_;
  assign new_n6629_ = new_n6624_ & ~new_n6628_;
  assign new_n6630_ = pi0142 & ~new_n6627_;
  assign new_n6631_ = ~new_n6214_ & new_n6504_;
  assign new_n6632_ = ~pi0142 & ~new_n6631_;
  assign new_n6633_ = new_n6180_ & ~new_n6185_;
  assign new_n6634_ = ~pi0587 & ~new_n6633_;
  assign new_n6635_ = ~pi0228 & ~new_n6634_;
  assign new_n6636_ = ~new_n6632_ & new_n6635_;
  assign new_n6637_ = ~new_n6630_ & new_n6636_;
  assign new_n6638_ = ~new_n6578_ & ~new_n6624_;
  assign new_n6639_ = ~new_n6637_ & new_n6638_;
  assign new_n6640_ = ~new_n6629_ & ~new_n6639_;
  assign new_n6641_ = ~pi0299 & ~new_n6640_;
  assign new_n6642_ = new_n2993_ & ~new_n6572_;
  assign new_n6643_ = new_n6631_ & new_n6642_;
  assign new_n6644_ = ~pi0947 & ~new_n6633_;
  assign new_n6645_ = ~new_n2993_ & ~new_n6644_;
  assign new_n6646_ = new_n6627_ & new_n6645_;
  assign new_n6647_ = ~new_n6643_ & ~new_n6646_;
  assign new_n6648_ = ~pi0228 & ~new_n6647_;
  assign new_n6649_ = new_n6588_ & ~new_n6648_;
  assign new_n6650_ = new_n3186_ & ~new_n6649_;
  assign new_n6651_ = ~new_n6641_ & new_n6650_;
  assign new_n6652_ = ~new_n3186_ & new_n6619_;
  assign new_n6653_ = pi0100 & ~new_n6652_;
  assign new_n6654_ = ~new_n6651_ & new_n6653_;
  assign new_n6655_ = ~pi0087 & ~new_n6654_;
  assign new_n6656_ = ~new_n6623_ & new_n6655_;
  assign new_n6657_ = pi0087 & new_n6619_;
  assign new_n6658_ = ~pi0075 & ~new_n6657_;
  assign new_n6659_ = ~new_n6656_ & new_n6658_;
  assign new_n6660_ = ~new_n3227_ & new_n6619_;
  assign new_n6661_ = new_n3246_ & new_n6618_;
  assign new_n6662_ = ~new_n6660_ & ~new_n6661_;
  assign new_n6663_ = pi0075 & new_n6662_;
  assign new_n6664_ = ~pi0092 & ~new_n6663_;
  assign new_n6665_ = ~new_n6659_ & new_n6664_;
  assign new_n6666_ = ~pi0075 & new_n6662_;
  assign new_n6667_ = pi0075 & ~new_n6619_;
  assign new_n6668_ = pi0092 & ~new_n6667_;
  assign new_n6669_ = ~new_n6666_ & new_n6668_;
  assign new_n6670_ = ~pi0054 & ~new_n6669_;
  assign new_n6671_ = ~new_n6665_ & new_n6670_;
  assign new_n6672_ = new_n3242_ & new_n6662_;
  assign new_n6673_ = ~new_n3242_ & ~new_n6619_;
  assign new_n6674_ = ~new_n6672_ & ~new_n6673_;
  assign new_n6675_ = pi0054 & ~new_n6674_;
  assign new_n6676_ = ~pi0074 & ~new_n6675_;
  assign new_n6677_ = ~new_n6671_ & new_n6676_;
  assign new_n6678_ = ~pi0054 & new_n6672_;
  assign new_n6679_ = ~new_n6554_ & ~new_n6619_;
  assign new_n6680_ = pi0074 & ~new_n6679_;
  assign new_n6681_ = ~new_n6678_ & new_n6680_;
  assign new_n6682_ = ~pi0055 & ~new_n6681_;
  assign new_n6683_ = ~new_n6677_ & new_n6682_;
  assign new_n6684_ = pi0055 & ~new_n6574_;
  assign new_n6685_ = new_n3298_ & ~new_n6684_;
  assign new_n6686_ = ~new_n6683_ & new_n6685_;
  assign new_n6687_ = ~new_n3298_ & new_n6587_;
  assign new_n6688_ = ~pi0059 & ~new_n6687_;
  assign new_n6689_ = ~new_n6686_ & new_n6688_;
  assign new_n6690_ = ~new_n6566_ & new_n6574_;
  assign new_n6691_ = pi0059 & ~new_n6690_;
  assign new_n6692_ = ~pi0057 & ~new_n6691_;
  assign new_n6693_ = ~new_n6689_ & new_n6692_;
  assign po0172 = ~new_n6575_ & ~new_n6693_;
  assign new_n6695_ = pi0030 & new_n6185_;
  assign new_n6696_ = pi0228 & new_n6695_;
  assign new_n6697_ = pi0970 & new_n6696_;
  assign new_n6698_ = ~pi0228 & pi0970;
  assign new_n6699_ = new_n6203_ & new_n6698_;
  assign new_n6700_ = new_n3273_ & new_n6699_;
  assign new_n6701_ = new_n6305_ & new_n6700_;
  assign new_n6702_ = ~new_n6697_ & ~new_n6701_;
  assign new_n6703_ = pi0057 & ~new_n6702_;
  assign new_n6704_ = pi0299 & ~new_n6697_;
  assign new_n6705_ = new_n6185_ & ~new_n6433_;
  assign new_n6706_ = new_n6698_ & new_n6705_;
  assign new_n6707_ = new_n6704_ & ~new_n6706_;
  assign new_n6708_ = pi0299 & new_n6429_;
  assign new_n6709_ = ~new_n6707_ & ~new_n6708_;
  assign new_n6710_ = new_n6430_ & ~new_n6436_;
  assign new_n6711_ = ~new_n6430_ & new_n6433_;
  assign new_n6712_ = ~new_n6710_ & ~new_n6711_;
  assign new_n6713_ = new_n6185_ & new_n6712_;
  assign new_n6714_ = new_n6698_ & new_n6713_;
  assign new_n6715_ = ~new_n6697_ & ~new_n6714_;
  assign new_n6716_ = new_n6429_ & ~new_n6715_;
  assign new_n6717_ = ~new_n6709_ & ~new_n6716_;
  assign new_n6718_ = new_n6185_ & ~new_n6391_;
  assign new_n6719_ = ~new_n6396_ & ~new_n6718_;
  assign new_n6720_ = ~pi0228 & new_n6420_;
  assign new_n6721_ = ~new_n6389_ & ~new_n6396_;
  assign new_n6722_ = ~new_n6696_ & ~new_n6721_;
  assign new_n6723_ = ~new_n6720_ & new_n6722_;
  assign new_n6724_ = ~new_n6719_ & ~new_n6723_;
  assign new_n6725_ = pi0967 & new_n6724_;
  assign new_n6726_ = ~pi0299 & ~new_n6725_;
  assign new_n6727_ = pi0232 & ~new_n6726_;
  assign new_n6728_ = ~new_n6717_ & new_n6727_;
  assign new_n6729_ = pi0967 & new_n6718_;
  assign new_n6730_ = ~pi0299 & ~new_n6729_;
  assign new_n6731_ = ~pi0232 & ~new_n6707_;
  assign new_n6732_ = ~new_n6730_ & new_n6731_;
  assign new_n6733_ = ~new_n6728_ & ~new_n6732_;
  assign new_n6734_ = ~pi0039 & ~new_n6733_;
  assign new_n6735_ = pi0299 & pi0970;
  assign new_n6736_ = new_n6453_ & ~new_n6472_;
  assign new_n6737_ = new_n6185_ & new_n6736_;
  assign new_n6738_ = ~pi0228 & ~new_n6737_;
  assign new_n6739_ = new_n6735_ & ~new_n6738_;
  assign new_n6740_ = ~pi0299 & pi0967;
  assign new_n6741_ = new_n6185_ & new_n6483_;
  assign new_n6742_ = ~pi0228 & ~new_n6741_;
  assign new_n6743_ = new_n6740_ & ~new_n6742_;
  assign new_n6744_ = ~new_n6739_ & ~new_n6743_;
  assign new_n6745_ = pi0228 & ~new_n6695_;
  assign new_n6746_ = pi0039 & ~new_n6745_;
  assign new_n6747_ = ~new_n6744_ & new_n6746_;
  assign new_n6748_ = ~pi0038 & ~new_n6747_;
  assign new_n6749_ = ~new_n6734_ & new_n6748_;
  assign new_n6750_ = ~pi0228 & ~new_n6203_;
  assign new_n6751_ = ~new_n6745_ & ~new_n6750_;
  assign new_n6752_ = pi0967 & new_n6751_;
  assign new_n6753_ = ~pi0299 & ~new_n6752_;
  assign new_n6754_ = ~new_n6699_ & new_n6704_;
  assign new_n6755_ = ~pi0039 & ~new_n6754_;
  assign new_n6756_ = ~new_n6753_ & new_n6755_;
  assign new_n6757_ = ~new_n6735_ & ~new_n6740_;
  assign new_n6758_ = new_n6696_ & ~new_n6757_;
  assign new_n6759_ = pi0039 & new_n6758_;
  assign new_n6760_ = pi0038 & ~new_n6759_;
  assign new_n6761_ = ~new_n6756_ & new_n6760_;
  assign new_n6762_ = ~new_n6749_ & ~new_n6761_;
  assign new_n6763_ = ~pi0100 & ~new_n6762_;
  assign new_n6764_ = new_n6185_ & new_n6504_;
  assign new_n6765_ = new_n6260_ & new_n6764_;
  assign new_n6766_ = ~new_n6260_ & new_n6508_;
  assign new_n6767_ = ~pi0228 & ~new_n6766_;
  assign new_n6768_ = ~new_n6765_ & new_n6767_;
  assign new_n6769_ = ~new_n6745_ & ~new_n6768_;
  assign new_n6770_ = pi0967 & new_n6769_;
  assign new_n6771_ = ~pi0299 & ~new_n6770_;
  assign new_n6772_ = new_n2993_ & ~new_n6764_;
  assign new_n6773_ = ~new_n2993_ & ~new_n6508_;
  assign new_n6774_ = ~pi0228 & ~new_n6773_;
  assign new_n6775_ = ~new_n6772_ & new_n6774_;
  assign new_n6776_ = pi0970 & new_n6775_;
  assign new_n6777_ = new_n6704_ & ~new_n6776_;
  assign new_n6778_ = new_n3186_ & ~new_n6777_;
  assign new_n6779_ = ~new_n6771_ & new_n6778_;
  assign new_n6780_ = ~new_n3186_ & new_n6758_;
  assign new_n6781_ = pi0100 & ~new_n6780_;
  assign new_n6782_ = ~new_n6779_ & new_n6781_;
  assign new_n6783_ = ~pi0087 & ~new_n6782_;
  assign new_n6784_ = ~new_n6763_ & new_n6783_;
  assign new_n6785_ = pi0087 & new_n6758_;
  assign new_n6786_ = ~pi0075 & ~new_n6785_;
  assign new_n6787_ = ~new_n6784_ & new_n6786_;
  assign new_n6788_ = ~new_n3227_ & new_n6758_;
  assign new_n6789_ = new_n3246_ & new_n6756_;
  assign new_n6790_ = ~new_n6788_ & ~new_n6789_;
  assign new_n6791_ = pi0075 & new_n6790_;
  assign new_n6792_ = ~pi0092 & ~new_n6791_;
  assign new_n6793_ = ~new_n6787_ & new_n6792_;
  assign new_n6794_ = ~pi0075 & new_n6790_;
  assign new_n6795_ = pi0075 & ~new_n6758_;
  assign new_n6796_ = pi0092 & ~new_n6795_;
  assign new_n6797_ = ~new_n6794_ & new_n6796_;
  assign new_n6798_ = ~pi0054 & ~new_n6797_;
  assign new_n6799_ = ~new_n6793_ & new_n6798_;
  assign new_n6800_ = new_n3242_ & new_n6790_;
  assign new_n6801_ = ~new_n3242_ & ~new_n6758_;
  assign new_n6802_ = ~new_n6800_ & ~new_n6801_;
  assign new_n6803_ = pi0054 & ~new_n6802_;
  assign new_n6804_ = ~pi0074 & ~new_n6803_;
  assign new_n6805_ = ~new_n6799_ & new_n6804_;
  assign new_n6806_ = ~pi0054 & new_n6800_;
  assign new_n6807_ = ~new_n6554_ & ~new_n6758_;
  assign new_n6808_ = pi0074 & ~new_n6807_;
  assign new_n6809_ = ~new_n6806_ & new_n6808_;
  assign new_n6810_ = ~pi0055 & ~new_n6809_;
  assign new_n6811_ = ~new_n6805_ & new_n6810_;
  assign new_n6812_ = pi0055 & ~new_n6697_;
  assign new_n6813_ = ~new_n6700_ & new_n6812_;
  assign new_n6814_ = new_n3298_ & ~new_n6813_;
  assign new_n6815_ = ~new_n6811_ & new_n6814_;
  assign new_n6816_ = ~new_n3298_ & new_n6697_;
  assign new_n6817_ = ~pi0059 & ~new_n6816_;
  assign new_n6818_ = ~new_n6815_ & new_n6817_;
  assign new_n6819_ = new_n6304_ & new_n6700_;
  assign new_n6820_ = pi0059 & ~new_n6697_;
  assign new_n6821_ = ~new_n6819_ & new_n6820_;
  assign new_n6822_ = ~pi0057 & ~new_n6821_;
  assign new_n6823_ = ~new_n6818_ & new_n6822_;
  assign po0173 = ~new_n6703_ & ~new_n6823_;
  assign new_n6825_ = pi0972 & new_n6696_;
  assign new_n6826_ = ~pi0228 & pi0972;
  assign new_n6827_ = new_n6203_ & new_n6826_;
  assign new_n6828_ = new_n3273_ & new_n6827_;
  assign new_n6829_ = new_n6305_ & new_n6828_;
  assign new_n6830_ = ~new_n6825_ & ~new_n6829_;
  assign new_n6831_ = pi0057 & ~new_n6830_;
  assign new_n6832_ = pi0299 & ~new_n6825_;
  assign new_n6833_ = new_n6705_ & new_n6826_;
  assign new_n6834_ = new_n6832_ & ~new_n6833_;
  assign new_n6835_ = ~new_n6708_ & ~new_n6834_;
  assign new_n6836_ = new_n6713_ & new_n6826_;
  assign new_n6837_ = ~new_n6825_ & ~new_n6836_;
  assign new_n6838_ = new_n6429_ & ~new_n6837_;
  assign new_n6839_ = ~new_n6835_ & ~new_n6838_;
  assign new_n6840_ = pi0961 & new_n6724_;
  assign new_n6841_ = ~pi0299 & ~new_n6840_;
  assign new_n6842_ = pi0232 & ~new_n6841_;
  assign new_n6843_ = ~new_n6839_ & new_n6842_;
  assign new_n6844_ = pi0961 & new_n6718_;
  assign new_n6845_ = ~pi0299 & ~new_n6844_;
  assign new_n6846_ = ~pi0232 & ~new_n6834_;
  assign new_n6847_ = ~new_n6845_ & new_n6846_;
  assign new_n6848_ = ~new_n6843_ & ~new_n6847_;
  assign new_n6849_ = ~pi0039 & ~new_n6848_;
  assign new_n6850_ = ~pi0299 & pi0961;
  assign new_n6851_ = ~new_n6742_ & new_n6850_;
  assign new_n6852_ = pi0299 & pi0972;
  assign new_n6853_ = ~new_n6738_ & new_n6852_;
  assign new_n6854_ = ~new_n6851_ & ~new_n6853_;
  assign new_n6855_ = new_n6746_ & ~new_n6854_;
  assign new_n6856_ = ~pi0038 & ~new_n6855_;
  assign new_n6857_ = ~new_n6849_ & new_n6856_;
  assign new_n6858_ = pi0961 & new_n6751_;
  assign new_n6859_ = ~pi0299 & ~new_n6858_;
  assign new_n6860_ = ~new_n6827_ & new_n6832_;
  assign new_n6861_ = ~pi0039 & ~new_n6860_;
  assign new_n6862_ = ~new_n6859_ & new_n6861_;
  assign new_n6863_ = ~new_n6850_ & ~new_n6852_;
  assign new_n6864_ = new_n6696_ & ~new_n6863_;
  assign new_n6865_ = pi0039 & new_n6864_;
  assign new_n6866_ = pi0038 & ~new_n6865_;
  assign new_n6867_ = ~new_n6862_ & new_n6866_;
  assign new_n6868_ = ~new_n6857_ & ~new_n6867_;
  assign new_n6869_ = ~pi0100 & ~new_n6868_;
  assign new_n6870_ = pi0961 & new_n6769_;
  assign new_n6871_ = ~pi0299 & ~new_n6870_;
  assign new_n6872_ = pi0972 & new_n6775_;
  assign new_n6873_ = new_n6832_ & ~new_n6872_;
  assign new_n6874_ = new_n3186_ & ~new_n6873_;
  assign new_n6875_ = ~new_n6871_ & new_n6874_;
  assign new_n6876_ = ~new_n3186_ & new_n6864_;
  assign new_n6877_ = pi0100 & ~new_n6876_;
  assign new_n6878_ = ~new_n6875_ & new_n6877_;
  assign new_n6879_ = ~pi0087 & ~new_n6878_;
  assign new_n6880_ = ~new_n6869_ & new_n6879_;
  assign new_n6881_ = pi0087 & new_n6864_;
  assign new_n6882_ = ~pi0075 & ~new_n6881_;
  assign new_n6883_ = ~new_n6880_ & new_n6882_;
  assign new_n6884_ = ~new_n3227_ & new_n6864_;
  assign new_n6885_ = new_n3246_ & new_n6862_;
  assign new_n6886_ = ~new_n6884_ & ~new_n6885_;
  assign new_n6887_ = pi0075 & new_n6886_;
  assign new_n6888_ = ~pi0092 & ~new_n6887_;
  assign new_n6889_ = ~new_n6883_ & new_n6888_;
  assign new_n6890_ = ~pi0075 & new_n6886_;
  assign new_n6891_ = pi0075 & ~new_n6864_;
  assign new_n6892_ = pi0092 & ~new_n6891_;
  assign new_n6893_ = ~new_n6890_ & new_n6892_;
  assign new_n6894_ = ~pi0054 & ~new_n6893_;
  assign new_n6895_ = ~new_n6889_ & new_n6894_;
  assign new_n6896_ = new_n3242_ & new_n6886_;
  assign new_n6897_ = ~new_n3242_ & ~new_n6864_;
  assign new_n6898_ = ~new_n6896_ & ~new_n6897_;
  assign new_n6899_ = pi0054 & ~new_n6898_;
  assign new_n6900_ = ~pi0074 & ~new_n6899_;
  assign new_n6901_ = ~new_n6895_ & new_n6900_;
  assign new_n6902_ = ~pi0054 & new_n6896_;
  assign new_n6903_ = ~new_n6554_ & ~new_n6864_;
  assign new_n6904_ = pi0074 & ~new_n6903_;
  assign new_n6905_ = ~new_n6902_ & new_n6904_;
  assign new_n6906_ = ~pi0055 & ~new_n6905_;
  assign new_n6907_ = ~new_n6901_ & new_n6906_;
  assign new_n6908_ = pi0055 & ~new_n6825_;
  assign new_n6909_ = ~new_n6828_ & new_n6908_;
  assign new_n6910_ = new_n3298_ & ~new_n6909_;
  assign new_n6911_ = ~new_n6907_ & new_n6910_;
  assign new_n6912_ = ~new_n3298_ & new_n6825_;
  assign new_n6913_ = ~pi0059 & ~new_n6912_;
  assign new_n6914_ = ~new_n6911_ & new_n6913_;
  assign new_n6915_ = new_n6304_ & new_n6828_;
  assign new_n6916_ = pi0059 & ~new_n6825_;
  assign new_n6917_ = ~new_n6915_ & new_n6916_;
  assign new_n6918_ = ~pi0057 & ~new_n6917_;
  assign new_n6919_ = ~new_n6914_ & new_n6918_;
  assign po0174 = ~new_n6831_ & ~new_n6919_;
  assign new_n6921_ = pi0960 & new_n6696_;
  assign new_n6922_ = ~pi0228 & pi0960;
  assign new_n6923_ = new_n6203_ & new_n6922_;
  assign new_n6924_ = new_n3273_ & new_n6923_;
  assign new_n6925_ = new_n6305_ & new_n6924_;
  assign new_n6926_ = ~new_n6921_ & ~new_n6925_;
  assign new_n6927_ = pi0057 & ~new_n6926_;
  assign new_n6928_ = pi0299 & ~new_n6921_;
  assign new_n6929_ = new_n6705_ & new_n6922_;
  assign new_n6930_ = new_n6928_ & ~new_n6929_;
  assign new_n6931_ = ~new_n6708_ & ~new_n6930_;
  assign new_n6932_ = new_n6713_ & new_n6922_;
  assign new_n6933_ = ~new_n6921_ & ~new_n6932_;
  assign new_n6934_ = new_n6429_ & ~new_n6933_;
  assign new_n6935_ = ~new_n6931_ & ~new_n6934_;
  assign new_n6936_ = pi0977 & new_n6724_;
  assign new_n6937_ = ~pi0299 & ~new_n6936_;
  assign new_n6938_ = pi0232 & ~new_n6937_;
  assign new_n6939_ = ~new_n6935_ & new_n6938_;
  assign new_n6940_ = pi0977 & new_n6718_;
  assign new_n6941_ = ~pi0299 & ~new_n6940_;
  assign new_n6942_ = ~pi0232 & ~new_n6930_;
  assign new_n6943_ = ~new_n6941_ & new_n6942_;
  assign new_n6944_ = ~new_n6939_ & ~new_n6943_;
  assign new_n6945_ = ~pi0039 & ~new_n6944_;
  assign new_n6946_ = ~pi0299 & pi0977;
  assign new_n6947_ = ~new_n6742_ & new_n6946_;
  assign new_n6948_ = pi0299 & pi0960;
  assign new_n6949_ = ~new_n6738_ & new_n6948_;
  assign new_n6950_ = ~new_n6947_ & ~new_n6949_;
  assign new_n6951_ = new_n6746_ & ~new_n6950_;
  assign new_n6952_ = ~pi0038 & ~new_n6951_;
  assign new_n6953_ = ~new_n6945_ & new_n6952_;
  assign new_n6954_ = pi0977 & new_n6751_;
  assign new_n6955_ = ~pi0299 & ~new_n6954_;
  assign new_n6956_ = ~new_n6923_ & new_n6928_;
  assign new_n6957_ = ~pi0039 & ~new_n6956_;
  assign new_n6958_ = ~new_n6955_ & new_n6957_;
  assign new_n6959_ = ~new_n6946_ & ~new_n6948_;
  assign new_n6960_ = new_n6696_ & ~new_n6959_;
  assign new_n6961_ = pi0039 & new_n6960_;
  assign new_n6962_ = pi0038 & ~new_n6961_;
  assign new_n6963_ = ~new_n6958_ & new_n6962_;
  assign new_n6964_ = ~new_n6953_ & ~new_n6963_;
  assign new_n6965_ = ~pi0100 & ~new_n6964_;
  assign new_n6966_ = pi0977 & new_n6769_;
  assign new_n6967_ = ~pi0299 & ~new_n6966_;
  assign new_n6968_ = pi0960 & new_n6775_;
  assign new_n6969_ = new_n6928_ & ~new_n6968_;
  assign new_n6970_ = new_n3186_ & ~new_n6969_;
  assign new_n6971_ = ~new_n6967_ & new_n6970_;
  assign new_n6972_ = ~new_n3186_ & new_n6960_;
  assign new_n6973_ = pi0100 & ~new_n6972_;
  assign new_n6974_ = ~new_n6971_ & new_n6973_;
  assign new_n6975_ = ~pi0087 & ~new_n6974_;
  assign new_n6976_ = ~new_n6965_ & new_n6975_;
  assign new_n6977_ = pi0087 & new_n6960_;
  assign new_n6978_ = ~pi0075 & ~new_n6977_;
  assign new_n6979_ = ~new_n6976_ & new_n6978_;
  assign new_n6980_ = ~new_n3227_ & new_n6960_;
  assign new_n6981_ = new_n3246_ & new_n6958_;
  assign new_n6982_ = ~new_n6980_ & ~new_n6981_;
  assign new_n6983_ = pi0075 & new_n6982_;
  assign new_n6984_ = ~pi0092 & ~new_n6983_;
  assign new_n6985_ = ~new_n6979_ & new_n6984_;
  assign new_n6986_ = ~pi0075 & new_n6982_;
  assign new_n6987_ = pi0075 & ~new_n6960_;
  assign new_n6988_ = pi0092 & ~new_n6987_;
  assign new_n6989_ = ~new_n6986_ & new_n6988_;
  assign new_n6990_ = ~pi0054 & ~new_n6989_;
  assign new_n6991_ = ~new_n6985_ & new_n6990_;
  assign new_n6992_ = new_n3242_ & new_n6982_;
  assign new_n6993_ = ~new_n3242_ & ~new_n6960_;
  assign new_n6994_ = ~new_n6992_ & ~new_n6993_;
  assign new_n6995_ = pi0054 & ~new_n6994_;
  assign new_n6996_ = ~pi0074 & ~new_n6995_;
  assign new_n6997_ = ~new_n6991_ & new_n6996_;
  assign new_n6998_ = ~pi0054 & new_n6992_;
  assign new_n6999_ = ~new_n6554_ & ~new_n6960_;
  assign new_n7000_ = pi0074 & ~new_n6999_;
  assign new_n7001_ = ~new_n6998_ & new_n7000_;
  assign new_n7002_ = ~pi0055 & ~new_n7001_;
  assign new_n7003_ = ~new_n6997_ & new_n7002_;
  assign new_n7004_ = pi0055 & ~new_n6921_;
  assign new_n7005_ = ~new_n6924_ & new_n7004_;
  assign new_n7006_ = new_n3298_ & ~new_n7005_;
  assign new_n7007_ = ~new_n7003_ & new_n7006_;
  assign new_n7008_ = ~new_n3298_ & new_n6921_;
  assign new_n7009_ = ~pi0059 & ~new_n7008_;
  assign new_n7010_ = ~new_n7007_ & new_n7009_;
  assign new_n7011_ = new_n6304_ & new_n6924_;
  assign new_n7012_ = pi0059 & ~new_n6921_;
  assign new_n7013_ = ~new_n7011_ & new_n7012_;
  assign new_n7014_ = ~pi0057 & ~new_n7013_;
  assign new_n7015_ = ~new_n7010_ & new_n7014_;
  assign po0175 = ~new_n6927_ & ~new_n7015_;
  assign new_n7017_ = pi0963 & new_n6696_;
  assign new_n7018_ = ~pi0228 & pi0963;
  assign new_n7019_ = new_n6203_ & new_n7018_;
  assign new_n7020_ = new_n3273_ & new_n7019_;
  assign new_n7021_ = new_n6305_ & new_n7020_;
  assign new_n7022_ = ~new_n7017_ & ~new_n7021_;
  assign new_n7023_ = pi0057 & ~new_n7022_;
  assign new_n7024_ = pi0299 & ~new_n7017_;
  assign new_n7025_ = new_n6705_ & new_n7018_;
  assign new_n7026_ = new_n7024_ & ~new_n7025_;
  assign new_n7027_ = ~new_n6708_ & ~new_n7026_;
  assign new_n7028_ = new_n6713_ & new_n7018_;
  assign new_n7029_ = ~new_n7017_ & ~new_n7028_;
  assign new_n7030_ = new_n6429_ & ~new_n7029_;
  assign new_n7031_ = ~new_n7027_ & ~new_n7030_;
  assign new_n7032_ = pi0969 & new_n6724_;
  assign new_n7033_ = ~pi0299 & ~new_n7032_;
  assign new_n7034_ = pi0232 & ~new_n7033_;
  assign new_n7035_ = ~new_n7031_ & new_n7034_;
  assign new_n7036_ = pi0969 & new_n6718_;
  assign new_n7037_ = ~pi0299 & ~new_n7036_;
  assign new_n7038_ = ~pi0232 & ~new_n7026_;
  assign new_n7039_ = ~new_n7037_ & new_n7038_;
  assign new_n7040_ = ~new_n7035_ & ~new_n7039_;
  assign new_n7041_ = ~pi0039 & ~new_n7040_;
  assign new_n7042_ = ~pi0299 & pi0969;
  assign new_n7043_ = ~new_n6742_ & new_n7042_;
  assign new_n7044_ = pi0299 & pi0963;
  assign new_n7045_ = ~new_n6738_ & new_n7044_;
  assign new_n7046_ = ~new_n7043_ & ~new_n7045_;
  assign new_n7047_ = new_n6746_ & ~new_n7046_;
  assign new_n7048_ = ~pi0038 & ~new_n7047_;
  assign new_n7049_ = ~new_n7041_ & new_n7048_;
  assign new_n7050_ = pi0969 & new_n6751_;
  assign new_n7051_ = ~pi0299 & ~new_n7050_;
  assign new_n7052_ = ~new_n7019_ & new_n7024_;
  assign new_n7053_ = ~pi0039 & ~new_n7052_;
  assign new_n7054_ = ~new_n7051_ & new_n7053_;
  assign new_n7055_ = ~new_n7042_ & ~new_n7044_;
  assign new_n7056_ = new_n6696_ & ~new_n7055_;
  assign new_n7057_ = pi0039 & new_n7056_;
  assign new_n7058_ = pi0038 & ~new_n7057_;
  assign new_n7059_ = ~new_n7054_ & new_n7058_;
  assign new_n7060_ = ~new_n7049_ & ~new_n7059_;
  assign new_n7061_ = ~pi0100 & ~new_n7060_;
  assign new_n7062_ = pi0969 & new_n6769_;
  assign new_n7063_ = ~pi0299 & ~new_n7062_;
  assign new_n7064_ = pi0963 & new_n6775_;
  assign new_n7065_ = new_n7024_ & ~new_n7064_;
  assign new_n7066_ = new_n3186_ & ~new_n7065_;
  assign new_n7067_ = ~new_n7063_ & new_n7066_;
  assign new_n7068_ = ~new_n3186_ & new_n7056_;
  assign new_n7069_ = pi0100 & ~new_n7068_;
  assign new_n7070_ = ~new_n7067_ & new_n7069_;
  assign new_n7071_ = ~pi0087 & ~new_n7070_;
  assign new_n7072_ = ~new_n7061_ & new_n7071_;
  assign new_n7073_ = pi0087 & new_n7056_;
  assign new_n7074_ = ~pi0075 & ~new_n7073_;
  assign new_n7075_ = ~new_n7072_ & new_n7074_;
  assign new_n7076_ = ~new_n3227_ & new_n7056_;
  assign new_n7077_ = new_n3246_ & new_n7054_;
  assign new_n7078_ = ~new_n7076_ & ~new_n7077_;
  assign new_n7079_ = pi0075 & new_n7078_;
  assign new_n7080_ = ~pi0092 & ~new_n7079_;
  assign new_n7081_ = ~new_n7075_ & new_n7080_;
  assign new_n7082_ = ~pi0075 & new_n7078_;
  assign new_n7083_ = pi0075 & ~new_n7056_;
  assign new_n7084_ = pi0092 & ~new_n7083_;
  assign new_n7085_ = ~new_n7082_ & new_n7084_;
  assign new_n7086_ = ~pi0054 & ~new_n7085_;
  assign new_n7087_ = ~new_n7081_ & new_n7086_;
  assign new_n7088_ = new_n3242_ & new_n7078_;
  assign new_n7089_ = ~new_n3242_ & ~new_n7056_;
  assign new_n7090_ = ~new_n7088_ & ~new_n7089_;
  assign new_n7091_ = pi0054 & ~new_n7090_;
  assign new_n7092_ = ~pi0074 & ~new_n7091_;
  assign new_n7093_ = ~new_n7087_ & new_n7092_;
  assign new_n7094_ = ~pi0054 & new_n7088_;
  assign new_n7095_ = ~new_n6554_ & ~new_n7056_;
  assign new_n7096_ = pi0074 & ~new_n7095_;
  assign new_n7097_ = ~new_n7094_ & new_n7096_;
  assign new_n7098_ = ~pi0055 & ~new_n7097_;
  assign new_n7099_ = ~new_n7093_ & new_n7098_;
  assign new_n7100_ = pi0055 & ~new_n7017_;
  assign new_n7101_ = ~new_n7020_ & new_n7100_;
  assign new_n7102_ = new_n3298_ & ~new_n7101_;
  assign new_n7103_ = ~new_n7099_ & new_n7102_;
  assign new_n7104_ = ~new_n3298_ & new_n7017_;
  assign new_n7105_ = ~pi0059 & ~new_n7104_;
  assign new_n7106_ = ~new_n7103_ & new_n7105_;
  assign new_n7107_ = new_n6304_ & new_n7020_;
  assign new_n7108_ = pi0059 & ~new_n7017_;
  assign new_n7109_ = ~new_n7107_ & new_n7108_;
  assign new_n7110_ = ~pi0057 & ~new_n7109_;
  assign new_n7111_ = ~new_n7106_ & new_n7110_;
  assign po0176 = ~new_n7023_ & ~new_n7111_;
  assign new_n7113_ = pi0975 & new_n6696_;
  assign new_n7114_ = ~pi0228 & pi0975;
  assign new_n7115_ = new_n6203_ & new_n7114_;
  assign new_n7116_ = new_n3273_ & new_n7115_;
  assign new_n7117_ = new_n6305_ & new_n7116_;
  assign new_n7118_ = ~new_n7113_ & ~new_n7117_;
  assign new_n7119_ = pi0057 & ~new_n7118_;
  assign new_n7120_ = pi0299 & ~new_n7113_;
  assign new_n7121_ = new_n6705_ & new_n7114_;
  assign new_n7122_ = new_n7120_ & ~new_n7121_;
  assign new_n7123_ = ~new_n6708_ & ~new_n7122_;
  assign new_n7124_ = new_n6713_ & new_n7114_;
  assign new_n7125_ = ~new_n7113_ & ~new_n7124_;
  assign new_n7126_ = new_n6429_ & ~new_n7125_;
  assign new_n7127_ = ~new_n7123_ & ~new_n7126_;
  assign new_n7128_ = pi0971 & new_n6724_;
  assign new_n7129_ = ~pi0299 & ~new_n7128_;
  assign new_n7130_ = pi0232 & ~new_n7129_;
  assign new_n7131_ = ~new_n7127_ & new_n7130_;
  assign new_n7132_ = pi0971 & new_n6718_;
  assign new_n7133_ = ~pi0299 & ~new_n7132_;
  assign new_n7134_ = ~pi0232 & ~new_n7122_;
  assign new_n7135_ = ~new_n7133_ & new_n7134_;
  assign new_n7136_ = ~new_n7131_ & ~new_n7135_;
  assign new_n7137_ = ~pi0039 & ~new_n7136_;
  assign new_n7138_ = ~pi0299 & pi0971;
  assign new_n7139_ = ~new_n6742_ & new_n7138_;
  assign new_n7140_ = pi0299 & pi0975;
  assign new_n7141_ = ~new_n6738_ & new_n7140_;
  assign new_n7142_ = ~new_n7139_ & ~new_n7141_;
  assign new_n7143_ = new_n6746_ & ~new_n7142_;
  assign new_n7144_ = ~pi0038 & ~new_n7143_;
  assign new_n7145_ = ~new_n7137_ & new_n7144_;
  assign new_n7146_ = pi0971 & new_n6751_;
  assign new_n7147_ = ~pi0299 & ~new_n7146_;
  assign new_n7148_ = ~new_n7115_ & new_n7120_;
  assign new_n7149_ = ~pi0039 & ~new_n7148_;
  assign new_n7150_ = ~new_n7147_ & new_n7149_;
  assign new_n7151_ = ~new_n7138_ & ~new_n7140_;
  assign new_n7152_ = new_n6696_ & ~new_n7151_;
  assign new_n7153_ = pi0039 & new_n7152_;
  assign new_n7154_ = pi0038 & ~new_n7153_;
  assign new_n7155_ = ~new_n7150_ & new_n7154_;
  assign new_n7156_ = ~new_n7145_ & ~new_n7155_;
  assign new_n7157_ = ~pi0100 & ~new_n7156_;
  assign new_n7158_ = pi0971 & new_n6769_;
  assign new_n7159_ = ~pi0299 & ~new_n7158_;
  assign new_n7160_ = pi0975 & new_n6775_;
  assign new_n7161_ = new_n7120_ & ~new_n7160_;
  assign new_n7162_ = new_n3186_ & ~new_n7161_;
  assign new_n7163_ = ~new_n7159_ & new_n7162_;
  assign new_n7164_ = ~new_n3186_ & new_n7152_;
  assign new_n7165_ = pi0100 & ~new_n7164_;
  assign new_n7166_ = ~new_n7163_ & new_n7165_;
  assign new_n7167_ = ~pi0087 & ~new_n7166_;
  assign new_n7168_ = ~new_n7157_ & new_n7167_;
  assign new_n7169_ = pi0087 & new_n7152_;
  assign new_n7170_ = ~pi0075 & ~new_n7169_;
  assign new_n7171_ = ~new_n7168_ & new_n7170_;
  assign new_n7172_ = ~new_n3227_ & new_n7152_;
  assign new_n7173_ = new_n3246_ & new_n7150_;
  assign new_n7174_ = ~new_n7172_ & ~new_n7173_;
  assign new_n7175_ = pi0075 & new_n7174_;
  assign new_n7176_ = ~pi0092 & ~new_n7175_;
  assign new_n7177_ = ~new_n7171_ & new_n7176_;
  assign new_n7178_ = ~pi0075 & new_n7174_;
  assign new_n7179_ = pi0075 & ~new_n7152_;
  assign new_n7180_ = pi0092 & ~new_n7179_;
  assign new_n7181_ = ~new_n7178_ & new_n7180_;
  assign new_n7182_ = ~pi0054 & ~new_n7181_;
  assign new_n7183_ = ~new_n7177_ & new_n7182_;
  assign new_n7184_ = new_n3242_ & new_n7174_;
  assign new_n7185_ = ~new_n3242_ & ~new_n7152_;
  assign new_n7186_ = ~new_n7184_ & ~new_n7185_;
  assign new_n7187_ = pi0054 & ~new_n7186_;
  assign new_n7188_ = ~pi0074 & ~new_n7187_;
  assign new_n7189_ = ~new_n7183_ & new_n7188_;
  assign new_n7190_ = ~pi0054 & new_n7184_;
  assign new_n7191_ = ~new_n6554_ & ~new_n7152_;
  assign new_n7192_ = pi0074 & ~new_n7191_;
  assign new_n7193_ = ~new_n7190_ & new_n7192_;
  assign new_n7194_ = ~pi0055 & ~new_n7193_;
  assign new_n7195_ = ~new_n7189_ & new_n7194_;
  assign new_n7196_ = pi0055 & ~new_n7113_;
  assign new_n7197_ = ~new_n7116_ & new_n7196_;
  assign new_n7198_ = new_n3298_ & ~new_n7197_;
  assign new_n7199_ = ~new_n7195_ & new_n7198_;
  assign new_n7200_ = ~new_n3298_ & new_n7113_;
  assign new_n7201_ = ~pi0059 & ~new_n7200_;
  assign new_n7202_ = ~new_n7199_ & new_n7201_;
  assign new_n7203_ = new_n6304_ & new_n7116_;
  assign new_n7204_ = pi0059 & ~new_n7113_;
  assign new_n7205_ = ~new_n7203_ & new_n7204_;
  assign new_n7206_ = ~pi0057 & ~new_n7205_;
  assign new_n7207_ = ~new_n7202_ & new_n7206_;
  assign po0177 = ~new_n7119_ & ~new_n7207_;
  assign new_n7209_ = pi0978 & new_n6696_;
  assign new_n7210_ = ~pi0228 & pi0978;
  assign new_n7211_ = new_n3273_ & new_n7210_;
  assign new_n7212_ = new_n6203_ & new_n7211_;
  assign new_n7213_ = new_n6305_ & new_n7212_;
  assign new_n7214_ = ~new_n7209_ & ~new_n7213_;
  assign new_n7215_ = pi0057 & ~new_n7214_;
  assign new_n7216_ = ~pi0299 & pi0974;
  assign new_n7217_ = pi0299 & pi0978;
  assign new_n7218_ = ~new_n7216_ & ~new_n7217_;
  assign new_n7219_ = new_n6751_ & ~new_n7218_;
  assign new_n7220_ = ~pi0039 & new_n7219_;
  assign new_n7221_ = new_n6696_ & ~new_n7218_;
  assign new_n7222_ = pi0039 & new_n7221_;
  assign new_n7223_ = pi0038 & ~new_n7222_;
  assign new_n7224_ = ~new_n7220_ & new_n7223_;
  assign new_n7225_ = pi0299 & ~new_n7209_;
  assign new_n7226_ = new_n6705_ & new_n7210_;
  assign new_n7227_ = new_n7225_ & ~new_n7226_;
  assign new_n7228_ = ~new_n6708_ & ~new_n7227_;
  assign new_n7229_ = new_n6713_ & new_n7210_;
  assign new_n7230_ = ~new_n7209_ & ~new_n7229_;
  assign new_n7231_ = new_n6429_ & ~new_n7230_;
  assign new_n7232_ = ~new_n7228_ & ~new_n7231_;
  assign new_n7233_ = pi0974 & new_n6724_;
  assign new_n7234_ = ~pi0299 & ~new_n7233_;
  assign new_n7235_ = pi0232 & ~new_n7234_;
  assign new_n7236_ = ~new_n7232_ & new_n7235_;
  assign new_n7237_ = pi0974 & new_n6718_;
  assign new_n7238_ = ~pi0299 & ~new_n7237_;
  assign new_n7239_ = ~pi0232 & ~new_n7227_;
  assign new_n7240_ = ~new_n7238_ & new_n7239_;
  assign new_n7241_ = ~new_n7236_ & ~new_n7240_;
  assign new_n7242_ = ~pi0039 & ~new_n7241_;
  assign new_n7243_ = ~new_n6742_ & new_n7216_;
  assign new_n7244_ = ~new_n6738_ & new_n7217_;
  assign new_n7245_ = ~new_n7243_ & ~new_n7244_;
  assign new_n7246_ = new_n6746_ & ~new_n7245_;
  assign new_n7247_ = ~pi0038 & ~new_n7246_;
  assign new_n7248_ = ~new_n7242_ & new_n7247_;
  assign new_n7249_ = ~new_n7224_ & ~new_n7248_;
  assign new_n7250_ = ~pi0100 & ~new_n7249_;
  assign new_n7251_ = pi0974 & new_n6769_;
  assign new_n7252_ = ~pi0299 & ~new_n7251_;
  assign new_n7253_ = pi0978 & new_n6775_;
  assign new_n7254_ = new_n7225_ & ~new_n7253_;
  assign new_n7255_ = new_n3186_ & ~new_n7254_;
  assign new_n7256_ = ~new_n7252_ & new_n7255_;
  assign new_n7257_ = ~new_n3186_ & new_n7221_;
  assign new_n7258_ = pi0100 & ~new_n7257_;
  assign new_n7259_ = ~new_n7256_ & new_n7258_;
  assign new_n7260_ = ~pi0087 & ~new_n7259_;
  assign new_n7261_ = ~new_n7250_ & new_n7260_;
  assign new_n7262_ = pi0087 & new_n7221_;
  assign new_n7263_ = ~pi0075 & ~new_n7262_;
  assign new_n7264_ = ~new_n7261_ & new_n7263_;
  assign new_n7265_ = ~pi0228 & ~new_n3227_;
  assign new_n7266_ = new_n7219_ & ~new_n7265_;
  assign new_n7267_ = pi0075 & ~new_n7266_;
  assign new_n7268_ = ~pi0092 & ~new_n7267_;
  assign new_n7269_ = ~new_n7264_ & new_n7268_;
  assign new_n7270_ = ~pi0075 & ~new_n7266_;
  assign new_n7271_ = pi0075 & ~new_n7221_;
  assign new_n7272_ = pi0092 & ~new_n7271_;
  assign new_n7273_ = ~new_n7270_ & new_n7272_;
  assign new_n7274_ = ~pi0054 & ~new_n7273_;
  assign new_n7275_ = ~new_n7269_ & new_n7274_;
  assign new_n7276_ = new_n3242_ & ~new_n7266_;
  assign new_n7277_ = ~new_n3242_ & ~new_n7221_;
  assign new_n7278_ = ~new_n7276_ & ~new_n7277_;
  assign new_n7279_ = pi0054 & ~new_n7278_;
  assign new_n7280_ = ~pi0074 & ~new_n7279_;
  assign new_n7281_ = ~new_n7275_ & new_n7280_;
  assign new_n7282_ = ~pi0054 & new_n7276_;
  assign new_n7283_ = ~new_n6554_ & ~new_n7221_;
  assign new_n7284_ = pi0074 & ~new_n7283_;
  assign new_n7285_ = ~new_n7282_ & new_n7284_;
  assign new_n7286_ = ~pi0055 & ~new_n7285_;
  assign new_n7287_ = ~new_n7281_ & new_n7286_;
  assign new_n7288_ = pi0055 & ~new_n7209_;
  assign new_n7289_ = ~new_n7212_ & new_n7288_;
  assign new_n7290_ = new_n3298_ & ~new_n7289_;
  assign new_n7291_ = ~new_n7287_ & new_n7290_;
  assign new_n7292_ = ~new_n3298_ & new_n7209_;
  assign new_n7293_ = ~pi0059 & ~new_n7292_;
  assign new_n7294_ = ~new_n7291_ & new_n7293_;
  assign new_n7295_ = new_n6304_ & new_n7212_;
  assign new_n7296_ = pi0059 & ~new_n7209_;
  assign new_n7297_ = ~new_n7295_ & new_n7296_;
  assign new_n7298_ = ~pi0057 & ~new_n7297_;
  assign new_n7299_ = ~new_n7294_ & new_n7298_;
  assign po0178 = ~new_n7215_ & ~new_n7299_;
  assign new_n7301_ = new_n3246_ & new_n6257_;
  assign new_n7302_ = pi0075 & ~new_n7301_;
  assign new_n7303_ = new_n3211_ & new_n3235_;
  assign new_n7304_ = new_n6257_ & new_n7303_;
  assign new_n7305_ = pi0092 & ~new_n7304_;
  assign new_n7306_ = ~new_n7302_ & ~new_n7305_;
  assign new_n7307_ = pi0299 & ~new_n6223_;
  assign new_n7308_ = new_n6736_ & new_n7307_;
  assign new_n7309_ = ~pi0299 & ~new_n6244_;
  assign new_n7310_ = new_n6483_ & new_n7309_;
  assign new_n7311_ = pi0039 & ~new_n7310_;
  assign new_n7312_ = ~new_n7308_ & new_n7311_;
  assign new_n7313_ = ~new_n6434_ & new_n6708_;
  assign new_n7314_ = ~new_n6712_ & new_n7313_;
  assign new_n7315_ = new_n6396_ & new_n6420_;
  assign new_n7316_ = ~pi0299 & ~new_n6400_;
  assign new_n7317_ = ~new_n6721_ & new_n7316_;
  assign new_n7318_ = ~new_n7315_ & new_n7317_;
  assign new_n7319_ = pi0299 & new_n6433_;
  assign new_n7320_ = ~new_n6429_ & new_n7319_;
  assign new_n7321_ = pi0232 & ~new_n7320_;
  assign new_n7322_ = ~new_n7318_ & new_n7321_;
  assign new_n7323_ = ~new_n7314_ & new_n7322_;
  assign new_n7324_ = ~pi0299 & new_n6389_;
  assign new_n7325_ = ~pi0232 & ~new_n7319_;
  assign new_n7326_ = ~new_n7324_ & new_n7325_;
  assign new_n7327_ = ~pi0039 & ~new_n7326_;
  assign new_n7328_ = ~new_n7323_ & new_n7327_;
  assign new_n7329_ = ~new_n7312_ & ~new_n7328_;
  assign new_n7330_ = ~pi0038 & ~new_n7329_;
  assign new_n7331_ = ~new_n6133_ & ~new_n7330_;
  assign new_n7332_ = ~pi0100 & ~new_n7331_;
  assign new_n7333_ = ~pi0038 & new_n6257_;
  assign new_n7334_ = pi0100 & ~new_n7333_;
  assign new_n7335_ = new_n6286_ & ~new_n7334_;
  assign new_n7336_ = ~new_n7332_ & new_n7335_;
  assign new_n7337_ = new_n3242_ & ~new_n7336_;
  assign new_n7338_ = new_n7306_ & ~new_n7337_;
  assign new_n7339_ = ~pi0054 & ~new_n7338_;
  assign new_n7340_ = ~pi0092 & new_n7304_;
  assign new_n7341_ = pi0054 & ~new_n7340_;
  assign new_n7342_ = ~new_n7339_ & ~new_n7341_;
  assign new_n7343_ = ~pi0074 & ~new_n7342_;
  assign new_n7344_ = ~new_n6130_ & ~new_n7343_;
  assign new_n7345_ = ~pi0055 & ~new_n7344_;
  assign new_n7346_ = new_n3283_ & new_n6125_;
  assign new_n7347_ = pi0055 & ~new_n7346_;
  assign new_n7348_ = ~pi0056 & ~new_n7347_;
  assign new_n7349_ = ~pi0062 & new_n7348_;
  assign new_n7350_ = ~new_n7345_ & new_n7349_;
  assign new_n7351_ = new_n3436_ & ~new_n7350_;
  assign po0195 = new_n6123_ & ~new_n7351_;
  assign new_n7353_ = ~pi0954 & ~po0195;
  assign new_n7354_ = pi0024 & pi0954;
  assign po0182 = ~new_n7353_ & ~new_n7354_;
  assign new_n7356_ = new_n3281_ & new_n3326_;
  assign new_n7357_ = new_n3437_ & new_n7356_;
  assign new_n7358_ = ~new_n3131_ & ~new_n7357_;
  assign new_n7359_ = pi0062 & ~new_n7358_;
  assign new_n7360_ = ~pi0100 & new_n4686_;
  assign new_n7361_ = new_n3100_ & ~new_n6507_;
  assign new_n7362_ = ~pi0299 & ~new_n7361_;
  assign new_n7363_ = pi0299 & ~new_n3395_;
  assign new_n7364_ = ~new_n7362_ & ~new_n7363_;
  assign new_n7365_ = pi0100 & new_n3326_;
  assign new_n7366_ = new_n7364_ & new_n7365_;
  assign new_n7367_ = ~pi0039 & ~new_n7366_;
  assign new_n7368_ = ~new_n7360_ & new_n7367_;
  assign new_n7369_ = ~pi0100 & new_n3326_;
  assign new_n7370_ = pi0039 & ~new_n7369_;
  assign new_n7371_ = ~pi0038 & ~new_n7370_;
  assign new_n7372_ = ~new_n7368_ & new_n7371_;
  assign new_n7373_ = ~new_n3131_ & ~new_n7372_;
  assign new_n7374_ = ~pi0087 & ~new_n7373_;
  assign new_n7375_ = ~new_n3131_ & ~new_n7356_;
  assign new_n7376_ = pi0087 & ~new_n7375_;
  assign new_n7377_ = ~pi0075 & ~new_n7376_;
  assign new_n7378_ = ~new_n7374_ & new_n7377_;
  assign new_n7379_ = pi0075 & ~new_n3131_;
  assign new_n7380_ = ~pi0092 & ~new_n7379_;
  assign new_n7381_ = ~new_n7378_ & new_n7380_;
  assign new_n7382_ = new_n3326_ & new_n3413_;
  assign new_n7383_ = ~new_n3131_ & ~new_n7382_;
  assign new_n7384_ = pi0092 & ~new_n7383_;
  assign new_n7385_ = new_n3270_ & ~new_n7384_;
  assign new_n7386_ = ~new_n7381_ & new_n7385_;
  assign new_n7387_ = ~new_n3131_ & ~new_n3270_;
  assign new_n7388_ = ~pi0055 & ~new_n7387_;
  assign new_n7389_ = ~new_n7386_ & new_n7388_;
  assign new_n7390_ = new_n3281_ & new_n6128_;
  assign new_n7391_ = new_n3326_ & new_n7390_;
  assign new_n7392_ = ~pi0074 & new_n7391_;
  assign new_n7393_ = ~new_n3131_ & ~new_n7392_;
  assign new_n7394_ = pi0055 & ~new_n7393_;
  assign new_n7395_ = ~pi0056 & ~new_n7394_;
  assign new_n7396_ = ~new_n7389_ & new_n7395_;
  assign new_n7397_ = new_n3285_ & new_n3326_;
  assign new_n7398_ = pi0056 & ~new_n3131_;
  assign new_n7399_ = ~new_n7397_ & new_n7398_;
  assign new_n7400_ = ~pi0062 & ~new_n7399_;
  assign new_n7401_ = ~new_n7396_ & new_n7400_;
  assign new_n7402_ = ~new_n7359_ & ~new_n7401_;
  assign new_n7403_ = new_n3436_ & ~new_n7402_;
  assign new_n7404_ = new_n3131_ & ~new_n3436_;
  assign po0183 = new_n7403_ | new_n7404_;
  assign new_n7406_ = pi0119 & pi1056;
  assign new_n7407_ = ~pi0228 & pi0252;
  assign new_n7408_ = ~pi0119 & ~new_n7407_;
  assign new_n7409_ = ~pi0468 & ~new_n7408_;
  assign po0184 = new_n7406_ | ~new_n7409_;
  assign new_n7411_ = pi0119 & pi1077;
  assign po0185 = ~new_n7409_ | new_n7411_;
  assign new_n7413_ = pi0119 & pi1073;
  assign po0186 = ~new_n7409_ | new_n7413_;
  assign new_n7415_ = pi0119 & pi1041;
  assign po0187 = ~new_n7409_ | new_n7415_;
  assign new_n7417_ = pi0360 & ~pi0462;
  assign new_n7418_ = ~pi0360 & pi0462;
  assign new_n7419_ = ~new_n7417_ & ~new_n7418_;
  assign new_n7420_ = pi0352 & ~pi0353;
  assign new_n7421_ = ~pi0352 & pi0353;
  assign new_n7422_ = ~new_n7420_ & ~new_n7421_;
  assign new_n7423_ = new_n7419_ & new_n7422_;
  assign new_n7424_ = ~new_n7419_ & ~new_n7422_;
  assign new_n7425_ = ~new_n7423_ & ~new_n7424_;
  assign new_n7426_ = pi0354 & ~new_n7425_;
  assign new_n7427_ = ~pi0354 & new_n7425_;
  assign new_n7428_ = ~new_n7426_ & ~new_n7427_;
  assign new_n7429_ = pi0351 & pi1199;
  assign new_n7430_ = pi0345 & ~pi0346;
  assign new_n7431_ = ~pi0345 & pi0346;
  assign new_n7432_ = ~new_n7430_ & ~new_n7431_;
  assign new_n7433_ = pi0323 & ~new_n7432_;
  assign new_n7434_ = ~pi0323 & new_n7432_;
  assign new_n7435_ = ~new_n7433_ & ~new_n7434_;
  assign new_n7436_ = pi0358 & ~pi0450;
  assign new_n7437_ = ~pi0358 & pi0450;
  assign new_n7438_ = ~new_n7436_ & ~new_n7437_;
  assign new_n7439_ = new_n7435_ & ~new_n7438_;
  assign new_n7440_ = ~new_n7435_ & new_n7438_;
  assign new_n7441_ = ~new_n7439_ & ~new_n7440_;
  assign new_n7442_ = ~pi0327 & ~pi0362;
  assign new_n7443_ = pi0327 & pi0362;
  assign new_n7444_ = ~new_n7442_ & ~new_n7443_;
  assign new_n7445_ = pi0343 & ~pi0344;
  assign new_n7446_ = ~pi0343 & pi0344;
  assign new_n7447_ = ~new_n7445_ & ~new_n7446_;
  assign new_n7448_ = new_n7444_ & ~new_n7447_;
  assign new_n7449_ = ~new_n7444_ & new_n7447_;
  assign new_n7450_ = ~new_n7448_ & ~new_n7449_;
  assign new_n7451_ = ~new_n7441_ & ~new_n7450_;
  assign new_n7452_ = new_n7441_ & new_n7450_;
  assign new_n7453_ = pi1197 & ~new_n7452_;
  assign new_n7454_ = ~new_n7451_ & new_n7453_;
  assign new_n7455_ = ~pi0074 & new_n6290_;
  assign new_n7456_ = ~pi0122 & pi0829;
  assign new_n7457_ = new_n2534_ & ~new_n6154_;
  assign new_n7458_ = ~pi0841 & new_n2492_;
  assign new_n7459_ = pi0090 & new_n7458_;
  assign new_n7460_ = ~pi0093 & ~new_n7459_;
  assign new_n7461_ = new_n7457_ & ~new_n7460_;
  assign new_n7462_ = ~pi0051 & ~new_n7461_;
  assign new_n7463_ = ~pi0050 & ~pi0077;
  assign new_n7464_ = ~pi0094 & new_n7463_;
  assign new_n7465_ = new_n2576_ & new_n7464_;
  assign new_n7466_ = ~pi0088 & pi0098;
  assign new_n7467_ = new_n2484_ & new_n7466_;
  assign new_n7468_ = new_n7465_ & new_n7467_;
  assign new_n7469_ = ~pi0097 & ~new_n7468_;
  assign new_n7470_ = new_n2514_ & ~new_n7469_;
  assign new_n7471_ = ~pi0035 & new_n2493_;
  assign new_n7472_ = ~pi0070 & new_n7471_;
  assign new_n7473_ = new_n7470_ & new_n7472_;
  assign new_n7474_ = new_n7462_ & ~new_n7473_;
  assign new_n7475_ = ~new_n2558_ & ~new_n7474_;
  assign new_n7476_ = ~pi0096 & new_n3098_;
  assign new_n7477_ = new_n7475_ & new_n7476_;
  assign new_n7478_ = new_n6277_ & new_n7477_;
  assign new_n7479_ = ~new_n7456_ & new_n7478_;
  assign new_n7480_ = ~pi0096 & ~new_n7475_;
  assign new_n7481_ = pi0096 & ~new_n6384_;
  assign new_n7482_ = new_n3098_ & ~new_n7481_;
  assign new_n7483_ = new_n2799_ & new_n7456_;
  assign new_n7484_ = new_n7482_ & new_n7483_;
  assign new_n7485_ = ~new_n7480_ & new_n7484_;
  assign new_n7486_ = ~new_n7479_ & ~new_n7485_;
  assign new_n7487_ = ~pi1093 & ~new_n7486_;
  assign new_n7488_ = ~pi0087 & ~new_n7487_;
  assign new_n7489_ = new_n3100_ & po0740;
  assign new_n7490_ = pi0087 & ~new_n7489_;
  assign new_n7491_ = ~pi0075 & new_n3281_;
  assign new_n7492_ = ~new_n7490_ & new_n7491_;
  assign new_n7493_ = ~new_n7488_ & new_n7492_;
  assign new_n7494_ = ~pi0567 & ~new_n7493_;
  assign new_n7495_ = new_n7455_ & ~new_n7494_;
  assign new_n7496_ = ~pi0299 & ~new_n3068_;
  assign new_n7497_ = pi0299 & ~new_n2448_;
  assign new_n7498_ = ~new_n7496_ & ~new_n7497_;
  assign new_n7499_ = pi0232 & new_n6185_;
  assign new_n7500_ = new_n7498_ & new_n7499_;
  assign new_n7501_ = new_n3227_ & ~new_n7500_;
  assign new_n7502_ = ~pi0024 & new_n6510_;
  assign new_n7503_ = ~new_n2732_ & po1057;
  assign new_n7504_ = pi1091 & new_n7503_;
  assign new_n7505_ = new_n7483_ & new_n7504_;
  assign new_n7506_ = new_n7502_ & new_n7505_;
  assign new_n7507_ = pi1093 & new_n7506_;
  assign new_n7508_ = new_n7501_ & new_n7507_;
  assign new_n7509_ = pi0075 & ~new_n7508_;
  assign new_n7510_ = pi1093 & ~new_n2732_;
  assign new_n7511_ = pi0824 & new_n2799_;
  assign new_n7512_ = ~new_n2558_ & new_n7476_;
  assign new_n7513_ = ~new_n7462_ & new_n7512_;
  assign new_n7514_ = new_n7511_ & new_n7513_;
  assign new_n7515_ = ~pi0829 & new_n7514_;
  assign new_n7516_ = ~pi0024 & new_n2565_;
  assign new_n7517_ = ~pi0046 & pi0097;
  assign new_n7518_ = ~pi0108 & new_n7517_;
  assign new_n7519_ = new_n6401_ & new_n7518_;
  assign new_n7520_ = new_n2581_ & new_n7519_;
  assign new_n7521_ = ~pi0091 & new_n7520_;
  assign new_n7522_ = ~new_n7516_ & ~new_n7521_;
  assign new_n7523_ = new_n2518_ & new_n7457_;
  assign new_n7524_ = ~new_n7522_ & new_n7523_;
  assign new_n7525_ = new_n7462_ & ~new_n7524_;
  assign new_n7526_ = ~new_n2558_ & ~new_n7525_;
  assign new_n7527_ = ~pi0096 & ~new_n7526_;
  assign new_n7528_ = new_n2800_ & new_n7482_;
  assign new_n7529_ = ~new_n7527_ & new_n7528_;
  assign new_n7530_ = ~new_n7515_ & ~new_n7529_;
  assign new_n7531_ = ~pi0122 & ~new_n7530_;
  assign new_n7532_ = pi0122 & new_n6277_;
  assign new_n7533_ = new_n7513_ & new_n7532_;
  assign new_n7534_ = ~new_n7531_ & ~new_n7533_;
  assign new_n7535_ = new_n7510_ & ~new_n7534_;
  assign new_n7536_ = pi1091 & ~new_n7535_;
  assign new_n7537_ = ~new_n7487_ & new_n7536_;
  assign new_n7538_ = ~pi1091 & ~new_n7487_;
  assign new_n7539_ = ~new_n7537_ & ~new_n7538_;
  assign new_n7540_ = ~pi0039 & ~new_n7539_;
  assign new_n7541_ = ~new_n2732_ & new_n2753_;
  assign new_n7542_ = new_n6456_ & new_n7541_;
  assign new_n7543_ = new_n2754_ & new_n7542_;
  assign new_n7544_ = pi1091 & new_n7543_;
  assign new_n7545_ = ~new_n6244_ & new_n7544_;
  assign new_n7546_ = ~pi0299 & new_n6480_;
  assign new_n7547_ = ~pi0224 & new_n7546_;
  assign new_n7548_ = new_n7545_ & new_n7547_;
  assign new_n7549_ = ~new_n6223_ & new_n7544_;
  assign new_n7550_ = ~pi0216 & new_n6605_;
  assign new_n7551_ = new_n7549_ & new_n7550_;
  assign new_n7552_ = pi0039 & ~new_n7551_;
  assign new_n7553_ = ~new_n7548_ & new_n7552_;
  assign new_n7554_ = ~pi0038 & ~new_n7553_;
  assign new_n7555_ = ~new_n7540_ & new_n7554_;
  assign new_n7556_ = ~pi0100 & ~new_n7555_;
  assign new_n7557_ = new_n6458_ & new_n7513_;
  assign new_n7558_ = new_n7554_ & new_n7557_;
  assign new_n7559_ = ~new_n7536_ & new_n7558_;
  assign new_n7560_ = new_n7556_ & ~new_n7559_;
  assign new_n7561_ = pi1093 & new_n7483_;
  assign new_n7562_ = new_n7503_ & new_n7561_;
  assign new_n7563_ = new_n3100_ & new_n7562_;
  assign new_n7564_ = pi1091 & new_n7563_;
  assign new_n7565_ = pi0228 & new_n7564_;
  assign new_n7566_ = new_n3186_ & ~new_n7500_;
  assign new_n7567_ = new_n7565_ & new_n7566_;
  assign new_n7568_ = pi0100 & ~new_n7567_;
  assign new_n7569_ = ~new_n7560_ & ~new_n7568_;
  assign new_n7570_ = ~pi0087 & ~new_n7569_;
  assign new_n7571_ = new_n3100_ & new_n7511_;
  assign new_n7572_ = ~pi1091 & pi1093;
  assign new_n7573_ = ~new_n7571_ & new_n7572_;
  assign new_n7574_ = pi1093 & new_n2732_;
  assign new_n7575_ = new_n6277_ & ~new_n7574_;
  assign new_n7576_ = new_n3100_ & new_n7575_;
  assign new_n7577_ = ~new_n7572_ & ~new_n7576_;
  assign new_n7578_ = new_n3212_ & ~new_n7577_;
  assign new_n7579_ = ~new_n7573_ & new_n7578_;
  assign new_n7580_ = pi0087 & ~new_n7579_;
  assign new_n7581_ = ~new_n7570_ & ~new_n7580_;
  assign new_n7582_ = ~pi0075 & ~new_n7581_;
  assign new_n7583_ = ~new_n7509_ & ~new_n7582_;
  assign new_n7584_ = pi0567 & ~new_n7583_;
  assign new_n7585_ = new_n7495_ & ~new_n7584_;
  assign new_n7586_ = pi0350 & ~pi0592;
  assign new_n7587_ = ~new_n7585_ & ~new_n7586_;
  assign new_n7588_ = pi0321 & ~pi0347;
  assign new_n7589_ = ~pi0321 & pi0347;
  assign new_n7590_ = ~new_n7588_ & ~new_n7589_;
  assign new_n7591_ = pi0316 & ~pi0349;
  assign new_n7592_ = ~pi0316 & pi0349;
  assign new_n7593_ = ~new_n7591_ & ~new_n7592_;
  assign new_n7594_ = pi0348 & new_n7593_;
  assign new_n7595_ = ~pi0348 & ~new_n7593_;
  assign new_n7596_ = ~new_n7594_ & ~new_n7595_;
  assign new_n7597_ = pi0315 & ~pi0359;
  assign new_n7598_ = ~pi0315 & pi0359;
  assign new_n7599_ = ~new_n7597_ & ~new_n7598_;
  assign new_n7600_ = pi0322 & new_n7599_;
  assign new_n7601_ = ~pi0322 & ~new_n7599_;
  assign new_n7602_ = ~new_n7600_ & ~new_n7601_;
  assign new_n7603_ = new_n7596_ & ~new_n7602_;
  assign new_n7604_ = ~new_n7596_ & new_n7602_;
  assign new_n7605_ = ~new_n7603_ & ~new_n7604_;
  assign new_n7606_ = new_n7590_ & new_n7605_;
  assign new_n7607_ = ~new_n7590_ & ~new_n7605_;
  assign new_n7608_ = ~new_n7606_ & ~new_n7607_;
  assign new_n7609_ = ~pi0087 & ~new_n7568_;
  assign new_n7610_ = ~new_n7556_ & new_n7609_;
  assign new_n7611_ = ~pi1091 & ~new_n7489_;
  assign new_n7612_ = pi1091 & ~new_n7576_;
  assign new_n7613_ = pi0087 & ~pi0100;
  assign new_n7614_ = new_n3186_ & new_n7613_;
  assign new_n7615_ = ~new_n7612_ & new_n7614_;
  assign new_n7616_ = ~new_n7611_ & new_n7615_;
  assign new_n7617_ = ~pi0075 & ~new_n7616_;
  assign new_n7618_ = ~new_n7610_ & new_n7617_;
  assign new_n7619_ = ~new_n7509_ & ~new_n7618_;
  assign new_n7620_ = pi0567 & ~new_n7619_;
  assign new_n7621_ = new_n7495_ & ~new_n7620_;
  assign new_n7622_ = new_n7586_ & ~new_n7621_;
  assign new_n7623_ = ~new_n7608_ & ~new_n7622_;
  assign new_n7624_ = ~new_n7587_ & new_n7623_;
  assign new_n7625_ = pi0452 & ~pi0455;
  assign new_n7626_ = ~pi0452 & pi0455;
  assign new_n7627_ = ~new_n7625_ & ~new_n7626_;
  assign new_n7628_ = pi0355 & new_n7627_;
  assign new_n7629_ = ~pi0355 & ~new_n7627_;
  assign new_n7630_ = ~new_n7628_ & ~new_n7629_;
  assign new_n7631_ = pi0320 & ~pi0460;
  assign new_n7632_ = ~pi0320 & pi0460;
  assign new_n7633_ = ~new_n7631_ & ~new_n7632_;
  assign new_n7634_ = pi0342 & ~new_n7633_;
  assign new_n7635_ = ~pi0342 & new_n7633_;
  assign new_n7636_ = ~new_n7634_ & ~new_n7635_;
  assign new_n7637_ = pi0361 & ~pi0441;
  assign new_n7638_ = ~pi0361 & pi0441;
  assign new_n7639_ = ~new_n7637_ & ~new_n7638_;
  assign new_n7640_ = new_n7636_ & new_n7639_;
  assign new_n7641_ = ~new_n7636_ & ~new_n7639_;
  assign new_n7642_ = ~new_n7640_ & ~new_n7641_;
  assign new_n7643_ = pi0458 & new_n7642_;
  assign new_n7644_ = ~pi0458 & ~new_n7642_;
  assign new_n7645_ = ~new_n7643_ & ~new_n7644_;
  assign new_n7646_ = new_n7630_ & new_n7645_;
  assign new_n7647_ = ~new_n7630_ & ~new_n7645_;
  assign new_n7648_ = ~new_n7646_ & ~new_n7647_;
  assign new_n7649_ = pi1196 & new_n7648_;
  assign new_n7650_ = ~pi0350 & ~pi0592;
  assign new_n7651_ = ~new_n7585_ & ~new_n7650_;
  assign new_n7652_ = ~new_n7621_ & new_n7650_;
  assign new_n7653_ = new_n7608_ & ~new_n7652_;
  assign new_n7654_ = ~new_n7651_ & new_n7653_;
  assign new_n7655_ = ~new_n7649_ & ~new_n7654_;
  assign new_n7656_ = ~new_n7624_ & new_n7655_;
  assign new_n7657_ = ~pi0592 & ~new_n7621_;
  assign new_n7658_ = pi0592 & ~new_n7585_;
  assign new_n7659_ = ~new_n7657_ & ~new_n7658_;
  assign new_n7660_ = new_n7649_ & ~new_n7659_;
  assign new_n7661_ = pi1198 & ~new_n7660_;
  assign new_n7662_ = ~new_n7656_ & new_n7661_;
  assign new_n7663_ = ~pi0455 & ~new_n7659_;
  assign new_n7664_ = pi0455 & ~new_n7585_;
  assign new_n7665_ = ~new_n7663_ & ~new_n7664_;
  assign new_n7666_ = ~pi0452 & ~new_n7665_;
  assign new_n7667_ = pi0455 & ~new_n7659_;
  assign new_n7668_ = ~pi0455 & ~new_n7585_;
  assign new_n7669_ = ~new_n7667_ & ~new_n7668_;
  assign new_n7670_ = pi0452 & ~new_n7669_;
  assign new_n7671_ = ~new_n7666_ & ~new_n7670_;
  assign new_n7672_ = ~pi0355 & ~new_n7671_;
  assign new_n7673_ = ~pi0452 & ~new_n7669_;
  assign new_n7674_ = pi0452 & ~new_n7665_;
  assign new_n7675_ = ~new_n7673_ & ~new_n7674_;
  assign new_n7676_ = pi0355 & ~new_n7675_;
  assign new_n7677_ = ~new_n7672_ & ~new_n7676_;
  assign new_n7678_ = ~pi0458 & ~new_n7677_;
  assign new_n7679_ = ~pi0355 & ~new_n7675_;
  assign new_n7680_ = pi0355 & ~new_n7671_;
  assign new_n7681_ = ~new_n7679_ & ~new_n7680_;
  assign new_n7682_ = pi0458 & ~new_n7681_;
  assign new_n7683_ = ~new_n7642_ & ~new_n7682_;
  assign new_n7684_ = ~new_n7678_ & new_n7683_;
  assign new_n7685_ = ~pi0458 & ~new_n7681_;
  assign new_n7686_ = pi0458 & ~new_n7677_;
  assign new_n7687_ = new_n7642_ & ~new_n7686_;
  assign new_n7688_ = ~new_n7685_ & new_n7687_;
  assign new_n7689_ = pi1196 & ~new_n7688_;
  assign new_n7690_ = ~new_n7684_ & new_n7689_;
  assign new_n7691_ = ~pi1196 & ~new_n7585_;
  assign new_n7692_ = ~pi1198 & ~new_n7691_;
  assign new_n7693_ = ~new_n7690_ & new_n7692_;
  assign new_n7694_ = ~new_n7662_ & ~new_n7693_;
  assign new_n7695_ = ~new_n7454_ & ~new_n7694_;
  assign new_n7696_ = new_n7454_ & new_n7659_;
  assign new_n7697_ = ~new_n7695_ & ~new_n7696_;
  assign new_n7698_ = ~new_n7429_ & new_n7697_;
  assign new_n7699_ = pi1199 & ~new_n7659_;
  assign new_n7700_ = pi0351 & new_n7699_;
  assign new_n7701_ = ~new_n7698_ & ~new_n7700_;
  assign new_n7702_ = ~pi0461 & ~new_n7701_;
  assign new_n7703_ = ~pi0351 & pi1199;
  assign new_n7704_ = new_n7697_ & ~new_n7703_;
  assign new_n7705_ = ~pi0351 & new_n7699_;
  assign new_n7706_ = ~new_n7704_ & ~new_n7705_;
  assign new_n7707_ = pi0461 & ~new_n7706_;
  assign new_n7708_ = ~new_n7702_ & ~new_n7707_;
  assign new_n7709_ = ~pi0357 & ~new_n7708_;
  assign new_n7710_ = ~pi0461 & ~new_n7706_;
  assign new_n7711_ = pi0461 & ~new_n7701_;
  assign new_n7712_ = ~new_n7710_ & ~new_n7711_;
  assign new_n7713_ = pi0357 & ~new_n7712_;
  assign new_n7714_ = ~new_n7709_ & ~new_n7713_;
  assign new_n7715_ = ~pi0356 & ~new_n7714_;
  assign new_n7716_ = ~pi0357 & ~new_n7712_;
  assign new_n7717_ = pi0357 & ~new_n7708_;
  assign new_n7718_ = ~new_n7716_ & ~new_n7717_;
  assign new_n7719_ = pi0356 & ~new_n7718_;
  assign new_n7720_ = ~new_n7715_ & ~new_n7719_;
  assign new_n7721_ = new_n7428_ & ~new_n7720_;
  assign new_n7722_ = ~pi0356 & ~new_n7718_;
  assign new_n7723_ = pi0356 & ~new_n7714_;
  assign new_n7724_ = ~new_n7722_ & ~new_n7723_;
  assign new_n7725_ = ~new_n7428_ & ~new_n7724_;
  assign new_n7726_ = ~pi0591 & ~new_n7725_;
  assign new_n7727_ = ~new_n7721_ & new_n7726_;
  assign new_n7728_ = pi0591 & new_n7585_;
  assign new_n7729_ = pi0590 & ~new_n7728_;
  assign new_n7730_ = ~new_n7727_ & new_n7729_;
  assign new_n7731_ = ~pi0285 & ~pi0286;
  assign new_n7732_ = ~pi0289 & new_n7731_;
  assign new_n7733_ = ~pi0288 & new_n7732_;
  assign new_n7734_ = ~pi0363 & ~pi0372;
  assign new_n7735_ = pi0363 & pi0372;
  assign new_n7736_ = ~new_n7734_ & ~new_n7735_;
  assign new_n7737_ = pi0386 & ~new_n7736_;
  assign new_n7738_ = ~pi0386 & new_n7736_;
  assign new_n7739_ = ~new_n7737_ & ~new_n7738_;
  assign new_n7740_ = pi0338 & ~pi0388;
  assign new_n7741_ = ~pi0338 & pi0388;
  assign new_n7742_ = ~new_n7740_ & ~new_n7741_;
  assign new_n7743_ = pi0337 & ~pi0339;
  assign new_n7744_ = ~pi0337 & pi0339;
  assign new_n7745_ = ~new_n7743_ & ~new_n7744_;
  assign new_n7746_ = pi0387 & new_n7745_;
  assign new_n7747_ = ~pi0387 & ~new_n7745_;
  assign new_n7748_ = ~new_n7746_ & ~new_n7747_;
  assign new_n7749_ = pi0380 & ~new_n7748_;
  assign new_n7750_ = ~pi0380 & new_n7748_;
  assign new_n7751_ = ~new_n7749_ & ~new_n7750_;
  assign new_n7752_ = new_n7742_ & ~new_n7751_;
  assign new_n7753_ = ~new_n7742_ & new_n7751_;
  assign new_n7754_ = ~new_n7752_ & ~new_n7753_;
  assign new_n7755_ = new_n7739_ & new_n7754_;
  assign new_n7756_ = ~new_n7739_ & ~new_n7754_;
  assign new_n7757_ = ~new_n7755_ & ~new_n7756_;
  assign new_n7758_ = pi1196 & ~new_n7757_;
  assign new_n7759_ = ~pi0368 & ~pi0389;
  assign new_n7760_ = pi0368 & pi0389;
  assign new_n7761_ = ~new_n7759_ & ~new_n7760_;
  assign new_n7762_ = pi0365 & ~pi0447;
  assign new_n7763_ = ~pi0365 & pi0447;
  assign new_n7764_ = ~new_n7762_ & ~new_n7763_;
  assign new_n7765_ = pi0336 & ~pi0383;
  assign new_n7766_ = ~pi0336 & pi0383;
  assign new_n7767_ = ~new_n7765_ & ~new_n7766_;
  assign new_n7768_ = pi0364 & ~pi0366;
  assign new_n7769_ = ~pi0364 & pi0366;
  assign new_n7770_ = ~new_n7768_ & ~new_n7769_;
  assign new_n7771_ = new_n7767_ & new_n7770_;
  assign new_n7772_ = ~new_n7767_ & ~new_n7770_;
  assign new_n7773_ = ~new_n7771_ & ~new_n7772_;
  assign new_n7774_ = new_n7764_ & new_n7773_;
  assign new_n7775_ = ~new_n7764_ & ~new_n7773_;
  assign new_n7776_ = ~new_n7774_ & ~new_n7775_;
  assign new_n7777_ = pi0367 & ~new_n7776_;
  assign new_n7778_ = ~pi0367 & new_n7776_;
  assign new_n7779_ = ~new_n7777_ & ~new_n7778_;
  assign new_n7780_ = ~new_n7761_ & ~new_n7779_;
  assign new_n7781_ = new_n7761_ & new_n7779_;
  assign new_n7782_ = pi1197 & ~new_n7781_;
  assign new_n7783_ = ~new_n7780_ & new_n7782_;
  assign new_n7784_ = ~new_n7758_ & ~new_n7783_;
  assign new_n7785_ = pi0377 & pi0592;
  assign new_n7786_ = ~new_n7585_ & ~new_n7785_;
  assign new_n7787_ = pi0379 & ~pi0382;
  assign new_n7788_ = ~pi0379 & pi0382;
  assign new_n7789_ = ~new_n7787_ & ~new_n7788_;
  assign new_n7790_ = pi0376 & ~pi0439;
  assign new_n7791_ = ~pi0376 & pi0439;
  assign new_n7792_ = ~new_n7790_ & ~new_n7791_;
  assign new_n7793_ = pi0381 & new_n7792_;
  assign new_n7794_ = ~pi0381 & ~new_n7792_;
  assign new_n7795_ = ~new_n7793_ & ~new_n7794_;
  assign new_n7796_ = pi0317 & ~pi0385;
  assign new_n7797_ = ~pi0317 & pi0385;
  assign new_n7798_ = ~new_n7796_ & ~new_n7797_;
  assign new_n7799_ = pi0378 & new_n7798_;
  assign new_n7800_ = ~pi0378 & ~new_n7798_;
  assign new_n7801_ = ~new_n7799_ & ~new_n7800_;
  assign new_n7802_ = new_n7795_ & ~new_n7801_;
  assign new_n7803_ = ~new_n7795_ & new_n7801_;
  assign new_n7804_ = ~new_n7802_ & ~new_n7803_;
  assign new_n7805_ = new_n7789_ & new_n7804_;
  assign new_n7806_ = ~new_n7789_ & ~new_n7804_;
  assign new_n7807_ = ~new_n7805_ & ~new_n7806_;
  assign new_n7808_ = ~new_n7621_ & new_n7785_;
  assign new_n7809_ = ~new_n7807_ & ~new_n7808_;
  assign new_n7810_ = ~new_n7786_ & new_n7809_;
  assign new_n7811_ = ~pi0377 & pi0592;
  assign new_n7812_ = ~new_n7585_ & ~new_n7811_;
  assign new_n7813_ = ~new_n7621_ & new_n7811_;
  assign new_n7814_ = new_n7807_ & ~new_n7813_;
  assign new_n7815_ = ~new_n7812_ & new_n7814_;
  assign new_n7816_ = ~new_n7810_ & ~new_n7815_;
  assign new_n7817_ = new_n7784_ & ~new_n7816_;
  assign new_n7818_ = pi0592 & ~new_n7621_;
  assign new_n7819_ = ~pi0592 & ~new_n7585_;
  assign new_n7820_ = ~new_n7818_ & ~new_n7819_;
  assign new_n7821_ = ~new_n7784_ & new_n7820_;
  assign new_n7822_ = ~new_n7817_ & ~new_n7821_;
  assign new_n7823_ = pi1199 & new_n7822_;
  assign new_n7824_ = ~pi1196 & ~new_n7783_;
  assign new_n7825_ = new_n7820_ & ~new_n7824_;
  assign new_n7826_ = new_n7585_ & ~new_n7783_;
  assign new_n7827_ = ~pi1196 & new_n7826_;
  assign new_n7828_ = ~new_n7825_ & ~new_n7827_;
  assign new_n7829_ = ~new_n7757_ & ~new_n7828_;
  assign new_n7830_ = new_n7783_ & new_n7820_;
  assign new_n7831_ = ~new_n7826_ & ~new_n7830_;
  assign new_n7832_ = new_n7757_ & ~new_n7831_;
  assign new_n7833_ = ~pi1199 & ~new_n7832_;
  assign new_n7834_ = ~new_n7829_ & new_n7833_;
  assign new_n7835_ = ~new_n7823_ & ~new_n7834_;
  assign new_n7836_ = ~pi0374 & ~new_n7835_;
  assign new_n7837_ = ~pi1198 & new_n7834_;
  assign new_n7838_ = ~pi1198 & pi1199;
  assign new_n7839_ = new_n7822_ & new_n7838_;
  assign new_n7840_ = pi1198 & ~new_n7820_;
  assign new_n7841_ = ~new_n7839_ & ~new_n7840_;
  assign new_n7842_ = ~new_n7837_ & new_n7841_;
  assign new_n7843_ = pi0374 & ~new_n7842_;
  assign new_n7844_ = ~new_n7836_ & ~new_n7843_;
  assign new_n7845_ = ~pi0369 & ~new_n7844_;
  assign new_n7846_ = ~pi0374 & ~new_n7842_;
  assign new_n7847_ = pi0374 & ~new_n7835_;
  assign new_n7848_ = ~new_n7846_ & ~new_n7847_;
  assign new_n7849_ = pi0369 & ~new_n7848_;
  assign new_n7850_ = ~new_n7845_ & ~new_n7849_;
  assign new_n7851_ = ~pi0370 & ~new_n7850_;
  assign new_n7852_ = pi0369 & ~new_n7844_;
  assign new_n7853_ = ~pi0369 & ~new_n7848_;
  assign new_n7854_ = ~new_n7852_ & ~new_n7853_;
  assign new_n7855_ = pi0370 & ~new_n7854_;
  assign new_n7856_ = ~new_n7851_ & ~new_n7855_;
  assign new_n7857_ = ~pi0371 & ~new_n7856_;
  assign new_n7858_ = ~pi0370 & ~new_n7854_;
  assign new_n7859_ = pi0370 & ~new_n7850_;
  assign new_n7860_ = ~new_n7858_ & ~new_n7859_;
  assign new_n7861_ = pi0371 & ~new_n7860_;
  assign new_n7862_ = ~new_n7857_ & ~new_n7861_;
  assign new_n7863_ = ~pi0373 & ~new_n7862_;
  assign new_n7864_ = ~pi0371 & ~new_n7860_;
  assign new_n7865_ = pi0371 & ~new_n7856_;
  assign new_n7866_ = ~new_n7864_ & ~new_n7865_;
  assign new_n7867_ = pi0373 & ~new_n7866_;
  assign new_n7868_ = ~new_n7863_ & ~new_n7867_;
  assign new_n7869_ = ~pi0375 & new_n7868_;
  assign new_n7870_ = pi0384 & ~pi0442;
  assign new_n7871_ = ~pi0384 & pi0442;
  assign new_n7872_ = ~new_n7870_ & ~new_n7871_;
  assign new_n7873_ = pi0440 & ~new_n7872_;
  assign new_n7874_ = ~pi0440 & new_n7872_;
  assign new_n7875_ = ~new_n7873_ & ~new_n7874_;
  assign new_n7876_ = ~pi0373 & ~new_n7866_;
  assign new_n7877_ = pi0373 & ~new_n7862_;
  assign new_n7878_ = ~new_n7876_ & ~new_n7877_;
  assign new_n7879_ = pi0375 & new_n7878_;
  assign new_n7880_ = ~new_n7875_ & ~new_n7879_;
  assign new_n7881_ = ~new_n7869_ & new_n7880_;
  assign new_n7882_ = pi0375 & new_n7868_;
  assign new_n7883_ = ~pi0375 & new_n7878_;
  assign new_n7884_ = new_n7875_ & ~new_n7883_;
  assign new_n7885_ = ~new_n7882_ & new_n7884_;
  assign new_n7886_ = ~pi0591 & ~new_n7885_;
  assign new_n7887_ = ~new_n7881_ & new_n7886_;
  assign new_n7888_ = pi1197 & ~new_n7659_;
  assign new_n7889_ = pi0328 & ~pi0408;
  assign new_n7890_ = ~pi0328 & pi0408;
  assign new_n7891_ = ~new_n7889_ & ~new_n7890_;
  assign new_n7892_ = ~pi0394 & ~pi0396;
  assign new_n7893_ = pi0394 & pi0396;
  assign new_n7894_ = ~new_n7892_ & ~new_n7893_;
  assign new_n7895_ = new_n7891_ & ~new_n7894_;
  assign new_n7896_ = ~new_n7891_ & new_n7894_;
  assign new_n7897_ = ~new_n7895_ & ~new_n7896_;
  assign new_n7898_ = pi0398 & ~pi0399;
  assign new_n7899_ = ~pi0398 & pi0399;
  assign new_n7900_ = ~new_n7898_ & ~new_n7899_;
  assign new_n7901_ = pi0395 & new_n7900_;
  assign new_n7902_ = ~pi0395 & ~new_n7900_;
  assign new_n7903_ = ~new_n7901_ & ~new_n7902_;
  assign new_n7904_ = pi0329 & ~new_n7903_;
  assign new_n7905_ = ~pi0329 & new_n7903_;
  assign new_n7906_ = ~new_n7904_ & ~new_n7905_;
  assign new_n7907_ = pi0400 & ~new_n7906_;
  assign new_n7908_ = ~pi0400 & new_n7906_;
  assign new_n7909_ = ~new_n7907_ & ~new_n7908_;
  assign new_n7910_ = new_n7897_ & new_n7909_;
  assign new_n7911_ = ~new_n7897_ & ~new_n7909_;
  assign new_n7912_ = ~new_n7910_ & ~new_n7911_;
  assign new_n7913_ = pi1198 & ~new_n7912_;
  assign new_n7914_ = new_n7659_ & new_n7913_;
  assign new_n7915_ = pi0390 & ~pi0410;
  assign new_n7916_ = ~pi0390 & pi0410;
  assign new_n7917_ = ~new_n7915_ & ~new_n7916_;
  assign new_n7918_ = pi0397 & ~pi0412;
  assign new_n7919_ = ~pi0397 & pi0412;
  assign new_n7920_ = ~new_n7918_ & ~new_n7919_;
  assign new_n7921_ = pi0404 & new_n7920_;
  assign new_n7922_ = ~pi0404 & ~new_n7920_;
  assign new_n7923_ = ~new_n7921_ & ~new_n7922_;
  assign new_n7924_ = pi0319 & ~pi0324;
  assign new_n7925_ = ~pi0319 & pi0324;
  assign new_n7926_ = ~new_n7924_ & ~new_n7925_;
  assign new_n7927_ = pi0456 & ~new_n7926_;
  assign new_n7928_ = ~pi0456 & new_n7926_;
  assign new_n7929_ = ~new_n7927_ & ~new_n7928_;
  assign new_n7930_ = new_n7923_ & ~new_n7929_;
  assign new_n7931_ = ~new_n7923_ & new_n7929_;
  assign new_n7932_ = ~new_n7930_ & ~new_n7931_;
  assign new_n7933_ = new_n7917_ & new_n7932_;
  assign new_n7934_ = ~new_n7917_ & ~new_n7932_;
  assign new_n7935_ = ~new_n7933_ & ~new_n7934_;
  assign new_n7936_ = pi0411 & new_n7935_;
  assign new_n7937_ = ~pi0411 & ~new_n7935_;
  assign new_n7938_ = ~new_n7936_ & ~new_n7937_;
  assign new_n7939_ = new_n7559_ & new_n7938_;
  assign new_n7940_ = new_n7556_ & ~new_n7939_;
  assign new_n7941_ = new_n7609_ & ~new_n7940_;
  assign new_n7942_ = ~new_n7577_ & new_n7614_;
  assign new_n7943_ = new_n7571_ & new_n7938_;
  assign new_n7944_ = new_n7572_ & ~new_n7943_;
  assign new_n7945_ = new_n7942_ & ~new_n7944_;
  assign new_n7946_ = ~pi0075 & ~pi0592;
  assign new_n7947_ = pi1196 & new_n7946_;
  assign new_n7948_ = ~new_n7945_ & new_n7947_;
  assign new_n7949_ = ~new_n7941_ & new_n7948_;
  assign new_n7950_ = ~pi1196 & new_n7582_;
  assign new_n7951_ = ~new_n7949_ & ~new_n7950_;
  assign new_n7952_ = ~pi1199 & ~new_n7951_;
  assign new_n7953_ = pi0318 & ~pi0409;
  assign new_n7954_ = ~pi0318 & pi0409;
  assign new_n7955_ = ~new_n7953_ & ~new_n7954_;
  assign new_n7956_ = pi0401 & ~pi0402;
  assign new_n7957_ = ~pi0401 & pi0402;
  assign new_n7958_ = ~new_n7956_ & ~new_n7957_;
  assign new_n7959_ = pi0406 & new_n7958_;
  assign new_n7960_ = ~pi0406 & ~new_n7958_;
  assign new_n7961_ = ~new_n7959_ & ~new_n7960_;
  assign new_n7962_ = ~pi0403 & ~pi0405;
  assign new_n7963_ = pi0403 & pi0405;
  assign new_n7964_ = ~new_n7962_ & ~new_n7963_;
  assign new_n7965_ = pi0325 & ~pi0326;
  assign new_n7966_ = ~pi0325 & pi0326;
  assign new_n7967_ = ~new_n7965_ & ~new_n7966_;
  assign new_n7968_ = new_n7964_ & new_n7967_;
  assign new_n7969_ = ~new_n7964_ & ~new_n7967_;
  assign new_n7970_ = ~new_n7968_ & ~new_n7969_;
  assign new_n7971_ = new_n7961_ & ~new_n7970_;
  assign new_n7972_ = ~new_n7961_ & new_n7970_;
  assign new_n7973_ = ~new_n7971_ & ~new_n7972_;
  assign new_n7974_ = new_n7955_ & new_n7973_;
  assign new_n7975_ = ~new_n7955_ & ~new_n7973_;
  assign new_n7976_ = ~new_n7974_ & ~new_n7975_;
  assign new_n7977_ = pi1196 & ~new_n7938_;
  assign new_n7978_ = ~pi0075 & new_n7977_;
  assign new_n7979_ = ~new_n7976_ & ~new_n7978_;
  assign new_n7980_ = new_n7559_ & new_n7979_;
  assign new_n7981_ = new_n7556_ & ~new_n7980_;
  assign new_n7982_ = new_n7609_ & ~new_n7981_;
  assign new_n7983_ = new_n7571_ & ~new_n7976_;
  assign new_n7984_ = new_n7572_ & ~new_n7983_;
  assign new_n7985_ = new_n7942_ & ~new_n7984_;
  assign new_n7986_ = ~new_n7944_ & new_n7985_;
  assign new_n7987_ = ~pi1196 & new_n7985_;
  assign new_n7988_ = pi1199 & new_n7946_;
  assign new_n7989_ = ~new_n7987_ & new_n7988_;
  assign new_n7990_ = ~new_n7986_ & new_n7989_;
  assign new_n7991_ = ~new_n7982_ & new_n7990_;
  assign new_n7992_ = ~new_n7583_ & ~new_n7946_;
  assign new_n7993_ = ~new_n7991_ & ~new_n7992_;
  assign new_n7994_ = ~new_n7952_ & new_n7993_;
  assign new_n7995_ = pi0567 & ~new_n7994_;
  assign new_n7996_ = new_n7495_ & ~new_n7913_;
  assign new_n7997_ = ~new_n7995_ & new_n7996_;
  assign new_n7998_ = ~new_n7914_ & ~new_n7997_;
  assign new_n7999_ = ~pi1197 & new_n7998_;
  assign new_n8000_ = ~new_n7888_ & ~new_n7999_;
  assign new_n8001_ = pi0333 & ~new_n8000_;
  assign new_n8002_ = ~pi0333 & new_n7998_;
  assign new_n8003_ = ~new_n8001_ & ~new_n8002_;
  assign new_n8004_ = pi0391 & ~new_n8003_;
  assign new_n8005_ = pi0333 & ~new_n7998_;
  assign new_n8006_ = ~pi0333 & new_n8000_;
  assign new_n8007_ = ~new_n8005_ & ~new_n8006_;
  assign new_n8008_ = ~pi0391 & new_n8007_;
  assign new_n8009_ = ~new_n8004_ & ~new_n8008_;
  assign new_n8010_ = ~pi0392 & ~new_n8009_;
  assign new_n8011_ = ~pi0391 & ~new_n8003_;
  assign new_n8012_ = pi0391 & new_n8007_;
  assign new_n8013_ = ~new_n8011_ & ~new_n8012_;
  assign new_n8014_ = pi0392 & ~new_n8013_;
  assign new_n8015_ = ~new_n8010_ & ~new_n8014_;
  assign new_n8016_ = ~pi0393 & ~new_n8015_;
  assign new_n8017_ = ~pi0392 & ~new_n8013_;
  assign new_n8018_ = pi0392 & ~new_n8009_;
  assign new_n8019_ = ~new_n8017_ & ~new_n8018_;
  assign new_n8020_ = pi0393 & ~new_n8019_;
  assign new_n8021_ = ~new_n8016_ & ~new_n8020_;
  assign new_n8022_ = pi0334 & new_n8021_;
  assign new_n8023_ = pi0407 & ~pi0463;
  assign new_n8024_ = ~pi0407 & pi0463;
  assign new_n8025_ = ~new_n8023_ & ~new_n8024_;
  assign new_n8026_ = pi0335 & ~pi0413;
  assign new_n8027_ = ~pi0335 & pi0413;
  assign new_n8028_ = ~new_n8026_ & ~new_n8027_;
  assign new_n8029_ = new_n8025_ & new_n8028_;
  assign new_n8030_ = ~new_n8025_ & ~new_n8028_;
  assign new_n8031_ = ~new_n8029_ & ~new_n8030_;
  assign new_n8032_ = ~pi0393 & ~new_n8019_;
  assign new_n8033_ = pi0393 & ~new_n8015_;
  assign new_n8034_ = ~new_n8032_ & ~new_n8033_;
  assign new_n8035_ = ~pi0334 & new_n8034_;
  assign new_n8036_ = ~new_n8031_ & ~new_n8035_;
  assign new_n8037_ = ~new_n8022_ & new_n8036_;
  assign new_n8038_ = pi0334 & new_n8034_;
  assign new_n8039_ = ~pi0334 & new_n8021_;
  assign new_n8040_ = new_n8031_ & ~new_n8039_;
  assign new_n8041_ = ~new_n8038_ & new_n8040_;
  assign new_n8042_ = pi0591 & ~new_n8041_;
  assign new_n8043_ = ~new_n8037_ & new_n8042_;
  assign new_n8044_ = ~pi0590 & ~new_n8043_;
  assign new_n8045_ = ~new_n7887_ & new_n8044_;
  assign new_n8046_ = new_n7733_ & ~new_n8045_;
  assign new_n8047_ = ~new_n7730_ & new_n8046_;
  assign new_n8048_ = new_n7502_ & new_n7562_;
  assign new_n8049_ = pi1091 & ~new_n8048_;
  assign new_n8050_ = new_n7501_ & ~new_n8049_;
  assign new_n8051_ = ~pi0122 & pi1093;
  assign new_n8052_ = ~pi0098 & new_n7511_;
  assign new_n8053_ = new_n8051_ & new_n8052_;
  assign new_n8054_ = ~pi1091 & ~new_n8053_;
  assign new_n8055_ = new_n8050_ & ~new_n8054_;
  assign new_n8056_ = new_n7511_ & new_n8051_;
  assign new_n8057_ = ~pi1091 & new_n8056_;
  assign new_n8058_ = ~pi0098 & new_n8057_;
  assign new_n8059_ = ~new_n7501_ & new_n8058_;
  assign new_n8060_ = pi0075 & ~new_n8059_;
  assign new_n8061_ = ~new_n8055_ & new_n8060_;
  assign new_n8062_ = ~pi0039 & ~new_n7537_;
  assign new_n8063_ = ~pi0122 & new_n8052_;
  assign new_n8064_ = pi0122 & new_n7514_;
  assign new_n8065_ = ~new_n8063_ & ~new_n8064_;
  assign new_n8066_ = pi1093 & ~new_n8065_;
  assign new_n8067_ = new_n7538_ & ~new_n8066_;
  assign new_n8068_ = new_n8062_ & ~new_n8067_;
  assign new_n8069_ = pi1091 & ~new_n7543_;
  assign new_n8070_ = ~new_n8054_ & ~new_n8069_;
  assign new_n8071_ = ~new_n6215_ & new_n8070_;
  assign new_n8072_ = new_n6215_ & new_n8058_;
  assign new_n8073_ = ~new_n8071_ & ~new_n8072_;
  assign new_n8074_ = ~new_n6212_ & new_n8073_;
  assign new_n8075_ = ~pi0216 & new_n6453_;
  assign new_n8076_ = new_n6221_ & new_n8070_;
  assign new_n8077_ = ~new_n6221_ & new_n8058_;
  assign new_n8078_ = ~new_n8076_ & ~new_n8077_;
  assign new_n8079_ = new_n6212_ & new_n8078_;
  assign new_n8080_ = new_n8075_ & ~new_n8079_;
  assign new_n8081_ = ~new_n8074_ & new_n8080_;
  assign new_n8082_ = new_n8058_ & ~new_n8075_;
  assign new_n8083_ = pi0299 & ~new_n8082_;
  assign new_n8084_ = ~new_n8081_ & new_n8083_;
  assign new_n8085_ = ~new_n6238_ & new_n8073_;
  assign new_n8086_ = ~pi0223 & new_n5791_;
  assign new_n8087_ = new_n6238_ & new_n8078_;
  assign new_n8088_ = new_n8086_ & ~new_n8087_;
  assign new_n8089_ = ~new_n8085_ & new_n8088_;
  assign new_n8090_ = new_n8058_ & ~new_n8086_;
  assign new_n8091_ = ~pi0299 & ~new_n8090_;
  assign new_n8092_ = ~new_n8089_ & new_n8091_;
  assign new_n8093_ = pi0039 & ~new_n8092_;
  assign new_n8094_ = ~new_n8084_ & new_n8093_;
  assign new_n8095_ = ~new_n8068_ & ~new_n8094_;
  assign new_n8096_ = ~pi0038 & ~new_n8095_;
  assign new_n8097_ = pi0038 & new_n8058_;
  assign new_n8098_ = ~pi0100 & ~new_n8097_;
  assign new_n8099_ = ~new_n8096_ & new_n8098_;
  assign new_n8100_ = pi0228 & ~new_n7500_;
  assign new_n8101_ = pi1091 & ~new_n7563_;
  assign new_n8102_ = ~new_n8054_ & ~new_n8101_;
  assign new_n8103_ = new_n8100_ & ~new_n8102_;
  assign new_n8104_ = ~new_n8058_ & ~new_n8100_;
  assign new_n8105_ = new_n3186_ & ~new_n8104_;
  assign new_n8106_ = ~new_n8103_ & new_n8105_;
  assign new_n8107_ = ~new_n3186_ & new_n8058_;
  assign new_n8108_ = pi0100 & ~new_n8107_;
  assign new_n8109_ = ~new_n8106_ & new_n8108_;
  assign new_n8110_ = ~pi0087 & ~new_n8109_;
  assign new_n8111_ = ~new_n8099_ & new_n8110_;
  assign new_n8112_ = pi0122 & new_n7571_;
  assign new_n8113_ = ~new_n8063_ & ~new_n8112_;
  assign new_n8114_ = pi1093 & ~new_n8113_;
  assign new_n8115_ = new_n7611_ & ~new_n8114_;
  assign new_n8116_ = new_n3212_ & ~new_n7612_;
  assign new_n8117_ = ~new_n8115_ & new_n8116_;
  assign new_n8118_ = ~new_n8058_ & ~new_n8117_;
  assign new_n8119_ = pi0087 & ~new_n8118_;
  assign new_n8120_ = ~pi0075 & ~new_n8119_;
  assign new_n8121_ = ~new_n8111_ & new_n8120_;
  assign new_n8122_ = ~new_n8061_ & ~new_n8121_;
  assign new_n8123_ = pi0567 & ~new_n8122_;
  assign new_n8124_ = new_n7495_ & ~new_n8123_;
  assign new_n8125_ = pi0567 & new_n8058_;
  assign new_n8126_ = ~new_n7455_ & new_n8125_;
  assign new_n8127_ = ~new_n8124_ & ~new_n8126_;
  assign new_n8128_ = pi0592 & new_n8127_;
  assign new_n8129_ = ~new_n7657_ & ~new_n8128_;
  assign new_n8130_ = new_n7454_ & ~new_n8129_;
  assign new_n8131_ = pi0455 & ~new_n8129_;
  assign new_n8132_ = ~pi0455 & new_n8127_;
  assign new_n8133_ = ~new_n8131_ & ~new_n8132_;
  assign new_n8134_ = pi0452 & ~new_n8133_;
  assign new_n8135_ = pi0355 & ~new_n7645_;
  assign new_n8136_ = ~pi0355 & new_n7645_;
  assign new_n8137_ = ~new_n8135_ & ~new_n8136_;
  assign new_n8138_ = ~pi0455 & ~new_n8129_;
  assign new_n8139_ = pi0455 & new_n8127_;
  assign new_n8140_ = ~new_n8138_ & ~new_n8139_;
  assign new_n8141_ = ~pi0452 & ~new_n8140_;
  assign new_n8142_ = new_n8137_ & ~new_n8141_;
  assign new_n8143_ = ~new_n8134_ & new_n8142_;
  assign new_n8144_ = pi0452 & ~new_n8140_;
  assign new_n8145_ = ~pi0452 & ~new_n8133_;
  assign new_n8146_ = ~new_n8137_ & ~new_n8145_;
  assign new_n8147_ = ~new_n8144_ & new_n8146_;
  assign new_n8148_ = pi1196 & ~new_n8147_;
  assign new_n8149_ = ~new_n8143_ & new_n8148_;
  assign new_n8150_ = ~pi1196 & new_n8127_;
  assign new_n8151_ = ~pi1198 & ~new_n8150_;
  assign new_n8152_ = ~new_n8149_ & new_n8151_;
  assign new_n8153_ = ~new_n7650_ & new_n8127_;
  assign new_n8154_ = new_n7653_ & ~new_n8153_;
  assign new_n8155_ = ~new_n7586_ & new_n8127_;
  assign new_n8156_ = new_n7623_ & ~new_n8155_;
  assign new_n8157_ = ~new_n7649_ & ~new_n8156_;
  assign new_n8158_ = ~new_n8154_ & new_n8157_;
  assign new_n8159_ = new_n7649_ & ~new_n8129_;
  assign new_n8160_ = pi1198 & ~new_n8159_;
  assign new_n8161_ = ~new_n8158_ & new_n8160_;
  assign new_n8162_ = ~new_n7454_ & ~new_n8161_;
  assign new_n8163_ = ~new_n8152_ & new_n8162_;
  assign new_n8164_ = ~new_n8130_ & ~new_n8163_;
  assign new_n8165_ = ~new_n7429_ & ~new_n8164_;
  assign new_n8166_ = pi1199 & ~new_n8129_;
  assign new_n8167_ = pi0351 & new_n8166_;
  assign new_n8168_ = ~new_n8165_ & ~new_n8167_;
  assign new_n8169_ = ~pi0461 & ~new_n8168_;
  assign new_n8170_ = ~new_n7703_ & ~new_n8164_;
  assign new_n8171_ = ~pi0351 & new_n8166_;
  assign new_n8172_ = ~new_n8170_ & ~new_n8171_;
  assign new_n8173_ = pi0461 & ~new_n8172_;
  assign new_n8174_ = ~new_n8169_ & ~new_n8173_;
  assign new_n8175_ = ~pi0357 & ~new_n8174_;
  assign new_n8176_ = ~pi0461 & ~new_n8172_;
  assign new_n8177_ = pi0461 & ~new_n8168_;
  assign new_n8178_ = ~new_n8176_ & ~new_n8177_;
  assign new_n8179_ = pi0357 & ~new_n8178_;
  assign new_n8180_ = ~new_n8175_ & ~new_n8179_;
  assign new_n8181_ = ~pi0356 & ~new_n8180_;
  assign new_n8182_ = ~pi0357 & ~new_n8178_;
  assign new_n8183_ = pi0357 & ~new_n8174_;
  assign new_n8184_ = ~new_n8182_ & ~new_n8183_;
  assign new_n8185_ = pi0356 & ~new_n8184_;
  assign new_n8186_ = ~new_n8181_ & ~new_n8185_;
  assign new_n8187_ = new_n7428_ & ~new_n8186_;
  assign new_n8188_ = ~pi0356 & ~new_n8184_;
  assign new_n8189_ = pi0356 & ~new_n8180_;
  assign new_n8190_ = ~new_n8188_ & ~new_n8189_;
  assign new_n8191_ = ~new_n7428_ & ~new_n8190_;
  assign new_n8192_ = ~pi0591 & ~new_n8191_;
  assign new_n8193_ = ~new_n8187_ & new_n8192_;
  assign new_n8194_ = pi0591 & ~new_n8127_;
  assign new_n8195_ = pi0590 & ~new_n8194_;
  assign new_n8196_ = ~new_n8193_ & new_n8195_;
  assign new_n8197_ = pi0375 & new_n7875_;
  assign new_n8198_ = ~pi0375 & ~new_n7875_;
  assign new_n8199_ = ~new_n8197_ & ~new_n8198_;
  assign new_n8200_ = pi0373 & ~new_n8199_;
  assign new_n8201_ = ~pi0373 & new_n8199_;
  assign new_n8202_ = ~new_n8200_ & ~new_n8201_;
  assign new_n8203_ = ~pi0592 & new_n8127_;
  assign new_n8204_ = ~new_n7818_ & ~new_n8203_;
  assign new_n8205_ = ~new_n7784_ & new_n8204_;
  assign new_n8206_ = new_n7784_ & ~new_n8127_;
  assign new_n8207_ = ~pi1199 & ~new_n8206_;
  assign new_n8208_ = ~new_n8205_ & new_n8207_;
  assign new_n8209_ = ~new_n7811_ & new_n8127_;
  assign new_n8210_ = new_n7814_ & ~new_n8209_;
  assign new_n8211_ = ~new_n7785_ & new_n8127_;
  assign new_n8212_ = new_n7809_ & ~new_n8211_;
  assign new_n8213_ = ~new_n8210_ & ~new_n8212_;
  assign new_n8214_ = new_n7784_ & ~new_n8213_;
  assign new_n8215_ = pi1199 & ~new_n8205_;
  assign new_n8216_ = ~new_n8214_ & new_n8215_;
  assign new_n8217_ = ~new_n8208_ & ~new_n8216_;
  assign new_n8218_ = ~pi0374 & ~new_n8217_;
  assign new_n8219_ = ~pi1198 & ~new_n8217_;
  assign new_n8220_ = pi1198 & ~new_n8204_;
  assign new_n8221_ = ~new_n8219_ & ~new_n8220_;
  assign new_n8222_ = pi0374 & ~new_n8221_;
  assign new_n8223_ = ~new_n8218_ & ~new_n8222_;
  assign new_n8224_ = ~pi0369 & ~new_n8223_;
  assign new_n8225_ = ~pi0374 & ~new_n8221_;
  assign new_n8226_ = pi0374 & ~new_n8217_;
  assign new_n8227_ = ~new_n8225_ & ~new_n8226_;
  assign new_n8228_ = pi0369 & ~new_n8227_;
  assign new_n8229_ = ~new_n8224_ & ~new_n8228_;
  assign new_n8230_ = ~pi0370 & ~new_n8229_;
  assign new_n8231_ = pi0369 & ~new_n8223_;
  assign new_n8232_ = ~pi0369 & ~new_n8227_;
  assign new_n8233_ = ~new_n8231_ & ~new_n8232_;
  assign new_n8234_ = pi0370 & ~new_n8233_;
  assign new_n8235_ = ~new_n8230_ & ~new_n8234_;
  assign new_n8236_ = ~pi0371 & ~new_n8235_;
  assign new_n8237_ = ~pi0370 & ~new_n8233_;
  assign new_n8238_ = pi0370 & ~new_n8229_;
  assign new_n8239_ = ~new_n8237_ & ~new_n8238_;
  assign new_n8240_ = pi0371 & ~new_n8239_;
  assign new_n8241_ = ~new_n8236_ & ~new_n8240_;
  assign new_n8242_ = new_n8202_ & ~new_n8241_;
  assign new_n8243_ = ~pi0371 & ~new_n8239_;
  assign new_n8244_ = pi0371 & ~new_n8235_;
  assign new_n8245_ = ~new_n8243_ & ~new_n8244_;
  assign new_n8246_ = ~new_n8202_ & ~new_n8245_;
  assign new_n8247_ = ~pi0591 & ~new_n8246_;
  assign new_n8248_ = ~new_n8242_ & new_n8247_;
  assign new_n8249_ = pi0334 & ~new_n8031_;
  assign new_n8250_ = ~pi0334 & new_n8031_;
  assign new_n8251_ = ~new_n8249_ & ~new_n8250_;
  assign new_n8252_ = pi0393 & new_n8251_;
  assign new_n8253_ = ~pi0393 & ~new_n8251_;
  assign new_n8254_ = ~new_n8252_ & ~new_n8253_;
  assign new_n8255_ = ~pi0592 & pi1196;
  assign new_n8256_ = new_n7938_ & new_n8053_;
  assign new_n8257_ = ~pi1091 & new_n8256_;
  assign new_n8258_ = pi0567 & new_n8257_;
  assign new_n8259_ = ~new_n7455_ & new_n8258_;
  assign new_n8260_ = ~new_n7976_ & new_n8052_;
  assign new_n8261_ = new_n8259_ & new_n8260_;
  assign new_n8262_ = new_n8255_ & ~new_n8261_;
  assign new_n8263_ = ~new_n8086_ & new_n8257_;
  assign new_n8264_ = ~pi0299 & ~new_n8263_;
  assign new_n8265_ = ~new_n7976_ & new_n8053_;
  assign new_n8266_ = ~pi1091 & new_n8265_;
  assign new_n8267_ = ~new_n8086_ & new_n8266_;
  assign new_n8268_ = ~pi0299 & ~new_n8267_;
  assign new_n8269_ = ~new_n8264_ & ~new_n8268_;
  assign new_n8270_ = ~new_n6215_ & new_n7544_;
  assign new_n8271_ = ~new_n7976_ & new_n8257_;
  assign new_n8272_ = ~new_n8270_ & ~new_n8271_;
  assign new_n8273_ = ~new_n6238_ & new_n8272_;
  assign new_n8274_ = new_n6221_ & new_n7544_;
  assign new_n8275_ = ~new_n8271_ & ~new_n8274_;
  assign new_n8276_ = new_n6238_ & new_n8275_;
  assign new_n8277_ = new_n8086_ & ~new_n8276_;
  assign new_n8278_ = ~new_n8273_ & new_n8277_;
  assign new_n8279_ = ~new_n8269_ & ~new_n8278_;
  assign new_n8280_ = ~new_n8075_ & new_n8257_;
  assign new_n8281_ = pi0299 & ~new_n8280_;
  assign new_n8282_ = ~new_n8075_ & new_n8266_;
  assign new_n8283_ = pi0299 & ~new_n8282_;
  assign new_n8284_ = ~new_n8281_ & ~new_n8283_;
  assign new_n8285_ = ~new_n6212_ & new_n8272_;
  assign new_n8286_ = new_n6212_ & new_n8275_;
  assign new_n8287_ = new_n8075_ & ~new_n8286_;
  assign new_n8288_ = ~new_n8285_ & new_n8287_;
  assign new_n8289_ = ~new_n8284_ & ~new_n8288_;
  assign new_n8290_ = pi0039 & ~new_n8289_;
  assign new_n8291_ = ~new_n8279_ & new_n8290_;
  assign new_n8292_ = new_n7538_ & ~new_n7938_;
  assign new_n8293_ = new_n8068_ & ~new_n8292_;
  assign new_n8294_ = new_n7514_ & ~new_n7976_;
  assign new_n8295_ = pi0122 & ~new_n8294_;
  assign new_n8296_ = ~pi0122 & ~new_n8260_;
  assign new_n8297_ = pi1093 & ~new_n8296_;
  assign new_n8298_ = ~new_n8295_ & new_n8297_;
  assign new_n8299_ = new_n7538_ & ~new_n8298_;
  assign new_n8300_ = new_n8293_ & ~new_n8299_;
  assign new_n8301_ = ~new_n8291_ & ~new_n8300_;
  assign new_n8302_ = ~pi0038 & ~new_n8301_;
  assign new_n8303_ = pi0038 & new_n8257_;
  assign new_n8304_ = ~pi0100 & ~new_n8303_;
  assign new_n8305_ = pi0038 & new_n8266_;
  assign new_n8306_ = ~pi0100 & ~new_n8305_;
  assign new_n8307_ = ~new_n8304_ & ~new_n8306_;
  assign new_n8308_ = ~new_n8302_ & ~new_n8307_;
  assign new_n8309_ = new_n7496_ & new_n7564_;
  assign new_n8310_ = new_n6185_ & ~new_n7497_;
  assign new_n8311_ = ~new_n7496_ & ~new_n8310_;
  assign new_n8312_ = ~pi1091 & ~new_n8271_;
  assign new_n8313_ = new_n8311_ & ~new_n8312_;
  assign new_n8314_ = ~new_n8101_ & new_n8313_;
  assign new_n8315_ = ~new_n8309_ & ~new_n8314_;
  assign new_n8316_ = pi0228 & ~new_n8315_;
  assign new_n8317_ = pi0228 & new_n8311_;
  assign new_n8318_ = new_n8271_ & ~new_n8317_;
  assign new_n8319_ = pi0232 & ~new_n8318_;
  assign new_n8320_ = ~new_n8316_ & new_n8319_;
  assign new_n8321_ = ~pi0232 & ~new_n8271_;
  assign new_n8322_ = ~new_n7565_ & new_n8321_;
  assign new_n8323_ = new_n3186_ & ~new_n8322_;
  assign new_n8324_ = ~new_n8320_ & new_n8323_;
  assign new_n8325_ = ~new_n3186_ & new_n8271_;
  assign new_n8326_ = pi0100 & ~new_n8325_;
  assign new_n8327_ = ~new_n8324_ & new_n8326_;
  assign new_n8328_ = ~new_n8308_ & ~new_n8327_;
  assign new_n8329_ = ~pi0087 & ~new_n8328_;
  assign new_n8330_ = ~new_n3212_ & new_n8257_;
  assign new_n8331_ = pi0087 & ~new_n8330_;
  assign new_n8332_ = ~new_n3212_ & new_n8266_;
  assign new_n8333_ = pi0087 & ~new_n8332_;
  assign new_n8334_ = ~new_n8331_ & ~new_n8333_;
  assign new_n8335_ = new_n7611_ & ~new_n7938_;
  assign new_n8336_ = new_n7611_ & new_n7976_;
  assign new_n8337_ = new_n8117_ & ~new_n8336_;
  assign new_n8338_ = ~new_n8335_ & new_n8337_;
  assign new_n8339_ = ~new_n8334_ & ~new_n8338_;
  assign new_n8340_ = ~new_n8329_ & ~new_n8339_;
  assign new_n8341_ = ~pi0075 & ~new_n8340_;
  assign new_n8342_ = ~new_n7501_ & new_n8257_;
  assign new_n8343_ = pi0075 & ~new_n8342_;
  assign new_n8344_ = ~new_n7501_ & new_n8266_;
  assign new_n8345_ = pi0075 & ~new_n8344_;
  assign new_n8346_ = ~new_n8343_ & ~new_n8345_;
  assign new_n8347_ = new_n8050_ & ~new_n8312_;
  assign new_n8348_ = ~new_n8346_ & ~new_n8347_;
  assign new_n8349_ = ~new_n8341_ & ~new_n8348_;
  assign new_n8350_ = new_n8262_ & ~new_n8349_;
  assign new_n8351_ = pi0567 & new_n8266_;
  assign new_n8352_ = ~new_n7455_ & new_n8351_;
  assign new_n8353_ = ~pi0592 & ~pi1196;
  assign new_n8354_ = ~new_n8352_ & new_n8353_;
  assign new_n8355_ = new_n8333_ & ~new_n8337_;
  assign new_n8356_ = new_n7568_ & ~new_n8266_;
  assign new_n8357_ = new_n8062_ & ~new_n8299_;
  assign new_n8358_ = ~new_n8266_ & ~new_n8274_;
  assign new_n8359_ = new_n6238_ & new_n8358_;
  assign new_n8360_ = ~new_n8266_ & ~new_n8270_;
  assign new_n8361_ = ~new_n6238_ & new_n8360_;
  assign new_n8362_ = new_n8086_ & ~new_n8361_;
  assign new_n8363_ = ~new_n8359_ & new_n8362_;
  assign new_n8364_ = new_n8268_ & ~new_n8363_;
  assign new_n8365_ = new_n6212_ & new_n8358_;
  assign new_n8366_ = ~new_n6212_ & new_n8360_;
  assign new_n8367_ = new_n8075_ & ~new_n8366_;
  assign new_n8368_ = ~new_n8365_ & new_n8367_;
  assign new_n8369_ = new_n8283_ & ~new_n8368_;
  assign new_n8370_ = pi0039 & ~new_n8369_;
  assign new_n8371_ = ~new_n8364_ & new_n8370_;
  assign new_n8372_ = ~new_n8357_ & ~new_n8371_;
  assign new_n8373_ = ~pi0038 & ~new_n8372_;
  assign new_n8374_ = new_n8306_ & ~new_n8373_;
  assign new_n8375_ = ~new_n8356_ & ~new_n8374_;
  assign new_n8376_ = ~pi0087 & ~new_n8375_;
  assign new_n8377_ = ~new_n8355_ & ~new_n8376_;
  assign new_n8378_ = ~pi0075 & ~new_n8377_;
  assign new_n8379_ = ~pi1091 & ~new_n8265_;
  assign new_n8380_ = new_n8050_ & ~new_n8379_;
  assign new_n8381_ = new_n8345_ & ~new_n8380_;
  assign new_n8382_ = ~new_n8378_ & ~new_n8381_;
  assign new_n8383_ = new_n8354_ & ~new_n8382_;
  assign new_n8384_ = ~new_n8350_ & ~new_n8383_;
  assign new_n8385_ = pi0567 & ~new_n8384_;
  assign new_n8386_ = ~new_n8262_ & ~new_n8354_;
  assign new_n8387_ = ~new_n7495_ & ~new_n8386_;
  assign new_n8388_ = pi1199 & ~new_n8387_;
  assign new_n8389_ = ~new_n8385_ & new_n8388_;
  assign new_n8390_ = ~new_n8257_ & ~new_n8274_;
  assign new_n8391_ = new_n6238_ & new_n8390_;
  assign new_n8392_ = ~new_n8257_ & ~new_n8270_;
  assign new_n8393_ = ~new_n6238_ & new_n8392_;
  assign new_n8394_ = new_n8086_ & ~new_n8393_;
  assign new_n8395_ = ~new_n8391_ & new_n8394_;
  assign new_n8396_ = new_n8264_ & ~new_n8395_;
  assign new_n8397_ = new_n6212_ & new_n8390_;
  assign new_n8398_ = ~new_n6212_ & new_n8392_;
  assign new_n8399_ = new_n8075_ & ~new_n8398_;
  assign new_n8400_ = ~new_n8397_ & new_n8399_;
  assign new_n8401_ = new_n8281_ & ~new_n8400_;
  assign new_n8402_ = pi0039 & ~new_n8401_;
  assign new_n8403_ = ~new_n8396_ & new_n8402_;
  assign new_n8404_ = ~new_n8293_ & ~new_n8403_;
  assign new_n8405_ = ~pi0038 & ~new_n8404_;
  assign new_n8406_ = new_n8304_ & ~new_n8405_;
  assign new_n8407_ = new_n7568_ & ~new_n8257_;
  assign new_n8408_ = ~new_n8406_ & ~new_n8407_;
  assign new_n8409_ = ~pi0087 & ~new_n8408_;
  assign new_n8410_ = new_n8117_ & ~new_n8335_;
  assign new_n8411_ = new_n8331_ & ~new_n8410_;
  assign new_n8412_ = ~new_n8409_ & ~new_n8411_;
  assign new_n8413_ = ~pi0075 & ~new_n8412_;
  assign new_n8414_ = ~pi1091 & ~new_n8256_;
  assign new_n8415_ = new_n8050_ & ~new_n8414_;
  assign new_n8416_ = new_n8343_ & ~new_n8415_;
  assign new_n8417_ = ~new_n8413_ & ~new_n8416_;
  assign new_n8418_ = pi0567 & ~new_n8417_;
  assign new_n8419_ = new_n7495_ & ~new_n8418_;
  assign new_n8420_ = new_n8255_ & ~new_n8259_;
  assign new_n8421_ = ~new_n8419_ & new_n8420_;
  assign new_n8422_ = ~pi1199 & ~new_n8150_;
  assign new_n8423_ = ~new_n8421_ & new_n8422_;
  assign new_n8424_ = ~new_n7913_ & ~new_n8423_;
  assign new_n8425_ = ~new_n8389_ & new_n8424_;
  assign new_n8426_ = new_n7657_ & new_n7913_;
  assign new_n8427_ = ~new_n8128_ & ~new_n8426_;
  assign new_n8428_ = ~new_n8425_ & new_n8427_;
  assign new_n8429_ = ~pi0333 & ~new_n8428_;
  assign new_n8430_ = ~pi1197 & ~new_n8428_;
  assign new_n8431_ = pi1197 & ~new_n8129_;
  assign new_n8432_ = ~new_n8430_ & ~new_n8431_;
  assign new_n8433_ = pi0333 & ~new_n8432_;
  assign new_n8434_ = ~new_n8429_ & ~new_n8433_;
  assign new_n8435_ = ~pi0391 & ~new_n8434_;
  assign new_n8436_ = ~pi0333 & ~new_n8432_;
  assign new_n8437_ = pi0333 & ~new_n8428_;
  assign new_n8438_ = ~new_n8436_ & ~new_n8437_;
  assign new_n8439_ = pi0391 & ~new_n8438_;
  assign new_n8440_ = ~new_n8435_ & ~new_n8439_;
  assign new_n8441_ = ~pi0392 & ~new_n8440_;
  assign new_n8442_ = ~pi0391 & ~new_n8438_;
  assign new_n8443_ = pi0391 & ~new_n8434_;
  assign new_n8444_ = ~new_n8442_ & ~new_n8443_;
  assign new_n8445_ = pi0392 & ~new_n8444_;
  assign new_n8446_ = ~new_n8441_ & ~new_n8445_;
  assign new_n8447_ = new_n8254_ & ~new_n8446_;
  assign new_n8448_ = ~pi0392 & ~new_n8444_;
  assign new_n8449_ = pi0392 & ~new_n8440_;
  assign new_n8450_ = ~new_n8448_ & ~new_n8449_;
  assign new_n8451_ = ~new_n8254_ & ~new_n8450_;
  assign new_n8452_ = pi0591 & ~new_n8451_;
  assign new_n8453_ = ~new_n8447_ & new_n8452_;
  assign new_n8454_ = ~pi0590 & ~new_n8453_;
  assign new_n8455_ = ~new_n8248_ & new_n8454_;
  assign new_n8456_ = ~new_n7733_ & ~new_n8455_;
  assign new_n8457_ = ~new_n8196_ & new_n8456_;
  assign new_n8458_ = ~pi0588 & ~new_n8457_;
  assign new_n8459_ = ~new_n8047_ & new_n8458_;
  assign po1038 = pi0057 | ~new_n6305_;
  assign new_n8461_ = pi0433 & ~pi0451;
  assign new_n8462_ = ~pi0433 & pi0451;
  assign new_n8463_ = ~new_n8461_ & ~new_n8462_;
  assign new_n8464_ = pi0449 & new_n8463_;
  assign new_n8465_ = ~pi0449 & ~new_n8463_;
  assign new_n8466_ = ~new_n8464_ & ~new_n8465_;
  assign new_n8467_ = pi0448 & ~new_n8466_;
  assign new_n8468_ = ~pi0448 & new_n8466_;
  assign new_n8469_ = ~new_n8467_ & ~new_n8468_;
  assign new_n8470_ = ~pi0417 & ~pi0418;
  assign new_n8471_ = pi0417 & pi0418;
  assign new_n8472_ = ~new_n8470_ & ~new_n8471_;
  assign new_n8473_ = pi0437 & new_n8472_;
  assign new_n8474_ = ~pi0437 & ~new_n8472_;
  assign new_n8475_ = ~new_n8473_ & ~new_n8474_;
  assign new_n8476_ = pi0453 & ~pi0464;
  assign new_n8477_ = ~pi0453 & pi0464;
  assign new_n8478_ = ~new_n8476_ & ~new_n8477_;
  assign new_n8479_ = new_n8475_ & new_n8478_;
  assign new_n8480_ = ~new_n8475_ & ~new_n8478_;
  assign new_n8481_ = ~new_n8479_ & ~new_n8480_;
  assign new_n8482_ = pi0415 & ~pi0431;
  assign new_n8483_ = ~pi0415 & pi0431;
  assign new_n8484_ = ~new_n8482_ & ~new_n8483_;
  assign new_n8485_ = pi0416 & ~pi0438;
  assign new_n8486_ = ~pi0416 & pi0438;
  assign new_n8487_ = ~new_n8485_ & ~new_n8486_;
  assign new_n8488_ = new_n8484_ & new_n8487_;
  assign new_n8489_ = ~new_n8484_ & ~new_n8487_;
  assign new_n8490_ = ~new_n8488_ & ~new_n8489_;
  assign new_n8491_ = ~new_n8481_ & new_n8490_;
  assign new_n8492_ = new_n8481_ & ~new_n8490_;
  assign new_n8493_ = pi1197 & ~new_n8492_;
  assign new_n8494_ = ~new_n8491_ & new_n8493_;
  assign new_n8495_ = pi0421 & ~pi0454;
  assign new_n8496_ = ~pi0421 & pi0454;
  assign new_n8497_ = ~new_n8495_ & ~new_n8496_;
  assign new_n8498_ = pi0432 & ~pi0459;
  assign new_n8499_ = ~pi0432 & pi0459;
  assign new_n8500_ = ~new_n8498_ & ~new_n8499_;
  assign new_n8501_ = new_n8497_ & ~new_n8500_;
  assign new_n8502_ = ~new_n8497_ & new_n8500_;
  assign new_n8503_ = ~new_n8501_ & ~new_n8502_;
  assign new_n8504_ = ~pi0419 & ~pi0420;
  assign new_n8505_ = pi0419 & pi0420;
  assign new_n8506_ = ~new_n8504_ & ~new_n8505_;
  assign new_n8507_ = pi0423 & ~pi0424;
  assign new_n8508_ = ~pi0423 & pi0424;
  assign new_n8509_ = ~new_n8507_ & ~new_n8508_;
  assign new_n8510_ = new_n8506_ & ~new_n8509_;
  assign new_n8511_ = ~new_n8506_ & new_n8509_;
  assign new_n8512_ = ~new_n8510_ & ~new_n8511_;
  assign new_n8513_ = new_n8503_ & new_n8512_;
  assign new_n8514_ = ~new_n8503_ & ~new_n8512_;
  assign new_n8515_ = ~new_n8513_ & ~new_n8514_;
  assign new_n8516_ = ~pi0425 & new_n8515_;
  assign new_n8517_ = pi0425 & ~new_n8515_;
  assign new_n8518_ = pi1198 & ~new_n8517_;
  assign new_n8519_ = ~new_n8516_ & new_n8518_;
  assign new_n8520_ = ~new_n8494_ & ~new_n8519_;
  assign new_n8521_ = new_n7659_ & ~new_n8520_;
  assign new_n8522_ = ~pi0443 & ~pi0592;
  assign new_n8523_ = ~new_n7585_ & ~new_n8522_;
  assign new_n8524_ = ~new_n7621_ & new_n8522_;
  assign new_n8525_ = ~new_n8523_ & ~new_n8524_;
  assign new_n8526_ = ~pi0444 & ~new_n8525_;
  assign new_n8527_ = pi0443 & ~pi0592;
  assign new_n8528_ = ~new_n7585_ & ~new_n8527_;
  assign new_n8529_ = ~new_n7621_ & new_n8527_;
  assign new_n8530_ = ~new_n8528_ & ~new_n8529_;
  assign new_n8531_ = pi0444 & ~new_n8530_;
  assign new_n8532_ = ~new_n8526_ & ~new_n8531_;
  assign new_n8533_ = pi0436 & ~new_n8532_;
  assign new_n8534_ = ~pi0429 & ~pi0435;
  assign new_n8535_ = pi0429 & pi0435;
  assign new_n8536_ = ~new_n8534_ & ~new_n8535_;
  assign new_n8537_ = pi0434 & ~pi0446;
  assign new_n8538_ = ~pi0434 & pi0446;
  assign new_n8539_ = ~new_n8537_ & ~new_n8538_;
  assign new_n8540_ = pi0414 & ~pi0422;
  assign new_n8541_ = ~pi0414 & pi0422;
  assign new_n8542_ = ~new_n8540_ & ~new_n8541_;
  assign new_n8543_ = new_n8539_ & new_n8542_;
  assign new_n8544_ = ~new_n8539_ & ~new_n8542_;
  assign new_n8545_ = ~new_n8543_ & ~new_n8544_;
  assign new_n8546_ = new_n8536_ & new_n8545_;
  assign new_n8547_ = ~new_n8536_ & ~new_n8545_;
  assign new_n8548_ = ~new_n8546_ & ~new_n8547_;
  assign new_n8549_ = ~pi0444 & ~new_n8530_;
  assign new_n8550_ = pi0444 & ~new_n8525_;
  assign new_n8551_ = ~new_n8549_ & ~new_n8550_;
  assign new_n8552_ = ~pi0436 & ~new_n8551_;
  assign new_n8553_ = ~new_n8548_ & ~new_n8552_;
  assign new_n8554_ = ~new_n8533_ & new_n8553_;
  assign new_n8555_ = pi0436 & ~new_n8551_;
  assign new_n8556_ = ~pi0436 & ~new_n8532_;
  assign new_n8557_ = new_n8548_ & ~new_n8556_;
  assign new_n8558_ = ~new_n8555_ & new_n8557_;
  assign new_n8559_ = pi1196 & ~new_n8558_;
  assign new_n8560_ = ~new_n8554_ & new_n8559_;
  assign new_n8561_ = ~new_n7691_ & new_n8520_;
  assign new_n8562_ = ~new_n8560_ & new_n8561_;
  assign new_n8563_ = ~new_n8521_ & ~new_n8562_;
  assign new_n8564_ = ~pi0428 & ~new_n8563_;
  assign new_n8565_ = pi0428 & new_n7659_;
  assign new_n8566_ = ~new_n8564_ & ~new_n8565_;
  assign new_n8567_ = ~pi0427 & ~new_n8566_;
  assign new_n8568_ = pi0428 & ~new_n8563_;
  assign new_n8569_ = ~pi0428 & new_n7659_;
  assign new_n8570_ = ~new_n8568_ & ~new_n8569_;
  assign new_n8571_ = pi0427 & ~new_n8570_;
  assign new_n8572_ = ~new_n8567_ & ~new_n8571_;
  assign new_n8573_ = pi0430 & ~new_n8572_;
  assign new_n8574_ = ~pi0427 & ~new_n8570_;
  assign new_n8575_ = pi0427 & ~new_n8566_;
  assign new_n8576_ = ~new_n8574_ & ~new_n8575_;
  assign new_n8577_ = ~pi0430 & ~new_n8576_;
  assign new_n8578_ = ~new_n8573_ & ~new_n8577_;
  assign new_n8579_ = pi0426 & ~new_n8578_;
  assign new_n8580_ = pi0430 & ~new_n8576_;
  assign new_n8581_ = ~pi0430 & ~new_n8572_;
  assign new_n8582_ = ~new_n8580_ & ~new_n8581_;
  assign new_n8583_ = ~pi0426 & ~new_n8582_;
  assign new_n8584_ = ~new_n8579_ & ~new_n8583_;
  assign new_n8585_ = pi0445 & ~new_n8584_;
  assign new_n8586_ = pi0426 & ~new_n8582_;
  assign new_n8587_ = ~pi0426 & ~new_n8578_;
  assign new_n8588_ = ~new_n8586_ & ~new_n8587_;
  assign new_n8589_ = ~pi0445 & ~new_n8588_;
  assign new_n8590_ = ~new_n8585_ & ~new_n8589_;
  assign new_n8591_ = new_n8469_ & ~new_n8590_;
  assign new_n8592_ = pi0445 & ~new_n8588_;
  assign new_n8593_ = ~pi0445 & ~new_n8584_;
  assign new_n8594_ = ~new_n8592_ & ~new_n8593_;
  assign new_n8595_ = ~new_n8469_ & ~new_n8594_;
  assign new_n8596_ = pi1199 & ~new_n8595_;
  assign new_n8597_ = ~new_n8591_ & new_n8596_;
  assign new_n8598_ = ~pi0590 & ~pi0591;
  assign new_n8599_ = ~pi1199 & new_n8563_;
  assign new_n8600_ = new_n8598_ & ~new_n8599_;
  assign new_n8601_ = ~new_n8597_ & new_n8600_;
  assign new_n8602_ = new_n7585_ & ~new_n8598_;
  assign new_n8603_ = new_n7733_ & ~new_n8602_;
  assign new_n8604_ = ~new_n8601_ & new_n8603_;
  assign new_n8605_ = new_n8127_ & ~new_n8527_;
  assign new_n8606_ = ~pi0436 & pi0444;
  assign new_n8607_ = pi0436 & ~pi0444;
  assign new_n8608_ = ~new_n8606_ & ~new_n8607_;
  assign new_n8609_ = new_n8548_ & ~new_n8608_;
  assign new_n8610_ = ~new_n8548_ & new_n8608_;
  assign new_n8611_ = ~new_n8609_ & ~new_n8610_;
  assign new_n8612_ = ~new_n8529_ & ~new_n8611_;
  assign new_n8613_ = ~new_n8605_ & new_n8612_;
  assign new_n8614_ = new_n8127_ & ~new_n8522_;
  assign new_n8615_ = ~new_n8524_ & new_n8611_;
  assign new_n8616_ = ~new_n8614_ & new_n8615_;
  assign new_n8617_ = pi1196 & ~new_n8616_;
  assign new_n8618_ = ~new_n8613_ & new_n8617_;
  assign new_n8619_ = ~new_n8150_ & ~new_n8618_;
  assign new_n8620_ = new_n8520_ & ~new_n8619_;
  assign new_n8621_ = ~new_n8129_ & ~new_n8520_;
  assign new_n8622_ = ~new_n8620_ & ~new_n8621_;
  assign new_n8623_ = pi0428 & new_n8622_;
  assign new_n8624_ = ~pi0428 & new_n8129_;
  assign new_n8625_ = pi0427 & ~new_n8624_;
  assign new_n8626_ = ~new_n8623_ & new_n8625_;
  assign new_n8627_ = ~pi0428 & new_n8622_;
  assign new_n8628_ = pi0428 & new_n8129_;
  assign new_n8629_ = ~pi0427 & ~new_n8628_;
  assign new_n8630_ = ~new_n8627_ & new_n8629_;
  assign new_n8631_ = ~new_n8626_ & ~new_n8630_;
  assign new_n8632_ = pi0430 & ~new_n8631_;
  assign new_n8633_ = ~pi0427 & pi0428;
  assign new_n8634_ = pi0427 & ~pi0428;
  assign new_n8635_ = ~new_n8633_ & ~new_n8634_;
  assign new_n8636_ = new_n8129_ & new_n8635_;
  assign new_n8637_ = new_n8622_ & ~new_n8635_;
  assign new_n8638_ = ~new_n8636_ & ~new_n8637_;
  assign new_n8639_ = ~pi0430 & new_n8638_;
  assign new_n8640_ = ~new_n8632_ & ~new_n8639_;
  assign new_n8641_ = ~pi0426 & ~new_n8640_;
  assign new_n8642_ = ~pi0430 & ~new_n8631_;
  assign new_n8643_ = pi0430 & new_n8638_;
  assign new_n8644_ = ~new_n8642_ & ~new_n8643_;
  assign new_n8645_ = pi0426 & ~new_n8644_;
  assign new_n8646_ = ~new_n8641_ & ~new_n8645_;
  assign new_n8647_ = ~pi0445 & ~new_n8646_;
  assign new_n8648_ = ~pi0426 & ~new_n8644_;
  assign new_n8649_ = pi0426 & ~new_n8640_;
  assign new_n8650_ = ~new_n8648_ & ~new_n8649_;
  assign new_n8651_ = pi0445 & ~new_n8650_;
  assign new_n8652_ = ~new_n8647_ & ~new_n8651_;
  assign new_n8653_ = ~pi0448 & new_n8652_;
  assign new_n8654_ = ~pi0445 & ~new_n8650_;
  assign new_n8655_ = pi0445 & ~new_n8646_;
  assign new_n8656_ = ~new_n8654_ & ~new_n8655_;
  assign new_n8657_ = pi0448 & new_n8656_;
  assign new_n8658_ = ~new_n8466_ & ~new_n8657_;
  assign new_n8659_ = ~new_n8653_ & new_n8658_;
  assign new_n8660_ = pi0448 & new_n8652_;
  assign new_n8661_ = ~pi0448 & new_n8656_;
  assign new_n8662_ = new_n8466_ & ~new_n8661_;
  assign new_n8663_ = ~new_n8660_ & new_n8662_;
  assign new_n8664_ = ~new_n8659_ & ~new_n8663_;
  assign new_n8665_ = pi1199 & ~new_n8664_;
  assign new_n8666_ = ~pi1199 & ~new_n8622_;
  assign new_n8667_ = new_n8598_ & ~new_n8666_;
  assign new_n8668_ = ~new_n8665_ & new_n8667_;
  assign new_n8669_ = ~new_n8127_ & ~new_n8598_;
  assign new_n8670_ = ~new_n7733_ & ~new_n8669_;
  assign new_n8671_ = ~new_n8668_ & new_n8670_;
  assign new_n8672_ = ~new_n8604_ & ~new_n8671_;
  assign new_n8673_ = pi0588 & ~new_n8672_;
  assign new_n8674_ = ~po1038 & ~new_n8673_;
  assign new_n8675_ = ~new_n8459_ & new_n8674_;
  assign new_n8676_ = ~pi0592 & new_n7648_;
  assign new_n8677_ = ~new_n7636_ & new_n8125_;
  assign new_n8678_ = ~new_n8676_ & new_n8677_;
  assign new_n8679_ = pi0361 & ~pi0458;
  assign new_n8680_ = ~pi0361 & pi0458;
  assign new_n8681_ = ~new_n8679_ & ~new_n8680_;
  assign new_n8682_ = new_n7630_ & new_n8681_;
  assign new_n8683_ = ~new_n7630_ & ~new_n8681_;
  assign new_n8684_ = ~new_n8682_ & ~new_n8683_;
  assign new_n8685_ = pi0441 & ~new_n8684_;
  assign new_n8686_ = ~pi0441 & new_n8684_;
  assign new_n8687_ = ~pi0592 & ~new_n8686_;
  assign new_n8688_ = ~new_n8685_ & new_n8687_;
  assign new_n8689_ = new_n7636_ & new_n8125_;
  assign new_n8690_ = ~new_n8688_ & new_n8689_;
  assign new_n8691_ = pi1196 & ~new_n8690_;
  assign new_n8692_ = ~new_n8678_ & new_n8691_;
  assign new_n8693_ = ~pi1198 & ~new_n8692_;
  assign new_n8694_ = pi0350 & ~new_n7608_;
  assign new_n8695_ = ~pi0350 & new_n7608_;
  assign new_n8696_ = ~new_n8694_ & ~new_n8695_;
  assign new_n8697_ = ~new_n7649_ & new_n8696_;
  assign new_n8698_ = ~pi0592 & new_n8125_;
  assign new_n8699_ = pi1198 & new_n8698_;
  assign new_n8700_ = new_n8697_ & new_n8699_;
  assign new_n8701_ = ~new_n8693_ & ~new_n8700_;
  assign new_n8702_ = ~new_n7454_ & ~new_n8701_;
  assign new_n8703_ = ~pi0592 & ~new_n8702_;
  assign new_n8704_ = new_n8125_ & ~new_n8703_;
  assign new_n8705_ = ~new_n7703_ & ~new_n8704_;
  assign new_n8706_ = pi0592 & new_n8125_;
  assign new_n8707_ = pi1199 & ~new_n8706_;
  assign new_n8708_ = ~pi0351 & new_n8707_;
  assign new_n8709_ = ~new_n8705_ & ~new_n8708_;
  assign new_n8710_ = ~pi0461 & ~new_n8709_;
  assign new_n8711_ = ~new_n7429_ & ~new_n8704_;
  assign new_n8712_ = pi0351 & new_n8707_;
  assign new_n8713_ = ~new_n8711_ & ~new_n8712_;
  assign new_n8714_ = pi0461 & ~new_n8713_;
  assign new_n8715_ = ~new_n8710_ & ~new_n8714_;
  assign new_n8716_ = ~pi0357 & ~new_n8715_;
  assign new_n8717_ = ~pi0461 & ~new_n8713_;
  assign new_n8718_ = pi0461 & ~new_n8709_;
  assign new_n8719_ = ~new_n8717_ & ~new_n8718_;
  assign new_n8720_ = pi0357 & ~new_n8719_;
  assign new_n8721_ = ~new_n8716_ & ~new_n8720_;
  assign new_n8722_ = pi0356 & ~new_n8721_;
  assign new_n8723_ = ~pi0357 & ~new_n8719_;
  assign new_n8724_ = pi0357 & ~new_n8715_;
  assign new_n8725_ = ~new_n8723_ & ~new_n8724_;
  assign new_n8726_ = ~pi0356 & ~new_n8725_;
  assign new_n8727_ = new_n7428_ & ~new_n8726_;
  assign new_n8728_ = ~new_n8722_ & new_n8727_;
  assign new_n8729_ = pi0356 & ~new_n8725_;
  assign new_n8730_ = ~pi0356 & ~new_n8721_;
  assign new_n8731_ = ~new_n7428_ & ~new_n8730_;
  assign new_n8732_ = ~new_n8729_ & new_n8731_;
  assign new_n8733_ = ~new_n8728_ & ~new_n8732_;
  assign new_n8734_ = pi0590 & ~new_n8733_;
  assign new_n8735_ = pi0592 & ~new_n7784_;
  assign new_n8736_ = ~pi0377 & ~new_n7807_;
  assign new_n8737_ = pi0377 & new_n7807_;
  assign new_n8738_ = ~new_n8736_ & ~new_n8737_;
  assign new_n8739_ = new_n7784_ & ~new_n8738_;
  assign new_n8740_ = pi0592 & ~new_n8739_;
  assign new_n8741_ = new_n8125_ & ~new_n8740_;
  assign new_n8742_ = pi1199 & ~new_n8741_;
  assign new_n8743_ = ~new_n8735_ & ~new_n8742_;
  assign new_n8744_ = new_n8706_ & new_n8743_;
  assign new_n8745_ = ~pi0369 & ~pi0374;
  assign new_n8746_ = pi0369 & pi0374;
  assign new_n8747_ = ~new_n8745_ & ~new_n8746_;
  assign new_n8748_ = ~pi0370 & ~new_n8747_;
  assign new_n8749_ = pi0370 & new_n8747_;
  assign new_n8750_ = ~new_n8748_ & ~new_n8749_;
  assign new_n8751_ = ~pi0371 & ~new_n8750_;
  assign new_n8752_ = pi0371 & new_n8750_;
  assign new_n8753_ = ~new_n8751_ & ~new_n8752_;
  assign new_n8754_ = ~pi0373 & ~new_n8753_;
  assign new_n8755_ = pi0373 & new_n8753_;
  assign new_n8756_ = ~new_n8754_ & ~new_n8755_;
  assign new_n8757_ = pi0375 & ~new_n8756_;
  assign new_n8758_ = ~pi0375 & new_n8756_;
  assign new_n8759_ = ~new_n8757_ & ~new_n8758_;
  assign new_n8760_ = ~new_n7875_ & ~new_n8759_;
  assign new_n8761_ = new_n7875_ & new_n8759_;
  assign new_n8762_ = ~new_n8760_ & ~new_n8761_;
  assign new_n8763_ = new_n8744_ & new_n8762_;
  assign new_n8764_ = ~pi1198 & new_n8744_;
  assign new_n8765_ = ~new_n8698_ & ~new_n8764_;
  assign new_n8766_ = ~new_n8763_ & new_n8765_;
  assign new_n8767_ = ~pi0590 & ~new_n8766_;
  assign new_n8768_ = ~pi0591 & ~new_n8767_;
  assign new_n8769_ = ~new_n8734_ & new_n8768_;
  assign new_n8770_ = pi1197 & ~new_n8706_;
  assign new_n8771_ = ~pi0592 & new_n8351_;
  assign new_n8772_ = ~new_n7977_ & new_n8771_;
  assign new_n8773_ = new_n8707_ & ~new_n8772_;
  assign new_n8774_ = new_n8255_ & new_n8258_;
  assign new_n8775_ = new_n8125_ & ~new_n8255_;
  assign new_n8776_ = ~pi1199 & ~new_n8775_;
  assign new_n8777_ = ~new_n8774_ & new_n8776_;
  assign new_n8778_ = ~new_n8773_ & ~new_n8777_;
  assign new_n8779_ = ~pi1197 & ~new_n8778_;
  assign new_n8780_ = ~new_n8770_ & ~new_n8779_;
  assign new_n8781_ = ~pi0333 & ~new_n8780_;
  assign new_n8782_ = pi1198 & ~new_n8706_;
  assign new_n8783_ = new_n8778_ & ~new_n8782_;
  assign new_n8784_ = ~new_n7912_ & ~new_n8783_;
  assign new_n8785_ = new_n8778_ & ~new_n8784_;
  assign new_n8786_ = ~new_n8781_ & new_n8785_;
  assign new_n8787_ = ~pi0391 & ~new_n8786_;
  assign new_n8788_ = pi0333 & ~new_n8780_;
  assign new_n8789_ = ~pi0333 & ~new_n8778_;
  assign new_n8790_ = ~new_n8784_ & ~new_n8789_;
  assign new_n8791_ = ~new_n8788_ & new_n8790_;
  assign new_n8792_ = pi0391 & ~new_n8791_;
  assign new_n8793_ = ~new_n8787_ & ~new_n8792_;
  assign new_n8794_ = ~pi0392 & ~new_n8793_;
  assign new_n8795_ = ~pi0391 & ~new_n8791_;
  assign new_n8796_ = pi0391 & ~new_n8786_;
  assign new_n8797_ = ~new_n8795_ & ~new_n8796_;
  assign new_n8798_ = pi0392 & ~new_n8797_;
  assign new_n8799_ = ~new_n8794_ & ~new_n8798_;
  assign new_n8800_ = pi0393 & ~new_n8799_;
  assign new_n8801_ = ~pi0392 & ~new_n8797_;
  assign new_n8802_ = pi0392 & ~new_n8793_;
  assign new_n8803_ = ~new_n8801_ & ~new_n8802_;
  assign new_n8804_ = ~pi0393 & ~new_n8803_;
  assign new_n8805_ = new_n8251_ & ~new_n8804_;
  assign new_n8806_ = ~new_n8800_ & new_n8805_;
  assign new_n8807_ = pi0393 & ~new_n8803_;
  assign new_n8808_ = ~pi0393 & ~new_n8799_;
  assign new_n8809_ = ~new_n8251_ & ~new_n8808_;
  assign new_n8810_ = ~new_n8807_ & new_n8809_;
  assign new_n8811_ = ~new_n8806_ & ~new_n8810_;
  assign new_n8812_ = ~pi0590 & ~new_n8811_;
  assign new_n8813_ = pi0590 & new_n8125_;
  assign new_n8814_ = pi0591 & ~new_n8813_;
  assign new_n8815_ = ~new_n8812_ & new_n8814_;
  assign new_n8816_ = ~new_n8769_ & ~new_n8815_;
  assign new_n8817_ = ~pi0588 & ~new_n8816_;
  assign new_n8818_ = ~new_n7733_ & po1038;
  assign new_n8819_ = pi0436 & ~pi0443;
  assign new_n8820_ = ~pi0436 & pi0443;
  assign new_n8821_ = ~new_n8819_ & ~new_n8820_;
  assign new_n8822_ = ~pi0444 & new_n8821_;
  assign new_n8823_ = pi0444 & ~new_n8821_;
  assign new_n8824_ = ~new_n8822_ & ~new_n8823_;
  assign new_n8825_ = new_n8548_ & new_n8824_;
  assign new_n8826_ = ~new_n8548_ & ~new_n8824_;
  assign new_n8827_ = new_n8255_ & ~new_n8826_;
  assign new_n8828_ = ~new_n8825_ & new_n8827_;
  assign new_n8829_ = new_n8520_ & ~new_n8828_;
  assign new_n8830_ = new_n8698_ & new_n8829_;
  assign new_n8831_ = pi0430 & ~new_n8635_;
  assign new_n8832_ = ~pi0430 & new_n8635_;
  assign new_n8833_ = ~new_n8831_ & ~new_n8832_;
  assign new_n8834_ = ~pi0426 & ~new_n8833_;
  assign new_n8835_ = pi0426 & new_n8833_;
  assign new_n8836_ = ~new_n8834_ & ~new_n8835_;
  assign new_n8837_ = ~pi0445 & ~new_n8836_;
  assign new_n8838_ = pi0445 & new_n8836_;
  assign new_n8839_ = ~new_n8837_ & ~new_n8838_;
  assign new_n8840_ = ~pi0448 & ~new_n8839_;
  assign new_n8841_ = pi0448 & new_n8839_;
  assign new_n8842_ = ~new_n8840_ & ~new_n8841_;
  assign new_n8843_ = new_n8830_ & new_n8842_;
  assign new_n8844_ = ~new_n8706_ & ~new_n8843_;
  assign new_n8845_ = ~new_n8466_ & ~new_n8844_;
  assign new_n8846_ = new_n8830_ & ~new_n8842_;
  assign new_n8847_ = ~new_n8706_ & ~new_n8846_;
  assign new_n8848_ = new_n8466_ & ~new_n8847_;
  assign new_n8849_ = pi1199 & ~new_n8848_;
  assign new_n8850_ = ~new_n8845_ & new_n8849_;
  assign new_n8851_ = ~pi1199 & ~new_n8706_;
  assign new_n8852_ = ~new_n8830_ & new_n8851_;
  assign new_n8853_ = new_n8598_ & ~new_n8852_;
  assign new_n8854_ = ~new_n8850_ & new_n8853_;
  assign new_n8855_ = new_n8125_ & ~new_n8598_;
  assign new_n8856_ = pi0588 & ~new_n8855_;
  assign new_n8857_ = ~new_n8854_ & new_n8856_;
  assign new_n8858_ = new_n8818_ & ~new_n8857_;
  assign new_n8859_ = ~new_n8817_ & new_n8858_;
  assign new_n8860_ = ~pi0217 & ~new_n8859_;
  assign new_n8861_ = ~new_n8675_ & new_n8860_;
  assign new_n8862_ = ~new_n7585_ & new_n7733_;
  assign new_n8863_ = ~new_n7733_ & new_n8127_;
  assign new_n8864_ = ~po1038 & ~new_n8863_;
  assign new_n8865_ = ~new_n8862_ & new_n8864_;
  assign new_n8866_ = new_n8125_ & new_n8818_;
  assign new_n8867_ = pi0217 & ~new_n8866_;
  assign new_n8868_ = ~new_n8865_ & new_n8867_;
  assign new_n8869_ = ~pi1161 & ~pi1162;
  assign new_n8870_ = ~pi1163 & new_n8869_;
  assign new_n8871_ = ~new_n8868_ & new_n8870_;
  assign new_n8872_ = ~new_n8861_ & new_n8871_;
  assign new_n8873_ = pi1161 & ~pi1163;
  assign new_n8874_ = new_n2754_ & new_n8873_;
  assign new_n8875_ = ~pi0031 & pi1162;
  assign new_n8876_ = new_n8874_ & new_n8875_;
  assign po0189 = new_n8872_ | new_n8876_;
  assign new_n8878_ = new_n3298_ & new_n3436_;
  assign new_n8879_ = ~pi0055 & ~pi0074;
  assign new_n8880_ = new_n8878_ & new_n8879_;
  assign new_n8881_ = new_n6290_ & new_n8880_;
  assign new_n8882_ = pi0100 & new_n3186_;
  assign new_n8883_ = ~new_n6263_ & ~po1057;
  assign new_n8884_ = new_n6502_ & new_n8883_;
  assign new_n8885_ = ~pi0137 & new_n8884_;
  assign new_n8886_ = pi0129 & new_n3100_;
  assign new_n8887_ = ~pi0137 & pi0252;
  assign new_n8888_ = po1057 & ~new_n7500_;
  assign new_n8889_ = new_n6263_ & ~new_n8888_;
  assign new_n8890_ = new_n8887_ & new_n8889_;
  assign new_n8891_ = new_n8886_ & new_n8890_;
  assign new_n8892_ = ~new_n8885_ & ~new_n8891_;
  assign new_n8893_ = new_n8882_ & ~new_n8892_;
  assign new_n8894_ = ~pi0024 & ~pi0090;
  assign new_n8895_ = new_n6168_ & new_n8894_;
  assign new_n8896_ = pi0050 & new_n2586_;
  assign new_n8897_ = new_n2484_ & new_n8896_;
  assign new_n8898_ = new_n2482_ & new_n2510_;
  assign new_n8899_ = new_n2490_ & new_n8898_;
  assign new_n8900_ = ~pi0093 & new_n8899_;
  assign new_n8901_ = new_n8897_ & new_n8900_;
  assign new_n8902_ = new_n8895_ & new_n8901_;
  assign new_n8903_ = pi0829 & ~pi1093;
  assign new_n8904_ = new_n2799_ & new_n8903_;
  assign po0840 = new_n2795_ | new_n8904_;
  assign new_n8906_ = ~new_n7733_ & ~po0840;
  assign new_n8907_ = ~pi0137 & ~new_n8906_;
  assign new_n8908_ = new_n8902_ & ~new_n8907_;
  assign new_n8909_ = pi0076 & ~pi0084;
  assign new_n8910_ = new_n2468_ & new_n8909_;
  assign new_n8911_ = ~pi0068 & ~pi0073;
  assign new_n8912_ = ~pi0049 & ~pi0066;
  assign new_n8913_ = new_n8911_ & new_n8912_;
  assign new_n8914_ = new_n8910_ & new_n8913_;
  assign new_n8915_ = ~pi0089 & ~pi0102;
  assign new_n8916_ = new_n7463_ & new_n8915_;
  assign new_n8917_ = ~pi0064 & ~pi0081;
  assign new_n8918_ = new_n2476_ & new_n8917_;
  assign new_n8919_ = new_n8916_ & new_n8918_;
  assign new_n8920_ = new_n8914_ & new_n8919_;
  assign new_n8921_ = new_n2451_ & new_n2641_;
  assign new_n8922_ = ~pi0103 & new_n2460_;
  assign new_n8923_ = new_n8921_ & new_n8922_;
  assign new_n8924_ = new_n2455_ & new_n2606_;
  assign new_n8925_ = ~pi0045 & ~pi0048;
  assign new_n8926_ = ~pi0061 & ~pi0104;
  assign new_n8927_ = new_n8925_ & new_n8926_;
  assign new_n8928_ = new_n8924_ & new_n8927_;
  assign new_n8929_ = new_n8923_ & new_n8928_;
  assign new_n8930_ = new_n8920_ & new_n8929_;
  assign new_n8931_ = ~new_n8896_ & ~new_n8930_;
  assign new_n8932_ = new_n2486_ & new_n2491_;
  assign new_n8933_ = ~new_n8931_ & new_n8932_;
  assign new_n8934_ = ~pi0024 & ~new_n8933_;
  assign new_n8935_ = new_n2484_ & new_n8930_;
  assign new_n8936_ = new_n8899_ & new_n8935_;
  assign new_n8937_ = pi0024 & ~new_n8936_;
  assign new_n8938_ = new_n2550_ & new_n2782_;
  assign new_n8939_ = ~pi0137 & new_n7471_;
  assign new_n8940_ = new_n8938_ & new_n8939_;
  assign new_n8941_ = ~new_n8906_ & new_n8940_;
  assign new_n8942_ = ~new_n8937_ & new_n8941_;
  assign new_n8943_ = ~new_n8934_ & new_n8942_;
  assign new_n8944_ = ~new_n8908_ & ~new_n8943_;
  assign new_n8945_ = ~pi0032 & ~new_n8944_;
  assign new_n8946_ = ~pi0024 & ~pi0841;
  assign new_n8947_ = pi0032 & ~new_n8946_;
  assign new_n8948_ = new_n2499_ & new_n8947_;
  assign new_n8949_ = ~new_n8945_ & ~new_n8948_;
  assign new_n8950_ = ~new_n6166_ & ~new_n8949_;
  assign new_n8951_ = ~pi0032 & ~new_n8902_;
  assign new_n8952_ = new_n6166_ & ~new_n6170_;
  assign new_n8953_ = ~new_n8951_ & new_n8952_;
  assign new_n8954_ = ~new_n8950_ & ~new_n8953_;
  assign new_n8955_ = ~pi0095 & new_n3281_;
  assign new_n8956_ = ~new_n8954_ & new_n8955_;
  assign new_n8957_ = ~new_n8893_ & ~new_n8956_;
  assign new_n8958_ = new_n3235_ & ~new_n8957_;
  assign new_n8959_ = ~pi0024 & new_n2548_;
  assign new_n8960_ = new_n2494_ & new_n3098_;
  assign new_n8961_ = ~pi0051 & new_n8960_;
  assign new_n8962_ = new_n8959_ & new_n8961_;
  assign new_n8963_ = ~po0840 & new_n8962_;
  assign new_n8964_ = pi0252 & ~new_n8888_;
  assign new_n8965_ = ~pi0087 & new_n3186_;
  assign new_n8966_ = pi0075 & ~pi0100;
  assign new_n8967_ = new_n8965_ & new_n8966_;
  assign new_n8968_ = ~pi0137 & new_n8967_;
  assign new_n8969_ = ~new_n6282_ & new_n8968_;
  assign new_n8970_ = ~new_n8964_ & new_n8969_;
  assign new_n8971_ = new_n8963_ & new_n8970_;
  assign new_n8972_ = ~new_n8958_ & ~new_n8971_;
  assign po0190 = new_n8881_ & ~new_n8972_;
  assign new_n8974_ = ~pi0195 & ~pi0196;
  assign new_n8975_ = ~pi0138 & new_n8974_;
  assign new_n8976_ = ~pi0139 & new_n8975_;
  assign new_n8977_ = ~pi0118 & new_n8976_;
  assign new_n8978_ = ~pi0079 & new_n8977_;
  assign new_n8979_ = ~pi0034 & new_n8978_;
  assign new_n8980_ = ~pi0033 & ~new_n8979_;
  assign new_n8981_ = pi0149 & pi0157;
  assign new_n8982_ = ~pi0149 & ~pi0157;
  assign new_n8983_ = new_n6185_ & ~new_n8982_;
  assign new_n8984_ = ~new_n8981_ & new_n8983_;
  assign new_n8985_ = pi0232 & new_n8984_;
  assign new_n8986_ = pi0075 & ~new_n8985_;
  assign new_n8987_ = pi0100 & ~new_n8985_;
  assign new_n8988_ = ~new_n8986_ & ~new_n8987_;
  assign new_n8989_ = ~pi0075 & ~pi0100;
  assign new_n8990_ = new_n7499_ & new_n8989_;
  assign new_n8991_ = pi0169 & new_n8990_;
  assign new_n8992_ = new_n8988_ & ~new_n8991_;
  assign new_n8993_ = pi0074 & ~new_n8992_;
  assign new_n8994_ = pi0164 & new_n8990_;
  assign new_n8995_ = new_n8988_ & ~new_n8994_;
  assign new_n8996_ = ~pi0074 & ~new_n8995_;
  assign new_n8997_ = ~new_n3436_ & ~new_n8996_;
  assign new_n8998_ = ~new_n8993_ & new_n8997_;
  assign new_n8999_ = pi0178 & pi0183;
  assign new_n9000_ = ~pi0178 & ~pi0183;
  assign new_n9001_ = new_n6185_ & ~new_n9000_;
  assign new_n9002_ = ~new_n8999_ & new_n9001_;
  assign new_n9003_ = ~pi0299 & ~new_n9002_;
  assign new_n9004_ = pi0299 & ~new_n8984_;
  assign new_n9005_ = pi0232 & ~new_n9004_;
  assign new_n9006_ = ~new_n9003_ & new_n9005_;
  assign new_n9007_ = pi0100 & ~new_n9006_;
  assign new_n9008_ = pi0075 & ~new_n9006_;
  assign new_n9009_ = ~new_n9007_ & ~new_n9008_;
  assign new_n9010_ = pi0191 & ~pi0299;
  assign new_n9011_ = pi0169 & pi0299;
  assign new_n9012_ = ~new_n9010_ & ~new_n9011_;
  assign new_n9013_ = new_n8990_ & ~new_n9012_;
  assign new_n9014_ = new_n9009_ & ~new_n9013_;
  assign new_n9015_ = pi0074 & ~new_n9014_;
  assign new_n9016_ = ~pi0055 & ~new_n9015_;
  assign new_n9017_ = ~pi0186 & ~pi0299;
  assign new_n9018_ = ~pi0164 & pi0299;
  assign new_n9019_ = ~new_n9017_ & ~new_n9018_;
  assign new_n9020_ = new_n7499_ & new_n9019_;
  assign new_n9021_ = new_n8989_ & new_n9020_;
  assign new_n9022_ = new_n9009_ & ~new_n9021_;
  assign new_n9023_ = pi0054 & ~new_n9022_;
  assign new_n9024_ = pi0299 & new_n7499_;
  assign new_n9025_ = ~new_n6132_ & new_n9024_;
  assign new_n9026_ = ~pi0186 & ~new_n9025_;
  assign new_n9027_ = ~new_n6257_ & new_n7499_;
  assign new_n9028_ = pi0186 & ~new_n9027_;
  assign new_n9029_ = pi0164 & ~new_n9028_;
  assign new_n9030_ = ~new_n9026_ & new_n9029_;
  assign new_n9031_ = ~pi0299 & new_n7499_;
  assign new_n9032_ = ~new_n6132_ & new_n9031_;
  assign new_n9033_ = ~pi0164 & pi0186;
  assign new_n9034_ = new_n9032_ & new_n9033_;
  assign new_n9035_ = ~new_n9030_ & ~new_n9034_;
  assign new_n9036_ = pi0038 & ~new_n9035_;
  assign new_n9037_ = ~pi0176 & pi0232;
  assign new_n9038_ = ~pi0040 & new_n2476_;
  assign new_n9039_ = ~pi0102 & new_n8917_;
  assign new_n9040_ = new_n2455_ & new_n9039_;
  assign new_n9041_ = new_n2453_ & new_n9040_;
  assign new_n9042_ = new_n2474_ & new_n9041_;
  assign new_n9043_ = ~pi0060 & new_n9042_;
  assign new_n9044_ = new_n2505_ & new_n2513_;
  assign new_n9045_ = ~pi0053 & new_n9044_;
  assign new_n9046_ = new_n9043_ & new_n9045_;
  assign new_n9047_ = ~pi0058 & new_n9046_;
  assign new_n9048_ = new_n7471_ & new_n9047_;
  assign new_n9049_ = ~pi0032 & new_n2551_;
  assign new_n9050_ = new_n9048_ & new_n9049_;
  assign new_n9051_ = ~pi0095 & new_n9050_;
  assign new_n9052_ = new_n6457_ & ~new_n6469_;
  assign new_n9053_ = new_n6193_ & new_n9052_;
  assign new_n9054_ = ~new_n6224_ & ~new_n9053_;
  assign new_n9055_ = new_n9051_ & ~new_n9054_;
  assign new_n9056_ = new_n6221_ & new_n9055_;
  assign new_n9057_ = new_n9038_ & ~new_n9056_;
  assign new_n9058_ = pi0224 & new_n6480_;
  assign new_n9059_ = new_n9038_ & ~new_n9058_;
  assign new_n9060_ = ~new_n9057_ & ~new_n9059_;
  assign new_n9061_ = new_n9051_ & new_n9053_;
  assign new_n9062_ = new_n6185_ & new_n9061_;
  assign new_n9063_ = new_n9038_ & ~new_n9062_;
  assign new_n9064_ = ~new_n6238_ & ~new_n9063_;
  assign new_n9065_ = ~new_n9059_ & new_n9064_;
  assign new_n9066_ = pi0174 & new_n9065_;
  assign new_n9067_ = ~new_n9060_ & ~new_n9066_;
  assign new_n9068_ = ~pi0299 & ~new_n9067_;
  assign new_n9069_ = pi0216 & new_n6453_;
  assign new_n9070_ = new_n9038_ & ~new_n9069_;
  assign new_n9071_ = pi0299 & ~new_n9070_;
  assign new_n9072_ = new_n6224_ & new_n9051_;
  assign new_n9073_ = ~new_n6215_ & new_n9072_;
  assign new_n9074_ = new_n9038_ & ~new_n9073_;
  assign new_n9075_ = new_n6185_ & new_n9074_;
  assign new_n9076_ = ~pi0152 & new_n9075_;
  assign new_n9077_ = new_n6185_ & new_n9055_;
  assign new_n9078_ = new_n9038_ & ~new_n9077_;
  assign new_n9079_ = ~new_n6212_ & ~new_n9078_;
  assign new_n9080_ = new_n9057_ & ~new_n9079_;
  assign new_n9081_ = ~pi0154 & ~new_n9080_;
  assign new_n9082_ = ~new_n9076_ & new_n9081_;
  assign new_n9083_ = new_n9038_ & ~new_n9061_;
  assign new_n9084_ = new_n6222_ & ~new_n9083_;
  assign new_n9085_ = pi0152 & new_n9084_;
  assign new_n9086_ = new_n9057_ & ~new_n9085_;
  assign new_n9087_ = pi0154 & ~new_n9086_;
  assign new_n9088_ = new_n9069_ & ~new_n9087_;
  assign new_n9089_ = ~new_n9082_ & new_n9088_;
  assign new_n9090_ = new_n9071_ & ~new_n9089_;
  assign new_n9091_ = ~new_n9068_ & ~new_n9090_;
  assign new_n9092_ = new_n6243_ & new_n9072_;
  assign new_n9093_ = new_n9038_ & new_n9058_;
  assign new_n9094_ = ~new_n9092_ & new_n9093_;
  assign new_n9095_ = ~new_n9059_ & ~new_n9094_;
  assign new_n9096_ = ~pi0299 & new_n9095_;
  assign new_n9097_ = new_n9091_ & ~new_n9096_;
  assign new_n9098_ = new_n9037_ & ~new_n9097_;
  assign new_n9099_ = pi0176 & pi0232;
  assign new_n9100_ = ~new_n9091_ & new_n9099_;
  assign new_n9101_ = new_n9071_ & ~new_n9080_;
  assign new_n9102_ = ~new_n6238_ & ~new_n9078_;
  assign new_n9103_ = ~new_n9059_ & new_n9102_;
  assign new_n9104_ = ~new_n9060_ & ~new_n9103_;
  assign new_n9105_ = ~pi0299 & ~new_n9104_;
  assign new_n9106_ = ~new_n9101_ & ~new_n9105_;
  assign new_n9107_ = ~pi0232 & ~new_n9106_;
  assign new_n9108_ = pi0039 & ~new_n9107_;
  assign new_n9109_ = ~new_n9100_ & new_n9108_;
  assign new_n9110_ = ~new_n9098_ & new_n9109_;
  assign new_n9111_ = pi0095 & ~new_n9038_;
  assign new_n9112_ = ~new_n2449_ & ~new_n9111_;
  assign new_n9113_ = ~pi0040 & ~pi0479;
  assign new_n9114_ = new_n2476_ & ~new_n9050_;
  assign new_n9115_ = new_n9113_ & new_n9114_;
  assign new_n9116_ = ~new_n9112_ & ~new_n9115_;
  assign new_n9117_ = pi0032 & ~new_n9038_;
  assign new_n9118_ = new_n2476_ & ~new_n2549_;
  assign new_n9119_ = new_n2476_ & ~new_n9048_;
  assign new_n9120_ = pi0070 & ~new_n9119_;
  assign new_n9121_ = new_n2476_ & ~new_n9046_;
  assign new_n9122_ = pi0058 & ~new_n9121_;
  assign new_n9123_ = pi0053 & ~new_n9043_;
  assign new_n9124_ = ~pi0060 & new_n8896_;
  assign new_n9125_ = new_n2504_ & ~new_n9124_;
  assign new_n9126_ = ~new_n9123_ & ~new_n9125_;
  assign new_n9127_ = ~pi0111 & new_n2456_;
  assign new_n9128_ = ~pi0068 & new_n2457_;
  assign new_n9129_ = ~pi0036 & new_n9128_;
  assign new_n9130_ = new_n9127_ & new_n9129_;
  assign new_n9131_ = ~pi0066 & ~pi0084;
  assign new_n9132_ = pi0073 & ~pi0082;
  assign new_n9133_ = new_n9131_ & new_n9132_;
  assign new_n9134_ = new_n9130_ & new_n9133_;
  assign new_n9135_ = new_n9041_ & new_n9134_;
  assign new_n9136_ = new_n2466_ & new_n9135_;
  assign new_n9137_ = new_n2483_ & new_n9136_;
  assign new_n9138_ = new_n2476_ & ~new_n9137_;
  assign new_n9139_ = ~new_n9126_ & new_n9138_;
  assign new_n9140_ = new_n2505_ & ~new_n9139_;
  assign new_n9141_ = ~new_n2476_ & ~new_n2505_;
  assign new_n9142_ = new_n2513_ & ~new_n9141_;
  assign new_n9143_ = ~new_n9140_ & new_n9142_;
  assign new_n9144_ = new_n2476_ & ~new_n2513_;
  assign new_n9145_ = ~pi0058 & ~new_n9144_;
  assign new_n9146_ = ~new_n9143_ & new_n9145_;
  assign new_n9147_ = ~new_n9122_ & ~new_n9146_;
  assign new_n9148_ = ~pi0090 & ~new_n9147_;
  assign new_n9149_ = ~pi0841 & new_n9047_;
  assign new_n9150_ = new_n2476_ & ~new_n9149_;
  assign new_n9151_ = pi0090 & ~new_n9150_;
  assign new_n9152_ = new_n2547_ & ~new_n9151_;
  assign new_n9153_ = ~new_n9148_ & new_n9152_;
  assign new_n9154_ = new_n2476_ & ~new_n2547_;
  assign new_n9155_ = ~pi0070 & ~new_n9154_;
  assign new_n9156_ = ~new_n9153_ & new_n9155_;
  assign new_n9157_ = ~new_n9120_ & ~new_n9156_;
  assign new_n9158_ = ~pi0051 & ~new_n9157_;
  assign new_n9159_ = pi0051 & ~new_n2476_;
  assign new_n9160_ = new_n2549_ & ~new_n9159_;
  assign new_n9161_ = ~new_n9158_ & new_n9160_;
  assign new_n9162_ = ~new_n9118_ & ~new_n9161_;
  assign new_n9163_ = ~pi0040 & ~new_n9162_;
  assign new_n9164_ = ~pi0032 & ~new_n9163_;
  assign new_n9165_ = ~new_n9117_ & ~new_n9164_;
  assign new_n9166_ = ~pi0095 & ~new_n9165_;
  assign new_n9167_ = ~new_n9116_ & ~new_n9166_;
  assign new_n9168_ = ~pi0072 & ~pi0093;
  assign new_n9169_ = new_n2496_ & new_n9168_;
  assign new_n9170_ = ~pi0090 & new_n9169_;
  assign new_n9171_ = new_n9149_ & new_n9170_;
  assign new_n9172_ = new_n9038_ & ~new_n9171_;
  assign new_n9173_ = pi0032 & ~new_n9172_;
  assign new_n9174_ = ~new_n9164_ & ~new_n9173_;
  assign new_n9175_ = ~pi0095 & ~new_n9174_;
  assign new_n9176_ = ~pi0198 & new_n9175_;
  assign new_n9177_ = new_n9167_ & ~new_n9176_;
  assign new_n9178_ = ~new_n6185_ & new_n9177_;
  assign new_n9179_ = new_n9044_ & new_n9126_;
  assign new_n9180_ = new_n2476_ & ~new_n9179_;
  assign new_n9181_ = ~pi0058 & ~new_n9180_;
  assign new_n9182_ = ~new_n9122_ & ~new_n9181_;
  assign new_n9183_ = ~pi0090 & ~new_n9182_;
  assign new_n9184_ = new_n9152_ & ~new_n9183_;
  assign new_n9185_ = new_n9155_ & ~new_n9184_;
  assign new_n9186_ = ~new_n9120_ & ~new_n9185_;
  assign new_n9187_ = ~pi0051 & ~new_n9186_;
  assign new_n9188_ = new_n9160_ & ~new_n9187_;
  assign new_n9189_ = ~new_n9118_ & ~new_n9188_;
  assign new_n9190_ = ~pi0040 & ~new_n9189_;
  assign new_n9191_ = ~pi0032 & ~new_n9190_;
  assign new_n9192_ = ~new_n9173_ & ~new_n9191_;
  assign new_n9193_ = ~pi0095 & ~new_n9192_;
  assign new_n9194_ = ~pi0198 & new_n9193_;
  assign new_n9195_ = new_n6185_ & ~new_n9111_;
  assign new_n9196_ = ~new_n9117_ & ~new_n9191_;
  assign new_n9197_ = ~pi0095 & ~new_n9196_;
  assign new_n9198_ = new_n9195_ & ~new_n9197_;
  assign new_n9199_ = ~new_n9194_ & new_n9198_;
  assign new_n9200_ = ~new_n9178_ & ~new_n9199_;
  assign new_n9201_ = ~pi0183 & ~new_n9200_;
  assign new_n9202_ = ~pi0040 & ~new_n9117_;
  assign new_n9203_ = new_n2476_ & ~new_n6167_;
  assign new_n9204_ = ~pi0032 & ~new_n9203_;
  assign new_n9205_ = pi0093 & ~new_n2476_;
  assign new_n9206_ = new_n6167_ & ~new_n9205_;
  assign new_n9207_ = new_n2476_ & ~new_n9122_;
  assign new_n9208_ = ~pi0090 & ~new_n9207_;
  assign new_n9209_ = ~new_n9151_ & ~new_n9208_;
  assign new_n9210_ = ~pi0093 & ~new_n9209_;
  assign new_n9211_ = new_n9206_ & ~new_n9210_;
  assign new_n9212_ = new_n9204_ & ~new_n9211_;
  assign new_n9213_ = new_n9202_ & ~new_n9212_;
  assign new_n9214_ = ~pi0095 & ~new_n9213_;
  assign new_n9215_ = new_n9195_ & ~new_n9214_;
  assign new_n9216_ = ~new_n9178_ & ~new_n9215_;
  assign new_n9217_ = pi0183 & ~new_n9216_;
  assign new_n9218_ = ~new_n9201_ & ~new_n9217_;
  assign new_n9219_ = ~pi0095 & new_n9218_;
  assign new_n9220_ = ~pi0174 & ~new_n9116_;
  assign new_n9221_ = ~new_n9219_ & new_n9220_;
  assign new_n9222_ = pi0183 & new_n6185_;
  assign new_n9223_ = ~new_n9177_ & ~new_n9222_;
  assign new_n9224_ = new_n8932_ & new_n9136_;
  assign new_n9225_ = ~pi0090 & new_n9224_;
  assign new_n9226_ = new_n9209_ & ~new_n9225_;
  assign new_n9227_ = ~pi0093 & ~new_n9226_;
  assign new_n9228_ = new_n9206_ & ~new_n9227_;
  assign new_n9229_ = new_n9204_ & ~new_n9228_;
  assign new_n9230_ = new_n9202_ & ~new_n9229_;
  assign new_n9231_ = ~pi0095 & ~new_n9230_;
  assign new_n9232_ = ~new_n9116_ & ~new_n9231_;
  assign new_n9233_ = new_n6185_ & ~new_n9232_;
  assign new_n9234_ = pi0183 & new_n9233_;
  assign new_n9235_ = pi0174 & ~new_n9234_;
  assign new_n9236_ = ~new_n9223_ & new_n9235_;
  assign new_n9237_ = ~pi0180 & ~new_n9236_;
  assign new_n9238_ = ~new_n9221_ & new_n9237_;
  assign new_n9239_ = new_n9195_ & ~new_n9231_;
  assign new_n9240_ = ~new_n9178_ & ~new_n9239_;
  assign new_n9241_ = pi0183 & ~new_n9240_;
  assign new_n9242_ = ~pi0040 & new_n6185_;
  assign new_n9243_ = ~new_n9111_ & ~new_n9166_;
  assign new_n9244_ = ~new_n9176_ & new_n9243_;
  assign new_n9245_ = new_n9242_ & new_n9244_;
  assign new_n9246_ = ~new_n9178_ & ~new_n9245_;
  assign new_n9247_ = ~pi0183 & ~new_n9246_;
  assign new_n9248_ = ~new_n9241_ & ~new_n9247_;
  assign new_n9249_ = pi0174 & ~new_n9248_;
  assign new_n9250_ = ~pi0174 & ~new_n9218_;
  assign new_n9251_ = pi0180 & ~new_n9250_;
  assign new_n9252_ = ~new_n9249_ & new_n9251_;
  assign new_n9253_ = ~new_n9238_ & ~new_n9252_;
  assign new_n9254_ = ~pi0193 & ~new_n9253_;
  assign new_n9255_ = ~pi0040 & ~new_n2476_;
  assign new_n9256_ = pi0095 & ~new_n9255_;
  assign new_n9257_ = pi0032 & ~new_n9255_;
  assign new_n9258_ = new_n2518_ & new_n2547_;
  assign new_n9259_ = ~new_n2476_ & ~new_n9258_;
  assign new_n9260_ = new_n7471_ & new_n9181_;
  assign new_n9261_ = ~new_n9259_ & ~new_n9260_;
  assign new_n9262_ = ~pi0070 & ~new_n9261_;
  assign new_n9263_ = ~new_n9120_ & ~new_n9262_;
  assign new_n9264_ = ~pi0051 & ~new_n9263_;
  assign new_n9265_ = new_n9160_ & ~new_n9264_;
  assign new_n9266_ = ~new_n9118_ & ~new_n9265_;
  assign new_n9267_ = ~pi0040 & new_n9266_;
  assign new_n9268_ = ~pi0032 & ~new_n9267_;
  assign new_n9269_ = ~new_n9257_ & ~new_n9268_;
  assign new_n9270_ = ~pi0095 & ~new_n9269_;
  assign new_n9271_ = ~new_n9256_ & ~new_n9270_;
  assign new_n9272_ = pi0198 & ~new_n9271_;
  assign new_n9273_ = ~pi0040 & ~new_n9172_;
  assign new_n9274_ = pi0032 & ~new_n9273_;
  assign new_n9275_ = ~new_n9268_ & ~new_n9274_;
  assign new_n9276_ = ~pi0095 & ~new_n9275_;
  assign new_n9277_ = ~new_n9256_ & ~new_n9276_;
  assign new_n9278_ = ~pi0198 & ~new_n9277_;
  assign new_n9279_ = ~new_n9272_ & ~new_n9278_;
  assign new_n9280_ = new_n9242_ & ~new_n9279_;
  assign new_n9281_ = ~new_n9178_ & ~new_n9280_;
  assign new_n9282_ = ~pi0183 & ~new_n9281_;
  assign new_n9283_ = new_n6185_ & ~new_n9038_;
  assign new_n9284_ = ~new_n6185_ & ~new_n9177_;
  assign new_n9285_ = ~new_n9283_ & ~new_n9284_;
  assign new_n9286_ = pi0183 & new_n9285_;
  assign new_n9287_ = ~pi0174 & ~new_n9286_;
  assign new_n9288_ = ~new_n9282_ & new_n9287_;
  assign new_n9289_ = new_n7471_ & new_n9146_;
  assign new_n9290_ = ~new_n9259_ & ~new_n9289_;
  assign new_n9291_ = ~pi0070 & ~new_n9290_;
  assign new_n9292_ = ~new_n9120_ & ~new_n9291_;
  assign new_n9293_ = ~pi0051 & ~new_n9292_;
  assign new_n9294_ = new_n9160_ & ~new_n9293_;
  assign new_n9295_ = ~pi0040 & ~new_n9118_;
  assign new_n9296_ = ~new_n9294_ & new_n9295_;
  assign new_n9297_ = ~pi0032 & ~new_n9296_;
  assign new_n9298_ = ~new_n9257_ & ~new_n9297_;
  assign new_n9299_ = ~new_n2782_ & ~new_n9038_;
  assign new_n9300_ = ~new_n9298_ & ~new_n9299_;
  assign new_n9301_ = ~pi0095 & ~new_n9300_;
  assign new_n9302_ = ~new_n9111_ & ~new_n9301_;
  assign new_n9303_ = ~new_n9274_ & ~new_n9297_;
  assign new_n9304_ = ~pi0095 & ~new_n9303_;
  assign new_n9305_ = ~new_n9256_ & ~new_n9304_;
  assign new_n9306_ = new_n9302_ & ~new_n9305_;
  assign new_n9307_ = ~pi0198 & ~new_n9306_;
  assign new_n9308_ = new_n6185_ & ~new_n9307_;
  assign new_n9309_ = new_n9302_ & new_n9308_;
  assign new_n9310_ = ~new_n9178_ & ~new_n9309_;
  assign new_n9311_ = ~pi0183 & ~new_n9310_;
  assign new_n9312_ = new_n2493_ & new_n6167_;
  assign new_n9313_ = new_n8932_ & new_n9312_;
  assign new_n9314_ = ~pi0032 & new_n9313_;
  assign new_n9315_ = new_n9136_ & new_n9314_;
  assign new_n9316_ = new_n9038_ & ~new_n9315_;
  assign new_n9317_ = ~pi0095 & ~new_n9316_;
  assign new_n9318_ = new_n9195_ & ~new_n9317_;
  assign new_n9319_ = ~new_n9178_ & ~new_n9318_;
  assign new_n9320_ = pi0183 & ~new_n9319_;
  assign new_n9321_ = pi0174 & ~new_n9320_;
  assign new_n9322_ = ~new_n9311_ & new_n9321_;
  assign new_n9323_ = pi0180 & ~new_n9322_;
  assign new_n9324_ = ~new_n9288_ & new_n9323_;
  assign new_n9325_ = ~new_n9116_ & ~new_n9301_;
  assign new_n9326_ = ~new_n9283_ & ~new_n9308_;
  assign new_n9327_ = new_n9325_ & ~new_n9326_;
  assign new_n9328_ = ~new_n9178_ & ~new_n9327_;
  assign new_n9329_ = ~pi0183 & ~new_n9328_;
  assign new_n9330_ = new_n6185_ & ~new_n9317_;
  assign new_n9331_ = ~new_n9116_ & new_n9330_;
  assign new_n9332_ = ~new_n9178_ & ~new_n9331_;
  assign new_n9333_ = pi0183 & ~new_n9332_;
  assign new_n9334_ = pi0174 & ~new_n9333_;
  assign new_n9335_ = ~new_n9329_ & new_n9334_;
  assign new_n9336_ = ~pi0095 & ~new_n9038_;
  assign new_n9337_ = ~new_n9116_ & ~new_n9336_;
  assign new_n9338_ = new_n6185_ & new_n9337_;
  assign new_n9339_ = ~new_n9178_ & ~new_n9338_;
  assign new_n9340_ = pi0183 & ~new_n9339_;
  assign new_n9341_ = ~pi0040 & ~new_n9266_;
  assign new_n9342_ = ~pi0032 & ~new_n9341_;
  assign new_n9343_ = ~new_n9117_ & ~new_n9342_;
  assign new_n9344_ = ~pi0095 & ~new_n9343_;
  assign new_n9345_ = ~new_n9116_ & ~new_n9344_;
  assign new_n9346_ = ~new_n9173_ & ~new_n9342_;
  assign new_n9347_ = ~pi0095 & ~new_n9346_;
  assign new_n9348_ = ~pi0198 & new_n9347_;
  assign new_n9349_ = new_n9345_ & ~new_n9348_;
  assign new_n9350_ = new_n6185_ & ~new_n9349_;
  assign new_n9351_ = ~new_n9284_ & ~new_n9350_;
  assign new_n9352_ = ~pi0183 & new_n9351_;
  assign new_n9353_ = ~pi0174 & ~new_n9352_;
  assign new_n9354_ = ~new_n9340_ & new_n9353_;
  assign new_n9355_ = ~pi0180 & ~new_n9354_;
  assign new_n9356_ = ~new_n9335_ & new_n9355_;
  assign new_n9357_ = pi0193 & ~new_n9356_;
  assign new_n9358_ = ~new_n9324_ & new_n9357_;
  assign new_n9359_ = ~new_n9254_ & ~new_n9358_;
  assign new_n9360_ = ~pi0299 & ~new_n9359_;
  assign new_n9361_ = pi0158 & pi0299;
  assign new_n9362_ = ~pi0210 & new_n9175_;
  assign new_n9363_ = new_n9167_ & ~new_n9362_;
  assign new_n9364_ = ~new_n6185_ & ~new_n9363_;
  assign new_n9365_ = new_n9243_ & ~new_n9362_;
  assign new_n9366_ = new_n6185_ & ~new_n9365_;
  assign new_n9367_ = ~new_n9364_ & ~new_n9366_;
  assign new_n9368_ = pi0152 & new_n9367_;
  assign new_n9369_ = ~new_n6185_ & new_n9363_;
  assign new_n9370_ = ~pi0210 & new_n9193_;
  assign new_n9371_ = new_n9198_ & ~new_n9370_;
  assign new_n9372_ = ~new_n9369_ & ~new_n9371_;
  assign new_n9373_ = ~pi0152 & ~new_n9372_;
  assign new_n9374_ = ~pi0172 & ~new_n9373_;
  assign new_n9375_ = ~new_n9368_ & new_n9374_;
  assign new_n9376_ = ~pi0210 & ~new_n9306_;
  assign new_n9377_ = new_n6185_ & ~new_n9376_;
  assign new_n9378_ = new_n9302_ & new_n9377_;
  assign new_n9379_ = ~new_n9369_ & ~new_n9378_;
  assign new_n9380_ = pi0152 & ~new_n9379_;
  assign new_n9381_ = ~new_n9111_ & ~new_n9347_;
  assign new_n9382_ = ~pi0210 & ~new_n9381_;
  assign new_n9383_ = new_n6185_ & ~new_n9382_;
  assign new_n9384_ = ~new_n9111_ & ~new_n9344_;
  assign new_n9385_ = new_n9383_ & new_n9384_;
  assign new_n9386_ = ~new_n9369_ & ~new_n9385_;
  assign new_n9387_ = ~pi0152 & ~new_n9386_;
  assign new_n9388_ = pi0172 & ~new_n9387_;
  assign new_n9389_ = ~new_n9380_ & new_n9388_;
  assign new_n9390_ = ~new_n9375_ & ~new_n9389_;
  assign new_n9391_ = new_n9361_ & ~new_n9390_;
  assign new_n9392_ = ~new_n9283_ & ~new_n9377_;
  assign new_n9393_ = new_n9325_ & ~new_n9392_;
  assign new_n9394_ = pi0152 & ~new_n9393_;
  assign new_n9395_ = ~new_n9283_ & ~new_n9383_;
  assign new_n9396_ = new_n9345_ & ~new_n9395_;
  assign new_n9397_ = ~pi0152 & ~new_n9396_;
  assign new_n9398_ = pi0172 & ~new_n9397_;
  assign new_n9399_ = ~new_n9394_ & new_n9398_;
  assign new_n9400_ = pi0152 & ~new_n9363_;
  assign new_n9401_ = ~new_n9116_ & ~new_n9197_;
  assign new_n9402_ = ~new_n9370_ & new_n9401_;
  assign new_n9403_ = new_n6185_ & new_n9402_;
  assign new_n9404_ = ~pi0152 & ~new_n9403_;
  assign new_n9405_ = ~pi0172 & ~new_n9404_;
  assign new_n9406_ = ~new_n9400_ & new_n9405_;
  assign new_n9407_ = ~pi0158 & pi0299;
  assign new_n9408_ = ~new_n9369_ & new_n9407_;
  assign new_n9409_ = ~new_n9406_ & new_n9408_;
  assign new_n9410_ = ~new_n9399_ & new_n9409_;
  assign new_n9411_ = ~pi0149 & ~new_n9410_;
  assign new_n9412_ = ~new_n9391_ & new_n9411_;
  assign new_n9413_ = ~new_n9338_ & ~new_n9369_;
  assign new_n9414_ = ~pi0152 & ~new_n9413_;
  assign new_n9415_ = ~new_n9331_ & ~new_n9369_;
  assign new_n9416_ = pi0152 & ~new_n9415_;
  assign new_n9417_ = pi0172 & ~new_n9416_;
  assign new_n9418_ = ~new_n9414_ & new_n9417_;
  assign new_n9419_ = ~new_n9233_ & ~new_n9364_;
  assign new_n9420_ = pi0152 & new_n9419_;
  assign new_n9421_ = ~new_n9116_ & ~new_n9214_;
  assign new_n9422_ = new_n6185_ & ~new_n9421_;
  assign new_n9423_ = ~new_n9364_ & ~new_n9422_;
  assign new_n9424_ = ~pi0152 & new_n9423_;
  assign new_n9425_ = ~pi0172 & ~new_n9424_;
  assign new_n9426_ = ~new_n9420_ & new_n9425_;
  assign new_n9427_ = ~new_n9418_ & ~new_n9426_;
  assign new_n9428_ = new_n9407_ & ~new_n9427_;
  assign new_n9429_ = ~new_n9215_ & ~new_n9369_;
  assign new_n9430_ = ~pi0152 & ~new_n9429_;
  assign new_n9431_ = ~new_n9239_ & ~new_n9369_;
  assign new_n9432_ = pi0152 & ~new_n9431_;
  assign new_n9433_ = ~pi0172 & ~new_n9432_;
  assign new_n9434_ = ~new_n9430_ & new_n9433_;
  assign new_n9435_ = ~new_n9283_ & ~new_n9364_;
  assign new_n9436_ = ~pi0152 & new_n9435_;
  assign new_n9437_ = ~new_n9318_ & ~new_n9369_;
  assign new_n9438_ = pi0152 & ~new_n9437_;
  assign new_n9439_ = pi0172 & ~new_n9438_;
  assign new_n9440_ = ~new_n9436_ & new_n9439_;
  assign new_n9441_ = ~new_n9434_ & ~new_n9440_;
  assign new_n9442_ = new_n9361_ & ~new_n9441_;
  assign new_n9443_ = pi0149 & ~new_n9442_;
  assign new_n9444_ = ~new_n9428_ & new_n9443_;
  assign new_n9445_ = ~new_n9412_ & ~new_n9444_;
  assign new_n9446_ = ~new_n9360_ & ~new_n9445_;
  assign new_n9447_ = pi0232 & ~new_n9446_;
  assign new_n9448_ = ~new_n6166_ & new_n9175_;
  assign new_n9449_ = new_n9167_ & ~new_n9448_;
  assign new_n9450_ = ~pi0232 & ~new_n9449_;
  assign new_n9451_ = ~pi0039 & ~new_n9450_;
  assign new_n9452_ = ~new_n9447_ & new_n9451_;
  assign new_n9453_ = ~new_n9110_ & ~new_n9452_;
  assign new_n9454_ = ~pi0038 & ~new_n9453_;
  assign new_n9455_ = ~new_n9036_ & ~new_n9454_;
  assign new_n9456_ = ~pi0100 & ~new_n9455_;
  assign new_n9457_ = ~pi0087 & ~new_n9007_;
  assign new_n9458_ = ~new_n9456_ & new_n9457_;
  assign new_n9459_ = pi0038 & new_n9020_;
  assign new_n9460_ = ~pi0100 & new_n9459_;
  assign new_n9461_ = ~new_n9007_ & ~new_n9460_;
  assign new_n9462_ = new_n3211_ & new_n9038_;
  assign new_n9463_ = pi0087 & ~new_n9462_;
  assign new_n9464_ = new_n9461_ & new_n9463_;
  assign new_n9465_ = new_n3242_ & ~new_n9464_;
  assign new_n9466_ = ~new_n9458_ & new_n9465_;
  assign new_n9467_ = ~pi0075 & pi0092;
  assign new_n9468_ = pi0232 & ~new_n3398_;
  assign new_n9469_ = ~pi0176 & ~pi0299;
  assign new_n9470_ = new_n6185_ & ~new_n9469_;
  assign new_n9471_ = new_n9468_ & new_n9470_;
  assign new_n9472_ = new_n3226_ & new_n9051_;
  assign new_n9473_ = ~new_n9471_ & new_n9472_;
  assign new_n9474_ = new_n9462_ & ~new_n9473_;
  assign new_n9475_ = new_n9461_ & ~new_n9474_;
  assign new_n9476_ = new_n9467_ & ~new_n9475_;
  assign new_n9477_ = ~new_n9008_ & ~new_n9476_;
  assign new_n9478_ = ~new_n9466_ & new_n9477_;
  assign new_n9479_ = ~pi0054 & ~new_n9478_;
  assign new_n9480_ = ~new_n9023_ & ~new_n9479_;
  assign new_n9481_ = ~pi0074 & ~new_n9480_;
  assign new_n9482_ = new_n9016_ & ~new_n9481_;
  assign new_n9483_ = pi0055 & ~new_n8993_;
  assign new_n9484_ = pi0054 & ~new_n8995_;
  assign new_n9485_ = ~pi0092 & ~new_n8986_;
  assign new_n9486_ = pi0164 & new_n7499_;
  assign new_n9487_ = pi0038 & ~new_n9486_;
  assign new_n9488_ = new_n3245_ & ~new_n9487_;
  assign new_n9489_ = pi0149 & new_n7499_;
  assign new_n9490_ = ~pi0039 & ~new_n9489_;
  assign new_n9491_ = new_n9051_ & new_n9490_;
  assign new_n9492_ = new_n9038_ & ~new_n9491_;
  assign new_n9493_ = ~pi0038 & ~new_n9492_;
  assign new_n9494_ = new_n9488_ & ~new_n9493_;
  assign new_n9495_ = ~pi0038 & ~new_n9038_;
  assign new_n9496_ = ~pi0100 & ~new_n9495_;
  assign new_n9497_ = ~new_n9487_ & new_n9496_;
  assign new_n9498_ = pi0087 & new_n9497_;
  assign new_n9499_ = ~new_n8987_ & ~new_n9498_;
  assign new_n9500_ = ~new_n9494_ & new_n9499_;
  assign new_n9501_ = ~pi0075 & ~new_n9500_;
  assign new_n9502_ = new_n9485_ & ~new_n9501_;
  assign new_n9503_ = ~pi0075 & new_n9497_;
  assign new_n9504_ = pi0092 & new_n8988_;
  assign new_n9505_ = ~new_n9503_ & new_n9504_;
  assign new_n9506_ = ~pi0054 & ~new_n9505_;
  assign new_n9507_ = ~new_n9502_ & new_n9506_;
  assign new_n9508_ = ~new_n9484_ & ~new_n9507_;
  assign new_n9509_ = ~pi0074 & ~new_n9508_;
  assign new_n9510_ = new_n9483_ & ~new_n9509_;
  assign new_n9511_ = new_n3298_ & ~new_n9510_;
  assign new_n9512_ = ~new_n9482_ & new_n9511_;
  assign new_n9513_ = pi0038 & new_n9486_;
  assign new_n9514_ = new_n8989_ & new_n9513_;
  assign new_n9515_ = new_n8988_ & ~new_n9514_;
  assign new_n9516_ = ~new_n9484_ & new_n9515_;
  assign new_n9517_ = ~pi0074 & ~new_n9516_;
  assign new_n9518_ = ~new_n8993_ & ~new_n9517_;
  assign new_n9519_ = ~new_n3298_ & ~new_n9518_;
  assign new_n9520_ = new_n3436_ & ~new_n9519_;
  assign new_n9521_ = ~pi0038 & new_n9038_;
  assign new_n9522_ = new_n8989_ & new_n9521_;
  assign new_n9523_ = new_n3270_ & new_n9522_;
  assign new_n9524_ = ~new_n3298_ & new_n9523_;
  assign new_n9525_ = new_n9520_ & ~new_n9524_;
  assign new_n9526_ = ~new_n9512_ & new_n9525_;
  assign new_n9527_ = ~new_n8998_ & ~new_n9526_;
  assign new_n9528_ = ~new_n8980_ & ~new_n9527_;
  assign new_n9529_ = new_n6243_ & new_n6470_;
  assign new_n9530_ = new_n9058_ & new_n9529_;
  assign new_n9531_ = ~pi0174 & new_n9530_;
  assign new_n9532_ = ~pi0299 & ~new_n9531_;
  assign new_n9533_ = new_n9037_ & ~new_n9532_;
  assign new_n9534_ = ~new_n6466_ & new_n9058_;
  assign new_n9535_ = new_n6243_ & new_n9534_;
  assign new_n9536_ = ~pi0174 & new_n9535_;
  assign new_n9537_ = new_n6243_ & new_n9058_;
  assign new_n9538_ = new_n7544_ & new_n9537_;
  assign new_n9539_ = pi0174 & new_n9538_;
  assign new_n9540_ = ~pi0299 & ~new_n9539_;
  assign new_n9541_ = ~new_n9536_ & new_n9540_;
  assign new_n9542_ = new_n9099_ & ~new_n9541_;
  assign new_n9543_ = ~new_n9533_ & ~new_n9542_;
  assign new_n9544_ = new_n6222_ & ~new_n6466_;
  assign new_n9545_ = pi0154 & ~new_n9544_;
  assign new_n9546_ = new_n6222_ & new_n6470_;
  assign new_n9547_ = ~pi0154 & ~new_n9546_;
  assign new_n9548_ = ~pi0152 & ~new_n9547_;
  assign new_n9549_ = ~new_n9545_ & new_n9548_;
  assign new_n9550_ = new_n6185_ & new_n7544_;
  assign new_n9551_ = ~new_n6212_ & new_n9550_;
  assign new_n9552_ = pi0152 & pi0154;
  assign new_n9553_ = new_n9551_ & new_n9552_;
  assign new_n9554_ = ~new_n9549_ & ~new_n9553_;
  assign new_n9555_ = new_n9069_ & ~new_n9554_;
  assign new_n9556_ = pi0299 & ~new_n9555_;
  assign new_n9557_ = pi0039 & ~new_n9556_;
  assign new_n9558_ = ~new_n9543_ & new_n9557_;
  assign new_n9559_ = pi0090 & ~new_n7458_;
  assign new_n9560_ = new_n2547_ & ~new_n6136_;
  assign new_n9561_ = ~new_n9559_ & new_n9560_;
  assign new_n9562_ = ~pi0090 & new_n2514_;
  assign new_n9563_ = new_n2547_ & new_n9562_;
  assign new_n9564_ = new_n2508_ & new_n9563_;
  assign new_n9565_ = new_n2476_ & new_n9564_;
  assign new_n9566_ = new_n9140_ & new_n9565_;
  assign new_n9567_ = ~pi0070 & ~new_n9566_;
  assign new_n9568_ = ~new_n9561_ & new_n9567_;
  assign new_n9569_ = new_n2849_ & new_n3098_;
  assign new_n9570_ = ~new_n9568_ & new_n9569_;
  assign new_n9571_ = ~new_n9567_ & new_n9569_;
  assign new_n9572_ = ~new_n6387_ & ~new_n9571_;
  assign new_n9573_ = ~pi0198 & ~new_n9572_;
  assign new_n9574_ = ~new_n9570_ & ~new_n9573_;
  assign new_n9575_ = new_n9222_ & ~new_n9574_;
  assign new_n9576_ = new_n9169_ & ~new_n9559_;
  assign new_n9577_ = new_n2476_ & new_n9224_;
  assign new_n9578_ = new_n6136_ & ~new_n9577_;
  assign new_n9579_ = new_n9576_ & ~new_n9578_;
  assign new_n9580_ = new_n3097_ & new_n6185_;
  assign new_n9581_ = ~pi0040 & new_n9580_;
  assign new_n9582_ = new_n9579_ & new_n9581_;
  assign new_n9583_ = ~pi0183 & new_n9582_;
  assign new_n9584_ = ~pi0174 & ~new_n9583_;
  assign new_n9585_ = ~new_n9575_ & new_n9584_;
  assign new_n9586_ = ~new_n9125_ & new_n9564_;
  assign new_n9587_ = ~pi0070 & ~new_n9586_;
  assign new_n9588_ = ~new_n9561_ & new_n9587_;
  assign new_n9589_ = new_n9569_ & ~new_n9588_;
  assign new_n9590_ = ~new_n6388_ & ~new_n9589_;
  assign new_n9591_ = new_n6185_ & ~new_n9590_;
  assign new_n9592_ = pi0183 & new_n9591_;
  assign new_n9593_ = ~new_n6136_ & new_n9576_;
  assign new_n9594_ = new_n9581_ & new_n9593_;
  assign new_n9595_ = ~pi0183 & new_n9594_;
  assign new_n9596_ = pi0174 & ~new_n9595_;
  assign new_n9597_ = ~new_n9592_ & new_n9596_;
  assign new_n9598_ = ~new_n9585_ & ~new_n9597_;
  assign new_n9599_ = pi0193 & ~new_n9598_;
  assign new_n9600_ = ~new_n6388_ & ~new_n9571_;
  assign new_n9601_ = ~pi0174 & new_n9600_;
  assign new_n9602_ = new_n9569_ & ~new_n9587_;
  assign new_n9603_ = ~new_n6388_ & ~new_n9602_;
  assign new_n9604_ = pi0174 & new_n9603_;
  assign new_n9605_ = new_n9222_ & ~new_n9604_;
  assign new_n9606_ = ~new_n9601_ & new_n9605_;
  assign new_n9607_ = new_n9170_ & new_n9577_;
  assign new_n9608_ = new_n3097_ & new_n9607_;
  assign new_n9609_ = new_n9242_ & new_n9608_;
  assign new_n9610_ = ~pi0174 & ~pi0183;
  assign new_n9611_ = new_n9609_ & new_n9610_;
  assign new_n9612_ = ~pi0193 & ~new_n9611_;
  assign new_n9613_ = ~new_n9606_ & new_n9612_;
  assign new_n9614_ = ~new_n9599_ & ~new_n9613_;
  assign new_n9615_ = new_n2943_ & new_n6185_;
  assign new_n9616_ = pi0180 & new_n9615_;
  assign new_n9617_ = ~pi0299 & ~new_n9616_;
  assign new_n9618_ = ~new_n9614_ & new_n9617_;
  assign new_n9619_ = ~pi0039 & pi0232;
  assign new_n9620_ = pi0172 & new_n9570_;
  assign new_n9621_ = ~new_n6432_ & ~new_n9571_;
  assign new_n9622_ = ~pi0152 & new_n9621_;
  assign new_n9623_ = ~new_n9620_ & new_n9622_;
  assign new_n9624_ = ~new_n6432_ & ~new_n9602_;
  assign new_n9625_ = pi0172 & new_n9589_;
  assign new_n9626_ = pi0152 & ~new_n9625_;
  assign new_n9627_ = new_n9624_ & new_n9626_;
  assign new_n9628_ = pi0149 & new_n6185_;
  assign new_n9629_ = ~new_n9627_ & new_n9628_;
  assign new_n9630_ = ~new_n9623_ & new_n9629_;
  assign new_n9631_ = ~pi0152 & new_n9582_;
  assign new_n9632_ = ~new_n9594_ & ~new_n9631_;
  assign new_n9633_ = pi0172 & ~new_n9632_;
  assign new_n9634_ = ~pi0152 & ~pi0172;
  assign new_n9635_ = new_n9609_ & new_n9634_;
  assign new_n9636_ = ~new_n9633_ & ~new_n9635_;
  assign new_n9637_ = ~pi0149 & ~new_n9636_;
  assign new_n9638_ = pi0158 & new_n9615_;
  assign new_n9639_ = pi0299 & ~new_n9638_;
  assign new_n9640_ = ~new_n9637_ & new_n9639_;
  assign new_n9641_ = ~new_n9630_ & new_n9640_;
  assign new_n9642_ = new_n9619_ & ~new_n9641_;
  assign new_n9643_ = ~new_n9618_ & new_n9642_;
  assign new_n9644_ = ~new_n9558_ & ~new_n9643_;
  assign new_n9645_ = ~pi0038 & ~new_n9644_;
  assign new_n9646_ = ~pi0087 & ~new_n9036_;
  assign new_n9647_ = ~new_n9645_ & new_n9646_;
  assign new_n9648_ = pi0087 & ~new_n9459_;
  assign new_n9649_ = ~pi0100 & ~new_n9648_;
  assign new_n9650_ = ~new_n9647_ & new_n9649_;
  assign new_n9651_ = ~new_n9007_ & ~new_n9650_;
  assign new_n9652_ = new_n3242_ & ~new_n9651_;
  assign new_n9653_ = ~pi0038 & ~pi0087;
  assign new_n9654_ = ~pi0100 & new_n9653_;
  assign new_n9655_ = new_n9471_ & new_n9654_;
  assign new_n9656_ = new_n6132_ & new_n9655_;
  assign new_n9657_ = new_n9461_ & ~new_n9656_;
  assign new_n9658_ = new_n9467_ & ~new_n9657_;
  assign new_n9659_ = ~new_n9008_ & ~new_n9658_;
  assign new_n9660_ = ~new_n9652_ & new_n9659_;
  assign new_n9661_ = ~pi0054 & ~new_n9660_;
  assign new_n9662_ = ~new_n9023_ & ~new_n9661_;
  assign new_n9663_ = ~pi0074 & ~new_n9662_;
  assign new_n9664_ = new_n9016_ & ~new_n9663_;
  assign new_n9665_ = new_n6132_ & new_n9489_;
  assign new_n9666_ = ~pi0038 & ~new_n9665_;
  assign new_n9667_ = new_n9488_ & ~new_n9666_;
  assign new_n9668_ = new_n7613_ & new_n9513_;
  assign new_n9669_ = ~new_n8987_ & ~new_n9668_;
  assign new_n9670_ = ~new_n9667_ & new_n9669_;
  assign new_n9671_ = ~pi0075 & ~new_n9670_;
  assign new_n9672_ = new_n9485_ & ~new_n9671_;
  assign new_n9673_ = pi0092 & new_n9515_;
  assign new_n9674_ = ~pi0054 & ~new_n9673_;
  assign new_n9675_ = ~new_n9672_ & new_n9674_;
  assign new_n9676_ = ~new_n9484_ & ~new_n9675_;
  assign new_n9677_ = ~pi0074 & ~new_n9676_;
  assign new_n9678_ = new_n9483_ & ~new_n9677_;
  assign new_n9679_ = new_n3298_ & ~new_n9678_;
  assign new_n9680_ = ~new_n9664_ & new_n9679_;
  assign new_n9681_ = new_n9520_ & ~new_n9680_;
  assign new_n9682_ = ~new_n8998_ & ~new_n9681_;
  assign new_n9683_ = new_n8980_ & ~new_n9682_;
  assign new_n9684_ = ~pi0954 & ~new_n9683_;
  assign new_n9685_ = ~new_n9528_ & new_n9684_;
  assign new_n9686_ = ~pi0033 & ~new_n9527_;
  assign new_n9687_ = pi0033 & ~new_n9682_;
  assign new_n9688_ = pi0954 & ~new_n9687_;
  assign new_n9689_ = ~new_n9686_ & new_n9688_;
  assign po0191 = ~new_n9685_ & ~new_n9689_;
  assign new_n9691_ = pi0197 & new_n8982_;
  assign new_n9692_ = ~pi0197 & ~new_n8982_;
  assign new_n9693_ = ~new_n9691_ & ~new_n9692_;
  assign new_n9694_ = pi0162 & new_n6185_;
  assign new_n9695_ = new_n9693_ & ~new_n9694_;
  assign new_n9696_ = new_n9691_ & new_n9694_;
  assign new_n9697_ = ~pi0162 & ~pi0197;
  assign new_n9698_ = new_n8983_ & ~new_n9697_;
  assign new_n9699_ = new_n6185_ & ~new_n9698_;
  assign new_n9700_ = ~new_n9696_ & new_n9699_;
  assign new_n9701_ = ~new_n9693_ & ~new_n9700_;
  assign new_n9702_ = ~new_n9695_ & ~new_n9701_;
  assign new_n9703_ = pi0232 & new_n9702_;
  assign new_n9704_ = ~new_n8989_ & new_n9703_;
  assign new_n9705_ = pi0167 & new_n7499_;
  assign new_n9706_ = new_n8989_ & new_n9705_;
  assign new_n9707_ = ~new_n9704_ & ~new_n9706_;
  assign new_n9708_ = ~pi0074 & new_n9707_;
  assign new_n9709_ = pi0148 & new_n8990_;
  assign new_n9710_ = pi0074 & ~new_n9709_;
  assign new_n9711_ = ~new_n9704_ & new_n9710_;
  assign new_n9712_ = ~new_n9708_ & ~new_n9711_;
  assign new_n9713_ = ~new_n3436_ & new_n9712_;
  assign new_n9714_ = ~pi0054 & ~new_n9704_;
  assign new_n9715_ = pi0038 & new_n9706_;
  assign new_n9716_ = new_n9714_ & ~new_n9715_;
  assign new_n9717_ = ~pi0074 & new_n9716_;
  assign new_n9718_ = new_n9712_ & ~new_n9717_;
  assign new_n9719_ = ~new_n3298_ & ~new_n9718_;
  assign new_n9720_ = new_n3436_ & ~new_n9719_;
  assign new_n9721_ = ~new_n3298_ & ~new_n9523_;
  assign new_n9722_ = new_n3436_ & ~new_n9721_;
  assign new_n9723_ = ~new_n9720_ & ~new_n9722_;
  assign new_n9724_ = pi0299 & ~new_n9702_;
  assign new_n9725_ = pi0140 & pi0145;
  assign new_n9726_ = ~pi0140 & ~pi0145;
  assign new_n9727_ = ~new_n9725_ & ~new_n9726_;
  assign new_n9728_ = new_n9001_ & ~new_n9727_;
  assign new_n9729_ = new_n9000_ & ~new_n9725_;
  assign new_n9730_ = new_n6185_ & ~new_n9726_;
  assign new_n9731_ = new_n9729_ & new_n9730_;
  assign new_n9732_ = ~pi0299 & ~new_n9731_;
  assign new_n9733_ = ~new_n9728_ & new_n9732_;
  assign new_n9734_ = pi0232 & ~new_n9733_;
  assign new_n9735_ = ~new_n9724_ & new_n9734_;
  assign new_n9736_ = pi0100 & ~new_n9735_;
  assign new_n9737_ = pi0075 & ~new_n9735_;
  assign new_n9738_ = ~new_n9736_ & ~new_n9737_;
  assign new_n9739_ = pi0141 & ~pi0299;
  assign new_n9740_ = pi0148 & pi0299;
  assign new_n9741_ = ~new_n9739_ & ~new_n9740_;
  assign new_n9742_ = new_n7499_ & ~new_n9741_;
  assign new_n9743_ = new_n8989_ & ~new_n9742_;
  assign new_n9744_ = new_n9738_ & ~new_n9743_;
  assign new_n9745_ = pi0074 & ~new_n9744_;
  assign new_n9746_ = ~pi0055 & ~new_n9745_;
  assign new_n9747_ = pi0188 & ~pi0299;
  assign new_n9748_ = pi0167 & pi0299;
  assign new_n9749_ = ~new_n9747_ & ~new_n9748_;
  assign new_n9750_ = new_n7499_ & ~new_n9749_;
  assign new_n9751_ = ~pi0100 & ~new_n9750_;
  assign new_n9752_ = ~pi0075 & new_n9751_;
  assign new_n9753_ = new_n9738_ & ~new_n9752_;
  assign new_n9754_ = pi0054 & ~new_n9753_;
  assign new_n9755_ = ~pi0142 & ~new_n9328_;
  assign new_n9756_ = pi0142 & new_n9177_;
  assign new_n9757_ = ~pi0140 & ~new_n9756_;
  assign new_n9758_ = ~new_n9755_ & new_n9757_;
  assign new_n9759_ = ~pi0142 & ~new_n9332_;
  assign new_n9760_ = pi0142 & ~new_n9233_;
  assign new_n9761_ = ~new_n9284_ & new_n9760_;
  assign new_n9762_ = pi0140 & ~new_n9761_;
  assign new_n9763_ = ~new_n9759_ & new_n9762_;
  assign new_n9764_ = ~new_n9758_ & ~new_n9763_;
  assign new_n9765_ = ~pi0181 & ~new_n9764_;
  assign new_n9766_ = ~pi0142 & ~new_n9310_;
  assign new_n9767_ = pi0142 & ~new_n9246_;
  assign new_n9768_ = ~pi0140 & ~new_n9767_;
  assign new_n9769_ = ~new_n9766_ & new_n9768_;
  assign new_n9770_ = ~pi0142 & ~new_n9319_;
  assign new_n9771_ = pi0142 & ~new_n9240_;
  assign new_n9772_ = pi0140 & ~new_n9771_;
  assign new_n9773_ = ~new_n9770_ & new_n9772_;
  assign new_n9774_ = ~new_n9769_ & ~new_n9773_;
  assign new_n9775_ = pi0181 & ~new_n9774_;
  assign new_n9776_ = pi0144 & ~new_n9775_;
  assign new_n9777_ = ~new_n9765_ & new_n9776_;
  assign new_n9778_ = ~pi0142 & ~new_n9281_;
  assign new_n9779_ = pi0142 & ~new_n9200_;
  assign new_n9780_ = ~pi0140 & ~new_n9779_;
  assign new_n9781_ = ~new_n9778_ & new_n9780_;
  assign new_n9782_ = pi0142 & ~new_n9216_;
  assign new_n9783_ = ~pi0142 & new_n9285_;
  assign new_n9784_ = pi0140 & ~new_n9783_;
  assign new_n9785_ = ~new_n9782_ & new_n9784_;
  assign new_n9786_ = ~new_n9781_ & ~new_n9785_;
  assign new_n9787_ = pi0181 & ~new_n9786_;
  assign new_n9788_ = ~pi0142 & new_n9351_;
  assign new_n9789_ = ~new_n9194_ & new_n9401_;
  assign new_n9790_ = new_n6185_ & ~new_n9789_;
  assign new_n9791_ = pi0142 & ~new_n9790_;
  assign new_n9792_ = ~new_n9284_ & new_n9791_;
  assign new_n9793_ = ~pi0140 & ~new_n9792_;
  assign new_n9794_ = ~new_n9788_ & new_n9793_;
  assign new_n9795_ = ~pi0142 & ~new_n9339_;
  assign new_n9796_ = pi0142 & ~new_n9422_;
  assign new_n9797_ = ~new_n9284_ & new_n9796_;
  assign new_n9798_ = pi0140 & ~new_n9797_;
  assign new_n9799_ = ~new_n9795_ & new_n9798_;
  assign new_n9800_ = ~new_n9794_ & ~new_n9799_;
  assign new_n9801_ = ~pi0181 & ~new_n9800_;
  assign new_n9802_ = ~pi0144 & ~new_n9801_;
  assign new_n9803_ = ~new_n9787_ & new_n9802_;
  assign new_n9804_ = ~pi0299 & ~new_n9803_;
  assign new_n9805_ = ~new_n9777_ & new_n9804_;
  assign new_n9806_ = ~pi0159 & pi0299;
  assign new_n9807_ = ~pi0146 & ~new_n9413_;
  assign new_n9808_ = pi0146 & new_n9423_;
  assign new_n9809_ = ~pi0161 & ~new_n9808_;
  assign new_n9810_ = ~new_n9807_ & new_n9809_;
  assign new_n9811_ = ~pi0146 & ~new_n9415_;
  assign new_n9812_ = pi0146 & new_n9419_;
  assign new_n9813_ = pi0161 & ~new_n9812_;
  assign new_n9814_ = ~new_n9811_ & new_n9813_;
  assign new_n9815_ = ~new_n9810_ & ~new_n9814_;
  assign new_n9816_ = pi0162 & ~new_n9815_;
  assign new_n9817_ = pi0161 & ~new_n9393_;
  assign new_n9818_ = ~pi0161 & ~new_n9396_;
  assign new_n9819_ = ~pi0146 & ~new_n9818_;
  assign new_n9820_ = ~new_n9817_ & new_n9819_;
  assign new_n9821_ = pi0161 & ~new_n9363_;
  assign new_n9822_ = ~pi0161 & ~new_n9403_;
  assign new_n9823_ = pi0146 & ~new_n9822_;
  assign new_n9824_ = ~new_n9821_ & new_n9823_;
  assign new_n9825_ = ~pi0162 & ~new_n9369_;
  assign new_n9826_ = ~new_n9824_ & new_n9825_;
  assign new_n9827_ = ~new_n9820_ & new_n9826_;
  assign new_n9828_ = ~new_n9816_ & ~new_n9827_;
  assign new_n9829_ = new_n9806_ & ~new_n9828_;
  assign new_n9830_ = ~pi0146 & ~new_n9437_;
  assign new_n9831_ = pi0146 & ~new_n9431_;
  assign new_n9832_ = pi0161 & ~new_n9831_;
  assign new_n9833_ = ~new_n9830_ & new_n9832_;
  assign new_n9834_ = pi0146 & ~new_n9429_;
  assign new_n9835_ = ~pi0146 & new_n9435_;
  assign new_n9836_ = ~pi0161 & ~new_n9835_;
  assign new_n9837_ = ~new_n9834_ & new_n9836_;
  assign new_n9838_ = pi0162 & ~new_n9837_;
  assign new_n9839_ = ~new_n9833_ & new_n9838_;
  assign new_n9840_ = pi0159 & pi0299;
  assign new_n9841_ = ~pi0146 & ~new_n9386_;
  assign new_n9842_ = pi0146 & ~new_n9372_;
  assign new_n9843_ = ~pi0161 & ~new_n9842_;
  assign new_n9844_ = ~new_n9841_ & new_n9843_;
  assign new_n9845_ = ~pi0146 & ~new_n9379_;
  assign new_n9846_ = pi0146 & new_n9367_;
  assign new_n9847_ = pi0161 & ~new_n9846_;
  assign new_n9848_ = ~new_n9845_ & new_n9847_;
  assign new_n9849_ = ~pi0162 & ~new_n9848_;
  assign new_n9850_ = ~new_n9844_ & new_n9849_;
  assign new_n9851_ = new_n9840_ & ~new_n9850_;
  assign new_n9852_ = ~new_n9839_ & new_n9851_;
  assign new_n9853_ = ~new_n9829_ & ~new_n9852_;
  assign new_n9854_ = ~new_n9805_ & new_n9853_;
  assign new_n9855_ = pi0232 & ~new_n9854_;
  assign new_n9856_ = ~new_n9450_ & ~new_n9855_;
  assign new_n9857_ = new_n3186_ & ~new_n9856_;
  assign new_n9858_ = pi0144 & new_n9104_;
  assign new_n9859_ = ~pi0177 & ~pi0299;
  assign new_n9860_ = ~pi0144 & ~new_n9060_;
  assign new_n9861_ = ~new_n9095_ & new_n9860_;
  assign new_n9862_ = new_n9859_ & ~new_n9861_;
  assign new_n9863_ = ~new_n9858_ & new_n9862_;
  assign new_n9864_ = ~new_n9060_ & ~new_n9065_;
  assign new_n9865_ = pi0177 & ~pi0299;
  assign new_n9866_ = ~new_n9860_ & new_n9865_;
  assign new_n9867_ = ~new_n9864_ & new_n9866_;
  assign new_n9868_ = ~new_n9863_ & ~new_n9867_;
  assign new_n9869_ = pi0232 & ~new_n9868_;
  assign new_n9870_ = ~new_n9107_ & ~new_n9869_;
  assign new_n9871_ = ~pi0038 & ~new_n9870_;
  assign new_n9872_ = ~pi0161 & new_n9075_;
  assign new_n9873_ = ~new_n9080_ & ~new_n9872_;
  assign new_n9874_ = new_n9069_ & ~new_n9873_;
  assign new_n9875_ = ~pi0038 & ~pi0155;
  assign new_n9876_ = new_n9071_ & new_n9875_;
  assign new_n9877_ = ~new_n9874_ & new_n9876_;
  assign new_n9878_ = pi0161 & new_n9084_;
  assign new_n9879_ = new_n9057_ & new_n9069_;
  assign new_n9880_ = ~new_n9878_ & new_n9879_;
  assign new_n9881_ = ~pi0038 & pi0155;
  assign new_n9882_ = new_n9071_ & new_n9881_;
  assign new_n9883_ = ~new_n9880_ & new_n9882_;
  assign new_n9884_ = ~new_n9877_ & ~new_n9883_;
  assign new_n9885_ = pi0232 & ~new_n9884_;
  assign new_n9886_ = ~new_n9871_ & ~new_n9885_;
  assign new_n9887_ = pi0039 & ~new_n9886_;
  assign new_n9888_ = pi0188 & new_n9032_;
  assign new_n9889_ = ~pi0167 & ~new_n9888_;
  assign new_n9890_ = ~pi0188 & ~new_n9025_;
  assign new_n9891_ = pi0167 & pi0188;
  assign new_n9892_ = ~new_n9027_ & new_n9891_;
  assign new_n9893_ = ~new_n9890_ & ~new_n9892_;
  assign new_n9894_ = ~new_n9889_ & new_n9893_;
  assign new_n9895_ = pi0038 & ~new_n9894_;
  assign new_n9896_ = ~pi0087 & ~new_n9895_;
  assign new_n9897_ = ~new_n9887_ & new_n9896_;
  assign new_n9898_ = ~new_n9857_ & new_n9897_;
  assign new_n9899_ = pi0038 & ~new_n9750_;
  assign new_n9900_ = ~new_n9495_ & ~new_n9899_;
  assign new_n9901_ = pi0087 & new_n9900_;
  assign new_n9902_ = ~pi0100 & ~new_n9901_;
  assign new_n9903_ = ~new_n9898_ & new_n9902_;
  assign new_n9904_ = ~new_n9736_ & ~new_n9903_;
  assign new_n9905_ = new_n3242_ & ~new_n9904_;
  assign new_n9906_ = pi0155 & pi0299;
  assign new_n9907_ = ~new_n9865_ & ~new_n9906_;
  assign new_n9908_ = ~pi0038 & new_n9907_;
  assign new_n9909_ = new_n7499_ & ~new_n9908_;
  assign new_n9910_ = new_n9472_ & ~new_n9909_;
  assign new_n9911_ = new_n9900_ & ~new_n9910_;
  assign new_n9912_ = ~pi0100 & ~new_n9911_;
  assign new_n9913_ = ~new_n9736_ & ~new_n9912_;
  assign new_n9914_ = new_n9467_ & ~new_n9913_;
  assign new_n9915_ = ~new_n9737_ & ~new_n9914_;
  assign new_n9916_ = ~new_n9905_ & new_n9915_;
  assign new_n9917_ = ~pi0054 & ~new_n9916_;
  assign new_n9918_ = ~new_n9754_ & ~new_n9917_;
  assign new_n9919_ = ~pi0074 & ~new_n9918_;
  assign new_n9920_ = new_n9746_ & ~new_n9919_;
  assign new_n9921_ = pi0055 & ~new_n9711_;
  assign new_n9922_ = pi0054 & new_n9707_;
  assign new_n9923_ = ~new_n9522_ & new_n9716_;
  assign new_n9924_ = ~new_n6290_ & ~new_n9923_;
  assign new_n9925_ = pi0100 & ~new_n9703_;
  assign new_n9926_ = pi0038 & new_n9705_;
  assign new_n9927_ = new_n9472_ & ~new_n9694_;
  assign new_n9928_ = new_n9521_ & ~new_n9927_;
  assign new_n9929_ = ~pi0100 & ~new_n9928_;
  assign new_n9930_ = ~pi0232 & new_n9472_;
  assign new_n9931_ = ~new_n9929_ & ~new_n9930_;
  assign new_n9932_ = ~new_n9926_ & ~new_n9931_;
  assign new_n9933_ = ~new_n9925_ & ~new_n9932_;
  assign new_n9934_ = ~pi0075 & ~new_n9933_;
  assign new_n9935_ = pi0075 & ~new_n9703_;
  assign new_n9936_ = ~pi0092 & ~new_n9935_;
  assign new_n9937_ = ~new_n9934_ & new_n9936_;
  assign new_n9938_ = ~new_n9924_ & ~new_n9937_;
  assign new_n9939_ = ~new_n9922_ & ~new_n9938_;
  assign new_n9940_ = ~pi0074 & ~new_n9939_;
  assign new_n9941_ = new_n9921_ & ~new_n9940_;
  assign new_n9942_ = new_n3298_ & ~new_n9941_;
  assign new_n9943_ = ~new_n9920_ & new_n9942_;
  assign new_n9944_ = ~new_n9723_ & ~new_n9943_;
  assign new_n9945_ = ~new_n9713_ & ~new_n9944_;
  assign new_n9946_ = ~pi0034 & new_n9945_;
  assign new_n9947_ = ~pi0142 & new_n9582_;
  assign new_n9948_ = pi0142 & new_n9609_;
  assign new_n9949_ = ~pi0140 & ~new_n9948_;
  assign new_n9950_ = ~new_n9947_ & new_n9949_;
  assign new_n9951_ = ~pi0142 & new_n9570_;
  assign new_n9952_ = pi0140 & new_n9600_;
  assign new_n9953_ = ~new_n9951_ & new_n9952_;
  assign new_n9954_ = ~new_n9950_ & ~new_n9953_;
  assign new_n9955_ = ~pi0144 & ~new_n9954_;
  assign new_n9956_ = pi0140 & ~new_n6185_;
  assign new_n9957_ = ~pi0142 & new_n9594_;
  assign new_n9958_ = ~pi0140 & ~new_n9957_;
  assign new_n9959_ = ~pi0142 & new_n9589_;
  assign new_n9960_ = pi0140 & ~new_n9959_;
  assign new_n9961_ = new_n9603_ & new_n9960_;
  assign new_n9962_ = ~new_n9958_ & ~new_n9961_;
  assign new_n9963_ = pi0144 & ~new_n9962_;
  assign new_n9964_ = ~new_n9956_ & ~new_n9963_;
  assign new_n9965_ = ~new_n9955_ & new_n9964_;
  assign new_n9966_ = pi0181 & new_n9615_;
  assign new_n9967_ = ~pi0299 & ~new_n9966_;
  assign new_n9968_ = ~new_n9965_ & new_n9967_;
  assign new_n9969_ = ~pi0146 & ~new_n9582_;
  assign new_n9970_ = pi0146 & ~new_n9609_;
  assign new_n9971_ = ~pi0161 & ~new_n9970_;
  assign new_n9972_ = ~new_n9969_ & new_n9971_;
  assign new_n9973_ = ~pi0146 & pi0161;
  assign new_n9974_ = new_n9594_ & new_n9973_;
  assign new_n9975_ = ~new_n9972_ & ~new_n9974_;
  assign new_n9976_ = ~pi0162 & ~new_n9975_;
  assign new_n9977_ = ~pi0162 & new_n9615_;
  assign new_n9978_ = new_n9840_ & ~new_n9977_;
  assign new_n9979_ = ~new_n9806_ & ~new_n9978_;
  assign new_n9980_ = ~new_n9694_ & ~new_n9979_;
  assign new_n9981_ = ~pi0146 & new_n9570_;
  assign new_n9982_ = new_n9621_ & ~new_n9981_;
  assign new_n9983_ = ~pi0161 & ~new_n9982_;
  assign new_n9984_ = ~pi0146 & new_n9589_;
  assign new_n9985_ = new_n9624_ & ~new_n9984_;
  assign new_n9986_ = pi0161 & ~new_n9985_;
  assign new_n9987_ = pi0159 & new_n2943_;
  assign new_n9988_ = pi0299 & ~new_n9987_;
  assign new_n9989_ = ~new_n9986_ & new_n9988_;
  assign new_n9990_ = ~new_n9983_ & new_n9989_;
  assign new_n9991_ = ~new_n9980_ & ~new_n9990_;
  assign new_n9992_ = ~new_n9976_ & ~new_n9991_;
  assign new_n9993_ = pi0232 & ~new_n9992_;
  assign new_n9994_ = ~new_n9968_ & new_n9993_;
  assign new_n9995_ = new_n3186_ & ~new_n9994_;
  assign new_n9996_ = pi0161 & ~new_n9551_;
  assign new_n9997_ = ~pi0161 & ~new_n9544_;
  assign new_n9998_ = new_n9069_ & ~new_n9997_;
  assign new_n9999_ = ~new_n9996_ & new_n9998_;
  assign new_n10000_ = new_n9881_ & ~new_n9999_;
  assign new_n10001_ = ~pi0161 & new_n9069_;
  assign new_n10002_ = new_n9546_ & new_n10001_;
  assign new_n10003_ = new_n9875_ & ~new_n10002_;
  assign new_n10004_ = ~new_n10000_ & ~new_n10003_;
  assign new_n10005_ = pi0299 & ~new_n10004_;
  assign new_n10006_ = ~pi0144 & new_n9535_;
  assign new_n10007_ = pi0144 & new_n9538_;
  assign new_n10008_ = new_n9865_ & ~new_n10007_;
  assign new_n10009_ = ~new_n10006_ & new_n10008_;
  assign new_n10010_ = ~pi0144 & new_n9530_;
  assign new_n10011_ = new_n9859_ & ~new_n10010_;
  assign new_n10012_ = pi0232 & ~new_n10011_;
  assign new_n10013_ = ~new_n10009_ & new_n10012_;
  assign new_n10014_ = ~pi0038 & ~new_n10013_;
  assign new_n10015_ = ~new_n10005_ & ~new_n10014_;
  assign new_n10016_ = pi0039 & ~new_n10015_;
  assign new_n10017_ = ~new_n9895_ & ~new_n10016_;
  assign new_n10018_ = ~new_n9995_ & new_n10017_;
  assign new_n10019_ = ~pi0100 & ~new_n10018_;
  assign new_n10020_ = ~new_n9736_ & ~new_n10019_;
  assign new_n10021_ = ~pi0087 & ~new_n10020_;
  assign new_n10022_ = ~new_n3211_ & ~new_n9751_;
  assign new_n10023_ = ~new_n9736_ & new_n10022_;
  assign new_n10024_ = pi0087 & ~new_n10023_;
  assign new_n10025_ = ~new_n10021_ & ~new_n10024_;
  assign new_n10026_ = new_n3242_ & ~new_n10025_;
  assign new_n10027_ = pi0038 & ~new_n9749_;
  assign new_n10028_ = new_n3186_ & ~new_n9907_;
  assign new_n10029_ = new_n3094_ & new_n10028_;
  assign new_n10030_ = ~new_n10027_ & ~new_n10029_;
  assign new_n10031_ = new_n7499_ & ~new_n10030_;
  assign new_n10032_ = ~pi0100 & ~new_n10031_;
  assign new_n10033_ = ~new_n9736_ & ~new_n10032_;
  assign new_n10034_ = ~pi0087 & ~new_n10033_;
  assign new_n10035_ = ~new_n10024_ & ~new_n10034_;
  assign new_n10036_ = new_n9467_ & ~new_n10035_;
  assign new_n10037_ = ~new_n9737_ & ~new_n10036_;
  assign new_n10038_ = ~new_n10026_ & new_n10037_;
  assign new_n10039_ = ~pi0054 & ~new_n10038_;
  assign new_n10040_ = ~new_n9754_ & ~new_n10039_;
  assign new_n10041_ = ~pi0074 & ~new_n10040_;
  assign new_n10042_ = new_n9746_ & ~new_n10041_;
  assign new_n10043_ = ~pi0092 & pi0162;
  assign new_n10044_ = new_n9619_ & new_n10043_;
  assign new_n10045_ = new_n9653_ & new_n10044_;
  assign new_n10046_ = new_n6203_ & new_n10045_;
  assign new_n10047_ = ~new_n9926_ & ~new_n10046_;
  assign new_n10048_ = new_n8989_ & ~new_n10047_;
  assign new_n10049_ = new_n9714_ & ~new_n10048_;
  assign new_n10050_ = ~new_n9922_ & ~new_n10049_;
  assign new_n10051_ = ~pi0074 & ~new_n10050_;
  assign new_n10052_ = new_n9921_ & ~new_n10051_;
  assign new_n10053_ = new_n3298_ & ~new_n10052_;
  assign new_n10054_ = ~new_n10042_ & new_n10053_;
  assign new_n10055_ = new_n9720_ & ~new_n10054_;
  assign new_n10056_ = ~new_n9713_ & ~new_n10055_;
  assign new_n10057_ = pi0034 & new_n10056_;
  assign new_n10058_ = ~pi0033 & ~pi0954;
  assign new_n10059_ = ~new_n10057_ & ~new_n10058_;
  assign new_n10060_ = ~new_n9946_ & new_n10059_;
  assign new_n10061_ = ~pi0034 & ~new_n8978_;
  assign new_n10062_ = new_n9945_ & ~new_n10061_;
  assign new_n10063_ = new_n10056_ & new_n10061_;
  assign new_n10064_ = new_n10058_ & ~new_n10063_;
  assign new_n10065_ = ~new_n10062_ & new_n10064_;
  assign po0192 = ~new_n10060_ & ~new_n10065_;
  assign new_n10067_ = pi0137 & new_n8884_;
  assign new_n10068_ = new_n2732_ & new_n2797_;
  assign new_n10069_ = new_n7511_ & ~new_n10068_;
  assign new_n10070_ = pi0683 & new_n10069_;
  assign new_n10071_ = pi0252 & po1057;
  assign new_n10072_ = ~new_n10070_ & new_n10071_;
  assign new_n10073_ = pi0146 & new_n7497_;
  assign new_n10074_ = pi0142 & new_n7496_;
  assign new_n10075_ = ~new_n10073_ & ~new_n10074_;
  assign new_n10076_ = ~new_n7498_ & new_n10075_;
  assign new_n10077_ = ~new_n10072_ & ~new_n10076_;
  assign new_n10078_ = ~new_n7500_ & ~new_n10077_;
  assign new_n10079_ = ~new_n8887_ & ~new_n10078_;
  assign new_n10080_ = new_n6263_ & ~new_n8889_;
  assign new_n10081_ = ~new_n10072_ & new_n10080_;
  assign new_n10082_ = ~new_n10079_ & ~new_n10081_;
  assign new_n10083_ = new_n8886_ & ~new_n10082_;
  assign new_n10084_ = ~new_n10067_ & ~new_n10083_;
  assign new_n10085_ = new_n8882_ & ~new_n10084_;
  assign new_n10086_ = ~pi0090 & new_n6135_;
  assign new_n10087_ = ~pi0093 & ~new_n10086_;
  assign new_n10088_ = ~new_n6154_ & ~new_n10087_;
  assign new_n10089_ = ~pi0035 & ~new_n10088_;
  assign new_n10090_ = pi0035 & ~new_n2735_;
  assign new_n10091_ = new_n8938_ & ~new_n10090_;
  assign new_n10092_ = ~new_n10089_ & new_n10091_;
  assign new_n10093_ = ~pi0032 & new_n10092_;
  assign new_n10094_ = pi0032 & ~pi0093;
  assign new_n10095_ = new_n8895_ & new_n10094_;
  assign new_n10096_ = new_n7458_ & new_n10095_;
  assign new_n10097_ = ~new_n10093_ & ~new_n10096_;
  assign new_n10098_ = ~pi0095 & ~new_n6166_;
  assign new_n10099_ = ~new_n10097_ & new_n10098_;
  assign new_n10100_ = ~new_n2553_ & ~new_n10092_;
  assign new_n10101_ = pi1082 & new_n3097_;
  assign new_n10102_ = ~new_n10100_ & new_n10101_;
  assign new_n10103_ = new_n6166_ & ~new_n10089_;
  assign new_n10104_ = new_n2733_ & new_n7561_;
  assign new_n10105_ = ~pi0137 & ~new_n6166_;
  assign new_n10106_ = ~new_n7733_ & ~new_n10105_;
  assign new_n10107_ = new_n10104_ & new_n10106_;
  assign new_n10108_ = ~pi0122 & ~po0740;
  assign new_n10109_ = new_n7733_ & ~new_n10105_;
  assign new_n10110_ = new_n10108_ & new_n10109_;
  assign new_n10111_ = ~new_n10107_ & ~new_n10110_;
  assign new_n10112_ = ~new_n10103_ & new_n10111_;
  assign new_n10113_ = new_n2493_ & new_n8936_;
  assign new_n10114_ = new_n10089_ & ~new_n10113_;
  assign new_n10115_ = new_n3097_ & new_n10091_;
  assign new_n10116_ = ~new_n10114_ & new_n10115_;
  assign new_n10117_ = ~new_n10112_ & new_n10116_;
  assign new_n10118_ = ~pi0038 & ~new_n10117_;
  assign new_n10119_ = ~new_n10102_ & new_n10118_;
  assign new_n10120_ = ~new_n10099_ & new_n10119_;
  assign new_n10121_ = pi0038 & ~new_n8962_;
  assign new_n10122_ = ~pi0039 & ~pi0100;
  assign new_n10123_ = ~new_n10121_ & new_n10122_;
  assign new_n10124_ = ~new_n10120_ & new_n10123_;
  assign new_n10125_ = ~new_n10085_ & ~new_n10124_;
  assign new_n10126_ = new_n3235_ & ~new_n10125_;
  assign new_n10127_ = pi0137 & ~po0840;
  assign new_n10128_ = ~new_n6282_ & new_n10127_;
  assign new_n10129_ = ~new_n8964_ & ~new_n10128_;
  assign new_n10130_ = new_n8967_ & ~new_n10129_;
  assign new_n10131_ = new_n8962_ & new_n10130_;
  assign new_n10132_ = ~new_n10126_ & ~new_n10131_;
  assign new_n10133_ = ~pi0092 & ~new_n10132_;
  assign new_n10134_ = ~pi0054 & ~new_n10133_;
  assign new_n10135_ = ~pi0024 & new_n7340_;
  assign new_n10136_ = pi0054 & ~new_n10135_;
  assign new_n10137_ = new_n3298_ & new_n8879_;
  assign new_n10138_ = ~new_n10136_ & new_n10137_;
  assign new_n10139_ = ~new_n10134_ & new_n10138_;
  assign new_n10140_ = ~pi0059 & ~new_n10139_;
  assign new_n10141_ = new_n3273_ & new_n3298_;
  assign new_n10142_ = new_n8962_ & new_n10141_;
  assign new_n10143_ = ~pi0055 & new_n10142_;
  assign new_n10144_ = pi0059 & ~new_n10143_;
  assign new_n10145_ = ~pi0057 & ~new_n10144_;
  assign po0193 = ~new_n10140_ & new_n10145_;
  assign new_n10147_ = new_n2514_ & new_n2580_;
  assign new_n10148_ = ~pi0083 & new_n2647_;
  assign new_n10149_ = ~pi0065 & new_n2451_;
  assign new_n10150_ = new_n2476_ & new_n10149_;
  assign new_n10151_ = new_n9039_ & new_n10150_;
  assign new_n10152_ = ~pi0069 & new_n10151_;
  assign new_n10153_ = ~pi0067 & ~pi0071;
  assign new_n10154_ = pi0036 & ~pi0103;
  assign new_n10155_ = new_n10153_ & new_n10154_;
  assign new_n10156_ = new_n10152_ & new_n10155_;
  assign new_n10157_ = new_n10148_ & new_n10156_;
  assign new_n10158_ = new_n10147_ & new_n10157_;
  assign new_n10159_ = ~pi0058 & new_n7516_;
  assign new_n10160_ = ~new_n10158_ & ~new_n10159_;
  assign new_n10161_ = new_n2493_ & new_n6379_;
  assign new_n10162_ = new_n6167_ & new_n10161_;
  assign new_n10163_ = new_n3270_ & ~po1038;
  assign new_n10164_ = new_n3413_ & new_n10163_;
  assign new_n10165_ = ~pi0092 & new_n10164_;
  assign new_n10166_ = new_n10162_ & new_n10165_;
  assign new_n10167_ = po0740 & new_n10166_;
  assign po0194 = ~new_n10160_ & new_n10167_;
  assign new_n10169_ = ~pi0039 & new_n3098_;
  assign new_n10170_ = pi0024 & new_n10169_;
  assign new_n10171_ = new_n2498_ & new_n10170_;
  assign new_n10172_ = pi0038 & ~new_n10171_;
  assign new_n10173_ = ~pi0081 & ~new_n2598_;
  assign new_n10174_ = new_n6379_ & new_n9258_;
  assign new_n10175_ = new_n2520_ & new_n10174_;
  assign new_n10176_ = new_n2551_ & new_n10175_;
  assign new_n10177_ = ~pi0071 & new_n2476_;
  assign new_n10178_ = ~pi0104 & new_n2461_;
  assign new_n10179_ = new_n10177_ & new_n10178_;
  assign new_n10180_ = ~pi0045 & ~pi0073;
  assign new_n10181_ = new_n8912_ & new_n10180_;
  assign new_n10182_ = ~pi0048 & ~pi0065;
  assign new_n10183_ = ~pi0082 & ~pi0084;
  assign new_n10184_ = pi0089 & new_n10183_;
  assign new_n10185_ = new_n10182_ & new_n10184_;
  assign new_n10186_ = new_n10181_ & new_n10185_;
  assign new_n10187_ = new_n9130_ & new_n10186_;
  assign new_n10188_ = new_n10179_ & new_n10187_;
  assign new_n10189_ = pi0332 & new_n10188_;
  assign new_n10190_ = ~pi0064 & ~new_n10189_;
  assign new_n10191_ = ~pi0039 & ~pi0841;
  assign new_n10192_ = new_n2454_ & new_n10191_;
  assign new_n10193_ = ~new_n10190_ & new_n10192_;
  assign new_n10194_ = new_n10176_ & new_n10193_;
  assign new_n10195_ = new_n10173_ & new_n10194_;
  assign new_n10196_ = ~pi0038 & ~new_n10195_;
  assign new_n10197_ = new_n3272_ & ~po1038;
  assign new_n10198_ = ~new_n10196_ & new_n10197_;
  assign po0196 = ~new_n10172_ & new_n10198_;
  assign new_n10200_ = ~pi0038 & new_n10197_;
  assign new_n10201_ = ~pi0984 & ~new_n2799_;
  assign new_n10202_ = pi0835 & ~new_n10201_;
  assign new_n10203_ = new_n6188_ & ~new_n10202_;
  assign new_n10204_ = new_n6198_ & ~new_n10203_;
  assign new_n10205_ = pi1093 & new_n10204_;
  assign new_n10206_ = new_n6189_ & new_n6454_;
  assign new_n10207_ = ~new_n10205_ & new_n10206_;
  assign new_n10208_ = ~pi0215 & new_n10207_;
  assign new_n10209_ = ~new_n6215_ & new_n10204_;
  assign new_n10210_ = new_n10206_ & ~new_n10209_;
  assign new_n10211_ = ~new_n6212_ & new_n10210_;
  assign new_n10212_ = new_n6221_ & new_n10204_;
  assign new_n10213_ = new_n10206_ & ~new_n10212_;
  assign new_n10214_ = new_n6212_ & new_n10213_;
  assign new_n10215_ = pi0299 & ~new_n10214_;
  assign new_n10216_ = ~new_n10211_ & new_n10215_;
  assign new_n10217_ = ~new_n10208_ & new_n10216_;
  assign new_n10218_ = pi0786 & ~pi1082;
  assign new_n10219_ = ~pi0223 & new_n10207_;
  assign new_n10220_ = ~new_n6238_ & new_n10210_;
  assign new_n10221_ = new_n6238_ & new_n10213_;
  assign new_n10222_ = ~pi0299 & ~new_n10221_;
  assign new_n10223_ = ~new_n10220_ & new_n10222_;
  assign new_n10224_ = ~new_n10219_ & new_n10223_;
  assign new_n10225_ = ~new_n10218_ & ~new_n10224_;
  assign new_n10226_ = ~new_n10217_ & new_n10225_;
  assign new_n10227_ = new_n5788_ & ~new_n6223_;
  assign new_n10228_ = new_n3489_ & ~new_n6244_;
  assign new_n10229_ = ~new_n10227_ & ~new_n10228_;
  assign new_n10230_ = po0740 & new_n10218_;
  assign new_n10231_ = ~new_n10229_ & new_n10230_;
  assign new_n10232_ = new_n6456_ & new_n10231_;
  assign new_n10233_ = ~new_n10226_ & ~new_n10232_;
  assign new_n10234_ = pi0039 & ~new_n10233_;
  assign new_n10235_ = ~pi0039 & ~pi0095;
  assign new_n10236_ = new_n6166_ & new_n6386_;
  assign new_n10237_ = new_n2510_ & ~new_n2583_;
  assign new_n10238_ = new_n8916_ & new_n8921_;
  assign new_n10239_ = new_n9127_ & new_n10238_;
  assign new_n10240_ = new_n8917_ & new_n9131_;
  assign new_n10241_ = ~pi0065 & ~pi0069;
  assign new_n10242_ = new_n10240_ & new_n10241_;
  assign new_n10243_ = pi0048 & ~pi0049;
  assign new_n10244_ = ~pi0068 & ~pi0082;
  assign new_n10245_ = new_n10243_ & new_n10244_;
  assign new_n10246_ = new_n10180_ & new_n10245_;
  assign new_n10247_ = new_n10242_ & new_n10246_;
  assign new_n10248_ = new_n10239_ & new_n10247_;
  assign new_n10249_ = new_n10179_ & new_n10248_;
  assign new_n10250_ = ~pi0841 & new_n2483_;
  assign new_n10251_ = new_n2505_ & new_n10250_;
  assign new_n10252_ = ~pi0097 & new_n10251_;
  assign new_n10253_ = new_n10249_ & new_n10252_;
  assign new_n10254_ = new_n10237_ & new_n10253_;
  assign new_n10255_ = pi0108 & new_n2510_;
  assign new_n10256_ = new_n2582_ & new_n10255_;
  assign new_n10257_ = ~pi0047 & ~new_n10256_;
  assign new_n10258_ = ~new_n10254_ & new_n10257_;
  assign new_n10259_ = ~pi0986 & ~po0740;
  assign new_n10260_ = pi0252 & ~new_n10259_;
  assign new_n10261_ = pi0314 & ~new_n10260_;
  assign new_n10262_ = new_n6148_ & new_n10261_;
  assign new_n10263_ = ~new_n10258_ & new_n10262_;
  assign new_n10264_ = ~pi0047 & ~pi0841;
  assign new_n10265_ = new_n10249_ & new_n10264_;
  assign new_n10266_ = ~new_n2569_ & ~new_n10265_;
  assign new_n10267_ = new_n2489_ & new_n2519_;
  assign new_n10268_ = ~new_n10261_ & new_n10267_;
  assign new_n10269_ = ~new_n10266_ & new_n10268_;
  assign new_n10270_ = ~new_n10263_ & ~new_n10269_;
  assign new_n10271_ = new_n2493_ & ~new_n10270_;
  assign new_n10272_ = ~pi0035 & ~new_n10271_;
  assign new_n10273_ = pi0035 & ~new_n6383_;
  assign new_n10274_ = new_n2551_ & ~new_n10273_;
  assign new_n10275_ = new_n2724_ & new_n10274_;
  assign new_n10276_ = ~new_n10272_ & new_n10275_;
  assign new_n10277_ = ~new_n10236_ & ~new_n10276_;
  assign new_n10278_ = new_n10235_ & ~new_n10277_;
  assign new_n10279_ = ~new_n10234_ & ~new_n10278_;
  assign po0197 = new_n10200_ & ~new_n10279_;
  assign new_n10281_ = new_n3097_ & ~new_n3366_;
  assign new_n10282_ = ~pi0093 & pi0102;
  assign new_n10283_ = new_n2518_ & new_n10282_;
  assign new_n10284_ = new_n2453_ & new_n10283_;
  assign new_n10285_ = new_n6167_ & new_n10284_;
  assign new_n10286_ = new_n2520_ & new_n10285_;
  assign new_n10287_ = new_n2479_ & new_n10286_;
  assign new_n10288_ = ~pi0040 & ~new_n10287_;
  assign new_n10289_ = new_n10281_ & ~new_n10288_;
  assign new_n10290_ = ~pi1082 & ~new_n10289_;
  assign new_n10291_ = new_n6379_ & new_n10287_;
  assign new_n10292_ = pi1082 & ~new_n10291_;
  assign new_n10293_ = new_n10165_ & ~new_n10292_;
  assign po0198 = ~new_n10290_ & new_n10293_;
  assign new_n10295_ = ~pi0041 & ~pi0072;
  assign new_n10296_ = ~new_n8100_ & ~new_n10295_;
  assign new_n10297_ = ~new_n2733_ & new_n10295_;
  assign new_n10298_ = new_n8100_ & ~new_n10297_;
  assign new_n10299_ = ~pi0044 & new_n3100_;
  assign new_n10300_ = ~pi0101 & new_n10299_;
  assign new_n10301_ = new_n7561_ & new_n10300_;
  assign new_n10302_ = new_n7502_ & new_n10301_;
  assign new_n10303_ = pi0041 & ~new_n10302_;
  assign new_n10304_ = ~pi0041 & pi0072;
  assign new_n10305_ = new_n2733_ & ~new_n10304_;
  assign new_n10306_ = ~pi0099 & new_n6272_;
  assign new_n10307_ = ~pi0072 & pi0101;
  assign new_n10308_ = ~pi0041 & ~new_n10307_;
  assign new_n10309_ = ~pi0024 & new_n2498_;
  assign new_n10310_ = pi0252 & new_n6379_;
  assign new_n10311_ = new_n7561_ & new_n10310_;
  assign new_n10312_ = new_n10309_ & new_n10311_;
  assign new_n10313_ = ~pi0044 & new_n10312_;
  assign new_n10314_ = new_n10308_ & new_n10313_;
  assign new_n10315_ = ~new_n10306_ & new_n10314_;
  assign new_n10316_ = new_n10305_ & ~new_n10315_;
  assign new_n10317_ = ~new_n10303_ & new_n10316_;
  assign new_n10318_ = new_n10298_ & ~new_n10317_;
  assign new_n10319_ = ~new_n10296_ & ~new_n10318_;
  assign new_n10320_ = ~pi0039 & ~new_n10319_;
  assign new_n10321_ = ~pi0166 & new_n6185_;
  assign new_n10322_ = pi0161 & new_n10321_;
  assign new_n10323_ = ~pi0152 & new_n10322_;
  assign new_n10324_ = ~new_n7496_ & ~new_n10323_;
  assign new_n10325_ = ~pi0189 & new_n6185_;
  assign new_n10326_ = pi0144 & new_n10325_;
  assign new_n10327_ = ~pi0174 & new_n10326_;
  assign new_n10328_ = ~pi0299 & ~new_n10327_;
  assign new_n10329_ = pi0232 & ~new_n10328_;
  assign new_n10330_ = ~new_n10324_ & new_n10329_;
  assign new_n10331_ = ~pi0072 & ~new_n10330_;
  assign new_n10332_ = pi0039 & ~new_n10331_;
  assign new_n10333_ = new_n3246_ & ~new_n10332_;
  assign new_n10334_ = ~new_n10320_ & new_n10333_;
  assign new_n10335_ = ~pi0039 & ~new_n10295_;
  assign new_n10336_ = ~new_n10332_ & ~new_n10335_;
  assign new_n10337_ = ~new_n3246_ & new_n10336_;
  assign new_n10338_ = pi0075 & ~new_n10337_;
  assign new_n10339_ = ~new_n10334_ & new_n10338_;
  assign new_n10340_ = new_n7477_ & ~new_n7483_;
  assign new_n10341_ = ~pi1093 & ~new_n7485_;
  assign new_n10342_ = ~new_n10340_ & new_n10341_;
  assign new_n10343_ = ~pi0044 & ~new_n10342_;
  assign new_n10344_ = new_n2761_ & ~new_n7469_;
  assign new_n10345_ = new_n2759_ & new_n10344_;
  assign new_n10346_ = ~new_n7516_ & ~new_n10345_;
  assign new_n10347_ = new_n2518_ & ~new_n10346_;
  assign new_n10348_ = new_n7460_ & ~new_n10347_;
  assign new_n10349_ = new_n7457_ & ~new_n10348_;
  assign new_n10350_ = ~pi0051 & ~new_n10349_;
  assign new_n10351_ = ~new_n2558_ & ~new_n10350_;
  assign new_n10352_ = ~pi0096 & ~new_n10351_;
  assign new_n10353_ = new_n6379_ & ~new_n7481_;
  assign new_n10354_ = ~pi0072 & new_n7483_;
  assign new_n10355_ = new_n10353_ & new_n10354_;
  assign new_n10356_ = ~new_n10352_ & new_n10355_;
  assign new_n10357_ = ~new_n10340_ & ~new_n10356_;
  assign new_n10358_ = pi1093 & new_n10357_;
  assign new_n10359_ = new_n10343_ & ~new_n10358_;
  assign new_n10360_ = ~pi0101 & new_n10359_;
  assign new_n10361_ = pi0041 & ~new_n10360_;
  assign new_n10362_ = pi0044 & pi0072;
  assign new_n10363_ = ~new_n7480_ & new_n10353_;
  assign new_n10364_ = new_n10354_ & ~new_n10363_;
  assign new_n10365_ = ~pi0072 & ~new_n7477_;
  assign new_n10366_ = ~new_n7483_ & new_n10365_;
  assign new_n10367_ = ~pi1093 & ~new_n10366_;
  assign new_n10368_ = ~new_n10364_ & new_n10367_;
  assign new_n10369_ = ~pi0072 & new_n10357_;
  assign new_n10370_ = pi1093 & ~new_n10369_;
  assign new_n10371_ = ~new_n10368_ & ~new_n10370_;
  assign new_n10372_ = ~pi0044 & ~new_n10371_;
  assign new_n10373_ = ~new_n10362_ & ~new_n10372_;
  assign new_n10374_ = ~pi0101 & new_n10373_;
  assign new_n10375_ = new_n10308_ & ~new_n10374_;
  assign new_n10376_ = new_n2733_ & ~new_n10375_;
  assign new_n10377_ = ~new_n10361_ & new_n10376_;
  assign new_n10378_ = new_n10365_ & ~new_n10368_;
  assign new_n10379_ = ~pi0044 & ~new_n10378_;
  assign new_n10380_ = ~new_n10362_ & ~new_n10379_;
  assign new_n10381_ = ~pi0101 & new_n10380_;
  assign new_n10382_ = new_n10308_ & ~new_n10381_;
  assign new_n10383_ = pi1093 & ~new_n7477_;
  assign new_n10384_ = new_n10343_ & ~new_n10383_;
  assign new_n10385_ = ~pi0101 & new_n10384_;
  assign new_n10386_ = pi0041 & ~new_n10385_;
  assign new_n10387_ = ~new_n2733_ & ~new_n10386_;
  assign new_n10388_ = ~new_n10382_ & new_n10387_;
  assign new_n10389_ = pi0228 & ~new_n10388_;
  assign new_n10390_ = ~new_n10377_ & new_n10389_;
  assign new_n10391_ = ~pi0109 & new_n6349_;
  assign new_n10392_ = new_n2589_ & new_n10391_;
  assign new_n10393_ = ~pi0110 & ~new_n10392_;
  assign new_n10394_ = new_n2489_ & ~new_n2568_;
  assign new_n10395_ = ~pi0480 & pi0949;
  assign new_n10396_ = new_n2497_ & new_n10395_;
  assign new_n10397_ = ~pi0047 & new_n10396_;
  assign new_n10398_ = new_n10394_ & new_n10397_;
  assign new_n10399_ = ~new_n10393_ & new_n10398_;
  assign new_n10400_ = pi0901 & ~pi0959;
  assign new_n10401_ = new_n2514_ & new_n2589_;
  assign new_n10402_ = new_n2497_ & new_n10401_;
  assign new_n10403_ = ~new_n10395_ & new_n10402_;
  assign new_n10404_ = new_n10400_ & ~new_n10403_;
  assign new_n10405_ = ~new_n10399_ & new_n10404_;
  assign new_n10406_ = new_n2490_ & new_n2567_;
  assign new_n10407_ = pi0110 & new_n10406_;
  assign new_n10408_ = new_n10396_ & new_n10407_;
  assign new_n10409_ = ~new_n10400_ & ~new_n10408_;
  assign new_n10410_ = ~pi0250 & pi0252;
  assign new_n10411_ = new_n6379_ & new_n10410_;
  assign new_n10412_ = ~new_n10409_ & new_n10411_;
  assign new_n10413_ = ~new_n10405_ & new_n10412_;
  assign new_n10414_ = ~pi0072 & new_n10413_;
  assign new_n10415_ = new_n10162_ & new_n10407_;
  assign new_n10416_ = new_n10395_ & ~new_n10410_;
  assign new_n10417_ = new_n10415_ & new_n10416_;
  assign new_n10418_ = ~new_n10414_ & ~new_n10417_;
  assign new_n10419_ = ~pi0044 & ~new_n10418_;
  assign new_n10420_ = ~pi0101 & new_n10419_;
  assign new_n10421_ = pi0041 & ~new_n10420_;
  assign new_n10422_ = new_n6379_ & ~new_n10410_;
  assign new_n10423_ = new_n10408_ & new_n10422_;
  assign new_n10424_ = ~pi0072 & ~new_n10423_;
  assign new_n10425_ = ~new_n10413_ & new_n10424_;
  assign new_n10426_ = ~pi0044 & ~new_n10425_;
  assign new_n10427_ = ~new_n10362_ & ~new_n10426_;
  assign new_n10428_ = ~pi0101 & new_n10427_;
  assign new_n10429_ = new_n10308_ & ~new_n10428_;
  assign new_n10430_ = ~new_n10421_ & ~new_n10429_;
  assign new_n10431_ = ~pi0228 & ~new_n10430_;
  assign new_n10432_ = ~pi0039 & ~new_n10431_;
  assign new_n10433_ = ~new_n10390_ & new_n10432_;
  assign new_n10434_ = pi0287 & new_n3100_;
  assign new_n10435_ = new_n10330_ & new_n10434_;
  assign new_n10436_ = ~new_n10331_ & ~new_n10435_;
  assign new_n10437_ = pi0039 & ~new_n10436_;
  assign new_n10438_ = new_n3211_ & ~new_n10437_;
  assign new_n10439_ = ~new_n10433_ & new_n10438_;
  assign new_n10440_ = new_n2498_ & new_n6379_;
  assign new_n10441_ = ~pi0044 & new_n10440_;
  assign new_n10442_ = new_n10308_ & new_n10441_;
  assign new_n10443_ = ~new_n10304_ & ~new_n10442_;
  assign new_n10444_ = ~pi0072 & ~new_n7561_;
  assign new_n10445_ = ~new_n10443_ & ~new_n10444_;
  assign new_n10446_ = ~new_n10306_ & new_n10445_;
  assign new_n10447_ = pi0041 & ~new_n10301_;
  assign new_n10448_ = new_n2733_ & ~new_n10306_;
  assign new_n10449_ = ~new_n10305_ & ~new_n10448_;
  assign new_n10450_ = ~new_n10447_ & ~new_n10449_;
  assign new_n10451_ = ~new_n10446_ & new_n10450_;
  assign new_n10452_ = new_n10298_ & ~new_n10451_;
  assign new_n10453_ = ~new_n10296_ & ~new_n10452_;
  assign new_n10454_ = ~pi0039 & ~new_n10453_;
  assign new_n10455_ = ~new_n10332_ & ~new_n10454_;
  assign new_n10456_ = new_n6258_ & ~new_n10455_;
  assign new_n10457_ = pi0038 & ~new_n10336_;
  assign new_n10458_ = ~pi0087 & ~new_n10457_;
  assign new_n10459_ = ~new_n10456_ & new_n10458_;
  assign new_n10460_ = ~new_n10439_ & new_n10459_;
  assign new_n10461_ = pi0041 & ~new_n10300_;
  assign new_n10462_ = pi0228 & new_n10443_;
  assign new_n10463_ = ~new_n10461_ & new_n10462_;
  assign new_n10464_ = ~pi0228 & new_n10295_;
  assign new_n10465_ = new_n3212_ & ~new_n10464_;
  assign new_n10466_ = ~new_n10463_ & new_n10465_;
  assign new_n10467_ = ~new_n3211_ & new_n10335_;
  assign new_n10468_ = pi0087 & ~new_n10467_;
  assign new_n10469_ = ~new_n10332_ & new_n10468_;
  assign new_n10470_ = ~new_n10466_ & new_n10469_;
  assign new_n10471_ = ~pi0075 & ~new_n10470_;
  assign new_n10472_ = ~new_n10460_ & new_n10471_;
  assign new_n10473_ = ~new_n10339_ & ~new_n10472_;
  assign new_n10474_ = new_n7455_ & ~new_n10473_;
  assign new_n10475_ = ~new_n7455_ & ~new_n10336_;
  assign new_n10476_ = ~po1038 & ~new_n10475_;
  assign new_n10477_ = ~new_n10474_ & new_n10476_;
  assign new_n10478_ = pi0039 & pi0232;
  assign new_n10479_ = new_n10323_ & new_n10478_;
  assign new_n10480_ = ~pi0072 & ~new_n10335_;
  assign new_n10481_ = po1038 & new_n10480_;
  assign new_n10482_ = ~new_n10479_ & new_n10481_;
  assign po0199 = ~new_n10477_ & ~new_n10482_;
  assign new_n10484_ = pi0211 & pi0214;
  assign new_n10485_ = pi0212 & new_n10484_;
  assign new_n10486_ = ~pi0219 & ~new_n10485_;
  assign new_n10487_ = ~pi0115 & new_n2733_;
  assign new_n10488_ = pi0042 & ~pi0114;
  assign new_n10489_ = pi0072 & pi0116;
  assign new_n10490_ = pi0072 & pi0113;
  assign new_n10491_ = pi0072 & ~new_n6265_;
  assign new_n10492_ = ~pi0099 & new_n10375_;
  assign new_n10493_ = ~new_n10491_ & ~new_n10492_;
  assign new_n10494_ = ~pi0113 & ~new_n10493_;
  assign new_n10495_ = ~new_n10490_ & ~new_n10494_;
  assign new_n10496_ = ~pi0116 & ~new_n10495_;
  assign new_n10497_ = ~new_n10489_ & ~new_n10496_;
  assign new_n10498_ = new_n10488_ & ~new_n10497_;
  assign new_n10499_ = pi0042 & ~pi0072;
  assign new_n10500_ = pi0114 & ~new_n10499_;
  assign new_n10501_ = new_n6265_ & new_n10360_;
  assign new_n10502_ = new_n6269_ & new_n10501_;
  assign new_n10503_ = ~pi0042 & ~new_n10502_;
  assign new_n10504_ = ~new_n10500_ & ~new_n10503_;
  assign new_n10505_ = ~new_n10498_ & new_n10504_;
  assign new_n10506_ = new_n10487_ & ~new_n10505_;
  assign new_n10507_ = ~pi0115 & ~new_n2733_;
  assign new_n10508_ = ~pi0099 & new_n10382_;
  assign new_n10509_ = ~new_n10491_ & ~new_n10508_;
  assign new_n10510_ = ~pi0113 & ~new_n10509_;
  assign new_n10511_ = ~new_n10490_ & ~new_n10510_;
  assign new_n10512_ = ~pi0116 & ~new_n10511_;
  assign new_n10513_ = ~new_n10489_ & ~new_n10512_;
  assign new_n10514_ = pi0042 & new_n10513_;
  assign new_n10515_ = new_n6265_ & new_n10385_;
  assign new_n10516_ = new_n6269_ & new_n10515_;
  assign new_n10517_ = ~pi0042 & new_n10516_;
  assign new_n10518_ = ~pi0114 & ~new_n10517_;
  assign new_n10519_ = ~new_n10514_ & new_n10518_;
  assign new_n10520_ = ~new_n10500_ & ~new_n10519_;
  assign new_n10521_ = new_n10507_ & ~new_n10520_;
  assign new_n10522_ = pi0115 & ~new_n10499_;
  assign new_n10523_ = pi0228 & ~new_n10522_;
  assign new_n10524_ = ~new_n10521_ & new_n10523_;
  assign new_n10525_ = ~new_n10506_ & new_n10524_;
  assign new_n10526_ = ~pi0099 & new_n10429_;
  assign new_n10527_ = ~new_n10491_ & ~new_n10526_;
  assign new_n10528_ = ~pi0113 & ~new_n10527_;
  assign new_n10529_ = ~new_n10490_ & ~new_n10528_;
  assign new_n10530_ = ~pi0116 & ~new_n10529_;
  assign new_n10531_ = ~new_n10489_ & ~new_n10530_;
  assign new_n10532_ = new_n10488_ & ~new_n10531_;
  assign new_n10533_ = new_n6265_ & new_n10420_;
  assign new_n10534_ = ~pi0113 & new_n10533_;
  assign new_n10535_ = ~pi0116 & new_n10534_;
  assign new_n10536_ = ~pi0042 & ~new_n10535_;
  assign new_n10537_ = ~new_n10500_ & ~new_n10536_;
  assign new_n10538_ = ~new_n10532_ & new_n10537_;
  assign new_n10539_ = ~pi0115 & ~new_n10538_;
  assign new_n10540_ = ~pi0228 & ~new_n10522_;
  assign new_n10541_ = ~new_n10539_ & new_n10540_;
  assign new_n10542_ = ~pi0039 & ~new_n10541_;
  assign new_n10543_ = ~new_n10525_ & new_n10542_;
  assign new_n10544_ = ~pi0072 & pi0199;
  assign new_n10545_ = ~pi0232 & ~new_n10544_;
  assign new_n10546_ = ~pi0299 & ~new_n10545_;
  assign new_n10547_ = ~pi0072 & ~new_n10325_;
  assign new_n10548_ = new_n6185_ & new_n10434_;
  assign new_n10549_ = ~pi0189 & new_n10548_;
  assign new_n10550_ = ~new_n10547_ & ~new_n10549_;
  assign new_n10551_ = pi0199 & ~new_n10550_;
  assign new_n10552_ = pi0232 & ~new_n10551_;
  assign new_n10553_ = new_n10546_ & ~new_n10552_;
  assign new_n10554_ = pi0039 & ~new_n10553_;
  assign new_n10555_ = ~new_n10543_ & ~new_n10554_;
  assign new_n10556_ = new_n3211_ & ~new_n10555_;
  assign new_n10557_ = ~new_n8100_ & ~new_n10499_;
  assign new_n10558_ = ~new_n10487_ & new_n10499_;
  assign new_n10559_ = new_n8100_ & ~new_n10558_;
  assign new_n10560_ = new_n10487_ & ~new_n10500_;
  assign new_n10561_ = new_n6265_ & new_n10300_;
  assign new_n10562_ = new_n6269_ & new_n10561_;
  assign new_n10563_ = new_n7561_ & new_n10562_;
  assign new_n10564_ = ~pi0114 & ~new_n6268_;
  assign new_n10565_ = new_n10563_ & new_n10564_;
  assign new_n10566_ = ~pi0042 & new_n10565_;
  assign new_n10567_ = new_n6266_ & new_n10441_;
  assign new_n10568_ = new_n6269_ & new_n10567_;
  assign new_n10569_ = ~pi0072 & ~new_n10568_;
  assign new_n10570_ = ~new_n10444_ & ~new_n10569_;
  assign new_n10571_ = pi0042 & ~new_n10570_;
  assign new_n10572_ = ~pi0114 & ~new_n10571_;
  assign new_n10573_ = ~new_n10566_ & new_n10572_;
  assign new_n10574_ = new_n10560_ & ~new_n10573_;
  assign new_n10575_ = new_n10559_ & ~new_n10574_;
  assign new_n10576_ = ~new_n10557_ & ~new_n10575_;
  assign new_n10577_ = ~pi0039 & ~new_n10576_;
  assign new_n10578_ = pi0199 & new_n10547_;
  assign new_n10579_ = pi0232 & ~new_n10578_;
  assign new_n10580_ = new_n10546_ & ~new_n10579_;
  assign new_n10581_ = pi0039 & ~new_n10580_;
  assign new_n10582_ = ~new_n10577_ & ~new_n10581_;
  assign new_n10583_ = new_n6258_ & ~new_n10582_;
  assign new_n10584_ = ~pi0039 & ~new_n10499_;
  assign new_n10585_ = ~new_n10581_ & ~new_n10584_;
  assign new_n10586_ = pi0038 & ~new_n10585_;
  assign new_n10587_ = ~pi0087 & ~new_n10586_;
  assign new_n10588_ = ~new_n10583_ & new_n10587_;
  assign new_n10589_ = ~new_n10556_ & new_n10588_;
  assign new_n10590_ = pi0228 & new_n10562_;
  assign new_n10591_ = ~pi0115 & new_n10590_;
  assign new_n10592_ = ~pi0114 & new_n10591_;
  assign new_n10593_ = ~pi0042 & new_n10592_;
  assign new_n10594_ = pi0228 & new_n10567_;
  assign new_n10595_ = new_n6271_ & new_n10594_;
  assign new_n10596_ = new_n10499_ & ~new_n10595_;
  assign new_n10597_ = new_n3212_ & ~new_n10596_;
  assign new_n10598_ = ~new_n10593_ & new_n10597_;
  assign new_n10599_ = ~new_n3211_ & new_n10584_;
  assign new_n10600_ = pi0087 & ~new_n10599_;
  assign new_n10601_ = ~new_n10598_ & new_n10600_;
  assign new_n10602_ = ~new_n10581_ & new_n10601_;
  assign new_n10603_ = ~pi0075 & ~new_n10602_;
  assign new_n10604_ = ~new_n10589_ & new_n10603_;
  assign new_n10605_ = new_n7502_ & new_n10565_;
  assign new_n10606_ = ~pi0042 & new_n10605_;
  assign new_n10607_ = new_n6266_ & new_n10313_;
  assign new_n10608_ = ~pi0113 & new_n10607_;
  assign new_n10609_ = ~pi0116 & new_n10608_;
  assign new_n10610_ = new_n10499_ & ~new_n10609_;
  assign new_n10611_ = ~pi0114 & ~new_n10610_;
  assign new_n10612_ = ~new_n10606_ & new_n10611_;
  assign new_n10613_ = new_n10560_ & ~new_n10612_;
  assign new_n10614_ = new_n10559_ & ~new_n10613_;
  assign new_n10615_ = new_n3246_ & ~new_n10557_;
  assign new_n10616_ = ~new_n10614_ & new_n10615_;
  assign new_n10617_ = ~new_n3246_ & new_n10499_;
  assign new_n10618_ = ~pi0039 & ~new_n10617_;
  assign new_n10619_ = ~new_n10616_ & new_n10618_;
  assign new_n10620_ = ~new_n10581_ & ~new_n10619_;
  assign new_n10621_ = pi0075 & ~new_n10620_;
  assign new_n10622_ = new_n7455_ & ~new_n10621_;
  assign new_n10623_ = ~new_n10604_ & new_n10622_;
  assign new_n10624_ = pi0207 & pi0208;
  assign new_n10625_ = ~new_n7455_ & new_n10585_;
  assign new_n10626_ = ~new_n10624_ & ~new_n10625_;
  assign new_n10627_ = ~new_n10623_ & new_n10626_;
  assign new_n10628_ = ~pi0072 & pi0200;
  assign new_n10629_ = ~pi0232 & ~new_n10628_;
  assign new_n10630_ = ~pi0299 & ~new_n10629_;
  assign new_n10631_ = pi0200 & new_n10547_;
  assign new_n10632_ = pi0232 & ~new_n10631_;
  assign new_n10633_ = new_n10630_ & ~new_n10632_;
  assign new_n10634_ = pi0039 & ~new_n10633_;
  assign new_n10635_ = ~new_n10580_ & new_n10634_;
  assign new_n10636_ = ~new_n10584_ & ~new_n10635_;
  assign new_n10637_ = ~new_n7455_ & new_n10636_;
  assign new_n10638_ = new_n10624_ & ~new_n10637_;
  assign new_n10639_ = pi0200 & ~new_n10550_;
  assign new_n10640_ = new_n10552_ & ~new_n10639_;
  assign new_n10641_ = ~new_n10546_ & ~new_n10630_;
  assign new_n10642_ = ~new_n10640_ & ~new_n10641_;
  assign new_n10643_ = pi0039 & ~new_n10642_;
  assign new_n10644_ = ~new_n10543_ & ~new_n10643_;
  assign new_n10645_ = new_n3211_ & ~new_n10644_;
  assign new_n10646_ = pi0038 & ~new_n10636_;
  assign new_n10647_ = ~pi0087 & ~new_n10646_;
  assign new_n10648_ = ~new_n10577_ & ~new_n10635_;
  assign new_n10649_ = new_n6258_ & ~new_n10648_;
  assign new_n10650_ = new_n10647_ & ~new_n10649_;
  assign new_n10651_ = ~new_n10645_ & new_n10650_;
  assign new_n10652_ = new_n10601_ & ~new_n10635_;
  assign new_n10653_ = ~pi0075 & ~new_n10652_;
  assign new_n10654_ = ~new_n10651_ & new_n10653_;
  assign new_n10655_ = ~new_n10619_ & ~new_n10635_;
  assign new_n10656_ = pi0075 & ~new_n10655_;
  assign new_n10657_ = new_n7455_ & ~new_n10656_;
  assign new_n10658_ = ~new_n10654_ & new_n10657_;
  assign new_n10659_ = new_n10638_ & ~new_n10658_;
  assign new_n10660_ = ~new_n10627_ & ~new_n10659_;
  assign new_n10661_ = new_n10486_ & ~new_n10660_;
  assign new_n10662_ = pi0232 & ~pi0299;
  assign new_n10663_ = ~new_n10551_ & new_n10662_;
  assign new_n10664_ = new_n10321_ & new_n10434_;
  assign new_n10665_ = ~pi0166 & new_n7499_;
  assign new_n10666_ = ~pi0072 & ~new_n10665_;
  assign new_n10667_ = pi0232 & pi0299;
  assign new_n10668_ = ~new_n10666_ & new_n10667_;
  assign new_n10669_ = ~new_n10664_ & new_n10668_;
  assign new_n10670_ = pi0072 & ~pi0232;
  assign new_n10671_ = pi0299 & ~new_n10670_;
  assign new_n10672_ = new_n10545_ & ~new_n10671_;
  assign new_n10673_ = ~new_n10669_ & ~new_n10672_;
  assign new_n10674_ = ~new_n10663_ & new_n10673_;
  assign new_n10675_ = pi0039 & ~new_n10674_;
  assign new_n10676_ = ~new_n10543_ & ~new_n10675_;
  assign new_n10677_ = new_n3211_ & ~new_n10676_;
  assign new_n10678_ = pi0299 & new_n10666_;
  assign new_n10679_ = pi0039 & ~new_n10678_;
  assign new_n10680_ = ~new_n10580_ & new_n10679_;
  assign new_n10681_ = ~new_n10577_ & ~new_n10680_;
  assign new_n10682_ = new_n6258_ & ~new_n10681_;
  assign new_n10683_ = ~new_n10584_ & ~new_n10680_;
  assign new_n10684_ = pi0038 & ~new_n10683_;
  assign new_n10685_ = ~pi0087 & ~new_n10684_;
  assign new_n10686_ = ~new_n10682_ & new_n10685_;
  assign new_n10687_ = ~new_n10677_ & new_n10686_;
  assign new_n10688_ = new_n10601_ & ~new_n10680_;
  assign new_n10689_ = ~pi0075 & ~new_n10688_;
  assign new_n10690_ = ~new_n10687_ & new_n10689_;
  assign new_n10691_ = ~new_n10619_ & ~new_n10680_;
  assign new_n10692_ = pi0075 & ~new_n10691_;
  assign new_n10693_ = new_n7455_ & ~new_n10692_;
  assign new_n10694_ = ~new_n10690_ & new_n10693_;
  assign new_n10695_ = ~new_n10624_ & ~new_n10694_;
  assign new_n10696_ = ~pi0299 & new_n10640_;
  assign new_n10697_ = ~new_n10628_ & new_n10672_;
  assign new_n10698_ = ~new_n10669_ & ~new_n10697_;
  assign new_n10699_ = ~new_n10696_ & new_n10698_;
  assign new_n10700_ = pi0039 & ~new_n10699_;
  assign new_n10701_ = ~new_n10543_ & ~new_n10700_;
  assign new_n10702_ = new_n3211_ & ~new_n10701_;
  assign new_n10703_ = new_n10634_ & new_n10680_;
  assign new_n10704_ = ~new_n10577_ & ~new_n10703_;
  assign new_n10705_ = new_n6258_ & ~new_n10704_;
  assign new_n10706_ = ~new_n10647_ & ~new_n10685_;
  assign new_n10707_ = ~new_n10705_ & ~new_n10706_;
  assign new_n10708_ = ~new_n10702_ & new_n10707_;
  assign new_n10709_ = new_n10600_ & ~new_n10703_;
  assign new_n10710_ = ~new_n10598_ & new_n10709_;
  assign new_n10711_ = ~pi0075 & ~new_n10710_;
  assign new_n10712_ = ~new_n10708_ & new_n10711_;
  assign new_n10713_ = ~new_n10619_ & ~new_n10703_;
  assign new_n10714_ = pi0075 & ~new_n10713_;
  assign new_n10715_ = new_n7455_ & ~new_n10714_;
  assign new_n10716_ = ~new_n10712_ & new_n10715_;
  assign new_n10717_ = new_n10638_ & ~new_n10716_;
  assign new_n10718_ = ~new_n10695_ & ~new_n10717_;
  assign new_n10719_ = ~new_n7455_ & new_n10683_;
  assign new_n10720_ = ~new_n10486_ & ~new_n10719_;
  assign new_n10721_ = ~new_n10718_ & new_n10720_;
  assign new_n10722_ = ~po1038 & ~new_n10721_;
  assign new_n10723_ = ~new_n10661_ & new_n10722_;
  assign new_n10724_ = ~new_n10486_ & new_n10666_;
  assign new_n10725_ = pi0039 & ~new_n10724_;
  assign new_n10726_ = po1038 & ~new_n10584_;
  assign new_n10727_ = ~new_n10725_ & new_n10726_;
  assign po0200 = new_n10723_ | new_n10727_;
  assign new_n10729_ = pi0212 & pi0214;
  assign new_n10730_ = ~pi0211 & ~pi0219;
  assign new_n10731_ = new_n10729_ & ~new_n10730_;
  assign new_n10732_ = ~pi0211 & ~new_n10729_;
  assign new_n10733_ = ~new_n10731_ & ~new_n10732_;
  assign new_n10734_ = ~new_n2733_ & ~new_n10513_;
  assign new_n10735_ = new_n2733_ & ~new_n10497_;
  assign new_n10736_ = ~new_n10734_ & ~new_n10735_;
  assign new_n10737_ = pi0228 & ~new_n10736_;
  assign new_n10738_ = ~pi0228 & ~new_n10531_;
  assign new_n10739_ = ~new_n10737_ & ~new_n10738_;
  assign new_n10740_ = ~pi0042 & new_n6270_;
  assign new_n10741_ = pi0043 & new_n10740_;
  assign new_n10742_ = ~new_n10739_ & new_n10741_;
  assign new_n10743_ = ~pi0228 & ~new_n10535_;
  assign new_n10744_ = ~new_n2733_ & ~new_n10515_;
  assign new_n10745_ = new_n2733_ & ~new_n10501_;
  assign new_n10746_ = ~new_n10744_ & ~new_n10745_;
  assign new_n10747_ = new_n6269_ & new_n10746_;
  assign new_n10748_ = pi0228 & ~new_n10747_;
  assign new_n10749_ = ~new_n10743_ & ~new_n10748_;
  assign new_n10750_ = ~pi0043 & ~new_n10749_;
  assign new_n10751_ = pi0043 & ~pi0072;
  assign new_n10752_ = ~new_n10740_ & ~new_n10751_;
  assign new_n10753_ = ~new_n10750_ & ~new_n10752_;
  assign new_n10754_ = ~new_n10742_ & new_n10753_;
  assign new_n10755_ = ~pi0039 & ~new_n10754_;
  assign new_n10756_ = ~new_n10639_ & new_n10662_;
  assign new_n10757_ = new_n10629_ & ~new_n10671_;
  assign new_n10758_ = ~new_n10669_ & ~new_n10757_;
  assign new_n10759_ = ~new_n10756_ & new_n10758_;
  assign new_n10760_ = pi0039 & ~new_n10759_;
  assign new_n10761_ = ~new_n10755_ & ~new_n10760_;
  assign new_n10762_ = new_n3211_ & ~new_n10761_;
  assign new_n10763_ = ~new_n8100_ & ~new_n10751_;
  assign new_n10764_ = new_n2733_ & new_n10740_;
  assign new_n10765_ = new_n10751_ & ~new_n10764_;
  assign new_n10766_ = new_n8100_ & ~new_n10765_;
  assign new_n10767_ = ~pi0043 & pi0052;
  assign new_n10768_ = new_n10563_ & new_n10767_;
  assign new_n10769_ = pi0043 & ~new_n10570_;
  assign new_n10770_ = ~new_n10768_ & ~new_n10769_;
  assign new_n10771_ = new_n10764_ & ~new_n10770_;
  assign new_n10772_ = new_n10766_ & ~new_n10771_;
  assign new_n10773_ = ~new_n10763_ & ~new_n10772_;
  assign new_n10774_ = ~pi0039 & ~new_n10773_;
  assign new_n10775_ = ~new_n10633_ & new_n10679_;
  assign new_n10776_ = ~new_n10774_ & ~new_n10775_;
  assign new_n10777_ = new_n6258_ & ~new_n10776_;
  assign new_n10778_ = ~pi0039 & ~new_n10751_;
  assign new_n10779_ = ~new_n10775_ & ~new_n10778_;
  assign new_n10780_ = pi0038 & ~new_n10779_;
  assign new_n10781_ = ~pi0087 & ~new_n10780_;
  assign new_n10782_ = ~new_n10777_ & new_n10781_;
  assign new_n10783_ = ~new_n10762_ & new_n10782_;
  assign new_n10784_ = ~pi0043 & ~new_n10562_;
  assign new_n10785_ = pi0043 & ~new_n10569_;
  assign new_n10786_ = pi0228 & new_n10740_;
  assign new_n10787_ = ~new_n10785_ & new_n10786_;
  assign new_n10788_ = ~new_n10784_ & new_n10787_;
  assign new_n10789_ = new_n10751_ & ~new_n10786_;
  assign new_n10790_ = new_n3212_ & ~new_n10789_;
  assign new_n10791_ = ~new_n10788_ & new_n10790_;
  assign new_n10792_ = ~new_n3211_ & new_n10778_;
  assign new_n10793_ = pi0087 & ~new_n10792_;
  assign new_n10794_ = ~new_n10791_ & new_n10793_;
  assign new_n10795_ = ~new_n10775_ & new_n10794_;
  assign new_n10796_ = ~pi0075 & ~new_n10795_;
  assign new_n10797_ = ~new_n10783_ & new_n10796_;
  assign new_n10798_ = ~pi0072 & ~new_n10609_;
  assign new_n10799_ = pi0043 & new_n10798_;
  assign new_n10800_ = new_n7502_ & new_n10563_;
  assign new_n10801_ = new_n10767_ & new_n10800_;
  assign new_n10802_ = ~new_n10799_ & ~new_n10801_;
  assign new_n10803_ = new_n10764_ & ~new_n10802_;
  assign new_n10804_ = new_n10766_ & ~new_n10803_;
  assign new_n10805_ = ~new_n10763_ & ~new_n10804_;
  assign new_n10806_ = ~pi0039 & ~new_n10805_;
  assign new_n10807_ = new_n3246_ & ~new_n10806_;
  assign new_n10808_ = ~new_n3246_ & ~new_n10778_;
  assign new_n10809_ = ~new_n10807_ & ~new_n10808_;
  assign new_n10810_ = ~new_n10775_ & ~new_n10809_;
  assign new_n10811_ = pi0075 & ~new_n10810_;
  assign new_n10812_ = new_n7455_ & ~new_n10811_;
  assign new_n10813_ = ~new_n10797_ & new_n10812_;
  assign new_n10814_ = ~new_n7455_ & new_n10779_;
  assign new_n10815_ = ~new_n10624_ & ~new_n10814_;
  assign new_n10816_ = ~new_n10813_ & new_n10815_;
  assign new_n10817_ = ~pi0199 & ~pi0200;
  assign new_n10818_ = ~new_n10550_ & new_n10817_;
  assign new_n10819_ = new_n10662_ & ~new_n10818_;
  assign new_n10820_ = ~pi0299 & ~new_n10817_;
  assign new_n10821_ = ~pi0072 & ~new_n10820_;
  assign new_n10822_ = ~pi0232 & ~new_n10821_;
  assign new_n10823_ = ~new_n10669_ & ~new_n10822_;
  assign new_n10824_ = ~new_n10819_ & new_n10823_;
  assign new_n10825_ = pi0039 & ~new_n10824_;
  assign new_n10826_ = ~new_n10755_ & ~new_n10825_;
  assign new_n10827_ = new_n3211_ & ~new_n10826_;
  assign new_n10828_ = ~pi0299 & ~new_n10822_;
  assign new_n10829_ = new_n10547_ & new_n10817_;
  assign new_n10830_ = pi0232 & ~new_n10829_;
  assign new_n10831_ = new_n10828_ & ~new_n10830_;
  assign new_n10832_ = pi0039 & ~new_n10831_;
  assign new_n10833_ = ~new_n10678_ & new_n10832_;
  assign new_n10834_ = ~new_n10774_ & ~new_n10833_;
  assign new_n10835_ = new_n6258_ & ~new_n10834_;
  assign new_n10836_ = ~new_n10778_ & ~new_n10833_;
  assign new_n10837_ = pi0038 & ~new_n10836_;
  assign new_n10838_ = ~pi0087 & ~new_n10837_;
  assign new_n10839_ = ~new_n10835_ & new_n10838_;
  assign new_n10840_ = ~new_n10827_ & new_n10839_;
  assign new_n10841_ = new_n10794_ & ~new_n10833_;
  assign new_n10842_ = ~pi0075 & ~new_n10841_;
  assign new_n10843_ = ~new_n10840_ & new_n10842_;
  assign new_n10844_ = ~new_n10809_ & ~new_n10833_;
  assign new_n10845_ = pi0075 & ~new_n10844_;
  assign new_n10846_ = new_n7455_ & ~new_n10845_;
  assign new_n10847_ = ~new_n10843_ & new_n10846_;
  assign new_n10848_ = ~new_n7455_ & new_n10836_;
  assign new_n10849_ = new_n10624_ & ~new_n10848_;
  assign new_n10850_ = ~new_n10847_ & new_n10849_;
  assign new_n10851_ = ~new_n10816_ & ~new_n10850_;
  assign new_n10852_ = new_n10733_ & ~new_n10851_;
  assign new_n10853_ = pi0232 & ~new_n10639_;
  assign new_n10854_ = new_n10630_ & ~new_n10853_;
  assign new_n10855_ = pi0039 & ~new_n10854_;
  assign new_n10856_ = ~new_n10755_ & ~new_n10855_;
  assign new_n10857_ = new_n3211_ & ~new_n10856_;
  assign new_n10858_ = ~new_n10634_ & ~new_n10774_;
  assign new_n10859_ = new_n6258_ & ~new_n10858_;
  assign new_n10860_ = ~new_n10634_ & ~new_n10778_;
  assign new_n10861_ = pi0038 & ~new_n10860_;
  assign new_n10862_ = ~pi0087 & ~new_n10861_;
  assign new_n10863_ = ~new_n10859_ & new_n10862_;
  assign new_n10864_ = ~new_n10857_ & new_n10863_;
  assign new_n10865_ = ~new_n10634_ & new_n10794_;
  assign new_n10866_ = ~pi0075 & ~new_n10865_;
  assign new_n10867_ = ~new_n10864_ & new_n10866_;
  assign new_n10868_ = ~new_n10634_ & ~new_n10809_;
  assign new_n10869_ = pi0075 & ~new_n10868_;
  assign new_n10870_ = new_n7455_ & ~new_n10869_;
  assign new_n10871_ = ~new_n10867_ & new_n10870_;
  assign new_n10872_ = ~new_n7455_ & new_n10860_;
  assign new_n10873_ = ~new_n10624_ & ~new_n10872_;
  assign new_n10874_ = ~new_n10871_ & new_n10873_;
  assign new_n10875_ = pi0232 & ~new_n10818_;
  assign new_n10876_ = new_n10828_ & ~new_n10875_;
  assign new_n10877_ = pi0039 & ~new_n10876_;
  assign new_n10878_ = ~new_n10755_ & ~new_n10877_;
  assign new_n10879_ = new_n3211_ & ~new_n10878_;
  assign new_n10880_ = ~new_n10774_ & ~new_n10832_;
  assign new_n10881_ = new_n6258_ & ~new_n10880_;
  assign new_n10882_ = ~new_n10778_ & ~new_n10832_;
  assign new_n10883_ = pi0038 & ~new_n10882_;
  assign new_n10884_ = ~pi0087 & ~new_n10883_;
  assign new_n10885_ = ~new_n10881_ & new_n10884_;
  assign new_n10886_ = ~new_n10879_ & new_n10885_;
  assign new_n10887_ = ~new_n3281_ & ~new_n10882_;
  assign new_n10888_ = new_n10794_ & ~new_n10887_;
  assign new_n10889_ = ~pi0075 & ~new_n10888_;
  assign new_n10890_ = ~new_n10886_ & new_n10889_;
  assign new_n10891_ = ~new_n10809_ & ~new_n10832_;
  assign new_n10892_ = pi0075 & ~new_n10891_;
  assign new_n10893_ = new_n7455_ & ~new_n10892_;
  assign new_n10894_ = ~new_n10890_ & new_n10893_;
  assign new_n10895_ = ~new_n7455_ & new_n10882_;
  assign new_n10896_ = new_n10624_ & ~new_n10895_;
  assign new_n10897_ = ~new_n10894_ & new_n10896_;
  assign new_n10898_ = ~new_n10874_ & ~new_n10897_;
  assign new_n10899_ = ~new_n10733_ & ~new_n10898_;
  assign new_n10900_ = ~po1038 & ~new_n10899_;
  assign new_n10901_ = ~new_n10852_ & new_n10900_;
  assign new_n10902_ = new_n10666_ & new_n10733_;
  assign new_n10903_ = pi0039 & ~new_n10902_;
  assign new_n10904_ = po1038 & ~new_n10778_;
  assign new_n10905_ = ~new_n10903_ & new_n10904_;
  assign po0201 = new_n10901_ | new_n10905_;
  assign new_n10907_ = pi0044 & ~pi0072;
  assign new_n10908_ = ~new_n8100_ & ~new_n10907_;
  assign new_n10909_ = ~pi0039 & ~new_n10908_;
  assign new_n10910_ = ~new_n2733_ & new_n10907_;
  assign new_n10911_ = new_n8100_ & ~new_n10910_;
  assign new_n10912_ = new_n7504_ & ~new_n10362_;
  assign new_n10913_ = new_n7561_ & new_n10299_;
  assign new_n10914_ = new_n7502_ & new_n10913_;
  assign new_n10915_ = pi0044 & ~new_n10312_;
  assign new_n10916_ = ~new_n10914_ & ~new_n10915_;
  assign new_n10917_ = new_n10912_ & ~new_n10916_;
  assign new_n10918_ = new_n10911_ & ~new_n10917_;
  assign new_n10919_ = new_n10909_ & ~new_n10918_;
  assign new_n10920_ = pi0039 & new_n7500_;
  assign new_n10921_ = ~pi0072 & new_n10920_;
  assign new_n10922_ = ~new_n10919_ & ~new_n10921_;
  assign new_n10923_ = new_n3246_ & ~new_n10922_;
  assign new_n10924_ = ~pi0072 & new_n7500_;
  assign new_n10925_ = pi0039 & ~new_n10924_;
  assign new_n10926_ = ~pi0039 & ~new_n10907_;
  assign new_n10927_ = ~new_n10925_ & ~new_n10926_;
  assign new_n10928_ = ~new_n3246_ & new_n10927_;
  assign new_n10929_ = pi0075 & ~new_n10928_;
  assign new_n10930_ = ~new_n10923_ & new_n10929_;
  assign new_n10931_ = pi0044 & new_n10371_;
  assign new_n10932_ = new_n2733_ & ~new_n10359_;
  assign new_n10933_ = ~new_n10931_ & new_n10932_;
  assign new_n10934_ = pi0044 & new_n10378_;
  assign new_n10935_ = ~new_n2733_ & ~new_n10384_;
  assign new_n10936_ = ~new_n10934_ & new_n10935_;
  assign new_n10937_ = ~new_n10933_ & ~new_n10936_;
  assign new_n10938_ = pi0228 & ~new_n10937_;
  assign new_n10939_ = pi0044 & new_n10425_;
  assign new_n10940_ = ~pi0228 & ~new_n10939_;
  assign new_n10941_ = ~new_n10419_ & new_n10940_;
  assign new_n10942_ = ~pi0039 & ~new_n10941_;
  assign new_n10943_ = ~new_n10938_ & new_n10942_;
  assign new_n10944_ = pi0287 & new_n10440_;
  assign new_n10945_ = ~pi0072 & ~new_n10944_;
  assign new_n10946_ = new_n10920_ & new_n10945_;
  assign new_n10947_ = new_n3211_ & ~new_n10946_;
  assign new_n10948_ = ~new_n10943_ & new_n10947_;
  assign new_n10949_ = new_n7561_ & new_n10440_;
  assign new_n10950_ = pi0044 & ~new_n10949_;
  assign new_n10951_ = ~new_n10913_ & ~new_n10950_;
  assign new_n10952_ = new_n10912_ & ~new_n10951_;
  assign new_n10953_ = new_n10911_ & ~new_n10952_;
  assign new_n10954_ = new_n10909_ & ~new_n10953_;
  assign new_n10955_ = new_n6258_ & ~new_n10921_;
  assign new_n10956_ = ~new_n10954_ & new_n10955_;
  assign new_n10957_ = pi0038 & ~new_n10927_;
  assign new_n10958_ = ~pi0087 & ~new_n10957_;
  assign new_n10959_ = ~new_n10956_ & new_n10958_;
  assign new_n10960_ = ~new_n10948_ & new_n10959_;
  assign new_n10961_ = pi0228 & new_n3211_;
  assign new_n10962_ = new_n10299_ & new_n10961_;
  assign new_n10963_ = new_n10440_ & new_n10961_;
  assign new_n10964_ = new_n10907_ & ~new_n10963_;
  assign new_n10965_ = ~pi0039 & ~new_n10964_;
  assign new_n10966_ = ~new_n10962_ & new_n10965_;
  assign new_n10967_ = pi0087 & ~new_n10925_;
  assign new_n10968_ = ~new_n10966_ & new_n10967_;
  assign new_n10969_ = ~pi0075 & ~new_n10968_;
  assign new_n10970_ = ~new_n10960_ & new_n10969_;
  assign new_n10971_ = ~new_n10930_ & ~new_n10970_;
  assign new_n10972_ = new_n7455_ & ~new_n10971_;
  assign new_n10973_ = ~new_n7455_ & ~new_n10927_;
  assign new_n10974_ = ~po1038 & ~new_n10973_;
  assign new_n10975_ = ~new_n10972_ & new_n10974_;
  assign new_n10976_ = new_n2448_ & new_n7499_;
  assign new_n10977_ = ~pi0072 & new_n10976_;
  assign new_n10978_ = pi0039 & ~new_n10977_;
  assign new_n10979_ = po1038 & ~new_n10926_;
  assign new_n10980_ = ~new_n10978_ & new_n10979_;
  assign po0202 = new_n10975_ | new_n10980_;
  assign new_n10982_ = ~pi0038 & pi0039;
  assign new_n10983_ = new_n10197_ & new_n10982_;
  assign new_n10984_ = pi0979 & new_n10983_;
  assign po0203 = new_n6454_ & new_n10984_;
  assign new_n10986_ = ~pi0049 & ~pi0076;
  assign new_n10987_ = new_n8911_ & new_n10986_;
  assign new_n10988_ = ~pi0102 & ~pi0104;
  assign new_n10989_ = ~pi0111 & new_n10988_;
  assign new_n10990_ = new_n10177_ & new_n10989_;
  assign new_n10991_ = new_n10987_ & new_n10990_;
  assign new_n10992_ = pi0061 & ~pi0082;
  assign new_n10993_ = ~pi0083 & ~pi0089;
  assign new_n10994_ = new_n10992_ & new_n10993_;
  assign new_n10995_ = new_n7463_ & new_n8925_;
  assign new_n10996_ = new_n10994_ & new_n10995_;
  assign new_n10997_ = new_n8923_ & new_n10996_;
  assign new_n10998_ = new_n10242_ & new_n10997_;
  assign new_n10999_ = new_n10991_ & new_n10998_;
  assign new_n11000_ = new_n8932_ & new_n10999_;
  assign new_n11001_ = ~pi0841 & new_n11000_;
  assign new_n11002_ = new_n2491_ & new_n2697_;
  assign new_n11003_ = pi0024 & new_n11002_;
  assign new_n11004_ = ~new_n11001_ & ~new_n11003_;
  assign po0204 = new_n10166_ & ~new_n11004_;
  assign new_n11006_ = ~new_n2679_ & new_n7463_;
  assign new_n11007_ = ~pi0082 & new_n2463_;
  assign new_n11008_ = ~pi0084 & pi0104;
  assign new_n11009_ = new_n2607_ & new_n11008_;
  assign new_n11010_ = new_n10181_ & new_n11009_;
  assign new_n11011_ = new_n11007_ & new_n11010_;
  assign new_n11012_ = ~pi0036 & ~new_n11011_;
  assign new_n11013_ = new_n8924_ & new_n9039_;
  assign new_n11014_ = ~pi0067 & ~pi0103;
  assign new_n11015_ = new_n2476_ & new_n11014_;
  assign new_n11016_ = ~pi0098 & new_n11015_;
  assign new_n11017_ = new_n11013_ & new_n11016_;
  assign new_n11018_ = ~new_n11012_ & new_n11017_;
  assign new_n11019_ = ~new_n2648_ & new_n11018_;
  assign new_n11020_ = ~pi0088 & ~new_n11019_;
  assign new_n11021_ = new_n2532_ & ~new_n11020_;
  assign new_n11022_ = new_n11006_ & new_n11021_;
  assign new_n11023_ = new_n2489_ & new_n11022_;
  assign new_n11024_ = ~new_n10159_ & ~new_n11023_;
  assign new_n11025_ = new_n10162_ & ~new_n11024_;
  assign new_n11026_ = new_n7574_ & ~new_n11025_;
  assign new_n11027_ = ~new_n2799_ & new_n11025_;
  assign new_n11028_ = ~pi0036 & new_n11018_;
  assign new_n11029_ = ~pi0088 & ~new_n11028_;
  assign new_n11030_ = new_n11006_ & ~new_n11029_;
  assign new_n11031_ = new_n10176_ & new_n11030_;
  assign new_n11032_ = ~pi0824 & new_n2799_;
  assign new_n11033_ = new_n11031_ & new_n11032_;
  assign new_n11034_ = pi0829 & ~new_n11033_;
  assign new_n11035_ = ~new_n11027_ & new_n11034_;
  assign new_n11036_ = ~new_n2732_ & new_n11035_;
  assign new_n11037_ = ~new_n11026_ & ~new_n11036_;
  assign new_n11038_ = pi1091 & ~new_n11037_;
  assign new_n11039_ = ~new_n7511_ & new_n11025_;
  assign new_n11040_ = ~pi0829 & ~new_n11039_;
  assign new_n11041_ = ~new_n11035_ & ~new_n11040_;
  assign new_n11042_ = ~pi1093 & ~new_n11041_;
  assign new_n11043_ = new_n7511_ & new_n10162_;
  assign new_n11044_ = ~new_n10160_ & new_n11043_;
  assign new_n11045_ = ~new_n6468_ & ~new_n7572_;
  assign new_n11046_ = ~new_n11044_ & ~new_n11045_;
  assign new_n11047_ = ~new_n11039_ & new_n11046_;
  assign new_n11048_ = new_n10165_ & ~new_n11047_;
  assign new_n11049_ = ~new_n11042_ & new_n11048_;
  assign po0205 = ~new_n11038_ & new_n11049_;
  assign new_n11051_ = ~pi0072 & pi0841;
  assign new_n11052_ = new_n2494_ & new_n11051_;
  assign new_n11053_ = ~pi0051 & new_n11052_;
  assign new_n11054_ = new_n10249_ & new_n11053_;
  assign new_n11055_ = new_n10165_ & new_n11054_;
  assign po0206 = new_n10175_ & new_n11055_;
  assign new_n11057_ = pi0074 & ~new_n8962_;
  assign new_n11058_ = ~pi0103 & new_n2641_;
  assign new_n11059_ = new_n10240_ & new_n11058_;
  assign new_n11060_ = new_n8911_ & new_n8924_;
  assign new_n11061_ = new_n11059_ & new_n11060_;
  assign new_n11062_ = new_n2453_ & new_n2476_;
  assign new_n11063_ = ~pi0045 & pi0049;
  assign new_n11064_ = new_n10989_ & new_n11063_;
  assign new_n11065_ = new_n11062_ & new_n11064_;
  assign new_n11066_ = new_n11061_ & new_n11065_;
  assign new_n11067_ = new_n11007_ & new_n11066_;
  assign new_n11068_ = new_n2495_ & new_n8932_;
  assign new_n11069_ = new_n11067_ & new_n11068_;
  assign new_n11070_ = new_n10161_ & new_n11052_;
  assign new_n11071_ = new_n11069_ & new_n11070_;
  assign new_n11072_ = ~pi0074 & ~new_n11071_;
  assign new_n11073_ = new_n7390_ & ~po1038;
  assign new_n11074_ = ~new_n11072_ & new_n11073_;
  assign po0207 = ~new_n11057_ & new_n11074_;
  assign new_n11076_ = pi0024 & new_n8899_;
  assign new_n11077_ = ~new_n10401_ & ~new_n11076_;
  assign new_n11078_ = pi0024 & ~pi0094;
  assign new_n11079_ = ~new_n8897_ & new_n11078_;
  assign new_n11080_ = ~pi0252 & ~new_n8888_;
  assign new_n11081_ = pi0252 & ~po0840;
  assign new_n11082_ = ~new_n11080_ & ~new_n11081_;
  assign new_n11083_ = new_n10162_ & new_n11082_;
  assign new_n11084_ = ~new_n11079_ & new_n11083_;
  assign new_n11085_ = ~new_n11077_ & new_n11084_;
  assign new_n11086_ = new_n2535_ & new_n7476_;
  assign new_n11087_ = pi0024 & ~pi0090;
  assign new_n11088_ = new_n11086_ & new_n11087_;
  assign new_n11089_ = ~new_n11082_ & new_n11088_;
  assign new_n11090_ = new_n8901_ & new_n11089_;
  assign new_n11091_ = ~new_n11085_ & ~new_n11090_;
  assign new_n11092_ = ~pi0100 & ~new_n11091_;
  assign new_n11093_ = pi0100 & ~new_n6263_;
  assign new_n11094_ = new_n6504_ & new_n11093_;
  assign new_n11095_ = ~new_n11092_ & ~new_n11094_;
  assign new_n11096_ = new_n3186_ & new_n3235_;
  assign new_n11097_ = ~new_n11095_ & new_n11096_;
  assign new_n11098_ = new_n6282_ & new_n8967_;
  assign new_n11099_ = new_n8963_ & new_n11098_;
  assign new_n11100_ = ~new_n11097_ & ~new_n11099_;
  assign po0208 = new_n8881_ & ~new_n11100_;
  assign new_n11102_ = new_n2489_ & new_n10166_;
  assign new_n11103_ = new_n2532_ & new_n11102_;
  assign new_n11104_ = new_n9040_ & new_n11062_;
  assign new_n11105_ = new_n2456_ & new_n11104_;
  assign new_n11106_ = ~pi0069 & new_n11105_;
  assign new_n11107_ = new_n2641_ & new_n11106_;
  assign new_n11108_ = new_n2643_ & new_n11107_;
  assign po0209 = new_n11103_ & new_n11108_;
  assign new_n11110_ = ~pi0219 & new_n10732_;
  assign new_n11111_ = pi0052 & ~pi0072;
  assign new_n11112_ = ~pi0039 & new_n11111_;
  assign new_n11113_ = pi0038 & ~new_n11112_;
  assign new_n11114_ = new_n6267_ & new_n6270_;
  assign new_n11115_ = pi0228 & new_n11114_;
  assign new_n11116_ = ~pi0052 & new_n10562_;
  assign new_n11117_ = pi0052 & new_n10569_;
  assign new_n11118_ = ~new_n11116_ & ~new_n11117_;
  assign new_n11119_ = new_n11115_ & ~new_n11118_;
  assign new_n11120_ = new_n11111_ & ~new_n11115_;
  assign new_n11121_ = ~new_n11119_ & ~new_n11120_;
  assign new_n11122_ = ~pi0038 & new_n11121_;
  assign new_n11123_ = ~new_n11113_ & ~new_n11122_;
  assign new_n11124_ = ~pi0100 & ~new_n11123_;
  assign new_n11125_ = pi0100 & ~new_n11112_;
  assign new_n11126_ = ~pi0100 & new_n10982_;
  assign new_n11127_ = pi0087 & ~new_n11126_;
  assign new_n11128_ = ~new_n11125_ & new_n11127_;
  assign new_n11129_ = ~new_n11124_ & new_n11128_;
  assign new_n11130_ = ~pi0114 & new_n6267_;
  assign new_n11131_ = pi0052 & new_n10497_;
  assign new_n11132_ = ~pi0052 & new_n10502_;
  assign new_n11133_ = new_n10487_ & ~new_n11132_;
  assign new_n11134_ = ~new_n11131_ & new_n11133_;
  assign new_n11135_ = pi0052 & new_n10513_;
  assign new_n11136_ = ~pi0052 & new_n10516_;
  assign new_n11137_ = new_n10507_ & ~new_n11136_;
  assign new_n11138_ = ~new_n11135_ & new_n11137_;
  assign new_n11139_ = ~new_n11134_ & ~new_n11138_;
  assign new_n11140_ = new_n11130_ & ~new_n11139_;
  assign new_n11141_ = ~new_n11111_ & ~new_n11114_;
  assign new_n11142_ = pi0228 & ~new_n11141_;
  assign new_n11143_ = ~new_n11140_ & new_n11142_;
  assign new_n11144_ = pi0052 & new_n10531_;
  assign new_n11145_ = ~pi0052 & new_n10535_;
  assign new_n11146_ = new_n11114_ & ~new_n11145_;
  assign new_n11147_ = ~new_n11144_ & new_n11146_;
  assign new_n11148_ = ~pi0228 & ~new_n11141_;
  assign new_n11149_ = ~new_n11147_ & new_n11148_;
  assign new_n11150_ = ~pi0039 & ~new_n11149_;
  assign new_n11151_ = ~new_n11143_ & new_n11150_;
  assign new_n11152_ = ~pi0100 & new_n11151_;
  assign new_n11153_ = new_n8100_ & new_n10487_;
  assign new_n11154_ = new_n11130_ & new_n11153_;
  assign new_n11155_ = new_n7561_ & new_n11154_;
  assign new_n11156_ = new_n10568_ & new_n11155_;
  assign new_n11157_ = new_n11111_ & ~new_n11156_;
  assign new_n11158_ = pi0100 & ~new_n11157_;
  assign new_n11159_ = ~pi0039 & ~new_n11158_;
  assign new_n11160_ = ~new_n11152_ & new_n11159_;
  assign new_n11161_ = ~pi0038 & ~new_n11160_;
  assign new_n11162_ = ~pi0087 & ~new_n11113_;
  assign new_n11163_ = ~new_n11161_ & new_n11162_;
  assign new_n11164_ = ~new_n11129_ & ~new_n11163_;
  assign new_n11165_ = ~pi0075 & ~new_n11164_;
  assign new_n11166_ = new_n10609_ & new_n11154_;
  assign new_n11167_ = new_n3246_ & new_n11166_;
  assign new_n11168_ = new_n11112_ & ~new_n11167_;
  assign new_n11169_ = pi0075 & new_n11168_;
  assign new_n11170_ = new_n7455_ & ~new_n11169_;
  assign new_n11171_ = ~new_n11165_ & new_n11170_;
  assign new_n11172_ = ~new_n7455_ & ~new_n11112_;
  assign new_n11173_ = new_n10624_ & ~new_n11172_;
  assign new_n11174_ = ~new_n11171_ & new_n11173_;
  assign new_n11175_ = ~new_n10877_ & ~new_n11151_;
  assign new_n11176_ = new_n3211_ & ~new_n11175_;
  assign new_n11177_ = ~pi0039 & ~new_n11157_;
  assign new_n11178_ = ~new_n10832_ & ~new_n11177_;
  assign new_n11179_ = new_n6258_ & ~new_n11178_;
  assign new_n11180_ = ~pi0039 & ~new_n11111_;
  assign new_n11181_ = ~new_n10832_ & ~new_n11180_;
  assign new_n11182_ = pi0038 & ~new_n11181_;
  assign new_n11183_ = ~pi0087 & ~new_n11182_;
  assign new_n11184_ = ~new_n11179_ & new_n11183_;
  assign new_n11185_ = ~new_n11176_ & new_n11184_;
  assign new_n11186_ = ~new_n3211_ & new_n11181_;
  assign new_n11187_ = ~pi0039 & new_n11121_;
  assign new_n11188_ = new_n3211_ & ~new_n10832_;
  assign new_n11189_ = ~new_n11187_ & new_n11188_;
  assign new_n11190_ = ~new_n11186_ & ~new_n11189_;
  assign new_n11191_ = pi0087 & ~new_n11190_;
  assign new_n11192_ = ~pi0075 & ~new_n11191_;
  assign new_n11193_ = ~new_n11185_ & new_n11192_;
  assign new_n11194_ = new_n11111_ & ~new_n11166_;
  assign new_n11195_ = ~pi0039 & ~new_n11194_;
  assign new_n11196_ = new_n3246_ & ~new_n10832_;
  assign new_n11197_ = ~new_n11195_ & new_n11196_;
  assign new_n11198_ = ~new_n3246_ & new_n11181_;
  assign new_n11199_ = pi0075 & ~new_n11198_;
  assign new_n11200_ = ~new_n11197_ & new_n11199_;
  assign new_n11201_ = new_n7455_ & ~new_n10624_;
  assign new_n11202_ = ~new_n11200_ & new_n11201_;
  assign new_n11203_ = ~new_n11193_ & new_n11202_;
  assign new_n11204_ = ~new_n11174_ & ~new_n11203_;
  assign new_n11205_ = ~new_n11110_ & ~new_n11204_;
  assign new_n11206_ = ~new_n10669_ & new_n10671_;
  assign new_n11207_ = pi0039 & ~new_n11206_;
  assign new_n11208_ = ~new_n11151_ & ~new_n11207_;
  assign new_n11209_ = new_n3211_ & ~new_n11208_;
  assign new_n11210_ = ~new_n10679_ & ~new_n11180_;
  assign new_n11211_ = pi0038 & ~new_n11210_;
  assign new_n11212_ = ~new_n10679_ & ~new_n11177_;
  assign new_n11213_ = new_n6258_ & ~new_n11212_;
  assign new_n11214_ = ~new_n11211_ & ~new_n11213_;
  assign new_n11215_ = ~new_n11209_ & new_n11214_;
  assign new_n11216_ = ~pi0087 & ~new_n11215_;
  assign new_n11217_ = ~new_n3211_ & new_n11210_;
  assign new_n11218_ = pi0087 & ~new_n11217_;
  assign new_n11219_ = new_n3211_ & ~new_n10679_;
  assign new_n11220_ = ~new_n11187_ & new_n11219_;
  assign new_n11221_ = new_n11218_ & ~new_n11220_;
  assign new_n11222_ = new_n10624_ & ~new_n11221_;
  assign new_n11223_ = ~new_n11216_ & new_n11222_;
  assign new_n11224_ = ~new_n10825_ & ~new_n11151_;
  assign new_n11225_ = new_n3211_ & ~new_n11224_;
  assign new_n11226_ = ~new_n10833_ & ~new_n11177_;
  assign new_n11227_ = new_n6258_ & ~new_n11226_;
  assign new_n11228_ = new_n11182_ & ~new_n11210_;
  assign new_n11229_ = ~new_n11227_ & ~new_n11228_;
  assign new_n11230_ = ~new_n11225_ & new_n11229_;
  assign new_n11231_ = ~pi0087 & ~new_n11230_;
  assign new_n11232_ = new_n3211_ & ~new_n10833_;
  assign new_n11233_ = ~new_n11187_ & new_n11232_;
  assign new_n11234_ = ~new_n11186_ & new_n11218_;
  assign new_n11235_ = ~new_n11233_ & new_n11234_;
  assign new_n11236_ = ~new_n10624_ & ~new_n11235_;
  assign new_n11237_ = ~new_n11231_ & new_n11236_;
  assign new_n11238_ = ~new_n11223_ & ~new_n11237_;
  assign new_n11239_ = ~pi0075 & ~new_n11238_;
  assign new_n11240_ = ~pi0039 & ~new_n11168_;
  assign new_n11241_ = ~new_n10624_ & new_n10833_;
  assign new_n11242_ = new_n10624_ & new_n10679_;
  assign new_n11243_ = pi0075 & ~new_n11242_;
  assign new_n11244_ = ~new_n11241_ & new_n11243_;
  assign new_n11245_ = ~new_n11240_ & new_n11244_;
  assign new_n11246_ = new_n7455_ & ~new_n11245_;
  assign new_n11247_ = ~new_n11239_ & new_n11246_;
  assign new_n11248_ = ~new_n7455_ & ~new_n11210_;
  assign new_n11249_ = new_n11110_ & ~new_n11248_;
  assign new_n11250_ = ~new_n11247_ & new_n11249_;
  assign new_n11251_ = ~new_n7455_ & ~new_n10624_;
  assign new_n11252_ = new_n11181_ & new_n11251_;
  assign new_n11253_ = ~po1038 & ~new_n11252_;
  assign new_n11254_ = ~new_n11250_ & new_n11253_;
  assign new_n11255_ = ~new_n11205_ & new_n11254_;
  assign new_n11256_ = pi0039 & new_n11110_;
  assign new_n11257_ = new_n10666_ & new_n11256_;
  assign new_n11258_ = po1038 & ~new_n11112_;
  assign new_n11259_ = ~new_n11257_ & new_n11258_;
  assign po0210 = ~new_n11255_ & ~new_n11259_;
  assign new_n11261_ = pi0024 & new_n10162_;
  assign new_n11262_ = pi0053 & new_n2505_;
  assign new_n11263_ = new_n2514_ & new_n11262_;
  assign new_n11264_ = new_n2506_ & new_n11263_;
  assign new_n11265_ = new_n11261_ & new_n11264_;
  assign new_n11266_ = ~pi0039 & ~new_n11265_;
  assign new_n11267_ = ~pi0287 & ~pi0979;
  assign new_n11268_ = new_n6186_ & new_n11267_;
  assign new_n11269_ = pi0039 & ~new_n11268_;
  assign new_n11270_ = new_n10200_ & ~new_n11269_;
  assign new_n11271_ = ~new_n11266_ & new_n11270_;
  assign po0211 = ~new_n3357_ & new_n11271_;
  assign new_n11273_ = new_n3247_ & new_n10171_;
  assign new_n11274_ = pi0054 & ~new_n11273_;
  assign new_n11275_ = new_n8899_ & new_n9045_;
  assign new_n11276_ = ~pi0060 & ~pi0085;
  assign new_n11277_ = pi0106 & new_n11276_;
  assign new_n11278_ = new_n2468_ & new_n8915_;
  assign new_n11279_ = new_n11277_ & new_n11278_;
  assign new_n11280_ = new_n10987_ & new_n11279_;
  assign new_n11281_ = new_n8928_ & new_n11059_;
  assign new_n11282_ = new_n11280_ & new_n11281_;
  assign new_n11283_ = new_n11062_ & new_n11282_;
  assign new_n11284_ = new_n11275_ & new_n11283_;
  assign new_n11285_ = ~pi0841 & new_n2493_;
  assign new_n11286_ = new_n8960_ & new_n11285_;
  assign new_n11287_ = new_n2495_ & new_n3243_;
  assign new_n11288_ = new_n11286_ & new_n11287_;
  assign new_n11289_ = new_n11284_ & new_n11288_;
  assign new_n11290_ = ~pi0054 & ~new_n11289_;
  assign new_n11291_ = new_n8880_ & ~new_n11290_;
  assign po0212 = ~new_n11274_ & new_n11291_;
  assign new_n11293_ = ~pi0054 & new_n11273_;
  assign new_n11294_ = ~pi0074 & new_n11293_;
  assign new_n11295_ = pi0055 & ~new_n11294_;
  assign new_n11296_ = pi0045 & new_n2468_;
  assign new_n11297_ = new_n2476_ & new_n11296_;
  assign new_n11298_ = new_n11061_ & new_n11297_;
  assign new_n11299_ = new_n2465_ & new_n11298_;
  assign new_n11300_ = new_n6379_ & new_n9313_;
  assign new_n11301_ = new_n2454_ & new_n3273_;
  assign new_n11302_ = new_n11300_ & new_n11301_;
  assign new_n11303_ = new_n11299_ & new_n11302_;
  assign new_n11304_ = ~pi0055 & ~new_n11303_;
  assign new_n11305_ = new_n8878_ & ~new_n11304_;
  assign po0213 = ~new_n11295_ & new_n11305_;
  assign new_n11307_ = pi0056 & ~pi0062;
  assign new_n11308_ = pi0055 & new_n10142_;
  assign new_n11309_ = ~new_n11307_ & ~new_n11308_;
  assign new_n11310_ = new_n3097_ & new_n3285_;
  assign new_n11311_ = new_n6169_ & new_n11310_;
  assign new_n11312_ = pi0056 & ~new_n11311_;
  assign new_n11313_ = new_n3436_ & ~new_n11312_;
  assign po0214 = ~new_n11309_ & new_n11313_;
  assign new_n11315_ = new_n6385_ & new_n11310_;
  assign new_n11316_ = ~pi0056 & pi0062;
  assign new_n11317_ = ~pi0924 & new_n11316_;
  assign new_n11318_ = ~new_n11307_ & ~new_n11317_;
  assign new_n11319_ = new_n11315_ & ~new_n11318_;
  assign new_n11320_ = ~pi0057 & ~new_n11319_;
  assign new_n11321_ = new_n6304_ & new_n11294_;
  assign new_n11322_ = pi0057 & ~new_n11321_;
  assign new_n11323_ = ~pi0059 & ~new_n11322_;
  assign po0215 = ~new_n11320_ & new_n11323_;
  assign new_n11325_ = ~pi0093 & new_n11086_;
  assign new_n11326_ = new_n10165_ & new_n11325_;
  assign po0216 = new_n7459_ & new_n11326_;
  assign new_n11328_ = pi0924 & new_n11316_;
  assign new_n11329_ = new_n11315_ & new_n11328_;
  assign new_n11330_ = ~pi0059 & ~new_n11329_;
  assign new_n11331_ = pi0059 & ~new_n11321_;
  assign new_n11332_ = ~pi0057 & ~new_n11331_;
  assign po0217 = ~new_n11330_ & new_n11332_;
  assign new_n11334_ = pi0039 & ~pi0979;
  assign new_n11335_ = ~new_n6186_ & new_n11334_;
  assign new_n11336_ = new_n6187_ & new_n11335_;
  assign new_n11337_ = new_n6454_ & new_n11336_;
  assign new_n11338_ = ~pi0039 & new_n11261_;
  assign new_n11339_ = new_n11275_ & new_n11338_;
  assign new_n11340_ = new_n2503_ & new_n11339_;
  assign new_n11341_ = ~new_n11337_ & ~new_n11340_;
  assign po0218 = new_n10200_ & ~new_n11341_;
  assign new_n11343_ = pi0841 & new_n11000_;
  assign new_n11344_ = ~pi0024 & new_n11275_;
  assign new_n11345_ = new_n2503_ & new_n11344_;
  assign new_n11346_ = ~new_n11343_ & ~new_n11345_;
  assign po0219 = new_n10166_ & ~new_n11346_;
  assign new_n11348_ = new_n11311_ & new_n11316_;
  assign new_n11349_ = ~pi0057 & ~new_n11348_;
  assign new_n11350_ = pi0057 & ~new_n10143_;
  assign new_n11351_ = ~pi0059 & ~new_n11350_;
  assign po0220 = ~new_n11349_ & new_n11351_;
  assign new_n11353_ = new_n2670_ & new_n8932_;
  assign new_n11354_ = new_n9042_ & new_n11353_;
  assign new_n11355_ = pi0999 & new_n11354_;
  assign new_n11356_ = ~pi0024 & new_n11002_;
  assign new_n11357_ = ~new_n11355_ & ~new_n11356_;
  assign po0221 = new_n10166_ & ~new_n11357_;
  assign new_n11359_ = ~pi0063 & pi0107;
  assign new_n11360_ = new_n2475_ & new_n11359_;
  assign new_n11361_ = ~pi0064 & ~new_n11360_;
  assign new_n11362_ = new_n2454_ & ~new_n11361_;
  assign new_n11363_ = new_n10173_ & new_n11362_;
  assign new_n11364_ = pi0841 & ~new_n11363_;
  assign new_n11365_ = new_n9042_ & new_n11359_;
  assign new_n11366_ = ~pi0841 & ~new_n11365_;
  assign new_n11367_ = new_n11103_ & ~new_n11366_;
  assign po0222 = ~new_n11364_ & new_n11367_;
  assign new_n11369_ = pi0039 & new_n10218_;
  assign new_n11370_ = new_n10200_ & new_n11369_;
  assign new_n11371_ = ~new_n10223_ & new_n11370_;
  assign po0223 = ~new_n10216_ & new_n11371_;
  assign new_n11373_ = ~pi0199 & ~pi0299;
  assign new_n11374_ = pi0314 & new_n2453_;
  assign new_n11375_ = new_n11300_ & new_n11374_;
  assign new_n11376_ = pi0081 & ~pi0102;
  assign new_n11377_ = new_n11375_ & new_n11376_;
  assign new_n11378_ = new_n2478_ & new_n11377_;
  assign new_n11379_ = new_n3273_ & new_n11378_;
  assign new_n11380_ = ~new_n11373_ & new_n11379_;
  assign new_n11381_ = pi0219 & ~new_n11380_;
  assign new_n11382_ = new_n3211_ & new_n3271_;
  assign new_n11383_ = pi0199 & ~pi0299;
  assign new_n11384_ = new_n3226_ & new_n11383_;
  assign new_n11385_ = new_n11382_ & new_n11384_;
  assign new_n11386_ = new_n11378_ & new_n11385_;
  assign new_n11387_ = ~pi0219 & ~new_n11386_;
  assign new_n11388_ = ~po1038 & ~new_n11387_;
  assign po0224 = ~new_n11381_ & new_n11388_;
  assign new_n11390_ = pi0083 & ~pi0103;
  assign new_n11391_ = new_n11104_ & new_n11390_;
  assign new_n11392_ = new_n10165_ & new_n11391_;
  assign new_n11393_ = new_n11375_ & new_n11392_;
  assign po0225 = new_n2473_ & new_n11393_;
  assign new_n11395_ = ~new_n6223_ & new_n6470_;
  assign new_n11396_ = new_n3329_ & new_n5788_;
  assign new_n11397_ = new_n11395_ & new_n11396_;
  assign new_n11398_ = ~new_n6244_ & new_n6470_;
  assign new_n11399_ = new_n3313_ & new_n3489_;
  assign new_n11400_ = new_n11398_ & new_n11399_;
  assign new_n11401_ = ~new_n11397_ & ~new_n11400_;
  assign po0226 = new_n10983_ & ~new_n11401_;
  assign new_n11403_ = pi0069 & new_n11058_;
  assign new_n11404_ = new_n10148_ & new_n11403_;
  assign new_n11405_ = ~pi0071 & ~new_n11404_;
  assign new_n11406_ = ~pi0081 & ~pi0314;
  assign new_n11407_ = new_n2454_ & new_n11406_;
  assign new_n11408_ = new_n6336_ & new_n11407_;
  assign new_n11409_ = ~new_n11405_ & new_n11408_;
  assign new_n11410_ = pi0071 & pi0314;
  assign new_n11411_ = new_n7463_ & new_n11410_;
  assign new_n11412_ = new_n10151_ & new_n11411_;
  assign new_n11413_ = new_n2474_ & new_n11412_;
  assign new_n11414_ = ~new_n11409_ & ~new_n11413_;
  assign po0227 = new_n11103_ & ~new_n11414_;
  assign new_n11416_ = new_n2548_ & new_n2560_;
  assign new_n11417_ = ~pi0096 & new_n11416_;
  assign new_n11418_ = new_n10170_ & new_n11417_;
  assign new_n11419_ = pi0198 & pi0589;
  assign new_n11420_ = new_n3490_ & ~new_n6244_;
  assign new_n11421_ = new_n11419_ & new_n11420_;
  assign new_n11422_ = pi0210 & pi0589;
  assign new_n11423_ = ~pi0221 & new_n5788_;
  assign new_n11424_ = ~pi0216 & new_n11423_;
  assign new_n11425_ = ~new_n6223_ & new_n11424_;
  assign new_n11426_ = new_n11422_ & new_n11425_;
  assign new_n11427_ = ~new_n11421_ & ~new_n11426_;
  assign new_n11428_ = ~pi0593 & new_n6455_;
  assign new_n11429_ = ~new_n6463_ & new_n11428_;
  assign new_n11430_ = ~new_n11427_ & new_n11429_;
  assign new_n11431_ = ~pi0287 & ~new_n11430_;
  assign new_n11432_ = pi0039 & ~new_n11431_;
  assign new_n11433_ = new_n3100_ & new_n11432_;
  assign new_n11434_ = ~new_n11418_ & ~new_n11433_;
  assign po0228 = new_n10200_ & ~new_n11434_;
  assign new_n11436_ = ~pi0050 & new_n8932_;
  assign new_n11437_ = new_n6342_ & new_n11436_;
  assign new_n11438_ = new_n2458_ & new_n2470_;
  assign new_n11439_ = new_n6321_ & new_n11438_;
  assign new_n11440_ = new_n11015_ & new_n11439_;
  assign new_n11441_ = ~pi0064 & new_n8924_;
  assign new_n11442_ = new_n11440_ & new_n11441_;
  assign new_n11443_ = ~pi0081 & ~new_n11442_;
  assign new_n11444_ = ~pi0199 & pi0200;
  assign new_n11445_ = ~pi0299 & new_n11444_;
  assign new_n11446_ = pi0211 & ~pi0219;
  assign new_n11447_ = pi0299 & new_n11446_;
  assign new_n11448_ = ~new_n11445_ & ~new_n11447_;
  assign new_n11449_ = pi0314 & ~new_n11448_;
  assign new_n11450_ = new_n10162_ & new_n11449_;
  assign new_n11451_ = ~new_n11443_ & new_n11450_;
  assign new_n11452_ = new_n11437_ & new_n11451_;
  assign new_n11453_ = new_n11013_ & new_n11448_;
  assign new_n11454_ = new_n11375_ & new_n11453_;
  assign new_n11455_ = new_n11440_ & new_n11454_;
  assign new_n11456_ = ~new_n11452_ & ~new_n11455_;
  assign po0229 = new_n10165_ & ~new_n11456_;
  assign new_n11458_ = pi0024 & new_n2498_;
  assign new_n11459_ = pi0072 & new_n11458_;
  assign new_n11460_ = pi0088 & new_n10147_;
  assign new_n11461_ = new_n6462_ & new_n9170_;
  assign new_n11462_ = new_n11460_ & new_n11461_;
  assign new_n11463_ = new_n2678_ & new_n11462_;
  assign new_n11464_ = ~new_n11459_ & ~new_n11463_;
  assign new_n11465_ = new_n6379_ & ~new_n11464_;
  assign new_n11466_ = ~pi0039 & ~new_n11465_;
  assign new_n11467_ = new_n7547_ & new_n11398_;
  assign new_n11468_ = new_n7550_ & new_n11395_;
  assign new_n11469_ = pi0039 & ~new_n11468_;
  assign new_n11470_ = ~new_n11467_ & new_n11469_;
  assign new_n11471_ = new_n10200_ & ~new_n11470_;
  assign po0230 = ~new_n11466_ & new_n11471_;
  assign new_n11473_ = new_n9058_ & new_n11398_;
  assign new_n11474_ = ~pi0299 & ~new_n11473_;
  assign new_n11475_ = new_n9069_ & new_n11395_;
  assign new_n11476_ = pi0299 & ~new_n11475_;
  assign new_n11477_ = ~new_n11474_ & ~new_n11476_;
  assign new_n11478_ = pi0039 & ~new_n11477_;
  assign new_n11479_ = ~pi0314 & pi1050;
  assign new_n11480_ = new_n9577_ & new_n10162_;
  assign new_n11481_ = new_n11479_ & new_n11480_;
  assign new_n11482_ = ~pi0039 & ~new_n11481_;
  assign new_n11483_ = new_n10200_ & ~new_n11482_;
  assign po0231 = ~new_n11478_ & new_n11483_;
  assign new_n11485_ = pi0074 & new_n11293_;
  assign new_n11486_ = new_n2538_ & new_n7520_;
  assign new_n11487_ = ~pi0096 & ~new_n11486_;
  assign new_n11488_ = ~pi0096 & ~pi1093;
  assign new_n11489_ = new_n7511_ & new_n11488_;
  assign new_n11490_ = new_n3413_ & new_n7455_;
  assign new_n11491_ = ~new_n11489_ & new_n11490_;
  assign new_n11492_ = ~pi0096 & ~new_n6166_;
  assign new_n11493_ = pi0479 & ~new_n11492_;
  assign new_n11494_ = ~po0840 & ~new_n11493_;
  assign new_n11495_ = new_n11491_ & new_n11494_;
  assign new_n11496_ = ~new_n11487_ & new_n11495_;
  assign new_n11497_ = new_n7482_ & new_n11496_;
  assign new_n11498_ = ~new_n11485_ & ~new_n11497_;
  assign po0232 = ~po1038 & ~new_n11498_;
  assign new_n11500_ = pi0096 & ~pi1093;
  assign new_n11501_ = new_n2798_ & ~new_n11487_;
  assign new_n11502_ = ~new_n11500_ & ~new_n11501_;
  assign new_n11503_ = new_n3227_ & ~new_n11502_;
  assign new_n11504_ = new_n7528_ & new_n11503_;
  assign new_n11505_ = ~pi0075 & ~new_n11504_;
  assign new_n11506_ = new_n3246_ & new_n10171_;
  assign new_n11507_ = pi0075 & ~new_n11506_;
  assign new_n11508_ = new_n8881_ & ~new_n11507_;
  assign po0233 = ~new_n11505_ & new_n11508_;
  assign new_n11510_ = new_n3098_ & new_n10402_;
  assign new_n11511_ = pi0252 & new_n2800_;
  assign new_n11512_ = new_n11510_ & ~new_n11511_;
  assign new_n11513_ = ~pi0137 & new_n11512_;
  assign new_n11514_ = ~pi0137 & new_n2733_;
  assign new_n11515_ = ~new_n8899_ & ~new_n10401_;
  assign new_n11516_ = ~pi0094 & ~new_n8935_;
  assign new_n11517_ = new_n10162_ & ~new_n11516_;
  assign new_n11518_ = ~new_n11515_ & new_n11517_;
  assign new_n11519_ = ~new_n2800_ & ~new_n11518_;
  assign new_n11520_ = ~pi0252 & new_n11518_;
  assign new_n11521_ = new_n8930_ & new_n10176_;
  assign new_n11522_ = pi0252 & new_n11521_;
  assign new_n11523_ = new_n2800_ & ~new_n11522_;
  assign new_n11524_ = ~new_n11520_ & new_n11523_;
  assign new_n11525_ = ~new_n11519_ & ~new_n11524_;
  assign new_n11526_ = pi0122 & ~new_n11525_;
  assign new_n11527_ = new_n7511_ & new_n11519_;
  assign new_n11528_ = ~new_n6277_ & ~new_n11510_;
  assign new_n11529_ = ~new_n11524_ & ~new_n11528_;
  assign new_n11530_ = ~new_n11527_ & new_n11529_;
  assign new_n11531_ = ~pi0122 & ~new_n11530_;
  assign new_n11532_ = ~new_n11526_ & ~new_n11531_;
  assign new_n11533_ = ~pi1093 & ~new_n11532_;
  assign new_n11534_ = ~pi0122 & ~new_n11512_;
  assign new_n11535_ = ~new_n11526_ & ~new_n11534_;
  assign new_n11536_ = pi1093 & ~new_n11535_;
  assign new_n11537_ = ~new_n11533_ & ~new_n11536_;
  assign new_n11538_ = new_n2733_ & ~new_n11537_;
  assign new_n11539_ = ~new_n11514_ & ~new_n11538_;
  assign new_n11540_ = ~new_n11513_ & ~new_n11539_;
  assign new_n11541_ = ~pi0122 & new_n11510_;
  assign new_n11542_ = pi1093 & ~new_n11518_;
  assign new_n11543_ = ~new_n8051_ & ~new_n11542_;
  assign new_n11544_ = ~new_n11541_ & ~new_n11543_;
  assign new_n11545_ = ~new_n11533_ & ~new_n11544_;
  assign new_n11546_ = ~new_n2733_ & ~new_n11545_;
  assign new_n11547_ = ~pi0137 & ~new_n2733_;
  assign new_n11548_ = ~new_n11546_ & ~new_n11547_;
  assign new_n11549_ = pi0252 & pi1092;
  assign new_n11550_ = ~pi1093 & new_n11549_;
  assign new_n11551_ = new_n2753_ & new_n11550_;
  assign new_n11552_ = ~pi0137 & ~new_n11551_;
  assign new_n11553_ = new_n11510_ & new_n11552_;
  assign new_n11554_ = ~new_n11548_ & ~new_n11553_;
  assign new_n11555_ = ~new_n11540_ & ~new_n11554_;
  assign new_n11556_ = ~po1057 & ~new_n11555_;
  assign new_n11557_ = ~new_n10108_ & new_n11521_;
  assign new_n11558_ = po1057 & ~new_n11557_;
  assign new_n11559_ = ~pi0137 & po1057;
  assign new_n11560_ = ~new_n11558_ & ~new_n11559_;
  assign new_n11561_ = ~new_n11556_ & new_n11560_;
  assign new_n11562_ = ~pi0210 & ~new_n11561_;
  assign new_n11563_ = ~new_n11538_ & ~new_n11546_;
  assign new_n11564_ = ~po1057 & ~new_n11563_;
  assign new_n11565_ = ~new_n11558_ & ~new_n11564_;
  assign new_n11566_ = pi0210 & ~new_n11565_;
  assign new_n11567_ = ~new_n11562_ & ~new_n11566_;
  assign new_n11568_ = new_n2447_ & new_n10321_;
  assign new_n11569_ = ~new_n11567_ & ~new_n11568_;
  assign new_n11570_ = ~pi0210 & ~new_n11555_;
  assign new_n11571_ = pi0210 & ~new_n11563_;
  assign new_n11572_ = ~new_n11570_ & ~new_n11571_;
  assign new_n11573_ = new_n11568_ & ~new_n11572_;
  assign new_n11574_ = pi0299 & ~new_n11573_;
  assign new_n11575_ = ~new_n11569_ & new_n11574_;
  assign new_n11576_ = ~pi0198 & ~new_n11561_;
  assign new_n11577_ = pi0198 & ~new_n11565_;
  assign new_n11578_ = ~new_n11576_ & ~new_n11577_;
  assign new_n11579_ = new_n3068_ & new_n6185_;
  assign new_n11580_ = ~new_n11578_ & ~new_n11579_;
  assign new_n11581_ = pi0198 & ~new_n11563_;
  assign new_n11582_ = ~pi0198 & ~new_n11555_;
  assign new_n11583_ = ~new_n11581_ & ~new_n11582_;
  assign new_n11584_ = new_n11579_ & ~new_n11583_;
  assign new_n11585_ = ~pi0299 & ~new_n11584_;
  assign new_n11586_ = ~new_n11580_ & new_n11585_;
  assign new_n11587_ = ~new_n11575_ & ~new_n11586_;
  assign new_n11588_ = pi0232 & ~new_n11587_;
  assign new_n11589_ = ~pi0299 & ~new_n11578_;
  assign new_n11590_ = pi0299 & ~new_n11567_;
  assign new_n11591_ = ~pi0232 & ~new_n11590_;
  assign new_n11592_ = ~new_n11589_ & new_n11591_;
  assign new_n11593_ = ~new_n11588_ & ~new_n11592_;
  assign new_n11594_ = new_n7733_ & ~new_n11593_;
  assign new_n11595_ = new_n2800_ & ~new_n11510_;
  assign new_n11596_ = ~new_n11511_ & ~new_n11519_;
  assign new_n11597_ = ~new_n11595_ & new_n11596_;
  assign new_n11598_ = new_n8051_ & ~new_n11597_;
  assign new_n11599_ = ~new_n11526_ & ~new_n11598_;
  assign new_n11600_ = new_n2733_ & ~new_n11599_;
  assign new_n11601_ = ~new_n2733_ & new_n11542_;
  assign new_n11602_ = ~pi1093 & ~new_n11525_;
  assign new_n11603_ = ~new_n11601_ & ~new_n11602_;
  assign new_n11604_ = ~new_n11600_ & new_n11603_;
  assign new_n11605_ = ~po1057 & new_n11604_;
  assign new_n11606_ = po1057 & new_n11521_;
  assign new_n11607_ = ~new_n10104_ & new_n11606_;
  assign new_n11608_ = ~new_n11605_ & ~new_n11607_;
  assign new_n11609_ = pi0210 & ~new_n11608_;
  assign new_n11610_ = ~pi0137 & ~new_n11597_;
  assign new_n11611_ = ~pi1093 & new_n11610_;
  assign new_n11612_ = pi0137 & new_n11602_;
  assign new_n11613_ = ~new_n11542_ & ~new_n11612_;
  assign new_n11614_ = ~new_n11611_ & new_n11613_;
  assign new_n11615_ = ~po1057 & new_n11614_;
  assign new_n11616_ = ~new_n11606_ & ~new_n11615_;
  assign new_n11617_ = new_n8904_ & new_n11559_;
  assign new_n11618_ = ~new_n2733_ & ~new_n11617_;
  assign new_n11619_ = ~new_n11616_ & new_n11618_;
  assign new_n11620_ = pi0137 & ~new_n11599_;
  assign new_n11621_ = ~new_n11610_ & ~new_n11612_;
  assign new_n11622_ = ~new_n11620_ & new_n11621_;
  assign new_n11623_ = ~po1057 & ~new_n11622_;
  assign new_n11624_ = pi0137 & ~new_n8051_;
  assign new_n11625_ = new_n2800_ & ~new_n11624_;
  assign new_n11626_ = new_n11521_ & ~new_n11625_;
  assign new_n11627_ = po1057 & ~new_n11626_;
  assign new_n11628_ = new_n2733_ & ~new_n11627_;
  assign new_n11629_ = ~new_n11623_ & new_n11628_;
  assign new_n11630_ = ~new_n11619_ & ~new_n11629_;
  assign new_n11631_ = ~pi0210 & ~new_n11630_;
  assign new_n11632_ = ~new_n11609_ & ~new_n11631_;
  assign new_n11633_ = ~new_n11568_ & ~new_n11632_;
  assign new_n11634_ = ~new_n2733_ & new_n11614_;
  assign new_n11635_ = new_n2733_ & new_n11622_;
  assign new_n11636_ = ~new_n11634_ & ~new_n11635_;
  assign new_n11637_ = ~pi0210 & new_n11636_;
  assign new_n11638_ = pi0210 & ~new_n11604_;
  assign new_n11639_ = new_n11568_ & ~new_n11638_;
  assign new_n11640_ = ~new_n11637_ & new_n11639_;
  assign new_n11641_ = pi0299 & ~new_n11640_;
  assign new_n11642_ = ~new_n11633_ & new_n11641_;
  assign new_n11643_ = pi0198 & ~new_n11608_;
  assign new_n11644_ = ~pi0198 & ~new_n11630_;
  assign new_n11645_ = ~new_n11643_ & ~new_n11644_;
  assign new_n11646_ = ~new_n11579_ & ~new_n11645_;
  assign new_n11647_ = ~pi0198 & ~new_n11636_;
  assign new_n11648_ = pi0198 & new_n11604_;
  assign new_n11649_ = ~new_n11647_ & ~new_n11648_;
  assign new_n11650_ = new_n11579_ & ~new_n11649_;
  assign new_n11651_ = ~pi0299 & ~new_n11650_;
  assign new_n11652_ = ~new_n11646_ & new_n11651_;
  assign new_n11653_ = ~new_n11642_ & ~new_n11652_;
  assign new_n11654_ = pi0232 & ~new_n11653_;
  assign new_n11655_ = pi0299 & ~new_n11632_;
  assign new_n11656_ = ~pi0299 & ~new_n11645_;
  assign new_n11657_ = ~pi0232 & ~new_n11656_;
  assign new_n11658_ = ~new_n11655_ & new_n11657_;
  assign new_n11659_ = ~new_n7733_ & ~new_n11658_;
  assign new_n11660_ = ~new_n11654_ & new_n11659_;
  assign new_n11661_ = ~new_n11594_ & ~new_n11660_;
  assign po0234 = new_n10165_ & ~new_n11661_;
  assign new_n11663_ = new_n2578_ & new_n2593_;
  assign new_n11664_ = ~pi0086 & ~new_n11663_;
  assign new_n11665_ = new_n6350_ & ~new_n11664_;
  assign new_n11666_ = new_n2491_ & new_n11665_;
  assign new_n11667_ = ~pi0314 & ~new_n11666_;
  assign new_n11668_ = pi0086 & new_n8899_;
  assign new_n11669_ = new_n2587_ & new_n11668_;
  assign new_n11670_ = pi0314 & ~new_n11669_;
  assign new_n11671_ = new_n10166_ & ~new_n11670_;
  assign po0235 = ~new_n11667_ & new_n11671_;
  assign new_n11673_ = pi0119 & pi0232;
  assign po0236 = ~pi0468 & new_n11673_;
  assign new_n11675_ = pi0163 & ~new_n9700_;
  assign new_n11676_ = ~pi0163 & ~new_n9696_;
  assign new_n11677_ = ~new_n9698_ & new_n11676_;
  assign new_n11678_ = ~new_n11675_ & ~new_n11677_;
  assign new_n11679_ = pi0232 & new_n11678_;
  assign new_n11680_ = pi0075 & ~new_n11679_;
  assign new_n11681_ = pi0100 & ~new_n11679_;
  assign new_n11682_ = ~new_n11680_ & ~new_n11681_;
  assign new_n11683_ = pi0147 & new_n7499_;
  assign new_n11684_ = new_n8989_ & new_n11683_;
  assign new_n11685_ = new_n11682_ & ~new_n11684_;
  assign new_n11686_ = ~new_n8989_ & new_n11679_;
  assign new_n11687_ = pi0074 & ~new_n11686_;
  assign new_n11688_ = ~new_n3436_ & ~new_n11687_;
  assign new_n11689_ = new_n11685_ & new_n11688_;
  assign new_n11690_ = pi0299 & ~new_n11678_;
  assign new_n11691_ = ~new_n9729_ & new_n9730_;
  assign new_n11692_ = pi0184 & new_n6185_;
  assign new_n11693_ = ~new_n11691_ & new_n11692_;
  assign new_n11694_ = ~pi0184 & new_n11691_;
  assign new_n11695_ = ~pi0299 & ~new_n11694_;
  assign new_n11696_ = ~new_n11693_ & new_n11695_;
  assign new_n11697_ = pi0232 & ~new_n11696_;
  assign new_n11698_ = ~new_n11690_ & new_n11697_;
  assign new_n11699_ = ~new_n8989_ & new_n11698_;
  assign new_n11700_ = pi0074 & ~new_n11699_;
  assign new_n11701_ = ~pi0055 & ~new_n11700_;
  assign new_n11702_ = ~pi0187 & ~pi0299;
  assign new_n11703_ = ~pi0147 & pi0299;
  assign new_n11704_ = ~new_n11702_ & ~new_n11703_;
  assign new_n11705_ = new_n7499_ & new_n11704_;
  assign new_n11706_ = new_n8989_ & ~new_n11705_;
  assign new_n11707_ = pi0054 & ~new_n11706_;
  assign new_n11708_ = ~new_n11699_ & new_n11707_;
  assign new_n11709_ = ~pi0187 & ~new_n9025_;
  assign new_n11710_ = pi0187 & ~new_n9027_;
  assign new_n11711_ = pi0147 & ~new_n11710_;
  assign new_n11712_ = ~new_n11709_ & new_n11711_;
  assign new_n11713_ = ~pi0147 & pi0187;
  assign new_n11714_ = new_n9032_ & new_n11713_;
  assign new_n11715_ = ~new_n11712_ & ~new_n11714_;
  assign new_n11716_ = pi0038 & ~new_n11715_;
  assign new_n11717_ = ~pi0040 & ~new_n9213_;
  assign new_n11718_ = ~pi0095 & ~new_n11717_;
  assign new_n11719_ = ~pi0040 & ~new_n9230_;
  assign new_n11720_ = pi0166 & new_n11719_;
  assign new_n11721_ = new_n11718_ & ~new_n11720_;
  assign new_n11722_ = new_n6185_ & ~new_n9256_;
  assign new_n11723_ = ~new_n11721_ & new_n11722_;
  assign new_n11724_ = ~pi0153 & ~new_n11723_;
  assign new_n11725_ = ~pi0040 & ~new_n9316_;
  assign new_n11726_ = ~pi0095 & ~new_n11725_;
  assign new_n11727_ = pi0166 & ~new_n11726_;
  assign new_n11728_ = new_n11722_ & new_n11727_;
  assign new_n11729_ = new_n9255_ & new_n10321_;
  assign new_n11730_ = pi0153 & ~new_n11729_;
  assign new_n11731_ = ~new_n11728_ & new_n11730_;
  assign new_n11732_ = pi0160 & ~new_n11731_;
  assign new_n11733_ = ~new_n11724_ & new_n11732_;
  assign new_n11734_ = ~pi0153 & new_n11721_;
  assign new_n11735_ = ~new_n2449_ & ~new_n9256_;
  assign new_n11736_ = new_n9113_ & ~new_n9114_;
  assign new_n11737_ = ~new_n11735_ & ~new_n11736_;
  assign new_n11738_ = ~new_n11480_ & ~new_n11726_;
  assign new_n11739_ = pi0153 & ~new_n11727_;
  assign new_n11740_ = ~new_n11738_ & new_n11739_;
  assign new_n11741_ = ~pi0160 & new_n6185_;
  assign new_n11742_ = ~new_n11740_ & new_n11741_;
  assign new_n11743_ = ~new_n11737_ & new_n11742_;
  assign new_n11744_ = ~new_n11734_ & new_n11743_;
  assign new_n11745_ = pi0163 & ~new_n11744_;
  assign new_n11746_ = ~new_n11733_ & new_n11745_;
  assign new_n11747_ = ~pi0040 & ~new_n9365_;
  assign new_n11748_ = ~pi0095 & ~new_n11747_;
  assign new_n11749_ = ~new_n11737_ & ~new_n11748_;
  assign new_n11750_ = pi0166 & new_n11749_;
  assign new_n11751_ = ~pi0040 & new_n9189_;
  assign new_n11752_ = ~pi0032 & ~new_n11751_;
  assign new_n11753_ = ~new_n9274_ & ~new_n11752_;
  assign new_n11754_ = ~pi0095 & ~new_n11753_;
  assign new_n11755_ = ~new_n11737_ & ~new_n11754_;
  assign new_n11756_ = ~pi0210 & ~new_n11755_;
  assign new_n11757_ = ~new_n9257_ & ~new_n11752_;
  assign new_n11758_ = ~pi0095 & ~new_n11757_;
  assign new_n11759_ = ~new_n11737_ & ~new_n11758_;
  assign new_n11760_ = pi0210 & ~new_n11759_;
  assign new_n11761_ = new_n10321_ & ~new_n11760_;
  assign new_n11762_ = ~new_n11756_ & new_n11761_;
  assign new_n11763_ = ~pi0153 & ~new_n11762_;
  assign new_n11764_ = ~new_n11750_ & new_n11763_;
  assign new_n11765_ = ~new_n9270_ & ~new_n11737_;
  assign new_n11766_ = pi0210 & ~new_n11765_;
  assign new_n11767_ = ~new_n9276_ & ~new_n11737_;
  assign new_n11768_ = ~pi0210 & ~new_n11767_;
  assign new_n11769_ = new_n10321_ & ~new_n11768_;
  assign new_n11770_ = ~new_n11766_ & new_n11769_;
  assign new_n11771_ = ~new_n9304_ & ~new_n11737_;
  assign new_n11772_ = ~pi0210 & ~new_n11771_;
  assign new_n11773_ = pi0166 & new_n6185_;
  assign new_n11774_ = ~pi0095 & ~new_n9298_;
  assign new_n11775_ = ~new_n11737_ & ~new_n11774_;
  assign new_n11776_ = pi0210 & ~new_n11775_;
  assign new_n11777_ = new_n11773_ & ~new_n11776_;
  assign new_n11778_ = ~new_n11772_ & new_n11777_;
  assign new_n11779_ = pi0153 & ~new_n11778_;
  assign new_n11780_ = ~new_n11770_ & new_n11779_;
  assign new_n11781_ = ~pi0160 & ~new_n11780_;
  assign new_n11782_ = ~new_n11764_ & new_n11781_;
  assign new_n11783_ = new_n11747_ & new_n11773_;
  assign new_n11784_ = ~new_n9256_ & ~new_n11758_;
  assign new_n11785_ = pi0210 & ~new_n11784_;
  assign new_n11786_ = ~new_n9256_ & ~new_n11754_;
  assign new_n11787_ = ~pi0210 & ~new_n11786_;
  assign new_n11788_ = new_n10321_ & ~new_n11787_;
  assign new_n11789_ = ~new_n11785_ & new_n11788_;
  assign new_n11790_ = ~pi0153 & ~new_n11789_;
  assign new_n11791_ = ~new_n11783_ & new_n11790_;
  assign new_n11792_ = ~new_n9256_ & ~new_n11774_;
  assign new_n11793_ = pi0210 & ~new_n11792_;
  assign new_n11794_ = ~pi0210 & ~new_n9305_;
  assign new_n11795_ = new_n11773_ & ~new_n11794_;
  assign new_n11796_ = ~new_n11793_ & new_n11795_;
  assign new_n11797_ = ~pi0210 & ~new_n9277_;
  assign new_n11798_ = pi0210 & ~new_n9271_;
  assign new_n11799_ = new_n10321_ & ~new_n11798_;
  assign new_n11800_ = ~new_n11797_ & new_n11799_;
  assign new_n11801_ = pi0153 & ~new_n11800_;
  assign new_n11802_ = ~new_n11796_ & new_n11801_;
  assign new_n11803_ = pi0160 & ~new_n11802_;
  assign new_n11804_ = ~new_n11791_ & new_n11803_;
  assign new_n11805_ = ~pi0163 & ~new_n11804_;
  assign new_n11806_ = ~new_n11782_ & new_n11805_;
  assign new_n11807_ = ~new_n11746_ & ~new_n11806_;
  assign new_n11808_ = ~new_n6185_ & new_n11749_;
  assign new_n11809_ = pi0299 & ~new_n11808_;
  assign new_n11810_ = ~new_n11807_ & new_n11809_;
  assign new_n11811_ = ~pi0040 & ~new_n9244_;
  assign new_n11812_ = ~pi0095 & ~new_n11811_;
  assign new_n11813_ = ~new_n11737_ & ~new_n11812_;
  assign new_n11814_ = ~new_n6185_ & new_n11813_;
  assign new_n11815_ = ~pi0175 & ~pi0299;
  assign new_n11816_ = pi0189 & new_n11719_;
  assign new_n11817_ = new_n11718_ & ~new_n11816_;
  assign new_n11818_ = ~pi0182 & new_n11737_;
  assign new_n11819_ = pi0182 & new_n9256_;
  assign new_n11820_ = new_n6185_ & ~new_n11819_;
  assign new_n11821_ = ~new_n11818_ & new_n11820_;
  assign new_n11822_ = ~new_n11817_ & new_n11821_;
  assign new_n11823_ = pi0184 & ~new_n11822_;
  assign new_n11824_ = pi0189 & new_n6185_;
  assign new_n11825_ = new_n11811_ & new_n11824_;
  assign new_n11826_ = pi0198 & ~new_n11784_;
  assign new_n11827_ = ~pi0198 & ~new_n11786_;
  assign new_n11828_ = new_n10325_ & ~new_n11827_;
  assign new_n11829_ = ~new_n11826_ & new_n11828_;
  assign new_n11830_ = pi0182 & ~pi0184;
  assign new_n11831_ = ~new_n11829_ & new_n11830_;
  assign new_n11832_ = ~new_n11825_ & new_n11831_;
  assign new_n11833_ = ~new_n11823_ & ~new_n11832_;
  assign new_n11834_ = new_n11815_ & ~new_n11833_;
  assign new_n11835_ = pi0198 & ~new_n11792_;
  assign new_n11836_ = ~pi0198 & ~new_n9305_;
  assign new_n11837_ = new_n11824_ & ~new_n11836_;
  assign new_n11838_ = ~new_n11835_ & new_n11837_;
  assign new_n11839_ = new_n9279_ & new_n10325_;
  assign new_n11840_ = pi0182 & ~new_n11839_;
  assign new_n11841_ = ~new_n11838_ & new_n11840_;
  assign new_n11842_ = pi0198 & ~new_n11775_;
  assign new_n11843_ = ~pi0198 & ~new_n11771_;
  assign new_n11844_ = new_n11824_ & ~new_n11843_;
  assign new_n11845_ = ~new_n11842_ & new_n11844_;
  assign new_n11846_ = ~pi0182 & ~new_n11845_;
  assign new_n11847_ = ~new_n11841_ & ~new_n11846_;
  assign new_n11848_ = pi0095 & ~pi0182;
  assign new_n11849_ = ~new_n9279_ & ~new_n11848_;
  assign new_n11850_ = new_n10325_ & ~new_n11737_;
  assign new_n11851_ = ~new_n11849_ & new_n11850_;
  assign new_n11852_ = ~new_n11847_ & ~new_n11851_;
  assign new_n11853_ = ~pi0184 & ~new_n11852_;
  assign new_n11854_ = pi0175 & ~pi0299;
  assign new_n11855_ = ~pi0095 & pi0189;
  assign new_n11856_ = new_n2476_ & ~new_n11855_;
  assign new_n11857_ = new_n11725_ & ~new_n11856_;
  assign new_n11858_ = ~new_n11848_ & ~new_n11857_;
  assign new_n11859_ = new_n11692_ & ~new_n11858_;
  assign new_n11860_ = ~new_n11818_ & new_n11859_;
  assign new_n11861_ = new_n11854_ & ~new_n11860_;
  assign new_n11862_ = ~new_n11853_ & new_n11861_;
  assign new_n11863_ = ~new_n11834_ & ~new_n11862_;
  assign new_n11864_ = ~new_n11814_ & ~new_n11863_;
  assign new_n11865_ = ~new_n10325_ & new_n11813_;
  assign new_n11866_ = ~pi0198 & ~new_n11755_;
  assign new_n11867_ = pi0198 & ~new_n11759_;
  assign new_n11868_ = new_n10325_ & ~new_n11867_;
  assign new_n11869_ = ~new_n11866_ & new_n11868_;
  assign new_n11870_ = ~pi0182 & ~pi0184;
  assign new_n11871_ = new_n11815_ & new_n11870_;
  assign new_n11872_ = ~new_n11869_ & new_n11871_;
  assign new_n11873_ = ~new_n11865_ & new_n11872_;
  assign new_n11874_ = ~new_n11864_ & ~new_n11873_;
  assign new_n11875_ = ~new_n11810_ & new_n11874_;
  assign new_n11876_ = pi0232 & ~new_n11875_;
  assign new_n11877_ = pi0299 & new_n11749_;
  assign new_n11878_ = ~pi0299 & new_n11813_;
  assign new_n11879_ = ~pi0232 & ~new_n11878_;
  assign new_n11880_ = ~new_n11877_ & new_n11879_;
  assign new_n11881_ = ~pi0039 & ~new_n11880_;
  assign new_n11882_ = ~new_n11876_ & new_n11881_;
  assign new_n11883_ = ~new_n9058_ & ~new_n9255_;
  assign new_n11884_ = ~pi0040 & ~new_n9057_;
  assign new_n11885_ = ~pi0189 & ~new_n11884_;
  assign new_n11886_ = new_n2476_ & ~new_n9061_;
  assign new_n11887_ = new_n9242_ & ~new_n11886_;
  assign new_n11888_ = new_n6215_ & new_n9255_;
  assign new_n11889_ = new_n2476_ & ~new_n9055_;
  assign new_n11890_ = ~pi0040 & ~new_n11889_;
  assign new_n11891_ = new_n6221_ & new_n11890_;
  assign new_n11892_ = ~new_n11888_ & ~new_n11891_;
  assign new_n11893_ = ~new_n11887_ & new_n11892_;
  assign new_n11894_ = pi0189 & ~new_n6238_;
  assign new_n11895_ = new_n11893_ & new_n11894_;
  assign new_n11896_ = ~new_n11885_ & ~new_n11895_;
  assign new_n11897_ = pi0179 & ~new_n11896_;
  assign new_n11898_ = new_n6238_ & ~new_n11884_;
  assign new_n11899_ = new_n9072_ & new_n9242_;
  assign new_n11900_ = ~new_n2476_ & new_n9242_;
  assign new_n11901_ = ~new_n11899_ & ~new_n11900_;
  assign new_n11902_ = new_n11892_ & new_n11901_;
  assign new_n11903_ = ~pi0189 & ~new_n11902_;
  assign new_n11904_ = ~new_n6215_ & new_n11890_;
  assign new_n11905_ = ~new_n11888_ & ~new_n11904_;
  assign new_n11906_ = pi0189 & ~new_n11905_;
  assign new_n11907_ = ~pi0179 & ~new_n6238_;
  assign new_n11908_ = ~new_n11906_ & new_n11907_;
  assign new_n11909_ = ~new_n11903_ & new_n11908_;
  assign new_n11910_ = ~new_n11898_ & ~new_n11909_;
  assign new_n11911_ = ~new_n11897_ & new_n11910_;
  assign new_n11912_ = new_n9058_ & ~new_n11911_;
  assign new_n11913_ = ~new_n11883_ & ~new_n11912_;
  assign new_n11914_ = ~pi0299 & ~new_n11913_;
  assign new_n11915_ = ~new_n9069_ & new_n9255_;
  assign new_n11916_ = pi0299 & ~new_n11915_;
  assign new_n11917_ = pi0166 & ~new_n6212_;
  assign new_n11918_ = new_n11893_ & new_n11917_;
  assign new_n11919_ = ~new_n11884_ & ~new_n11917_;
  assign new_n11920_ = new_n9069_ & ~new_n11919_;
  assign new_n11921_ = ~new_n11918_ & new_n11920_;
  assign new_n11922_ = new_n11916_ & ~new_n11921_;
  assign new_n11923_ = ~new_n11914_ & ~new_n11922_;
  assign new_n11924_ = pi0156 & pi0232;
  assign new_n11925_ = ~new_n11923_ & new_n11924_;
  assign new_n11926_ = new_n6212_ & ~new_n11884_;
  assign new_n11927_ = ~new_n6212_ & new_n11905_;
  assign new_n11928_ = ~new_n11926_ & ~new_n11927_;
  assign new_n11929_ = ~pi0166 & ~new_n6212_;
  assign new_n11930_ = ~new_n11928_ & ~new_n11929_;
  assign new_n11931_ = new_n11902_ & new_n11929_;
  assign new_n11932_ = new_n9069_ & ~new_n11931_;
  assign new_n11933_ = ~new_n11930_ & new_n11932_;
  assign new_n11934_ = new_n11916_ & ~new_n11933_;
  assign new_n11935_ = ~new_n11914_ & ~new_n11934_;
  assign new_n11936_ = ~pi0156 & pi0232;
  assign new_n11937_ = ~new_n11935_ & new_n11936_;
  assign new_n11938_ = ~new_n6238_ & new_n11905_;
  assign new_n11939_ = ~new_n11898_ & ~new_n11938_;
  assign new_n11940_ = new_n9058_ & ~new_n11939_;
  assign new_n11941_ = ~pi0299 & ~new_n11883_;
  assign new_n11942_ = ~new_n11940_ & new_n11941_;
  assign new_n11943_ = new_n9071_ & new_n11928_;
  assign new_n11944_ = ~pi0232 & ~new_n11943_;
  assign new_n11945_ = ~new_n11942_ & new_n11944_;
  assign new_n11946_ = pi0039 & ~new_n11945_;
  assign new_n11947_ = ~new_n11937_ & new_n11946_;
  assign new_n11948_ = ~new_n11925_ & new_n11947_;
  assign new_n11949_ = ~pi0038 & ~new_n11948_;
  assign new_n11950_ = ~new_n11882_ & new_n11949_;
  assign new_n11951_ = ~new_n11716_ & ~new_n11950_;
  assign new_n11952_ = new_n3245_ & ~new_n11951_;
  assign new_n11953_ = pi0100 & ~new_n11698_;
  assign new_n11954_ = pi0038 & ~new_n11705_;
  assign new_n11955_ = ~pi0100 & ~new_n11954_;
  assign new_n11956_ = ~pi0038 & ~pi0040;
  assign new_n11957_ = pi0087 & ~new_n2476_;
  assign new_n11958_ = new_n11956_ & new_n11957_;
  assign new_n11959_ = new_n11955_ & ~new_n11958_;
  assign new_n11960_ = pi0087 & new_n11959_;
  assign new_n11961_ = ~new_n11953_ & ~new_n11960_;
  assign new_n11962_ = ~new_n11952_ & new_n11961_;
  assign new_n11963_ = new_n3242_ & ~new_n11962_;
  assign new_n11964_ = pi0075 & ~new_n11698_;
  assign new_n11965_ = pi0039 & ~new_n9255_;
  assign new_n11966_ = new_n9653_ & ~new_n11965_;
  assign new_n11967_ = new_n2476_ & ~new_n9051_;
  assign new_n11968_ = ~pi0040 & ~new_n11967_;
  assign new_n11969_ = ~pi0179 & ~pi0299;
  assign new_n11970_ = ~pi0156 & pi0299;
  assign new_n11971_ = ~new_n11969_ & ~new_n11970_;
  assign new_n11972_ = new_n7499_ & new_n11971_;
  assign new_n11973_ = new_n2476_ & new_n11972_;
  assign new_n11974_ = new_n11968_ & ~new_n11973_;
  assign new_n11975_ = ~pi0039 & ~new_n11974_;
  assign new_n11976_ = new_n11966_ & ~new_n11975_;
  assign new_n11977_ = new_n11959_ & ~new_n11976_;
  assign new_n11978_ = ~new_n11953_ & ~new_n11977_;
  assign new_n11979_ = new_n9467_ & ~new_n11978_;
  assign new_n11980_ = ~new_n11964_ & ~new_n11979_;
  assign new_n11981_ = ~new_n11963_ & new_n11980_;
  assign new_n11982_ = ~pi0054 & ~new_n11981_;
  assign new_n11983_ = ~new_n11708_ & ~new_n11982_;
  assign new_n11984_ = ~pi0074 & ~new_n11983_;
  assign new_n11985_ = new_n11701_ & ~new_n11984_;
  assign new_n11986_ = pi0055 & ~new_n11687_;
  assign new_n11987_ = pi0054 & ~new_n11685_;
  assign new_n11988_ = pi0163 & pi0232;
  assign new_n11989_ = ~new_n6185_ & new_n9051_;
  assign new_n11990_ = new_n9038_ & ~new_n11989_;
  assign new_n11991_ = new_n11988_ & new_n11990_;
  assign new_n11992_ = new_n11968_ & ~new_n11991_;
  assign new_n11993_ = ~pi0039 & ~new_n11992_;
  assign new_n11994_ = new_n11966_ & ~new_n11993_;
  assign new_n11995_ = pi0038 & ~new_n11683_;
  assign new_n11996_ = ~pi0100 & ~new_n11995_;
  assign new_n11997_ = ~new_n11958_ & new_n11996_;
  assign new_n11998_ = ~new_n11994_ & new_n11997_;
  assign new_n11999_ = ~new_n11681_ & ~new_n11998_;
  assign new_n12000_ = new_n3242_ & ~new_n11999_;
  assign new_n12001_ = ~new_n11956_ & new_n11996_;
  assign new_n12002_ = ~new_n11681_ & ~new_n12001_;
  assign new_n12003_ = ~new_n9462_ & new_n12002_;
  assign new_n12004_ = new_n9467_ & ~new_n12003_;
  assign new_n12005_ = ~new_n11680_ & ~new_n12004_;
  assign new_n12006_ = ~new_n12000_ & new_n12005_;
  assign new_n12007_ = ~pi0054 & ~new_n12006_;
  assign new_n12008_ = ~new_n11987_ & ~new_n12007_;
  assign new_n12009_ = ~pi0074 & ~new_n12008_;
  assign new_n12010_ = new_n11986_ & ~new_n12009_;
  assign new_n12011_ = new_n3298_ & ~new_n12010_;
  assign new_n12012_ = ~new_n11985_ & new_n12011_;
  assign new_n12013_ = ~pi0075 & ~new_n12002_;
  assign new_n12014_ = ~new_n11680_ & ~new_n12013_;
  assign new_n12015_ = ~pi0054 & ~new_n12014_;
  assign new_n12016_ = ~new_n11987_ & ~new_n12015_;
  assign new_n12017_ = ~pi0074 & ~new_n12016_;
  assign new_n12018_ = ~new_n11687_ & ~new_n12017_;
  assign new_n12019_ = ~new_n3298_ & ~new_n12018_;
  assign new_n12020_ = new_n3436_ & ~new_n12019_;
  assign new_n12021_ = ~new_n9524_ & new_n12020_;
  assign new_n12022_ = ~new_n12012_ & new_n12021_;
  assign new_n12023_ = ~new_n11689_ & ~new_n12022_;
  assign new_n12024_ = ~pi0079 & new_n12023_;
  assign new_n12025_ = ~pi0032 & pi0095;
  assign new_n12026_ = ~pi0479 & new_n12025_;
  assign new_n12027_ = new_n2552_ & new_n12026_;
  assign new_n12028_ = ~pi0040 & ~new_n12027_;
  assign new_n12029_ = new_n9621_ & new_n12028_;
  assign new_n12030_ = new_n10321_ & ~new_n12029_;
  assign new_n12031_ = new_n9624_ & new_n12028_;
  assign new_n12032_ = new_n11773_ & ~new_n12031_;
  assign new_n12033_ = ~pi0153 & ~new_n12032_;
  assign new_n12034_ = ~new_n12030_ & new_n12033_;
  assign new_n12035_ = ~pi0210 & ~new_n9572_;
  assign new_n12036_ = ~new_n9570_ & new_n12028_;
  assign new_n12037_ = ~new_n12035_ & new_n12036_;
  assign new_n12038_ = new_n10321_ & ~new_n12037_;
  assign new_n12039_ = ~new_n9589_ & new_n12031_;
  assign new_n12040_ = new_n11773_ & ~new_n12039_;
  assign new_n12041_ = pi0153 & ~new_n12040_;
  assign new_n12042_ = ~new_n12038_ & new_n12041_;
  assign new_n12043_ = ~new_n12034_ & ~new_n12042_;
  assign new_n12044_ = pi0040 & ~new_n6185_;
  assign new_n12045_ = pi0163 & ~new_n12044_;
  assign new_n12046_ = ~new_n12043_ & new_n12045_;
  assign new_n12047_ = pi0160 & ~new_n12046_;
  assign new_n12048_ = pi0153 & new_n9570_;
  assign new_n12049_ = new_n9621_ & ~new_n12048_;
  assign new_n12050_ = new_n10321_ & ~new_n12049_;
  assign new_n12051_ = pi0153 & new_n9589_;
  assign new_n12052_ = new_n9624_ & ~new_n12051_;
  assign new_n12053_ = new_n11773_ & ~new_n12052_;
  assign new_n12054_ = ~pi0040 & pi0163;
  assign new_n12055_ = ~new_n12053_ & new_n12054_;
  assign new_n12056_ = ~new_n12050_ & new_n12055_;
  assign new_n12057_ = pi0153 & new_n9580_;
  assign new_n12058_ = new_n9593_ & new_n12057_;
  assign new_n12059_ = new_n9608_ & new_n10321_;
  assign new_n12060_ = ~pi0040 & ~pi0163;
  assign new_n12061_ = ~new_n12059_ & new_n12060_;
  assign new_n12062_ = ~new_n12058_ & new_n12061_;
  assign new_n12063_ = ~pi0160 & ~new_n12062_;
  assign new_n12064_ = ~new_n12056_ & new_n12063_;
  assign new_n12065_ = ~new_n12047_ & ~new_n12064_;
  assign new_n12066_ = new_n6185_ & new_n12027_;
  assign new_n12067_ = new_n12062_ & ~new_n12066_;
  assign new_n12068_ = pi0299 & ~new_n12067_;
  assign new_n12069_ = ~new_n12065_ & new_n12068_;
  assign new_n12070_ = pi0184 & new_n9600_;
  assign new_n12071_ = ~pi0184 & ~new_n9608_;
  assign new_n12072_ = ~pi0189 & ~new_n12071_;
  assign new_n12073_ = ~new_n12070_ & new_n12072_;
  assign new_n12074_ = pi0182 & new_n12027_;
  assign new_n12075_ = pi0184 & pi0189;
  assign new_n12076_ = ~new_n9603_ & new_n12075_;
  assign new_n12077_ = ~new_n12074_ & ~new_n12076_;
  assign new_n12078_ = ~new_n12073_ & new_n12077_;
  assign new_n12079_ = new_n6185_ & ~new_n12078_;
  assign new_n12080_ = ~pi0040 & ~new_n12079_;
  assign new_n12081_ = new_n11815_ & ~new_n12080_;
  assign new_n12082_ = ~pi0189 & ~new_n9579_;
  assign new_n12083_ = pi0189 & ~new_n9593_;
  assign new_n12084_ = new_n3097_ & ~new_n12083_;
  assign new_n12085_ = ~new_n12082_ & new_n12084_;
  assign new_n12086_ = ~new_n12074_ & ~new_n12085_;
  assign new_n12087_ = new_n6185_ & ~new_n12086_;
  assign new_n12088_ = ~pi0184 & ~new_n12087_;
  assign new_n12089_ = ~new_n9574_ & new_n10325_;
  assign new_n12090_ = pi0189 & new_n9591_;
  assign new_n12091_ = ~pi0182 & pi0184;
  assign new_n12092_ = ~new_n12090_ & new_n12091_;
  assign new_n12093_ = ~new_n12089_ & new_n12092_;
  assign new_n12094_ = ~new_n12088_ & ~new_n12093_;
  assign new_n12095_ = ~pi0040 & ~new_n12094_;
  assign new_n12096_ = ~new_n9573_ & new_n12036_;
  assign new_n12097_ = new_n10325_ & ~new_n12096_;
  assign new_n12098_ = new_n9590_ & new_n12028_;
  assign new_n12099_ = new_n11824_ & ~new_n12098_;
  assign new_n12100_ = pi0182 & pi0184;
  assign new_n12101_ = ~new_n12044_ & new_n12100_;
  assign new_n12102_ = ~new_n12099_ & new_n12101_;
  assign new_n12103_ = ~new_n12097_ & new_n12102_;
  assign new_n12104_ = new_n11854_ & ~new_n12103_;
  assign new_n12105_ = ~new_n12095_ & new_n12104_;
  assign new_n12106_ = ~new_n12081_ & ~new_n12105_;
  assign new_n12107_ = ~new_n12069_ & new_n12106_;
  assign new_n12108_ = ~pi0039 & ~new_n12107_;
  assign new_n12109_ = new_n2552_ & new_n9580_;
  assign new_n12110_ = ~pi0189 & new_n9053_;
  assign new_n12111_ = pi0179 & new_n6224_;
  assign new_n12112_ = ~new_n12110_ & ~new_n12111_;
  assign new_n12113_ = ~new_n6238_ & new_n9058_;
  assign new_n12114_ = ~new_n12112_ & new_n12113_;
  assign new_n12115_ = new_n12109_ & new_n12114_;
  assign new_n12116_ = ~pi0040 & ~pi0299;
  assign new_n12117_ = ~new_n12115_ & new_n12116_;
  assign new_n12118_ = ~new_n6212_ & new_n9069_;
  assign new_n12119_ = pi0156 & new_n6224_;
  assign new_n12120_ = ~pi0166 & new_n9053_;
  assign new_n12121_ = ~new_n12119_ & ~new_n12120_;
  assign new_n12122_ = new_n12118_ & ~new_n12121_;
  assign new_n12123_ = new_n12109_ & new_n12122_;
  assign new_n12124_ = ~pi0040 & pi0299;
  assign new_n12125_ = ~new_n12123_ & new_n12124_;
  assign new_n12126_ = pi0039 & ~new_n12125_;
  assign new_n12127_ = ~new_n12117_ & new_n12126_;
  assign new_n12128_ = pi0232 & ~new_n12127_;
  assign new_n12129_ = ~new_n12108_ & new_n12128_;
  assign new_n12130_ = ~pi0040 & ~pi0232;
  assign new_n12131_ = ~pi0038 & ~new_n12130_;
  assign new_n12132_ = ~new_n12129_ & new_n12131_;
  assign new_n12133_ = ~new_n11716_ & ~new_n12132_;
  assign new_n12134_ = new_n3245_ & ~new_n12133_;
  assign new_n12135_ = pi0087 & ~new_n11956_;
  assign new_n12136_ = new_n11955_ & new_n12135_;
  assign new_n12137_ = ~new_n11953_ & ~new_n12136_;
  assign new_n12138_ = ~new_n12134_ & new_n12137_;
  assign new_n12139_ = new_n3242_ & ~new_n12138_;
  assign new_n12140_ = new_n3097_ & new_n3226_;
  assign new_n12141_ = new_n11972_ & new_n12140_;
  assign new_n12142_ = new_n2552_ & new_n12141_;
  assign new_n12143_ = new_n11956_ & ~new_n12142_;
  assign new_n12144_ = new_n11955_ & ~new_n12143_;
  assign new_n12145_ = ~new_n11953_ & ~new_n12144_;
  assign new_n12146_ = new_n9467_ & ~new_n12145_;
  assign new_n12147_ = ~new_n11964_ & ~new_n12146_;
  assign new_n12148_ = ~new_n12139_ & new_n12147_;
  assign new_n12149_ = ~pi0054 & ~new_n12148_;
  assign new_n12150_ = ~new_n11708_ & ~new_n12149_;
  assign new_n12151_ = ~pi0074 & ~new_n12150_;
  assign new_n12152_ = new_n11701_ & ~new_n12151_;
  assign new_n12153_ = ~pi0092 & new_n3226_;
  assign new_n12154_ = new_n11988_ & new_n12153_;
  assign new_n12155_ = new_n12109_ & new_n12154_;
  assign new_n12156_ = new_n11956_ & ~new_n12155_;
  assign new_n12157_ = ~pi0075 & new_n11996_;
  assign new_n12158_ = ~new_n12156_ & new_n12157_;
  assign new_n12159_ = new_n11682_ & ~new_n12158_;
  assign new_n12160_ = ~pi0054 & ~new_n12159_;
  assign new_n12161_ = ~new_n11987_ & ~new_n12160_;
  assign new_n12162_ = ~pi0074 & ~new_n12161_;
  assign new_n12163_ = new_n11986_ & ~new_n12162_;
  assign new_n12164_ = new_n3298_ & ~new_n12163_;
  assign new_n12165_ = ~new_n12152_ & new_n12164_;
  assign new_n12166_ = new_n12020_ & ~new_n12165_;
  assign new_n12167_ = ~new_n11689_ & ~new_n12166_;
  assign new_n12168_ = pi0079 & new_n12167_;
  assign new_n12169_ = ~pi0034 & new_n10058_;
  assign new_n12170_ = ~new_n12168_ & ~new_n12169_;
  assign new_n12171_ = ~new_n12024_ & new_n12170_;
  assign new_n12172_ = ~pi0079 & ~new_n8977_;
  assign new_n12173_ = new_n12023_ & ~new_n12172_;
  assign new_n12174_ = new_n12167_ & new_n12172_;
  assign new_n12175_ = new_n12169_ & ~new_n12174_;
  assign new_n12176_ = ~new_n12173_ & new_n12175_;
  assign po0237 = new_n12171_ | new_n12176_;
  assign new_n12178_ = pi0098 & pi1092;
  assign new_n12179_ = pi1093 & new_n12178_;
  assign new_n12180_ = ~pi0567 & new_n2754_;
  assign new_n12181_ = ~new_n12179_ & ~new_n12180_;
  assign new_n12182_ = ~new_n8598_ & new_n12181_;
  assign new_n12183_ = pi0588 & ~new_n12182_;
  assign new_n12184_ = pi0592 & ~new_n12181_;
  assign new_n12185_ = ~new_n7455_ & new_n12181_;
  assign new_n12186_ = new_n7455_ & ~new_n12180_;
  assign new_n12187_ = pi0075 & new_n12179_;
  assign new_n12188_ = pi1091 & new_n12179_;
  assign new_n12189_ = ~pi0110 & new_n2490_;
  assign new_n12190_ = ~pi0088 & new_n2484_;
  assign new_n12191_ = new_n10391_ & new_n12190_;
  assign new_n12192_ = new_n12189_ & new_n12191_;
  assign new_n12193_ = new_n7465_ & new_n12192_;
  assign new_n12194_ = new_n7472_ & new_n12193_;
  assign new_n12195_ = pi0051 & new_n12194_;
  assign new_n12196_ = pi0090 & pi0093;
  assign new_n12197_ = ~pi0841 & ~new_n2493_;
  assign new_n12198_ = ~new_n12196_ & new_n12197_;
  assign new_n12199_ = new_n2535_ & new_n12198_;
  assign new_n12200_ = new_n12193_ & new_n12199_;
  assign new_n12201_ = ~new_n12195_ & ~new_n12200_;
  assign new_n12202_ = pi0824 & pi0950;
  assign new_n12203_ = new_n7476_ & new_n12202_;
  assign new_n12204_ = ~new_n12201_ & new_n12203_;
  assign new_n12205_ = ~pi0098 & ~new_n12204_;
  assign new_n12206_ = pi1092 & ~new_n12205_;
  assign new_n12207_ = ~new_n12188_ & ~new_n12206_;
  assign new_n12208_ = ~new_n7572_ & ~new_n12188_;
  assign new_n12209_ = new_n3227_ & ~new_n12208_;
  assign new_n12210_ = ~new_n12207_ & new_n12209_;
  assign new_n12211_ = new_n3099_ & new_n12202_;
  assign new_n12212_ = new_n12194_ & new_n12211_;
  assign new_n12213_ = ~pi0098 & ~new_n12212_;
  assign new_n12214_ = pi1092 & ~new_n12213_;
  assign new_n12215_ = ~new_n12188_ & ~new_n12214_;
  assign new_n12216_ = new_n7614_ & ~new_n12208_;
  assign new_n12217_ = ~new_n12215_ & new_n12216_;
  assign new_n12218_ = ~new_n3212_ & new_n12179_;
  assign new_n12219_ = ~new_n12217_ & ~new_n12218_;
  assign new_n12220_ = ~new_n12210_ & new_n12219_;
  assign new_n12221_ = ~pi0075 & ~new_n12220_;
  assign new_n12222_ = ~new_n12187_ & ~new_n12221_;
  assign new_n12223_ = pi0567 & ~new_n12222_;
  assign new_n12224_ = new_n12186_ & ~new_n12223_;
  assign new_n12225_ = ~new_n12185_ & ~new_n12224_;
  assign new_n12226_ = ~pi0592 & new_n12225_;
  assign new_n12227_ = ~new_n12184_ & ~new_n12226_;
  assign new_n12228_ = ~new_n8520_ & new_n12227_;
  assign new_n12229_ = ~pi1196 & ~new_n12181_;
  assign new_n12230_ = new_n8520_ & ~new_n12229_;
  assign new_n12231_ = ~pi0443 & ~new_n12181_;
  assign new_n12232_ = pi0443 & ~new_n12227_;
  assign new_n12233_ = ~new_n12231_ & ~new_n12232_;
  assign new_n12234_ = new_n8608_ & new_n12233_;
  assign new_n12235_ = pi0443 & ~new_n12181_;
  assign new_n12236_ = ~pi0443 & ~new_n12227_;
  assign new_n12237_ = ~new_n12235_ & ~new_n12236_;
  assign new_n12238_ = ~new_n8608_ & new_n12237_;
  assign new_n12239_ = ~new_n12234_ & ~new_n12238_;
  assign new_n12240_ = pi0435 & ~new_n12239_;
  assign new_n12241_ = pi0444 & new_n12233_;
  assign new_n12242_ = ~pi0444 & new_n12237_;
  assign new_n12243_ = ~pi0436 & ~new_n12242_;
  assign new_n12244_ = ~new_n12241_ & new_n12243_;
  assign new_n12245_ = pi0444 & new_n12237_;
  assign new_n12246_ = ~pi0444 & new_n12233_;
  assign new_n12247_ = pi0436 & ~new_n12246_;
  assign new_n12248_ = ~new_n12245_ & new_n12247_;
  assign new_n12249_ = ~new_n12244_ & ~new_n12248_;
  assign new_n12250_ = ~pi0435 & new_n12249_;
  assign new_n12251_ = ~new_n12240_ & ~new_n12250_;
  assign new_n12252_ = pi0429 & new_n12251_;
  assign new_n12253_ = ~pi0435 & ~new_n12239_;
  assign new_n12254_ = pi0435 & new_n12249_;
  assign new_n12255_ = ~new_n12253_ & ~new_n12254_;
  assign new_n12256_ = ~pi0429 & new_n12255_;
  assign new_n12257_ = ~new_n8545_ & ~new_n12256_;
  assign new_n12258_ = ~new_n12252_ & new_n12257_;
  assign new_n12259_ = pi0429 & new_n12255_;
  assign new_n12260_ = ~pi0429 & new_n12251_;
  assign new_n12261_ = new_n8545_ & ~new_n12260_;
  assign new_n12262_ = ~new_n12259_ & new_n12261_;
  assign new_n12263_ = pi1196 & ~new_n12262_;
  assign new_n12264_ = ~new_n12258_ & new_n12263_;
  assign new_n12265_ = new_n12230_ & ~new_n12264_;
  assign new_n12266_ = ~new_n12228_ & ~new_n12265_;
  assign new_n12267_ = ~pi0428 & ~new_n12266_;
  assign new_n12268_ = pi0428 & new_n12227_;
  assign new_n12269_ = ~new_n12267_ & ~new_n12268_;
  assign new_n12270_ = ~pi0427 & ~new_n12269_;
  assign new_n12271_ = pi0428 & ~new_n12266_;
  assign new_n12272_ = ~pi0428 & new_n12227_;
  assign new_n12273_ = ~new_n12271_ & ~new_n12272_;
  assign new_n12274_ = pi0427 & ~new_n12273_;
  assign new_n12275_ = ~new_n12270_ & ~new_n12274_;
  assign new_n12276_ = pi0430 & ~new_n12275_;
  assign new_n12277_ = ~pi0427 & ~new_n12273_;
  assign new_n12278_ = pi0427 & ~new_n12269_;
  assign new_n12279_ = ~new_n12277_ & ~new_n12278_;
  assign new_n12280_ = ~pi0430 & ~new_n12279_;
  assign new_n12281_ = ~new_n12276_ & ~new_n12280_;
  assign new_n12282_ = pi0426 & ~new_n12281_;
  assign new_n12283_ = pi0430 & ~new_n12279_;
  assign new_n12284_ = ~pi0430 & ~new_n12275_;
  assign new_n12285_ = ~new_n12283_ & ~new_n12284_;
  assign new_n12286_ = ~pi0426 & ~new_n12285_;
  assign new_n12287_ = ~new_n12282_ & ~new_n12286_;
  assign new_n12288_ = pi0445 & ~new_n12287_;
  assign new_n12289_ = pi0426 & ~new_n12285_;
  assign new_n12290_ = ~pi0426 & ~new_n12281_;
  assign new_n12291_ = ~new_n12289_ & ~new_n12290_;
  assign new_n12292_ = ~pi0445 & ~new_n12291_;
  assign new_n12293_ = ~new_n12288_ & ~new_n12292_;
  assign new_n12294_ = ~pi0448 & new_n12293_;
  assign new_n12295_ = pi0445 & ~new_n12291_;
  assign new_n12296_ = ~pi0445 & ~new_n12287_;
  assign new_n12297_ = ~new_n12295_ & ~new_n12296_;
  assign new_n12298_ = pi0448 & new_n12297_;
  assign new_n12299_ = ~new_n8466_ & ~new_n12298_;
  assign new_n12300_ = ~new_n12294_ & new_n12299_;
  assign new_n12301_ = ~pi0448 & new_n12297_;
  assign new_n12302_ = pi0448 & new_n12293_;
  assign new_n12303_ = new_n8466_ & ~new_n12302_;
  assign new_n12304_ = ~new_n12301_ & new_n12303_;
  assign new_n12305_ = pi1199 & ~new_n12304_;
  assign new_n12306_ = ~new_n12300_ & new_n12305_;
  assign new_n12307_ = ~pi1199 & new_n12266_;
  assign new_n12308_ = new_n8598_ & ~new_n12307_;
  assign new_n12309_ = ~new_n12306_ & new_n12308_;
  assign new_n12310_ = new_n12183_ & ~new_n12309_;
  assign new_n12311_ = pi0591 & ~new_n12181_;
  assign new_n12312_ = pi0590 & ~new_n12311_;
  assign new_n12313_ = new_n8697_ & new_n12181_;
  assign new_n12314_ = ~new_n8697_ & new_n12227_;
  assign new_n12315_ = ~new_n12313_ & ~new_n12314_;
  assign new_n12316_ = pi1198 & ~new_n12315_;
  assign new_n12317_ = ~pi1198 & ~new_n12229_;
  assign new_n12318_ = new_n7627_ & new_n12181_;
  assign new_n12319_ = ~new_n7627_ & new_n12227_;
  assign new_n12320_ = ~new_n12318_ & ~new_n12319_;
  assign new_n12321_ = pi0355 & ~new_n12320_;
  assign new_n12322_ = pi0455 & ~new_n12181_;
  assign new_n12323_ = ~pi0455 & ~new_n12227_;
  assign new_n12324_ = ~new_n12322_ & ~new_n12323_;
  assign new_n12325_ = ~pi0452 & ~new_n12324_;
  assign new_n12326_ = ~pi0455 & ~new_n12181_;
  assign new_n12327_ = pi0455 & ~new_n12227_;
  assign new_n12328_ = ~new_n12326_ & ~new_n12327_;
  assign new_n12329_ = pi0452 & ~new_n12328_;
  assign new_n12330_ = ~new_n12325_ & ~new_n12329_;
  assign new_n12331_ = ~pi0355 & new_n12330_;
  assign new_n12332_ = ~new_n12321_ & ~new_n12331_;
  assign new_n12333_ = pi0458 & new_n12332_;
  assign new_n12334_ = ~pi0355 & ~new_n12320_;
  assign new_n12335_ = pi0355 & new_n12330_;
  assign new_n12336_ = ~new_n12334_ & ~new_n12335_;
  assign new_n12337_ = ~pi0458 & new_n12336_;
  assign new_n12338_ = new_n7642_ & ~new_n12337_;
  assign new_n12339_ = ~new_n12333_ & new_n12338_;
  assign new_n12340_ = pi0458 & new_n12336_;
  assign new_n12341_ = ~pi0458 & new_n12332_;
  assign new_n12342_ = ~new_n7642_ & ~new_n12341_;
  assign new_n12343_ = ~new_n12340_ & new_n12342_;
  assign new_n12344_ = pi1196 & ~new_n12343_;
  assign new_n12345_ = ~new_n12339_ & new_n12344_;
  assign new_n12346_ = new_n12317_ & ~new_n12345_;
  assign new_n12347_ = ~new_n12316_ & ~new_n12346_;
  assign new_n12348_ = ~new_n7454_ & ~new_n12347_;
  assign new_n12349_ = new_n7454_ & new_n12227_;
  assign new_n12350_ = ~new_n12348_ & ~new_n12349_;
  assign new_n12351_ = ~new_n7429_ & new_n12350_;
  assign new_n12352_ = pi1199 & ~new_n12227_;
  assign new_n12353_ = pi0351 & new_n12352_;
  assign new_n12354_ = ~new_n12351_ & ~new_n12353_;
  assign new_n12355_ = ~pi0461 & ~new_n12354_;
  assign new_n12356_ = ~new_n7703_ & new_n12350_;
  assign new_n12357_ = ~pi0351 & new_n12352_;
  assign new_n12358_ = ~new_n12356_ & ~new_n12357_;
  assign new_n12359_ = pi0461 & ~new_n12358_;
  assign new_n12360_ = ~new_n12355_ & ~new_n12359_;
  assign new_n12361_ = ~pi0357 & ~new_n12360_;
  assign new_n12362_ = ~pi0461 & ~new_n12358_;
  assign new_n12363_ = pi0461 & ~new_n12354_;
  assign new_n12364_ = ~new_n12362_ & ~new_n12363_;
  assign new_n12365_ = pi0357 & ~new_n12364_;
  assign new_n12366_ = ~new_n12361_ & ~new_n12365_;
  assign new_n12367_ = ~pi0356 & ~new_n12366_;
  assign new_n12368_ = ~pi0357 & ~new_n12364_;
  assign new_n12369_ = pi0357 & ~new_n12360_;
  assign new_n12370_ = ~new_n12368_ & ~new_n12369_;
  assign new_n12371_ = pi0356 & ~new_n12370_;
  assign new_n12372_ = ~new_n12367_ & ~new_n12371_;
  assign new_n12373_ = pi0354 & ~new_n12372_;
  assign new_n12374_ = ~pi0356 & ~new_n12370_;
  assign new_n12375_ = pi0356 & ~new_n12366_;
  assign new_n12376_ = ~new_n12374_ & ~new_n12375_;
  assign new_n12377_ = ~pi0354 & ~new_n12376_;
  assign new_n12378_ = new_n7425_ & ~new_n12377_;
  assign new_n12379_ = ~new_n12373_ & new_n12378_;
  assign new_n12380_ = pi0354 & ~new_n12376_;
  assign new_n12381_ = ~pi0354 & ~new_n12372_;
  assign new_n12382_ = ~new_n7425_ & ~new_n12381_;
  assign new_n12383_ = ~new_n12380_ & new_n12382_;
  assign new_n12384_ = ~pi0591 & ~new_n12383_;
  assign new_n12385_ = ~new_n12379_ & new_n12384_;
  assign new_n12386_ = new_n12312_ & ~new_n12385_;
  assign new_n12387_ = ~pi1197 & ~new_n7913_;
  assign new_n12388_ = ~new_n12227_ & ~new_n12387_;
  assign new_n12389_ = new_n8255_ & ~new_n12185_;
  assign new_n12390_ = ~pi0411 & new_n12178_;
  assign new_n12391_ = new_n7935_ & ~new_n12390_;
  assign new_n12392_ = pi0411 & new_n12206_;
  assign new_n12393_ = new_n12391_ & ~new_n12392_;
  assign new_n12394_ = ~new_n7935_ & ~new_n12178_;
  assign new_n12395_ = ~new_n7937_ & ~new_n12394_;
  assign new_n12396_ = ~pi0411 & new_n12206_;
  assign new_n12397_ = ~new_n12395_ & ~new_n12396_;
  assign new_n12398_ = ~new_n12393_ & ~new_n12397_;
  assign new_n12399_ = ~new_n12188_ & ~new_n12398_;
  assign new_n12400_ = new_n12209_ & ~new_n12399_;
  assign new_n12401_ = pi0411 & new_n12214_;
  assign new_n12402_ = new_n12391_ & ~new_n12401_;
  assign new_n12403_ = ~pi0411 & new_n12214_;
  assign new_n12404_ = ~new_n12395_ & ~new_n12403_;
  assign new_n12405_ = ~new_n12402_ & ~new_n12404_;
  assign new_n12406_ = ~new_n12188_ & ~new_n12405_;
  assign new_n12407_ = new_n12216_ & ~new_n12406_;
  assign new_n12408_ = ~new_n12218_ & ~new_n12407_;
  assign new_n12409_ = ~new_n12400_ & new_n12408_;
  assign new_n12410_ = ~pi0075 & ~new_n12409_;
  assign new_n12411_ = ~new_n12187_ & ~new_n12410_;
  assign new_n12412_ = pi0567 & ~new_n12411_;
  assign new_n12413_ = new_n12186_ & ~new_n12412_;
  assign new_n12414_ = new_n12389_ & ~new_n12413_;
  assign new_n12415_ = ~new_n12184_ & ~new_n12229_;
  assign new_n12416_ = ~pi1199 & new_n12415_;
  assign new_n12417_ = ~new_n12414_ & new_n12416_;
  assign new_n12418_ = new_n7976_ & new_n12217_;
  assign new_n12419_ = new_n7976_ & new_n12206_;
  assign new_n12420_ = ~new_n7976_ & new_n12178_;
  assign new_n12421_ = ~new_n12419_ & ~new_n12420_;
  assign new_n12422_ = new_n12210_ & ~new_n12421_;
  assign new_n12423_ = ~new_n12418_ & ~new_n12422_;
  assign new_n12424_ = new_n12409_ & new_n12423_;
  assign new_n12425_ = new_n12389_ & ~new_n12424_;
  assign new_n12426_ = new_n7976_ & new_n12214_;
  assign new_n12427_ = ~new_n12420_ & ~new_n12426_;
  assign new_n12428_ = new_n12217_ & ~new_n12427_;
  assign new_n12429_ = ~new_n12218_ & ~new_n12428_;
  assign new_n12430_ = ~new_n12422_ & new_n12429_;
  assign new_n12431_ = new_n8353_ & ~new_n12185_;
  assign new_n12432_ = ~new_n12430_ & new_n12431_;
  assign new_n12433_ = ~new_n12425_ & ~new_n12432_;
  assign new_n12434_ = ~pi0075 & pi0567;
  assign new_n12435_ = ~new_n12433_ & new_n12434_;
  assign new_n12436_ = new_n7946_ & new_n12186_;
  assign new_n12437_ = ~new_n12181_ & ~new_n12436_;
  assign new_n12438_ = pi1199 & ~new_n12437_;
  assign new_n12439_ = ~new_n12435_ & new_n12438_;
  assign new_n12440_ = ~new_n7913_ & ~new_n12439_;
  assign new_n12441_ = ~new_n12417_ & new_n12440_;
  assign new_n12442_ = ~pi1197 & new_n12441_;
  assign new_n12443_ = ~new_n12388_ & ~new_n12442_;
  assign new_n12444_ = ~pi0333 & ~new_n12443_;
  assign new_n12445_ = new_n7913_ & ~new_n12227_;
  assign new_n12446_ = ~new_n12441_ & ~new_n12445_;
  assign new_n12447_ = pi0333 & ~new_n12446_;
  assign new_n12448_ = ~new_n12444_ & ~new_n12447_;
  assign new_n12449_ = ~pi0391 & ~new_n12448_;
  assign new_n12450_ = pi0333 & ~new_n12443_;
  assign new_n12451_ = ~pi0333 & ~new_n12446_;
  assign new_n12452_ = ~new_n12450_ & ~new_n12451_;
  assign new_n12453_ = pi0391 & ~new_n12452_;
  assign new_n12454_ = ~new_n12449_ & ~new_n12453_;
  assign new_n12455_ = ~pi0392 & ~new_n12454_;
  assign new_n12456_ = ~pi0391 & ~new_n12452_;
  assign new_n12457_ = pi0391 & ~new_n12448_;
  assign new_n12458_ = ~new_n12456_ & ~new_n12457_;
  assign new_n12459_ = pi0392 & ~new_n12458_;
  assign new_n12460_ = ~new_n12455_ & ~new_n12459_;
  assign new_n12461_ = pi0393 & ~new_n12460_;
  assign new_n12462_ = ~pi0392 & ~new_n12458_;
  assign new_n12463_ = pi0392 & ~new_n12454_;
  assign new_n12464_ = ~new_n12462_ & ~new_n12463_;
  assign new_n12465_ = ~pi0393 & ~new_n12464_;
  assign new_n12466_ = new_n8251_ & ~new_n12465_;
  assign new_n12467_ = ~new_n12461_ & new_n12466_;
  assign new_n12468_ = pi0393 & ~new_n12464_;
  assign new_n12469_ = ~pi0393 & ~new_n12460_;
  assign new_n12470_ = ~new_n8251_ & ~new_n12469_;
  assign new_n12471_ = ~new_n12468_ & new_n12470_;
  assign new_n12472_ = pi0591 & ~new_n12471_;
  assign new_n12473_ = ~new_n12467_ & new_n12472_;
  assign new_n12474_ = ~pi0592 & ~new_n12181_;
  assign new_n12475_ = pi0592 & new_n12225_;
  assign new_n12476_ = ~new_n12474_ & ~new_n12475_;
  assign new_n12477_ = ~new_n8739_ & new_n12476_;
  assign new_n12478_ = new_n8739_ & new_n12181_;
  assign new_n12479_ = pi1199 & ~new_n12478_;
  assign new_n12480_ = ~new_n12477_ & new_n12479_;
  assign new_n12481_ = ~pi1197 & ~new_n12181_;
  assign new_n12482_ = ~new_n7758_ & ~new_n12481_;
  assign new_n12483_ = new_n7761_ & new_n7776_;
  assign new_n12484_ = ~new_n7761_ & ~new_n7776_;
  assign new_n12485_ = ~new_n12483_ & ~new_n12484_;
  assign new_n12486_ = pi0367 & ~new_n12485_;
  assign new_n12487_ = ~pi0367 & new_n12485_;
  assign new_n12488_ = ~new_n12486_ & ~new_n12487_;
  assign new_n12489_ = new_n12476_ & new_n12488_;
  assign new_n12490_ = new_n12181_ & ~new_n12488_;
  assign new_n12491_ = pi1197 & ~new_n12490_;
  assign new_n12492_ = ~new_n12489_ & new_n12491_;
  assign new_n12493_ = new_n12482_ & ~new_n12492_;
  assign new_n12494_ = new_n7758_ & new_n12476_;
  assign new_n12495_ = ~pi1199 & ~new_n12494_;
  assign new_n12496_ = ~new_n12493_ & new_n12495_;
  assign new_n12497_ = ~new_n12480_ & ~new_n12496_;
  assign new_n12498_ = ~pi1198 & ~new_n12497_;
  assign new_n12499_ = pi1198 & ~new_n12476_;
  assign new_n12500_ = ~new_n12498_ & ~new_n12499_;
  assign new_n12501_ = ~pi0374 & ~new_n12500_;
  assign new_n12502_ = pi0374 & ~new_n12497_;
  assign new_n12503_ = ~new_n12501_ & ~new_n12502_;
  assign new_n12504_ = ~pi0369 & ~new_n12503_;
  assign new_n12505_ = pi0371 & new_n8202_;
  assign new_n12506_ = ~pi0371 & ~new_n8202_;
  assign new_n12507_ = ~new_n12505_ & ~new_n12506_;
  assign new_n12508_ = pi0370 & ~new_n12507_;
  assign new_n12509_ = ~pi0370 & new_n12507_;
  assign new_n12510_ = ~new_n12508_ & ~new_n12509_;
  assign new_n12511_ = ~pi0374 & ~new_n12497_;
  assign new_n12512_ = pi0374 & ~new_n12500_;
  assign new_n12513_ = ~new_n12511_ & ~new_n12512_;
  assign new_n12514_ = pi0369 & ~new_n12513_;
  assign new_n12515_ = new_n12510_ & ~new_n12514_;
  assign new_n12516_ = ~new_n12504_ & new_n12515_;
  assign new_n12517_ = pi0369 & ~new_n12503_;
  assign new_n12518_ = ~pi0369 & ~new_n12513_;
  assign new_n12519_ = ~new_n12510_ & ~new_n12518_;
  assign new_n12520_ = ~new_n12517_ & new_n12519_;
  assign new_n12521_ = ~pi0591 & ~new_n12520_;
  assign new_n12522_ = ~new_n12516_ & new_n12521_;
  assign new_n12523_ = ~pi0590 & ~new_n12522_;
  assign new_n12524_ = ~new_n12473_ & new_n12523_;
  assign new_n12525_ = ~pi0588 & ~new_n12524_;
  assign new_n12526_ = ~new_n12386_ & new_n12525_;
  assign new_n12527_ = new_n7733_ & ~new_n12526_;
  assign new_n12528_ = ~new_n12310_ & new_n12527_;
  assign new_n12529_ = ~new_n8057_ & ~new_n12179_;
  assign new_n12530_ = ~pi0122 & new_n12529_;
  assign new_n12531_ = new_n7572_ & ~new_n12530_;
  assign new_n12532_ = new_n3212_ & ~new_n12188_;
  assign new_n12533_ = ~new_n12531_ & new_n12532_;
  assign new_n12534_ = ~pi0087 & new_n12532_;
  assign new_n12535_ = ~new_n12206_ & new_n12534_;
  assign new_n12536_ = pi0087 & new_n12532_;
  assign new_n12537_ = ~new_n12214_ & new_n12536_;
  assign new_n12538_ = ~new_n12535_ & ~new_n12537_;
  assign new_n12539_ = pi0122 & ~new_n12538_;
  assign new_n12540_ = ~new_n12533_ & ~new_n12539_;
  assign new_n12541_ = ~pi0075 & ~new_n12540_;
  assign new_n12542_ = pi0567 & new_n7455_;
  assign new_n12543_ = ~new_n7491_ & new_n12529_;
  assign new_n12544_ = new_n12542_ & ~new_n12543_;
  assign new_n12545_ = ~new_n12541_ & new_n12544_;
  assign new_n12546_ = ~new_n7455_ & ~new_n12529_;
  assign new_n12547_ = ~new_n12180_ & ~new_n12546_;
  assign new_n12548_ = ~new_n12545_ & new_n12547_;
  assign new_n12549_ = ~pi0592 & ~new_n12548_;
  assign new_n12550_ = ~new_n12184_ & ~new_n12549_;
  assign new_n12551_ = ~new_n8520_ & new_n12550_;
  assign new_n12552_ = pi0443 & ~new_n12550_;
  assign new_n12553_ = ~new_n12231_ & ~new_n12552_;
  assign new_n12554_ = new_n8608_ & new_n12553_;
  assign new_n12555_ = ~pi0443 & ~new_n12550_;
  assign new_n12556_ = ~new_n12235_ & ~new_n12555_;
  assign new_n12557_ = ~new_n8608_ & new_n12556_;
  assign new_n12558_ = ~new_n12554_ & ~new_n12557_;
  assign new_n12559_ = pi0435 & ~new_n12558_;
  assign new_n12560_ = pi0444 & new_n12553_;
  assign new_n12561_ = ~pi0444 & new_n12556_;
  assign new_n12562_ = ~pi0436 & ~new_n12561_;
  assign new_n12563_ = ~new_n12560_ & new_n12562_;
  assign new_n12564_ = pi0444 & new_n12556_;
  assign new_n12565_ = ~pi0444 & new_n12553_;
  assign new_n12566_ = pi0436 & ~new_n12565_;
  assign new_n12567_ = ~new_n12564_ & new_n12566_;
  assign new_n12568_ = ~new_n12563_ & ~new_n12567_;
  assign new_n12569_ = ~pi0435 & new_n12568_;
  assign new_n12570_ = ~new_n12559_ & ~new_n12569_;
  assign new_n12571_ = pi0429 & new_n12570_;
  assign new_n12572_ = ~pi0435 & ~new_n12558_;
  assign new_n12573_ = pi0435 & new_n12568_;
  assign new_n12574_ = ~new_n12572_ & ~new_n12573_;
  assign new_n12575_ = ~pi0429 & new_n12574_;
  assign new_n12576_ = ~new_n8545_ & ~new_n12575_;
  assign new_n12577_ = ~new_n12571_ & new_n12576_;
  assign new_n12578_ = pi0429 & new_n12574_;
  assign new_n12579_ = ~pi0429 & new_n12570_;
  assign new_n12580_ = new_n8545_ & ~new_n12579_;
  assign new_n12581_ = ~new_n12578_ & new_n12580_;
  assign new_n12582_ = pi1196 & ~new_n12581_;
  assign new_n12583_ = ~new_n12577_ & new_n12582_;
  assign new_n12584_ = new_n12230_ & ~new_n12583_;
  assign new_n12585_ = ~new_n12551_ & ~new_n12584_;
  assign new_n12586_ = ~pi0428 & ~new_n12585_;
  assign new_n12587_ = pi0428 & new_n12550_;
  assign new_n12588_ = ~new_n12586_ & ~new_n12587_;
  assign new_n12589_ = ~pi0427 & ~new_n12588_;
  assign new_n12590_ = pi0428 & ~new_n12585_;
  assign new_n12591_ = ~pi0428 & new_n12550_;
  assign new_n12592_ = ~new_n12590_ & ~new_n12591_;
  assign new_n12593_ = pi0427 & ~new_n12592_;
  assign new_n12594_ = ~new_n12589_ & ~new_n12593_;
  assign new_n12595_ = pi0430 & ~new_n12594_;
  assign new_n12596_ = ~pi0427 & ~new_n12592_;
  assign new_n12597_ = pi0427 & ~new_n12588_;
  assign new_n12598_ = ~new_n12596_ & ~new_n12597_;
  assign new_n12599_ = ~pi0430 & ~new_n12598_;
  assign new_n12600_ = ~new_n12595_ & ~new_n12599_;
  assign new_n12601_ = pi0426 & ~new_n12600_;
  assign new_n12602_ = pi0430 & ~new_n12598_;
  assign new_n12603_ = ~pi0430 & ~new_n12594_;
  assign new_n12604_ = ~new_n12602_ & ~new_n12603_;
  assign new_n12605_ = ~pi0426 & ~new_n12604_;
  assign new_n12606_ = ~new_n12601_ & ~new_n12605_;
  assign new_n12607_ = pi0445 & ~new_n12606_;
  assign new_n12608_ = pi0426 & ~new_n12604_;
  assign new_n12609_ = ~pi0426 & ~new_n12600_;
  assign new_n12610_ = ~new_n12608_ & ~new_n12609_;
  assign new_n12611_ = ~pi0445 & ~new_n12610_;
  assign new_n12612_ = ~new_n12607_ & ~new_n12611_;
  assign new_n12613_ = pi0448 & new_n12612_;
  assign new_n12614_ = pi0445 & ~new_n12610_;
  assign new_n12615_ = ~pi0445 & ~new_n12606_;
  assign new_n12616_ = ~new_n12614_ & ~new_n12615_;
  assign new_n12617_ = ~pi0448 & new_n12616_;
  assign new_n12618_ = new_n8466_ & ~new_n12617_;
  assign new_n12619_ = ~new_n12613_ & new_n12618_;
  assign new_n12620_ = ~pi0448 & new_n12612_;
  assign new_n12621_ = pi0448 & new_n12616_;
  assign new_n12622_ = ~new_n8466_ & ~new_n12621_;
  assign new_n12623_ = ~new_n12620_ & new_n12622_;
  assign new_n12624_ = pi1199 & ~new_n12623_;
  assign new_n12625_ = ~new_n12619_ & new_n12624_;
  assign new_n12626_ = ~pi1199 & new_n12585_;
  assign new_n12627_ = new_n8598_ & ~new_n12626_;
  assign new_n12628_ = ~new_n12625_ & new_n12627_;
  assign new_n12629_ = new_n12183_ & ~new_n12628_;
  assign new_n12630_ = ~new_n8697_ & new_n12550_;
  assign new_n12631_ = ~new_n12313_ & ~new_n12630_;
  assign new_n12632_ = pi1198 & ~new_n12631_;
  assign new_n12633_ = ~new_n7627_ & new_n12550_;
  assign new_n12634_ = ~new_n12318_ & ~new_n12633_;
  assign new_n12635_ = ~pi0355 & ~new_n12634_;
  assign new_n12636_ = ~pi0455 & ~new_n12550_;
  assign new_n12637_ = ~new_n12322_ & ~new_n12636_;
  assign new_n12638_ = ~pi0452 & ~new_n12637_;
  assign new_n12639_ = pi0455 & ~new_n12550_;
  assign new_n12640_ = ~new_n12326_ & ~new_n12639_;
  assign new_n12641_ = pi0452 & ~new_n12640_;
  assign new_n12642_ = ~new_n12638_ & ~new_n12641_;
  assign new_n12643_ = pi0355 & new_n12642_;
  assign new_n12644_ = ~new_n12635_ & ~new_n12643_;
  assign new_n12645_ = pi0458 & new_n12644_;
  assign new_n12646_ = pi0355 & ~new_n12634_;
  assign new_n12647_ = ~pi0355 & new_n12642_;
  assign new_n12648_ = ~new_n12646_ & ~new_n12647_;
  assign new_n12649_ = ~pi0458 & new_n12648_;
  assign new_n12650_ = ~new_n7642_ & ~new_n12649_;
  assign new_n12651_ = ~new_n12645_ & new_n12650_;
  assign new_n12652_ = pi0458 & new_n12648_;
  assign new_n12653_ = ~pi0458 & new_n12644_;
  assign new_n12654_ = new_n7642_ & ~new_n12653_;
  assign new_n12655_ = ~new_n12652_ & new_n12654_;
  assign new_n12656_ = pi1196 & ~new_n12655_;
  assign new_n12657_ = ~new_n12651_ & new_n12656_;
  assign new_n12658_ = new_n12317_ & ~new_n12657_;
  assign new_n12659_ = ~new_n12632_ & ~new_n12658_;
  assign new_n12660_ = ~new_n7454_ & ~new_n12659_;
  assign new_n12661_ = new_n7454_ & new_n12550_;
  assign new_n12662_ = ~new_n12660_ & ~new_n12661_;
  assign new_n12663_ = ~new_n7429_ & new_n12662_;
  assign new_n12664_ = pi1199 & ~new_n12550_;
  assign new_n12665_ = pi0351 & new_n12664_;
  assign new_n12666_ = ~new_n12663_ & ~new_n12665_;
  assign new_n12667_ = ~pi0461 & ~new_n12666_;
  assign new_n12668_ = ~new_n7703_ & new_n12662_;
  assign new_n12669_ = ~pi0351 & new_n12664_;
  assign new_n12670_ = ~new_n12668_ & ~new_n12669_;
  assign new_n12671_ = pi0461 & ~new_n12670_;
  assign new_n12672_ = ~new_n12667_ & ~new_n12671_;
  assign new_n12673_ = ~pi0357 & ~new_n12672_;
  assign new_n12674_ = ~pi0461 & ~new_n12670_;
  assign new_n12675_ = pi0461 & ~new_n12666_;
  assign new_n12676_ = ~new_n12674_ & ~new_n12675_;
  assign new_n12677_ = pi0357 & ~new_n12676_;
  assign new_n12678_ = ~new_n12673_ & ~new_n12677_;
  assign new_n12679_ = ~pi0356 & ~new_n12678_;
  assign new_n12680_ = ~pi0357 & ~new_n12676_;
  assign new_n12681_ = pi0357 & ~new_n12672_;
  assign new_n12682_ = ~new_n12680_ & ~new_n12681_;
  assign new_n12683_ = pi0356 & ~new_n12682_;
  assign new_n12684_ = ~new_n12679_ & ~new_n12683_;
  assign new_n12685_ = pi0354 & ~new_n12684_;
  assign new_n12686_ = ~pi0356 & ~new_n12682_;
  assign new_n12687_ = pi0356 & ~new_n12678_;
  assign new_n12688_ = ~new_n12686_ & ~new_n12687_;
  assign new_n12689_ = ~pi0354 & ~new_n12688_;
  assign new_n12690_ = new_n7425_ & ~new_n12689_;
  assign new_n12691_ = ~new_n12685_ & new_n12690_;
  assign new_n12692_ = pi0354 & ~new_n12688_;
  assign new_n12693_ = ~pi0354 & ~new_n12684_;
  assign new_n12694_ = ~new_n7425_ & ~new_n12693_;
  assign new_n12695_ = ~new_n12692_ & new_n12694_;
  assign new_n12696_ = ~pi0591 & ~new_n12695_;
  assign new_n12697_ = ~new_n12691_ & new_n12696_;
  assign new_n12698_ = new_n12312_ & ~new_n12697_;
  assign new_n12699_ = pi0367 & ~new_n12181_;
  assign new_n12700_ = pi0592 & ~new_n12548_;
  assign new_n12701_ = ~new_n12474_ & ~new_n12700_;
  assign new_n12702_ = ~pi0367 & ~new_n12701_;
  assign new_n12703_ = ~new_n12699_ & ~new_n12702_;
  assign new_n12704_ = ~new_n7761_ & new_n12703_;
  assign new_n12705_ = ~pi0367 & ~new_n12181_;
  assign new_n12706_ = pi0367 & ~new_n12701_;
  assign new_n12707_ = ~new_n12705_ & ~new_n12706_;
  assign new_n12708_ = new_n7761_ & new_n12707_;
  assign new_n12709_ = ~new_n12704_ & ~new_n12708_;
  assign new_n12710_ = new_n7764_ & new_n12709_;
  assign new_n12711_ = new_n7761_ & ~new_n12703_;
  assign new_n12712_ = ~new_n7761_ & ~new_n12707_;
  assign new_n12713_ = ~new_n12711_ & ~new_n12712_;
  assign new_n12714_ = ~new_n7764_ & ~new_n12713_;
  assign new_n12715_ = new_n7773_ & ~new_n12714_;
  assign new_n12716_ = ~new_n12710_ & new_n12715_;
  assign new_n12717_ = ~new_n7764_ & new_n12709_;
  assign new_n12718_ = new_n7764_ & ~new_n12713_;
  assign new_n12719_ = ~new_n7773_ & ~new_n12718_;
  assign new_n12720_ = ~new_n12717_ & new_n12719_;
  assign new_n12721_ = pi1197 & ~new_n12720_;
  assign new_n12722_ = ~new_n12716_ & new_n12721_;
  assign new_n12723_ = new_n12482_ & ~new_n12722_;
  assign new_n12724_ = new_n7758_ & new_n12701_;
  assign new_n12725_ = ~pi1199 & ~new_n12724_;
  assign new_n12726_ = ~new_n12723_ & new_n12725_;
  assign new_n12727_ = ~pi1198 & new_n12726_;
  assign new_n12728_ = ~new_n8739_ & new_n12701_;
  assign new_n12729_ = ~new_n12478_ & ~new_n12728_;
  assign new_n12730_ = new_n7838_ & new_n12729_;
  assign new_n12731_ = pi1198 & ~new_n12701_;
  assign new_n12732_ = ~new_n12730_ & ~new_n12731_;
  assign new_n12733_ = ~new_n12727_ & new_n12732_;
  assign new_n12734_ = ~pi0374 & ~new_n12733_;
  assign new_n12735_ = pi1199 & new_n12729_;
  assign new_n12736_ = ~new_n12726_ & ~new_n12735_;
  assign new_n12737_ = pi0374 & ~new_n12736_;
  assign new_n12738_ = ~new_n12734_ & ~new_n12737_;
  assign new_n12739_ = pi0369 & ~new_n12738_;
  assign new_n12740_ = ~pi0374 & ~new_n12736_;
  assign new_n12741_ = pi0374 & ~new_n12733_;
  assign new_n12742_ = ~new_n12740_ & ~new_n12741_;
  assign new_n12743_ = ~pi0369 & ~new_n12742_;
  assign new_n12744_ = ~new_n12510_ & ~new_n12743_;
  assign new_n12745_ = ~new_n12739_ & new_n12744_;
  assign new_n12746_ = ~pi0369 & ~new_n12738_;
  assign new_n12747_ = pi0369 & ~new_n12742_;
  assign new_n12748_ = new_n12510_ & ~new_n12747_;
  assign new_n12749_ = ~new_n12746_ & new_n12748_;
  assign new_n12750_ = ~pi0591 & ~new_n12749_;
  assign new_n12751_ = ~new_n12745_ & new_n12750_;
  assign new_n12752_ = ~new_n12387_ & new_n12550_;
  assign new_n12753_ = pi0397 & ~pi0404;
  assign new_n12754_ = ~pi0397 & pi0404;
  assign new_n12755_ = ~new_n12753_ & ~new_n12754_;
  assign new_n12756_ = pi0411 & ~new_n12755_;
  assign new_n12757_ = ~pi0411 & new_n12755_;
  assign new_n12758_ = ~new_n12756_ & ~new_n12757_;
  assign new_n12759_ = ~new_n7917_ & new_n12758_;
  assign new_n12760_ = new_n7917_ & ~new_n12758_;
  assign new_n12761_ = ~new_n12759_ & ~new_n12760_;
  assign new_n12762_ = new_n7511_ & new_n12761_;
  assign new_n12763_ = ~new_n12178_ & ~new_n12762_;
  assign new_n12764_ = ~pi0412 & ~new_n12763_;
  assign new_n12765_ = new_n7511_ & ~new_n12761_;
  assign new_n12766_ = ~new_n12178_ & ~new_n12765_;
  assign new_n12767_ = pi0412 & ~new_n12766_;
  assign new_n12768_ = ~new_n7929_ & ~new_n12767_;
  assign new_n12769_ = ~new_n12764_ & new_n12768_;
  assign new_n12770_ = pi0412 & ~new_n12763_;
  assign new_n12771_ = ~pi0412 & ~new_n12766_;
  assign new_n12772_ = new_n7929_ & ~new_n12771_;
  assign new_n12773_ = ~new_n12770_ & new_n12772_;
  assign new_n12774_ = ~pi0122 & ~new_n12773_;
  assign new_n12775_ = ~new_n12769_ & new_n12774_;
  assign new_n12776_ = ~new_n12178_ & ~new_n12775_;
  assign new_n12777_ = new_n7572_ & ~new_n12776_;
  assign new_n12778_ = ~new_n12188_ & ~new_n12777_;
  assign new_n12779_ = pi0567 & ~new_n12778_;
  assign new_n12780_ = ~new_n12180_ & ~new_n12779_;
  assign new_n12781_ = ~new_n12186_ & ~new_n12780_;
  assign new_n12782_ = pi0122 & new_n12398_;
  assign new_n12783_ = ~new_n12775_ & ~new_n12782_;
  assign new_n12784_ = new_n7572_ & ~new_n12783_;
  assign new_n12785_ = new_n12534_ & ~new_n12784_;
  assign new_n12786_ = pi0122 & new_n12405_;
  assign new_n12787_ = ~new_n12775_ & ~new_n12786_;
  assign new_n12788_ = new_n7572_ & ~new_n12787_;
  assign new_n12789_ = new_n12536_ & ~new_n12788_;
  assign new_n12790_ = ~new_n3212_ & new_n12778_;
  assign new_n12791_ = ~new_n12789_ & ~new_n12790_;
  assign new_n12792_ = ~new_n12785_ & new_n12791_;
  assign new_n12793_ = ~pi0075 & ~new_n12792_;
  assign new_n12794_ = pi0075 & new_n12778_;
  assign new_n12795_ = new_n12542_ & ~new_n12794_;
  assign new_n12796_ = ~new_n12793_ & new_n12795_;
  assign new_n12797_ = ~new_n12781_ & ~new_n12796_;
  assign new_n12798_ = new_n8255_ & ~new_n12797_;
  assign new_n12799_ = ~new_n12229_ & ~new_n12798_;
  assign new_n12800_ = ~pi1199 & ~new_n12799_;
  assign new_n12801_ = ~pi0122 & new_n7511_;
  assign new_n12802_ = ~new_n12178_ & ~new_n12801_;
  assign new_n12803_ = new_n7511_ & new_n7976_;
  assign new_n12804_ = ~pi0122 & ~new_n12178_;
  assign new_n12805_ = ~new_n12803_ & new_n12804_;
  assign new_n12806_ = ~new_n12208_ & ~new_n12805_;
  assign new_n12807_ = ~new_n12802_ & new_n12806_;
  assign new_n12808_ = pi0567 & new_n12807_;
  assign new_n12809_ = ~new_n12180_ & ~new_n12808_;
  assign new_n12810_ = ~new_n12779_ & new_n12809_;
  assign new_n12811_ = ~new_n12186_ & ~new_n12810_;
  assign new_n12812_ = new_n3212_ & ~new_n12806_;
  assign new_n12813_ = ~new_n12777_ & new_n12812_;
  assign new_n12814_ = new_n12421_ & new_n12534_;
  assign new_n12815_ = ~new_n7935_ & ~new_n12396_;
  assign new_n12816_ = ~new_n12393_ & ~new_n12815_;
  assign new_n12817_ = new_n12814_ & ~new_n12816_;
  assign new_n12818_ = ~new_n12426_ & new_n12536_;
  assign new_n12819_ = ~new_n12405_ & new_n12818_;
  assign new_n12820_ = ~new_n12817_ & ~new_n12819_;
  assign new_n12821_ = ~pi0122 & new_n12803_;
  assign new_n12822_ = ~new_n12775_ & ~new_n12821_;
  assign new_n12823_ = ~new_n12820_ & new_n12822_;
  assign new_n12824_ = ~new_n12813_ & ~new_n12823_;
  assign new_n12825_ = ~pi0075 & ~new_n12824_;
  assign new_n12826_ = ~new_n7491_ & ~new_n12807_;
  assign new_n12827_ = ~new_n12777_ & new_n12826_;
  assign new_n12828_ = new_n12542_ & ~new_n12827_;
  assign new_n12829_ = ~new_n12825_ & new_n12828_;
  assign new_n12830_ = ~new_n12811_ & ~new_n12829_;
  assign new_n12831_ = new_n8255_ & ~new_n12830_;
  assign new_n12832_ = ~new_n12186_ & ~new_n12809_;
  assign new_n12833_ = new_n12427_ & new_n12536_;
  assign new_n12834_ = ~new_n12814_ & ~new_n12833_;
  assign new_n12835_ = pi0122 & ~new_n12834_;
  assign new_n12836_ = ~new_n12812_ & ~new_n12835_;
  assign new_n12837_ = ~pi0075 & ~new_n12836_;
  assign new_n12838_ = new_n12542_ & ~new_n12826_;
  assign new_n12839_ = ~new_n12837_ & new_n12838_;
  assign new_n12840_ = ~new_n12832_ & ~new_n12839_;
  assign new_n12841_ = new_n8353_ & ~new_n12840_;
  assign new_n12842_ = ~new_n12831_ & ~new_n12841_;
  assign new_n12843_ = pi1199 & ~new_n12842_;
  assign new_n12844_ = ~new_n12184_ & ~new_n12843_;
  assign new_n12845_ = ~new_n12800_ & new_n12844_;
  assign new_n12846_ = new_n12387_ & new_n12845_;
  assign new_n12847_ = ~new_n12752_ & ~new_n12846_;
  assign new_n12848_ = pi0333 & ~new_n12847_;
  assign new_n12849_ = new_n7913_ & ~new_n12550_;
  assign new_n12850_ = ~new_n7913_ & ~new_n12845_;
  assign new_n12851_ = ~new_n12849_ & ~new_n12850_;
  assign new_n12852_ = ~pi0333 & new_n12851_;
  assign new_n12853_ = ~new_n12848_ & ~new_n12852_;
  assign new_n12854_ = pi0391 & ~new_n12853_;
  assign new_n12855_ = pi0333 & ~new_n12851_;
  assign new_n12856_ = ~pi0333 & new_n12847_;
  assign new_n12857_ = ~new_n12855_ & ~new_n12856_;
  assign new_n12858_ = ~pi0391 & new_n12857_;
  assign new_n12859_ = ~new_n12854_ & ~new_n12858_;
  assign new_n12860_ = ~pi0392 & ~new_n12859_;
  assign new_n12861_ = ~pi0391 & new_n12853_;
  assign new_n12862_ = pi0391 & ~new_n12857_;
  assign new_n12863_ = ~new_n12861_ & ~new_n12862_;
  assign new_n12864_ = pi0392 & new_n12863_;
  assign new_n12865_ = ~new_n12860_ & ~new_n12864_;
  assign new_n12866_ = pi0393 & ~new_n12865_;
  assign new_n12867_ = pi0392 & ~new_n12859_;
  assign new_n12868_ = ~pi0392 & new_n12863_;
  assign new_n12869_ = ~new_n12867_ & ~new_n12868_;
  assign new_n12870_ = ~pi0393 & ~new_n12869_;
  assign new_n12871_ = ~new_n12866_ & ~new_n12870_;
  assign new_n12872_ = new_n8251_ & ~new_n12871_;
  assign new_n12873_ = pi0393 & ~new_n12869_;
  assign new_n12874_ = ~pi0393 & ~new_n12865_;
  assign new_n12875_ = ~new_n12873_ & ~new_n12874_;
  assign new_n12876_ = ~new_n8251_ & ~new_n12875_;
  assign new_n12877_ = pi0591 & ~new_n12876_;
  assign new_n12878_ = ~new_n12872_ & new_n12877_;
  assign new_n12879_ = ~pi0590 & ~new_n12878_;
  assign new_n12880_ = ~new_n12751_ & new_n12879_;
  assign new_n12881_ = ~pi0588 & ~new_n12880_;
  assign new_n12882_ = ~new_n12698_ & new_n12881_;
  assign new_n12883_ = ~new_n7733_ & ~new_n12882_;
  assign new_n12884_ = ~new_n12629_ & new_n12883_;
  assign new_n12885_ = ~pi0080 & ~po1038;
  assign new_n12886_ = ~new_n12884_ & new_n12885_;
  assign new_n12887_ = ~new_n12528_ & new_n12886_;
  assign new_n12888_ = ~new_n8698_ & new_n12181_;
  assign new_n12889_ = ~new_n12387_ & ~new_n12888_;
  assign new_n12890_ = new_n8255_ & ~new_n12780_;
  assign new_n12891_ = new_n12415_ & ~new_n12890_;
  assign new_n12892_ = ~pi1199 & ~new_n12891_;
  assign new_n12893_ = new_n8255_ & ~new_n12810_;
  assign new_n12894_ = new_n8353_ & ~new_n12809_;
  assign new_n12895_ = ~new_n12184_ & ~new_n12894_;
  assign new_n12896_ = ~new_n12893_ & new_n12895_;
  assign new_n12897_ = pi1199 & ~new_n12896_;
  assign new_n12898_ = ~new_n12892_ & ~new_n12897_;
  assign new_n12899_ = new_n12387_ & ~new_n12898_;
  assign new_n12900_ = ~new_n12889_ & ~new_n12899_;
  assign new_n12901_ = pi0333 & ~new_n12900_;
  assign new_n12902_ = new_n7913_ & ~new_n12888_;
  assign new_n12903_ = ~new_n7913_ & ~new_n12898_;
  assign new_n12904_ = ~new_n12902_ & ~new_n12903_;
  assign new_n12905_ = ~pi0333 & ~new_n12904_;
  assign new_n12906_ = ~new_n12901_ & ~new_n12905_;
  assign new_n12907_ = ~pi0391 & ~new_n12906_;
  assign new_n12908_ = pi0392 & new_n8254_;
  assign new_n12909_ = ~pi0392 & ~new_n8254_;
  assign new_n12910_ = ~new_n12908_ & ~new_n12909_;
  assign new_n12911_ = ~pi0333 & ~new_n12900_;
  assign new_n12912_ = pi0333 & ~new_n12904_;
  assign new_n12913_ = ~new_n12911_ & ~new_n12912_;
  assign new_n12914_ = pi0391 & ~new_n12913_;
  assign new_n12915_ = new_n12910_ & ~new_n12914_;
  assign new_n12916_ = ~new_n12907_ & new_n12915_;
  assign new_n12917_ = ~pi0391 & ~new_n12913_;
  assign new_n12918_ = pi0391 & ~new_n12906_;
  assign new_n12919_ = ~new_n12910_ & ~new_n12918_;
  assign new_n12920_ = ~new_n12917_ & new_n12919_;
  assign new_n12921_ = pi0591 & ~new_n12920_;
  assign new_n12922_ = ~new_n12916_ & new_n12921_;
  assign new_n12923_ = ~new_n8698_ & ~new_n8766_;
  assign new_n12924_ = new_n8125_ & ~new_n8743_;
  assign new_n12925_ = ~pi1198 & ~new_n12924_;
  assign new_n12926_ = ~new_n8782_ & ~new_n12925_;
  assign new_n12927_ = ~new_n12923_ & new_n12926_;
  assign new_n12928_ = new_n12181_ & ~new_n12927_;
  assign new_n12929_ = ~pi0591 & ~new_n12928_;
  assign new_n12930_ = ~pi0590 & ~new_n12929_;
  assign new_n12931_ = ~new_n12922_ & new_n12930_;
  assign new_n12932_ = ~new_n8706_ & new_n12181_;
  assign new_n12933_ = new_n8702_ & new_n12932_;
  assign new_n12934_ = ~new_n7429_ & new_n12933_;
  assign new_n12935_ = ~new_n12888_ & ~new_n12934_;
  assign new_n12936_ = pi0461 & ~new_n12935_;
  assign new_n12937_ = ~new_n7703_ & new_n12933_;
  assign new_n12938_ = ~new_n12888_ & ~new_n12937_;
  assign new_n12939_ = ~pi0461 & ~new_n12938_;
  assign new_n12940_ = ~new_n12936_ & ~new_n12939_;
  assign new_n12941_ = pi0357 & ~new_n12940_;
  assign new_n12942_ = pi0461 & ~new_n12938_;
  assign new_n12943_ = ~pi0461 & ~new_n12935_;
  assign new_n12944_ = ~new_n12942_ & ~new_n12943_;
  assign new_n12945_ = ~pi0357 & ~new_n12944_;
  assign new_n12946_ = ~new_n12941_ & ~new_n12945_;
  assign new_n12947_ = pi0356 & ~new_n12946_;
  assign new_n12948_ = pi0357 & ~new_n12944_;
  assign new_n12949_ = ~pi0357 & ~new_n12940_;
  assign new_n12950_ = ~new_n12948_ & ~new_n12949_;
  assign new_n12951_ = ~pi0356 & ~new_n12950_;
  assign new_n12952_ = ~new_n12947_ & ~new_n12951_;
  assign new_n12953_ = ~pi0354 & new_n12952_;
  assign new_n12954_ = pi0356 & ~new_n12950_;
  assign new_n12955_ = ~pi0356 & ~new_n12946_;
  assign new_n12956_ = ~new_n12954_ & ~new_n12955_;
  assign new_n12957_ = pi0354 & new_n12956_;
  assign new_n12958_ = new_n7425_ & ~new_n12957_;
  assign new_n12959_ = ~new_n12953_ & new_n12958_;
  assign new_n12960_ = ~pi0354 & new_n12956_;
  assign new_n12961_ = pi0354 & new_n12952_;
  assign new_n12962_ = ~new_n7425_ & ~new_n12961_;
  assign new_n12963_ = ~new_n12960_ & new_n12962_;
  assign new_n12964_ = ~pi0591 & ~new_n12963_;
  assign new_n12965_ = ~new_n12959_ & new_n12964_;
  assign new_n12966_ = new_n12312_ & ~new_n12965_;
  assign new_n12967_ = ~pi0588 & ~new_n12966_;
  assign new_n12968_ = ~new_n12931_ & new_n12967_;
  assign new_n12969_ = pi0592 & ~new_n8520_;
  assign new_n12970_ = new_n8125_ & ~new_n8829_;
  assign new_n12971_ = ~new_n12969_ & new_n12970_;
  assign new_n12972_ = new_n12181_ & ~new_n12971_;
  assign new_n12973_ = ~pi0428 & ~new_n12972_;
  assign new_n12974_ = pi0428 & ~new_n12888_;
  assign new_n12975_ = ~new_n12973_ & ~new_n12974_;
  assign new_n12976_ = ~pi0427 & ~new_n12975_;
  assign new_n12977_ = pi0428 & ~new_n12972_;
  assign new_n12978_ = ~pi0428 & ~new_n12888_;
  assign new_n12979_ = ~new_n12977_ & ~new_n12978_;
  assign new_n12980_ = pi0427 & ~new_n12979_;
  assign new_n12981_ = ~new_n12976_ & ~new_n12980_;
  assign new_n12982_ = ~pi0430 & ~new_n12981_;
  assign new_n12983_ = ~pi0427 & ~new_n12979_;
  assign new_n12984_ = pi0427 & ~new_n12975_;
  assign new_n12985_ = ~new_n12983_ & ~new_n12984_;
  assign new_n12986_ = pi0430 & ~new_n12985_;
  assign new_n12987_ = ~new_n12982_ & ~new_n12986_;
  assign new_n12988_ = ~pi0426 & ~new_n12987_;
  assign new_n12989_ = ~pi0430 & ~new_n12985_;
  assign new_n12990_ = pi0430 & ~new_n12981_;
  assign new_n12991_ = ~new_n12989_ & ~new_n12990_;
  assign new_n12992_ = pi0426 & ~new_n12991_;
  assign new_n12993_ = ~new_n12988_ & ~new_n12992_;
  assign new_n12994_ = ~pi0445 & ~new_n12993_;
  assign new_n12995_ = ~pi0426 & ~new_n12991_;
  assign new_n12996_ = pi0426 & ~new_n12987_;
  assign new_n12997_ = ~new_n12995_ & ~new_n12996_;
  assign new_n12998_ = pi0445 & ~new_n12997_;
  assign new_n12999_ = ~new_n12994_ & ~new_n12998_;
  assign new_n13000_ = pi0448 & ~new_n12999_;
  assign new_n13001_ = ~pi0445 & ~new_n12997_;
  assign new_n13002_ = pi0445 & ~new_n12993_;
  assign new_n13003_ = ~new_n13001_ & ~new_n13002_;
  assign new_n13004_ = ~pi0448 & ~new_n13003_;
  assign new_n13005_ = ~new_n8466_ & ~new_n13004_;
  assign new_n13006_ = ~new_n13000_ & new_n13005_;
  assign new_n13007_ = ~pi0448 & ~new_n12999_;
  assign new_n13008_ = pi0448 & ~new_n13003_;
  assign new_n13009_ = new_n8466_ & ~new_n13008_;
  assign new_n13010_ = ~new_n13007_ & new_n13009_;
  assign new_n13011_ = pi1199 & ~new_n13010_;
  assign new_n13012_ = ~new_n13006_ & new_n13011_;
  assign new_n13013_ = ~pi1199 & ~new_n12972_;
  assign new_n13014_ = new_n8598_ & ~new_n13013_;
  assign new_n13015_ = ~new_n13012_ & new_n13014_;
  assign new_n13016_ = new_n12183_ & ~new_n13015_;
  assign new_n13017_ = ~new_n7733_ & ~new_n13016_;
  assign new_n13018_ = ~new_n12968_ & new_n13017_;
  assign new_n13019_ = new_n7733_ & new_n12181_;
  assign new_n13020_ = ~pi0080 & po1038;
  assign new_n13021_ = ~new_n13019_ & new_n13020_;
  assign new_n13022_ = ~new_n13018_ & new_n13021_;
  assign new_n13023_ = ~pi0217 & ~new_n13022_;
  assign new_n13024_ = ~new_n12887_ & new_n13023_;
  assign new_n13025_ = ~pi0080 & ~new_n12181_;
  assign new_n13026_ = pi0217 & ~new_n13025_;
  assign new_n13027_ = new_n8870_ & ~new_n13026_;
  assign po0238 = ~new_n13024_ & new_n13027_;
  assign new_n13029_ = ~po1038 & new_n11302_;
  assign new_n13030_ = pi0081 & ~pi0314;
  assign new_n13031_ = new_n2478_ & new_n13030_;
  assign new_n13032_ = pi0068 & ~pi0081;
  assign new_n13033_ = new_n2469_ & new_n13032_;
  assign new_n13034_ = new_n11015_ & new_n13033_;
  assign new_n13035_ = new_n11441_ & new_n13034_;
  assign new_n13036_ = new_n2634_ & new_n13035_;
  assign new_n13037_ = ~new_n13031_ & ~new_n13036_;
  assign po0239 = new_n13029_ & ~new_n13037_;
  assign new_n13039_ = pi0069 & pi0314;
  assign new_n13040_ = new_n2601_ & new_n13039_;
  assign new_n13041_ = pi0066 & ~pi0073;
  assign new_n13042_ = new_n2457_ & new_n13041_;
  assign new_n13043_ = new_n2471_ & new_n13042_;
  assign new_n13044_ = ~new_n13040_ & ~new_n13043_;
  assign new_n13045_ = new_n11103_ & new_n11105_;
  assign po0240 = ~new_n13044_ & new_n13045_;
  assign new_n13047_ = new_n2486_ & new_n11104_;
  assign new_n13048_ = new_n2491_ & new_n13047_;
  assign new_n13049_ = new_n2469_ & new_n2608_;
  assign new_n13050_ = pi0084 & new_n9128_;
  assign new_n13051_ = new_n13049_ & new_n13050_;
  assign new_n13052_ = ~pi0083 & ~new_n13051_;
  assign new_n13053_ = new_n13048_ & ~new_n13052_;
  assign new_n13054_ = new_n2604_ & new_n13053_;
  assign new_n13055_ = ~pi0314 & ~new_n13054_;
  assign new_n13056_ = new_n2456_ & new_n13051_;
  assign new_n13057_ = new_n13048_ & new_n13056_;
  assign new_n13058_ = pi0314 & ~new_n13057_;
  assign new_n13059_ = new_n10166_ & ~new_n13058_;
  assign po0241 = ~new_n13055_ & new_n13059_;
  assign new_n13061_ = pi0211 & pi0299;
  assign new_n13062_ = pi0219 & pi0299;
  assign new_n13063_ = ~new_n13061_ & ~new_n13062_;
  assign new_n13064_ = ~new_n10820_ & new_n13063_;
  assign new_n13065_ = ~po1038 & new_n13064_;
  assign po0242 = new_n11379_ & new_n13065_;
  assign new_n13067_ = new_n6330_ & new_n11106_;
  assign new_n13068_ = ~pi0314 & new_n11107_;
  assign new_n13069_ = new_n11439_ & new_n13068_;
  assign new_n13070_ = ~new_n13067_ & ~new_n13069_;
  assign po0243 = new_n11103_ & ~new_n13070_;
  assign new_n13072_ = new_n7549_ & new_n11396_;
  assign new_n13073_ = new_n7545_ & new_n11399_;
  assign new_n13074_ = ~new_n13072_ & ~new_n13073_;
  assign po0244 = new_n10983_ & ~new_n13074_;
  assign new_n13076_ = new_n2654_ & new_n13047_;
  assign new_n13077_ = pi0314 & new_n10166_;
  assign new_n13078_ = new_n2491_ & new_n13077_;
  assign po0245 = new_n13076_ & new_n13078_;
  assign new_n13080_ = new_n7511_ & new_n11031_;
  assign new_n13081_ = ~pi1093 & ~new_n13080_;
  assign new_n13082_ = new_n7464_ & new_n12191_;
  assign new_n13083_ = new_n11028_ & new_n13082_;
  assign new_n13084_ = new_n11043_ & new_n12189_;
  assign new_n13085_ = new_n13083_ & new_n13084_;
  assign new_n13086_ = pi1093 & ~new_n13085_;
  assign new_n13087_ = new_n3273_ & ~new_n10068_;
  assign new_n13088_ = ~new_n13086_ & new_n13087_;
  assign new_n13089_ = ~new_n13081_ & new_n13088_;
  assign new_n13090_ = new_n7733_ & ~new_n13089_;
  assign new_n13091_ = new_n2497_ & new_n7511_;
  assign new_n13092_ = ~pi1093 & new_n3098_;
  assign new_n13093_ = new_n3273_ & new_n13092_;
  assign new_n13094_ = new_n13091_ & new_n13093_;
  assign new_n13095_ = new_n11460_ & new_n13094_;
  assign new_n13096_ = new_n2678_ & new_n13095_;
  assign new_n13097_ = ~new_n7733_ & ~new_n13096_;
  assign new_n13098_ = ~po1038 & ~new_n13097_;
  assign po0246 = ~new_n13090_ & new_n13098_;
  assign new_n13100_ = pi0070 & ~new_n8959_;
  assign new_n13101_ = new_n2454_ & new_n8917_;
  assign new_n13102_ = new_n8932_ & new_n13101_;
  assign new_n13103_ = new_n10188_ & new_n13102_;
  assign new_n13104_ = pi0841 & new_n7471_;
  assign new_n13105_ = new_n13103_ & new_n13104_;
  assign new_n13106_ = ~pi0070 & ~new_n13105_;
  assign new_n13107_ = new_n3099_ & new_n10165_;
  assign new_n13108_ = ~new_n13106_ & new_n13107_;
  assign po0247 = ~new_n13100_ & new_n13108_;
  assign new_n13110_ = ~pi1050 & new_n9577_;
  assign new_n13111_ = ~pi0090 & ~new_n13110_;
  assign new_n13112_ = new_n11326_ & ~new_n13111_;
  assign new_n13113_ = ~new_n2705_ & new_n13112_;
  assign po0248 = ~new_n7459_ & new_n13113_;
  assign new_n13115_ = ~pi0058 & new_n2565_;
  assign new_n13116_ = ~new_n10158_ & ~new_n13115_;
  assign new_n13117_ = new_n2795_ & new_n10162_;
  assign new_n13118_ = ~new_n13116_ & new_n13117_;
  assign new_n13119_ = pi0024 & new_n2536_;
  assign new_n13120_ = ~new_n2795_ & new_n13119_;
  assign new_n13121_ = new_n11086_ & new_n13120_;
  assign new_n13122_ = new_n2565_ & new_n13121_;
  assign new_n13123_ = ~pi0039 & ~new_n13122_;
  assign new_n13124_ = ~new_n13118_ & new_n13123_;
  assign new_n13125_ = new_n10197_ & ~new_n13124_;
  assign po0249 = new_n7554_ & new_n13125_;
  assign new_n13127_ = pi0092 & new_n3100_;
  assign new_n13128_ = new_n3413_ & new_n11479_;
  assign new_n13129_ = new_n13127_ & new_n13128_;
  assign new_n13130_ = new_n5788_ & new_n6225_;
  assign new_n13131_ = new_n7549_ & new_n13130_;
  assign new_n13132_ = new_n3489_ & new_n6245_;
  assign new_n13133_ = new_n7545_ & new_n13132_;
  assign new_n13134_ = ~new_n13131_ & ~new_n13133_;
  assign new_n13135_ = new_n3282_ & new_n11126_;
  assign new_n13136_ = ~new_n13134_ & new_n13135_;
  assign new_n13137_ = ~new_n13129_ & ~new_n13136_;
  assign po0250 = new_n10163_ & ~new_n13137_;
  assign new_n13139_ = ~pi1050 & new_n3100_;
  assign new_n13140_ = pi0092 & ~new_n13139_;
  assign new_n13141_ = pi0093 & new_n11086_;
  assign new_n13142_ = new_n2734_ & new_n13141_;
  assign new_n13143_ = ~pi0092 & ~new_n13142_;
  assign new_n13144_ = new_n10164_ & ~new_n13143_;
  assign po0251 = ~new_n13140_ & new_n13144_;
  assign new_n13146_ = new_n11069_ & new_n11286_;
  assign new_n13147_ = new_n2733_ & new_n13146_;
  assign new_n13148_ = pi1093 & ~new_n13147_;
  assign new_n13149_ = new_n2800_ & ~new_n13148_;
  assign new_n13150_ = new_n10251_ & new_n11067_;
  assign new_n13151_ = ~new_n2589_ & ~new_n13150_;
  assign new_n13152_ = new_n2514_ & new_n10162_;
  assign new_n13153_ = pi0252 & new_n13152_;
  assign new_n13154_ = ~new_n13151_ & new_n13153_;
  assign new_n13155_ = ~new_n13149_ & ~new_n13154_;
  assign new_n13156_ = ~po0840 & ~new_n13155_;
  assign new_n13157_ = ~new_n13146_ & ~new_n13156_;
  assign new_n13158_ = pi0252 & new_n13155_;
  assign new_n13159_ = ~new_n13157_ & ~new_n13158_;
  assign new_n13160_ = new_n8888_ & ~new_n13159_;
  assign new_n13161_ = ~new_n8888_ & ~new_n13146_;
  assign new_n13162_ = new_n10165_ & ~new_n13161_;
  assign po0252 = ~new_n13160_ & new_n13162_;
  assign new_n13164_ = ~new_n6244_ & ~new_n6466_;
  assign new_n13165_ = new_n3490_ & ~new_n11419_;
  assign new_n13166_ = new_n13164_ & new_n13165_;
  assign new_n13167_ = ~new_n11422_ & new_n11425_;
  assign new_n13168_ = ~new_n6466_ & new_n13167_;
  assign new_n13169_ = pi0039 & ~new_n13168_;
  assign new_n13170_ = ~new_n13166_ & new_n13169_;
  assign new_n13171_ = new_n2450_ & new_n12025_;
  assign new_n13172_ = new_n11458_ & new_n13171_;
  assign new_n13173_ = ~pi0332 & new_n10162_;
  assign new_n13174_ = new_n11285_ & new_n13173_;
  assign new_n13175_ = new_n13103_ & new_n13174_;
  assign new_n13176_ = ~pi0039 & ~new_n13175_;
  assign new_n13177_ = ~new_n13172_ & new_n13176_;
  assign new_n13178_ = new_n10200_ & ~new_n13177_;
  assign po0253 = ~new_n13170_ & new_n13178_;
  assign new_n13180_ = new_n10309_ & new_n13171_;
  assign new_n13181_ = pi0479 & ~po0840;
  assign new_n13182_ = new_n2940_ & new_n13181_;
  assign new_n13183_ = pi0096 & new_n2724_;
  assign new_n13184_ = new_n2534_ & new_n13183_;
  assign new_n13185_ = ~new_n13181_ & new_n13184_;
  assign new_n13186_ = new_n2736_ & new_n13185_;
  assign new_n13187_ = ~new_n13182_ & ~new_n13186_;
  assign new_n13188_ = ~pi0095 & ~new_n13187_;
  assign new_n13189_ = ~new_n13180_ & ~new_n13188_;
  assign po0254 = new_n10165_ & ~new_n13189_;
  assign new_n13191_ = pi0039 & pi0593;
  assign new_n13192_ = ~new_n11427_ & new_n13191_;
  assign new_n13193_ = ~new_n6466_ & new_n13192_;
  assign new_n13194_ = new_n6166_ & new_n13181_;
  assign new_n13195_ = ~po0740 & ~new_n13194_;
  assign new_n13196_ = ~pi0096 & new_n10169_;
  assign new_n13197_ = ~new_n13195_ & new_n13196_;
  assign new_n13198_ = new_n11486_ & new_n13197_;
  assign new_n13199_ = ~new_n13193_ & ~new_n13198_;
  assign po0255 = new_n10200_ & ~new_n13199_;
  assign new_n13201_ = ~pi0092 & new_n11480_;
  assign new_n13202_ = ~new_n13127_ & ~new_n13201_;
  assign new_n13203_ = pi0314 & pi1050;
  assign new_n13204_ = new_n10164_ & new_n13203_;
  assign po0256 = ~new_n13202_ & new_n13204_;
  assign new_n13206_ = ~pi0072 & pi0099;
  assign new_n13207_ = ~new_n8100_ & ~new_n13206_;
  assign new_n13208_ = ~new_n2733_ & new_n13206_;
  assign new_n13209_ = new_n8100_ & ~new_n13208_;
  assign new_n13210_ = ~new_n10314_ & new_n13206_;
  assign new_n13211_ = new_n6266_ & new_n10914_;
  assign new_n13212_ = ~new_n13210_ & ~new_n13211_;
  assign new_n13213_ = new_n10448_ & ~new_n13212_;
  assign new_n13214_ = new_n13209_ & ~new_n13213_;
  assign new_n13215_ = ~new_n13207_ & ~new_n13214_;
  assign new_n13216_ = ~pi0039 & ~new_n13215_;
  assign new_n13217_ = ~pi0072 & pi0152;
  assign new_n13218_ = new_n10322_ & new_n13217_;
  assign new_n13219_ = pi0299 & new_n13218_;
  assign new_n13220_ = ~pi0072 & pi0174;
  assign new_n13221_ = ~pi0299 & new_n13220_;
  assign new_n13222_ = new_n10326_ & new_n13221_;
  assign new_n13223_ = ~new_n13219_ & ~new_n13222_;
  assign new_n13224_ = pi0232 & ~new_n13223_;
  assign new_n13225_ = pi0039 & ~new_n13224_;
  assign new_n13226_ = new_n3246_ & ~new_n13225_;
  assign new_n13227_ = ~new_n13216_ & new_n13226_;
  assign new_n13228_ = ~pi0039 & ~new_n13206_;
  assign new_n13229_ = ~new_n13225_ & ~new_n13228_;
  assign new_n13230_ = ~new_n3246_ & new_n13229_;
  assign new_n13231_ = pi0075 & ~new_n13230_;
  assign new_n13232_ = ~new_n13227_ & new_n13231_;
  assign new_n13233_ = pi0041 & pi0072;
  assign new_n13234_ = pi0099 & ~new_n13233_;
  assign new_n13235_ = ~new_n10375_ & new_n13234_;
  assign new_n13236_ = new_n10745_ & ~new_n13235_;
  assign new_n13237_ = ~new_n10382_ & new_n13234_;
  assign new_n13238_ = new_n10744_ & ~new_n13237_;
  assign new_n13239_ = ~new_n13236_ & ~new_n13238_;
  assign new_n13240_ = pi0228 & ~new_n13239_;
  assign new_n13241_ = ~new_n10429_ & new_n13234_;
  assign new_n13242_ = ~pi0228 & ~new_n10533_;
  assign new_n13243_ = ~new_n13241_ & new_n13242_;
  assign new_n13244_ = ~pi0039 & ~new_n13243_;
  assign new_n13245_ = ~new_n13240_ & new_n13244_;
  assign new_n13246_ = new_n10478_ & ~new_n13223_;
  assign new_n13247_ = ~new_n10944_ & new_n13246_;
  assign new_n13248_ = new_n3211_ & ~new_n13247_;
  assign new_n13249_ = ~new_n13245_ & new_n13248_;
  assign new_n13250_ = ~new_n10445_ & new_n13206_;
  assign new_n13251_ = new_n6265_ & new_n10301_;
  assign new_n13252_ = ~new_n13250_ & ~new_n13251_;
  assign new_n13253_ = new_n10448_ & ~new_n13252_;
  assign new_n13254_ = new_n13209_ & ~new_n13253_;
  assign new_n13255_ = ~new_n13207_ & ~new_n13254_;
  assign new_n13256_ = ~pi0039 & ~new_n13255_;
  assign new_n13257_ = ~new_n13225_ & ~new_n13256_;
  assign new_n13258_ = new_n6258_ & ~new_n13257_;
  assign new_n13259_ = pi0038 & ~new_n13229_;
  assign new_n13260_ = ~pi0087 & ~new_n13259_;
  assign new_n13261_ = ~new_n13258_ & new_n13260_;
  assign new_n13262_ = ~new_n13249_ & new_n13261_;
  assign new_n13263_ = pi0228 & new_n10561_;
  assign new_n13264_ = pi0228 & new_n10442_;
  assign new_n13265_ = new_n13206_ & ~new_n13264_;
  assign new_n13266_ = new_n3281_ & ~new_n13265_;
  assign new_n13267_ = ~new_n13263_ & new_n13266_;
  assign new_n13268_ = ~new_n3281_ & ~new_n13229_;
  assign new_n13269_ = pi0087 & ~new_n13268_;
  assign new_n13270_ = ~new_n13267_ & new_n13269_;
  assign new_n13271_ = ~pi0075 & ~new_n13270_;
  assign new_n13272_ = ~new_n13262_ & new_n13271_;
  assign new_n13273_ = ~new_n13232_ & ~new_n13272_;
  assign new_n13274_ = new_n7455_ & ~new_n13273_;
  assign new_n13275_ = ~new_n7455_ & ~new_n13229_;
  assign new_n13276_ = ~po1038 & ~new_n13275_;
  assign new_n13277_ = ~new_n13274_ & new_n13276_;
  assign new_n13278_ = pi0232 & new_n13218_;
  assign new_n13279_ = pi0039 & ~new_n13278_;
  assign new_n13280_ = po1038 & ~new_n13228_;
  assign new_n13281_ = ~new_n13279_ & new_n13280_;
  assign po0257 = new_n13277_ | new_n13281_;
  assign new_n13283_ = ~new_n7499_ & new_n10072_;
  assign new_n13284_ = pi0129 & ~new_n13283_;
  assign new_n13285_ = new_n7498_ & ~new_n13284_;
  assign new_n13286_ = ~new_n6263_ & ~new_n6281_;
  assign new_n13287_ = pi0129 & ~new_n10072_;
  assign new_n13288_ = ~new_n10075_ & ~new_n13287_;
  assign new_n13289_ = ~new_n13286_ & ~new_n13288_;
  assign new_n13290_ = ~new_n13285_ & new_n13289_;
  assign new_n13291_ = ~pi0075 & new_n3226_;
  assign new_n13292_ = new_n6258_ & new_n13291_;
  assign new_n13293_ = ~new_n13290_ & new_n13292_;
  assign new_n13294_ = ~pi0024 & new_n8967_;
  assign new_n13295_ = po0840 & new_n13294_;
  assign new_n13296_ = ~new_n8964_ & new_n13295_;
  assign new_n13297_ = ~new_n13293_ & ~new_n13296_;
  assign new_n13298_ = new_n8881_ & ~new_n13297_;
  assign po0258 = new_n3100_ & new_n13298_;
  assign new_n13300_ = ~new_n8100_ & ~new_n10307_;
  assign new_n13301_ = ~new_n2733_ & new_n10307_;
  assign new_n13302_ = new_n8100_ & ~new_n13301_;
  assign new_n13303_ = new_n2733_ & ~new_n6273_;
  assign new_n13304_ = new_n10307_ & ~new_n10313_;
  assign new_n13305_ = ~new_n10302_ & ~new_n13304_;
  assign new_n13306_ = new_n13303_ & ~new_n13305_;
  assign new_n13307_ = new_n13302_ & ~new_n13306_;
  assign new_n13308_ = ~new_n13300_ & ~new_n13307_;
  assign new_n13309_ = ~pi0039 & ~new_n13308_;
  assign new_n13310_ = ~pi0144 & pi0174;
  assign new_n13311_ = new_n10325_ & new_n13310_;
  assign new_n13312_ = ~pi0072 & new_n13311_;
  assign new_n13313_ = ~pi0299 & ~new_n13312_;
  assign new_n13314_ = pi0152 & new_n3390_;
  assign new_n13315_ = new_n6185_ & new_n13314_;
  assign new_n13316_ = ~pi0072 & new_n13315_;
  assign new_n13317_ = pi0299 & ~new_n13316_;
  assign new_n13318_ = pi0232 & ~new_n13317_;
  assign new_n13319_ = ~new_n13313_ & new_n13318_;
  assign new_n13320_ = pi0039 & ~new_n13319_;
  assign new_n13321_ = new_n3246_ & ~new_n13320_;
  assign new_n13322_ = ~new_n13309_ & new_n13321_;
  assign new_n13323_ = ~pi0039 & ~new_n10307_;
  assign new_n13324_ = ~new_n13320_ & ~new_n13323_;
  assign new_n13325_ = ~new_n3246_ & new_n13324_;
  assign new_n13326_ = pi0075 & ~new_n13325_;
  assign new_n13327_ = ~new_n13322_ & new_n13326_;
  assign new_n13328_ = pi0101 & new_n10373_;
  assign new_n13329_ = new_n2733_ & ~new_n10360_;
  assign new_n13330_ = ~new_n13328_ & new_n13329_;
  assign new_n13331_ = pi0101 & new_n10380_;
  assign new_n13332_ = ~new_n2733_ & ~new_n10385_;
  assign new_n13333_ = ~new_n13331_ & new_n13332_;
  assign new_n13334_ = ~new_n13330_ & ~new_n13333_;
  assign new_n13335_ = pi0228 & ~new_n13334_;
  assign new_n13336_ = pi0101 & new_n10427_;
  assign new_n13337_ = ~pi0228 & ~new_n10420_;
  assign new_n13338_ = ~new_n13336_ & new_n13337_;
  assign new_n13339_ = ~pi0039 & ~new_n13338_;
  assign new_n13340_ = ~new_n13335_ & new_n13339_;
  assign new_n13341_ = new_n10945_ & new_n13311_;
  assign new_n13342_ = ~pi0299 & ~new_n13341_;
  assign new_n13343_ = new_n10945_ & new_n13315_;
  assign new_n13344_ = pi0299 & ~new_n13343_;
  assign new_n13345_ = new_n10478_ & ~new_n13344_;
  assign new_n13346_ = ~new_n13342_ & new_n13345_;
  assign new_n13347_ = new_n3211_ & ~new_n13346_;
  assign new_n13348_ = ~new_n13340_ & new_n13347_;
  assign new_n13349_ = ~pi0044 & new_n10949_;
  assign new_n13350_ = new_n10307_ & ~new_n13349_;
  assign new_n13351_ = ~new_n10301_ & ~new_n13350_;
  assign new_n13352_ = new_n13303_ & ~new_n13351_;
  assign new_n13353_ = new_n13302_ & ~new_n13352_;
  assign new_n13354_ = ~new_n13300_ & ~new_n13353_;
  assign new_n13355_ = ~pi0039 & ~new_n13354_;
  assign new_n13356_ = ~new_n13320_ & ~new_n13355_;
  assign new_n13357_ = new_n6258_ & ~new_n13356_;
  assign new_n13358_ = pi0038 & ~new_n13324_;
  assign new_n13359_ = ~pi0087 & ~new_n13358_;
  assign new_n13360_ = ~new_n13357_ & new_n13359_;
  assign new_n13361_ = ~new_n13348_ & new_n13360_;
  assign new_n13362_ = ~pi0101 & new_n10962_;
  assign new_n13363_ = new_n10441_ & new_n10961_;
  assign new_n13364_ = new_n10307_ & ~new_n13363_;
  assign new_n13365_ = ~pi0039 & ~new_n13364_;
  assign new_n13366_ = ~new_n13362_ & new_n13365_;
  assign new_n13367_ = pi0087 & ~new_n13320_;
  assign new_n13368_ = ~new_n13366_ & new_n13367_;
  assign new_n13369_ = ~pi0075 & ~new_n13368_;
  assign new_n13370_ = ~new_n13361_ & new_n13369_;
  assign new_n13371_ = ~new_n13327_ & ~new_n13370_;
  assign new_n13372_ = new_n7455_ & ~new_n13371_;
  assign new_n13373_ = ~new_n7455_ & ~new_n13324_;
  assign new_n13374_ = ~po1038 & ~new_n13373_;
  assign new_n13375_ = ~new_n13372_ & new_n13374_;
  assign new_n13376_ = pi0232 & new_n13316_;
  assign new_n13377_ = pi0039 & ~new_n13376_;
  assign new_n13378_ = po1038 & ~new_n13323_;
  assign new_n13379_ = ~new_n13377_ & new_n13378_;
  assign po0259 = new_n13375_ | new_n13379_;
  assign new_n13381_ = new_n2660_ & new_n8918_;
  assign po0260 = new_n13029_ & new_n13381_;
  assign new_n13383_ = ~pi0109 & ~new_n13076_;
  assign new_n13384_ = new_n6320_ & ~new_n13383_;
  assign new_n13385_ = ~pi0314 & ~new_n13384_;
  assign new_n13386_ = pi0109 & new_n2574_;
  assign new_n13387_ = new_n2487_ & new_n13386_;
  assign new_n13388_ = pi0314 & ~new_n13387_;
  assign new_n13389_ = new_n11102_ & ~new_n13388_;
  assign po0261 = ~new_n13385_ & new_n13389_;
  assign new_n13391_ = new_n7733_ & ~new_n8888_;
  assign new_n13392_ = new_n10069_ & ~new_n13391_;
  assign new_n13393_ = new_n10415_ & ~new_n13392_;
  assign new_n13394_ = ~pi0110 & ~new_n13083_;
  assign new_n13395_ = ~pi0047 & new_n11043_;
  assign new_n13396_ = ~new_n13394_ & new_n13395_;
  assign new_n13397_ = new_n10394_ & new_n13396_;
  assign new_n13398_ = ~po1057 & ~new_n13397_;
  assign new_n13399_ = po1057 & ~new_n13085_;
  assign new_n13400_ = ~new_n7500_ & ~new_n10068_;
  assign new_n13401_ = ~new_n13399_ & new_n13400_;
  assign new_n13402_ = ~new_n13398_ & new_n13401_;
  assign new_n13403_ = new_n7500_ & ~new_n10068_;
  assign new_n13404_ = new_n13397_ & new_n13403_;
  assign new_n13405_ = ~new_n13402_ & ~new_n13404_;
  assign new_n13406_ = ~new_n7733_ & ~new_n13405_;
  assign new_n13407_ = ~new_n13393_ & ~new_n13406_;
  assign po0262 = new_n10165_ & ~new_n13407_;
  assign new_n13409_ = pi0024 & new_n11284_;
  assign new_n13410_ = ~pi0053 & ~new_n11283_;
  assign new_n13411_ = new_n2508_ & ~new_n13410_;
  assign new_n13412_ = ~pi0024 & new_n2514_;
  assign new_n13413_ = new_n13411_ & new_n13412_;
  assign new_n13414_ = ~new_n13409_ & ~new_n13413_;
  assign new_n13415_ = pi0841 & ~new_n13414_;
  assign new_n13416_ = new_n8946_ & new_n11264_;
  assign new_n13417_ = ~new_n13415_ & ~new_n13416_;
  assign po0264 = new_n10166_ & ~new_n13417_;
  assign new_n13419_ = ~pi0999 & new_n10166_;
  assign po0265 = new_n11354_ & new_n13419_;
  assign new_n13421_ = ~pi0097 & new_n7468_;
  assign new_n13422_ = ~pi0108 & ~new_n13421_;
  assign new_n13423_ = new_n2490_ & ~new_n13422_;
  assign new_n13424_ = new_n10237_ & new_n13423_;
  assign new_n13425_ = ~pi0314 & ~new_n13424_;
  assign new_n13426_ = pi0314 & ~new_n7470_;
  assign new_n13427_ = new_n7472_ & ~new_n10260_;
  assign new_n13428_ = ~new_n13426_ & new_n13427_;
  assign new_n13429_ = ~new_n13425_ & new_n13428_;
  assign new_n13430_ = new_n7472_ & new_n10260_;
  assign new_n13431_ = new_n13424_ & new_n13430_;
  assign new_n13432_ = ~pi0051 & ~new_n13431_;
  assign new_n13433_ = ~new_n13429_ & new_n13432_;
  assign new_n13434_ = new_n3212_ & new_n7512_;
  assign new_n13435_ = ~new_n13433_ & new_n13434_;
  assign new_n13436_ = ~pi0087 & ~new_n13435_;
  assign new_n13437_ = new_n6289_ & new_n8881_;
  assign po0266 = ~new_n13436_ & new_n13437_;
  assign new_n13439_ = new_n2593_ & new_n11436_;
  assign po0267 = new_n13077_ & new_n13439_;
  assign new_n13441_ = ~pi0082 & ~pi0109;
  assign new_n13442_ = pi0111 & new_n13441_;
  assign new_n13443_ = new_n12189_ & new_n13442_;
  assign new_n13444_ = new_n2486_ & new_n13443_;
  assign new_n13445_ = new_n11107_ & new_n13444_;
  assign new_n13446_ = new_n2635_ & new_n13445_;
  assign new_n13447_ = pi0314 & new_n13446_;
  assign new_n13448_ = new_n8888_ & new_n10069_;
  assign new_n13449_ = new_n10407_ & new_n13448_;
  assign new_n13450_ = ~new_n13447_ & ~new_n13449_;
  assign po0268 = new_n10166_ & ~new_n13450_;
  assign new_n13452_ = pi0072 & new_n10309_;
  assign new_n13453_ = ~pi0314 & new_n13446_;
  assign new_n13454_ = new_n9170_ & new_n13453_;
  assign new_n13455_ = ~new_n13452_ & ~new_n13454_;
  assign new_n13456_ = new_n6379_ & new_n10165_;
  assign po0269 = ~new_n13455_ & new_n13456_;
  assign po0270 = ~pi0124 | pi0468;
  assign new_n13459_ = ~new_n2733_ & ~new_n10382_;
  assign new_n13460_ = ~pi0099 & ~new_n13459_;
  assign new_n13461_ = ~new_n10376_ & new_n13460_;
  assign new_n13462_ = pi0113 & ~new_n10491_;
  assign new_n13463_ = ~new_n13461_ & new_n13462_;
  assign new_n13464_ = ~pi0113 & new_n10746_;
  assign new_n13465_ = pi0228 & ~new_n13464_;
  assign new_n13466_ = ~new_n13463_ & new_n13465_;
  assign new_n13467_ = pi0113 & new_n10527_;
  assign new_n13468_ = ~pi0228 & ~new_n10534_;
  assign new_n13469_ = ~new_n13467_ & new_n13468_;
  assign new_n13470_ = ~pi0039 & ~new_n13469_;
  assign new_n13471_ = ~new_n13466_ & new_n13470_;
  assign new_n13472_ = new_n3211_ & ~new_n13471_;
  assign new_n13473_ = ~pi0072 & pi0113;
  assign new_n13474_ = ~pi0039 & new_n13473_;
  assign new_n13475_ = pi0038 & ~new_n13474_;
  assign new_n13476_ = new_n2733_ & new_n8100_;
  assign new_n13477_ = new_n7561_ & new_n10567_;
  assign new_n13478_ = ~new_n6272_ & ~new_n13477_;
  assign new_n13479_ = new_n13476_ & ~new_n13478_;
  assign new_n13480_ = new_n13473_ & ~new_n13479_;
  assign new_n13481_ = ~new_n6272_ & new_n13476_;
  assign new_n13482_ = ~pi0113 & new_n13481_;
  assign new_n13483_ = new_n13251_ & new_n13482_;
  assign new_n13484_ = ~new_n13480_ & ~new_n13483_;
  assign new_n13485_ = ~pi0039 & ~new_n13484_;
  assign new_n13486_ = new_n6258_ & ~new_n13485_;
  assign new_n13487_ = ~new_n13475_ & ~new_n13486_;
  assign new_n13488_ = ~new_n13472_ & new_n13487_;
  assign new_n13489_ = ~pi0087 & ~new_n13488_;
  assign new_n13490_ = ~new_n10594_ & new_n13473_;
  assign new_n13491_ = ~pi0113 & new_n13263_;
  assign new_n13492_ = ~new_n13490_ & ~new_n13491_;
  assign new_n13493_ = new_n3281_ & ~new_n13492_;
  assign new_n13494_ = ~new_n3211_ & new_n13474_;
  assign new_n13495_ = pi0087 & ~new_n13494_;
  assign new_n13496_ = ~new_n13493_ & new_n13495_;
  assign new_n13497_ = ~new_n13489_ & ~new_n13496_;
  assign new_n13498_ = ~pi0075 & ~new_n13497_;
  assign new_n13499_ = new_n7502_ & new_n13483_;
  assign new_n13500_ = ~new_n6272_ & ~new_n10607_;
  assign new_n13501_ = new_n13476_ & ~new_n13500_;
  assign new_n13502_ = new_n13473_ & ~new_n13501_;
  assign new_n13503_ = ~new_n13499_ & ~new_n13502_;
  assign new_n13504_ = new_n3227_ & ~new_n13503_;
  assign new_n13505_ = ~new_n3246_ & new_n13474_;
  assign new_n13506_ = pi0075 & ~new_n13505_;
  assign new_n13507_ = ~new_n13504_ & new_n13506_;
  assign new_n13508_ = ~new_n13498_ & ~new_n13507_;
  assign new_n13509_ = new_n8881_ & ~new_n13508_;
  assign new_n13510_ = ~new_n8881_ & ~new_n13474_;
  assign po0271 = ~new_n13509_ & ~new_n13510_;
  assign new_n13512_ = pi0114 & new_n10798_;
  assign new_n13513_ = new_n11153_ & ~new_n13512_;
  assign new_n13514_ = ~new_n10605_ & new_n13513_;
  assign new_n13515_ = ~pi0072 & pi0114;
  assign new_n13516_ = ~new_n11153_ & ~new_n13515_;
  assign new_n13517_ = new_n3227_ & ~new_n13516_;
  assign new_n13518_ = ~new_n13514_ & new_n13517_;
  assign new_n13519_ = ~pi0039 & new_n13515_;
  assign new_n13520_ = ~new_n3246_ & new_n13519_;
  assign new_n13521_ = pi0075 & ~new_n13520_;
  assign new_n13522_ = ~new_n13518_ & new_n13521_;
  assign new_n13523_ = ~pi0114 & ~new_n10749_;
  assign new_n13524_ = pi0114 & ~new_n10739_;
  assign new_n13525_ = ~new_n13523_ & ~new_n13524_;
  assign new_n13526_ = ~pi0115 & ~new_n13525_;
  assign new_n13527_ = pi0115 & ~new_n13515_;
  assign new_n13528_ = ~pi0039 & ~new_n13527_;
  assign new_n13529_ = ~new_n13526_ & new_n13528_;
  assign new_n13530_ = new_n3211_ & ~new_n13529_;
  assign new_n13531_ = pi0114 & ~new_n10570_;
  assign new_n13532_ = new_n11153_ & ~new_n13531_;
  assign new_n13533_ = ~new_n10565_ & new_n13532_;
  assign new_n13534_ = ~pi0039 & ~new_n13516_;
  assign new_n13535_ = ~new_n13533_ & new_n13534_;
  assign new_n13536_ = new_n6258_ & ~new_n13535_;
  assign new_n13537_ = pi0038 & ~new_n13519_;
  assign new_n13538_ = ~pi0087 & ~new_n13537_;
  assign new_n13539_ = ~new_n13536_ & new_n13538_;
  assign new_n13540_ = ~new_n13530_ & new_n13539_;
  assign new_n13541_ = pi0228 & new_n10568_;
  assign new_n13542_ = ~pi0115 & new_n13541_;
  assign new_n13543_ = new_n13515_ & ~new_n13542_;
  assign new_n13544_ = new_n3211_ & ~new_n13543_;
  assign new_n13545_ = ~new_n10592_ & new_n13544_;
  assign new_n13546_ = ~new_n3211_ & ~new_n13519_;
  assign new_n13547_ = new_n11127_ & ~new_n13546_;
  assign new_n13548_ = ~new_n13545_ & new_n13547_;
  assign new_n13549_ = ~pi0075 & ~new_n13548_;
  assign new_n13550_ = ~new_n13540_ & new_n13549_;
  assign new_n13551_ = ~new_n13522_ & ~new_n13550_;
  assign new_n13552_ = new_n8881_ & ~new_n13551_;
  assign new_n13553_ = ~new_n8881_ & ~new_n13519_;
  assign po0272 = ~new_n13552_ & ~new_n13553_;
  assign new_n13555_ = ~pi0052 & new_n11130_;
  assign new_n13556_ = ~pi0115 & ~new_n13555_;
  assign new_n13557_ = new_n10563_ & new_n13556_;
  assign new_n13558_ = new_n7502_ & new_n13557_;
  assign new_n13559_ = pi0115 & new_n10798_;
  assign new_n13560_ = new_n13476_ & ~new_n13559_;
  assign new_n13561_ = ~new_n13558_ & new_n13560_;
  assign new_n13562_ = ~pi0072 & pi0115;
  assign new_n13563_ = ~new_n13476_ & ~new_n13562_;
  assign new_n13564_ = new_n3227_ & ~new_n13563_;
  assign new_n13565_ = ~new_n13561_ & new_n13564_;
  assign new_n13566_ = ~pi0039 & new_n13562_;
  assign new_n13567_ = ~new_n3246_ & new_n13566_;
  assign new_n13568_ = pi0075 & ~new_n13567_;
  assign new_n13569_ = ~new_n13565_ & new_n13568_;
  assign new_n13570_ = pi0115 & ~new_n10739_;
  assign new_n13571_ = ~pi0115 & ~new_n10749_;
  assign new_n13572_ = ~pi0039 & ~new_n13571_;
  assign new_n13573_ = ~new_n13570_ & new_n13572_;
  assign new_n13574_ = new_n3211_ & ~new_n13573_;
  assign new_n13575_ = pi0115 & ~new_n10570_;
  assign new_n13576_ = new_n13476_ & ~new_n13575_;
  assign new_n13577_ = ~new_n13557_ & new_n13576_;
  assign new_n13578_ = ~pi0039 & ~new_n13563_;
  assign new_n13579_ = ~new_n13577_ & new_n13578_;
  assign new_n13580_ = new_n6258_ & ~new_n13579_;
  assign new_n13581_ = pi0038 & ~new_n13566_;
  assign new_n13582_ = ~pi0087 & ~new_n13581_;
  assign new_n13583_ = ~new_n13580_ & new_n13582_;
  assign new_n13584_ = ~new_n13574_ & new_n13583_;
  assign new_n13585_ = ~new_n13541_ & new_n13562_;
  assign new_n13586_ = new_n3211_ & ~new_n13585_;
  assign new_n13587_ = ~new_n10591_ & new_n13586_;
  assign new_n13588_ = ~new_n3211_ & ~new_n13566_;
  assign new_n13589_ = new_n11127_ & ~new_n13588_;
  assign new_n13590_ = ~new_n13587_ & new_n13589_;
  assign new_n13591_ = ~pi0075 & ~new_n13590_;
  assign new_n13592_ = ~new_n13584_ & new_n13591_;
  assign new_n13593_ = ~new_n13569_ & ~new_n13592_;
  assign new_n13594_ = new_n8881_ & ~new_n13593_;
  assign new_n13595_ = ~new_n8881_ & ~new_n13566_;
  assign po0273 = ~new_n13594_ & ~new_n13595_;
  assign new_n13597_ = pi0116 & new_n10511_;
  assign new_n13598_ = ~new_n2733_ & ~new_n13597_;
  assign new_n13599_ = new_n2733_ & ~new_n10495_;
  assign new_n13600_ = pi0116 & ~new_n13599_;
  assign new_n13601_ = ~new_n10502_ & ~new_n13600_;
  assign new_n13602_ = ~new_n13598_ & ~new_n13601_;
  assign new_n13603_ = ~new_n2733_ & new_n10516_;
  assign new_n13604_ = pi0228 & ~new_n13603_;
  assign new_n13605_ = ~new_n13602_ & new_n13604_;
  assign new_n13606_ = pi0116 & new_n10529_;
  assign new_n13607_ = new_n10743_ & ~new_n13606_;
  assign new_n13608_ = ~pi0039 & ~new_n13607_;
  assign new_n13609_ = ~new_n13605_ & new_n13608_;
  assign new_n13610_ = new_n3211_ & ~new_n13609_;
  assign new_n13611_ = ~pi0072 & pi0116;
  assign new_n13612_ = ~new_n13476_ & new_n13611_;
  assign new_n13613_ = ~pi0113 & new_n13477_;
  assign new_n13614_ = new_n13611_ & ~new_n13613_;
  assign new_n13615_ = ~new_n10563_ & ~new_n13614_;
  assign new_n13616_ = new_n13481_ & ~new_n13615_;
  assign new_n13617_ = ~new_n13612_ & ~new_n13616_;
  assign new_n13618_ = ~pi0039 & ~new_n13617_;
  assign new_n13619_ = new_n6258_ & ~new_n13618_;
  assign new_n13620_ = ~pi0039 & new_n13611_;
  assign new_n13621_ = pi0038 & ~new_n13620_;
  assign new_n13622_ = ~pi0087 & ~new_n13621_;
  assign new_n13623_ = ~new_n13619_ & new_n13622_;
  assign new_n13624_ = ~new_n13610_ & new_n13623_;
  assign new_n13625_ = ~pi0113 & new_n10594_;
  assign new_n13626_ = new_n13611_ & ~new_n13625_;
  assign new_n13627_ = ~pi0038 & ~new_n13626_;
  assign new_n13628_ = ~new_n10590_ & new_n13627_;
  assign new_n13629_ = ~new_n13621_ & ~new_n13628_;
  assign new_n13630_ = ~pi0100 & ~new_n13629_;
  assign new_n13631_ = pi0100 & ~new_n13620_;
  assign new_n13632_ = new_n11127_ & ~new_n13631_;
  assign new_n13633_ = ~new_n13630_ & new_n13632_;
  assign new_n13634_ = ~pi0075 & ~new_n13633_;
  assign new_n13635_ = ~new_n13624_ & new_n13634_;
  assign new_n13636_ = ~new_n10608_ & new_n13611_;
  assign new_n13637_ = ~new_n10800_ & ~new_n13636_;
  assign new_n13638_ = new_n13481_ & ~new_n13637_;
  assign new_n13639_ = ~new_n13612_ & ~new_n13638_;
  assign new_n13640_ = new_n3227_ & ~new_n13639_;
  assign new_n13641_ = ~new_n3246_ & new_n13620_;
  assign new_n13642_ = pi0075 & ~new_n13641_;
  assign new_n13643_ = ~new_n13640_ & new_n13642_;
  assign new_n13644_ = ~new_n13635_ & ~new_n13643_;
  assign new_n13645_ = new_n8881_ & ~new_n13644_;
  assign new_n13646_ = ~new_n8881_ & ~new_n13620_;
  assign po0274 = ~new_n13645_ & ~new_n13646_;
  assign new_n13648_ = new_n3671_ & new_n7364_;
  assign new_n13649_ = ~new_n3670_ & ~new_n13648_;
  assign new_n13650_ = ~pi0038 & ~new_n13649_;
  assign new_n13651_ = ~pi0087 & ~new_n13650_;
  assign new_n13652_ = new_n6289_ & ~new_n13651_;
  assign new_n13653_ = ~pi0092 & ~new_n13652_;
  assign new_n13654_ = ~pi0054 & ~new_n7305_;
  assign new_n13655_ = ~pi0074 & new_n13654_;
  assign new_n13656_ = ~new_n13653_ & new_n13655_;
  assign new_n13657_ = ~pi0055 & ~new_n13656_;
  assign new_n13658_ = ~new_n7347_ & ~new_n13657_;
  assign new_n13659_ = ~pi0056 & ~new_n13658_;
  assign new_n13660_ = ~new_n6127_ & ~new_n13659_;
  assign new_n13661_ = ~pi0062 & ~new_n13660_;
  assign new_n13662_ = ~pi0057 & new_n6300_;
  assign po0275 = ~new_n13661_ & new_n13662_;
  assign new_n13664_ = pi0163 & new_n6185_;
  assign new_n13665_ = ~new_n11678_ & ~new_n13664_;
  assign new_n13666_ = ~pi0150 & ~new_n13665_;
  assign new_n13667_ = pi0150 & new_n9699_;
  assign new_n13668_ = new_n11676_ & new_n13667_;
  assign new_n13669_ = ~new_n13666_ & ~new_n13668_;
  assign new_n13670_ = pi0232 & ~new_n13669_;
  assign new_n13671_ = ~new_n8989_ & new_n13670_;
  assign new_n13672_ = pi0074 & ~new_n13671_;
  assign new_n13673_ = pi0165 & new_n7499_;
  assign new_n13674_ = ~pi0038 & ~pi0054;
  assign new_n13675_ = ~new_n13673_ & ~new_n13674_;
  assign new_n13676_ = new_n8989_ & new_n13675_;
  assign new_n13677_ = ~pi0074 & ~new_n13671_;
  assign new_n13678_ = ~new_n13676_ & new_n13677_;
  assign new_n13679_ = ~new_n13672_ & ~new_n13678_;
  assign new_n13680_ = ~new_n3298_ & ~new_n13679_;
  assign new_n13681_ = new_n3436_ & ~new_n13680_;
  assign new_n13682_ = ~new_n9722_ & ~new_n13681_;
  assign new_n13683_ = pi0299 & new_n13669_;
  assign new_n13684_ = ~pi0184 & ~new_n11691_;
  assign new_n13685_ = ~pi0185 & new_n13684_;
  assign new_n13686_ = pi0185 & ~new_n13684_;
  assign new_n13687_ = new_n6185_ & ~new_n13686_;
  assign new_n13688_ = ~new_n13685_ & new_n13687_;
  assign new_n13689_ = ~pi0299 & ~new_n13688_;
  assign new_n13690_ = pi0232 & ~new_n13689_;
  assign new_n13691_ = ~new_n13683_ & new_n13690_;
  assign new_n13692_ = ~new_n8989_ & new_n13691_;
  assign new_n13693_ = pi0074 & ~new_n13692_;
  assign new_n13694_ = ~pi0055 & ~new_n13693_;
  assign new_n13695_ = ~pi0143 & ~pi0299;
  assign new_n13696_ = ~pi0165 & pi0299;
  assign new_n13697_ = ~new_n13695_ & ~new_n13696_;
  assign new_n13698_ = new_n7499_ & new_n13697_;
  assign new_n13699_ = new_n8989_ & ~new_n13698_;
  assign new_n13700_ = pi0054 & ~new_n13699_;
  assign new_n13701_ = ~new_n13692_ & new_n13700_;
  assign new_n13702_ = ~pi0143 & ~new_n9025_;
  assign new_n13703_ = pi0143 & ~new_n9027_;
  assign new_n13704_ = pi0165 & ~new_n13703_;
  assign new_n13705_ = ~new_n13702_ & new_n13704_;
  assign new_n13706_ = pi0143 & ~pi0165;
  assign new_n13707_ = new_n9032_ & new_n13706_;
  assign new_n13708_ = pi0038 & ~new_n13707_;
  assign new_n13709_ = ~new_n13705_ & new_n13708_;
  assign new_n13710_ = new_n3245_ & ~new_n13709_;
  assign new_n13711_ = ~new_n6185_ & new_n9337_;
  assign new_n13712_ = pi0151 & ~pi0168;
  assign new_n13713_ = ~new_n9403_ & new_n13712_;
  assign new_n13714_ = pi0168 & new_n9393_;
  assign new_n13715_ = ~pi0168 & new_n9396_;
  assign new_n13716_ = ~pi0151 & ~new_n13715_;
  assign new_n13717_ = ~new_n13714_ & new_n13716_;
  assign new_n13718_ = ~new_n13713_ & ~new_n13717_;
  assign new_n13719_ = ~new_n13711_ & ~new_n13718_;
  assign new_n13720_ = ~new_n6185_ & ~new_n9337_;
  assign new_n13721_ = new_n6185_ & ~new_n9363_;
  assign new_n13722_ = ~new_n13720_ & ~new_n13721_;
  assign new_n13723_ = pi0151 & pi0168;
  assign new_n13724_ = ~new_n13722_ & new_n13723_;
  assign new_n13725_ = pi0150 & ~new_n13724_;
  assign new_n13726_ = ~new_n13719_ & new_n13725_;
  assign new_n13727_ = ~new_n9233_ & ~new_n13720_;
  assign new_n13728_ = pi0168 & new_n13727_;
  assign new_n13729_ = ~new_n9422_ & ~new_n13720_;
  assign new_n13730_ = ~pi0168 & new_n13729_;
  assign new_n13731_ = pi0151 & ~new_n13730_;
  assign new_n13732_ = ~new_n13728_ & new_n13731_;
  assign new_n13733_ = pi0168 & new_n9331_;
  assign new_n13734_ = pi0168 & new_n6185_;
  assign new_n13735_ = new_n9337_ & ~new_n13734_;
  assign new_n13736_ = ~pi0151 & ~new_n13735_;
  assign new_n13737_ = ~new_n13733_ & new_n13736_;
  assign new_n13738_ = ~pi0150 & ~new_n13737_;
  assign new_n13739_ = ~new_n13732_ & new_n13738_;
  assign new_n13740_ = pi0299 & ~new_n13739_;
  assign new_n13741_ = ~new_n13726_ & new_n13740_;
  assign new_n13742_ = ~new_n9327_ & ~new_n13711_;
  assign new_n13743_ = ~pi0173 & ~new_n13742_;
  assign new_n13744_ = new_n6185_ & ~new_n9177_;
  assign new_n13745_ = pi0173 & ~new_n13720_;
  assign new_n13746_ = ~new_n13744_ & new_n13745_;
  assign new_n13747_ = pi0185 & ~new_n13746_;
  assign new_n13748_ = ~new_n13743_ & new_n13747_;
  assign new_n13749_ = pi0173 & new_n13727_;
  assign new_n13750_ = ~new_n9331_ & ~new_n13711_;
  assign new_n13751_ = ~pi0173 & ~new_n13750_;
  assign new_n13752_ = ~pi0185 & ~new_n13751_;
  assign new_n13753_ = ~new_n13749_ & new_n13752_;
  assign new_n13754_ = pi0190 & ~new_n13753_;
  assign new_n13755_ = ~new_n13748_ & new_n13754_;
  assign new_n13756_ = pi0173 & ~new_n9789_;
  assign new_n13757_ = ~pi0173 & ~new_n9349_;
  assign new_n13758_ = new_n6185_ & ~new_n13757_;
  assign new_n13759_ = ~new_n13756_ & new_n13758_;
  assign new_n13760_ = pi0185 & ~new_n13711_;
  assign new_n13761_ = ~new_n13759_ & new_n13760_;
  assign new_n13762_ = pi0173 & new_n13729_;
  assign new_n13763_ = ~pi0173 & new_n9337_;
  assign new_n13764_ = ~pi0185 & ~new_n13763_;
  assign new_n13765_ = ~new_n13762_ & new_n13764_;
  assign new_n13766_ = ~pi0190 & ~new_n13765_;
  assign new_n13767_ = ~new_n13761_ & new_n13766_;
  assign new_n13768_ = ~pi0299 & ~new_n13767_;
  assign new_n13769_ = ~new_n13755_ & new_n13768_;
  assign new_n13770_ = pi0232 & ~new_n13769_;
  assign new_n13771_ = ~new_n13741_ & new_n13770_;
  assign new_n13772_ = ~pi0232 & new_n9337_;
  assign new_n13773_ = ~pi0039 & ~new_n13772_;
  assign new_n13774_ = ~new_n13771_ & new_n13773_;
  assign new_n13775_ = ~pi0178 & ~pi0299;
  assign new_n13776_ = pi0168 & new_n9061_;
  assign new_n13777_ = pi0157 & new_n9072_;
  assign new_n13778_ = ~new_n13776_ & ~new_n13777_;
  assign new_n13779_ = new_n6185_ & new_n12118_;
  assign new_n13780_ = ~new_n13778_ & new_n13779_;
  assign new_n13781_ = pi0299 & ~new_n13780_;
  assign new_n13782_ = ~new_n13775_ & ~new_n13781_;
  assign new_n13783_ = new_n9038_ & ~new_n13782_;
  assign new_n13784_ = pi0178 & ~new_n9095_;
  assign new_n13785_ = ~pi0190 & ~new_n13784_;
  assign new_n13786_ = ~pi0299 & ~new_n13785_;
  assign new_n13787_ = ~new_n13783_ & ~new_n13786_;
  assign new_n13788_ = new_n6238_ & ~new_n9038_;
  assign new_n13789_ = new_n9058_ & ~new_n13788_;
  assign new_n13790_ = pi0178 & new_n13789_;
  assign new_n13791_ = ~new_n9102_ & new_n13790_;
  assign new_n13792_ = ~pi0178 & new_n13789_;
  assign new_n13793_ = ~new_n9064_ & new_n13792_;
  assign new_n13794_ = ~pi0299 & ~new_n9059_;
  assign new_n13795_ = pi0190 & new_n13794_;
  assign new_n13796_ = ~new_n13793_ & new_n13795_;
  assign new_n13797_ = ~new_n13791_ & new_n13796_;
  assign new_n13798_ = pi0232 & ~new_n13797_;
  assign new_n13799_ = ~new_n13787_ & new_n13798_;
  assign new_n13800_ = ~pi0232 & new_n9038_;
  assign new_n13801_ = pi0039 & ~new_n13800_;
  assign new_n13802_ = ~new_n13799_ & new_n13801_;
  assign new_n13803_ = ~pi0038 & ~new_n13802_;
  assign new_n13804_ = ~new_n13774_ & new_n13803_;
  assign new_n13805_ = new_n13710_ & ~new_n13804_;
  assign new_n13806_ = pi0100 & ~new_n13691_;
  assign new_n13807_ = pi0038 & ~new_n13698_;
  assign new_n13808_ = new_n7613_ & ~new_n13807_;
  assign new_n13809_ = ~new_n9521_ & new_n13808_;
  assign new_n13810_ = ~new_n13806_ & ~new_n13809_;
  assign new_n13811_ = ~new_n13805_ & new_n13810_;
  assign new_n13812_ = new_n3242_ & ~new_n13811_;
  assign new_n13813_ = pi0075 & ~new_n13691_;
  assign new_n13814_ = ~pi0100 & ~new_n13807_;
  assign new_n13815_ = ~pi0157 & pi0299;
  assign new_n13816_ = ~new_n13775_ & ~new_n13815_;
  assign new_n13817_ = new_n7499_ & new_n13816_;
  assign new_n13818_ = new_n9472_ & new_n13817_;
  assign new_n13819_ = new_n9521_ & ~new_n13818_;
  assign new_n13820_ = new_n13814_ & ~new_n13819_;
  assign new_n13821_ = ~new_n13806_ & ~new_n13820_;
  assign new_n13822_ = new_n9467_ & ~new_n13821_;
  assign new_n13823_ = ~new_n13813_ & ~new_n13822_;
  assign new_n13824_ = ~new_n13812_ & new_n13823_;
  assign new_n13825_ = ~pi0054 & ~new_n13824_;
  assign new_n13826_ = ~new_n13701_ & ~new_n13825_;
  assign new_n13827_ = ~pi0074 & ~new_n13826_;
  assign new_n13828_ = new_n13694_ & ~new_n13827_;
  assign new_n13829_ = pi0055 & ~new_n13672_;
  assign new_n13830_ = pi0150 & new_n7499_;
  assign new_n13831_ = ~pi0092 & new_n9472_;
  assign new_n13832_ = new_n13830_ & new_n13831_;
  assign new_n13833_ = new_n9038_ & new_n13674_;
  assign new_n13834_ = ~new_n13832_ & new_n13833_;
  assign new_n13835_ = ~new_n13675_ & ~new_n13834_;
  assign new_n13836_ = new_n8989_ & ~new_n13835_;
  assign new_n13837_ = new_n13677_ & ~new_n13836_;
  assign new_n13838_ = new_n13829_ & ~new_n13837_;
  assign new_n13839_ = new_n3298_ & ~new_n13838_;
  assign new_n13840_ = ~new_n13828_ & new_n13839_;
  assign new_n13841_ = ~new_n13682_ & ~new_n13840_;
  assign new_n13842_ = ~new_n8989_ & ~new_n13670_;
  assign new_n13843_ = new_n8989_ & new_n13673_;
  assign new_n13844_ = ~new_n3436_ & ~new_n13843_;
  assign new_n13845_ = ~new_n13842_ & new_n13844_;
  assign new_n13846_ = ~new_n13672_ & new_n13845_;
  assign new_n13847_ = ~new_n13841_ & ~new_n13846_;
  assign new_n13848_ = pi0118 & new_n13847_;
  assign new_n13849_ = ~pi0079 & new_n12169_;
  assign new_n13850_ = new_n6221_ & ~new_n6466_;
  assign new_n13851_ = ~pi0157 & new_n9551_;
  assign new_n13852_ = pi0168 & ~new_n13851_;
  assign new_n13853_ = pi0157 & ~new_n9546_;
  assign new_n13854_ = ~pi0157 & ~pi0168;
  assign new_n13855_ = ~new_n9544_ & new_n13854_;
  assign new_n13856_ = ~new_n13853_ & ~new_n13855_;
  assign new_n13857_ = ~new_n13852_ & new_n13856_;
  assign new_n13858_ = ~new_n13850_ & ~new_n13857_;
  assign new_n13859_ = new_n13130_ & ~new_n13858_;
  assign new_n13860_ = ~pi0178 & ~new_n6238_;
  assign new_n13861_ = new_n9550_ & new_n13860_;
  assign new_n13862_ = ~new_n13850_ & ~new_n13861_;
  assign new_n13863_ = pi0190 & ~new_n13862_;
  assign new_n13864_ = ~pi0178 & ~new_n13164_;
  assign new_n13865_ = pi0178 & ~new_n9529_;
  assign new_n13866_ = ~new_n13850_ & new_n13865_;
  assign new_n13867_ = ~pi0190 & ~new_n13866_;
  assign new_n13868_ = ~new_n13864_ & new_n13867_;
  assign new_n13869_ = ~new_n13863_ & ~new_n13868_;
  assign new_n13870_ = new_n13132_ & ~new_n13869_;
  assign new_n13871_ = pi0232 & ~new_n13870_;
  assign new_n13872_ = ~new_n13859_ & new_n13871_;
  assign new_n13873_ = new_n7309_ & new_n9534_;
  assign new_n13874_ = ~new_n6223_ & new_n13130_;
  assign new_n13875_ = ~new_n6466_ & new_n13874_;
  assign new_n13876_ = ~pi0232 & ~new_n13875_;
  assign new_n13877_ = ~new_n13873_ & new_n13876_;
  assign new_n13878_ = pi0039 & ~new_n13877_;
  assign new_n13879_ = ~new_n13872_ & new_n13878_;
  assign new_n13880_ = new_n9607_ & new_n13712_;
  assign new_n13881_ = ~pi0168 & ~new_n9579_;
  assign new_n13882_ = pi0168 & ~new_n9593_;
  assign new_n13883_ = ~pi0151 & ~new_n13882_;
  assign new_n13884_ = ~new_n13881_ & new_n13883_;
  assign new_n13885_ = ~new_n13880_ & ~new_n13884_;
  assign new_n13886_ = new_n9581_ & ~new_n13885_;
  assign new_n13887_ = pi0150 & ~new_n13886_;
  assign new_n13888_ = ~pi0151 & new_n9570_;
  assign new_n13889_ = new_n9621_ & ~new_n13888_;
  assign new_n13890_ = ~pi0168 & ~new_n13889_;
  assign new_n13891_ = ~pi0151 & new_n9589_;
  assign new_n13892_ = new_n9624_ & ~new_n13891_;
  assign new_n13893_ = new_n13734_ & ~new_n13892_;
  assign new_n13894_ = ~pi0150 & ~new_n13893_;
  assign new_n13895_ = ~new_n13890_ & new_n13894_;
  assign new_n13896_ = ~new_n13887_ & ~new_n13895_;
  assign new_n13897_ = ~new_n9570_ & ~new_n12035_;
  assign new_n13898_ = ~new_n6185_ & ~new_n13897_;
  assign new_n13899_ = pi0299 & ~new_n13898_;
  assign new_n13900_ = ~new_n13896_ & new_n13899_;
  assign new_n13901_ = new_n6379_ & new_n9607_;
  assign new_n13902_ = pi0173 & new_n13901_;
  assign new_n13903_ = ~pi0173 & new_n6379_;
  assign new_n13904_ = new_n9579_ & new_n13903_;
  assign new_n13905_ = ~new_n13902_ & ~new_n13904_;
  assign new_n13906_ = ~pi0190 & new_n6185_;
  assign new_n13907_ = ~new_n13905_ & new_n13906_;
  assign new_n13908_ = ~pi0173 & pi0190;
  assign new_n13909_ = new_n9594_ & new_n13908_;
  assign new_n13910_ = pi0185 & ~new_n13909_;
  assign new_n13911_ = ~new_n13907_ & new_n13910_;
  assign new_n13912_ = ~pi0173 & new_n9570_;
  assign new_n13913_ = new_n9600_ & ~new_n13912_;
  assign new_n13914_ = ~pi0190 & ~new_n13913_;
  assign new_n13915_ = pi0173 & new_n9603_;
  assign new_n13916_ = pi0190 & new_n9591_;
  assign new_n13917_ = ~new_n13915_ & new_n13916_;
  assign new_n13918_ = ~pi0185 & ~new_n13917_;
  assign new_n13919_ = ~new_n13914_ & new_n13918_;
  assign new_n13920_ = ~new_n13911_ & ~new_n13919_;
  assign new_n13921_ = ~new_n6185_ & ~new_n9574_;
  assign new_n13922_ = ~pi0299 & ~new_n13921_;
  assign new_n13923_ = ~new_n13920_ & new_n13922_;
  assign new_n13924_ = ~new_n13900_ & ~new_n13923_;
  assign new_n13925_ = pi0232 & ~new_n13924_;
  assign new_n13926_ = ~new_n6166_ & ~new_n9572_;
  assign new_n13927_ = ~pi0232 & ~new_n9570_;
  assign new_n13928_ = ~new_n13926_ & new_n13927_;
  assign new_n13929_ = ~pi0039 & ~new_n13928_;
  assign new_n13930_ = ~new_n13925_ & new_n13929_;
  assign new_n13931_ = ~new_n13879_ & ~new_n13930_;
  assign new_n13932_ = ~pi0038 & ~new_n13931_;
  assign new_n13933_ = new_n13710_ & ~new_n13932_;
  assign new_n13934_ = ~new_n13806_ & ~new_n13808_;
  assign new_n13935_ = ~new_n13933_ & new_n13934_;
  assign new_n13936_ = new_n3242_ & ~new_n13935_;
  assign new_n13937_ = new_n8965_ & ~new_n13817_;
  assign new_n13938_ = new_n3100_ & new_n13937_;
  assign new_n13939_ = new_n13814_ & ~new_n13938_;
  assign new_n13940_ = ~new_n13806_ & ~new_n13939_;
  assign new_n13941_ = new_n9467_ & ~new_n13940_;
  assign new_n13942_ = ~new_n13813_ & ~new_n13941_;
  assign new_n13943_ = ~new_n13936_ & new_n13942_;
  assign new_n13944_ = ~pi0054 & ~new_n13943_;
  assign new_n13945_ = ~new_n13701_ & ~new_n13944_;
  assign new_n13946_ = ~pi0074 & ~new_n13945_;
  assign new_n13947_ = new_n13694_ & ~new_n13946_;
  assign new_n13948_ = pi0054 & new_n13673_;
  assign new_n13949_ = ~pi0092 & new_n8989_;
  assign new_n13950_ = new_n8965_ & new_n13949_;
  assign new_n13951_ = ~new_n13830_ & new_n13950_;
  assign new_n13952_ = ~new_n13948_ & new_n13951_;
  assign new_n13953_ = new_n3100_ & new_n13952_;
  assign new_n13954_ = new_n13678_ & ~new_n13953_;
  assign new_n13955_ = new_n13829_ & ~new_n13954_;
  assign new_n13956_ = new_n3298_ & ~new_n13955_;
  assign new_n13957_ = ~new_n13947_ & new_n13956_;
  assign new_n13958_ = new_n13681_ & ~new_n13957_;
  assign new_n13959_ = ~new_n13846_ & ~new_n13958_;
  assign new_n13960_ = ~pi0118 & new_n13959_;
  assign new_n13961_ = ~new_n13849_ & ~new_n13960_;
  assign new_n13962_ = ~new_n13848_ & new_n13961_;
  assign new_n13963_ = ~pi0118 & ~new_n8976_;
  assign new_n13964_ = new_n13847_ & new_n13963_;
  assign new_n13965_ = new_n13959_ & ~new_n13963_;
  assign new_n13966_ = new_n13849_ & ~new_n13965_;
  assign new_n13967_ = ~new_n13964_ & new_n13966_;
  assign po0276 = new_n13962_ | new_n13967_;
  assign new_n13969_ = pi0128 & pi0228;
  assign new_n13970_ = ~new_n10163_ & new_n13969_;
  assign new_n13971_ = ~new_n3057_ & new_n3489_;
  assign new_n13972_ = new_n7545_ & new_n13971_;
  assign new_n13973_ = ~new_n3467_ & new_n5788_;
  assign new_n13974_ = new_n7549_ & new_n13973_;
  assign new_n13975_ = ~new_n13972_ & ~new_n13974_;
  assign new_n13976_ = pi0039 & ~new_n13975_;
  assign new_n13977_ = new_n2579_ & new_n10157_;
  assign new_n13978_ = new_n11664_ & ~new_n13977_;
  assign new_n13979_ = new_n2592_ & ~new_n13978_;
  assign new_n13980_ = ~pi0097 & ~new_n13979_;
  assign new_n13981_ = ~pi0046 & new_n2795_;
  assign new_n13982_ = new_n2758_ & new_n13981_;
  assign new_n13983_ = ~new_n13980_ & new_n13982_;
  assign new_n13984_ = pi0299 & new_n6431_;
  assign new_n13985_ = ~new_n6397_ & ~new_n13984_;
  assign new_n13986_ = new_n7499_ & ~new_n13985_;
  assign new_n13987_ = pi0109 & ~new_n13986_;
  assign new_n13988_ = ~new_n2795_ & new_n11665_;
  assign new_n13989_ = ~new_n13987_ & ~new_n13988_;
  assign new_n13990_ = ~new_n13983_ & new_n13989_;
  assign new_n13991_ = ~new_n6320_ & ~new_n13986_;
  assign new_n13992_ = ~new_n6401_ & new_n13986_;
  assign new_n13993_ = ~new_n13991_ & ~new_n13992_;
  assign new_n13994_ = ~new_n13990_ & new_n13993_;
  assign new_n13995_ = ~pi0091 & ~new_n13994_;
  assign new_n13996_ = new_n2536_ & ~new_n6355_;
  assign new_n13997_ = ~new_n13995_ & new_n13996_;
  assign new_n13998_ = ~new_n2563_ & ~new_n13997_;
  assign new_n13999_ = ~pi0039 & new_n11086_;
  assign new_n14000_ = ~new_n13998_ & new_n13999_;
  assign new_n14001_ = ~new_n13976_ & ~new_n14000_;
  assign new_n14002_ = ~pi0038 & ~new_n14001_;
  assign new_n14003_ = ~pi0228 & new_n14002_;
  assign new_n14004_ = ~new_n13969_ & ~new_n14003_;
  assign new_n14005_ = ~pi0100 & ~new_n14004_;
  assign new_n14006_ = new_n3186_ & new_n3326_;
  assign new_n14007_ = ~new_n13969_ & ~new_n14006_;
  assign new_n14008_ = pi0100 & ~new_n14007_;
  assign new_n14009_ = ~pi0087 & ~new_n14008_;
  assign new_n14010_ = ~new_n14005_ & new_n14009_;
  assign new_n14011_ = pi0087 & ~new_n13969_;
  assign new_n14012_ = ~pi0075 & ~new_n14011_;
  assign new_n14013_ = ~new_n14010_ & new_n14012_;
  assign new_n14014_ = new_n7369_ & new_n8965_;
  assign new_n14015_ = ~new_n13969_ & ~new_n14014_;
  assign new_n14016_ = pi0075 & ~new_n14015_;
  assign new_n14017_ = ~pi0092 & ~new_n14016_;
  assign new_n14018_ = ~new_n14013_ & new_n14017_;
  assign new_n14019_ = pi0092 & ~new_n13969_;
  assign new_n14020_ = ~new_n7382_ & new_n14019_;
  assign new_n14021_ = new_n10163_ & ~new_n14020_;
  assign new_n14022_ = ~new_n14018_ & new_n14021_;
  assign po0277 = new_n13970_ | new_n14022_;
  assign new_n14024_ = ~pi0031 & ~pi0080;
  assign new_n14025_ = pi0818 & new_n14024_;
  assign new_n14026_ = ~new_n7455_ & new_n8057_;
  assign new_n14027_ = ~new_n7733_ & ~new_n14026_;
  assign new_n14028_ = ~pi0120 & ~new_n7455_;
  assign new_n14029_ = ~pi1093 & new_n14028_;
  assign new_n14030_ = new_n14027_ & ~new_n14029_;
  assign new_n14031_ = new_n3100_ & new_n7505_;
  assign new_n14032_ = pi0120 & ~new_n8057_;
  assign new_n14033_ = ~new_n7564_ & new_n14032_;
  assign new_n14034_ = new_n14031_ & ~new_n14033_;
  assign new_n14035_ = ~pi0120 & pi1093;
  assign new_n14036_ = new_n7564_ & ~new_n14035_;
  assign new_n14037_ = ~new_n14034_ & ~new_n14036_;
  assign new_n14038_ = new_n3186_ & new_n8100_;
  assign new_n14039_ = ~new_n14037_ & new_n14038_;
  assign new_n14040_ = ~pi1091 & new_n12801_;
  assign new_n14041_ = new_n14035_ & ~new_n14040_;
  assign new_n14042_ = ~new_n14032_ & ~new_n14041_;
  assign new_n14043_ = pi0100 & ~new_n14042_;
  assign new_n14044_ = ~new_n14039_ & new_n14043_;
  assign new_n14045_ = ~pi1093 & new_n7486_;
  assign new_n14046_ = pi0120 & new_n14045_;
  assign new_n14047_ = ~pi0039 & ~new_n14046_;
  assign new_n14048_ = new_n7528_ & ~new_n10352_;
  assign new_n14049_ = new_n7477_ & new_n7511_;
  assign new_n14050_ = ~pi0829 & new_n14049_;
  assign new_n14051_ = ~pi0122 & ~new_n14050_;
  assign new_n14052_ = ~new_n14048_ & new_n14051_;
  assign new_n14053_ = pi0122 & ~new_n7478_;
  assign new_n14054_ = ~new_n2732_ & ~new_n14053_;
  assign new_n14055_ = ~new_n14052_ & new_n14054_;
  assign new_n14056_ = new_n2797_ & ~new_n14055_;
  assign new_n14057_ = new_n7572_ & ~new_n14049_;
  assign new_n14058_ = ~new_n12801_ & new_n14057_;
  assign new_n14059_ = ~new_n14056_ & ~new_n14058_;
  assign new_n14060_ = new_n14047_ & new_n14059_;
  assign new_n14061_ = new_n6215_ & ~new_n14042_;
  assign new_n14062_ = ~new_n7544_ & new_n14032_;
  assign new_n14063_ = pi1091 & pi1092;
  assign new_n14064_ = new_n7542_ & new_n14063_;
  assign new_n14065_ = new_n14041_ & ~new_n14064_;
  assign new_n14066_ = ~new_n14062_ & ~new_n14065_;
  assign new_n14067_ = ~new_n6215_ & ~new_n14066_;
  assign new_n14068_ = ~new_n14061_ & ~new_n14067_;
  assign new_n14069_ = ~new_n6238_ & ~new_n14068_;
  assign new_n14070_ = ~new_n6221_ & new_n14042_;
  assign new_n14071_ = new_n6221_ & new_n14066_;
  assign new_n14072_ = ~new_n14070_ & ~new_n14071_;
  assign new_n14073_ = new_n6238_ & new_n14072_;
  assign new_n14074_ = new_n8086_ & ~new_n14073_;
  assign new_n14075_ = ~new_n14069_ & new_n14074_;
  assign new_n14076_ = ~new_n8086_ & new_n14042_;
  assign new_n14077_ = ~pi0299 & ~new_n14076_;
  assign new_n14078_ = ~new_n14075_ & new_n14077_;
  assign new_n14079_ = ~new_n6212_ & ~new_n14068_;
  assign new_n14080_ = new_n6212_ & new_n14072_;
  assign new_n14081_ = new_n8075_ & ~new_n14080_;
  assign new_n14082_ = ~new_n14079_ & new_n14081_;
  assign new_n14083_ = ~new_n8075_ & new_n14042_;
  assign new_n14084_ = pi0299 & ~new_n14083_;
  assign new_n14085_ = ~new_n14082_ & new_n14084_;
  assign new_n14086_ = pi0039 & ~new_n14085_;
  assign new_n14087_ = ~new_n14078_ & new_n14086_;
  assign new_n14088_ = ~new_n14060_ & ~new_n14087_;
  assign new_n14089_ = ~pi0038 & ~new_n14088_;
  assign new_n14090_ = pi0038 & new_n8057_;
  assign new_n14091_ = ~pi0120 & ~pi1093;
  assign new_n14092_ = pi0038 & new_n14091_;
  assign new_n14093_ = ~pi0100 & ~new_n14092_;
  assign new_n14094_ = ~new_n14090_ & new_n14093_;
  assign new_n14095_ = ~new_n14089_ & new_n14094_;
  assign new_n14096_ = ~new_n14044_ & ~new_n14095_;
  assign new_n14097_ = ~pi0087 & ~new_n14096_;
  assign new_n14098_ = new_n7580_ & ~new_n14091_;
  assign new_n14099_ = new_n7572_ & ~new_n12801_;
  assign new_n14100_ = ~new_n8112_ & new_n14099_;
  assign new_n14101_ = new_n7578_ & ~new_n14100_;
  assign new_n14102_ = ~new_n3212_ & new_n8057_;
  assign new_n14103_ = pi0087 & ~new_n14102_;
  assign new_n14104_ = ~new_n14101_ & new_n14103_;
  assign new_n14105_ = new_n14098_ & new_n14104_;
  assign new_n14106_ = ~new_n14097_ & ~new_n14105_;
  assign new_n14107_ = ~pi0075 & ~new_n14106_;
  assign new_n14108_ = new_n7500_ & new_n14042_;
  assign new_n14109_ = ~new_n7506_ & new_n14041_;
  assign new_n14110_ = ~pi1091 & ~new_n8056_;
  assign new_n14111_ = ~new_n8049_ & ~new_n14110_;
  assign new_n14112_ = pi0120 & ~new_n14111_;
  assign new_n14113_ = ~new_n7500_ & ~new_n14112_;
  assign new_n14114_ = ~new_n14109_ & new_n14113_;
  assign new_n14115_ = ~new_n14108_ & ~new_n14114_;
  assign new_n14116_ = new_n3227_ & ~new_n14115_;
  assign new_n14117_ = ~new_n3227_ & new_n14042_;
  assign new_n14118_ = pi0075 & ~new_n14117_;
  assign new_n14119_ = ~new_n14116_ & new_n14118_;
  assign new_n14120_ = new_n7455_ & ~new_n14119_;
  assign new_n14121_ = ~new_n14107_ & new_n14120_;
  assign new_n14122_ = new_n14030_ & ~new_n14121_;
  assign new_n14123_ = ~new_n14056_ & ~new_n14057_;
  assign new_n14124_ = new_n14047_ & new_n14123_;
  assign new_n14125_ = pi1093 & ~new_n6221_;
  assign new_n14126_ = new_n6238_ & new_n14125_;
  assign new_n14127_ = new_n6215_ & ~new_n6238_;
  assign new_n14128_ = new_n8086_ & ~new_n14127_;
  assign new_n14129_ = ~new_n14126_ & new_n14128_;
  assign new_n14130_ = new_n7544_ & new_n14129_;
  assign new_n14131_ = ~pi0299 & ~new_n14091_;
  assign new_n14132_ = ~new_n14130_ & new_n14131_;
  assign new_n14133_ = new_n6212_ & new_n14125_;
  assign new_n14134_ = ~new_n6212_ & new_n6215_;
  assign new_n14135_ = new_n8075_ & ~new_n14134_;
  assign new_n14136_ = ~new_n14133_ & new_n14135_;
  assign new_n14137_ = new_n7544_ & new_n14136_;
  assign new_n14138_ = pi0299 & ~new_n14091_;
  assign new_n14139_ = ~new_n14137_ & new_n14138_;
  assign new_n14140_ = pi0039 & ~new_n14139_;
  assign new_n14141_ = ~new_n14132_ & new_n14140_;
  assign new_n14142_ = ~new_n14124_ & ~new_n14141_;
  assign new_n14143_ = ~pi0038 & ~new_n14142_;
  assign new_n14144_ = new_n14093_ & ~new_n14143_;
  assign new_n14145_ = pi0120 & new_n7564_;
  assign new_n14146_ = ~pi0120 & new_n14031_;
  assign new_n14147_ = ~new_n14145_ & ~new_n14146_;
  assign new_n14148_ = new_n14038_ & ~new_n14147_;
  assign new_n14149_ = pi0100 & ~new_n14091_;
  assign new_n14150_ = ~new_n14148_ & new_n14149_;
  assign new_n14151_ = ~new_n14144_ & ~new_n14150_;
  assign new_n14152_ = ~pi0087 & ~new_n14151_;
  assign new_n14153_ = ~new_n14098_ & ~new_n14152_;
  assign new_n14154_ = ~pi0075 & ~new_n14153_;
  assign new_n14155_ = new_n7509_ & ~new_n14091_;
  assign new_n14156_ = new_n7455_ & ~new_n14155_;
  assign new_n14157_ = ~new_n14154_ & new_n14156_;
  assign new_n14158_ = new_n7733_ & ~new_n14029_;
  assign new_n14159_ = ~new_n14157_ & new_n14158_;
  assign new_n14160_ = ~new_n14122_ & ~new_n14159_;
  assign new_n14161_ = new_n14025_ & ~new_n14160_;
  assign new_n14162_ = ~po1038 & ~new_n14161_;
  assign new_n14163_ = ~new_n7733_ & new_n14042_;
  assign new_n14164_ = pi0120 & ~new_n14163_;
  assign new_n14165_ = new_n14025_ & ~new_n14091_;
  assign new_n14166_ = ~new_n14163_ & new_n14165_;
  assign new_n14167_ = po1038 & ~new_n14166_;
  assign new_n14168_ = ~new_n14164_ & new_n14167_;
  assign new_n14169_ = ~new_n8870_ & ~new_n14168_;
  assign new_n14170_ = pi0951 & pi0982;
  assign new_n14171_ = pi1092 & new_n14170_;
  assign new_n14172_ = pi1093 & new_n14171_;
  assign new_n14173_ = ~pi0120 & ~new_n14172_;
  assign new_n14174_ = ~new_n14163_ & ~new_n14173_;
  assign new_n14175_ = new_n14167_ & ~new_n14174_;
  assign new_n14176_ = new_n8870_ & ~new_n14175_;
  assign new_n14177_ = ~new_n14169_ & ~new_n14176_;
  assign new_n14178_ = ~new_n14162_ & ~new_n14177_;
  assign new_n14179_ = pi0120 & new_n7507_;
  assign new_n14180_ = ~pi1091 & new_n14172_;
  assign new_n14181_ = ~pi0120 & ~new_n14180_;
  assign new_n14182_ = new_n2797_ & new_n14171_;
  assign new_n14183_ = ~pi0093 & ~pi0122;
  assign new_n14184_ = new_n2549_ & new_n14183_;
  assign new_n14185_ = new_n2753_ & new_n8894_;
  assign new_n14186_ = new_n14184_ & new_n14185_;
  assign new_n14187_ = new_n2535_ & new_n14186_;
  assign new_n14188_ = new_n10310_ & new_n14187_;
  assign new_n14189_ = new_n7503_ & new_n14188_;
  assign new_n14190_ = new_n2492_ & new_n14189_;
  assign new_n14191_ = new_n14182_ & ~new_n14190_;
  assign new_n14192_ = new_n14181_ & ~new_n14191_;
  assign new_n14193_ = ~new_n14179_ & ~new_n14192_;
  assign new_n14194_ = ~new_n7500_ & ~new_n14193_;
  assign new_n14195_ = new_n7500_ & new_n14173_;
  assign new_n14196_ = new_n3227_ & ~new_n14195_;
  assign new_n14197_ = ~new_n14194_ & new_n14196_;
  assign new_n14198_ = ~new_n3227_ & ~new_n14173_;
  assign new_n14199_ = pi0075 & ~new_n14198_;
  assign new_n14200_ = ~new_n14197_ & new_n14199_;
  assign new_n14201_ = pi0950 & new_n3100_;
  assign new_n14202_ = new_n7456_ & new_n7503_;
  assign new_n14203_ = new_n14201_ & new_n14202_;
  assign new_n14204_ = new_n14182_ & ~new_n14203_;
  assign new_n14205_ = new_n14181_ & ~new_n14204_;
  assign new_n14206_ = ~new_n14145_ & ~new_n14205_;
  assign new_n14207_ = ~pi0039 & new_n8100_;
  assign new_n14208_ = ~new_n14206_ & new_n14207_;
  assign new_n14209_ = pi0100 & ~new_n14208_;
  assign new_n14210_ = ~pi0038 & ~new_n14209_;
  assign new_n14211_ = ~new_n14038_ & new_n14173_;
  assign new_n14212_ = ~new_n14210_ & ~new_n14211_;
  assign new_n14213_ = ~new_n8086_ & new_n14173_;
  assign new_n14214_ = ~pi0299 & ~new_n14213_;
  assign new_n14215_ = ~new_n8274_ & ~new_n14173_;
  assign new_n14216_ = new_n6238_ & new_n14215_;
  assign new_n14217_ = ~new_n8270_ & ~new_n14173_;
  assign new_n14218_ = ~new_n6238_ & new_n14217_;
  assign new_n14219_ = new_n8086_ & ~new_n14218_;
  assign new_n14220_ = ~new_n14216_ & new_n14219_;
  assign new_n14221_ = new_n14214_ & ~new_n14220_;
  assign new_n14222_ = ~new_n8075_ & new_n14173_;
  assign new_n14223_ = pi0299 & ~new_n14222_;
  assign new_n14224_ = new_n6212_ & new_n14215_;
  assign new_n14225_ = ~new_n6212_ & new_n14217_;
  assign new_n14226_ = new_n8075_ & ~new_n14225_;
  assign new_n14227_ = ~new_n14224_ & new_n14226_;
  assign new_n14228_ = new_n14223_ & ~new_n14227_;
  assign new_n14229_ = ~new_n14221_ & ~new_n14228_;
  assign new_n14230_ = pi0039 & ~new_n14229_;
  assign new_n14231_ = ~new_n14045_ & new_n14123_;
  assign new_n14232_ = pi0120 & new_n14231_;
  assign new_n14233_ = new_n2580_ & new_n7466_;
  assign new_n14234_ = new_n2576_ & new_n14233_;
  assign new_n14235_ = ~pi0097 & ~new_n14234_;
  assign new_n14236_ = new_n2761_ & ~new_n14235_;
  assign new_n14237_ = new_n2759_ & new_n14236_;
  assign new_n14238_ = ~new_n7516_ & ~new_n14237_;
  assign new_n14239_ = new_n2518_ & ~new_n14238_;
  assign new_n14240_ = new_n7460_ & ~new_n14239_;
  assign new_n14241_ = new_n7457_ & ~new_n14240_;
  assign new_n14242_ = ~pi0051 & ~new_n14241_;
  assign new_n14243_ = ~new_n2558_ & ~new_n14242_;
  assign new_n14244_ = ~pi0096 & ~new_n14243_;
  assign new_n14245_ = ~pi0072 & pi0950;
  assign new_n14246_ = new_n10353_ & new_n14245_;
  assign new_n14247_ = ~new_n14244_ & new_n14246_;
  assign new_n14248_ = new_n7456_ & new_n14171_;
  assign new_n14249_ = ~new_n14247_ & new_n14248_;
  assign new_n14250_ = new_n9562_ & new_n14234_;
  assign new_n14251_ = new_n7457_ & new_n14250_;
  assign new_n14252_ = new_n7462_ & ~new_n14251_;
  assign new_n14253_ = pi0950 & new_n7512_;
  assign new_n14254_ = ~new_n14252_ & new_n14253_;
  assign new_n14255_ = pi0824 & new_n14254_;
  assign new_n14256_ = new_n14171_ & ~new_n14255_;
  assign new_n14257_ = ~pi0829 & new_n14256_;
  assign new_n14258_ = pi0829 & pi1092;
  assign new_n14259_ = pi0122 & new_n14170_;
  assign new_n14260_ = new_n14258_ & new_n14259_;
  assign new_n14261_ = ~new_n14254_ & new_n14260_;
  assign new_n14262_ = ~new_n14257_ & ~new_n14261_;
  assign new_n14263_ = ~new_n14249_ & new_n14262_;
  assign new_n14264_ = new_n7510_ & ~new_n14263_;
  assign new_n14265_ = new_n2732_ & new_n14172_;
  assign new_n14266_ = ~new_n14264_ & ~new_n14265_;
  assign new_n14267_ = pi1091 & ~new_n14266_;
  assign new_n14268_ = new_n14180_ & ~new_n14255_;
  assign new_n14269_ = ~pi0120 & ~new_n14268_;
  assign new_n14270_ = ~new_n14267_ & new_n14269_;
  assign new_n14271_ = ~pi0039 & ~new_n14270_;
  assign new_n14272_ = ~new_n14232_ & new_n14271_;
  assign new_n14273_ = ~new_n14230_ & ~new_n14272_;
  assign new_n14274_ = new_n3211_ & ~new_n14273_;
  assign new_n14275_ = ~new_n14212_ & ~new_n14274_;
  assign new_n14276_ = ~pi0087 & ~new_n14275_;
  assign new_n14277_ = ~new_n3212_ & new_n14173_;
  assign new_n14278_ = pi0087 & ~new_n14277_;
  assign new_n14279_ = ~new_n2732_ & ~new_n6194_;
  assign new_n14280_ = new_n14201_ & new_n14279_;
  assign new_n14281_ = new_n14182_ & ~new_n14280_;
  assign new_n14282_ = pi0824 & new_n14201_;
  assign new_n14283_ = new_n14180_ & ~new_n14282_;
  assign new_n14284_ = ~new_n14281_ & ~new_n14283_;
  assign new_n14285_ = ~pi0120 & ~new_n14284_;
  assign new_n14286_ = ~new_n7573_ & ~new_n7577_;
  assign new_n14287_ = pi0120 & ~new_n14286_;
  assign new_n14288_ = new_n3212_ & ~new_n14287_;
  assign new_n14289_ = ~new_n14285_ & new_n14288_;
  assign new_n14290_ = new_n14278_ & ~new_n14289_;
  assign new_n14291_ = ~pi0075 & ~new_n14290_;
  assign new_n14292_ = ~new_n14276_ & new_n14291_;
  assign new_n14293_ = ~new_n14200_ & ~new_n14292_;
  assign new_n14294_ = new_n7455_ & ~new_n14293_;
  assign new_n14295_ = new_n7733_ & ~new_n14294_;
  assign new_n14296_ = ~new_n12801_ & new_n14180_;
  assign new_n14297_ = ~new_n14204_ & ~new_n14296_;
  assign new_n14298_ = ~pi0120 & ~new_n14297_;
  assign new_n14299_ = ~new_n14033_ & ~new_n14298_;
  assign new_n14300_ = new_n8100_ & ~new_n14299_;
  assign new_n14301_ = ~new_n14042_ & ~new_n14173_;
  assign new_n14302_ = ~new_n8100_ & new_n14301_;
  assign new_n14303_ = new_n3186_ & ~new_n14302_;
  assign new_n14304_ = ~new_n14300_ & new_n14303_;
  assign new_n14305_ = ~new_n3186_ & ~new_n14301_;
  assign new_n14306_ = pi0100 & ~new_n14305_;
  assign new_n14307_ = ~new_n14304_ & new_n14306_;
  assign new_n14308_ = ~new_n14045_ & new_n14059_;
  assign new_n14309_ = pi0120 & new_n14308_;
  assign new_n14310_ = new_n14099_ & new_n14256_;
  assign new_n14311_ = ~pi0120 & ~new_n14310_;
  assign new_n14312_ = ~new_n14267_ & new_n14311_;
  assign new_n14313_ = ~new_n14309_ & ~new_n14312_;
  assign new_n14314_ = ~pi0039 & ~new_n14313_;
  assign new_n14315_ = ~new_n7542_ & new_n14182_;
  assign new_n14316_ = ~new_n14296_ & ~new_n14315_;
  assign new_n14317_ = ~pi0120 & ~new_n14316_;
  assign new_n14318_ = ~new_n14062_ & ~new_n14317_;
  assign new_n14319_ = ~new_n6215_ & ~new_n14318_;
  assign new_n14320_ = new_n6215_ & new_n14301_;
  assign new_n14321_ = ~new_n14319_ & ~new_n14320_;
  assign new_n14322_ = ~new_n6212_ & ~new_n14321_;
  assign new_n14323_ = new_n6221_ & ~new_n14318_;
  assign new_n14324_ = ~new_n6221_ & new_n14301_;
  assign new_n14325_ = ~new_n14323_ & ~new_n14324_;
  assign new_n14326_ = new_n6212_ & ~new_n14325_;
  assign new_n14327_ = new_n8075_ & ~new_n14326_;
  assign new_n14328_ = ~new_n14322_ & new_n14327_;
  assign new_n14329_ = new_n8057_ & ~new_n8075_;
  assign new_n14330_ = new_n14223_ & ~new_n14329_;
  assign new_n14331_ = ~new_n14328_ & new_n14330_;
  assign new_n14332_ = ~new_n6238_ & ~new_n14321_;
  assign new_n14333_ = new_n6238_ & ~new_n14325_;
  assign new_n14334_ = new_n8086_ & ~new_n14333_;
  assign new_n14335_ = ~new_n14332_ & new_n14334_;
  assign new_n14336_ = ~new_n14076_ & new_n14214_;
  assign new_n14337_ = ~new_n14335_ & new_n14336_;
  assign new_n14338_ = pi0039 & ~new_n14337_;
  assign new_n14339_ = ~new_n14331_ & new_n14338_;
  assign new_n14340_ = ~new_n14314_ & ~new_n14339_;
  assign new_n14341_ = ~pi0038 & ~new_n14340_;
  assign new_n14342_ = pi0038 & ~new_n14301_;
  assign new_n14343_ = ~pi0100 & ~new_n14342_;
  assign new_n14344_ = ~new_n14341_ & new_n14343_;
  assign new_n14345_ = ~new_n14307_ & ~new_n14344_;
  assign new_n14346_ = ~pi0087 & ~new_n14345_;
  assign new_n14347_ = ~new_n14101_ & ~new_n14288_;
  assign new_n14348_ = ~new_n14281_ & ~new_n14296_;
  assign new_n14349_ = new_n14285_ & ~new_n14348_;
  assign new_n14350_ = ~new_n14347_ & ~new_n14349_;
  assign new_n14351_ = ~new_n14102_ & new_n14278_;
  assign new_n14352_ = ~new_n14350_ & new_n14351_;
  assign new_n14353_ = ~new_n14346_ & ~new_n14352_;
  assign new_n14354_ = ~pi0075 & ~new_n14353_;
  assign new_n14355_ = new_n7500_ & ~new_n14301_;
  assign new_n14356_ = ~new_n14191_ & ~new_n14296_;
  assign new_n14357_ = ~pi0120 & ~new_n14356_;
  assign new_n14358_ = new_n14113_ & ~new_n14357_;
  assign new_n14359_ = ~new_n14355_ & ~new_n14358_;
  assign new_n14360_ = new_n3227_ & ~new_n14359_;
  assign new_n14361_ = ~new_n3227_ & ~new_n14301_;
  assign new_n14362_ = pi0075 & ~new_n14361_;
  assign new_n14363_ = ~new_n14360_ & new_n14362_;
  assign new_n14364_ = new_n7455_ & ~new_n14363_;
  assign new_n14365_ = ~new_n14354_ & new_n14364_;
  assign new_n14366_ = new_n14030_ & ~new_n14365_;
  assign new_n14367_ = ~new_n14295_ & ~new_n14366_;
  assign new_n14368_ = new_n14028_ & ~new_n14172_;
  assign new_n14369_ = new_n14176_ & ~new_n14368_;
  assign new_n14370_ = ~new_n14367_ & new_n14369_;
  assign new_n14371_ = ~pi0039 & ~new_n14231_;
  assign new_n14372_ = new_n7554_ & ~new_n14371_;
  assign new_n14373_ = ~pi0100 & ~new_n14372_;
  assign new_n14374_ = ~new_n7568_ & ~new_n14373_;
  assign new_n14375_ = ~pi0087 & ~new_n14374_;
  assign new_n14376_ = ~new_n7580_ & ~new_n14375_;
  assign new_n14377_ = ~pi0075 & ~new_n14376_;
  assign new_n14378_ = ~new_n7509_ & ~new_n14377_;
  assign new_n14379_ = new_n7733_ & ~new_n14028_;
  assign new_n14380_ = ~new_n14378_ & new_n14379_;
  assign new_n14381_ = new_n7568_ & ~new_n8057_;
  assign new_n14382_ = ~pi0039 & ~new_n14308_;
  assign new_n14383_ = ~new_n8069_ & ~new_n14110_;
  assign new_n14384_ = ~new_n6215_ & ~new_n14383_;
  assign new_n14385_ = new_n6215_ & ~new_n8057_;
  assign new_n14386_ = ~new_n14384_ & ~new_n14385_;
  assign new_n14387_ = ~new_n6238_ & ~new_n14386_;
  assign new_n14388_ = new_n6221_ & ~new_n14383_;
  assign new_n14389_ = ~new_n6221_ & ~new_n8057_;
  assign new_n14390_ = ~new_n14388_ & ~new_n14389_;
  assign new_n14391_ = new_n6238_ & ~new_n14390_;
  assign new_n14392_ = new_n8086_ & ~new_n14391_;
  assign new_n14393_ = ~new_n14387_ & new_n14392_;
  assign new_n14394_ = new_n8057_ & ~new_n8086_;
  assign new_n14395_ = ~pi0299 & ~new_n14394_;
  assign new_n14396_ = ~new_n14393_ & new_n14395_;
  assign new_n14397_ = ~new_n6212_ & ~new_n14386_;
  assign new_n14398_ = new_n6212_ & ~new_n14390_;
  assign new_n14399_ = new_n8075_ & ~new_n14398_;
  assign new_n14400_ = ~new_n14397_ & new_n14399_;
  assign new_n14401_ = pi0299 & ~new_n14329_;
  assign new_n14402_ = ~new_n14400_ & new_n14401_;
  assign new_n14403_ = ~new_n14396_ & ~new_n14402_;
  assign new_n14404_ = pi0039 & ~new_n14403_;
  assign new_n14405_ = ~pi0038 & ~new_n14404_;
  assign new_n14406_ = ~new_n14382_ & new_n14405_;
  assign new_n14407_ = ~pi0100 & ~new_n14090_;
  assign new_n14408_ = ~new_n14406_ & new_n14407_;
  assign new_n14409_ = ~new_n14381_ & ~new_n14408_;
  assign new_n14410_ = ~pi0087 & ~new_n14409_;
  assign new_n14411_ = ~new_n14104_ & ~new_n14410_;
  assign new_n14412_ = ~pi0075 & ~new_n14411_;
  assign new_n14413_ = new_n7501_ & new_n14111_;
  assign new_n14414_ = ~new_n7501_ & new_n8057_;
  assign new_n14415_ = pi0075 & ~new_n14414_;
  assign new_n14416_ = ~new_n14413_ & new_n14415_;
  assign new_n14417_ = ~new_n14412_ & ~new_n14416_;
  assign new_n14418_ = new_n14027_ & ~new_n14417_;
  assign new_n14419_ = ~new_n7455_ & ~new_n14163_;
  assign new_n14420_ = ~new_n14418_ & ~new_n14419_;
  assign new_n14421_ = ~new_n14380_ & new_n14420_;
  assign new_n14422_ = pi0120 & new_n14169_;
  assign new_n14423_ = ~new_n14421_ & new_n14422_;
  assign new_n14424_ = ~new_n14370_ & ~new_n14423_;
  assign new_n14425_ = ~new_n14025_ & ~new_n14424_;
  assign po0278 = new_n14178_ | new_n14425_;
  assign new_n14427_ = new_n2467_ & new_n10153_;
  assign new_n14428_ = ~pi0051 & new_n14427_;
  assign new_n14429_ = new_n6185_ & ~new_n14428_;
  assign new_n14430_ = pi0051 & pi0146;
  assign new_n14431_ = pi0051 & new_n6185_;
  assign new_n14432_ = ~pi0146 & new_n14431_;
  assign new_n14433_ = pi0161 & ~new_n14432_;
  assign new_n14434_ = ~new_n14430_ & ~new_n14433_;
  assign new_n14435_ = new_n14429_ & new_n14434_;
  assign new_n14436_ = ~pi0087 & ~new_n14435_;
  assign new_n14437_ = pi0087 & ~new_n13664_;
  assign new_n14438_ = pi0232 & ~new_n14437_;
  assign new_n14439_ = ~new_n14436_ & new_n14438_;
  assign new_n14440_ = ~pi0134 & ~pi0135;
  assign new_n14441_ = ~pi0136 & new_n14440_;
  assign new_n14442_ = ~pi0130 & new_n14441_;
  assign new_n14443_ = ~pi0132 & new_n14442_;
  assign new_n14444_ = ~pi0126 & new_n14443_;
  assign new_n14445_ = ~pi0121 & new_n14444_;
  assign new_n14446_ = ~pi0125 & ~pi0133;
  assign new_n14447_ = pi0121 & ~new_n14446_;
  assign new_n14448_ = ~pi0121 & new_n14446_;
  assign new_n14449_ = ~new_n14447_ & ~new_n14448_;
  assign new_n14450_ = ~new_n14445_ & ~new_n14449_;
  assign new_n14451_ = ~pi0087 & new_n14428_;
  assign new_n14452_ = ~new_n14450_ & new_n14451_;
  assign new_n14453_ = po1038 & ~new_n14452_;
  assign new_n14454_ = ~new_n14439_ & new_n14453_;
  assign new_n14455_ = pi0299 & ~new_n14435_;
  assign new_n14456_ = ~pi0142 & new_n14431_;
  assign new_n14457_ = pi0144 & ~new_n14456_;
  assign new_n14458_ = pi0051 & pi0142;
  assign new_n14459_ = new_n14429_ & ~new_n14458_;
  assign new_n14460_ = ~new_n14457_ & new_n14459_;
  assign new_n14461_ = ~pi0299 & ~new_n14460_;
  assign new_n14462_ = pi0232 & ~new_n14461_;
  assign new_n14463_ = ~new_n14455_ & new_n14462_;
  assign new_n14464_ = pi0038 & ~new_n14463_;
  assign new_n14465_ = ~pi0100 & ~new_n14464_;
  assign new_n14466_ = pi0038 & ~new_n14428_;
  assign new_n14467_ = ~pi0100 & ~new_n14466_;
  assign new_n14468_ = ~new_n14465_ & ~new_n14467_;
  assign new_n14469_ = new_n2456_ & new_n10152_;
  assign new_n14470_ = new_n13049_ & new_n14469_;
  assign new_n14471_ = ~pi0050 & pi0077;
  assign new_n14472_ = new_n2484_ & new_n14471_;
  assign new_n14473_ = new_n14470_ & new_n14472_;
  assign new_n14474_ = new_n2494_ & new_n7471_;
  assign new_n14475_ = ~pi0024 & pi0314;
  assign new_n14476_ = new_n14474_ & new_n14475_;
  assign new_n14477_ = new_n8899_ & new_n14476_;
  assign new_n14478_ = new_n14473_ & new_n14477_;
  assign new_n14479_ = new_n3098_ & new_n14478_;
  assign new_n14480_ = new_n2579_ & new_n14470_;
  assign new_n14481_ = ~pi0058 & new_n14474_;
  assign new_n14482_ = new_n9044_ & new_n14481_;
  assign new_n14483_ = new_n14480_ & new_n14482_;
  assign new_n14484_ = pi0072 & new_n6379_;
  assign new_n14485_ = new_n14483_ & new_n14484_;
  assign new_n14486_ = new_n14427_ & ~new_n14474_;
  assign new_n14487_ = ~pi0051 & ~new_n14486_;
  assign new_n14488_ = pi0086 & new_n14480_;
  assign new_n14489_ = ~new_n14473_ & ~new_n14488_;
  assign new_n14490_ = new_n11076_ & ~new_n14489_;
  assign new_n14491_ = ~pi0024 & new_n11668_;
  assign new_n14492_ = new_n14480_ & new_n14491_;
  assign new_n14493_ = new_n14427_ & ~new_n14492_;
  assign new_n14494_ = ~new_n14490_ & new_n14493_;
  assign new_n14495_ = new_n14487_ & ~new_n14494_;
  assign new_n14496_ = new_n3098_ & new_n14495_;
  assign new_n14497_ = new_n14428_ & ~new_n14496_;
  assign new_n14498_ = ~new_n14485_ & new_n14497_;
  assign new_n14499_ = ~new_n14479_ & new_n14498_;
  assign new_n14500_ = ~new_n6185_ & ~new_n14499_;
  assign new_n14501_ = pi0072 & new_n10440_;
  assign new_n14502_ = ~new_n14431_ & ~new_n14501_;
  assign new_n14503_ = new_n6185_ & ~new_n14502_;
  assign new_n14504_ = ~new_n14500_ & ~new_n14503_;
  assign new_n14505_ = ~pi0051 & new_n14476_;
  assign new_n14506_ = new_n13439_ & new_n14505_;
  assign new_n14507_ = new_n3098_ & new_n6185_;
  assign new_n14508_ = new_n14506_ & new_n14507_;
  assign new_n14509_ = new_n14504_ & ~new_n14508_;
  assign new_n14510_ = pi0142 & new_n14509_;
  assign new_n14511_ = ~new_n6185_ & new_n14499_;
  assign new_n14512_ = ~pi0072 & ~new_n14506_;
  assign new_n14513_ = new_n6380_ & ~new_n14512_;
  assign new_n14514_ = new_n6185_ & ~new_n14513_;
  assign new_n14515_ = ~new_n14511_ & ~new_n14514_;
  assign new_n14516_ = ~pi0142 & ~new_n14515_;
  assign new_n14517_ = ~pi0144 & ~new_n14516_;
  assign new_n14518_ = ~new_n14510_ & new_n14517_;
  assign new_n14519_ = new_n14428_ & ~new_n14479_;
  assign new_n14520_ = ~new_n14496_ & new_n14519_;
  assign new_n14521_ = ~new_n6185_ & ~new_n14520_;
  assign new_n14522_ = ~new_n14429_ & ~new_n14521_;
  assign new_n14523_ = ~new_n14485_ & new_n14522_;
  assign new_n14524_ = ~new_n14479_ & new_n14523_;
  assign new_n14525_ = new_n14457_ & ~new_n14524_;
  assign new_n14526_ = ~pi0180 & ~new_n14525_;
  assign new_n14527_ = ~new_n14518_ & new_n14526_;
  assign new_n14528_ = pi0144 & ~new_n14523_;
  assign new_n14529_ = ~pi0144 & ~new_n14504_;
  assign new_n14530_ = ~new_n14528_ & ~new_n14529_;
  assign new_n14531_ = ~new_n14456_ & ~new_n14530_;
  assign new_n14532_ = pi0180 & ~new_n14531_;
  assign new_n14533_ = pi0179 & ~new_n14532_;
  assign new_n14534_ = ~new_n14527_ & new_n14533_;
  assign new_n14535_ = ~pi0024 & ~new_n11669_;
  assign new_n14536_ = pi0024 & ~new_n11666_;
  assign new_n14537_ = ~new_n14535_ & ~new_n14536_;
  assign new_n14538_ = ~pi0314 & ~new_n14537_;
  assign new_n14539_ = pi0314 & ~new_n11666_;
  assign new_n14540_ = ~new_n14538_ & ~new_n14539_;
  assign new_n14541_ = new_n2497_ & new_n14540_;
  assign new_n14542_ = ~pi0072 & ~new_n14541_;
  assign new_n14543_ = new_n6380_ & ~new_n14542_;
  assign new_n14544_ = new_n6185_ & ~new_n14543_;
  assign new_n14545_ = ~new_n14511_ & ~new_n14544_;
  assign new_n14546_ = ~pi0142 & ~new_n14545_;
  assign new_n14547_ = new_n7471_ & new_n8960_;
  assign new_n14548_ = new_n14540_ & new_n14547_;
  assign new_n14549_ = ~pi0051 & ~new_n14548_;
  assign new_n14550_ = ~new_n14501_ & new_n14549_;
  assign new_n14551_ = new_n6185_ & ~new_n14550_;
  assign new_n14552_ = ~new_n14500_ & ~new_n14551_;
  assign new_n14553_ = pi0142 & new_n14552_;
  assign new_n14554_ = ~pi0144 & ~new_n14553_;
  assign new_n14555_ = ~new_n14546_ & new_n14554_;
  assign new_n14556_ = new_n14457_ & ~new_n14499_;
  assign new_n14557_ = ~pi0180 & ~new_n14556_;
  assign new_n14558_ = ~new_n14555_ & new_n14557_;
  assign new_n14559_ = new_n2497_ & new_n14537_;
  assign new_n14560_ = ~pi0072 & ~new_n14559_;
  assign new_n14561_ = new_n6380_ & ~new_n14560_;
  assign new_n14562_ = new_n6185_ & ~new_n14561_;
  assign new_n14563_ = ~new_n14511_ & ~new_n14562_;
  assign new_n14564_ = ~pi0142 & ~new_n14563_;
  assign new_n14565_ = new_n14507_ & new_n14559_;
  assign new_n14566_ = ~new_n14503_ & ~new_n14565_;
  assign new_n14567_ = ~new_n14500_ & new_n14566_;
  assign new_n14568_ = pi0142 & new_n14567_;
  assign new_n14569_ = ~pi0144 & ~new_n14568_;
  assign new_n14570_ = ~new_n14564_ & new_n14569_;
  assign new_n14571_ = ~pi0051 & new_n6185_;
  assign new_n14572_ = ~new_n14498_ & new_n14571_;
  assign new_n14573_ = ~new_n14500_ & ~new_n14572_;
  assign new_n14574_ = new_n6185_ & ~new_n14497_;
  assign new_n14575_ = ~pi0142 & ~new_n14574_;
  assign new_n14576_ = ~pi0051 & ~new_n14427_;
  assign new_n14577_ = new_n6185_ & new_n14576_;
  assign new_n14578_ = ~new_n14507_ & ~new_n14577_;
  assign new_n14579_ = new_n3098_ & ~new_n14495_;
  assign new_n14580_ = ~new_n14578_ & ~new_n14579_;
  assign new_n14581_ = pi0142 & ~new_n14580_;
  assign new_n14582_ = ~new_n14575_ & ~new_n14581_;
  assign new_n14583_ = ~new_n14522_ & ~new_n14582_;
  assign new_n14584_ = new_n14573_ & ~new_n14583_;
  assign new_n14585_ = pi0144 & ~new_n14584_;
  assign new_n14586_ = pi0180 & ~new_n14585_;
  assign new_n14587_ = ~new_n14570_ & new_n14586_;
  assign new_n14588_ = ~pi0179 & ~new_n14587_;
  assign new_n14589_ = ~new_n14558_ & new_n14588_;
  assign new_n14590_ = ~new_n14534_ & ~new_n14589_;
  assign new_n14591_ = ~pi0299 & ~new_n14590_;
  assign new_n14592_ = ~pi0161 & ~new_n14432_;
  assign new_n14593_ = ~new_n14504_ & new_n14592_;
  assign new_n14594_ = new_n14427_ & ~new_n14485_;
  assign new_n14595_ = new_n14571_ & ~new_n14594_;
  assign new_n14596_ = ~pi0146 & ~new_n14595_;
  assign new_n14597_ = ~new_n14500_ & new_n14596_;
  assign new_n14598_ = pi0146 & new_n14523_;
  assign new_n14599_ = pi0161 & ~new_n14598_;
  assign new_n14600_ = ~new_n14597_ & new_n14599_;
  assign new_n14601_ = ~new_n14593_ & ~new_n14600_;
  assign new_n14602_ = new_n9361_ & ~new_n14601_;
  assign new_n14603_ = pi0146 & new_n14509_;
  assign new_n14604_ = ~pi0146 & ~new_n14515_;
  assign new_n14605_ = ~pi0161 & ~new_n14604_;
  assign new_n14606_ = ~new_n14603_ & new_n14605_;
  assign new_n14607_ = new_n14571_ & new_n14594_;
  assign new_n14608_ = ~new_n14479_ & new_n14607_;
  assign new_n14609_ = ~new_n14431_ & ~new_n14608_;
  assign new_n14610_ = pi0146 & ~new_n14428_;
  assign new_n14611_ = ~new_n14609_ & ~new_n14610_;
  assign new_n14612_ = pi0161 & ~new_n14611_;
  assign new_n14613_ = ~new_n14511_ & new_n14612_;
  assign new_n14614_ = ~new_n14606_ & ~new_n14613_;
  assign new_n14615_ = new_n9407_ & ~new_n14614_;
  assign new_n14616_ = ~new_n14602_ & ~new_n14615_;
  assign new_n14617_ = pi0156 & ~new_n14616_;
  assign new_n14618_ = pi0146 & new_n14552_;
  assign new_n14619_ = ~pi0146 & ~new_n14545_;
  assign new_n14620_ = new_n9407_ & ~new_n14619_;
  assign new_n14621_ = ~new_n14618_ & new_n14620_;
  assign new_n14622_ = ~pi0146 & ~new_n14563_;
  assign new_n14623_ = pi0146 & new_n14567_;
  assign new_n14624_ = new_n9361_ & ~new_n14623_;
  assign new_n14625_ = ~new_n14622_ & new_n14624_;
  assign new_n14626_ = ~pi0161 & ~new_n14625_;
  assign new_n14627_ = ~new_n14621_ & new_n14626_;
  assign new_n14628_ = ~pi0146 & ~new_n14574_;
  assign new_n14629_ = pi0146 & ~new_n14580_;
  assign new_n14630_ = ~new_n14628_ & ~new_n14629_;
  assign new_n14631_ = ~new_n14522_ & ~new_n14630_;
  assign new_n14632_ = new_n14573_ & ~new_n14631_;
  assign new_n14633_ = new_n9361_ & ~new_n14632_;
  assign new_n14634_ = new_n9407_ & ~new_n14432_;
  assign new_n14635_ = ~new_n14499_ & new_n14634_;
  assign new_n14636_ = pi0161 & ~new_n14635_;
  assign new_n14637_ = ~new_n14633_ & new_n14636_;
  assign new_n14638_ = ~pi0156 & ~new_n14637_;
  assign new_n14639_ = ~new_n14627_ & new_n14638_;
  assign new_n14640_ = ~new_n14617_ & ~new_n14639_;
  assign new_n14641_ = ~new_n14591_ & new_n14640_;
  assign new_n14642_ = new_n9619_ & ~new_n14641_;
  assign new_n14643_ = new_n3098_ & new_n14483_;
  assign new_n14644_ = new_n14428_ & ~new_n14643_;
  assign new_n14645_ = ~new_n14432_ & ~new_n14644_;
  assign new_n14646_ = pi0161 & ~new_n14645_;
  assign new_n14647_ = ~new_n6185_ & ~new_n14644_;
  assign new_n14648_ = new_n2557_ & new_n7476_;
  assign new_n14649_ = ~pi0051 & ~new_n14648_;
  assign new_n14650_ = new_n6185_ & ~new_n14649_;
  assign new_n14651_ = ~new_n14647_ & ~new_n14650_;
  assign new_n14652_ = pi0146 & ~new_n14651_;
  assign new_n14653_ = ~new_n6203_ & ~new_n14647_;
  assign new_n14654_ = ~pi0146 & ~new_n14653_;
  assign new_n14655_ = ~pi0161 & ~new_n14654_;
  assign new_n14656_ = ~new_n14652_ & new_n14655_;
  assign new_n14657_ = ~new_n14646_ & ~new_n14656_;
  assign new_n14658_ = new_n6453_ & ~new_n14657_;
  assign new_n14659_ = ~new_n9069_ & ~new_n14658_;
  assign new_n14660_ = ~pi0287 & new_n6185_;
  assign new_n14661_ = ~pi0051 & new_n14660_;
  assign new_n14662_ = ~new_n14651_ & ~new_n14661_;
  assign new_n14663_ = new_n14592_ & new_n14662_;
  assign new_n14664_ = new_n14643_ & ~new_n14660_;
  assign new_n14665_ = new_n14428_ & ~new_n14664_;
  assign new_n14666_ = new_n14433_ & ~new_n14665_;
  assign new_n14667_ = ~new_n14663_ & ~new_n14666_;
  assign new_n14668_ = pi0216 & ~new_n14667_;
  assign new_n14669_ = ~new_n14659_ & ~new_n14668_;
  assign new_n14670_ = ~new_n14428_ & ~new_n14435_;
  assign new_n14671_ = ~new_n6453_ & ~new_n14670_;
  assign new_n14672_ = new_n9840_ & ~new_n14671_;
  assign new_n14673_ = ~new_n14669_ & new_n14672_;
  assign new_n14674_ = pi0142 & ~new_n14651_;
  assign new_n14675_ = ~pi0142 & ~new_n14653_;
  assign new_n14676_ = new_n6480_ & ~new_n14675_;
  assign new_n14677_ = ~new_n14674_ & new_n14676_;
  assign new_n14678_ = ~new_n9058_ & ~new_n14677_;
  assign new_n14679_ = pi0224 & ~new_n14456_;
  assign new_n14680_ = new_n14662_ & new_n14679_;
  assign new_n14681_ = ~new_n14678_ & ~new_n14680_;
  assign new_n14682_ = ~new_n14428_ & ~new_n14456_;
  assign new_n14683_ = ~new_n6480_ & ~new_n14682_;
  assign new_n14684_ = pi0144 & ~new_n14683_;
  assign new_n14685_ = ~new_n6480_ & new_n14577_;
  assign new_n14686_ = ~new_n14683_ & ~new_n14685_;
  assign new_n14687_ = ~new_n14684_ & new_n14686_;
  assign new_n14688_ = ~new_n14681_ & new_n14687_;
  assign new_n14689_ = ~pi0051 & ~new_n14644_;
  assign new_n14690_ = ~pi0287 & ~new_n14689_;
  assign new_n14691_ = ~new_n14577_ & ~new_n14660_;
  assign new_n14692_ = ~new_n14690_ & ~new_n14691_;
  assign new_n14693_ = ~new_n14459_ & ~new_n14692_;
  assign new_n14694_ = new_n9058_ & ~new_n14693_;
  assign new_n14695_ = new_n14427_ & new_n14694_;
  assign new_n14696_ = pi0051 & ~new_n6185_;
  assign new_n14697_ = ~new_n14689_ & ~new_n14696_;
  assign new_n14698_ = new_n6480_ & ~new_n14458_;
  assign new_n14699_ = new_n14697_ & new_n14698_;
  assign new_n14700_ = new_n14684_ & ~new_n14699_;
  assign new_n14701_ = ~new_n14695_ & new_n14700_;
  assign new_n14702_ = pi0181 & ~new_n14701_;
  assign new_n14703_ = ~new_n14688_ & new_n14702_;
  assign new_n14704_ = ~new_n14677_ & new_n14687_;
  assign new_n14705_ = ~pi0181 & ~new_n14700_;
  assign new_n14706_ = ~new_n14704_ & new_n14705_;
  assign new_n14707_ = ~pi0299 & ~new_n14706_;
  assign new_n14708_ = ~new_n14703_ & new_n14707_;
  assign new_n14709_ = new_n9806_ & ~new_n14671_;
  assign new_n14710_ = ~new_n14658_ & new_n14709_;
  assign new_n14711_ = pi0232 & ~new_n14710_;
  assign new_n14712_ = ~new_n14708_ & new_n14711_;
  assign new_n14713_ = ~new_n14673_ & new_n14712_;
  assign new_n14714_ = ~new_n6605_ & ~new_n7546_;
  assign new_n14715_ = new_n14643_ & ~new_n14714_;
  assign new_n14716_ = ~pi0232 & new_n14428_;
  assign new_n14717_ = ~new_n14715_ & new_n14716_;
  assign new_n14718_ = pi0039 & ~new_n14717_;
  assign new_n14719_ = ~new_n14713_ & new_n14718_;
  assign new_n14720_ = ~pi0039 & ~pi0232;
  assign new_n14721_ = ~new_n14499_ & new_n14720_;
  assign new_n14722_ = ~new_n14719_ & ~new_n14721_;
  assign new_n14723_ = ~new_n14642_ & new_n14722_;
  assign new_n14724_ = ~pi0038 & ~new_n14723_;
  assign new_n14725_ = ~new_n14468_ & ~new_n14724_;
  assign new_n14726_ = pi0100 & new_n14428_;
  assign new_n14727_ = new_n3283_ & ~new_n14726_;
  assign new_n14728_ = pi0100 & new_n14463_;
  assign new_n14729_ = new_n14727_ & ~new_n14728_;
  assign new_n14730_ = ~new_n14725_ & new_n14729_;
  assign new_n14731_ = ~pi0087 & ~new_n3271_;
  assign new_n14732_ = ~new_n14428_ & new_n14731_;
  assign new_n14733_ = ~new_n14463_ & new_n14732_;
  assign new_n14734_ = ~pi0184 & ~pi0299;
  assign new_n14735_ = ~pi0163 & pi0299;
  assign new_n14736_ = ~new_n14734_ & ~new_n14735_;
  assign new_n14737_ = new_n7499_ & new_n14736_;
  assign new_n14738_ = pi0087 & ~new_n14737_;
  assign new_n14739_ = ~new_n14450_ & ~new_n14738_;
  assign new_n14740_ = ~new_n14733_ & new_n14739_;
  assign new_n14741_ = ~new_n14730_ & new_n14740_;
  assign new_n14742_ = new_n6185_ & ~new_n14549_;
  assign new_n14743_ = ~new_n14458_ & new_n14742_;
  assign new_n14744_ = pi0144 & ~new_n14743_;
  assign new_n14745_ = new_n14427_ & ~new_n14478_;
  assign new_n14746_ = new_n14474_ & new_n14745_;
  assign new_n14747_ = new_n14494_ & new_n14746_;
  assign new_n14748_ = new_n14487_ & ~new_n14747_;
  assign new_n14749_ = new_n3098_ & ~new_n14748_;
  assign new_n14750_ = ~new_n14578_ & ~new_n14749_;
  assign new_n14751_ = pi0142 & new_n14750_;
  assign new_n14752_ = new_n6185_ & ~new_n14520_;
  assign new_n14753_ = ~pi0142 & new_n14752_;
  assign new_n14754_ = ~pi0144 & ~new_n14753_;
  assign new_n14755_ = ~new_n14751_ & new_n14754_;
  assign new_n14756_ = pi0180 & ~new_n14755_;
  assign new_n14757_ = ~new_n14744_ & new_n14756_;
  assign new_n14758_ = new_n14457_ & ~new_n14565_;
  assign new_n14759_ = ~pi0144 & ~new_n14582_;
  assign new_n14760_ = ~pi0180 & ~new_n14759_;
  assign new_n14761_ = ~new_n14758_ & new_n14760_;
  assign new_n14762_ = pi0179 & ~new_n14761_;
  assign new_n14763_ = ~new_n14757_ & new_n14762_;
  assign new_n14764_ = new_n14457_ & ~new_n14508_;
  assign new_n14765_ = ~pi0051 & ~new_n14745_;
  assign new_n14766_ = new_n3098_ & ~new_n14765_;
  assign new_n14767_ = ~new_n14578_ & ~new_n14766_;
  assign new_n14768_ = pi0142 & new_n14767_;
  assign new_n14769_ = new_n6185_ & ~new_n14519_;
  assign new_n14770_ = ~pi0142 & new_n14769_;
  assign new_n14771_ = ~pi0144 & ~new_n14770_;
  assign new_n14772_ = ~new_n14768_ & new_n14771_;
  assign new_n14773_ = pi0180 & ~new_n14772_;
  assign new_n14774_ = ~new_n14764_ & new_n14773_;
  assign new_n14775_ = ~pi0180 & new_n14460_;
  assign new_n14776_ = ~pi0179 & ~new_n14775_;
  assign new_n14777_ = ~new_n14774_ & new_n14776_;
  assign new_n14778_ = ~new_n14763_ & ~new_n14777_;
  assign new_n14779_ = ~pi0299 & ~new_n14778_;
  assign new_n14780_ = ~new_n14430_ & new_n14742_;
  assign new_n14781_ = pi0161 & ~new_n14780_;
  assign new_n14782_ = pi0146 & new_n14750_;
  assign new_n14783_ = ~pi0146 & new_n14752_;
  assign new_n14784_ = ~pi0161 & ~new_n14783_;
  assign new_n14785_ = ~new_n14782_ & new_n14784_;
  assign new_n14786_ = ~new_n14781_ & ~new_n14785_;
  assign new_n14787_ = new_n9361_ & ~new_n14786_;
  assign new_n14788_ = new_n14433_ & ~new_n14565_;
  assign new_n14789_ = ~pi0161 & ~new_n14630_;
  assign new_n14790_ = ~new_n14788_ & ~new_n14789_;
  assign new_n14791_ = new_n9407_ & ~new_n14790_;
  assign new_n14792_ = pi0232 & ~new_n14791_;
  assign new_n14793_ = ~new_n14787_ & new_n14792_;
  assign new_n14794_ = pi0156 & ~new_n14793_;
  assign new_n14795_ = ~pi0039 & ~new_n14794_;
  assign new_n14796_ = ~new_n14779_ & new_n14795_;
  assign new_n14797_ = ~pi0142 & ~new_n14648_;
  assign new_n14798_ = new_n9058_ & new_n14660_;
  assign new_n14799_ = pi0142 & ~new_n3100_;
  assign new_n14800_ = new_n14798_ & ~new_n14799_;
  assign new_n14801_ = ~new_n14797_ & new_n14800_;
  assign new_n14802_ = new_n14457_ & ~new_n14801_;
  assign new_n14803_ = ~pi0144 & ~new_n14459_;
  assign new_n14804_ = ~new_n14694_ & new_n14803_;
  assign new_n14805_ = pi0181 & ~new_n14804_;
  assign new_n14806_ = ~new_n14802_ & new_n14805_;
  assign new_n14807_ = ~pi0181 & new_n14460_;
  assign new_n14808_ = ~pi0299 & ~new_n14807_;
  assign new_n14809_ = ~new_n14806_ & new_n14808_;
  assign new_n14810_ = new_n6185_ & new_n6454_;
  assign new_n14811_ = new_n14433_ & ~new_n14810_;
  assign new_n14812_ = new_n14592_ & ~new_n14692_;
  assign new_n14813_ = new_n9069_ & ~new_n14812_;
  assign new_n14814_ = ~new_n14811_ & new_n14813_;
  assign new_n14815_ = ~new_n9069_ & new_n14435_;
  assign new_n14816_ = new_n9840_ & ~new_n14815_;
  assign new_n14817_ = ~new_n14814_ & new_n14816_;
  assign new_n14818_ = ~pi0159 & new_n14455_;
  assign new_n14819_ = new_n10478_ & ~new_n14818_;
  assign new_n14820_ = ~new_n14817_ & new_n14819_;
  assign new_n14821_ = ~new_n14809_ & new_n14820_;
  assign new_n14822_ = ~pi0038 & ~new_n14821_;
  assign new_n14823_ = ~new_n14796_ & new_n14822_;
  assign new_n14824_ = new_n14433_ & ~new_n14508_;
  assign new_n14825_ = pi0146 & new_n14767_;
  assign new_n14826_ = ~pi0146 & new_n14769_;
  assign new_n14827_ = ~pi0161 & ~new_n14826_;
  assign new_n14828_ = ~new_n14825_ & new_n14827_;
  assign new_n14829_ = ~new_n14824_ & ~new_n14828_;
  assign new_n14830_ = new_n9361_ & ~new_n14829_;
  assign new_n14831_ = ~pi0158 & new_n14455_;
  assign new_n14832_ = pi0232 & ~new_n14831_;
  assign new_n14833_ = ~new_n14830_ & new_n14832_;
  assign new_n14834_ = ~pi0156 & new_n3186_;
  assign new_n14835_ = ~new_n14833_ & new_n14834_;
  assign new_n14836_ = new_n14465_ & ~new_n14835_;
  assign new_n14837_ = ~new_n14823_ & new_n14836_;
  assign new_n14838_ = new_n3283_ & ~new_n14728_;
  assign new_n14839_ = ~new_n14837_ & new_n14838_;
  assign new_n14840_ = ~new_n14463_ & new_n14731_;
  assign new_n14841_ = new_n14450_ & ~new_n14738_;
  assign new_n14842_ = ~new_n14840_ & new_n14841_;
  assign new_n14843_ = ~new_n14839_ & new_n14842_;
  assign new_n14844_ = ~po1038 & ~new_n14843_;
  assign new_n14845_ = ~new_n14741_ & new_n14844_;
  assign po0279 = new_n14454_ | new_n14845_;
  assign new_n14847_ = new_n8057_ & new_n8818_;
  assign new_n14848_ = new_n7455_ & new_n14378_;
  assign new_n14849_ = new_n7733_ & ~new_n14848_;
  assign new_n14850_ = new_n7455_ & new_n14417_;
  assign new_n14851_ = new_n14027_ & ~new_n14850_;
  assign new_n14852_ = ~po1038 & ~new_n14851_;
  assign new_n14853_ = ~new_n14849_ & new_n14852_;
  assign po0280 = new_n14847_ | new_n14853_;
  assign new_n14855_ = ~pi0110 & new_n9053_;
  assign new_n14856_ = ~new_n6223_ & new_n6453_;
  assign new_n14857_ = new_n14855_ & new_n14856_;
  assign new_n14858_ = pi0039 & ~new_n14857_;
  assign new_n14859_ = pi0110 & new_n10069_;
  assign new_n14860_ = ~new_n10976_ & new_n14859_;
  assign new_n14861_ = po1057 & new_n14860_;
  assign new_n14862_ = ~pi0039 & ~new_n14861_;
  assign new_n14863_ = po1038 & ~new_n14862_;
  assign new_n14864_ = ~new_n14858_ & new_n14863_;
  assign new_n14865_ = ~pi0038 & new_n3272_;
  assign new_n14866_ = pi0299 & new_n14857_;
  assign new_n14867_ = ~new_n6244_ & new_n7546_;
  assign new_n14868_ = new_n14855_ & new_n14867_;
  assign new_n14869_ = pi0039 & ~new_n14868_;
  assign new_n14870_ = ~new_n14866_ & new_n14869_;
  assign new_n14871_ = ~pi0111 & ~new_n6326_;
  assign new_n14872_ = ~pi0036 & new_n2637_;
  assign new_n14873_ = ~new_n14871_ & new_n14872_;
  assign new_n14874_ = new_n2457_ & ~new_n14873_;
  assign new_n14875_ = ~new_n2602_ & ~new_n2646_;
  assign new_n14876_ = ~new_n14874_ & new_n14875_;
  assign new_n14877_ = ~pi0083 & ~new_n14876_;
  assign new_n14878_ = new_n2604_ & ~new_n14877_;
  assign new_n14879_ = ~pi0071 & ~new_n14878_;
  assign new_n14880_ = new_n6336_ & ~new_n14879_;
  assign new_n14881_ = ~pi0081 & ~new_n14880_;
  assign new_n14882_ = new_n11437_ & ~new_n14881_;
  assign new_n14883_ = ~pi0090 & ~new_n14882_;
  assign new_n14884_ = new_n2496_ & ~new_n14883_;
  assign new_n14885_ = pi0090 & ~new_n10406_;
  assign new_n14886_ = new_n9168_ & ~new_n14885_;
  assign new_n14887_ = new_n14884_ & new_n14886_;
  assign new_n14888_ = pi0072 & new_n2497_;
  assign new_n14889_ = new_n10406_ & new_n14888_;
  assign new_n14890_ = ~new_n14887_ & ~new_n14889_;
  assign new_n14891_ = new_n6379_ & ~new_n14890_;
  assign new_n14892_ = ~pi0110 & ~new_n14891_;
  assign new_n14893_ = new_n13448_ & ~new_n14892_;
  assign new_n14894_ = new_n2706_ & new_n14884_;
  assign new_n14895_ = ~pi0072 & ~new_n14894_;
  assign new_n14896_ = new_n6380_ & ~new_n13448_;
  assign new_n14897_ = ~new_n14895_ & new_n14896_;
  assign new_n14898_ = ~pi0039 & ~new_n14897_;
  assign new_n14899_ = ~new_n14893_ & new_n14898_;
  assign new_n14900_ = ~new_n14870_ & ~new_n14899_;
  assign new_n14901_ = new_n14865_ & ~new_n14900_;
  assign new_n14902_ = pi0110 & new_n13448_;
  assign new_n14903_ = ~pi0039 & ~new_n14902_;
  assign new_n14904_ = ~new_n14870_ & ~new_n14903_;
  assign new_n14905_ = ~new_n14865_ & ~new_n14904_;
  assign new_n14906_ = ~po1038 & ~new_n14905_;
  assign new_n14907_ = ~new_n14901_ & new_n14906_;
  assign po0281 = ~new_n14864_ & ~new_n14907_;
  assign new_n14909_ = ~pi0125 & new_n14445_;
  assign new_n14910_ = pi0125 & pi0133;
  assign new_n14911_ = ~new_n14446_ & ~new_n14910_;
  assign new_n14912_ = ~new_n14909_ & ~new_n14911_;
  assign new_n14913_ = new_n14428_ & ~new_n14912_;
  assign new_n14914_ = pi0172 & new_n14431_;
  assign new_n14915_ = ~pi0152 & new_n14577_;
  assign new_n14916_ = ~new_n14914_ & ~new_n14915_;
  assign new_n14917_ = pi0232 & ~new_n14916_;
  assign new_n14918_ = ~new_n14913_ & ~new_n14917_;
  assign new_n14919_ = ~pi0087 & ~new_n14918_;
  assign new_n14920_ = pi0087 & new_n7499_;
  assign new_n14921_ = pi0162 & new_n14920_;
  assign new_n14922_ = po1038 & ~new_n14921_;
  assign new_n14923_ = ~new_n14919_ & new_n14922_;
  assign new_n14924_ = ~pi0152 & new_n6185_;
  assign new_n14925_ = new_n14501_ & ~new_n14924_;
  assign new_n14926_ = ~pi0152 & new_n14595_;
  assign new_n14927_ = ~pi0197 & ~new_n14926_;
  assign new_n14928_ = ~new_n14925_ & new_n14927_;
  assign new_n14929_ = ~new_n6185_ & new_n14501_;
  assign new_n14930_ = ~new_n14571_ & ~new_n14929_;
  assign new_n14931_ = ~new_n14608_ & ~new_n14930_;
  assign new_n14932_ = ~pi0152 & pi0197;
  assign new_n14933_ = ~new_n14931_ & new_n14932_;
  assign new_n14934_ = ~new_n14928_ & ~new_n14933_;
  assign new_n14935_ = ~new_n14914_ & ~new_n14934_;
  assign new_n14936_ = ~new_n6185_ & ~new_n14501_;
  assign new_n14937_ = ~new_n14514_ & ~new_n14936_;
  assign new_n14938_ = ~pi0172 & new_n14937_;
  assign new_n14939_ = ~new_n14431_ & ~new_n14508_;
  assign new_n14940_ = ~new_n14501_ & new_n14939_;
  assign new_n14941_ = pi0172 & ~new_n14940_;
  assign new_n14942_ = pi0152 & pi0197;
  assign new_n14943_ = ~new_n14941_ & new_n14942_;
  assign new_n14944_ = ~new_n14938_ & new_n14943_;
  assign new_n14945_ = ~new_n14935_ & ~new_n14944_;
  assign new_n14946_ = new_n9875_ & ~new_n14945_;
  assign new_n14947_ = ~new_n14544_ & ~new_n14936_;
  assign new_n14948_ = ~pi0172 & new_n14947_;
  assign new_n14949_ = ~new_n14550_ & ~new_n14936_;
  assign new_n14950_ = pi0172 & new_n14949_;
  assign new_n14951_ = pi0152 & ~new_n14950_;
  assign new_n14952_ = ~new_n14948_ & new_n14951_;
  assign new_n14953_ = new_n6185_ & new_n14499_;
  assign new_n14954_ = ~new_n14930_ & ~new_n14953_;
  assign new_n14955_ = ~pi0152 & ~new_n14914_;
  assign new_n14956_ = ~new_n14954_ & new_n14955_;
  assign new_n14957_ = pi0197 & ~new_n14956_;
  assign new_n14958_ = ~new_n14952_ & new_n14957_;
  assign new_n14959_ = ~new_n14562_ & ~new_n14936_;
  assign new_n14960_ = pi0152 & new_n14959_;
  assign new_n14961_ = ~new_n14572_ & ~new_n14929_;
  assign new_n14962_ = ~pi0152 & ~new_n14961_;
  assign new_n14963_ = ~pi0172 & ~new_n14962_;
  assign new_n14964_ = ~new_n14960_ & new_n14963_;
  assign new_n14965_ = new_n14502_ & ~new_n14565_;
  assign new_n14966_ = pi0152 & ~new_n14965_;
  assign new_n14967_ = new_n14498_ & new_n14607_;
  assign new_n14968_ = ~new_n14936_ & ~new_n14967_;
  assign new_n14969_ = ~pi0152 & new_n14968_;
  assign new_n14970_ = pi0172 & ~new_n14969_;
  assign new_n14971_ = ~new_n14966_ & new_n14970_;
  assign new_n14972_ = ~pi0197 & ~new_n14971_;
  assign new_n14973_ = ~new_n14964_ & new_n14972_;
  assign new_n14974_ = new_n9881_ & ~new_n14973_;
  assign new_n14975_ = ~new_n14958_ & new_n14974_;
  assign new_n14976_ = ~new_n14946_ & ~new_n14975_;
  assign new_n14977_ = pi0299 & ~new_n14976_;
  assign new_n14978_ = pi0145 & new_n14937_;
  assign new_n14979_ = ~pi0145 & new_n14501_;
  assign new_n14980_ = pi0174 & ~new_n14979_;
  assign new_n14981_ = ~new_n14978_ & new_n14980_;
  assign new_n14982_ = pi0145 & new_n14931_;
  assign new_n14983_ = ~new_n14595_ & ~new_n14929_;
  assign new_n14984_ = ~pi0145 & ~new_n14983_;
  assign new_n14985_ = ~pi0174 & ~new_n14984_;
  assign new_n14986_ = ~new_n14982_ & new_n14985_;
  assign new_n14987_ = ~new_n14981_ & ~new_n14986_;
  assign new_n14988_ = ~pi0193 & ~new_n14987_;
  assign new_n14989_ = ~pi0145 & new_n14508_;
  assign new_n14990_ = ~new_n14939_ & ~new_n14989_;
  assign new_n14991_ = ~new_n14501_ & ~new_n14990_;
  assign new_n14992_ = pi0174 & ~new_n14991_;
  assign new_n14993_ = ~new_n14431_ & ~new_n14479_;
  assign new_n14994_ = pi0145 & ~new_n14993_;
  assign new_n14995_ = new_n14607_ & ~new_n14994_;
  assign new_n14996_ = ~pi0174 & ~new_n14995_;
  assign new_n14997_ = ~new_n14936_ & new_n14996_;
  assign new_n14998_ = pi0193 & ~new_n14997_;
  assign new_n14999_ = ~new_n14992_ & new_n14998_;
  assign new_n15000_ = ~new_n14988_ & ~new_n14999_;
  assign new_n15001_ = new_n9859_ & ~new_n15000_;
  assign new_n15002_ = pi0145 & new_n14947_;
  assign new_n15003_ = ~pi0145 & new_n14959_;
  assign new_n15004_ = ~pi0193 & ~new_n15003_;
  assign new_n15005_ = ~new_n15002_ & new_n15004_;
  assign new_n15006_ = pi0145 & new_n14949_;
  assign new_n15007_ = ~pi0145 & ~new_n14965_;
  assign new_n15008_ = pi0193 & ~new_n15007_;
  assign new_n15009_ = ~new_n15006_ & new_n15008_;
  assign new_n15010_ = pi0174 & ~new_n15009_;
  assign new_n15011_ = ~new_n15005_ & new_n15010_;
  assign new_n15012_ = ~pi0193 & ~new_n14961_;
  assign new_n15013_ = pi0193 & new_n14968_;
  assign new_n15014_ = ~pi0145 & ~new_n15013_;
  assign new_n15015_ = ~new_n15012_ & new_n15014_;
  assign new_n15016_ = pi0193 & new_n14431_;
  assign new_n15017_ = pi0145 & ~new_n15016_;
  assign new_n15018_ = ~new_n14954_ & new_n15017_;
  assign new_n15019_ = ~pi0174 & ~new_n15018_;
  assign new_n15020_ = ~new_n15015_ & new_n15019_;
  assign new_n15021_ = new_n9865_ & ~new_n15020_;
  assign new_n15022_ = ~new_n15011_ & new_n15021_;
  assign new_n15023_ = ~new_n15001_ & ~new_n15022_;
  assign new_n15024_ = ~pi0038 & ~new_n15023_;
  assign new_n15025_ = ~new_n14977_ & ~new_n15024_;
  assign new_n15026_ = new_n9619_ & ~new_n15025_;
  assign new_n15027_ = ~pi0299 & ~new_n8086_;
  assign new_n15028_ = pi0299 & ~new_n8075_;
  assign new_n15029_ = ~new_n15027_ & ~new_n15028_;
  assign new_n15030_ = new_n3100_ & new_n15029_;
  assign new_n15031_ = ~pi0232 & ~new_n15030_;
  assign new_n15032_ = pi0039 & ~new_n15031_;
  assign new_n15033_ = new_n14648_ & new_n14660_;
  assign new_n15034_ = ~new_n14431_ & ~new_n15033_;
  assign new_n15035_ = pi0224 & new_n15034_;
  assign new_n15036_ = new_n6480_ & ~new_n15035_;
  assign new_n15037_ = new_n3100_ & ~new_n6185_;
  assign new_n15038_ = ~new_n14650_ & ~new_n15037_;
  assign new_n15039_ = new_n8086_ & new_n15038_;
  assign new_n15040_ = new_n15036_ & ~new_n15039_;
  assign new_n15041_ = ~new_n14431_ & ~new_n15040_;
  assign new_n15042_ = pi0174 & ~new_n15041_;
  assign new_n15043_ = new_n6185_ & ~new_n14644_;
  assign new_n15044_ = ~new_n15037_ & ~new_n15043_;
  assign new_n15045_ = new_n8086_ & new_n15044_;
  assign new_n15046_ = new_n14643_ & new_n14660_;
  assign new_n15047_ = pi0224 & ~new_n15046_;
  assign new_n15048_ = new_n6480_ & ~new_n15047_;
  assign new_n15049_ = ~new_n14429_ & ~new_n15048_;
  assign new_n15050_ = ~new_n15045_ & ~new_n15049_;
  assign new_n15051_ = ~pi0174 & new_n15050_;
  assign new_n15052_ = pi0193 & ~new_n15051_;
  assign new_n15053_ = ~new_n15042_ & new_n15052_;
  assign new_n15054_ = new_n6185_ & new_n14689_;
  assign new_n15055_ = ~new_n15037_ & ~new_n15054_;
  assign new_n15056_ = ~pi0224 & new_n15055_;
  assign new_n15057_ = pi0224 & ~new_n14692_;
  assign new_n15058_ = new_n6480_ & ~new_n15057_;
  assign new_n15059_ = ~new_n15056_ & new_n15058_;
  assign new_n15060_ = ~new_n14685_ & ~new_n15059_;
  assign new_n15061_ = ~pi0174 & ~new_n15060_;
  assign new_n15062_ = ~new_n8086_ & ~new_n14798_;
  assign new_n15063_ = new_n3100_ & ~new_n15062_;
  assign new_n15064_ = pi0174 & new_n15063_;
  assign new_n15065_ = ~pi0193 & ~new_n15064_;
  assign new_n15066_ = ~new_n15061_ & new_n15065_;
  assign new_n15067_ = pi0180 & ~new_n15066_;
  assign new_n15068_ = ~new_n15053_ & new_n15067_;
  assign new_n15069_ = ~new_n8086_ & ~new_n14429_;
  assign new_n15070_ = ~new_n15055_ & ~new_n15069_;
  assign new_n15071_ = ~pi0174 & new_n15070_;
  assign new_n15072_ = new_n3100_ & new_n8086_;
  assign new_n15073_ = pi0174 & new_n15072_;
  assign new_n15074_ = ~new_n15016_ & ~new_n15073_;
  assign new_n15075_ = ~new_n15071_ & new_n15074_;
  assign new_n15076_ = ~pi0180 & ~new_n15075_;
  assign new_n15077_ = ~pi0299 & ~new_n15076_;
  assign new_n15078_ = ~new_n15068_ & new_n15077_;
  assign new_n15079_ = ~new_n8075_ & new_n14916_;
  assign new_n15080_ = ~pi0152 & ~new_n15044_;
  assign new_n15081_ = pi0152 & ~new_n15038_;
  assign new_n15082_ = ~new_n15080_ & ~new_n15081_;
  assign new_n15083_ = pi0051 & ~pi0172;
  assign new_n15084_ = ~new_n15082_ & ~new_n15083_;
  assign new_n15085_ = ~pi0216 & ~new_n15084_;
  assign new_n15086_ = new_n6453_ & new_n15085_;
  assign new_n15087_ = ~new_n15079_ & ~new_n15086_;
  assign new_n15088_ = new_n9407_ & ~new_n15087_;
  assign new_n15089_ = pi0152 & ~new_n14810_;
  assign new_n15090_ = ~pi0152 & ~new_n14692_;
  assign new_n15091_ = ~pi0172 & ~new_n15090_;
  assign new_n15092_ = ~new_n15089_ & new_n15091_;
  assign new_n15093_ = pi0152 & new_n15034_;
  assign new_n15094_ = ~new_n14429_ & ~new_n15046_;
  assign new_n15095_ = ~pi0152 & new_n15094_;
  assign new_n15096_ = pi0172 & ~new_n15095_;
  assign new_n15097_ = ~new_n15093_ & new_n15096_;
  assign new_n15098_ = pi0216 & ~new_n15097_;
  assign new_n15099_ = ~new_n15092_ & new_n15098_;
  assign new_n15100_ = new_n6453_ & ~new_n15099_;
  assign new_n15101_ = ~new_n15085_ & new_n15100_;
  assign new_n15102_ = ~new_n6453_ & ~new_n14916_;
  assign new_n15103_ = new_n9361_ & ~new_n15102_;
  assign new_n15104_ = ~new_n15101_ & new_n15103_;
  assign new_n15105_ = ~new_n15088_ & ~new_n15104_;
  assign new_n15106_ = ~new_n15078_ & new_n15105_;
  assign new_n15107_ = pi0232 & ~new_n15106_;
  assign new_n15108_ = new_n15032_ & ~new_n15107_;
  assign new_n15109_ = ~pi0232 & ~new_n14501_;
  assign new_n15110_ = ~pi0039 & ~new_n15109_;
  assign new_n15111_ = ~pi0038 & ~new_n15110_;
  assign new_n15112_ = ~new_n15108_ & new_n15111_;
  assign new_n15113_ = pi0299 & new_n14916_;
  assign new_n15114_ = ~pi0174 & new_n14577_;
  assign new_n15115_ = ~pi0299 & ~new_n15016_;
  assign new_n15116_ = ~new_n15114_ & new_n15115_;
  assign new_n15117_ = pi0232 & ~new_n15116_;
  assign new_n15118_ = ~new_n15113_ & new_n15117_;
  assign new_n15119_ = pi0038 & ~new_n15118_;
  assign new_n15120_ = ~pi0100 & ~new_n15119_;
  assign new_n15121_ = ~new_n15112_ & new_n15120_;
  assign new_n15122_ = ~new_n15026_ & new_n15121_;
  assign new_n15123_ = pi0100 & new_n15118_;
  assign new_n15124_ = new_n3283_ & ~new_n15123_;
  assign new_n15125_ = ~new_n15122_ & new_n15124_;
  assign new_n15126_ = new_n14731_ & ~new_n15118_;
  assign new_n15127_ = pi0140 & ~pi0299;
  assign new_n15128_ = pi0162 & pi0299;
  assign new_n15129_ = ~new_n15127_ & ~new_n15128_;
  assign new_n15130_ = new_n7499_ & ~new_n15129_;
  assign new_n15131_ = pi0087 & ~new_n15130_;
  assign new_n15132_ = new_n14912_ & ~new_n15131_;
  assign new_n15133_ = ~new_n15126_ & new_n15132_;
  assign new_n15134_ = ~new_n15125_ & new_n15133_;
  assign new_n15135_ = ~pi0145 & ~new_n14521_;
  assign new_n15136_ = ~new_n14742_ & new_n15135_;
  assign new_n15137_ = ~new_n14521_ & ~new_n14565_;
  assign new_n15138_ = pi0145 & new_n15137_;
  assign new_n15139_ = ~pi0051 & new_n15138_;
  assign new_n15140_ = ~pi0174 & ~new_n15139_;
  assign new_n15141_ = ~new_n15136_ & new_n15140_;
  assign new_n15142_ = ~pi0145 & ~new_n14519_;
  assign new_n15143_ = ~new_n6185_ & ~new_n14519_;
  assign new_n15144_ = ~new_n14429_ & ~new_n15143_;
  assign new_n15145_ = ~new_n14496_ & new_n15144_;
  assign new_n15146_ = ~new_n15142_ & new_n15145_;
  assign new_n15147_ = pi0174 & ~new_n15146_;
  assign new_n15148_ = ~pi0193 & ~new_n15147_;
  assign new_n15149_ = ~new_n15141_ & new_n15148_;
  assign new_n15150_ = new_n14507_ & new_n14541_;
  assign new_n15151_ = ~new_n14521_ & ~new_n15150_;
  assign new_n15152_ = ~pi0145 & new_n15151_;
  assign new_n15153_ = ~pi0174 & ~new_n15138_;
  assign new_n15154_ = ~new_n15152_ & new_n15153_;
  assign new_n15155_ = new_n3098_ & new_n15146_;
  assign new_n15156_ = ~new_n14521_ & ~new_n14750_;
  assign new_n15157_ = pi0174 & ~new_n15156_;
  assign new_n15158_ = ~new_n15155_ & new_n15157_;
  assign new_n15159_ = pi0193 & ~new_n15158_;
  assign new_n15160_ = ~new_n15154_ & new_n15159_;
  assign new_n15161_ = new_n9859_ & ~new_n15160_;
  assign new_n15162_ = ~new_n15149_ & new_n15161_;
  assign new_n15163_ = ~new_n14431_ & ~new_n14521_;
  assign new_n15164_ = ~pi0174 & ~new_n14989_;
  assign new_n15165_ = pi0145 & new_n14427_;
  assign new_n15166_ = ~new_n15164_ & ~new_n15165_;
  assign new_n15167_ = new_n15163_ & ~new_n15166_;
  assign new_n15168_ = ~new_n14521_ & ~new_n14769_;
  assign new_n15169_ = pi0174 & new_n15168_;
  assign new_n15170_ = ~new_n15167_ & ~new_n15169_;
  assign new_n15171_ = ~pi0193 & ~new_n15170_;
  assign new_n15172_ = pi0145 & ~new_n14577_;
  assign new_n15173_ = ~pi0145 & pi0174;
  assign new_n15174_ = ~new_n14767_ & new_n15173_;
  assign new_n15175_ = ~new_n15172_ & ~new_n15174_;
  assign new_n15176_ = ~new_n15164_ & new_n15175_;
  assign new_n15177_ = pi0193 & ~new_n14521_;
  assign new_n15178_ = ~new_n15176_ & new_n15177_;
  assign new_n15179_ = new_n9865_ & ~new_n15178_;
  assign new_n15180_ = ~new_n15171_ & new_n15179_;
  assign new_n15181_ = ~new_n15162_ & ~new_n15180_;
  assign new_n15182_ = ~pi0038 & ~new_n15181_;
  assign new_n15183_ = ~pi0152 & ~new_n15151_;
  assign new_n15184_ = pi0152 & ~new_n15156_;
  assign new_n15185_ = pi0172 & ~new_n15184_;
  assign new_n15186_ = ~new_n15183_ & new_n15185_;
  assign new_n15187_ = ~pi0152 & new_n14742_;
  assign new_n15188_ = ~new_n14520_ & ~new_n14924_;
  assign new_n15189_ = ~pi0172 & ~new_n15188_;
  assign new_n15190_ = ~new_n15187_ & new_n15189_;
  assign new_n15191_ = ~new_n15186_ & ~new_n15190_;
  assign new_n15192_ = ~pi0197 & ~new_n15191_;
  assign new_n15193_ = ~pi0152 & ~new_n15137_;
  assign new_n15194_ = ~new_n14521_ & ~new_n14580_;
  assign new_n15195_ = pi0172 & new_n15194_;
  assign new_n15196_ = ~pi0172 & new_n15145_;
  assign new_n15197_ = pi0152 & ~new_n15196_;
  assign new_n15198_ = ~new_n15195_ & new_n15197_;
  assign new_n15199_ = ~pi0172 & new_n14431_;
  assign new_n15200_ = pi0197 & ~new_n15199_;
  assign new_n15201_ = ~new_n15198_ & new_n15200_;
  assign new_n15202_ = ~new_n15193_ & new_n15201_;
  assign new_n15203_ = pi0299 & new_n9875_;
  assign new_n15204_ = ~new_n15202_ & new_n15203_;
  assign new_n15205_ = ~new_n15192_ & new_n15204_;
  assign new_n15206_ = ~new_n14508_ & ~new_n14521_;
  assign new_n15207_ = ~pi0152 & new_n15206_;
  assign new_n15208_ = ~new_n14431_ & new_n15207_;
  assign new_n15209_ = pi0152 & new_n15168_;
  assign new_n15210_ = ~pi0172 & ~new_n15209_;
  assign new_n15211_ = ~new_n15208_ & new_n15210_;
  assign new_n15212_ = ~new_n14521_ & ~new_n14767_;
  assign new_n15213_ = pi0152 & new_n15212_;
  assign new_n15214_ = pi0172 & ~new_n15213_;
  assign new_n15215_ = ~new_n15207_ & new_n15214_;
  assign new_n15216_ = ~pi0197 & ~new_n15215_;
  assign new_n15217_ = ~new_n15211_ & new_n15216_;
  assign new_n15218_ = ~pi0172 & ~new_n14915_;
  assign new_n15219_ = ~new_n14522_ & new_n15218_;
  assign new_n15220_ = pi0152 & new_n14577_;
  assign new_n15221_ = ~new_n14521_ & ~new_n15220_;
  assign new_n15222_ = pi0172 & ~new_n15221_;
  assign new_n15223_ = pi0197 & ~new_n15222_;
  assign new_n15224_ = ~new_n15219_ & new_n15223_;
  assign new_n15225_ = pi0299 & new_n9881_;
  assign new_n15226_ = ~new_n15224_ & new_n15225_;
  assign new_n15227_ = ~new_n15217_ & new_n15226_;
  assign new_n15228_ = ~new_n15205_ & ~new_n15227_;
  assign new_n15229_ = ~new_n15182_ & new_n15228_;
  assign new_n15230_ = new_n9619_ & ~new_n15229_;
  assign new_n15231_ = ~new_n14467_ & ~new_n15120_;
  assign new_n15232_ = ~new_n14428_ & new_n14916_;
  assign new_n15233_ = ~new_n9069_ & ~new_n15232_;
  assign new_n15234_ = ~pi0152 & new_n14653_;
  assign new_n15235_ = pi0152 & new_n14697_;
  assign new_n15236_ = pi0172 & ~new_n15235_;
  assign new_n15237_ = ~new_n15234_ & new_n15236_;
  assign new_n15238_ = ~new_n14644_ & ~new_n14924_;
  assign new_n15239_ = ~pi0152 & new_n14650_;
  assign new_n15240_ = ~new_n15238_ & ~new_n15239_;
  assign new_n15241_ = ~pi0172 & ~new_n15240_;
  assign new_n15242_ = new_n9069_ & ~new_n15241_;
  assign new_n15243_ = ~new_n15237_ & new_n15242_;
  assign new_n15244_ = new_n9407_ & ~new_n15243_;
  assign new_n15245_ = new_n14662_ & new_n14955_;
  assign new_n15246_ = pi0152 & ~new_n14914_;
  assign new_n15247_ = ~new_n14665_ & new_n15246_;
  assign new_n15248_ = new_n9069_ & ~new_n15247_;
  assign new_n15249_ = ~new_n15245_ & new_n15248_;
  assign new_n15250_ = new_n9361_ & ~new_n15249_;
  assign new_n15251_ = ~new_n15244_ & ~new_n15250_;
  assign new_n15252_ = ~new_n15233_ & ~new_n15251_;
  assign new_n15253_ = ~new_n6185_ & ~new_n14427_;
  assign new_n15254_ = ~new_n9058_ & ~new_n15253_;
  assign new_n15255_ = ~new_n14696_ & new_n15254_;
  assign new_n15256_ = new_n9058_ & new_n14653_;
  assign new_n15257_ = ~new_n15255_ & ~new_n15256_;
  assign new_n15258_ = ~pi0174 & ~new_n15257_;
  assign new_n15259_ = new_n9058_ & new_n14643_;
  assign new_n15260_ = new_n14428_ & ~new_n15259_;
  assign new_n15261_ = ~new_n14431_ & ~new_n15260_;
  assign new_n15262_ = pi0174 & ~new_n15261_;
  assign new_n15263_ = ~pi0180 & ~new_n15262_;
  assign new_n15264_ = ~new_n15258_ & new_n15263_;
  assign new_n15265_ = new_n9058_ & ~new_n14647_;
  assign new_n15266_ = ~new_n10548_ & new_n15265_;
  assign new_n15267_ = ~new_n15255_ & ~new_n15266_;
  assign new_n15268_ = ~pi0174 & ~new_n15267_;
  assign new_n15269_ = ~pi0051 & ~new_n14665_;
  assign new_n15270_ = new_n6185_ & ~new_n15269_;
  assign new_n15271_ = ~new_n15260_ & ~new_n15270_;
  assign new_n15272_ = pi0174 & ~new_n15271_;
  assign new_n15273_ = pi0180 & ~new_n15272_;
  assign new_n15274_ = ~new_n15268_ & new_n15273_;
  assign new_n15275_ = pi0193 & ~new_n15274_;
  assign new_n15276_ = ~new_n15264_ & new_n15275_;
  assign new_n15277_ = new_n9058_ & new_n14651_;
  assign new_n15278_ = ~pi0051 & new_n15254_;
  assign new_n15279_ = ~new_n15277_ & ~new_n15278_;
  assign new_n15280_ = pi0180 & new_n14661_;
  assign new_n15281_ = ~pi0174 & ~new_n15280_;
  assign new_n15282_ = new_n15279_ & new_n15281_;
  assign new_n15283_ = pi0180 & new_n14665_;
  assign new_n15284_ = pi0174 & ~new_n15260_;
  assign new_n15285_ = ~new_n15283_ & new_n15284_;
  assign new_n15286_ = ~pi0193 & ~new_n15285_;
  assign new_n15287_ = ~new_n15282_ & new_n15286_;
  assign new_n15288_ = ~pi0299 & ~new_n15287_;
  assign new_n15289_ = ~new_n15276_ & new_n15288_;
  assign new_n15290_ = ~new_n15252_ & ~new_n15289_;
  assign new_n15291_ = pi0232 & ~new_n15290_;
  assign new_n15292_ = ~pi0299 & ~new_n15260_;
  assign new_n15293_ = new_n9069_ & new_n14643_;
  assign new_n15294_ = new_n14428_ & ~new_n15293_;
  assign new_n15295_ = pi0299 & ~new_n15294_;
  assign new_n15296_ = ~new_n15292_ & ~new_n15295_;
  assign new_n15297_ = ~pi0232 & ~new_n15296_;
  assign new_n15298_ = pi0039 & ~new_n15297_;
  assign new_n15299_ = ~new_n15291_ & new_n15298_;
  assign new_n15300_ = ~pi0232 & ~new_n14520_;
  assign new_n15301_ = ~pi0039 & ~new_n15300_;
  assign new_n15302_ = ~pi0038 & ~new_n15301_;
  assign new_n15303_ = ~new_n15299_ & new_n15302_;
  assign new_n15304_ = ~new_n15231_ & ~new_n15303_;
  assign new_n15305_ = ~new_n15230_ & new_n15304_;
  assign new_n15306_ = new_n14727_ & ~new_n15123_;
  assign new_n15307_ = ~new_n15305_ & new_n15306_;
  assign new_n15308_ = new_n14732_ & ~new_n15118_;
  assign new_n15309_ = ~new_n14912_ & ~new_n15131_;
  assign new_n15310_ = ~new_n15308_ & new_n15309_;
  assign new_n15311_ = ~new_n15307_ & new_n15310_;
  assign new_n15312_ = ~po1038 & ~new_n15311_;
  assign new_n15313_ = ~new_n15134_ & new_n15312_;
  assign po0282 = new_n14923_ | new_n15313_;
  assign new_n15315_ = ~pi0189 & new_n14954_;
  assign new_n15316_ = pi0189 & new_n14947_;
  assign new_n15317_ = ~new_n15315_ & ~new_n15316_;
  assign new_n15318_ = pi0178 & ~new_n15317_;
  assign new_n15319_ = pi0189 & ~new_n14937_;
  assign new_n15320_ = ~pi0189 & ~new_n14931_;
  assign new_n15321_ = ~pi0178 & ~new_n15320_;
  assign new_n15322_ = ~new_n15319_ & new_n15321_;
  assign new_n15323_ = ~new_n15318_ & ~new_n15322_;
  assign new_n15324_ = pi0181 & ~new_n15323_;
  assign new_n15325_ = pi0189 & new_n14959_;
  assign new_n15326_ = ~pi0189 & ~new_n14961_;
  assign new_n15327_ = pi0178 & ~new_n15326_;
  assign new_n15328_ = ~new_n15325_ & new_n15327_;
  assign new_n15329_ = ~pi0189 & ~new_n14983_;
  assign new_n15330_ = pi0189 & new_n14501_;
  assign new_n15331_ = ~pi0178 & ~new_n15330_;
  assign new_n15332_ = ~new_n14431_ & new_n15331_;
  assign new_n15333_ = ~new_n15329_ & new_n15332_;
  assign new_n15334_ = ~pi0181 & ~new_n15333_;
  assign new_n15335_ = new_n14983_ & new_n15331_;
  assign new_n15336_ = new_n15334_ & ~new_n15335_;
  assign new_n15337_ = ~new_n15328_ & new_n15336_;
  assign new_n15338_ = new_n11815_ & ~new_n15337_;
  assign new_n15339_ = ~new_n15324_ & new_n15338_;
  assign new_n15340_ = ~pi0153 & new_n14947_;
  assign new_n15341_ = pi0153 & new_n14949_;
  assign new_n15342_ = pi0157 & ~new_n15341_;
  assign new_n15343_ = ~new_n15340_ & new_n15342_;
  assign new_n15344_ = ~pi0153 & new_n14937_;
  assign new_n15345_ = pi0153 & ~new_n14940_;
  assign new_n15346_ = ~pi0157 & ~new_n15345_;
  assign new_n15347_ = ~new_n15344_ & new_n15346_;
  assign new_n15348_ = ~new_n15343_ & ~new_n15347_;
  assign new_n15349_ = pi0166 & ~new_n15348_;
  assign new_n15350_ = ~pi0157 & new_n14931_;
  assign new_n15351_ = pi0157 & new_n14954_;
  assign new_n15352_ = pi0153 & new_n14431_;
  assign new_n15353_ = ~pi0166 & ~new_n15352_;
  assign new_n15354_ = ~new_n15351_ & new_n15353_;
  assign new_n15355_ = ~new_n15350_ & new_n15354_;
  assign new_n15356_ = ~new_n15349_ & ~new_n15355_;
  assign new_n15357_ = new_n9840_ & ~new_n15356_;
  assign new_n15358_ = pi0166 & ~new_n14965_;
  assign new_n15359_ = ~pi0166 & new_n14968_;
  assign new_n15360_ = pi0153 & ~new_n15359_;
  assign new_n15361_ = ~new_n15358_ & new_n15360_;
  assign new_n15362_ = pi0166 & new_n14959_;
  assign new_n15363_ = ~pi0166 & ~new_n14961_;
  assign new_n15364_ = ~pi0153 & ~new_n15363_;
  assign new_n15365_ = ~new_n15362_ & new_n15364_;
  assign new_n15366_ = ~new_n15361_ & ~new_n15365_;
  assign new_n15367_ = pi0157 & ~new_n15366_;
  assign new_n15368_ = ~pi0166 & ~new_n14983_;
  assign new_n15369_ = pi0166 & new_n14501_;
  assign new_n15370_ = ~pi0157 & ~new_n15352_;
  assign new_n15371_ = ~new_n15369_ & new_n15370_;
  assign new_n15372_ = ~new_n15368_ & new_n15371_;
  assign new_n15373_ = ~new_n15367_ & ~new_n15372_;
  assign new_n15374_ = new_n9806_ & ~new_n15373_;
  assign new_n15375_ = ~pi0189 & new_n15163_;
  assign new_n15376_ = new_n14949_ & ~new_n15375_;
  assign new_n15377_ = pi0178 & ~new_n15315_;
  assign new_n15378_ = ~new_n15376_ & new_n15377_;
  assign new_n15379_ = pi0189 & new_n14940_;
  assign new_n15380_ = ~new_n14431_ & new_n15320_;
  assign new_n15381_ = ~new_n15379_ & ~new_n15380_;
  assign new_n15382_ = ~pi0178 & ~new_n15381_;
  assign new_n15383_ = pi0181 & ~new_n15382_;
  assign new_n15384_ = ~new_n15378_ & new_n15383_;
  assign new_n15385_ = pi0189 & ~new_n14965_;
  assign new_n15386_ = ~pi0189 & new_n14968_;
  assign new_n15387_ = pi0178 & ~new_n15386_;
  assign new_n15388_ = ~new_n15385_ & new_n15387_;
  assign new_n15389_ = new_n15334_ & ~new_n15388_;
  assign new_n15390_ = new_n11854_ & ~new_n15389_;
  assign new_n15391_ = ~new_n15384_ & new_n15390_;
  assign new_n15392_ = ~new_n15374_ & ~new_n15391_;
  assign new_n15393_ = ~new_n15357_ & new_n15392_;
  assign new_n15394_ = ~new_n15339_ & new_n15393_;
  assign new_n15395_ = pi0232 & ~new_n15394_;
  assign new_n15396_ = new_n15110_ & ~new_n15395_;
  assign new_n15397_ = ~pi0126 & new_n14448_;
  assign new_n15398_ = pi0126 & ~new_n14448_;
  assign new_n15399_ = ~new_n15397_ & ~new_n15398_;
  assign new_n15400_ = ~new_n14444_ & ~new_n15399_;
  assign new_n15401_ = ~pi0166 & ~new_n15044_;
  assign new_n15402_ = pi0166 & ~new_n15038_;
  assign new_n15403_ = ~new_n15401_ & ~new_n15402_;
  assign new_n15404_ = pi0051 & ~pi0153;
  assign new_n15405_ = ~new_n15403_ & ~new_n15404_;
  assign new_n15406_ = ~pi0216 & ~new_n15405_;
  assign new_n15407_ = pi0166 & ~new_n15034_;
  assign new_n15408_ = ~pi0166 & ~new_n15094_;
  assign new_n15409_ = pi0153 & ~new_n15408_;
  assign new_n15410_ = ~new_n15407_ & new_n15409_;
  assign new_n15411_ = pi0166 & new_n14810_;
  assign new_n15412_ = ~pi0166 & new_n14692_;
  assign new_n15413_ = ~pi0153 & ~new_n15412_;
  assign new_n15414_ = ~new_n15411_ & new_n15413_;
  assign new_n15415_ = pi0160 & ~new_n15414_;
  assign new_n15416_ = ~new_n15410_ & new_n15415_;
  assign new_n15417_ = pi0216 & ~new_n15416_;
  assign new_n15418_ = new_n6453_ & ~new_n15417_;
  assign new_n15419_ = ~new_n15406_ & new_n15418_;
  assign new_n15420_ = ~pi0051 & ~new_n14577_;
  assign new_n15421_ = ~new_n10321_ & ~new_n14427_;
  assign new_n15422_ = ~pi0051 & ~new_n15421_;
  assign new_n15423_ = ~new_n15352_ & ~new_n15422_;
  assign new_n15424_ = ~new_n15420_ & ~new_n15423_;
  assign new_n15425_ = ~pi0160 & pi0216;
  assign new_n15426_ = new_n6453_ & ~new_n15425_;
  assign new_n15427_ = new_n15424_ & ~new_n15426_;
  assign new_n15428_ = pi0299 & ~new_n15427_;
  assign new_n15429_ = ~new_n15419_ & new_n15428_;
  assign new_n15430_ = ~pi0189 & new_n15070_;
  assign new_n15431_ = pi0189 & new_n15072_;
  assign new_n15432_ = ~pi0182 & ~new_n15431_;
  assign new_n15433_ = ~new_n15430_ & new_n15432_;
  assign new_n15434_ = ~new_n14431_ & new_n15433_;
  assign new_n15435_ = pi0189 & ~new_n15041_;
  assign new_n15436_ = ~pi0189 & new_n15050_;
  assign new_n15437_ = pi0182 & ~new_n15436_;
  assign new_n15438_ = ~new_n15435_ & new_n15437_;
  assign new_n15439_ = ~new_n15434_ & ~new_n15438_;
  assign new_n15440_ = new_n11854_ & ~new_n15439_;
  assign new_n15441_ = ~pi0189 & ~new_n15060_;
  assign new_n15442_ = pi0189 & new_n15063_;
  assign new_n15443_ = pi0182 & ~new_n15442_;
  assign new_n15444_ = ~new_n15441_ & new_n15443_;
  assign new_n15445_ = ~new_n15433_ & ~new_n15444_;
  assign new_n15446_ = new_n11815_ & ~new_n15445_;
  assign new_n15447_ = ~new_n15440_ & ~new_n15446_;
  assign new_n15448_ = ~new_n15429_ & new_n15447_;
  assign new_n15449_ = pi0232 & ~new_n15448_;
  assign new_n15450_ = new_n15032_ & ~new_n15449_;
  assign new_n15451_ = new_n15400_ & ~new_n15450_;
  assign new_n15452_ = ~new_n15396_ & new_n15451_;
  assign new_n15453_ = ~pi0166 & ~new_n15151_;
  assign new_n15454_ = pi0166 & ~new_n15156_;
  assign new_n15455_ = pi0153 & ~new_n15454_;
  assign new_n15456_ = ~new_n15453_ & new_n15455_;
  assign new_n15457_ = ~pi0166 & new_n14742_;
  assign new_n15458_ = ~new_n10321_ & ~new_n14520_;
  assign new_n15459_ = ~pi0153 & ~new_n15458_;
  assign new_n15460_ = ~new_n15457_ & new_n15459_;
  assign new_n15461_ = ~new_n15456_ & ~new_n15460_;
  assign new_n15462_ = ~pi0157 & ~new_n15461_;
  assign new_n15463_ = pi0051 & new_n10321_;
  assign new_n15464_ = pi0166 & ~new_n15168_;
  assign new_n15465_ = ~new_n15463_ & ~new_n15464_;
  assign new_n15466_ = ~pi0153 & ~new_n15465_;
  assign new_n15467_ = ~pi0166 & ~new_n15206_;
  assign new_n15468_ = pi0153 & pi0166;
  assign new_n15469_ = ~new_n15212_ & new_n15468_;
  assign new_n15470_ = pi0157 & ~new_n15469_;
  assign new_n15471_ = ~new_n15467_ & new_n15470_;
  assign new_n15472_ = ~new_n15466_ & new_n15471_;
  assign new_n15473_ = new_n9806_ & ~new_n15472_;
  assign new_n15474_ = ~new_n15462_ & new_n15473_;
  assign new_n15475_ = ~new_n10325_ & ~new_n14520_;
  assign new_n15476_ = ~pi0189 & new_n14742_;
  assign new_n15477_ = ~new_n15475_ & ~new_n15476_;
  assign new_n15478_ = ~pi0178 & ~new_n15477_;
  assign new_n15479_ = pi0189 & new_n15168_;
  assign new_n15480_ = pi0178 & ~new_n15375_;
  assign new_n15481_ = ~pi0189 & new_n15206_;
  assign new_n15482_ = pi0178 & ~new_n15481_;
  assign new_n15483_ = ~new_n15480_ & ~new_n15482_;
  assign new_n15484_ = ~new_n15479_ & ~new_n15483_;
  assign new_n15485_ = ~pi0181 & ~new_n15484_;
  assign new_n15486_ = ~new_n15478_ & new_n15485_;
  assign new_n15487_ = ~new_n14565_ & new_n15375_;
  assign new_n15488_ = pi0189 & new_n15145_;
  assign new_n15489_ = ~pi0178 & ~new_n15488_;
  assign new_n15490_ = ~new_n15487_ & new_n15489_;
  assign new_n15491_ = pi0189 & new_n14522_;
  assign new_n15492_ = new_n15480_ & ~new_n15491_;
  assign new_n15493_ = pi0181 & ~new_n15492_;
  assign new_n15494_ = ~new_n15490_ & new_n15493_;
  assign new_n15495_ = new_n11815_ & ~new_n15494_;
  assign new_n15496_ = ~new_n15486_ & new_n15495_;
  assign new_n15497_ = ~pi0189 & new_n15151_;
  assign new_n15498_ = pi0189 & new_n15156_;
  assign new_n15499_ = ~pi0178 & ~new_n15498_;
  assign new_n15500_ = ~new_n15497_ & new_n15499_;
  assign new_n15501_ = pi0189 & new_n15212_;
  assign new_n15502_ = new_n15482_ & ~new_n15501_;
  assign new_n15503_ = ~pi0181 & ~new_n15502_;
  assign new_n15504_ = ~new_n15500_ & new_n15503_;
  assign new_n15505_ = ~pi0189 & ~new_n14565_;
  assign new_n15506_ = pi0189 & ~new_n14580_;
  assign new_n15507_ = ~pi0178 & ~new_n15506_;
  assign new_n15508_ = ~new_n15505_ & new_n15507_;
  assign new_n15509_ = pi0178 & new_n11824_;
  assign new_n15510_ = new_n14576_ & new_n15509_;
  assign new_n15511_ = pi0181 & ~new_n15510_;
  assign new_n15512_ = ~new_n14521_ & new_n15511_;
  assign new_n15513_ = ~new_n15508_ & new_n15512_;
  assign new_n15514_ = new_n11854_ & ~new_n15513_;
  assign new_n15515_ = ~new_n15504_ & new_n15514_;
  assign new_n15516_ = ~pi0166 & ~new_n15137_;
  assign new_n15517_ = pi0166 & ~new_n15145_;
  assign new_n15518_ = ~new_n15463_ & ~new_n15517_;
  assign new_n15519_ = ~pi0153 & ~new_n15518_;
  assign new_n15520_ = ~new_n15194_ & new_n15468_;
  assign new_n15521_ = ~pi0157 & ~new_n15520_;
  assign new_n15522_ = ~new_n15519_ & new_n15521_;
  assign new_n15523_ = ~new_n15516_ & new_n15522_;
  assign new_n15524_ = ~pi0153 & ~new_n15424_;
  assign new_n15525_ = ~new_n14522_ & new_n15524_;
  assign new_n15526_ = pi0166 & new_n14577_;
  assign new_n15527_ = ~new_n14521_ & ~new_n15526_;
  assign new_n15528_ = pi0153 & ~new_n15527_;
  assign new_n15529_ = pi0157 & ~new_n15528_;
  assign new_n15530_ = ~new_n15525_ & new_n15529_;
  assign new_n15531_ = new_n9840_ & ~new_n15530_;
  assign new_n15532_ = ~new_n15523_ & new_n15531_;
  assign new_n15533_ = ~new_n15515_ & ~new_n15532_;
  assign new_n15534_ = ~new_n15496_ & new_n15533_;
  assign new_n15535_ = ~new_n15474_ & new_n15534_;
  assign new_n15536_ = pi0232 & ~new_n15535_;
  assign new_n15537_ = new_n15301_ & ~new_n15536_;
  assign new_n15538_ = ~new_n10321_ & ~new_n14644_;
  assign new_n15539_ = ~pi0166 & new_n14650_;
  assign new_n15540_ = ~new_n15538_ & ~new_n15539_;
  assign new_n15541_ = ~pi0153 & ~new_n15540_;
  assign new_n15542_ = ~pi0166 & new_n14653_;
  assign new_n15543_ = pi0166 & new_n14697_;
  assign new_n15544_ = pi0153 & ~new_n15543_;
  assign new_n15545_ = ~new_n15542_ & new_n15544_;
  assign new_n15546_ = ~new_n15541_ & ~new_n15545_;
  assign new_n15547_ = ~pi0160 & ~new_n15546_;
  assign new_n15548_ = ~pi0166 & new_n14662_;
  assign new_n15549_ = pi0166 & ~new_n14665_;
  assign new_n15550_ = ~new_n15548_ & ~new_n15549_;
  assign new_n15551_ = pi0160 & ~new_n15352_;
  assign new_n15552_ = ~new_n15550_ & new_n15551_;
  assign new_n15553_ = new_n9069_ & ~new_n15552_;
  assign new_n15554_ = ~new_n15547_ & new_n15553_;
  assign new_n15555_ = ~new_n9069_ & ~new_n15423_;
  assign new_n15556_ = pi0299 & ~new_n15555_;
  assign new_n15557_ = ~new_n15554_ & new_n15556_;
  assign new_n15558_ = pi0182 & new_n14665_;
  assign new_n15559_ = pi0189 & ~new_n15260_;
  assign new_n15560_ = ~new_n15558_ & new_n15559_;
  assign new_n15561_ = pi0182 & new_n14661_;
  assign new_n15562_ = ~pi0189 & ~new_n15561_;
  assign new_n15563_ = new_n15279_ & new_n15562_;
  assign new_n15564_ = ~new_n15560_ & ~new_n15563_;
  assign new_n15565_ = new_n11815_ & ~new_n15564_;
  assign new_n15566_ = ~pi0189 & ~new_n15257_;
  assign new_n15567_ = pi0189 & ~new_n15261_;
  assign new_n15568_ = ~pi0182 & ~new_n15567_;
  assign new_n15569_ = ~new_n15566_ & new_n15568_;
  assign new_n15570_ = ~pi0189 & ~new_n15267_;
  assign new_n15571_ = pi0189 & ~new_n15271_;
  assign new_n15572_ = pi0182 & ~new_n15571_;
  assign new_n15573_ = ~new_n15570_ & new_n15572_;
  assign new_n15574_ = ~new_n15569_ & ~new_n15573_;
  assign new_n15575_ = new_n11854_ & ~new_n15574_;
  assign new_n15576_ = ~new_n15565_ & ~new_n15575_;
  assign new_n15577_ = ~new_n15557_ & new_n15576_;
  assign new_n15578_ = pi0232 & ~new_n15577_;
  assign new_n15579_ = new_n15298_ & ~new_n15578_;
  assign new_n15580_ = ~new_n15400_ & ~new_n15579_;
  assign new_n15581_ = ~new_n15537_ & new_n15580_;
  assign new_n15582_ = new_n3211_ & ~new_n15581_;
  assign new_n15583_ = ~new_n15452_ & new_n15582_;
  assign new_n15584_ = pi0299 & ~new_n15424_;
  assign new_n15585_ = ~pi0189 & new_n14577_;
  assign new_n15586_ = pi0175 & new_n14431_;
  assign new_n15587_ = ~pi0299 & ~new_n15586_;
  assign new_n15588_ = ~new_n15585_ & new_n15587_;
  assign new_n15589_ = pi0232 & ~new_n15588_;
  assign new_n15590_ = ~new_n15584_ & new_n15589_;
  assign new_n15591_ = ~new_n3211_ & new_n15590_;
  assign new_n15592_ = ~new_n3211_ & new_n14428_;
  assign new_n15593_ = ~new_n15400_ & new_n15592_;
  assign new_n15594_ = new_n3283_ & ~new_n15593_;
  assign new_n15595_ = ~new_n15591_ & new_n15594_;
  assign new_n15596_ = ~new_n15583_ & new_n15595_;
  assign new_n15597_ = new_n14731_ & ~new_n15590_;
  assign new_n15598_ = ~pi0150 & pi0299;
  assign new_n15599_ = ~pi0185 & ~pi0299;
  assign new_n15600_ = ~new_n15598_ & ~new_n15599_;
  assign new_n15601_ = new_n7499_ & new_n15600_;
  assign new_n15602_ = pi0087 & ~new_n15601_;
  assign new_n15603_ = ~new_n15597_ & ~new_n15602_;
  assign new_n15604_ = new_n14451_ & ~new_n15400_;
  assign new_n15605_ = ~new_n15603_ & ~new_n15604_;
  assign new_n15606_ = ~po1038 & ~new_n15605_;
  assign new_n15607_ = ~new_n15596_ & new_n15606_;
  assign new_n15608_ = pi0232 & ~new_n15420_;
  assign new_n15609_ = new_n15400_ & ~new_n15608_;
  assign new_n15610_ = ~pi0232 & ~new_n14428_;
  assign new_n15611_ = ~new_n15423_ & ~new_n15610_;
  assign new_n15612_ = ~new_n15609_ & new_n15611_;
  assign new_n15613_ = ~pi0087 & ~new_n15612_;
  assign new_n15614_ = pi0087 & ~new_n13830_;
  assign new_n15615_ = po1038 & ~new_n15614_;
  assign new_n15616_ = ~new_n15613_ & new_n15615_;
  assign po0283 = ~new_n15607_ & ~new_n15616_;
  assign new_n15618_ = new_n3285_ & new_n8886_;
  assign new_n15619_ = ~new_n3298_ & ~new_n15618_;
  assign new_n15620_ = pi0129 & new_n6132_;
  assign new_n15621_ = pi0038 & ~new_n15620_;
  assign new_n15622_ = ~new_n2524_ & ~new_n2855_;
  assign new_n15623_ = new_n2597_ & ~new_n2668_;
  assign new_n15624_ = new_n2451_ & ~new_n15623_;
  assign new_n15625_ = new_n2682_ & ~new_n15624_;
  assign new_n15626_ = new_n2594_ & ~new_n15625_;
  assign new_n15627_ = new_n2686_ & ~new_n15626_;
  assign new_n15628_ = new_n2504_ & ~new_n15627_;
  assign new_n15629_ = ~new_n2507_ & ~new_n15628_;
  assign new_n15630_ = ~pi0086 & ~new_n15629_;
  assign new_n15631_ = new_n2592_ & ~new_n15630_;
  assign new_n15632_ = new_n2590_ & ~new_n15631_;
  assign new_n15633_ = ~new_n2585_ & ~new_n15632_;
  assign new_n15634_ = ~pi0108 & ~new_n15633_;
  assign new_n15635_ = new_n2584_ & ~new_n15634_;
  assign new_n15636_ = new_n2698_ & ~new_n15635_;
  assign new_n15637_ = ~new_n2575_ & ~new_n15636_;
  assign new_n15638_ = new_n2574_ & ~new_n15637_;
  assign new_n15639_ = new_n2573_ & ~new_n15638_;
  assign new_n15640_ = ~po0740 & new_n15639_;
  assign new_n15641_ = ~pi0097 & ~new_n15631_;
  assign new_n15642_ = ~new_n2585_ & ~new_n15641_;
  assign new_n15643_ = ~pi0108 & ~new_n15642_;
  assign new_n15644_ = new_n2584_ & ~new_n15643_;
  assign new_n15645_ = new_n2698_ & ~new_n15644_;
  assign new_n15646_ = ~new_n2575_ & ~new_n15645_;
  assign new_n15647_ = new_n2574_ & ~new_n15646_;
  assign new_n15648_ = new_n2573_ & ~new_n15647_;
  assign new_n15649_ = po0740 & new_n15648_;
  assign new_n15650_ = pi0250 & ~new_n7500_;
  assign new_n15651_ = new_n10071_ & new_n15650_;
  assign new_n15652_ = ~new_n15649_ & new_n15651_;
  assign new_n15653_ = ~new_n15640_ & new_n15652_;
  assign new_n15654_ = pi0127 & new_n15639_;
  assign new_n15655_ = ~pi0127 & new_n15648_;
  assign new_n15656_ = ~new_n15651_ & ~new_n15655_;
  assign new_n15657_ = ~new_n15654_ & new_n15656_;
  assign new_n15658_ = ~new_n15653_ & ~new_n15657_;
  assign new_n15659_ = new_n2566_ & ~new_n15658_;
  assign new_n15660_ = new_n2857_ & ~new_n15659_;
  assign new_n15661_ = new_n2547_ & ~new_n15660_;
  assign new_n15662_ = new_n15622_ & ~new_n15661_;
  assign new_n15663_ = ~pi0070 & ~new_n15662_;
  assign new_n15664_ = ~new_n2848_ & ~new_n15663_;
  assign new_n15665_ = ~pi0051 & ~new_n15664_;
  assign new_n15666_ = new_n2559_ & ~new_n15665_;
  assign new_n15667_ = new_n2926_ & ~new_n15666_;
  assign new_n15668_ = ~new_n2555_ & ~new_n15667_;
  assign new_n15669_ = new_n2724_ & ~new_n15668_;
  assign new_n15670_ = new_n3368_ & ~new_n15669_;
  assign new_n15671_ = ~pi0095 & ~new_n15670_;
  assign new_n15672_ = ~pi0039 & pi0129;
  assign new_n15673_ = ~new_n2726_ & new_n15672_;
  assign new_n15674_ = ~new_n15671_ & new_n15673_;
  assign new_n15675_ = pi0039 & new_n8886_;
  assign new_n15676_ = ~pi0038 & ~new_n15675_;
  assign new_n15677_ = ~new_n15674_ & new_n15676_;
  assign new_n15678_ = ~new_n15621_ & ~new_n15677_;
  assign new_n15679_ = new_n3245_ & ~new_n15678_;
  assign new_n15680_ = ~new_n3212_ & ~new_n8965_;
  assign new_n15681_ = new_n8886_ & ~new_n15680_;
  assign new_n15682_ = ~new_n3245_ & ~new_n15681_;
  assign new_n15683_ = ~pi0075 & ~new_n15682_;
  assign new_n15684_ = ~new_n15679_ & new_n15683_;
  assign new_n15685_ = pi0129 & new_n7301_;
  assign new_n15686_ = pi0075 & new_n15685_;
  assign new_n15687_ = ~pi0092 & ~new_n15686_;
  assign new_n15688_ = ~new_n15684_ & new_n15687_;
  assign new_n15689_ = pi0092 & ~pi0129;
  assign new_n15690_ = new_n13654_ & ~new_n15689_;
  assign new_n15691_ = ~new_n15688_ & new_n15690_;
  assign new_n15692_ = pi0054 & new_n3243_;
  assign new_n15693_ = new_n8886_ & new_n15692_;
  assign new_n15694_ = ~pi0074 & ~new_n15693_;
  assign new_n15695_ = ~new_n15691_ & new_n15694_;
  assign new_n15696_ = new_n6554_ & new_n15685_;
  assign new_n15697_ = pi0074 & ~new_n15696_;
  assign new_n15698_ = ~pi0055 & ~new_n15697_;
  assign new_n15699_ = ~new_n15695_ & new_n15698_;
  assign new_n15700_ = pi0055 & new_n3271_;
  assign new_n15701_ = new_n15685_ & new_n15700_;
  assign new_n15702_ = ~new_n15699_ & ~new_n15701_;
  assign new_n15703_ = ~pi0056 & ~new_n15702_;
  assign new_n15704_ = ~new_n11307_ & ~new_n11316_;
  assign new_n15705_ = ~new_n15703_ & new_n15704_;
  assign new_n15706_ = ~new_n15619_ & ~new_n15705_;
  assign new_n15707_ = new_n3436_ & ~new_n15706_;
  assign new_n15708_ = new_n3298_ & new_n15618_;
  assign new_n15709_ = ~new_n3436_ & ~new_n15708_;
  assign new_n15710_ = ~new_n6120_ & ~new_n15709_;
  assign po0284 = ~new_n15707_ & new_n15710_;
  assign new_n15712_ = ~new_n6130_ & ~new_n7347_;
  assign new_n15713_ = ~pi0038 & ~new_n3373_;
  assign new_n15714_ = new_n6134_ & ~new_n15713_;
  assign new_n15715_ = new_n6259_ & ~new_n6280_;
  assign new_n15716_ = ~pi0087 & ~new_n15715_;
  assign new_n15717_ = ~new_n15714_ & new_n15716_;
  assign new_n15718_ = new_n6289_ & ~new_n15717_;
  assign new_n15719_ = new_n8888_ & new_n10410_;
  assign new_n15720_ = ~pi0129 & ~new_n15719_;
  assign new_n15721_ = po0740 & new_n15719_;
  assign new_n15722_ = new_n8967_ & ~new_n15721_;
  assign new_n15723_ = ~new_n15720_ & new_n15722_;
  assign new_n15724_ = new_n3100_ & new_n15723_;
  assign new_n15725_ = new_n6290_ & ~new_n15724_;
  assign new_n15726_ = ~new_n15718_ & new_n15725_;
  assign new_n15727_ = ~new_n7305_ & ~new_n7341_;
  assign new_n15728_ = ~new_n15726_ & new_n15727_;
  assign new_n15729_ = new_n8879_ & ~new_n15728_;
  assign new_n15730_ = new_n15712_ & ~new_n15729_;
  assign new_n15731_ = ~pi0056 & ~new_n15730_;
  assign new_n15732_ = ~new_n6127_ & ~new_n15731_;
  assign new_n15733_ = ~pi0062 & ~new_n15732_;
  assign new_n15734_ = ~new_n6299_ & ~new_n15733_;
  assign new_n15735_ = new_n3436_ & ~new_n15734_;
  assign po0286 = new_n6123_ & ~new_n15735_;
  assign new_n15737_ = ~pi0051 & ~new_n15296_;
  assign new_n15738_ = ~pi0232 & ~new_n15737_;
  assign new_n15739_ = new_n10982_ & ~new_n15738_;
  assign new_n15740_ = ~pi0051 & ~new_n14651_;
  assign new_n15741_ = ~new_n14660_ & new_n15740_;
  assign new_n15742_ = pi0169 & ~new_n15741_;
  assign new_n15743_ = pi0162 & new_n9069_;
  assign new_n15744_ = ~pi0169 & ~new_n15269_;
  assign new_n15745_ = new_n15743_ & ~new_n15744_;
  assign new_n15746_ = ~new_n15742_ & new_n15745_;
  assign new_n15747_ = pi0169 & new_n6185_;
  assign new_n15748_ = ~new_n3100_ & new_n15747_;
  assign new_n15749_ = ~new_n14689_ & ~new_n15747_;
  assign new_n15750_ = ~pi0162 & new_n9069_;
  assign new_n15751_ = ~new_n15749_ & new_n15750_;
  assign new_n15752_ = ~new_n15748_ & new_n15751_;
  assign new_n15753_ = ~new_n9069_ & new_n14576_;
  assign new_n15754_ = ~new_n15747_ & new_n15753_;
  assign new_n15755_ = pi0299 & ~new_n15754_;
  assign new_n15756_ = ~new_n15752_ & new_n15755_;
  assign new_n15757_ = ~new_n15746_ & new_n15756_;
  assign new_n15758_ = ~pi0191 & ~pi0299;
  assign new_n15759_ = ~pi0051 & ~new_n15260_;
  assign new_n15760_ = pi0140 & new_n15270_;
  assign new_n15761_ = new_n15759_ & ~new_n15760_;
  assign new_n15762_ = new_n15758_ & ~new_n15761_;
  assign new_n15763_ = ~pi0051 & new_n15279_;
  assign new_n15764_ = pi0140 & new_n14660_;
  assign new_n15765_ = new_n15763_ & ~new_n15764_;
  assign new_n15766_ = new_n9010_ & ~new_n15765_;
  assign new_n15767_ = ~new_n15762_ & ~new_n15766_;
  assign new_n15768_ = ~new_n15757_ & new_n15767_;
  assign new_n15769_ = pi0232 & ~new_n15768_;
  assign new_n15770_ = new_n15739_ & ~new_n15769_;
  assign new_n15771_ = new_n7499_ & ~new_n9012_;
  assign new_n15772_ = new_n14576_ & ~new_n15771_;
  assign new_n15773_ = ~new_n10982_ & new_n15772_;
  assign new_n15774_ = ~pi0100 & ~new_n15773_;
  assign new_n15775_ = ~new_n15770_ & new_n15774_;
  assign new_n15776_ = ~new_n15420_ & ~new_n15772_;
  assign new_n15777_ = pi0100 & new_n15776_;
  assign new_n15778_ = new_n3283_ & ~new_n15777_;
  assign new_n15779_ = ~new_n14726_ & new_n15778_;
  assign new_n15780_ = ~new_n15775_ & new_n15779_;
  assign new_n15781_ = pi0087 & ~new_n9750_;
  assign new_n15782_ = new_n14731_ & ~new_n15776_;
  assign new_n15783_ = ~new_n15781_ & ~new_n15782_;
  assign new_n15784_ = ~new_n14451_ & ~new_n15783_;
  assign new_n15785_ = ~pi0132 & new_n15397_;
  assign new_n15786_ = pi0130 & ~new_n15785_;
  assign new_n15787_ = ~pi0130 & new_n15785_;
  assign new_n15788_ = ~new_n15786_ & ~new_n15787_;
  assign new_n15789_ = ~new_n14442_ & ~new_n15788_;
  assign new_n15790_ = ~new_n15784_ & ~new_n15789_;
  assign new_n15791_ = ~new_n15780_ & new_n15790_;
  assign new_n15792_ = ~new_n14696_ & new_n15094_;
  assign new_n15793_ = pi0224 & ~new_n15792_;
  assign new_n15794_ = ~new_n6185_ & ~new_n14649_;
  assign new_n15795_ = ~new_n15043_ & ~new_n15794_;
  assign new_n15796_ = ~pi0224 & ~new_n15795_;
  assign new_n15797_ = ~new_n15793_ & ~new_n15796_;
  assign new_n15798_ = new_n6480_ & ~new_n15797_;
  assign new_n15799_ = ~new_n6480_ & ~new_n15420_;
  assign new_n15800_ = ~new_n15798_ & ~new_n15799_;
  assign new_n15801_ = pi0140 & new_n15800_;
  assign new_n15802_ = new_n8086_ & ~new_n15795_;
  assign new_n15803_ = ~new_n8086_ & ~new_n15420_;
  assign new_n15804_ = ~new_n15802_ & ~new_n15803_;
  assign new_n15805_ = ~pi0140 & new_n15804_;
  assign new_n15806_ = new_n9010_ & ~new_n15805_;
  assign new_n15807_ = ~new_n15801_ & new_n15806_;
  assign new_n15808_ = ~new_n14649_ & ~new_n15747_;
  assign new_n15809_ = pi0169 & new_n15043_;
  assign new_n15810_ = ~new_n15808_ & ~new_n15809_;
  assign new_n15811_ = ~pi0216 & ~new_n15810_;
  assign new_n15812_ = ~pi0051 & ~new_n15033_;
  assign new_n15813_ = ~pi0169 & new_n15812_;
  assign new_n15814_ = pi0169 & new_n15792_;
  assign new_n15815_ = pi0162 & pi0216;
  assign new_n15816_ = ~new_n15814_ & new_n15815_;
  assign new_n15817_ = ~new_n15813_ & new_n15816_;
  assign new_n15818_ = ~new_n15811_ & ~new_n15817_;
  assign new_n15819_ = new_n6453_ & ~new_n15818_;
  assign new_n15820_ = pi0169 & new_n14577_;
  assign new_n15821_ = ~pi0051 & ~new_n15820_;
  assign new_n15822_ = ~new_n8075_ & ~new_n15743_;
  assign new_n15823_ = ~new_n15821_ & new_n15822_;
  assign new_n15824_ = ~new_n15819_ & ~new_n15823_;
  assign new_n15825_ = pi0299 & ~new_n15824_;
  assign new_n15826_ = new_n14648_ & new_n15036_;
  assign new_n15827_ = ~pi0051 & ~new_n15826_;
  assign new_n15828_ = pi0140 & new_n15827_;
  assign new_n15829_ = new_n8086_ & new_n14648_;
  assign new_n15830_ = ~pi0051 & ~new_n15829_;
  assign new_n15831_ = ~pi0140 & new_n15830_;
  assign new_n15832_ = new_n15758_ & ~new_n15831_;
  assign new_n15833_ = ~new_n15828_ & new_n15832_;
  assign new_n15834_ = ~new_n15825_ & ~new_n15833_;
  assign new_n15835_ = ~new_n15807_ & new_n15834_;
  assign new_n15836_ = pi0232 & ~new_n15835_;
  assign new_n15837_ = new_n14648_ & new_n15029_;
  assign new_n15838_ = ~pi0051 & ~new_n15837_;
  assign new_n15839_ = ~pi0232 & ~new_n15838_;
  assign new_n15840_ = pi0039 & ~new_n15839_;
  assign new_n15841_ = ~new_n15836_ & new_n15840_;
  assign new_n15842_ = ~pi0232 & ~new_n14550_;
  assign new_n15843_ = ~pi0039 & ~new_n15842_;
  assign new_n15844_ = ~new_n6185_ & new_n14550_;
  assign new_n15845_ = ~new_n14953_ & ~new_n15844_;
  assign new_n15846_ = ~new_n9012_ & ~new_n15845_;
  assign new_n15847_ = new_n9012_ & new_n14550_;
  assign new_n15848_ = pi0232 & ~new_n15847_;
  assign new_n15849_ = ~new_n15846_ & new_n15848_;
  assign new_n15850_ = new_n15843_ & ~new_n15849_;
  assign new_n15851_ = ~new_n15841_ & ~new_n15850_;
  assign new_n15852_ = ~pi0038 & ~new_n15851_;
  assign new_n15853_ = pi0038 & ~new_n15776_;
  assign new_n15854_ = ~pi0100 & ~new_n15853_;
  assign new_n15855_ = ~new_n15852_ & new_n15854_;
  assign new_n15856_ = new_n15778_ & ~new_n15855_;
  assign new_n15857_ = new_n15783_ & new_n15789_;
  assign new_n15858_ = ~new_n15856_ & new_n15857_;
  assign new_n15859_ = ~new_n15791_ & ~new_n15858_;
  assign new_n15860_ = ~po1038 & ~new_n15859_;
  assign new_n15861_ = ~pi0051 & ~pi0087;
  assign new_n15862_ = ~new_n15820_ & new_n15861_;
  assign new_n15863_ = new_n15789_ & new_n15862_;
  assign new_n15864_ = pi0169 & new_n7499_;
  assign new_n15865_ = ~pi0087 & new_n14576_;
  assign new_n15866_ = ~new_n15864_ & new_n15865_;
  assign new_n15867_ = pi0087 & ~new_n9705_;
  assign new_n15868_ = po1038 & ~new_n15867_;
  assign new_n15869_ = ~new_n15866_ & new_n15868_;
  assign new_n15870_ = ~new_n15863_ & new_n15869_;
  assign po0287 = ~new_n15860_ & ~new_n15870_;
  assign new_n15872_ = ~pi0100 & ~new_n14002_;
  assign new_n15873_ = ~pi0087 & ~new_n7334_;
  assign new_n15874_ = ~new_n15872_ & new_n15873_;
  assign new_n15875_ = ~pi0075 & ~new_n15874_;
  assign new_n15876_ = ~new_n7302_ & ~new_n15875_;
  assign new_n15877_ = ~pi0092 & ~new_n15876_;
  assign new_n15878_ = new_n8880_ & new_n13654_;
  assign po0288 = ~new_n15877_ & new_n15878_;
  assign new_n15880_ = pi0051 & ~pi0151;
  assign new_n15881_ = ~new_n13734_ & ~new_n14431_;
  assign new_n15882_ = ~new_n15880_ & ~new_n15881_;
  assign new_n15883_ = new_n14429_ & new_n15882_;
  assign new_n15884_ = pi0232 & new_n15883_;
  assign new_n15885_ = pi0132 & ~new_n15397_;
  assign new_n15886_ = ~new_n15785_ & ~new_n15885_;
  assign new_n15887_ = ~new_n14443_ & ~new_n15886_;
  assign new_n15888_ = new_n14428_ & ~new_n15887_;
  assign new_n15889_ = ~new_n15884_ & ~new_n15888_;
  assign new_n15890_ = ~pi0087 & ~new_n15889_;
  assign new_n15891_ = pi0164 & new_n14920_;
  assign new_n15892_ = po1038 & ~new_n15891_;
  assign new_n15893_ = ~new_n15890_ & new_n15892_;
  assign new_n15894_ = ~pi0190 & ~pi0299;
  assign new_n15895_ = ~new_n6185_ & ~new_n14561_;
  assign new_n15896_ = pi0182 & ~new_n15895_;
  assign new_n15897_ = ~new_n14544_ & new_n15896_;
  assign new_n15898_ = ~pi0182 & new_n14561_;
  assign new_n15899_ = ~pi0173 & ~new_n15898_;
  assign new_n15900_ = ~new_n15897_ & new_n15899_;
  assign new_n15901_ = ~new_n6185_ & new_n14561_;
  assign new_n15902_ = ~new_n14551_ & ~new_n15901_;
  assign new_n15903_ = pi0182 & ~new_n15902_;
  assign new_n15904_ = new_n14566_ & ~new_n15901_;
  assign new_n15905_ = ~pi0182 & ~new_n15904_;
  assign new_n15906_ = pi0173 & ~new_n15905_;
  assign new_n15907_ = ~new_n15903_ & new_n15906_;
  assign new_n15908_ = ~new_n15900_ & ~new_n15907_;
  assign new_n15909_ = new_n15894_ & ~new_n15908_;
  assign new_n15910_ = ~pi0151 & ~new_n14543_;
  assign new_n15911_ = pi0151 & new_n14550_;
  assign new_n15912_ = ~pi0168 & ~new_n15911_;
  assign new_n15913_ = ~new_n15910_ & new_n15912_;
  assign new_n15914_ = pi0168 & ~new_n15880_;
  assign new_n15915_ = ~new_n14499_ & new_n15914_;
  assign new_n15916_ = new_n6185_ & ~new_n15915_;
  assign new_n15917_ = ~new_n15913_ & new_n15916_;
  assign new_n15918_ = pi0160 & ~new_n15895_;
  assign new_n15919_ = ~new_n15917_ & new_n15918_;
  assign new_n15920_ = ~pi0168 & ~new_n15904_;
  assign new_n15921_ = pi0168 & ~new_n14967_;
  assign new_n15922_ = ~new_n15895_ & new_n15921_;
  assign new_n15923_ = pi0151 & ~new_n15922_;
  assign new_n15924_ = ~new_n15920_ & new_n15923_;
  assign new_n15925_ = ~new_n13734_ & new_n14561_;
  assign new_n15926_ = pi0168 & new_n14572_;
  assign new_n15927_ = ~pi0151 & ~new_n15926_;
  assign new_n15928_ = ~new_n15925_ & new_n15927_;
  assign new_n15929_ = ~pi0160 & ~new_n15928_;
  assign new_n15930_ = ~new_n15924_ & new_n15929_;
  assign new_n15931_ = pi0299 & ~new_n15930_;
  assign new_n15932_ = ~new_n15919_ & new_n15931_;
  assign new_n15933_ = pi0190 & ~pi0299;
  assign new_n15934_ = pi0182 & new_n14479_;
  assign new_n15935_ = new_n14498_ & ~new_n15934_;
  assign new_n15936_ = pi0051 & ~pi0173;
  assign new_n15937_ = new_n6185_ & ~new_n15936_;
  assign new_n15938_ = ~new_n15935_ & new_n15937_;
  assign new_n15939_ = new_n15933_ & ~new_n15938_;
  assign new_n15940_ = ~new_n15901_ & new_n15939_;
  assign new_n15941_ = pi0232 & ~new_n15940_;
  assign new_n15942_ = ~new_n15932_ & new_n15941_;
  assign new_n15943_ = ~new_n15909_ & new_n15942_;
  assign new_n15944_ = ~pi0232 & new_n14561_;
  assign new_n15945_ = ~new_n15943_ & ~new_n15944_;
  assign new_n15946_ = ~pi0039 & ~new_n15945_;
  assign new_n15947_ = pi0168 & ~new_n15044_;
  assign new_n15948_ = ~pi0168 & ~new_n15038_;
  assign new_n15949_ = ~new_n15947_ & ~new_n15948_;
  assign new_n15950_ = ~new_n15880_ & ~new_n15949_;
  assign new_n15951_ = ~pi0216 & ~new_n15950_;
  assign new_n15952_ = ~pi0168 & ~new_n15034_;
  assign new_n15953_ = pi0168 & ~new_n15094_;
  assign new_n15954_ = pi0151 & ~new_n15953_;
  assign new_n15955_ = ~new_n15952_ & new_n15954_;
  assign new_n15956_ = ~pi0168 & new_n14810_;
  assign new_n15957_ = pi0168 & new_n14692_;
  assign new_n15958_ = ~pi0151 & ~new_n15957_;
  assign new_n15959_ = ~new_n15956_ & new_n15958_;
  assign new_n15960_ = pi0149 & ~new_n15959_;
  assign new_n15961_ = ~new_n15955_ & new_n15960_;
  assign new_n15962_ = pi0216 & ~new_n15961_;
  assign new_n15963_ = new_n6453_ & ~new_n15962_;
  assign new_n15964_ = ~new_n15951_ & new_n15963_;
  assign new_n15965_ = ~pi0149 & pi0216;
  assign new_n15966_ = new_n6453_ & ~new_n15965_;
  assign new_n15967_ = new_n15883_ & ~new_n15966_;
  assign new_n15968_ = pi0299 & ~new_n15967_;
  assign new_n15969_ = ~new_n15964_ & new_n15968_;
  assign new_n15970_ = pi0183 & ~new_n15060_;
  assign new_n15971_ = ~pi0183 & ~new_n15055_;
  assign new_n15972_ = ~pi0173 & ~new_n15971_;
  assign new_n15973_ = ~new_n15970_ & new_n15972_;
  assign new_n15974_ = ~pi0183 & new_n15069_;
  assign new_n15975_ = ~pi0183 & ~new_n15045_;
  assign new_n15976_ = pi0173 & ~new_n15050_;
  assign new_n15977_ = ~new_n15975_ & new_n15976_;
  assign new_n15978_ = ~new_n15974_ & ~new_n15977_;
  assign new_n15979_ = ~new_n15973_ & new_n15978_;
  assign new_n15980_ = new_n15933_ & ~new_n15979_;
  assign new_n15981_ = pi0183 & new_n15041_;
  assign new_n15982_ = ~pi0183 & ~new_n14431_;
  assign new_n15983_ = ~new_n15072_ & new_n15982_;
  assign new_n15984_ = pi0173 & ~new_n15983_;
  assign new_n15985_ = ~new_n15981_ & new_n15984_;
  assign new_n15986_ = ~pi0183 & ~new_n8086_;
  assign new_n15987_ = ~pi0173 & ~new_n15986_;
  assign new_n15988_ = new_n15063_ & new_n15987_;
  assign new_n15989_ = new_n15894_ & ~new_n15988_;
  assign new_n15990_ = ~new_n15985_ & new_n15989_;
  assign new_n15991_ = ~new_n15980_ & ~new_n15990_;
  assign new_n15992_ = ~new_n15969_ & new_n15991_;
  assign new_n15993_ = pi0232 & ~new_n15992_;
  assign new_n15994_ = new_n15032_ & ~new_n15993_;
  assign new_n15995_ = ~new_n15946_ & ~new_n15994_;
  assign new_n15996_ = new_n3211_ & ~new_n15995_;
  assign new_n15997_ = pi0299 & ~new_n15883_;
  assign new_n15998_ = pi0190 & new_n14577_;
  assign new_n15999_ = pi0173 & new_n14431_;
  assign new_n16000_ = ~pi0299 & ~new_n15999_;
  assign new_n16001_ = ~new_n15998_ & new_n16000_;
  assign new_n16002_ = pi0232 & ~new_n16001_;
  assign new_n16003_ = ~new_n15997_ & new_n16002_;
  assign new_n16004_ = ~new_n3211_ & new_n16003_;
  assign new_n16005_ = new_n3283_ & ~new_n16004_;
  assign new_n16006_ = ~new_n15996_ & new_n16005_;
  assign new_n16007_ = new_n14731_ & ~new_n16003_;
  assign new_n16008_ = pi0087 & ~new_n9020_;
  assign new_n16009_ = new_n15887_ & ~new_n16008_;
  assign new_n16010_ = ~new_n16007_ & new_n16009_;
  assign new_n16011_ = ~new_n16006_ & new_n16010_;
  assign new_n16012_ = ~pi0183 & ~new_n15257_;
  assign new_n16013_ = pi0183 & ~new_n15267_;
  assign new_n16014_ = pi0173 & ~new_n16013_;
  assign new_n16015_ = ~new_n16012_ & new_n16014_;
  assign new_n16016_ = pi0183 & new_n14661_;
  assign new_n16017_ = ~pi0173 & ~new_n16016_;
  assign new_n16018_ = new_n15279_ & new_n16017_;
  assign new_n16019_ = ~new_n16015_ & ~new_n16018_;
  assign new_n16020_ = new_n15933_ & ~new_n16019_;
  assign new_n16021_ = ~new_n14428_ & new_n15997_;
  assign new_n16022_ = ~new_n13130_ & ~new_n16021_;
  assign new_n16023_ = ~new_n15034_ & ~new_n15880_;
  assign new_n16024_ = ~new_n14651_ & ~new_n16023_;
  assign new_n16025_ = pi0168 & ~new_n16024_;
  assign new_n16026_ = ~new_n14665_ & ~new_n15882_;
  assign new_n16027_ = ~pi0168 & ~new_n16026_;
  assign new_n16028_ = pi0149 & ~new_n16027_;
  assign new_n16029_ = ~new_n16025_ & new_n16028_;
  assign new_n16030_ = pi0168 & ~new_n14653_;
  assign new_n16031_ = ~pi0168 & ~new_n14697_;
  assign new_n16032_ = pi0151 & ~new_n16031_;
  assign new_n16033_ = ~new_n16030_ & new_n16032_;
  assign new_n16034_ = pi0168 & new_n14650_;
  assign new_n16035_ = ~new_n13734_ & ~new_n14644_;
  assign new_n16036_ = ~pi0151 & ~new_n16035_;
  assign new_n16037_ = ~new_n16034_ & new_n16036_;
  assign new_n16038_ = ~pi0149 & ~new_n16037_;
  assign new_n16039_ = ~new_n16033_ & new_n16038_;
  assign new_n16040_ = new_n9069_ & ~new_n16039_;
  assign new_n16041_ = ~new_n16029_ & new_n16040_;
  assign new_n16042_ = ~new_n16022_ & ~new_n16041_;
  assign new_n16043_ = pi0183 & new_n14665_;
  assign new_n16044_ = new_n15894_ & ~new_n15999_;
  assign new_n16045_ = ~new_n15260_ & new_n16044_;
  assign new_n16046_ = ~new_n16043_ & new_n16045_;
  assign new_n16047_ = ~new_n16042_ & ~new_n16046_;
  assign new_n16048_ = ~new_n16020_ & new_n16047_;
  assign new_n16049_ = pi0232 & ~new_n16048_;
  assign new_n16050_ = ~new_n15297_ & ~new_n16049_;
  assign new_n16051_ = pi0039 & ~new_n16050_;
  assign new_n16052_ = pi0151 & new_n14767_;
  assign new_n16053_ = ~pi0151 & ~new_n14519_;
  assign new_n16054_ = ~pi0168 & ~new_n16053_;
  assign new_n16055_ = ~new_n16052_ & new_n16054_;
  assign new_n16056_ = ~pi0151 & new_n14431_;
  assign new_n16057_ = pi0168 & ~new_n16056_;
  assign new_n16058_ = ~new_n14508_ & new_n16057_;
  assign new_n16059_ = ~new_n16055_ & ~new_n16058_;
  assign new_n16060_ = ~pi0160 & ~new_n15143_;
  assign new_n16061_ = ~new_n16059_ & new_n16060_;
  assign new_n16062_ = ~pi0151 & ~new_n15883_;
  assign new_n16063_ = ~new_n15144_ & new_n16062_;
  assign new_n16064_ = ~pi0168 & new_n14577_;
  assign new_n16065_ = ~new_n15143_ & ~new_n16064_;
  assign new_n16066_ = pi0151 & ~new_n16065_;
  assign new_n16067_ = pi0160 & ~new_n16066_;
  assign new_n16068_ = ~new_n16063_ & new_n16067_;
  assign new_n16069_ = pi0299 & ~new_n16068_;
  assign new_n16070_ = ~new_n16061_ & new_n16069_;
  assign new_n16071_ = ~pi0182 & new_n14508_;
  assign new_n16072_ = ~new_n15143_ & ~new_n15936_;
  assign new_n16073_ = ~new_n16071_ & new_n16072_;
  assign new_n16074_ = new_n15933_ & ~new_n16073_;
  assign new_n16075_ = pi0182 & new_n15144_;
  assign new_n16076_ = ~new_n14519_ & new_n16044_;
  assign new_n16077_ = ~new_n16075_ & new_n16076_;
  assign new_n16078_ = pi0232 & ~new_n16077_;
  assign new_n16079_ = ~new_n16074_ & new_n16078_;
  assign new_n16080_ = ~new_n16070_ & new_n16079_;
  assign new_n16081_ = ~pi0232 & new_n14519_;
  assign new_n16082_ = ~pi0039 & ~new_n16081_;
  assign new_n16083_ = ~new_n16080_ & new_n16082_;
  assign new_n16084_ = new_n3211_ & ~new_n16083_;
  assign new_n16085_ = ~new_n16051_ & new_n16084_;
  assign new_n16086_ = new_n3283_ & ~new_n15592_;
  assign new_n16087_ = ~new_n16004_ & new_n16086_;
  assign new_n16088_ = ~new_n16085_ & new_n16087_;
  assign new_n16089_ = new_n14732_ & ~new_n16003_;
  assign new_n16090_ = ~new_n15887_ & ~new_n16008_;
  assign new_n16091_ = ~new_n16089_ & new_n16090_;
  assign new_n16092_ = ~new_n16088_ & new_n16091_;
  assign new_n16093_ = ~po1038 & ~new_n16092_;
  assign new_n16094_ = ~new_n16011_ & new_n16093_;
  assign po0289 = new_n15893_ | new_n16094_;
  assign new_n16096_ = ~new_n6185_ & ~new_n14513_;
  assign new_n16097_ = ~new_n14544_ & ~new_n16096_;
  assign new_n16098_ = pi0154 & pi0232;
  assign new_n16099_ = pi0299 & new_n16098_;
  assign new_n16100_ = new_n16097_ & new_n16099_;
  assign new_n16101_ = new_n14513_ & ~new_n16099_;
  assign new_n16102_ = ~pi0039 & ~pi0176;
  assign new_n16103_ = ~new_n16101_ & new_n16102_;
  assign new_n16104_ = ~new_n16100_ & new_n16103_;
  assign new_n16105_ = new_n9468_ & new_n16097_;
  assign new_n16106_ = ~new_n9468_ & new_n14513_;
  assign new_n16107_ = ~pi0039 & pi0176;
  assign new_n16108_ = ~new_n16106_ & new_n16107_;
  assign new_n16109_ = ~new_n16105_ & new_n16108_;
  assign new_n16110_ = pi0197 & new_n14660_;
  assign new_n16111_ = ~new_n5766_ & ~new_n16110_;
  assign new_n16112_ = new_n6605_ & ~new_n16111_;
  assign new_n16113_ = ~pi0145 & ~new_n8086_;
  assign new_n16114_ = ~pi0299 & ~new_n16113_;
  assign new_n16115_ = ~new_n15062_ & new_n16114_;
  assign new_n16116_ = ~new_n16112_ & ~new_n16115_;
  assign new_n16117_ = new_n3100_ & ~new_n16116_;
  assign new_n16118_ = pi0232 & ~new_n16117_;
  assign new_n16119_ = ~new_n15031_ & ~new_n16118_;
  assign new_n16120_ = pi0039 & ~new_n16119_;
  assign new_n16121_ = new_n11382_ & ~new_n16120_;
  assign new_n16122_ = ~new_n16109_ & new_n16121_;
  assign new_n16123_ = ~new_n16104_ & new_n16122_;
  assign new_n16124_ = ~pi0133 & ~new_n14909_;
  assign new_n16125_ = ~pi0087 & new_n16124_;
  assign new_n16126_ = ~new_n16123_ & new_n16125_;
  assign new_n16127_ = pi0145 & new_n14665_;
  assign new_n16128_ = new_n15292_ & ~new_n16127_;
  assign new_n16129_ = new_n15293_ & ~new_n16110_;
  assign new_n16130_ = new_n14428_ & ~new_n16129_;
  assign new_n16131_ = pi0299 & ~new_n16130_;
  assign new_n16132_ = ~new_n16128_ & ~new_n16131_;
  assign new_n16133_ = pi0232 & ~new_n16132_;
  assign new_n16134_ = new_n15298_ & ~new_n16133_;
  assign new_n16135_ = ~new_n9471_ & new_n14496_;
  assign new_n16136_ = ~pi0039 & new_n14428_;
  assign new_n16137_ = ~new_n16135_ & new_n16136_;
  assign new_n16138_ = ~pi0038 & ~new_n16137_;
  assign new_n16139_ = ~new_n16134_ & new_n16138_;
  assign new_n16140_ = new_n14467_ & ~new_n16139_;
  assign new_n16141_ = new_n14727_ & ~new_n16140_;
  assign new_n16142_ = ~new_n14732_ & ~new_n16141_;
  assign new_n16143_ = ~new_n16124_ & ~new_n16142_;
  assign new_n16144_ = ~pi0183 & ~pi0299;
  assign new_n16145_ = ~pi0149 & pi0299;
  assign new_n16146_ = ~new_n16144_ & ~new_n16145_;
  assign new_n16147_ = new_n7499_ & new_n16146_;
  assign new_n16148_ = pi0087 & ~new_n16147_;
  assign new_n16149_ = ~new_n16143_ & ~new_n16148_;
  assign new_n16150_ = ~new_n16126_ & new_n16149_;
  assign new_n16151_ = ~po1038 & ~new_n16150_;
  assign new_n16152_ = new_n14451_ & ~new_n16124_;
  assign new_n16153_ = pi0149 & new_n14920_;
  assign new_n16154_ = po1038 & ~new_n16153_;
  assign new_n16155_ = ~new_n16152_ & new_n16154_;
  assign po0290 = new_n16151_ | new_n16155_;
  assign new_n16157_ = ~pi0136 & new_n15787_;
  assign new_n16158_ = ~pi0135 & new_n16157_;
  assign new_n16159_ = pi0134 & ~new_n16158_;
  assign new_n16160_ = new_n14427_ & ~new_n16159_;
  assign new_n16161_ = po1038 & new_n15861_;
  assign new_n16162_ = pi0171 & new_n6185_;
  assign new_n16163_ = ~new_n14427_ & new_n16162_;
  assign new_n16164_ = pi0232 & new_n16163_;
  assign new_n16165_ = new_n16161_ & ~new_n16164_;
  assign new_n16166_ = ~new_n16160_ & new_n16165_;
  assign new_n16167_ = pi0039 & pi0186;
  assign new_n16168_ = pi0192 & ~pi0299;
  assign new_n16169_ = ~new_n14660_ & new_n15763_;
  assign new_n16170_ = new_n16168_ & ~new_n16169_;
  assign new_n16171_ = ~pi0192 & ~pi0299;
  assign new_n16172_ = ~new_n15270_ & new_n15759_;
  assign new_n16173_ = new_n16171_ & ~new_n16172_;
  assign new_n16174_ = ~new_n16170_ & ~new_n16173_;
  assign new_n16175_ = new_n15753_ & ~new_n16162_;
  assign new_n16176_ = pi0299 & ~new_n16175_;
  assign new_n16177_ = pi0171 & ~new_n15741_;
  assign new_n16178_ = ~pi0171 & ~new_n15269_;
  assign new_n16179_ = new_n9069_ & ~new_n16178_;
  assign new_n16180_ = ~new_n16177_ & new_n16179_;
  assign new_n16181_ = new_n16176_ & ~new_n16180_;
  assign new_n16182_ = new_n16174_ & ~new_n16181_;
  assign new_n16183_ = pi0232 & ~new_n16182_;
  assign new_n16184_ = ~new_n15738_ & ~new_n16183_;
  assign new_n16185_ = new_n16167_ & ~new_n16184_;
  assign new_n16186_ = pi0039 & ~pi0186;
  assign new_n16187_ = ~new_n15763_ & new_n16168_;
  assign new_n16188_ = ~new_n15759_ & new_n16171_;
  assign new_n16189_ = ~new_n16187_ & ~new_n16188_;
  assign new_n16190_ = ~new_n16181_ & new_n16189_;
  assign new_n16191_ = pi0232 & ~new_n16190_;
  assign new_n16192_ = ~new_n15738_ & ~new_n16191_;
  assign new_n16193_ = new_n16186_ & ~new_n16192_;
  assign new_n16194_ = pi0171 & pi0299;
  assign new_n16195_ = ~new_n16168_ & ~new_n16194_;
  assign new_n16196_ = new_n7499_ & ~new_n16195_;
  assign new_n16197_ = new_n14576_ & ~new_n16196_;
  assign new_n16198_ = ~pi0039 & ~new_n16197_;
  assign new_n16199_ = pi0164 & ~new_n16198_;
  assign new_n16200_ = ~new_n16193_ & new_n16199_;
  assign new_n16201_ = ~new_n16185_ & new_n16200_;
  assign new_n16202_ = new_n4226_ & new_n6185_;
  assign new_n16203_ = ~new_n14689_ & ~new_n16162_;
  assign new_n16204_ = new_n9069_ & ~new_n16203_;
  assign new_n16205_ = ~new_n16202_ & new_n16204_;
  assign new_n16206_ = new_n16176_ & ~new_n16205_;
  assign new_n16207_ = new_n16174_ & ~new_n16206_;
  assign new_n16208_ = pi0232 & ~new_n16207_;
  assign new_n16209_ = ~new_n15738_ & ~new_n16208_;
  assign new_n16210_ = new_n16167_ & ~new_n16209_;
  assign new_n16211_ = new_n16189_ & ~new_n16206_;
  assign new_n16212_ = pi0232 & ~new_n16211_;
  assign new_n16213_ = ~new_n15738_ & ~new_n16212_;
  assign new_n16214_ = new_n16186_ & ~new_n16213_;
  assign new_n16215_ = ~pi0164 & ~new_n16198_;
  assign new_n16216_ = ~new_n16214_ & new_n16215_;
  assign new_n16217_ = ~new_n16210_ & new_n16216_;
  assign new_n16218_ = new_n3211_ & ~new_n16217_;
  assign new_n16219_ = ~new_n16201_ & new_n16218_;
  assign new_n16220_ = ~new_n15420_ & ~new_n16197_;
  assign new_n16221_ = ~new_n3211_ & new_n16220_;
  assign new_n16222_ = new_n3283_ & ~new_n16221_;
  assign new_n16223_ = ~new_n15592_ & new_n16222_;
  assign new_n16224_ = ~new_n16219_ & new_n16223_;
  assign new_n16225_ = new_n14731_ & new_n16197_;
  assign new_n16226_ = ~new_n16159_ & ~new_n16225_;
  assign new_n16227_ = ~new_n16224_ & new_n16226_;
  assign new_n16228_ = pi0232 & ~new_n16195_;
  assign new_n16229_ = new_n15845_ & new_n16228_;
  assign new_n16230_ = ~new_n14550_ & ~new_n16228_;
  assign new_n16231_ = ~pi0039 & ~new_n16230_;
  assign new_n16232_ = ~new_n16229_ & new_n16231_;
  assign new_n16233_ = ~pi0051 & ~new_n16163_;
  assign new_n16234_ = ~pi0164 & pi0216;
  assign new_n16235_ = new_n6453_ & ~new_n16234_;
  assign new_n16236_ = ~new_n16233_ & ~new_n16235_;
  assign new_n16237_ = ~new_n14649_ & ~new_n16162_;
  assign new_n16238_ = pi0171 & new_n15043_;
  assign new_n16239_ = ~new_n16237_ & ~new_n16238_;
  assign new_n16240_ = ~pi0216 & ~new_n16239_;
  assign new_n16241_ = ~pi0171 & new_n15812_;
  assign new_n16242_ = pi0171 & new_n15792_;
  assign new_n16243_ = pi0164 & pi0216;
  assign new_n16244_ = ~new_n16242_ & new_n16243_;
  assign new_n16245_ = ~new_n16241_ & new_n16244_;
  assign new_n16246_ = ~new_n16240_ & ~new_n16245_;
  assign new_n16247_ = new_n6453_ & ~new_n16246_;
  assign new_n16248_ = ~new_n16236_ & ~new_n16247_;
  assign new_n16249_ = pi0299 & ~new_n16248_;
  assign new_n16250_ = ~new_n15804_ & new_n16168_;
  assign new_n16251_ = ~new_n15830_ & new_n16171_;
  assign new_n16252_ = ~new_n16167_ & ~new_n16251_;
  assign new_n16253_ = ~new_n16250_ & new_n16252_;
  assign new_n16254_ = ~new_n15800_ & new_n16168_;
  assign new_n16255_ = ~new_n15827_ & new_n16171_;
  assign new_n16256_ = pi0186 & ~new_n16255_;
  assign new_n16257_ = ~new_n16254_ & new_n16256_;
  assign new_n16258_ = ~new_n16253_ & ~new_n16257_;
  assign new_n16259_ = ~new_n16249_ & ~new_n16258_;
  assign new_n16260_ = pi0232 & ~new_n16259_;
  assign new_n16261_ = new_n15840_ & ~new_n16260_;
  assign new_n16262_ = new_n3211_ & ~new_n16261_;
  assign new_n16263_ = ~new_n16232_ & new_n16262_;
  assign new_n16264_ = new_n16222_ & ~new_n16263_;
  assign new_n16265_ = new_n14731_ & ~new_n16220_;
  assign new_n16266_ = new_n16159_ & ~new_n16265_;
  assign new_n16267_ = ~new_n16264_ & new_n16266_;
  assign new_n16268_ = ~po1038 & ~new_n16267_;
  assign new_n16269_ = ~new_n16227_ & new_n16268_;
  assign po0291 = new_n16166_ | new_n16269_;
  assign new_n16271_ = pi0170 & new_n6185_;
  assign new_n16272_ = new_n10667_ & new_n16271_;
  assign new_n16273_ = new_n14576_ & ~new_n16272_;
  assign new_n16274_ = pi0194 & new_n9031_;
  assign new_n16275_ = new_n16273_ & ~new_n16274_;
  assign new_n16276_ = ~new_n15420_ & ~new_n16275_;
  assign new_n16277_ = pi0100 & new_n16276_;
  assign new_n16278_ = new_n3283_ & ~new_n16277_;
  assign new_n16279_ = ~new_n14649_ & ~new_n16271_;
  assign new_n16280_ = pi0170 & new_n15043_;
  assign new_n16281_ = new_n8075_ & ~new_n16280_;
  assign new_n16282_ = ~new_n16279_ & new_n16281_;
  assign new_n16283_ = ~new_n9069_ & ~new_n16282_;
  assign new_n16284_ = ~pi0170 & new_n15812_;
  assign new_n16285_ = pi0170 & new_n15792_;
  assign new_n16286_ = pi0216 & ~new_n16285_;
  assign new_n16287_ = ~new_n16284_ & new_n16286_;
  assign new_n16288_ = ~new_n16283_ & ~new_n16287_;
  assign new_n16289_ = pi0150 & pi0299;
  assign new_n16290_ = ~new_n14427_ & new_n16271_;
  assign new_n16291_ = ~pi0051 & ~new_n16290_;
  assign new_n16292_ = ~new_n6453_ & new_n16291_;
  assign new_n16293_ = new_n16289_ & ~new_n16292_;
  assign new_n16294_ = ~new_n16288_ & new_n16293_;
  assign new_n16295_ = ~new_n8075_ & new_n16291_;
  assign new_n16296_ = new_n15598_ & ~new_n16295_;
  assign new_n16297_ = ~new_n16282_ & new_n16296_;
  assign new_n16298_ = ~new_n16294_ & ~new_n16297_;
  assign new_n16299_ = pi0185 & new_n15827_;
  assign new_n16300_ = ~pi0185 & new_n15830_;
  assign new_n16301_ = ~pi0299 & ~new_n16300_;
  assign new_n16302_ = ~new_n16299_ & new_n16301_;
  assign new_n16303_ = new_n16298_ & ~new_n16302_;
  assign new_n16304_ = pi0232 & ~new_n16303_;
  assign new_n16305_ = new_n15840_ & ~new_n16304_;
  assign new_n16306_ = ~pi0299 & ~new_n14550_;
  assign new_n16307_ = pi0170 & ~new_n15845_;
  assign new_n16308_ = ~pi0170 & new_n14550_;
  assign new_n16309_ = new_n10667_ & ~new_n16308_;
  assign new_n16310_ = ~new_n16307_ & new_n16309_;
  assign new_n16311_ = new_n15843_ & ~new_n16310_;
  assign new_n16312_ = ~new_n16306_ & new_n16311_;
  assign new_n16313_ = ~new_n16305_ & ~new_n16312_;
  assign new_n16314_ = ~pi0038 & ~new_n16313_;
  assign new_n16315_ = ~new_n15420_ & ~new_n16273_;
  assign new_n16316_ = pi0038 & ~new_n16315_;
  assign new_n16317_ = ~pi0194 & ~new_n16316_;
  assign new_n16318_ = ~new_n16314_ & new_n16317_;
  assign new_n16319_ = pi0185 & new_n15800_;
  assign new_n16320_ = ~pi0185 & new_n15804_;
  assign new_n16321_ = ~pi0299 & ~new_n16320_;
  assign new_n16322_ = ~new_n16319_ & new_n16321_;
  assign new_n16323_ = new_n16298_ & ~new_n16322_;
  assign new_n16324_ = pi0232 & ~new_n16323_;
  assign new_n16325_ = new_n15840_ & ~new_n16324_;
  assign new_n16326_ = new_n10662_ & new_n15845_;
  assign new_n16327_ = new_n16311_ & ~new_n16326_;
  assign new_n16328_ = ~new_n16325_ & ~new_n16327_;
  assign new_n16329_ = ~pi0038 & ~new_n16328_;
  assign new_n16330_ = pi0170 & new_n7499_;
  assign new_n16331_ = ~new_n9031_ & ~new_n16330_;
  assign new_n16332_ = new_n14576_ & new_n16331_;
  assign new_n16333_ = ~new_n15420_ & ~new_n16332_;
  assign new_n16334_ = pi0038 & ~new_n16333_;
  assign new_n16335_ = pi0194 & ~new_n16334_;
  assign new_n16336_ = ~new_n16329_ & new_n16335_;
  assign new_n16337_ = ~new_n16318_ & ~new_n16336_;
  assign new_n16338_ = ~pi0100 & ~new_n16337_;
  assign new_n16339_ = new_n16278_ & ~new_n16338_;
  assign new_n16340_ = pi0135 & ~new_n16157_;
  assign new_n16341_ = pi0134 & new_n16158_;
  assign new_n16342_ = ~new_n16340_ & ~new_n16341_;
  assign new_n16343_ = new_n14731_ & ~new_n16276_;
  assign new_n16344_ = ~new_n16342_ & ~new_n16343_;
  assign new_n16345_ = ~new_n16339_ & new_n16344_;
  assign new_n16346_ = pi0185 & new_n15270_;
  assign new_n16347_ = new_n15759_ & ~new_n16346_;
  assign new_n16348_ = ~new_n10982_ & new_n16273_;
  assign new_n16349_ = ~pi0194 & ~new_n16348_;
  assign new_n16350_ = ~new_n16347_ & new_n16349_;
  assign new_n16351_ = ~pi0185 & new_n15763_;
  assign new_n16352_ = ~new_n10982_ & new_n16332_;
  assign new_n16353_ = pi0194 & ~new_n16352_;
  assign new_n16354_ = ~new_n16169_ & new_n16353_;
  assign new_n16355_ = ~new_n16351_ & new_n16354_;
  assign new_n16356_ = ~new_n16350_ & ~new_n16355_;
  assign new_n16357_ = ~pi0299 & ~new_n16356_;
  assign new_n16358_ = pi0170 & ~new_n15741_;
  assign new_n16359_ = ~pi0170 & ~new_n15269_;
  assign new_n16360_ = new_n9069_ & ~new_n16359_;
  assign new_n16361_ = ~new_n16358_ & new_n16360_;
  assign new_n16362_ = new_n16289_ & ~new_n16361_;
  assign new_n16363_ = new_n4449_ & new_n6185_;
  assign new_n16364_ = ~new_n14689_ & ~new_n16271_;
  assign new_n16365_ = new_n9069_ & ~new_n16364_;
  assign new_n16366_ = ~new_n16363_ & new_n16365_;
  assign new_n16367_ = new_n15598_ & ~new_n16366_;
  assign new_n16368_ = ~new_n16362_ & ~new_n16367_;
  assign new_n16369_ = new_n15753_ & ~new_n16271_;
  assign new_n16370_ = ~new_n16349_ & ~new_n16353_;
  assign new_n16371_ = ~new_n16369_ & ~new_n16370_;
  assign new_n16372_ = ~new_n16368_ & new_n16371_;
  assign new_n16373_ = ~new_n16357_ & ~new_n16372_;
  assign new_n16374_ = pi0232 & ~new_n16373_;
  assign new_n16375_ = ~new_n15739_ & ~new_n16370_;
  assign new_n16376_ = ~new_n16374_ & ~new_n16375_;
  assign new_n16377_ = ~pi0100 & ~new_n16376_;
  assign new_n16378_ = ~new_n14726_ & new_n16278_;
  assign new_n16379_ = ~new_n16377_ & new_n16378_;
  assign new_n16380_ = new_n14731_ & new_n16275_;
  assign new_n16381_ = new_n16342_ & ~new_n16380_;
  assign new_n16382_ = ~new_n16379_ & new_n16381_;
  assign new_n16383_ = ~po1038 & ~new_n16382_;
  assign new_n16384_ = ~new_n16345_ & new_n16383_;
  assign new_n16385_ = new_n14427_ & new_n16342_;
  assign new_n16386_ = ~new_n14427_ & new_n16330_;
  assign new_n16387_ = new_n16161_ & ~new_n16386_;
  assign new_n16388_ = ~new_n16385_ & new_n16387_;
  assign po0292 = new_n16384_ | new_n16388_;
  assign new_n16390_ = pi0136 & ~new_n15787_;
  assign new_n16391_ = ~new_n16157_ & ~new_n16390_;
  assign new_n16392_ = ~new_n14441_ & ~new_n16391_;
  assign new_n16393_ = ~new_n14576_ & new_n16392_;
  assign new_n16394_ = pi0148 & new_n7499_;
  assign new_n16395_ = ~new_n14427_ & ~new_n16394_;
  assign new_n16396_ = ~new_n16393_ & ~new_n16395_;
  assign new_n16397_ = new_n16161_ & ~new_n16396_;
  assign new_n16398_ = ~new_n9741_ & ~new_n15845_;
  assign new_n16399_ = new_n9741_ & new_n14550_;
  assign new_n16400_ = pi0232 & ~new_n16399_;
  assign new_n16401_ = ~new_n16398_ & new_n16400_;
  assign new_n16402_ = new_n15843_ & ~new_n16401_;
  assign new_n16403_ = pi0184 & new_n15800_;
  assign new_n16404_ = ~pi0184 & new_n15804_;
  assign new_n16405_ = new_n9739_ & ~new_n16404_;
  assign new_n16406_ = ~new_n16403_ & new_n16405_;
  assign new_n16407_ = pi0184 & new_n15827_;
  assign new_n16408_ = ~pi0141 & ~pi0299;
  assign new_n16409_ = ~pi0184 & new_n15830_;
  assign new_n16410_ = new_n16408_ & ~new_n16409_;
  assign new_n16411_ = ~new_n16407_ & new_n16410_;
  assign new_n16412_ = new_n8075_ & ~new_n15795_;
  assign new_n16413_ = pi0163 & new_n6453_;
  assign new_n16414_ = new_n15792_ & new_n16413_;
  assign new_n16415_ = ~new_n6453_ & new_n15420_;
  assign new_n16416_ = ~new_n8075_ & ~new_n15420_;
  assign new_n16417_ = ~pi0163 & ~new_n16416_;
  assign new_n16418_ = ~new_n16415_ & ~new_n16417_;
  assign new_n16419_ = ~new_n16414_ & new_n16418_;
  assign new_n16420_ = pi0148 & ~new_n16419_;
  assign new_n16421_ = ~new_n16412_ & new_n16420_;
  assign new_n16422_ = ~pi0287 & new_n13664_;
  assign new_n16423_ = pi0216 & ~new_n16422_;
  assign new_n16424_ = new_n6453_ & ~new_n16423_;
  assign new_n16425_ = new_n14648_ & new_n16424_;
  assign new_n16426_ = ~pi0051 & ~pi0148;
  assign new_n16427_ = ~new_n16425_ & new_n16426_;
  assign new_n16428_ = pi0299 & ~new_n16427_;
  assign new_n16429_ = ~new_n16421_ & new_n16428_;
  assign new_n16430_ = ~new_n16411_ & ~new_n16429_;
  assign new_n16431_ = ~new_n16406_ & new_n16430_;
  assign new_n16432_ = pi0232 & ~new_n16431_;
  assign new_n16433_ = new_n15840_ & ~new_n16432_;
  assign new_n16434_ = new_n3211_ & ~new_n16433_;
  assign new_n16435_ = ~new_n16402_ & new_n16434_;
  assign new_n16436_ = new_n9742_ & ~new_n14427_;
  assign new_n16437_ = ~pi0051 & ~new_n16436_;
  assign new_n16438_ = ~new_n3211_ & ~new_n16437_;
  assign new_n16439_ = new_n3283_ & ~new_n16438_;
  assign new_n16440_ = ~new_n16435_ & new_n16439_;
  assign new_n16441_ = new_n14731_ & new_n16437_;
  assign new_n16442_ = new_n16392_ & ~new_n16441_;
  assign new_n16443_ = ~new_n16440_ & new_n16442_;
  assign new_n16444_ = ~new_n11126_ & ~new_n14427_;
  assign new_n16445_ = new_n16437_ & new_n16444_;
  assign new_n16446_ = new_n9069_ & new_n15740_;
  assign new_n16447_ = ~new_n6185_ & new_n15753_;
  assign new_n16448_ = pi0148 & ~new_n16447_;
  assign new_n16449_ = ~new_n16446_ & new_n16448_;
  assign new_n16450_ = ~pi0051 & new_n15293_;
  assign new_n16451_ = ~pi0148 & ~new_n16450_;
  assign new_n16452_ = ~new_n16422_ & ~new_n16451_;
  assign new_n16453_ = ~pi0148 & new_n14576_;
  assign new_n16454_ = ~new_n16452_ & ~new_n16453_;
  assign new_n16455_ = ~new_n16449_ & ~new_n16454_;
  assign new_n16456_ = pi0299 & ~new_n16455_;
  assign new_n16457_ = pi0184 & new_n15270_;
  assign new_n16458_ = new_n15759_ & ~new_n16457_;
  assign new_n16459_ = new_n16408_ & ~new_n16458_;
  assign new_n16460_ = pi0184 & new_n14660_;
  assign new_n16461_ = new_n15763_ & ~new_n16460_;
  assign new_n16462_ = new_n9739_ & ~new_n16461_;
  assign new_n16463_ = ~new_n16459_ & ~new_n16462_;
  assign new_n16464_ = ~new_n16456_ & new_n16463_;
  assign new_n16465_ = pi0232 & ~new_n16464_;
  assign new_n16466_ = ~pi0100 & new_n15739_;
  assign new_n16467_ = ~new_n16465_ & new_n16466_;
  assign new_n16468_ = ~new_n16445_ & ~new_n16467_;
  assign new_n16469_ = new_n3283_ & ~new_n16468_;
  assign new_n16470_ = ~new_n14427_ & new_n16441_;
  assign new_n16471_ = ~new_n16392_ & ~new_n16470_;
  assign new_n16472_ = ~new_n16469_ & new_n16471_;
  assign new_n16473_ = ~po1038 & ~new_n16472_;
  assign new_n16474_ = ~new_n16443_ & new_n16473_;
  assign po0293 = new_n16397_ | new_n16474_;
  assign new_n16476_ = ~pi0039 & pi0137;
  assign new_n16477_ = new_n10434_ & new_n14865_;
  assign new_n16478_ = new_n6165_ & new_n11568_;
  assign new_n16479_ = ~pi0299 & ~po1038;
  assign new_n16480_ = ~pi0198 & new_n11579_;
  assign new_n16481_ = new_n16479_ & new_n16480_;
  assign new_n16482_ = ~new_n16478_ & ~new_n16481_;
  assign new_n16483_ = ~new_n16477_ & ~new_n16482_;
  assign new_n16484_ = ~pi0210 & new_n11568_;
  assign new_n16485_ = po1038 & new_n16484_;
  assign new_n16486_ = ~new_n16483_ & ~new_n16485_;
  assign new_n16487_ = new_n10478_ & ~new_n16486_;
  assign po0294 = new_n16476_ | new_n16487_;
  assign new_n16489_ = ~new_n9472_ & new_n9522_;
  assign new_n16490_ = pi0092 & ~new_n16489_;
  assign new_n16491_ = new_n3270_ & ~new_n16490_;
  assign new_n16492_ = ~pi0075 & ~new_n9463_;
  assign new_n16493_ = ~pi0299 & ~new_n9789_;
  assign new_n16494_ = pi0299 & ~new_n9402_;
  assign new_n16495_ = ~pi0232 & ~new_n16494_;
  assign new_n16496_ = ~new_n16493_ & new_n16495_;
  assign new_n16497_ = ~pi0039 & ~new_n16496_;
  assign new_n16498_ = pi0148 & new_n6185_;
  assign new_n16499_ = ~new_n9402_ & ~new_n16498_;
  assign new_n16500_ = pi0148 & new_n13721_;
  assign new_n16501_ = ~new_n16499_ & ~new_n16500_;
  assign new_n16502_ = pi0299 & ~new_n16501_;
  assign new_n16503_ = ~new_n6185_ & ~new_n9789_;
  assign new_n16504_ = ~new_n13744_ & ~new_n16503_;
  assign new_n16505_ = ~pi0299 & ~new_n16504_;
  assign new_n16506_ = pi0141 & new_n16505_;
  assign new_n16507_ = ~pi0141 & new_n16493_;
  assign new_n16508_ = pi0232 & ~new_n16507_;
  assign new_n16509_ = ~new_n16506_ & new_n16508_;
  assign new_n16510_ = ~new_n16502_ & new_n16509_;
  assign new_n16511_ = new_n16497_ & ~new_n16510_;
  assign new_n16512_ = ~new_n9074_ & ~new_n11990_;
  assign new_n16513_ = new_n9094_ & ~new_n16512_;
  assign new_n16514_ = new_n13794_ & ~new_n16513_;
  assign new_n16515_ = ~new_n6212_ & ~new_n9074_;
  assign new_n16516_ = new_n9069_ & ~new_n16512_;
  assign new_n16517_ = ~new_n16515_ & new_n16516_;
  assign new_n16518_ = new_n9071_ & ~new_n16517_;
  assign new_n16519_ = ~new_n16514_ & ~new_n16518_;
  assign new_n16520_ = ~pi0232 & ~new_n16519_;
  assign new_n16521_ = ~new_n9079_ & ~new_n16512_;
  assign new_n16522_ = ~new_n9070_ & ~new_n16521_;
  assign new_n16523_ = pi0148 & ~new_n16522_;
  assign new_n16524_ = ~new_n9740_ & ~new_n16518_;
  assign new_n16525_ = ~new_n16523_ & ~new_n16524_;
  assign new_n16526_ = ~pi0141 & new_n16514_;
  assign new_n16527_ = ~new_n9102_ & new_n16513_;
  assign new_n16528_ = new_n13794_ & ~new_n16527_;
  assign new_n16529_ = pi0141 & new_n16528_;
  assign new_n16530_ = ~new_n16526_ & ~new_n16529_;
  assign new_n16531_ = ~new_n16525_ & new_n16530_;
  assign new_n16532_ = pi0232 & ~new_n16531_;
  assign new_n16533_ = ~new_n16520_ & ~new_n16532_;
  assign new_n16534_ = pi0039 & ~new_n16533_;
  assign new_n16535_ = new_n3211_ & ~new_n16534_;
  assign new_n16536_ = ~new_n16511_ & new_n16535_;
  assign new_n16537_ = ~pi0087 & ~new_n16536_;
  assign new_n16538_ = new_n16492_ & ~new_n16537_;
  assign new_n16539_ = ~pi0092 & ~new_n16538_;
  assign new_n16540_ = new_n16491_ & ~new_n16539_;
  assign new_n16541_ = ~pi0055 & ~new_n16540_;
  assign new_n16542_ = new_n9523_ & ~new_n13831_;
  assign new_n16543_ = pi0055 & ~new_n16542_;
  assign new_n16544_ = ~new_n16541_ & ~new_n16543_;
  assign new_n16545_ = new_n3298_ & ~new_n16544_;
  assign new_n16546_ = new_n9722_ & ~new_n16545_;
  assign new_n16547_ = pi0138 & new_n16546_;
  assign new_n16548_ = ~pi0232 & ~new_n11477_;
  assign new_n16549_ = ~new_n9739_ & ~new_n11477_;
  assign new_n16550_ = new_n6221_ & new_n6470_;
  assign new_n16551_ = new_n9058_ & new_n16550_;
  assign new_n16552_ = new_n9739_ & ~new_n16551_;
  assign new_n16553_ = ~new_n6221_ & new_n9740_;
  assign new_n16554_ = ~new_n16552_ & ~new_n16553_;
  assign new_n16555_ = ~new_n16549_ & new_n16554_;
  assign new_n16556_ = pi0232 & ~new_n16555_;
  assign new_n16557_ = ~new_n16548_ & ~new_n16556_;
  assign new_n16558_ = pi0039 & ~new_n16557_;
  assign new_n16559_ = ~new_n9742_ & new_n13901_;
  assign new_n16560_ = ~pi0039 & ~new_n16559_;
  assign new_n16561_ = new_n10200_ & ~new_n16560_;
  assign new_n16562_ = ~new_n16558_ & new_n16561_;
  assign new_n16563_ = ~pi0138 & new_n16562_;
  assign new_n16564_ = ~pi0118 & new_n13849_;
  assign new_n16565_ = ~pi0139 & new_n16564_;
  assign new_n16566_ = ~new_n16563_ & ~new_n16565_;
  assign new_n16567_ = ~new_n16547_ & new_n16566_;
  assign new_n16568_ = ~pi0138 & ~new_n8974_;
  assign new_n16569_ = new_n16546_ & new_n16568_;
  assign new_n16570_ = new_n16562_ & ~new_n16568_;
  assign new_n16571_ = new_n16565_ & ~new_n16570_;
  assign new_n16572_ = ~new_n16569_ & new_n16571_;
  assign po0295 = ~new_n16567_ & ~new_n16572_;
  assign new_n16574_ = ~new_n9402_ & ~new_n15747_;
  assign new_n16575_ = pi0169 & new_n13721_;
  assign new_n16576_ = ~new_n16574_ & ~new_n16575_;
  assign new_n16577_ = pi0299 & ~new_n16576_;
  assign new_n16578_ = pi0191 & new_n16505_;
  assign new_n16579_ = ~pi0191 & new_n16493_;
  assign new_n16580_ = pi0232 & ~new_n16579_;
  assign new_n16581_ = ~new_n16578_ & new_n16580_;
  assign new_n16582_ = ~new_n16577_ & new_n16581_;
  assign new_n16583_ = new_n16497_ & ~new_n16582_;
  assign new_n16584_ = pi0191 & new_n16528_;
  assign new_n16585_ = ~pi0169 & new_n9074_;
  assign new_n16586_ = ~new_n16521_ & ~new_n16585_;
  assign new_n16587_ = new_n9069_ & ~new_n16586_;
  assign new_n16588_ = new_n9071_ & ~new_n16587_;
  assign new_n16589_ = ~pi0191 & new_n16514_;
  assign new_n16590_ = ~new_n16588_ & ~new_n16589_;
  assign new_n16591_ = ~new_n16584_ & new_n16590_;
  assign new_n16592_ = pi0232 & ~new_n16591_;
  assign new_n16593_ = ~new_n16520_ & ~new_n16592_;
  assign new_n16594_ = pi0039 & ~new_n16593_;
  assign new_n16595_ = new_n3211_ & ~new_n16594_;
  assign new_n16596_ = ~new_n16583_ & new_n16595_;
  assign new_n16597_ = ~pi0087 & ~new_n16596_;
  assign new_n16598_ = new_n16492_ & ~new_n16597_;
  assign new_n16599_ = ~pi0092 & ~new_n16598_;
  assign new_n16600_ = new_n16491_ & ~new_n16599_;
  assign new_n16601_ = ~pi0055 & ~new_n16600_;
  assign new_n16602_ = ~new_n16543_ & ~new_n16601_;
  assign new_n16603_ = new_n3298_ & ~new_n16602_;
  assign new_n16604_ = new_n9722_ & ~new_n16603_;
  assign new_n16605_ = pi0139 & new_n16604_;
  assign new_n16606_ = ~new_n6221_ & new_n9011_;
  assign new_n16607_ = ~new_n11476_ & ~new_n16606_;
  assign new_n16608_ = ~new_n11473_ & new_n15758_;
  assign new_n16609_ = new_n9010_ & ~new_n16551_;
  assign new_n16610_ = ~new_n16608_ & ~new_n16609_;
  assign new_n16611_ = new_n16607_ & new_n16610_;
  assign new_n16612_ = pi0232 & ~new_n16611_;
  assign new_n16613_ = ~new_n16548_ & ~new_n16612_;
  assign new_n16614_ = pi0039 & ~new_n16613_;
  assign new_n16615_ = new_n13901_ & ~new_n15771_;
  assign new_n16616_ = ~pi0039 & ~new_n16615_;
  assign new_n16617_ = new_n10200_ & ~new_n16616_;
  assign new_n16618_ = ~new_n16614_ & new_n16617_;
  assign new_n16619_ = ~pi0139 & new_n16618_;
  assign new_n16620_ = ~new_n16564_ & ~new_n16619_;
  assign new_n16621_ = ~new_n16605_ & new_n16620_;
  assign new_n16622_ = ~pi0139 & ~new_n8975_;
  assign new_n16623_ = new_n16604_ & new_n16622_;
  assign new_n16624_ = new_n16618_ & ~new_n16622_;
  assign new_n16625_ = new_n16564_ & ~new_n16624_;
  assign new_n16626_ = ~new_n16623_ & new_n16625_;
  assign po0296 = ~new_n16621_ & ~new_n16626_;
  assign new_n16628_ = pi0140 & ~new_n3272_;
  assign new_n16629_ = ~pi0661 & ~pi0681;
  assign new_n16630_ = ~pi0662 & new_n16629_;
  assign new_n16631_ = pi0680 & ~new_n16630_;
  assign new_n16632_ = ~new_n6189_ & new_n6454_;
  assign new_n16633_ = ~pi0120 & ~new_n16632_;
  assign new_n16634_ = pi0120 & ~new_n3100_;
  assign new_n16635_ = ~new_n16633_ & ~new_n16634_;
  assign new_n16636_ = new_n2754_ & new_n16635_;
  assign new_n16637_ = pi0665 & pi1091;
  assign new_n16638_ = pi0621 & pi1091;
  assign new_n16639_ = pi0603 & ~new_n16638_;
  assign new_n16640_ = ~new_n16637_ & ~new_n16639_;
  assign new_n16641_ = new_n16636_ & ~new_n16640_;
  assign new_n16642_ = pi0616 & ~new_n16641_;
  assign new_n16643_ = pi0614 & ~new_n16641_;
  assign new_n16644_ = pi0642 & ~new_n16641_;
  assign new_n16645_ = new_n2754_ & new_n16632_;
  assign new_n16646_ = ~pi0120 & ~new_n16645_;
  assign new_n16647_ = new_n2754_ & new_n3100_;
  assign new_n16648_ = new_n6192_ & new_n14279_;
  assign new_n16649_ = new_n16647_ & ~new_n16648_;
  assign new_n16650_ = pi0120 & ~new_n16649_;
  assign new_n16651_ = pi1091 & ~new_n16650_;
  assign new_n16652_ = ~new_n16646_ & new_n16651_;
  assign new_n16653_ = pi0665 & new_n16652_;
  assign new_n16654_ = pi0120 & ~new_n16647_;
  assign new_n16655_ = ~pi1091 & ~new_n16654_;
  assign new_n16656_ = pi0120 & pi0824;
  assign new_n16657_ = new_n6192_ & new_n16656_;
  assign new_n16658_ = new_n16655_ & ~new_n16657_;
  assign new_n16659_ = ~new_n16646_ & new_n16658_;
  assign new_n16660_ = ~new_n16652_ & ~new_n16659_;
  assign new_n16661_ = new_n16636_ & new_n16639_;
  assign new_n16662_ = ~new_n16660_ & new_n16661_;
  assign new_n16663_ = ~new_n16653_ & ~new_n16662_;
  assign new_n16664_ = ~new_n6185_ & new_n16636_;
  assign new_n16665_ = new_n16637_ & new_n16664_;
  assign new_n16666_ = ~pi0603 & new_n16665_;
  assign new_n16667_ = new_n16663_ & ~new_n16666_;
  assign new_n16668_ = ~new_n6185_ & new_n16660_;
  assign new_n16669_ = new_n16661_ & ~new_n16668_;
  assign new_n16670_ = new_n16636_ & new_n16637_;
  assign new_n16671_ = new_n6185_ & ~new_n16670_;
  assign new_n16672_ = ~new_n6185_ & ~new_n16653_;
  assign new_n16673_ = ~new_n16671_ & ~new_n16672_;
  assign new_n16674_ = ~pi0642 & ~new_n16673_;
  assign new_n16675_ = ~new_n16669_ & new_n16674_;
  assign new_n16676_ = new_n16667_ & new_n16675_;
  assign new_n16677_ = ~new_n16644_ & ~new_n16676_;
  assign new_n16678_ = ~pi0614 & ~new_n16677_;
  assign new_n16679_ = ~new_n16643_ & ~new_n16678_;
  assign new_n16680_ = ~pi0616 & ~new_n16679_;
  assign new_n16681_ = ~new_n16642_ & ~new_n16680_;
  assign new_n16682_ = new_n16631_ & ~new_n16681_;
  assign new_n16683_ = pi0616 & ~new_n16636_;
  assign new_n16684_ = pi0614 & ~new_n16636_;
  assign new_n16685_ = ~new_n6178_ & ~new_n16636_;
  assign new_n16686_ = new_n6185_ & ~new_n16636_;
  assign new_n16687_ = ~new_n16668_ & ~new_n16686_;
  assign new_n16688_ = new_n6178_ & ~new_n16687_;
  assign new_n16689_ = ~new_n16685_ & ~new_n16688_;
  assign new_n16690_ = ~pi0614 & ~new_n16689_;
  assign new_n16691_ = ~new_n16684_ & ~new_n16690_;
  assign new_n16692_ = ~pi0616 & ~new_n16691_;
  assign new_n16693_ = ~new_n16683_ & ~new_n16692_;
  assign new_n16694_ = ~pi0680 & ~new_n16693_;
  assign new_n16695_ = new_n6183_ & ~new_n16673_;
  assign new_n16696_ = ~new_n16669_ & new_n16695_;
  assign new_n16697_ = ~new_n16694_ & ~new_n16696_;
  assign new_n16698_ = ~new_n16682_ & new_n16697_;
  assign new_n16699_ = new_n6238_ & ~new_n16698_;
  assign new_n16700_ = new_n6185_ & ~new_n16660_;
  assign new_n16701_ = ~new_n16664_ & ~new_n16700_;
  assign new_n16702_ = ~pi0616 & new_n16690_;
  assign new_n16703_ = ~new_n16701_ & ~new_n16702_;
  assign new_n16704_ = ~pi0680 & ~new_n16703_;
  assign new_n16705_ = new_n6183_ & new_n16663_;
  assign new_n16706_ = ~pi0614 & ~pi0642;
  assign new_n16707_ = ~pi0616 & new_n16706_;
  assign new_n16708_ = new_n16661_ & ~new_n16701_;
  assign new_n16709_ = ~new_n16653_ & ~new_n16665_;
  assign new_n16710_ = ~new_n16708_ & new_n16709_;
  assign new_n16711_ = ~new_n16707_ & new_n16710_;
  assign new_n16712_ = new_n16667_ & new_n16707_;
  assign new_n16713_ = ~new_n16711_ & ~new_n16712_;
  assign new_n16714_ = new_n16631_ & ~new_n16713_;
  assign new_n16715_ = ~new_n16705_ & ~new_n16714_;
  assign new_n16716_ = ~new_n16704_ & new_n16715_;
  assign new_n16717_ = ~new_n6238_ & ~new_n16716_;
  assign new_n16718_ = pi0223 & ~new_n16717_;
  assign new_n16719_ = ~new_n16699_ & new_n16718_;
  assign new_n16720_ = ~pi0603 & ~new_n16636_;
  assign new_n16721_ = ~pi0824 & ~new_n16632_;
  assign new_n16722_ = new_n6454_ & ~new_n10203_;
  assign new_n16723_ = pi1092 & new_n16722_;
  assign new_n16724_ = ~new_n11032_ & ~new_n16723_;
  assign new_n16725_ = ~new_n16721_ & ~new_n16724_;
  assign new_n16726_ = pi1093 & new_n16725_;
  assign new_n16727_ = ~pi0120 & ~new_n16726_;
  assign new_n16728_ = new_n16655_ & ~new_n16727_;
  assign new_n16729_ = new_n2732_ & new_n16645_;
  assign new_n16730_ = ~pi0829 & ~new_n16725_;
  assign new_n16731_ = pi0829 & ~new_n16723_;
  assign new_n16732_ = new_n7510_ & ~new_n16731_;
  assign new_n16733_ = ~new_n16730_ & new_n16732_;
  assign new_n16734_ = ~new_n16729_ & ~new_n16733_;
  assign new_n16735_ = pi1091 & ~new_n16734_;
  assign new_n16736_ = ~pi0120 & ~new_n16735_;
  assign new_n16737_ = ~new_n16654_ & ~new_n16736_;
  assign new_n16738_ = ~new_n16728_ & ~new_n16737_;
  assign new_n16739_ = ~new_n6185_ & new_n16738_;
  assign new_n16740_ = ~new_n16686_ & ~new_n16739_;
  assign new_n16741_ = pi0603 & ~new_n16740_;
  assign new_n16742_ = ~new_n16720_ & ~new_n16741_;
  assign new_n16743_ = ~new_n16640_ & new_n16742_;
  assign new_n16744_ = ~pi0642 & ~new_n16743_;
  assign new_n16745_ = ~new_n16644_ & ~new_n16744_;
  assign new_n16746_ = ~pi0614 & ~new_n16745_;
  assign new_n16747_ = ~new_n16643_ & ~new_n16746_;
  assign new_n16748_ = ~pi0616 & ~new_n16747_;
  assign new_n16749_ = ~new_n16642_ & ~new_n16748_;
  assign new_n16750_ = new_n16631_ & ~new_n16749_;
  assign new_n16751_ = ~pi0642 & ~new_n16742_;
  assign new_n16752_ = ~new_n16685_ & ~new_n16751_;
  assign new_n16753_ = ~pi0614 & ~new_n16752_;
  assign new_n16754_ = ~new_n16684_ & ~new_n16753_;
  assign new_n16755_ = ~pi0616 & ~new_n16754_;
  assign new_n16756_ = ~new_n16683_ & ~new_n16755_;
  assign new_n16757_ = ~pi0680 & ~new_n16756_;
  assign new_n16758_ = new_n16637_ & new_n16737_;
  assign new_n16759_ = ~new_n6185_ & ~new_n16758_;
  assign new_n16760_ = ~new_n16671_ & ~new_n16759_;
  assign new_n16761_ = ~pi0603 & ~new_n16760_;
  assign new_n16762_ = pi0603 & ~pi0665;
  assign new_n16763_ = new_n16638_ & new_n16762_;
  assign new_n16764_ = ~new_n16741_ & ~new_n16763_;
  assign new_n16765_ = ~new_n16761_ & new_n16764_;
  assign new_n16766_ = new_n6183_ & ~new_n16765_;
  assign new_n16767_ = ~new_n16757_ & ~new_n16766_;
  assign new_n16768_ = ~new_n16750_ & new_n16767_;
  assign new_n16769_ = new_n6238_ & new_n16768_;
  assign new_n16770_ = new_n6185_ & ~new_n16738_;
  assign new_n16771_ = ~new_n16664_ & ~new_n16770_;
  assign new_n16772_ = ~new_n6180_ & new_n16771_;
  assign new_n16773_ = new_n6180_ & new_n16738_;
  assign new_n16774_ = ~new_n16772_ & ~new_n16773_;
  assign new_n16775_ = ~new_n16640_ & new_n16774_;
  assign new_n16776_ = new_n16631_ & ~new_n16775_;
  assign new_n16777_ = ~pi0680 & ~new_n16774_;
  assign new_n16778_ = pi0621 & ~new_n16728_;
  assign new_n16779_ = ~new_n16738_ & ~new_n16778_;
  assign new_n16780_ = pi0603 & new_n16779_;
  assign new_n16781_ = pi0603 & ~pi0621;
  assign new_n16782_ = new_n16758_ & ~new_n16781_;
  assign new_n16783_ = new_n6183_ & ~new_n16782_;
  assign new_n16784_ = ~new_n16780_ & new_n16783_;
  assign new_n16785_ = ~new_n16777_ & ~new_n16784_;
  assign new_n16786_ = ~new_n16776_ & new_n16785_;
  assign new_n16787_ = ~new_n6238_ & new_n16786_;
  assign new_n16788_ = ~new_n3057_ & ~new_n16787_;
  assign new_n16789_ = ~new_n16769_ & new_n16788_;
  assign new_n16790_ = pi0680 & new_n16640_;
  assign new_n16791_ = new_n16636_ & ~new_n16790_;
  assign new_n16792_ = new_n3057_ & ~new_n16791_;
  assign new_n16793_ = ~pi0223 & ~new_n16792_;
  assign new_n16794_ = ~new_n16789_ & new_n16793_;
  assign new_n16795_ = ~new_n16719_ & ~new_n16794_;
  assign new_n16796_ = ~pi0299 & ~new_n16795_;
  assign new_n16797_ = ~new_n6212_ & ~new_n16786_;
  assign new_n16798_ = new_n6212_ & ~new_n16768_;
  assign new_n16799_ = ~new_n16797_ & ~new_n16798_;
  assign new_n16800_ = ~new_n3467_ & ~new_n16799_;
  assign new_n16801_ = new_n3467_ & ~new_n16791_;
  assign new_n16802_ = ~pi0215 & ~new_n16801_;
  assign new_n16803_ = ~new_n16800_ & new_n16802_;
  assign new_n16804_ = new_n6212_ & ~new_n16698_;
  assign new_n16805_ = ~new_n6212_ & ~new_n16716_;
  assign new_n16806_ = pi0215 & ~new_n16805_;
  assign new_n16807_ = ~new_n16804_ & new_n16806_;
  assign new_n16808_ = ~new_n16803_ & ~new_n16807_;
  assign new_n16809_ = pi0299 & ~new_n16808_;
  assign new_n16810_ = ~new_n16796_ & ~new_n16809_;
  assign new_n16811_ = ~pi0140 & new_n16810_;
  assign new_n16812_ = new_n16636_ & ~new_n16637_;
  assign new_n16813_ = pi0665 & ~new_n16728_;
  assign new_n16814_ = ~new_n16738_ & ~new_n16813_;
  assign new_n16815_ = ~new_n16812_ & ~new_n16814_;
  assign new_n16816_ = ~pi0603 & new_n16771_;
  assign new_n16817_ = new_n16638_ & new_n16737_;
  assign new_n16818_ = new_n6185_ & new_n16817_;
  assign new_n16819_ = new_n16638_ & new_n16664_;
  assign new_n16820_ = pi0603 & ~new_n16819_;
  assign new_n16821_ = ~new_n16818_ & new_n16820_;
  assign new_n16822_ = ~new_n16816_ & ~new_n16821_;
  assign new_n16823_ = ~new_n16815_ & new_n16822_;
  assign new_n16824_ = pi0616 & ~new_n16823_;
  assign new_n16825_ = ~pi0665 & new_n16817_;
  assign new_n16826_ = pi0603 & ~new_n16825_;
  assign new_n16827_ = ~new_n16771_ & ~new_n16815_;
  assign new_n16828_ = ~pi0603 & ~new_n16827_;
  assign new_n16829_ = ~new_n16826_ & ~new_n16828_;
  assign new_n16830_ = new_n16707_ & ~new_n16829_;
  assign new_n16831_ = new_n16823_ & ~new_n16830_;
  assign new_n16832_ = new_n16706_ & new_n16829_;
  assign new_n16833_ = ~pi0616 & ~new_n16832_;
  assign new_n16834_ = ~new_n16831_ & new_n16833_;
  assign new_n16835_ = ~new_n16824_ & ~new_n16834_;
  assign new_n16836_ = ~new_n16630_ & ~new_n16835_;
  assign new_n16837_ = new_n6183_ & new_n16814_;
  assign new_n16838_ = ~new_n16826_ & new_n16837_;
  assign new_n16839_ = ~new_n16631_ & ~new_n16838_;
  assign new_n16840_ = ~new_n16836_ & ~new_n16839_;
  assign new_n16841_ = ~new_n6212_ & ~new_n16840_;
  assign new_n16842_ = new_n16636_ & ~new_n16639_;
  assign new_n16843_ = ~new_n16637_ & new_n16842_;
  assign new_n16844_ = pi0616 & ~new_n16843_;
  assign new_n16845_ = new_n16631_ & ~new_n16844_;
  assign new_n16846_ = new_n16636_ & new_n16638_;
  assign new_n16847_ = new_n6185_ & ~new_n16846_;
  assign new_n16848_ = ~new_n6185_ & ~new_n16817_;
  assign new_n16849_ = ~new_n16847_ & ~new_n16848_;
  assign new_n16850_ = pi0603 & ~new_n16849_;
  assign new_n16851_ = pi0603 & pi0665;
  assign new_n16852_ = ~pi0603 & ~new_n16812_;
  assign new_n16853_ = ~new_n16851_ & ~new_n16852_;
  assign new_n16854_ = ~new_n16850_ & new_n16853_;
  assign new_n16855_ = new_n16706_ & new_n16854_;
  assign new_n16856_ = ~new_n16706_ & new_n16843_;
  assign new_n16857_ = ~pi0616 & ~new_n16856_;
  assign new_n16858_ = ~new_n16855_ & new_n16857_;
  assign new_n16859_ = new_n16845_ & ~new_n16858_;
  assign new_n16860_ = new_n16740_ & new_n16766_;
  assign new_n16861_ = ~new_n16859_ & ~new_n16860_;
  assign new_n16862_ = new_n6212_ & new_n16861_;
  assign new_n16863_ = ~new_n3467_ & ~new_n16862_;
  assign new_n16864_ = ~new_n16841_ & new_n16863_;
  assign new_n16865_ = new_n3467_ & new_n16636_;
  assign new_n16866_ = new_n16790_ & new_n16865_;
  assign new_n16867_ = ~pi0215 & ~new_n16866_;
  assign new_n16868_ = ~new_n16864_ & new_n16867_;
  assign new_n16869_ = new_n2754_ & ~new_n16639_;
  assign new_n16870_ = ~new_n16701_ & new_n16869_;
  assign new_n16871_ = new_n16853_ & new_n16870_;
  assign new_n16872_ = pi0616 & ~new_n16871_;
  assign new_n16873_ = pi0614 & ~pi0616;
  assign new_n16874_ = ~new_n16871_ & new_n16873_;
  assign new_n16875_ = pi0621 & new_n16652_;
  assign new_n16876_ = ~new_n6185_ & ~new_n16875_;
  assign new_n16877_ = ~new_n16847_ & ~new_n16876_;
  assign new_n16878_ = pi0603 & ~new_n16877_;
  assign new_n16879_ = new_n16853_ & ~new_n16878_;
  assign new_n16880_ = ~pi0642 & ~new_n16879_;
  assign new_n16881_ = new_n16871_ & ~new_n16880_;
  assign new_n16882_ = new_n6179_ & ~new_n16881_;
  assign new_n16883_ = ~new_n16874_ & ~new_n16882_;
  assign new_n16884_ = ~new_n16872_ & new_n16883_;
  assign new_n16885_ = ~new_n16630_ & ~new_n16884_;
  assign new_n16886_ = ~new_n16660_ & new_n16790_;
  assign new_n16887_ = ~new_n16631_ & ~new_n16886_;
  assign new_n16888_ = ~new_n16885_ & ~new_n16887_;
  assign new_n16889_ = ~new_n6212_ & new_n16888_;
  assign new_n16890_ = ~new_n16707_ & new_n16842_;
  assign new_n16891_ = new_n16707_ & ~new_n16720_;
  assign new_n16892_ = ~new_n16878_ & new_n16891_;
  assign new_n16893_ = ~new_n16890_ & ~new_n16892_;
  assign new_n16894_ = ~new_n16637_ & ~new_n16893_;
  assign new_n16895_ = ~pi0616 & ~new_n16894_;
  assign new_n16896_ = new_n16845_ & ~new_n16895_;
  assign new_n16897_ = new_n6183_ & new_n16687_;
  assign new_n16898_ = ~new_n16878_ & new_n16897_;
  assign new_n16899_ = new_n16853_ & new_n16898_;
  assign new_n16900_ = ~new_n16896_ & ~new_n16899_;
  assign new_n16901_ = new_n6212_ & ~new_n16900_;
  assign new_n16902_ = pi0215 & ~new_n16901_;
  assign new_n16903_ = ~new_n16889_ & new_n16902_;
  assign new_n16904_ = ~new_n16868_ & ~new_n16903_;
  assign new_n16905_ = pi0299 & ~new_n16904_;
  assign new_n16906_ = ~new_n6238_ & new_n16840_;
  assign new_n16907_ = new_n6238_ & ~new_n16861_;
  assign new_n16908_ = ~new_n3057_ & ~new_n16907_;
  assign new_n16909_ = ~new_n16906_ & new_n16908_;
  assign new_n16910_ = new_n3057_ & new_n16636_;
  assign new_n16911_ = new_n16639_ & new_n16910_;
  assign new_n16912_ = ~pi0223 & ~new_n16911_;
  assign new_n16913_ = new_n2754_ & new_n16639_;
  assign new_n16914_ = pi0680 & ~new_n16637_;
  assign new_n16915_ = new_n2754_ & new_n16914_;
  assign new_n16916_ = ~new_n16639_ & new_n16915_;
  assign new_n16917_ = ~new_n16913_ & ~new_n16916_;
  assign new_n16918_ = new_n16636_ & ~new_n16917_;
  assign new_n16919_ = new_n3057_ & ~new_n16918_;
  assign new_n16920_ = new_n16912_ & ~new_n16919_;
  assign new_n16921_ = ~new_n16909_ & new_n16920_;
  assign new_n16922_ = ~new_n6238_ & ~new_n16888_;
  assign new_n16923_ = new_n6238_ & new_n16900_;
  assign new_n16924_ = pi0223 & ~new_n16923_;
  assign new_n16925_ = ~new_n16922_ & new_n16924_;
  assign new_n16926_ = ~pi0299 & ~new_n16925_;
  assign new_n16927_ = ~new_n16921_ & new_n16926_;
  assign new_n16928_ = ~new_n16905_ & ~new_n16927_;
  assign new_n16929_ = pi0140 & new_n16928_;
  assign new_n16930_ = pi0761 & ~new_n16929_;
  assign new_n16931_ = ~new_n16811_ & new_n16930_;
  assign new_n16932_ = ~new_n16780_ & ~new_n16829_;
  assign new_n16933_ = new_n16707_ & ~new_n16932_;
  assign new_n16934_ = new_n16639_ & ~new_n16771_;
  assign new_n16935_ = ~new_n16827_ & ~new_n16934_;
  assign new_n16936_ = ~new_n16707_ & ~new_n16935_;
  assign new_n16937_ = new_n16631_ & ~new_n16936_;
  assign new_n16938_ = ~new_n16933_ & new_n16937_;
  assign new_n16939_ = ~new_n6183_ & ~new_n16774_;
  assign new_n16940_ = new_n6183_ & new_n16738_;
  assign new_n16941_ = ~new_n16939_ & ~new_n16940_;
  assign new_n16942_ = new_n16639_ & new_n16941_;
  assign new_n16943_ = ~new_n16631_ & ~new_n16837_;
  assign new_n16944_ = ~new_n16942_ & new_n16943_;
  assign new_n16945_ = ~new_n16938_ & ~new_n16944_;
  assign new_n16946_ = ~new_n6238_ & new_n16945_;
  assign new_n16947_ = new_n16637_ & ~new_n16781_;
  assign new_n16948_ = new_n16636_ & ~new_n16947_;
  assign new_n16949_ = ~new_n16707_ & new_n16948_;
  assign new_n16950_ = new_n16631_ & ~new_n16949_;
  assign new_n16951_ = new_n16639_ & new_n16740_;
  assign new_n16952_ = ~new_n16854_ & ~new_n16951_;
  assign new_n16953_ = new_n16707_ & ~new_n16952_;
  assign new_n16954_ = new_n16950_ & ~new_n16953_;
  assign new_n16955_ = new_n16661_ & ~new_n16707_;
  assign new_n16956_ = new_n16707_ & new_n16951_;
  assign new_n16957_ = ~new_n16955_ & ~new_n16956_;
  assign new_n16958_ = ~pi0680 & new_n16957_;
  assign new_n16959_ = new_n16740_ & ~new_n16815_;
  assign new_n16960_ = new_n6183_ & ~new_n16959_;
  assign new_n16961_ = ~new_n16951_ & new_n16960_;
  assign new_n16962_ = ~new_n16958_ & ~new_n16961_;
  assign new_n16963_ = ~new_n16954_ & new_n16962_;
  assign new_n16964_ = new_n6238_ & new_n16963_;
  assign new_n16965_ = ~new_n3057_ & ~new_n16964_;
  assign new_n16966_ = ~new_n16946_ & new_n16965_;
  assign new_n16967_ = ~pi0223 & ~new_n16919_;
  assign new_n16968_ = ~new_n16966_ & new_n16967_;
  assign new_n16969_ = ~new_n6180_ & new_n16812_;
  assign new_n16970_ = ~new_n16668_ & new_n16812_;
  assign new_n16971_ = ~new_n16969_ & ~new_n16970_;
  assign new_n16972_ = ~new_n16669_ & new_n16971_;
  assign new_n16973_ = new_n16707_ & ~new_n16972_;
  assign new_n16974_ = new_n16950_ & ~new_n16973_;
  assign new_n16975_ = new_n16668_ & new_n16707_;
  assign new_n16976_ = new_n16708_ & ~new_n16975_;
  assign new_n16977_ = ~new_n6183_ & new_n16976_;
  assign new_n16978_ = ~new_n16669_ & ~new_n16977_;
  assign new_n16979_ = new_n16630_ & ~new_n16970_;
  assign new_n16980_ = pi0680 & ~new_n16979_;
  assign new_n16981_ = new_n16978_ & ~new_n16980_;
  assign new_n16982_ = ~new_n16974_ & ~new_n16981_;
  assign new_n16983_ = new_n6238_ & ~new_n16982_;
  assign new_n16984_ = ~new_n16662_ & ~new_n16977_;
  assign new_n16985_ = ~new_n16701_ & new_n16812_;
  assign new_n16986_ = ~new_n16971_ & new_n16980_;
  assign new_n16987_ = new_n16985_ & new_n16986_;
  assign new_n16988_ = new_n16984_ & ~new_n16987_;
  assign new_n16989_ = ~new_n6238_ & new_n16988_;
  assign new_n16990_ = pi0223 & ~new_n16989_;
  assign new_n16991_ = ~new_n16983_ & new_n16990_;
  assign new_n16992_ = ~pi0299 & ~new_n16991_;
  assign new_n16993_ = ~new_n16968_ & new_n16992_;
  assign new_n16994_ = ~new_n6212_ & new_n16945_;
  assign new_n16995_ = new_n6212_ & new_n16963_;
  assign new_n16996_ = ~new_n16994_ & ~new_n16995_;
  assign new_n16997_ = ~new_n3467_ & ~new_n16996_;
  assign new_n16998_ = new_n3467_ & new_n16918_;
  assign new_n16999_ = ~pi0215 & ~new_n16998_;
  assign new_n17000_ = ~new_n16997_ & new_n16999_;
  assign new_n17001_ = new_n6212_ & new_n16982_;
  assign new_n17002_ = ~new_n6212_ & ~new_n16988_;
  assign new_n17003_ = pi0215 & ~new_n17002_;
  assign new_n17004_ = ~new_n17001_ & new_n17003_;
  assign new_n17005_ = ~new_n17000_ & ~new_n17004_;
  assign new_n17006_ = pi0299 & ~new_n17005_;
  assign new_n17007_ = ~new_n16993_ & ~new_n17006_;
  assign new_n17008_ = pi0140 & new_n17007_;
  assign new_n17009_ = ~new_n16639_ & new_n16774_;
  assign new_n17010_ = ~pi0680 & ~new_n17009_;
  assign new_n17011_ = ~new_n6214_ & new_n16758_;
  assign new_n17012_ = ~new_n6180_ & new_n16665_;
  assign new_n17013_ = ~new_n17011_ & ~new_n17012_;
  assign new_n17014_ = new_n16947_ & ~new_n17013_;
  assign new_n17015_ = new_n16631_ & ~new_n17014_;
  assign new_n17016_ = ~new_n16783_ & ~new_n17015_;
  assign new_n17017_ = ~new_n17010_ & new_n17016_;
  assign new_n17018_ = ~new_n6238_ & new_n17017_;
  assign new_n17019_ = ~new_n16850_ & new_n16891_;
  assign new_n17020_ = new_n16637_ & new_n17019_;
  assign new_n17021_ = new_n16670_ & ~new_n16781_;
  assign new_n17022_ = ~new_n16707_ & new_n17021_;
  assign new_n17023_ = new_n16631_ & ~new_n17022_;
  assign new_n17024_ = ~new_n17020_ & new_n17023_;
  assign new_n17025_ = ~new_n16890_ & ~new_n17019_;
  assign new_n17026_ = ~pi0680 & new_n17025_;
  assign new_n17027_ = new_n16760_ & new_n16947_;
  assign new_n17028_ = new_n6183_ & ~new_n17027_;
  assign new_n17029_ = ~new_n17026_ & ~new_n17028_;
  assign new_n17030_ = ~new_n17024_ & new_n17029_;
  assign new_n17031_ = new_n6238_ & new_n17030_;
  assign new_n17032_ = ~new_n17018_ & ~new_n17031_;
  assign new_n17033_ = ~new_n3057_ & ~new_n17032_;
  assign new_n17034_ = ~new_n16639_ & ~new_n16914_;
  assign new_n17035_ = new_n16647_ & new_n17034_;
  assign new_n17036_ = ~new_n16633_ & new_n17035_;
  assign new_n17037_ = new_n3057_ & new_n17036_;
  assign new_n17038_ = ~pi0223 & ~new_n17037_;
  assign new_n17039_ = ~new_n17033_ & new_n17038_;
  assign new_n17040_ = ~new_n16709_ & ~new_n16893_;
  assign new_n17041_ = new_n16631_ & ~new_n17040_;
  assign new_n17042_ = new_n6180_ & ~new_n16652_;
  assign new_n17043_ = new_n16870_ & ~new_n17042_;
  assign new_n17044_ = ~pi0680 & ~new_n17043_;
  assign new_n17045_ = pi0680 & ~new_n16653_;
  assign new_n17046_ = ~new_n16781_ & ~new_n17045_;
  assign new_n17047_ = new_n6183_ & ~new_n17046_;
  assign new_n17048_ = ~new_n17044_ & ~new_n17047_;
  assign new_n17049_ = ~new_n17041_ & new_n17048_;
  assign new_n17050_ = ~new_n6238_ & new_n17049_;
  assign new_n17051_ = ~new_n6183_ & ~new_n16893_;
  assign new_n17052_ = ~new_n16914_ & new_n17051_;
  assign new_n17053_ = new_n6183_ & ~new_n16781_;
  assign new_n17054_ = new_n16673_ & new_n17053_;
  assign new_n17055_ = ~new_n17052_ & ~new_n17054_;
  assign new_n17056_ = new_n6238_ & ~new_n17055_;
  assign new_n17057_ = pi0223 & ~new_n17056_;
  assign new_n17058_ = ~new_n17050_ & new_n17057_;
  assign new_n17059_ = ~new_n17039_ & ~new_n17058_;
  assign new_n17060_ = ~pi0299 & ~new_n17059_;
  assign new_n17061_ = ~new_n6212_ & new_n17017_;
  assign new_n17062_ = new_n6212_ & new_n17030_;
  assign new_n17063_ = ~new_n17061_ & ~new_n17062_;
  assign new_n17064_ = ~new_n3467_ & ~new_n17063_;
  assign new_n17065_ = new_n3467_ & new_n17036_;
  assign new_n17066_ = ~pi0215 & ~new_n17065_;
  assign new_n17067_ = ~new_n17064_ & new_n17066_;
  assign new_n17068_ = ~new_n6212_ & new_n17049_;
  assign new_n17069_ = new_n6212_ & ~new_n17055_;
  assign new_n17070_ = pi0215 & ~new_n17069_;
  assign new_n17071_ = ~new_n17068_ & new_n17070_;
  assign new_n17072_ = ~new_n17067_ & ~new_n17071_;
  assign new_n17073_ = pi0299 & ~new_n17072_;
  assign new_n17074_ = ~new_n17060_ & ~new_n17073_;
  assign new_n17075_ = ~pi0140 & ~new_n17074_;
  assign new_n17076_ = ~pi0761 & ~new_n17075_;
  assign new_n17077_ = ~new_n17008_ & new_n17076_;
  assign new_n17078_ = ~new_n16931_ & ~new_n17077_;
  assign new_n17079_ = pi0039 & ~new_n17078_;
  assign new_n17080_ = ~pi0102 & ~new_n11299_;
  assign new_n17081_ = ~pi0098 & ~new_n2596_;
  assign new_n17082_ = ~new_n17080_ & new_n17081_;
  assign new_n17083_ = new_n7463_ & new_n12190_;
  assign new_n17084_ = new_n17082_ & new_n17083_;
  assign new_n17085_ = new_n8899_ & new_n9170_;
  assign new_n17086_ = new_n17084_ & new_n17085_;
  assign new_n17087_ = ~pi0040 & ~new_n17086_;
  assign new_n17088_ = new_n10281_ & ~new_n17087_;
  assign new_n17089_ = ~pi0252 & ~new_n17088_;
  assign new_n17090_ = new_n2536_ & new_n2572_;
  assign new_n17091_ = new_n8898_ & new_n17084_;
  assign new_n17092_ = ~pi0047 & ~new_n17091_;
  assign new_n17093_ = pi0314 & new_n10256_;
  assign new_n17094_ = new_n17092_ & ~new_n17093_;
  assign new_n17095_ = new_n17090_ & ~new_n17094_;
  assign new_n17096_ = ~pi0035 & ~new_n17095_;
  assign new_n17097_ = ~pi0040 & new_n10274_;
  assign new_n17098_ = ~new_n17096_ & new_n17097_;
  assign new_n17099_ = pi0252 & ~new_n2553_;
  assign new_n17100_ = ~new_n17098_ & new_n17099_;
  assign new_n17101_ = ~new_n17089_ & ~new_n17100_;
  assign new_n17102_ = new_n3097_ & new_n17101_;
  assign new_n17103_ = pi1092 & ~new_n12202_;
  assign new_n17104_ = new_n17102_ & new_n17103_;
  assign new_n17105_ = ~pi0088 & ~new_n17082_;
  assign new_n17106_ = new_n11006_ & ~new_n17105_;
  assign new_n17107_ = new_n2519_ & new_n17106_;
  assign new_n17108_ = ~pi0047 & ~new_n17093_;
  assign new_n17109_ = ~new_n17107_ & new_n17108_;
  assign new_n17110_ = new_n17090_ & ~new_n17109_;
  assign new_n17111_ = ~pi0035 & ~new_n17110_;
  assign new_n17112_ = pi0252 & new_n10274_;
  assign new_n17113_ = ~new_n17111_ & new_n17112_;
  assign new_n17114_ = ~pi0252 & new_n9313_;
  assign new_n17115_ = new_n17106_ & new_n17114_;
  assign new_n17116_ = ~pi0040 & ~new_n17115_;
  assign new_n17117_ = ~new_n17113_ & new_n17116_;
  assign new_n17118_ = new_n7511_ & new_n10281_;
  assign new_n17119_ = ~new_n17117_ & new_n17118_;
  assign new_n17120_ = ~new_n17104_ & ~new_n17119_;
  assign new_n17121_ = pi1093 & ~new_n17120_;
  assign new_n17122_ = ~new_n2732_ & ~new_n17121_;
  assign new_n17123_ = pi1092 & new_n2797_;
  assign po1106 = new_n2732_ & new_n17123_;
  assign new_n17125_ = new_n17102_ & po1106;
  assign new_n17126_ = ~new_n2733_ & ~new_n17125_;
  assign new_n17127_ = ~new_n17122_ & ~new_n17126_;
  assign new_n17128_ = ~pi1091 & new_n17121_;
  assign new_n17129_ = ~new_n17127_ & ~new_n17128_;
  assign new_n17130_ = pi0665 & ~new_n17128_;
  assign new_n17131_ = ~new_n17129_ & ~new_n17130_;
  assign new_n17132_ = ~pi0198 & ~new_n17131_;
  assign new_n17133_ = ~new_n3366_ & ~new_n17117_;
  assign new_n17134_ = ~pi0032 & ~new_n17133_;
  assign new_n17135_ = pi0032 & ~new_n6385_;
  assign new_n17136_ = ~pi0095 & new_n2799_;
  assign new_n17137_ = ~new_n17135_ & new_n17136_;
  assign new_n17138_ = ~new_n17134_ & new_n17137_;
  assign new_n17139_ = pi0824 & new_n17138_;
  assign new_n17140_ = ~new_n17104_ & ~new_n17139_;
  assign new_n17141_ = new_n7572_ & ~new_n17140_;
  assign new_n17142_ = ~pi0032 & ~new_n17101_;
  assign new_n17143_ = new_n17137_ & ~new_n17142_;
  assign new_n17144_ = ~pi0824 & pi0829;
  assign new_n17145_ = new_n17143_ & new_n17144_;
  assign new_n17146_ = new_n17140_ & ~new_n17145_;
  assign new_n17147_ = pi1093 & ~new_n17146_;
  assign new_n17148_ = ~new_n2732_ & ~new_n17147_;
  assign new_n17149_ = ~new_n17126_ & ~new_n17148_;
  assign new_n17150_ = ~new_n17141_ & ~new_n17149_;
  assign new_n17151_ = pi0665 & ~new_n17141_;
  assign new_n17152_ = ~new_n17150_ & ~new_n17151_;
  assign new_n17153_ = pi0198 & ~new_n17152_;
  assign new_n17154_ = ~new_n17132_ & ~new_n17153_;
  assign new_n17155_ = ~pi0603 & ~new_n17154_;
  assign new_n17156_ = pi0621 & new_n17127_;
  assign new_n17157_ = ~pi0198 & ~new_n17156_;
  assign new_n17158_ = pi0621 & new_n17149_;
  assign new_n17159_ = pi0198 & ~new_n17158_;
  assign new_n17160_ = ~new_n17157_ & ~new_n17159_;
  assign new_n17161_ = pi0603 & ~new_n17160_;
  assign new_n17162_ = ~new_n16851_ & ~new_n17161_;
  assign new_n17163_ = ~new_n17155_ & new_n17162_;
  assign new_n17164_ = pi0680 & new_n17163_;
  assign new_n17165_ = ~pi0299 & ~new_n17164_;
  assign new_n17166_ = pi0210 & ~new_n17152_;
  assign new_n17167_ = ~pi0210 & ~new_n17131_;
  assign new_n17168_ = ~new_n17166_ & ~new_n17167_;
  assign new_n17169_ = ~pi0603 & ~new_n17168_;
  assign new_n17170_ = ~pi0210 & ~new_n17156_;
  assign new_n17171_ = pi0210 & ~new_n17158_;
  assign new_n17172_ = ~new_n17170_ & ~new_n17171_;
  assign new_n17173_ = pi0603 & ~new_n17172_;
  assign new_n17174_ = ~new_n16851_ & ~new_n17173_;
  assign new_n17175_ = ~new_n17169_ & new_n17174_;
  assign new_n17176_ = pi0680 & new_n17175_;
  assign new_n17177_ = pi0299 & ~new_n17176_;
  assign new_n17178_ = ~new_n17165_ & ~new_n17177_;
  assign new_n17179_ = pi0140 & ~new_n17178_;
  assign new_n17180_ = ~pi0198 & new_n17129_;
  assign new_n17181_ = pi0198 & new_n17150_;
  assign new_n17182_ = ~new_n17180_ & ~new_n17181_;
  assign new_n17183_ = pi0665 & new_n17149_;
  assign new_n17184_ = pi0198 & ~new_n17183_;
  assign new_n17185_ = pi0665 & new_n17127_;
  assign new_n17186_ = ~pi0198 & ~new_n17185_;
  assign new_n17187_ = ~new_n17184_ & ~new_n17186_;
  assign new_n17188_ = pi0680 & ~new_n17187_;
  assign new_n17189_ = new_n17182_ & ~new_n17188_;
  assign new_n17190_ = ~pi0299 & ~new_n17189_;
  assign new_n17191_ = ~pi0210 & new_n17129_;
  assign new_n17192_ = pi0210 & new_n17150_;
  assign new_n17193_ = ~new_n17191_ & ~new_n17192_;
  assign new_n17194_ = ~pi0210 & ~new_n17185_;
  assign new_n17195_ = pi0210 & ~new_n17183_;
  assign new_n17196_ = ~new_n17194_ & ~new_n17195_;
  assign new_n17197_ = pi0680 & ~new_n17196_;
  assign new_n17198_ = new_n17193_ & ~new_n17197_;
  assign new_n17199_ = pi0299 & ~new_n17198_;
  assign new_n17200_ = ~new_n17190_ & ~new_n17199_;
  assign new_n17201_ = pi0621 & ~new_n17128_;
  assign new_n17202_ = ~new_n17129_ & ~new_n17201_;
  assign new_n17203_ = ~pi0198 & new_n17202_;
  assign new_n17204_ = pi0621 & ~new_n17141_;
  assign new_n17205_ = ~new_n17150_ & ~new_n17204_;
  assign new_n17206_ = pi0198 & new_n17205_;
  assign new_n17207_ = ~new_n17203_ & ~new_n17206_;
  assign new_n17208_ = pi0603 & ~new_n17207_;
  assign new_n17209_ = ~pi0299 & ~new_n17208_;
  assign new_n17210_ = ~pi0210 & ~new_n17202_;
  assign new_n17211_ = pi0210 & ~new_n17205_;
  assign new_n17212_ = ~new_n17210_ & ~new_n17211_;
  assign new_n17213_ = pi0603 & new_n17212_;
  assign new_n17214_ = pi0299 & ~new_n17213_;
  assign new_n17215_ = ~new_n17209_ & ~new_n17214_;
  assign new_n17216_ = pi0680 & new_n17215_;
  assign new_n17217_ = ~new_n17200_ & ~new_n17216_;
  assign new_n17218_ = ~pi0140 & ~new_n17217_;
  assign new_n17219_ = pi0761 & ~new_n17218_;
  assign new_n17220_ = ~new_n17179_ & new_n17219_;
  assign new_n17221_ = ~new_n17173_ & new_n17193_;
  assign new_n17222_ = pi0299 & ~new_n17221_;
  assign new_n17223_ = ~pi0603 & ~new_n17207_;
  assign new_n17224_ = ~new_n17160_ & ~new_n17223_;
  assign new_n17225_ = ~pi0299 & new_n17224_;
  assign new_n17226_ = ~new_n17222_ & ~new_n17225_;
  assign new_n17227_ = new_n17200_ & new_n17226_;
  assign new_n17228_ = ~pi0140 & new_n17227_;
  assign new_n17229_ = pi0680 & new_n17154_;
  assign new_n17230_ = ~pi0299 & ~new_n17229_;
  assign new_n17231_ = pi0680 & new_n17168_;
  assign new_n17232_ = pi0299 & ~new_n17231_;
  assign new_n17233_ = ~new_n17230_ & ~new_n17232_;
  assign new_n17234_ = ~new_n17215_ & ~new_n17233_;
  assign new_n17235_ = pi0140 & new_n17234_;
  assign new_n17236_ = ~pi0761 & ~new_n17235_;
  assign new_n17237_ = ~new_n17228_ & new_n17236_;
  assign new_n17238_ = ~pi0039 & ~new_n17237_;
  assign new_n17239_ = ~new_n17220_ & new_n17238_;
  assign new_n17240_ = ~pi0038 & ~new_n17239_;
  assign new_n17241_ = ~new_n17079_ & new_n17240_;
  assign new_n17242_ = ~pi0140 & ~new_n17035_;
  assign new_n17243_ = pi0140 & ~new_n16917_;
  assign new_n17244_ = new_n3100_ & new_n17243_;
  assign new_n17245_ = ~pi0761 & ~new_n17244_;
  assign new_n17246_ = ~new_n17242_ & new_n17245_;
  assign new_n17247_ = new_n16647_ & new_n16790_;
  assign new_n17248_ = ~pi0140 & ~new_n16647_;
  assign new_n17249_ = pi0761 & ~new_n17248_;
  assign new_n17250_ = ~new_n17247_ & new_n17249_;
  assign new_n17251_ = ~new_n17246_ & ~new_n17250_;
  assign new_n17252_ = ~pi0039 & ~new_n17251_;
  assign new_n17253_ = pi0039 & pi0140;
  assign new_n17254_ = pi0038 & ~new_n17253_;
  assign new_n17255_ = ~new_n17252_ & new_n17254_;
  assign new_n17256_ = ~new_n17241_ & ~new_n17255_;
  assign new_n17257_ = ~pi0738 & ~new_n17256_;
  assign new_n17258_ = pi0299 & ~new_n17193_;
  assign new_n17259_ = ~pi0299 & ~new_n17182_;
  assign new_n17260_ = ~new_n17258_ & ~new_n17259_;
  assign new_n17261_ = ~pi0039 & ~new_n17260_;
  assign new_n17262_ = pi0681 & ~new_n16703_;
  assign new_n17263_ = ~new_n6181_ & ~new_n16693_;
  assign new_n17264_ = new_n6181_ & new_n16660_;
  assign new_n17265_ = ~new_n6185_ & ~new_n17264_;
  assign new_n17266_ = ~new_n17263_ & new_n17265_;
  assign new_n17267_ = ~new_n16700_ & ~new_n17266_;
  assign new_n17268_ = ~pi0661 & ~new_n17267_;
  assign new_n17269_ = pi0661 & new_n16703_;
  assign new_n17270_ = ~pi0681 & ~new_n17269_;
  assign new_n17271_ = ~new_n17268_ & new_n17270_;
  assign new_n17272_ = ~new_n17262_ & ~new_n17271_;
  assign new_n17273_ = ~new_n6238_ & ~new_n17272_;
  assign new_n17274_ = pi0681 & ~new_n16693_;
  assign new_n17275_ = ~pi0616 & ~new_n16630_;
  assign new_n17276_ = new_n16691_ & new_n17275_;
  assign new_n17277_ = ~pi0680 & new_n16692_;
  assign new_n17278_ = pi0680 & ~new_n16687_;
  assign new_n17279_ = ~pi0616 & new_n16630_;
  assign new_n17280_ = ~new_n17278_ & new_n17279_;
  assign new_n17281_ = ~new_n17277_ & new_n17280_;
  assign new_n17282_ = ~new_n17276_ & ~new_n17281_;
  assign new_n17283_ = ~pi0680 & ~new_n16636_;
  assign new_n17284_ = pi0616 & new_n16630_;
  assign new_n17285_ = ~new_n17283_ & new_n17284_;
  assign new_n17286_ = ~new_n17278_ & new_n17285_;
  assign new_n17287_ = pi0616 & new_n16636_;
  assign new_n17288_ = ~new_n16630_ & new_n17287_;
  assign new_n17289_ = ~new_n17286_ & ~new_n17288_;
  assign new_n17290_ = ~pi0681 & new_n17289_;
  assign new_n17291_ = new_n17282_ & new_n17290_;
  assign new_n17292_ = ~new_n17274_ & ~new_n17291_;
  assign new_n17293_ = new_n6238_ & ~new_n17292_;
  assign new_n17294_ = ~new_n17273_ & ~new_n17293_;
  assign new_n17295_ = pi0223 & ~new_n17294_;
  assign new_n17296_ = pi0681 & ~new_n16756_;
  assign new_n17297_ = ~pi0616 & ~new_n16752_;
  assign new_n17298_ = ~pi0614 & ~new_n6183_;
  assign new_n17299_ = ~new_n16683_ & new_n17298_;
  assign new_n17300_ = ~new_n17297_ & new_n17299_;
  assign new_n17301_ = ~pi0614 & new_n6183_;
  assign new_n17302_ = new_n16740_ & new_n17301_;
  assign new_n17303_ = ~new_n17300_ & ~new_n17302_;
  assign new_n17304_ = pi0680 & ~new_n16740_;
  assign new_n17305_ = pi0614 & new_n16630_;
  assign new_n17306_ = ~new_n17283_ & new_n17305_;
  assign new_n17307_ = ~new_n17304_ & new_n17306_;
  assign new_n17308_ = pi0614 & new_n16636_;
  assign new_n17309_ = ~new_n16630_ & new_n17308_;
  assign new_n17310_ = ~new_n17307_ & ~new_n17309_;
  assign new_n17311_ = ~pi0681 & new_n17310_;
  assign new_n17312_ = new_n17303_ & new_n17311_;
  assign new_n17313_ = ~new_n17296_ & ~new_n17312_;
  assign new_n17314_ = new_n6238_ & ~new_n17313_;
  assign new_n17315_ = pi0681 & ~new_n16774_;
  assign new_n17316_ = ~new_n6182_ & new_n16774_;
  assign new_n17317_ = new_n6182_ & ~new_n16738_;
  assign new_n17318_ = ~pi0681 & ~new_n17317_;
  assign new_n17319_ = ~new_n17316_ & new_n17318_;
  assign new_n17320_ = ~new_n17315_ & ~new_n17319_;
  assign new_n17321_ = ~new_n6238_ & ~new_n17320_;
  assign new_n17322_ = ~new_n17314_ & ~new_n17321_;
  assign new_n17323_ = ~new_n3057_ & new_n17322_;
  assign new_n17324_ = ~pi0223 & ~new_n16910_;
  assign new_n17325_ = ~new_n17323_ & new_n17324_;
  assign new_n17326_ = ~new_n17295_ & ~new_n17325_;
  assign new_n17327_ = ~pi0299 & ~new_n17326_;
  assign new_n17328_ = new_n6211_ & ~new_n17313_;
  assign new_n17329_ = ~new_n6211_ & ~new_n17320_;
  assign new_n17330_ = new_n6206_ & ~new_n17329_;
  assign new_n17331_ = ~new_n17328_ & new_n17330_;
  assign new_n17332_ = ~new_n3467_ & new_n17331_;
  assign new_n17333_ = ~new_n6206_ & new_n17320_;
  assign new_n17334_ = ~new_n3467_ & new_n17333_;
  assign new_n17335_ = ~pi0215 & ~new_n16865_;
  assign new_n17336_ = ~new_n17334_ & new_n17335_;
  assign new_n17337_ = ~new_n17332_ & new_n17336_;
  assign new_n17338_ = ~new_n6206_ & new_n17272_;
  assign new_n17339_ = ~new_n6211_ & ~new_n17272_;
  assign new_n17340_ = new_n6211_ & ~new_n17292_;
  assign new_n17341_ = new_n6206_ & ~new_n17340_;
  assign new_n17342_ = ~new_n17339_ & new_n17341_;
  assign new_n17343_ = ~new_n17338_ & ~new_n17342_;
  assign new_n17344_ = pi0215 & new_n17343_;
  assign new_n17345_ = ~new_n17337_ & ~new_n17344_;
  assign new_n17346_ = pi0299 & ~new_n17345_;
  assign new_n17347_ = ~new_n17327_ & ~new_n17346_;
  assign new_n17348_ = pi0039 & ~new_n17347_;
  assign new_n17349_ = ~new_n17261_ & ~new_n17348_;
  assign new_n17350_ = pi0761 & new_n17349_;
  assign new_n17351_ = ~pi0039 & ~new_n17226_;
  assign new_n17352_ = new_n16740_ & ~new_n16850_;
  assign new_n17353_ = new_n6183_ & ~new_n17352_;
  assign new_n17354_ = ~new_n6183_ & new_n17025_;
  assign new_n17355_ = ~new_n17353_ & ~new_n17354_;
  assign new_n17356_ = new_n6212_ & ~new_n17355_;
  assign new_n17357_ = ~pi0603 & new_n16779_;
  assign new_n17358_ = ~new_n16817_ & ~new_n17357_;
  assign new_n17359_ = ~new_n16822_ & new_n17358_;
  assign new_n17360_ = new_n16941_ & ~new_n17359_;
  assign new_n17361_ = ~new_n6212_ & ~new_n17360_;
  assign new_n17362_ = ~new_n3467_ & ~new_n17361_;
  assign new_n17363_ = ~new_n17356_ & new_n17362_;
  assign new_n17364_ = new_n3467_ & new_n16842_;
  assign new_n17365_ = ~new_n17363_ & ~new_n17364_;
  assign new_n17366_ = ~pi0215 & ~new_n17365_;
  assign new_n17367_ = ~new_n16898_ & ~new_n17051_;
  assign new_n17368_ = new_n6212_ & new_n17367_;
  assign new_n17369_ = ~new_n6183_ & ~new_n17043_;
  assign new_n17370_ = ~new_n16660_ & new_n16869_;
  assign new_n17371_ = new_n6183_ & ~new_n17370_;
  assign new_n17372_ = ~new_n17369_ & ~new_n17371_;
  assign new_n17373_ = ~new_n6212_ & ~new_n17372_;
  assign new_n17374_ = pi0215 & ~new_n17373_;
  assign new_n17375_ = ~new_n17368_ & new_n17374_;
  assign new_n17376_ = ~new_n17366_ & ~new_n17375_;
  assign new_n17377_ = pi0299 & ~new_n17376_;
  assign new_n17378_ = new_n6238_ & ~new_n17355_;
  assign new_n17379_ = ~new_n6238_ & ~new_n17360_;
  assign new_n17380_ = ~new_n3057_ & ~new_n17379_;
  assign new_n17381_ = ~new_n17378_ & new_n17380_;
  assign new_n17382_ = new_n3057_ & new_n16842_;
  assign new_n17383_ = ~new_n17381_ & ~new_n17382_;
  assign new_n17384_ = ~pi0223 & ~new_n17383_;
  assign new_n17385_ = new_n6238_ & new_n17367_;
  assign new_n17386_ = ~new_n6238_ & ~new_n17372_;
  assign new_n17387_ = pi0223 & ~new_n17386_;
  assign new_n17388_ = ~new_n17385_ & new_n17387_;
  assign new_n17389_ = ~new_n17384_ & ~new_n17388_;
  assign new_n17390_ = ~pi0299 & ~new_n17389_;
  assign new_n17391_ = ~new_n17377_ & ~new_n17390_;
  assign new_n17392_ = pi0039 & new_n17391_;
  assign new_n17393_ = ~new_n17351_ & ~new_n17392_;
  assign new_n17394_ = ~pi0761 & new_n17393_;
  assign new_n17395_ = ~pi0140 & ~new_n17394_;
  assign new_n17396_ = ~new_n17350_ & new_n17395_;
  assign new_n17397_ = ~pi0039 & ~new_n17215_;
  assign new_n17398_ = ~new_n6212_ & ~new_n16942_;
  assign new_n17399_ = new_n6183_ & new_n16951_;
  assign new_n17400_ = ~new_n6183_ & ~new_n16957_;
  assign new_n17401_ = ~new_n17399_ & ~new_n17400_;
  assign new_n17402_ = new_n6212_ & new_n17401_;
  assign new_n17403_ = ~new_n3467_ & ~new_n17402_;
  assign new_n17404_ = ~new_n17398_ & new_n17403_;
  assign new_n17405_ = new_n3467_ & new_n16635_;
  assign new_n17406_ = new_n16913_ & new_n17405_;
  assign new_n17407_ = ~pi0215 & ~new_n17406_;
  assign new_n17408_ = ~new_n17404_ & new_n17407_;
  assign new_n17409_ = ~new_n6212_ & new_n16701_;
  assign new_n17410_ = ~new_n16978_ & ~new_n17409_;
  assign new_n17411_ = pi0215 & ~new_n17410_;
  assign new_n17412_ = pi0299 & ~new_n17411_;
  assign new_n17413_ = ~new_n17408_ & new_n17412_;
  assign new_n17414_ = ~new_n6238_ & ~new_n16942_;
  assign new_n17415_ = new_n6238_ & new_n17401_;
  assign new_n17416_ = ~new_n3057_ & ~new_n17415_;
  assign new_n17417_ = ~new_n17414_ & new_n17416_;
  assign new_n17418_ = new_n16912_ & ~new_n17417_;
  assign new_n17419_ = ~new_n6238_ & new_n16701_;
  assign new_n17420_ = ~new_n16978_ & ~new_n17419_;
  assign new_n17421_ = pi0223 & ~new_n17420_;
  assign new_n17422_ = ~pi0299 & ~new_n17421_;
  assign new_n17423_ = ~new_n17418_ & new_n17422_;
  assign new_n17424_ = ~new_n17413_ & ~new_n17423_;
  assign new_n17425_ = pi0039 & new_n17424_;
  assign new_n17426_ = ~new_n17397_ & ~new_n17425_;
  assign new_n17427_ = pi0140 & ~pi0761;
  assign new_n17428_ = new_n17426_ & new_n17427_;
  assign new_n17429_ = ~new_n17396_ & ~new_n17428_;
  assign new_n17430_ = ~pi0038 & ~new_n17429_;
  assign new_n17431_ = new_n2754_ & new_n6257_;
  assign new_n17432_ = ~pi0140 & ~new_n17431_;
  assign new_n17433_ = new_n6257_ & new_n16913_;
  assign new_n17434_ = ~pi0761 & new_n17433_;
  assign new_n17435_ = ~new_n17432_ & ~new_n17434_;
  assign new_n17436_ = pi0038 & ~new_n17435_;
  assign new_n17437_ = ~new_n17430_ & ~new_n17436_;
  assign new_n17438_ = pi0738 & ~new_n17437_;
  assign new_n17439_ = new_n3272_ & ~new_n17438_;
  assign new_n17440_ = ~new_n17257_ & new_n17439_;
  assign new_n17441_ = ~new_n16628_ & ~new_n17440_;
  assign new_n17442_ = ~pi0625 & new_n17441_;
  assign new_n17443_ = new_n3272_ & new_n17437_;
  assign new_n17444_ = ~new_n16628_ & ~new_n17443_;
  assign new_n17445_ = pi0625 & new_n17444_;
  assign new_n17446_ = ~pi1153 & ~new_n17445_;
  assign new_n17447_ = ~new_n17442_ & new_n17446_;
  assign new_n17448_ = new_n16910_ & new_n16914_;
  assign new_n17449_ = new_n16774_ & new_n16914_;
  assign new_n17450_ = ~new_n16630_ & new_n17449_;
  assign new_n17451_ = ~new_n16837_ & ~new_n17450_;
  assign new_n17452_ = ~new_n6238_ & new_n17451_;
  assign new_n17453_ = new_n6180_ & new_n16959_;
  assign new_n17454_ = ~new_n16969_ & ~new_n17453_;
  assign new_n17455_ = ~new_n16630_ & new_n17454_;
  assign new_n17456_ = new_n16630_ & ~new_n16959_;
  assign new_n17457_ = pi0680 & ~new_n17456_;
  assign new_n17458_ = ~new_n17455_ & new_n17457_;
  assign new_n17459_ = new_n6238_ & ~new_n17458_;
  assign new_n17460_ = ~new_n3057_ & ~new_n17459_;
  assign new_n17461_ = ~new_n17452_ & new_n17460_;
  assign new_n17462_ = ~new_n17448_ & ~new_n17461_;
  assign new_n17463_ = ~pi0223 & ~new_n17462_;
  assign new_n17464_ = pi0680 & ~new_n16971_;
  assign new_n17465_ = ~new_n17419_ & new_n17464_;
  assign new_n17466_ = pi0223 & ~new_n16979_;
  assign new_n17467_ = new_n17465_ & new_n17466_;
  assign new_n17468_ = ~new_n17463_ & ~new_n17467_;
  assign new_n17469_ = ~pi0299 & ~new_n17468_;
  assign new_n17470_ = new_n6212_ & ~new_n17458_;
  assign new_n17471_ = ~new_n6212_ & new_n17451_;
  assign new_n17472_ = ~new_n3467_ & ~new_n17471_;
  assign new_n17473_ = ~new_n17470_ & new_n17472_;
  assign new_n17474_ = new_n16636_ & new_n16914_;
  assign new_n17475_ = new_n3467_ & new_n17474_;
  assign new_n17476_ = ~new_n17473_ & ~new_n17475_;
  assign new_n17477_ = ~pi0215 & ~new_n17476_;
  assign new_n17478_ = ~new_n17409_ & new_n17464_;
  assign new_n17479_ = pi0215 & ~new_n16979_;
  assign new_n17480_ = new_n17478_ & new_n17479_;
  assign new_n17481_ = ~new_n17477_ & ~new_n17480_;
  assign new_n17482_ = pi0299 & ~new_n17481_;
  assign new_n17483_ = ~new_n17469_ & ~new_n17482_;
  assign new_n17484_ = pi0140 & ~new_n17483_;
  assign new_n17485_ = new_n6180_ & new_n16760_;
  assign new_n17486_ = ~new_n6180_ & new_n16670_;
  assign new_n17487_ = pi0680 & ~new_n17486_;
  assign new_n17488_ = ~new_n17485_ & new_n17487_;
  assign new_n17489_ = ~new_n16757_ & ~new_n17488_;
  assign new_n17490_ = ~new_n16630_ & new_n17489_;
  assign new_n17491_ = pi0680 & ~new_n16760_;
  assign new_n17492_ = new_n16630_ & ~new_n17491_;
  assign new_n17493_ = ~new_n16757_ & new_n17492_;
  assign new_n17494_ = ~new_n17490_ & ~new_n17493_;
  assign new_n17495_ = new_n6238_ & new_n17494_;
  assign new_n17496_ = ~new_n16630_ & ~new_n17013_;
  assign new_n17497_ = new_n16630_ & new_n16758_;
  assign new_n17498_ = pi0680 & ~new_n17497_;
  assign new_n17499_ = ~new_n17496_ & new_n17498_;
  assign new_n17500_ = ~new_n16777_ & ~new_n17499_;
  assign new_n17501_ = ~new_n6238_ & ~new_n17500_;
  assign new_n17502_ = ~new_n3057_ & ~new_n17501_;
  assign new_n17503_ = ~new_n17495_ & new_n17502_;
  assign new_n17504_ = new_n16910_ & ~new_n16914_;
  assign new_n17505_ = ~pi0223 & ~new_n17504_;
  assign new_n17506_ = ~new_n17503_ & new_n17505_;
  assign new_n17507_ = ~new_n16673_ & new_n17487_;
  assign new_n17508_ = ~new_n16695_ & ~new_n17507_;
  assign new_n17509_ = ~new_n17012_ & new_n17045_;
  assign new_n17510_ = ~new_n16704_ & ~new_n17509_;
  assign new_n17511_ = new_n17508_ & new_n17510_;
  assign new_n17512_ = ~new_n6238_ & new_n17511_;
  assign new_n17513_ = ~new_n16694_ & new_n17508_;
  assign new_n17514_ = new_n6238_ & new_n17513_;
  assign new_n17515_ = pi0223 & ~new_n17514_;
  assign new_n17516_ = ~new_n17512_ & new_n17515_;
  assign new_n17517_ = ~new_n17506_ & ~new_n17516_;
  assign new_n17518_ = ~pi0299 & ~new_n17517_;
  assign new_n17519_ = new_n6212_ & new_n17494_;
  assign new_n17520_ = ~new_n6212_ & ~new_n17500_;
  assign new_n17521_ = ~new_n3467_ & ~new_n17520_;
  assign new_n17522_ = ~new_n17519_ & new_n17521_;
  assign new_n17523_ = new_n2754_ & ~new_n16914_;
  assign new_n17524_ = new_n17405_ & new_n17523_;
  assign new_n17525_ = ~pi0215 & ~new_n17524_;
  assign new_n17526_ = ~new_n17522_ & new_n17525_;
  assign new_n17527_ = ~new_n6212_ & new_n17511_;
  assign new_n17528_ = new_n6212_ & new_n17513_;
  assign new_n17529_ = pi0215 & ~new_n17528_;
  assign new_n17530_ = ~new_n17527_ & new_n17529_;
  assign new_n17531_ = ~new_n17526_ & ~new_n17530_;
  assign new_n17532_ = pi0299 & ~new_n17531_;
  assign new_n17533_ = ~new_n17518_ & ~new_n17532_;
  assign new_n17534_ = pi0039 & new_n17533_;
  assign new_n17535_ = ~new_n17253_ & ~new_n17534_;
  assign new_n17536_ = ~new_n17484_ & ~new_n17535_;
  assign new_n17537_ = ~pi0140 & ~new_n17200_;
  assign new_n17538_ = pi0140 & new_n17233_;
  assign new_n17539_ = ~pi0039 & ~new_n17538_;
  assign new_n17540_ = ~new_n17537_ & new_n17539_;
  assign new_n17541_ = ~new_n17536_ & ~new_n17540_;
  assign new_n17542_ = ~pi0038 & ~new_n17541_;
  assign new_n17543_ = new_n6257_ & new_n16915_;
  assign new_n17544_ = pi0038 & ~new_n17543_;
  assign new_n17545_ = ~new_n17432_ & new_n17544_;
  assign new_n17546_ = ~pi0738 & ~new_n17545_;
  assign new_n17547_ = ~new_n17542_ & new_n17546_;
  assign new_n17548_ = ~pi0038 & ~new_n17349_;
  assign new_n17549_ = new_n2754_ & new_n6132_;
  assign new_n17550_ = pi0038 & ~new_n17549_;
  assign new_n17551_ = ~new_n17548_ & ~new_n17550_;
  assign new_n17552_ = ~pi0140 & pi0738;
  assign new_n17553_ = ~new_n17551_ & new_n17552_;
  assign new_n17554_ = new_n3272_ & ~new_n17553_;
  assign new_n17555_ = ~new_n17547_ & new_n17554_;
  assign new_n17556_ = ~new_n16628_ & ~new_n17555_;
  assign new_n17557_ = pi0625 & new_n17556_;
  assign new_n17558_ = new_n3272_ & new_n17551_;
  assign new_n17559_ = ~pi0140 & ~new_n17558_;
  assign new_n17560_ = ~pi0625 & new_n17559_;
  assign new_n17561_ = pi1153 & ~new_n17560_;
  assign new_n17562_ = ~new_n17557_ & new_n17561_;
  assign new_n17563_ = ~pi0608 & ~new_n17562_;
  assign new_n17564_ = ~new_n17447_ & new_n17563_;
  assign new_n17565_ = pi0625 & new_n17441_;
  assign new_n17566_ = ~pi0625 & new_n17444_;
  assign new_n17567_ = pi1153 & ~new_n17566_;
  assign new_n17568_ = ~new_n17565_ & new_n17567_;
  assign new_n17569_ = ~pi0625 & new_n17556_;
  assign new_n17570_ = pi0625 & new_n17559_;
  assign new_n17571_ = ~pi1153 & ~new_n17570_;
  assign new_n17572_ = ~new_n17569_ & new_n17571_;
  assign new_n17573_ = pi0608 & ~new_n17572_;
  assign new_n17574_ = ~new_n17568_ & new_n17573_;
  assign new_n17575_ = ~new_n17564_ & ~new_n17574_;
  assign new_n17576_ = pi0778 & ~new_n17575_;
  assign new_n17577_ = ~pi0778 & new_n17441_;
  assign new_n17578_ = ~new_n17576_ & ~new_n17577_;
  assign new_n17579_ = ~pi0609 & ~new_n17578_;
  assign new_n17580_ = ~pi0778 & ~new_n17556_;
  assign new_n17581_ = ~new_n17562_ & ~new_n17572_;
  assign new_n17582_ = pi0778 & ~new_n17581_;
  assign new_n17583_ = ~new_n17580_ & ~new_n17582_;
  assign new_n17584_ = pi0609 & new_n17583_;
  assign new_n17585_ = ~pi1155 & ~new_n17584_;
  assign new_n17586_ = ~new_n17579_ & new_n17585_;
  assign new_n17587_ = ~pi0608 & pi1153;
  assign new_n17588_ = pi0608 & ~pi1153;
  assign new_n17589_ = ~new_n17587_ & ~new_n17588_;
  assign new_n17590_ = pi0778 & ~new_n17589_;
  assign new_n17591_ = pi0609 & ~new_n17590_;
  assign new_n17592_ = ~new_n17559_ & ~new_n17591_;
  assign new_n17593_ = ~new_n17444_ & ~new_n17590_;
  assign new_n17594_ = pi0609 & new_n17593_;
  assign new_n17595_ = ~new_n17592_ & ~new_n17594_;
  assign new_n17596_ = pi1155 & ~new_n17595_;
  assign new_n17597_ = ~pi0660 & ~new_n17596_;
  assign new_n17598_ = ~new_n17586_ & new_n17597_;
  assign new_n17599_ = pi0609 & ~new_n17578_;
  assign new_n17600_ = ~pi0609 & new_n17583_;
  assign new_n17601_ = pi1155 & ~new_n17600_;
  assign new_n17602_ = ~new_n17599_ & new_n17601_;
  assign new_n17603_ = ~pi0609 & ~new_n17590_;
  assign new_n17604_ = ~new_n17559_ & ~new_n17603_;
  assign new_n17605_ = ~pi0609 & new_n17593_;
  assign new_n17606_ = ~new_n17604_ & ~new_n17605_;
  assign new_n17607_ = ~pi1155 & ~new_n17606_;
  assign new_n17608_ = pi0660 & ~new_n17607_;
  assign new_n17609_ = ~new_n17602_ & new_n17608_;
  assign new_n17610_ = ~new_n17598_ & ~new_n17609_;
  assign new_n17611_ = pi0785 & ~new_n17610_;
  assign new_n17612_ = ~pi0785 & ~new_n17578_;
  assign new_n17613_ = ~new_n17611_ & ~new_n17612_;
  assign new_n17614_ = ~pi0618 & ~new_n17613_;
  assign new_n17615_ = ~pi0660 & ~pi1155;
  assign new_n17616_ = pi0660 & pi1155;
  assign new_n17617_ = pi0785 & ~new_n17616_;
  assign new_n17618_ = ~new_n17615_ & new_n17617_;
  assign new_n17619_ = ~new_n17583_ & ~new_n17618_;
  assign new_n17620_ = ~new_n17559_ & new_n17618_;
  assign new_n17621_ = ~new_n17619_ & ~new_n17620_;
  assign new_n17622_ = pi0618 & new_n17621_;
  assign new_n17623_ = ~pi1154 & ~new_n17622_;
  assign new_n17624_ = ~new_n17614_ & new_n17623_;
  assign new_n17625_ = ~new_n17559_ & new_n17590_;
  assign new_n17626_ = ~new_n17593_ & ~new_n17625_;
  assign new_n17627_ = ~pi0785 & ~new_n17626_;
  assign new_n17628_ = ~new_n17596_ & ~new_n17607_;
  assign new_n17629_ = pi0785 & ~new_n17628_;
  assign new_n17630_ = ~new_n17627_ & ~new_n17629_;
  assign new_n17631_ = pi0618 & new_n17630_;
  assign new_n17632_ = ~pi0618 & new_n17559_;
  assign new_n17633_ = pi1154 & ~new_n17632_;
  assign new_n17634_ = ~new_n17631_ & new_n17633_;
  assign new_n17635_ = ~pi0627 & ~new_n17634_;
  assign new_n17636_ = ~new_n17624_ & new_n17635_;
  assign new_n17637_ = pi0618 & ~new_n17613_;
  assign new_n17638_ = ~pi0618 & new_n17621_;
  assign new_n17639_ = pi1154 & ~new_n17638_;
  assign new_n17640_ = ~new_n17637_ & new_n17639_;
  assign new_n17641_ = ~pi0618 & new_n17630_;
  assign new_n17642_ = pi0618 & new_n17559_;
  assign new_n17643_ = ~pi1154 & ~new_n17642_;
  assign new_n17644_ = ~new_n17641_ & new_n17643_;
  assign new_n17645_ = pi0627 & ~new_n17644_;
  assign new_n17646_ = ~new_n17640_ & new_n17645_;
  assign new_n17647_ = ~new_n17636_ & ~new_n17646_;
  assign new_n17648_ = pi0781 & ~new_n17647_;
  assign new_n17649_ = ~pi0781 & ~new_n17613_;
  assign new_n17650_ = ~new_n17648_ & ~new_n17649_;
  assign new_n17651_ = ~pi0619 & ~new_n17650_;
  assign new_n17652_ = ~pi0627 & ~pi1154;
  assign new_n17653_ = pi0627 & pi1154;
  assign new_n17654_ = pi0781 & ~new_n17653_;
  assign new_n17655_ = ~new_n17652_ & new_n17654_;
  assign new_n17656_ = new_n17621_ & ~new_n17655_;
  assign new_n17657_ = new_n17559_ & new_n17655_;
  assign new_n17658_ = ~new_n17656_ & ~new_n17657_;
  assign new_n17659_ = pi0619 & ~new_n17658_;
  assign new_n17660_ = ~pi1159 & ~new_n17659_;
  assign new_n17661_ = ~new_n17651_ & new_n17660_;
  assign new_n17662_ = ~pi0781 & ~new_n17630_;
  assign new_n17663_ = ~new_n17634_ & ~new_n17644_;
  assign new_n17664_ = pi0781 & ~new_n17663_;
  assign new_n17665_ = ~new_n17662_ & ~new_n17664_;
  assign new_n17666_ = pi0619 & new_n17665_;
  assign new_n17667_ = ~pi0619 & new_n17559_;
  assign new_n17668_ = pi1159 & ~new_n17667_;
  assign new_n17669_ = ~new_n17666_ & new_n17668_;
  assign new_n17670_ = ~pi0648 & ~new_n17669_;
  assign new_n17671_ = ~new_n17661_ & new_n17670_;
  assign new_n17672_ = pi0619 & ~new_n17650_;
  assign new_n17673_ = ~pi0619 & ~new_n17658_;
  assign new_n17674_ = pi1159 & ~new_n17673_;
  assign new_n17675_ = ~new_n17672_ & new_n17674_;
  assign new_n17676_ = ~pi0619 & new_n17665_;
  assign new_n17677_ = pi0619 & new_n17559_;
  assign new_n17678_ = ~pi1159 & ~new_n17677_;
  assign new_n17679_ = ~new_n17676_ & new_n17678_;
  assign new_n17680_ = pi0648 & ~new_n17679_;
  assign new_n17681_ = ~new_n17675_ & new_n17680_;
  assign new_n17682_ = ~new_n17671_ & ~new_n17681_;
  assign new_n17683_ = pi0789 & ~new_n17682_;
  assign new_n17684_ = ~pi0789 & ~new_n17650_;
  assign new_n17685_ = ~new_n17683_ & ~new_n17684_;
  assign new_n17686_ = ~pi0788 & new_n17685_;
  assign new_n17687_ = ~pi0626 & new_n17685_;
  assign new_n17688_ = ~pi0648 & pi1159;
  assign new_n17689_ = pi0648 & ~pi1159;
  assign new_n17690_ = ~new_n17688_ & ~new_n17689_;
  assign new_n17691_ = pi0789 & ~new_n17690_;
  assign new_n17692_ = new_n17658_ & ~new_n17691_;
  assign new_n17693_ = ~new_n17559_ & new_n17691_;
  assign new_n17694_ = ~new_n17692_ & ~new_n17693_;
  assign new_n17695_ = pi0626 & ~new_n17694_;
  assign new_n17696_ = ~pi0641 & ~new_n17695_;
  assign new_n17697_ = ~new_n17687_ & new_n17696_;
  assign new_n17698_ = ~pi0641 & ~pi1158;
  assign new_n17699_ = ~pi0789 & ~new_n17665_;
  assign new_n17700_ = ~new_n17669_ & ~new_n17679_;
  assign new_n17701_ = pi0789 & ~new_n17700_;
  assign new_n17702_ = ~new_n17699_ & ~new_n17701_;
  assign new_n17703_ = ~pi0626 & new_n17702_;
  assign new_n17704_ = pi0626 & new_n17559_;
  assign new_n17705_ = ~pi1158 & ~new_n17704_;
  assign new_n17706_ = ~new_n17703_ & new_n17705_;
  assign new_n17707_ = ~new_n17698_ & ~new_n17706_;
  assign new_n17708_ = ~new_n17697_ & ~new_n17707_;
  assign new_n17709_ = pi0626 & new_n17685_;
  assign new_n17710_ = ~pi0626 & ~new_n17694_;
  assign new_n17711_ = pi0641 & ~new_n17710_;
  assign new_n17712_ = ~new_n17709_ & new_n17711_;
  assign new_n17713_ = pi0641 & pi1158;
  assign new_n17714_ = pi0626 & new_n17702_;
  assign new_n17715_ = ~pi0626 & new_n17559_;
  assign new_n17716_ = pi1158 & ~new_n17715_;
  assign new_n17717_ = ~new_n17714_ & new_n17716_;
  assign new_n17718_ = ~new_n17713_ & ~new_n17717_;
  assign new_n17719_ = ~new_n17712_ & ~new_n17718_;
  assign new_n17720_ = ~new_n17708_ & ~new_n17719_;
  assign new_n17721_ = pi0788 & ~new_n17720_;
  assign new_n17722_ = ~new_n17686_ & ~new_n17721_;
  assign new_n17723_ = ~pi0628 & new_n17722_;
  assign new_n17724_ = ~new_n17706_ & ~new_n17717_;
  assign new_n17725_ = pi0788 & ~new_n17724_;
  assign new_n17726_ = ~pi0788 & ~new_n17702_;
  assign new_n17727_ = ~new_n17725_ & ~new_n17726_;
  assign new_n17728_ = pi0628 & new_n17727_;
  assign new_n17729_ = ~pi1156 & ~new_n17728_;
  assign new_n17730_ = ~new_n17723_ & new_n17729_;
  assign new_n17731_ = ~pi0641 & pi1158;
  assign new_n17732_ = pi0641 & ~pi1158;
  assign new_n17733_ = ~new_n17731_ & ~new_n17732_;
  assign new_n17734_ = pi0788 & ~new_n17733_;
  assign new_n17735_ = new_n17694_ & ~new_n17734_;
  assign new_n17736_ = new_n17559_ & new_n17734_;
  assign new_n17737_ = ~new_n17735_ & ~new_n17736_;
  assign new_n17738_ = pi0628 & ~new_n17737_;
  assign new_n17739_ = ~pi0628 & new_n17559_;
  assign new_n17740_ = pi1156 & ~new_n17739_;
  assign new_n17741_ = ~new_n17738_ & new_n17740_;
  assign new_n17742_ = ~pi0629 & ~new_n17741_;
  assign new_n17743_ = ~new_n17730_ & new_n17742_;
  assign new_n17744_ = pi0628 & new_n17722_;
  assign new_n17745_ = ~pi0628 & new_n17727_;
  assign new_n17746_ = pi1156 & ~new_n17745_;
  assign new_n17747_ = ~new_n17744_ & new_n17746_;
  assign new_n17748_ = ~pi0628 & ~new_n17737_;
  assign new_n17749_ = pi0628 & new_n17559_;
  assign new_n17750_ = ~pi1156 & ~new_n17749_;
  assign new_n17751_ = ~new_n17748_ & new_n17750_;
  assign new_n17752_ = pi0629 & ~new_n17751_;
  assign new_n17753_ = ~new_n17747_ & new_n17752_;
  assign new_n17754_ = ~new_n17743_ & ~new_n17753_;
  assign new_n17755_ = pi0792 & ~new_n17754_;
  assign new_n17756_ = ~pi0792 & new_n17722_;
  assign new_n17757_ = ~new_n17755_ & ~new_n17756_;
  assign new_n17758_ = ~pi0647 & ~new_n17757_;
  assign new_n17759_ = ~pi0629 & pi1156;
  assign new_n17760_ = pi0629 & ~pi1156;
  assign new_n17761_ = ~new_n17759_ & ~new_n17760_;
  assign new_n17762_ = pi0792 & ~new_n17761_;
  assign new_n17763_ = new_n17727_ & ~new_n17762_;
  assign new_n17764_ = new_n17559_ & new_n17762_;
  assign new_n17765_ = ~new_n17763_ & ~new_n17764_;
  assign new_n17766_ = pi0647 & ~new_n17765_;
  assign new_n17767_ = ~pi1157 & ~new_n17766_;
  assign new_n17768_ = ~new_n17758_ & new_n17767_;
  assign new_n17769_ = ~pi0792 & new_n17737_;
  assign new_n17770_ = ~new_n17741_ & ~new_n17751_;
  assign new_n17771_ = pi0792 & ~new_n17770_;
  assign new_n17772_ = ~new_n17769_ & ~new_n17771_;
  assign new_n17773_ = pi0647 & new_n17772_;
  assign new_n17774_ = ~pi0647 & new_n17559_;
  assign new_n17775_ = pi1157 & ~new_n17774_;
  assign new_n17776_ = ~new_n17773_ & new_n17775_;
  assign new_n17777_ = ~pi0630 & ~new_n17776_;
  assign new_n17778_ = ~new_n17768_ & new_n17777_;
  assign new_n17779_ = pi0647 & ~new_n17757_;
  assign new_n17780_ = ~pi0647 & ~new_n17765_;
  assign new_n17781_ = pi1157 & ~new_n17780_;
  assign new_n17782_ = ~new_n17779_ & new_n17781_;
  assign new_n17783_ = ~pi0647 & new_n17772_;
  assign new_n17784_ = pi0647 & new_n17559_;
  assign new_n17785_ = ~pi1157 & ~new_n17784_;
  assign new_n17786_ = ~new_n17783_ & new_n17785_;
  assign new_n17787_ = pi0630 & ~new_n17786_;
  assign new_n17788_ = ~new_n17782_ & new_n17787_;
  assign new_n17789_ = ~new_n17778_ & ~new_n17788_;
  assign new_n17790_ = pi0787 & ~new_n17789_;
  assign new_n17791_ = ~pi0787 & ~new_n17757_;
  assign new_n17792_ = ~new_n17790_ & ~new_n17791_;
  assign new_n17793_ = ~pi0644 & ~new_n17792_;
  assign new_n17794_ = ~pi0787 & ~new_n17772_;
  assign new_n17795_ = ~new_n17776_ & ~new_n17786_;
  assign new_n17796_ = pi0787 & ~new_n17795_;
  assign new_n17797_ = ~new_n17794_ & ~new_n17796_;
  assign new_n17798_ = pi0644 & new_n17797_;
  assign new_n17799_ = ~pi0715 & ~new_n17798_;
  assign new_n17800_ = ~new_n17793_ & new_n17799_;
  assign new_n17801_ = ~pi0630 & pi1157;
  assign new_n17802_ = pi0630 & ~pi1157;
  assign new_n17803_ = ~new_n17801_ & ~new_n17802_;
  assign new_n17804_ = pi0787 & ~new_n17803_;
  assign new_n17805_ = new_n17765_ & ~new_n17804_;
  assign new_n17806_ = ~new_n17559_ & new_n17804_;
  assign new_n17807_ = ~new_n17805_ & ~new_n17806_;
  assign new_n17808_ = ~pi0644 & new_n17807_;
  assign new_n17809_ = pi0644 & new_n17559_;
  assign new_n17810_ = pi0715 & ~new_n17809_;
  assign new_n17811_ = ~new_n17808_ & new_n17810_;
  assign new_n17812_ = ~pi1160 & ~new_n17811_;
  assign new_n17813_ = ~new_n17800_ & new_n17812_;
  assign new_n17814_ = pi0644 & ~new_n17792_;
  assign new_n17815_ = ~pi0644 & new_n17797_;
  assign new_n17816_ = pi0715 & ~new_n17815_;
  assign new_n17817_ = ~new_n17814_ & new_n17816_;
  assign new_n17818_ = pi0644 & new_n17807_;
  assign new_n17819_ = ~pi0644 & new_n17559_;
  assign new_n17820_ = ~pi0715 & ~new_n17819_;
  assign new_n17821_ = ~new_n17818_ & new_n17820_;
  assign new_n17822_ = pi1160 & ~new_n17821_;
  assign new_n17823_ = ~new_n17817_ & new_n17822_;
  assign new_n17824_ = pi0790 & ~new_n17823_;
  assign new_n17825_ = ~new_n17813_ & new_n17824_;
  assign new_n17826_ = ~pi0790 & new_n17792_;
  assign new_n17827_ = ~po1038 & ~new_n17826_;
  assign new_n17828_ = ~new_n17825_ & new_n17827_;
  assign new_n17829_ = ~pi0140 & po1038;
  assign new_n17830_ = ~pi0832 & ~new_n17829_;
  assign new_n17831_ = ~new_n17828_ & new_n17830_;
  assign new_n17832_ = ~pi0140 & ~new_n2754_;
  assign new_n17833_ = ~pi0738 & new_n16915_;
  assign new_n17834_ = ~new_n17832_ & ~new_n17833_;
  assign new_n17835_ = ~pi0778 & new_n17834_;
  assign new_n17836_ = ~pi0625 & new_n17833_;
  assign new_n17837_ = ~new_n17834_ & ~new_n17836_;
  assign new_n17838_ = pi1153 & ~new_n17837_;
  assign new_n17839_ = ~pi1153 & ~new_n17832_;
  assign new_n17840_ = ~new_n17836_ & new_n17839_;
  assign new_n17841_ = ~new_n17838_ & ~new_n17840_;
  assign new_n17842_ = pi0778 & ~new_n17841_;
  assign new_n17843_ = ~new_n17835_ & ~new_n17842_;
  assign new_n17844_ = new_n2754_ & new_n17618_;
  assign new_n17845_ = new_n17843_ & ~new_n17844_;
  assign new_n17846_ = new_n2754_ & new_n17655_;
  assign new_n17847_ = new_n17845_ & ~new_n17846_;
  assign new_n17848_ = new_n2754_ & new_n17691_;
  assign new_n17849_ = new_n17847_ & ~new_n17848_;
  assign new_n17850_ = ~pi0626 & pi1158;
  assign new_n17851_ = pi0626 & ~pi1158;
  assign new_n17852_ = ~new_n17850_ & ~new_n17851_;
  assign new_n17853_ = ~pi0626 & pi0641;
  assign new_n17854_ = pi0626 & ~pi0641;
  assign new_n17855_ = ~new_n17853_ & ~new_n17854_;
  assign new_n17856_ = ~new_n17852_ & ~new_n17855_;
  assign new_n17857_ = new_n17849_ & new_n17856_;
  assign new_n17858_ = new_n2754_ & new_n17590_;
  assign new_n17859_ = ~pi0761 & new_n16913_;
  assign new_n17860_ = ~new_n17832_ & ~new_n17859_;
  assign new_n17861_ = ~new_n17858_ & ~new_n17860_;
  assign new_n17862_ = ~pi0785 & ~new_n17861_;
  assign new_n17863_ = new_n2754_ & ~new_n17591_;
  assign new_n17864_ = ~new_n17860_ & ~new_n17863_;
  assign new_n17865_ = pi1155 & ~new_n17864_;
  assign new_n17866_ = pi0609 & new_n2754_;
  assign new_n17867_ = new_n17861_ & ~new_n17866_;
  assign new_n17868_ = ~pi1155 & ~new_n17867_;
  assign new_n17869_ = ~new_n17865_ & ~new_n17868_;
  assign new_n17870_ = pi0785 & ~new_n17869_;
  assign new_n17871_ = ~new_n17862_ & ~new_n17870_;
  assign new_n17872_ = ~pi0781 & ~new_n17871_;
  assign new_n17873_ = ~pi0618 & new_n2754_;
  assign new_n17874_ = new_n17871_ & ~new_n17873_;
  assign new_n17875_ = pi1154 & ~new_n17874_;
  assign new_n17876_ = pi0618 & new_n2754_;
  assign new_n17877_ = new_n17871_ & ~new_n17876_;
  assign new_n17878_ = ~pi1154 & ~new_n17877_;
  assign new_n17879_ = ~new_n17875_ & ~new_n17878_;
  assign new_n17880_ = pi0781 & ~new_n17879_;
  assign new_n17881_ = ~new_n17872_ & ~new_n17880_;
  assign new_n17882_ = ~pi0789 & ~new_n17881_;
  assign new_n17883_ = pi0619 & new_n17881_;
  assign new_n17884_ = ~pi0619 & new_n17832_;
  assign new_n17885_ = pi1159 & ~new_n17884_;
  assign new_n17886_ = ~new_n17883_ & new_n17885_;
  assign new_n17887_ = ~pi0619 & new_n17881_;
  assign new_n17888_ = pi0619 & new_n17832_;
  assign new_n17889_ = ~pi1159 & ~new_n17888_;
  assign new_n17890_ = ~new_n17887_ & new_n17889_;
  assign new_n17891_ = ~new_n17886_ & ~new_n17890_;
  assign new_n17892_ = pi0789 & ~new_n17891_;
  assign new_n17893_ = ~new_n17882_ & ~new_n17892_;
  assign new_n17894_ = pi0626 & new_n17893_;
  assign new_n17895_ = ~pi0626 & new_n17832_;
  assign new_n17896_ = pi1158 & ~new_n17895_;
  assign new_n17897_ = ~new_n17894_ & new_n17896_;
  assign new_n17898_ = ~pi0626 & new_n17893_;
  assign new_n17899_ = pi0626 & new_n17832_;
  assign new_n17900_ = ~pi1158 & ~new_n17899_;
  assign new_n17901_ = ~new_n17898_ & new_n17900_;
  assign new_n17902_ = ~new_n17897_ & ~new_n17901_;
  assign new_n17903_ = ~new_n17733_ & new_n17902_;
  assign new_n17904_ = ~new_n17857_ & ~new_n17903_;
  assign new_n17905_ = pi0788 & ~new_n17904_;
  assign new_n17906_ = ~new_n16639_ & ~new_n17834_;
  assign new_n17907_ = pi0625 & new_n17906_;
  assign new_n17908_ = new_n17860_ & ~new_n17906_;
  assign new_n17909_ = ~new_n17907_ & ~new_n17908_;
  assign new_n17910_ = new_n17839_ & ~new_n17909_;
  assign new_n17911_ = ~pi0608 & ~new_n17838_;
  assign new_n17912_ = ~new_n17910_ & new_n17911_;
  assign new_n17913_ = pi1153 & new_n17860_;
  assign new_n17914_ = ~new_n17907_ & new_n17913_;
  assign new_n17915_ = pi0608 & ~new_n17840_;
  assign new_n17916_ = ~new_n17914_ & new_n17915_;
  assign new_n17917_ = ~new_n17912_ & ~new_n17916_;
  assign new_n17918_ = pi0778 & ~new_n17917_;
  assign new_n17919_ = ~pi0778 & ~new_n17908_;
  assign new_n17920_ = ~new_n17918_ & ~new_n17919_;
  assign new_n17921_ = ~pi0609 & ~new_n17920_;
  assign new_n17922_ = pi0609 & new_n17843_;
  assign new_n17923_ = ~pi1155 & ~new_n17922_;
  assign new_n17924_ = ~new_n17921_ & new_n17923_;
  assign new_n17925_ = ~pi0660 & ~new_n17865_;
  assign new_n17926_ = ~new_n17924_ & new_n17925_;
  assign new_n17927_ = pi0609 & ~new_n17920_;
  assign new_n17928_ = ~pi0609 & new_n17843_;
  assign new_n17929_ = pi1155 & ~new_n17928_;
  assign new_n17930_ = ~new_n17927_ & new_n17929_;
  assign new_n17931_ = pi0660 & ~new_n17868_;
  assign new_n17932_ = ~new_n17930_ & new_n17931_;
  assign new_n17933_ = ~new_n17926_ & ~new_n17932_;
  assign new_n17934_ = pi0785 & ~new_n17933_;
  assign new_n17935_ = ~pi0785 & ~new_n17920_;
  assign new_n17936_ = ~new_n17934_ & ~new_n17935_;
  assign new_n17937_ = ~pi0618 & ~new_n17936_;
  assign new_n17938_ = pi0618 & new_n17845_;
  assign new_n17939_ = ~pi1154 & ~new_n17938_;
  assign new_n17940_ = ~new_n17937_ & new_n17939_;
  assign new_n17941_ = ~pi0627 & ~new_n17875_;
  assign new_n17942_ = ~new_n17940_ & new_n17941_;
  assign new_n17943_ = pi0618 & ~new_n17936_;
  assign new_n17944_ = ~pi0618 & new_n17845_;
  assign new_n17945_ = pi1154 & ~new_n17944_;
  assign new_n17946_ = ~new_n17943_ & new_n17945_;
  assign new_n17947_ = pi0627 & ~new_n17878_;
  assign new_n17948_ = ~new_n17946_ & new_n17947_;
  assign new_n17949_ = ~new_n17942_ & ~new_n17948_;
  assign new_n17950_ = pi0781 & ~new_n17949_;
  assign new_n17951_ = ~pi0781 & ~new_n17936_;
  assign new_n17952_ = ~new_n17950_ & ~new_n17951_;
  assign new_n17953_ = pi0619 & ~new_n17952_;
  assign new_n17954_ = ~pi0619 & new_n17847_;
  assign new_n17955_ = pi1159 & ~new_n17954_;
  assign new_n17956_ = ~new_n17953_ & new_n17955_;
  assign new_n17957_ = pi0648 & ~new_n17890_;
  assign new_n17958_ = ~new_n17956_ & new_n17957_;
  assign new_n17959_ = ~pi0619 & ~new_n17952_;
  assign new_n17960_ = pi0619 & new_n17847_;
  assign new_n17961_ = ~pi1159 & ~new_n17960_;
  assign new_n17962_ = ~new_n17959_ & new_n17961_;
  assign new_n17963_ = ~pi0648 & ~new_n17886_;
  assign new_n17964_ = ~new_n17962_ & new_n17963_;
  assign new_n17965_ = pi0789 & ~new_n17964_;
  assign new_n17966_ = ~new_n17958_ & new_n17965_;
  assign new_n17967_ = ~pi0789 & new_n17952_;
  assign new_n17968_ = pi0788 & ~new_n17852_;
  assign new_n17969_ = ~new_n17734_ & ~new_n17968_;
  assign new_n17970_ = ~new_n17967_ & new_n17969_;
  assign new_n17971_ = ~new_n17966_ & new_n17970_;
  assign new_n17972_ = ~new_n17905_ & ~new_n17971_;
  assign new_n17973_ = ~pi0628 & ~new_n17972_;
  assign new_n17974_ = ~pi0788 & ~new_n17893_;
  assign new_n17975_ = pi0788 & ~new_n17902_;
  assign new_n17976_ = ~new_n17974_ & ~new_n17975_;
  assign new_n17977_ = pi0628 & new_n17976_;
  assign new_n17978_ = ~pi1156 & ~new_n17977_;
  assign new_n17979_ = ~new_n17973_ & new_n17978_;
  assign new_n17980_ = new_n2754_ & new_n17734_;
  assign new_n17981_ = new_n17849_ & ~new_n17980_;
  assign new_n17982_ = ~pi0628 & new_n2754_;
  assign new_n17983_ = new_n17981_ & ~new_n17982_;
  assign new_n17984_ = pi1156 & ~new_n17983_;
  assign new_n17985_ = ~pi0629 & ~new_n17984_;
  assign new_n17986_ = ~new_n17979_ & new_n17985_;
  assign new_n17987_ = pi0628 & ~new_n17972_;
  assign new_n17988_ = ~pi0628 & new_n17976_;
  assign new_n17989_ = pi1156 & ~new_n17988_;
  assign new_n17990_ = ~new_n17987_ & new_n17989_;
  assign new_n17991_ = pi0628 & new_n2754_;
  assign new_n17992_ = new_n17981_ & ~new_n17991_;
  assign new_n17993_ = ~pi1156 & ~new_n17992_;
  assign new_n17994_ = pi0629 & ~new_n17993_;
  assign new_n17995_ = ~new_n17990_ & new_n17994_;
  assign new_n17996_ = ~new_n17986_ & ~new_n17995_;
  assign new_n17997_ = pi0792 & ~new_n17996_;
  assign new_n17998_ = ~pi0792 & ~new_n17972_;
  assign new_n17999_ = ~new_n17997_ & ~new_n17998_;
  assign new_n18000_ = ~pi0647 & ~new_n17999_;
  assign new_n18001_ = ~new_n17762_ & new_n17976_;
  assign new_n18002_ = new_n17762_ & new_n17832_;
  assign new_n18003_ = ~new_n18001_ & ~new_n18002_;
  assign new_n18004_ = pi0647 & ~new_n18003_;
  assign new_n18005_ = ~pi1157 & ~new_n18004_;
  assign new_n18006_ = ~new_n18000_ & new_n18005_;
  assign new_n18007_ = ~pi0628 & pi1156;
  assign new_n18008_ = pi0628 & ~pi1156;
  assign new_n18009_ = ~new_n18007_ & ~new_n18008_;
  assign new_n18010_ = pi0792 & ~new_n18009_;
  assign new_n18011_ = new_n2754_ & new_n18010_;
  assign new_n18012_ = new_n17981_ & ~new_n18011_;
  assign new_n18013_ = pi0647 & new_n18012_;
  assign new_n18014_ = ~pi0647 & new_n17832_;
  assign new_n18015_ = pi1157 & ~new_n18014_;
  assign new_n18016_ = ~new_n18013_ & new_n18015_;
  assign new_n18017_ = ~pi0630 & ~new_n18016_;
  assign new_n18018_ = ~new_n18006_ & new_n18017_;
  assign new_n18019_ = pi0647 & ~new_n17999_;
  assign new_n18020_ = ~pi0647 & ~new_n18003_;
  assign new_n18021_ = pi1157 & ~new_n18020_;
  assign new_n18022_ = ~new_n18019_ & new_n18021_;
  assign new_n18023_ = ~pi0647 & new_n18012_;
  assign new_n18024_ = pi0647 & new_n17832_;
  assign new_n18025_ = ~pi1157 & ~new_n18024_;
  assign new_n18026_ = ~new_n18023_ & new_n18025_;
  assign new_n18027_ = pi0630 & ~new_n18026_;
  assign new_n18028_ = ~new_n18022_ & new_n18027_;
  assign new_n18029_ = ~new_n18018_ & ~new_n18028_;
  assign new_n18030_ = pi0787 & ~new_n18029_;
  assign new_n18031_ = ~pi0787 & ~new_n17999_;
  assign new_n18032_ = ~new_n18030_ & ~new_n18031_;
  assign new_n18033_ = pi0644 & ~new_n18032_;
  assign new_n18034_ = ~pi0787 & ~new_n18012_;
  assign new_n18035_ = ~new_n18016_ & ~new_n18026_;
  assign new_n18036_ = pi0787 & ~new_n18035_;
  assign new_n18037_ = ~new_n18034_ & ~new_n18036_;
  assign new_n18038_ = ~pi0644 & new_n18037_;
  assign new_n18039_ = pi0715 & ~new_n18038_;
  assign new_n18040_ = ~new_n18033_ & new_n18039_;
  assign new_n18041_ = new_n17804_ & ~new_n17832_;
  assign new_n18042_ = ~new_n17804_ & new_n18003_;
  assign new_n18043_ = ~new_n18041_ & ~new_n18042_;
  assign new_n18044_ = pi0644 & new_n18043_;
  assign new_n18045_ = ~pi0644 & new_n17832_;
  assign new_n18046_ = ~pi0715 & ~new_n18045_;
  assign new_n18047_ = ~new_n18044_ & new_n18046_;
  assign new_n18048_ = pi1160 & ~new_n18047_;
  assign new_n18049_ = ~new_n18040_ & new_n18048_;
  assign new_n18050_ = ~pi0644 & ~new_n18032_;
  assign new_n18051_ = pi0644 & new_n18037_;
  assign new_n18052_ = ~pi0715 & ~new_n18051_;
  assign new_n18053_ = ~new_n18050_ & new_n18052_;
  assign new_n18054_ = ~pi0644 & new_n18043_;
  assign new_n18055_ = pi0644 & new_n17832_;
  assign new_n18056_ = pi0715 & ~new_n18055_;
  assign new_n18057_ = ~new_n18054_ & new_n18056_;
  assign new_n18058_ = ~pi1160 & ~new_n18057_;
  assign new_n18059_ = ~new_n18053_ & new_n18058_;
  assign new_n18060_ = ~new_n18049_ & ~new_n18059_;
  assign new_n18061_ = pi0790 & ~new_n18060_;
  assign new_n18062_ = ~pi0790 & ~new_n18032_;
  assign new_n18063_ = pi0832 & ~new_n18062_;
  assign new_n18064_ = ~new_n18061_ & new_n18063_;
  assign po0297 = ~new_n17831_ & ~new_n18064_;
  assign new_n18066_ = pi0141 & ~new_n3272_;
  assign new_n18067_ = ~pi0141 & new_n16810_;
  assign new_n18068_ = pi0141 & new_n16928_;
  assign new_n18069_ = ~pi0749 & ~new_n18068_;
  assign new_n18070_ = ~new_n18067_ & new_n18069_;
  assign new_n18071_ = pi0141 & new_n17007_;
  assign new_n18072_ = ~pi0141 & ~new_n17074_;
  assign new_n18073_ = pi0749 & ~new_n18072_;
  assign new_n18074_ = ~new_n18071_ & new_n18073_;
  assign new_n18075_ = pi0039 & ~new_n18074_;
  assign new_n18076_ = ~new_n18070_ & new_n18075_;
  assign new_n18077_ = pi0141 & new_n17178_;
  assign new_n18078_ = ~pi0141 & new_n17217_;
  assign new_n18079_ = ~pi0749 & ~new_n18078_;
  assign new_n18080_ = ~new_n18077_ & new_n18079_;
  assign new_n18081_ = ~pi0141 & ~new_n17227_;
  assign new_n18082_ = pi0141 & ~new_n17234_;
  assign new_n18083_ = pi0749 & ~new_n18082_;
  assign new_n18084_ = ~new_n18081_ & new_n18083_;
  assign new_n18085_ = ~pi0039 & ~new_n18084_;
  assign new_n18086_ = ~new_n18080_ & new_n18085_;
  assign new_n18087_ = ~pi0038 & ~new_n18086_;
  assign new_n18088_ = ~new_n18076_ & new_n18087_;
  assign new_n18089_ = ~pi0141 & ~new_n17431_;
  assign new_n18090_ = pi0749 & new_n17433_;
  assign new_n18091_ = ~new_n18089_ & ~new_n18090_;
  assign new_n18092_ = ~pi0039 & new_n17247_;
  assign new_n18093_ = pi0038 & ~new_n18092_;
  assign new_n18094_ = new_n18091_ & new_n18093_;
  assign new_n18095_ = pi0706 & ~new_n18094_;
  assign new_n18096_ = ~new_n18088_ & new_n18095_;
  assign new_n18097_ = pi0038 & ~new_n18091_;
  assign new_n18098_ = ~pi0749 & new_n17347_;
  assign new_n18099_ = pi0141 & new_n17424_;
  assign new_n18100_ = ~new_n18098_ & ~new_n18099_;
  assign new_n18101_ = pi0039 & ~new_n18100_;
  assign new_n18102_ = ~pi0141 & new_n17393_;
  assign new_n18103_ = pi0141 & new_n17397_;
  assign new_n18104_ = pi0749 & ~new_n18103_;
  assign new_n18105_ = ~new_n18102_ & new_n18104_;
  assign new_n18106_ = ~pi0039 & new_n17260_;
  assign new_n18107_ = ~pi0141 & ~pi0749;
  assign new_n18108_ = ~new_n18106_ & new_n18107_;
  assign new_n18109_ = ~new_n18105_ & ~new_n18108_;
  assign new_n18110_ = ~pi0038 & ~new_n18109_;
  assign new_n18111_ = ~new_n18101_ & new_n18110_;
  assign new_n18112_ = ~new_n18097_ & ~new_n18111_;
  assign new_n18113_ = ~pi0706 & ~new_n18112_;
  assign new_n18114_ = new_n3272_ & ~new_n18113_;
  assign new_n18115_ = ~new_n18096_ & new_n18114_;
  assign new_n18116_ = ~new_n18066_ & ~new_n18115_;
  assign new_n18117_ = ~pi0625 & new_n18116_;
  assign new_n18118_ = new_n3272_ & new_n18112_;
  assign new_n18119_ = ~new_n18066_ & ~new_n18118_;
  assign new_n18120_ = pi0625 & new_n18119_;
  assign new_n18121_ = ~pi1153 & ~new_n18120_;
  assign new_n18122_ = ~new_n18117_ & new_n18121_;
  assign new_n18123_ = ~pi0039 & new_n17200_;
  assign new_n18124_ = ~new_n17534_ & ~new_n18123_;
  assign new_n18125_ = ~pi0141 & new_n18124_;
  assign new_n18126_ = pi0039 & ~new_n17483_;
  assign new_n18127_ = ~pi0039 & new_n17233_;
  assign new_n18128_ = ~new_n18126_ & ~new_n18127_;
  assign new_n18129_ = pi0141 & ~new_n18128_;
  assign new_n18130_ = ~pi0038 & ~new_n18129_;
  assign new_n18131_ = ~new_n18125_ & new_n18130_;
  assign new_n18132_ = new_n17544_ & ~new_n18089_;
  assign new_n18133_ = pi0706 & ~new_n18132_;
  assign new_n18134_ = ~new_n18131_ & new_n18133_;
  assign new_n18135_ = ~pi0141 & ~pi0706;
  assign new_n18136_ = ~new_n17551_ & new_n18135_;
  assign new_n18137_ = new_n3272_ & ~new_n18136_;
  assign new_n18138_ = ~new_n18134_ & new_n18137_;
  assign new_n18139_ = ~new_n18066_ & ~new_n18138_;
  assign new_n18140_ = pi0625 & new_n18139_;
  assign new_n18141_ = ~pi0141 & ~new_n17558_;
  assign new_n18142_ = ~pi0625 & new_n18141_;
  assign new_n18143_ = pi1153 & ~new_n18142_;
  assign new_n18144_ = ~new_n18140_ & new_n18143_;
  assign new_n18145_ = ~pi0608 & ~new_n18144_;
  assign new_n18146_ = ~new_n18122_ & new_n18145_;
  assign new_n18147_ = pi0625 & new_n18116_;
  assign new_n18148_ = ~pi0625 & new_n18119_;
  assign new_n18149_ = pi1153 & ~new_n18148_;
  assign new_n18150_ = ~new_n18147_ & new_n18149_;
  assign new_n18151_ = ~pi0625 & new_n18139_;
  assign new_n18152_ = pi0625 & new_n18141_;
  assign new_n18153_ = ~pi1153 & ~new_n18152_;
  assign new_n18154_ = ~new_n18151_ & new_n18153_;
  assign new_n18155_ = pi0608 & ~new_n18154_;
  assign new_n18156_ = ~new_n18150_ & new_n18155_;
  assign new_n18157_ = ~new_n18146_ & ~new_n18156_;
  assign new_n18158_ = pi0778 & ~new_n18157_;
  assign new_n18159_ = ~pi0778 & new_n18116_;
  assign new_n18160_ = ~new_n18158_ & ~new_n18159_;
  assign new_n18161_ = ~pi0609 & ~new_n18160_;
  assign new_n18162_ = ~pi0778 & ~new_n18139_;
  assign new_n18163_ = ~new_n18144_ & ~new_n18154_;
  assign new_n18164_ = pi0778 & ~new_n18163_;
  assign new_n18165_ = ~new_n18162_ & ~new_n18164_;
  assign new_n18166_ = pi0609 & new_n18165_;
  assign new_n18167_ = ~pi1155 & ~new_n18166_;
  assign new_n18168_ = ~new_n18161_ & new_n18167_;
  assign new_n18169_ = ~new_n17591_ & ~new_n18141_;
  assign new_n18170_ = ~new_n17590_ & ~new_n18119_;
  assign new_n18171_ = pi0609 & new_n18170_;
  assign new_n18172_ = ~new_n18169_ & ~new_n18171_;
  assign new_n18173_ = pi1155 & ~new_n18172_;
  assign new_n18174_ = ~pi0660 & ~new_n18173_;
  assign new_n18175_ = ~new_n18168_ & new_n18174_;
  assign new_n18176_ = pi0609 & ~new_n18160_;
  assign new_n18177_ = ~pi0609 & new_n18165_;
  assign new_n18178_ = pi1155 & ~new_n18177_;
  assign new_n18179_ = ~new_n18176_ & new_n18178_;
  assign new_n18180_ = ~new_n17603_ & ~new_n18141_;
  assign new_n18181_ = ~pi0609 & new_n18170_;
  assign new_n18182_ = ~new_n18180_ & ~new_n18181_;
  assign new_n18183_ = ~pi1155 & ~new_n18182_;
  assign new_n18184_ = pi0660 & ~new_n18183_;
  assign new_n18185_ = ~new_n18179_ & new_n18184_;
  assign new_n18186_ = ~new_n18175_ & ~new_n18185_;
  assign new_n18187_ = pi0785 & ~new_n18186_;
  assign new_n18188_ = ~pi0785 & ~new_n18160_;
  assign new_n18189_ = ~new_n18187_ & ~new_n18188_;
  assign new_n18190_ = ~pi0618 & ~new_n18189_;
  assign new_n18191_ = ~new_n17618_ & ~new_n18165_;
  assign new_n18192_ = new_n17618_ & ~new_n18141_;
  assign new_n18193_ = ~new_n18191_ & ~new_n18192_;
  assign new_n18194_ = pi0618 & new_n18193_;
  assign new_n18195_ = ~pi1154 & ~new_n18194_;
  assign new_n18196_ = ~new_n18190_ & new_n18195_;
  assign new_n18197_ = new_n17590_ & ~new_n18141_;
  assign new_n18198_ = ~new_n18170_ & ~new_n18197_;
  assign new_n18199_ = ~pi0785 & ~new_n18198_;
  assign new_n18200_ = ~new_n18173_ & ~new_n18183_;
  assign new_n18201_ = pi0785 & ~new_n18200_;
  assign new_n18202_ = ~new_n18199_ & ~new_n18201_;
  assign new_n18203_ = pi0618 & new_n18202_;
  assign new_n18204_ = ~pi0618 & new_n18141_;
  assign new_n18205_ = pi1154 & ~new_n18204_;
  assign new_n18206_ = ~new_n18203_ & new_n18205_;
  assign new_n18207_ = ~pi0627 & ~new_n18206_;
  assign new_n18208_ = ~new_n18196_ & new_n18207_;
  assign new_n18209_ = pi0618 & ~new_n18189_;
  assign new_n18210_ = ~pi0618 & new_n18193_;
  assign new_n18211_ = pi1154 & ~new_n18210_;
  assign new_n18212_ = ~new_n18209_ & new_n18211_;
  assign new_n18213_ = ~pi0618 & new_n18202_;
  assign new_n18214_ = pi0618 & new_n18141_;
  assign new_n18215_ = ~pi1154 & ~new_n18214_;
  assign new_n18216_ = ~new_n18213_ & new_n18215_;
  assign new_n18217_ = pi0627 & ~new_n18216_;
  assign new_n18218_ = ~new_n18212_ & new_n18217_;
  assign new_n18219_ = ~new_n18208_ & ~new_n18218_;
  assign new_n18220_ = pi0781 & ~new_n18219_;
  assign new_n18221_ = ~pi0781 & ~new_n18189_;
  assign new_n18222_ = ~new_n18220_ & ~new_n18221_;
  assign new_n18223_ = ~pi0619 & ~new_n18222_;
  assign new_n18224_ = ~new_n17655_ & new_n18193_;
  assign new_n18225_ = new_n17655_ & new_n18141_;
  assign new_n18226_ = ~new_n18224_ & ~new_n18225_;
  assign new_n18227_ = pi0619 & ~new_n18226_;
  assign new_n18228_ = ~pi1159 & ~new_n18227_;
  assign new_n18229_ = ~new_n18223_ & new_n18228_;
  assign new_n18230_ = ~pi0781 & ~new_n18202_;
  assign new_n18231_ = ~new_n18206_ & ~new_n18216_;
  assign new_n18232_ = pi0781 & ~new_n18231_;
  assign new_n18233_ = ~new_n18230_ & ~new_n18232_;
  assign new_n18234_ = pi0619 & new_n18233_;
  assign new_n18235_ = ~pi0619 & new_n18141_;
  assign new_n18236_ = pi1159 & ~new_n18235_;
  assign new_n18237_ = ~new_n18234_ & new_n18236_;
  assign new_n18238_ = ~pi0648 & ~new_n18237_;
  assign new_n18239_ = ~new_n18229_ & new_n18238_;
  assign new_n18240_ = pi0619 & ~new_n18222_;
  assign new_n18241_ = ~pi0619 & ~new_n18226_;
  assign new_n18242_ = pi1159 & ~new_n18241_;
  assign new_n18243_ = ~new_n18240_ & new_n18242_;
  assign new_n18244_ = ~pi0619 & new_n18233_;
  assign new_n18245_ = pi0619 & new_n18141_;
  assign new_n18246_ = ~pi1159 & ~new_n18245_;
  assign new_n18247_ = ~new_n18244_ & new_n18246_;
  assign new_n18248_ = pi0648 & ~new_n18247_;
  assign new_n18249_ = ~new_n18243_ & new_n18248_;
  assign new_n18250_ = ~new_n18239_ & ~new_n18249_;
  assign new_n18251_ = pi0789 & ~new_n18250_;
  assign new_n18252_ = ~pi0789 & ~new_n18222_;
  assign new_n18253_ = ~new_n18251_ & ~new_n18252_;
  assign new_n18254_ = ~pi0788 & new_n18253_;
  assign new_n18255_ = ~pi0626 & new_n18253_;
  assign new_n18256_ = new_n17691_ & ~new_n18141_;
  assign new_n18257_ = ~new_n17691_ & new_n18226_;
  assign new_n18258_ = ~new_n18256_ & ~new_n18257_;
  assign new_n18259_ = pi0626 & ~new_n18258_;
  assign new_n18260_ = ~pi0641 & ~new_n18259_;
  assign new_n18261_ = ~new_n18255_ & new_n18260_;
  assign new_n18262_ = ~pi0789 & ~new_n18233_;
  assign new_n18263_ = ~new_n18237_ & ~new_n18247_;
  assign new_n18264_ = pi0789 & ~new_n18263_;
  assign new_n18265_ = ~new_n18262_ & ~new_n18264_;
  assign new_n18266_ = ~pi0626 & new_n18265_;
  assign new_n18267_ = pi0626 & new_n18141_;
  assign new_n18268_ = ~pi1158 & ~new_n18267_;
  assign new_n18269_ = ~new_n18266_ & new_n18268_;
  assign new_n18270_ = ~new_n17698_ & ~new_n18269_;
  assign new_n18271_ = ~new_n18261_ & ~new_n18270_;
  assign new_n18272_ = pi0626 & new_n18253_;
  assign new_n18273_ = ~pi0626 & ~new_n18258_;
  assign new_n18274_ = pi0641 & ~new_n18273_;
  assign new_n18275_ = ~new_n18272_ & new_n18274_;
  assign new_n18276_ = pi0626 & new_n18265_;
  assign new_n18277_ = ~pi0626 & new_n18141_;
  assign new_n18278_ = pi1158 & ~new_n18277_;
  assign new_n18279_ = ~new_n18276_ & new_n18278_;
  assign new_n18280_ = ~new_n17713_ & ~new_n18279_;
  assign new_n18281_ = ~new_n18275_ & ~new_n18280_;
  assign new_n18282_ = ~new_n18271_ & ~new_n18281_;
  assign new_n18283_ = pi0788 & ~new_n18282_;
  assign new_n18284_ = ~new_n18254_ & ~new_n18283_;
  assign new_n18285_ = ~pi0628 & new_n18284_;
  assign new_n18286_ = ~new_n18269_ & ~new_n18279_;
  assign new_n18287_ = pi0788 & ~new_n18286_;
  assign new_n18288_ = ~pi0788 & ~new_n18265_;
  assign new_n18289_ = ~new_n18287_ & ~new_n18288_;
  assign new_n18290_ = pi0628 & new_n18289_;
  assign new_n18291_ = ~pi1156 & ~new_n18290_;
  assign new_n18292_ = ~new_n18285_ & new_n18291_;
  assign new_n18293_ = ~new_n17734_ & new_n18258_;
  assign new_n18294_ = new_n17734_ & new_n18141_;
  assign new_n18295_ = ~new_n18293_ & ~new_n18294_;
  assign new_n18296_ = pi0628 & ~new_n18295_;
  assign new_n18297_ = ~pi0628 & new_n18141_;
  assign new_n18298_ = pi1156 & ~new_n18297_;
  assign new_n18299_ = ~new_n18296_ & new_n18298_;
  assign new_n18300_ = ~pi0629 & ~new_n18299_;
  assign new_n18301_ = ~new_n18292_ & new_n18300_;
  assign new_n18302_ = pi0628 & new_n18284_;
  assign new_n18303_ = ~pi0628 & new_n18289_;
  assign new_n18304_ = pi1156 & ~new_n18303_;
  assign new_n18305_ = ~new_n18302_ & new_n18304_;
  assign new_n18306_ = ~pi0628 & ~new_n18295_;
  assign new_n18307_ = pi0628 & new_n18141_;
  assign new_n18308_ = ~pi1156 & ~new_n18307_;
  assign new_n18309_ = ~new_n18306_ & new_n18308_;
  assign new_n18310_ = pi0629 & ~new_n18309_;
  assign new_n18311_ = ~new_n18305_ & new_n18310_;
  assign new_n18312_ = ~new_n18301_ & ~new_n18311_;
  assign new_n18313_ = pi0792 & ~new_n18312_;
  assign new_n18314_ = ~pi0792 & new_n18284_;
  assign new_n18315_ = ~new_n18313_ & ~new_n18314_;
  assign new_n18316_ = ~pi0647 & ~new_n18315_;
  assign new_n18317_ = ~new_n17762_ & new_n18289_;
  assign new_n18318_ = new_n17762_ & new_n18141_;
  assign new_n18319_ = ~new_n18317_ & ~new_n18318_;
  assign new_n18320_ = pi0647 & ~new_n18319_;
  assign new_n18321_ = ~pi1157 & ~new_n18320_;
  assign new_n18322_ = ~new_n18316_ & new_n18321_;
  assign new_n18323_ = ~pi0792 & new_n18295_;
  assign new_n18324_ = ~new_n18299_ & ~new_n18309_;
  assign new_n18325_ = pi0792 & ~new_n18324_;
  assign new_n18326_ = ~new_n18323_ & ~new_n18325_;
  assign new_n18327_ = pi0647 & new_n18326_;
  assign new_n18328_ = ~pi0647 & new_n18141_;
  assign new_n18329_ = pi1157 & ~new_n18328_;
  assign new_n18330_ = ~new_n18327_ & new_n18329_;
  assign new_n18331_ = ~pi0630 & ~new_n18330_;
  assign new_n18332_ = ~new_n18322_ & new_n18331_;
  assign new_n18333_ = pi0647 & ~new_n18315_;
  assign new_n18334_ = ~pi0647 & ~new_n18319_;
  assign new_n18335_ = pi1157 & ~new_n18334_;
  assign new_n18336_ = ~new_n18333_ & new_n18335_;
  assign new_n18337_ = ~pi0647 & new_n18326_;
  assign new_n18338_ = pi0647 & new_n18141_;
  assign new_n18339_ = ~pi1157 & ~new_n18338_;
  assign new_n18340_ = ~new_n18337_ & new_n18339_;
  assign new_n18341_ = pi0630 & ~new_n18340_;
  assign new_n18342_ = ~new_n18336_ & new_n18341_;
  assign new_n18343_ = ~new_n18332_ & ~new_n18342_;
  assign new_n18344_ = pi0787 & ~new_n18343_;
  assign new_n18345_ = ~pi0787 & ~new_n18315_;
  assign new_n18346_ = ~new_n18344_ & ~new_n18345_;
  assign new_n18347_ = ~pi0644 & ~new_n18346_;
  assign new_n18348_ = ~pi0787 & ~new_n18326_;
  assign new_n18349_ = ~new_n18330_ & ~new_n18340_;
  assign new_n18350_ = pi0787 & ~new_n18349_;
  assign new_n18351_ = ~new_n18348_ & ~new_n18350_;
  assign new_n18352_ = pi0644 & new_n18351_;
  assign new_n18353_ = ~pi0715 & ~new_n18352_;
  assign new_n18354_ = ~new_n18347_ & new_n18353_;
  assign new_n18355_ = new_n17804_ & ~new_n18141_;
  assign new_n18356_ = ~new_n17804_ & new_n18319_;
  assign new_n18357_ = ~new_n18355_ & ~new_n18356_;
  assign new_n18358_ = ~pi0644 & new_n18357_;
  assign new_n18359_ = pi0644 & new_n18141_;
  assign new_n18360_ = pi0715 & ~new_n18359_;
  assign new_n18361_ = ~new_n18358_ & new_n18360_;
  assign new_n18362_ = ~pi1160 & ~new_n18361_;
  assign new_n18363_ = ~new_n18354_ & new_n18362_;
  assign new_n18364_ = pi0644 & ~new_n18346_;
  assign new_n18365_ = ~pi0644 & new_n18351_;
  assign new_n18366_ = pi0715 & ~new_n18365_;
  assign new_n18367_ = ~new_n18364_ & new_n18366_;
  assign new_n18368_ = pi0644 & new_n18357_;
  assign new_n18369_ = ~pi0644 & new_n18141_;
  assign new_n18370_ = ~pi0715 & ~new_n18369_;
  assign new_n18371_ = ~new_n18368_ & new_n18370_;
  assign new_n18372_ = pi1160 & ~new_n18371_;
  assign new_n18373_ = ~new_n18367_ & new_n18372_;
  assign new_n18374_ = pi0790 & ~new_n18373_;
  assign new_n18375_ = ~new_n18363_ & new_n18374_;
  assign new_n18376_ = ~pi0790 & new_n18346_;
  assign new_n18377_ = ~po1038 & ~new_n18376_;
  assign new_n18378_ = ~new_n18375_ & new_n18377_;
  assign new_n18379_ = ~pi0141 & po1038;
  assign new_n18380_ = ~pi0832 & ~new_n18379_;
  assign new_n18381_ = ~new_n18378_ & new_n18380_;
  assign new_n18382_ = ~pi0141 & ~new_n2754_;
  assign new_n18383_ = pi0706 & new_n16915_;
  assign new_n18384_ = ~new_n18382_ & ~new_n18383_;
  assign new_n18385_ = ~pi0778 & new_n18384_;
  assign new_n18386_ = ~pi0625 & new_n18383_;
  assign new_n18387_ = ~new_n18384_ & ~new_n18386_;
  assign new_n18388_ = pi1153 & ~new_n18387_;
  assign new_n18389_ = ~pi1153 & ~new_n18382_;
  assign new_n18390_ = ~new_n18386_ & new_n18389_;
  assign new_n18391_ = ~new_n18388_ & ~new_n18390_;
  assign new_n18392_ = pi0778 & ~new_n18391_;
  assign new_n18393_ = ~new_n18385_ & ~new_n18392_;
  assign new_n18394_ = ~new_n17844_ & new_n18393_;
  assign new_n18395_ = ~new_n17846_ & new_n18394_;
  assign new_n18396_ = ~new_n17848_ & new_n18395_;
  assign new_n18397_ = new_n17856_ & new_n18396_;
  assign new_n18398_ = pi0749 & new_n16913_;
  assign new_n18399_ = ~new_n18382_ & ~new_n18398_;
  assign new_n18400_ = ~new_n17858_ & ~new_n18399_;
  assign new_n18401_ = ~pi0785 & ~new_n18400_;
  assign new_n18402_ = ~new_n17863_ & ~new_n18399_;
  assign new_n18403_ = pi1155 & ~new_n18402_;
  assign new_n18404_ = ~new_n17866_ & new_n18400_;
  assign new_n18405_ = ~pi1155 & ~new_n18404_;
  assign new_n18406_ = ~new_n18403_ & ~new_n18405_;
  assign new_n18407_ = pi0785 & ~new_n18406_;
  assign new_n18408_ = ~new_n18401_ & ~new_n18407_;
  assign new_n18409_ = ~pi0781 & ~new_n18408_;
  assign new_n18410_ = ~new_n17873_ & new_n18408_;
  assign new_n18411_ = pi1154 & ~new_n18410_;
  assign new_n18412_ = ~new_n17876_ & new_n18408_;
  assign new_n18413_ = ~pi1154 & ~new_n18412_;
  assign new_n18414_ = ~new_n18411_ & ~new_n18413_;
  assign new_n18415_ = pi0781 & ~new_n18414_;
  assign new_n18416_ = ~new_n18409_ & ~new_n18415_;
  assign new_n18417_ = ~pi0789 & ~new_n18416_;
  assign new_n18418_ = pi0619 & new_n18416_;
  assign new_n18419_ = ~pi0619 & new_n18382_;
  assign new_n18420_ = pi1159 & ~new_n18419_;
  assign new_n18421_ = ~new_n18418_ & new_n18420_;
  assign new_n18422_ = ~pi0619 & new_n18416_;
  assign new_n18423_ = pi0619 & new_n18382_;
  assign new_n18424_ = ~pi1159 & ~new_n18423_;
  assign new_n18425_ = ~new_n18422_ & new_n18424_;
  assign new_n18426_ = ~new_n18421_ & ~new_n18425_;
  assign new_n18427_ = pi0789 & ~new_n18426_;
  assign new_n18428_ = ~new_n18417_ & ~new_n18427_;
  assign new_n18429_ = pi0626 & new_n18428_;
  assign new_n18430_ = ~pi0626 & new_n18382_;
  assign new_n18431_ = pi1158 & ~new_n18430_;
  assign new_n18432_ = ~new_n18429_ & new_n18431_;
  assign new_n18433_ = ~pi0626 & new_n18428_;
  assign new_n18434_ = pi0626 & new_n18382_;
  assign new_n18435_ = ~pi1158 & ~new_n18434_;
  assign new_n18436_ = ~new_n18433_ & new_n18435_;
  assign new_n18437_ = ~new_n18432_ & ~new_n18436_;
  assign new_n18438_ = ~new_n17733_ & new_n18437_;
  assign new_n18439_ = ~new_n18397_ & ~new_n18438_;
  assign new_n18440_ = pi0788 & ~new_n18439_;
  assign new_n18441_ = ~new_n16639_ & ~new_n18384_;
  assign new_n18442_ = pi0625 & new_n18441_;
  assign new_n18443_ = new_n18399_ & ~new_n18441_;
  assign new_n18444_ = ~new_n18442_ & ~new_n18443_;
  assign new_n18445_ = new_n18389_ & ~new_n18444_;
  assign new_n18446_ = ~pi0608 & ~new_n18388_;
  assign new_n18447_ = ~new_n18445_ & new_n18446_;
  assign new_n18448_ = pi1153 & new_n18399_;
  assign new_n18449_ = ~new_n18442_ & new_n18448_;
  assign new_n18450_ = pi0608 & ~new_n18390_;
  assign new_n18451_ = ~new_n18449_ & new_n18450_;
  assign new_n18452_ = ~new_n18447_ & ~new_n18451_;
  assign new_n18453_ = pi0778 & ~new_n18452_;
  assign new_n18454_ = ~pi0778 & ~new_n18443_;
  assign new_n18455_ = ~new_n18453_ & ~new_n18454_;
  assign new_n18456_ = ~pi0609 & ~new_n18455_;
  assign new_n18457_ = pi0609 & new_n18393_;
  assign new_n18458_ = ~pi1155 & ~new_n18457_;
  assign new_n18459_ = ~new_n18456_ & new_n18458_;
  assign new_n18460_ = ~pi0660 & ~new_n18403_;
  assign new_n18461_ = ~new_n18459_ & new_n18460_;
  assign new_n18462_ = pi0609 & ~new_n18455_;
  assign new_n18463_ = ~pi0609 & new_n18393_;
  assign new_n18464_ = pi1155 & ~new_n18463_;
  assign new_n18465_ = ~new_n18462_ & new_n18464_;
  assign new_n18466_ = pi0660 & ~new_n18405_;
  assign new_n18467_ = ~new_n18465_ & new_n18466_;
  assign new_n18468_ = ~new_n18461_ & ~new_n18467_;
  assign new_n18469_ = pi0785 & ~new_n18468_;
  assign new_n18470_ = ~pi0785 & ~new_n18455_;
  assign new_n18471_ = ~new_n18469_ & ~new_n18470_;
  assign new_n18472_ = ~pi0618 & ~new_n18471_;
  assign new_n18473_ = pi0618 & new_n18394_;
  assign new_n18474_ = ~pi1154 & ~new_n18473_;
  assign new_n18475_ = ~new_n18472_ & new_n18474_;
  assign new_n18476_ = ~pi0627 & ~new_n18411_;
  assign new_n18477_ = ~new_n18475_ & new_n18476_;
  assign new_n18478_ = pi0618 & ~new_n18471_;
  assign new_n18479_ = ~pi0618 & new_n18394_;
  assign new_n18480_ = pi1154 & ~new_n18479_;
  assign new_n18481_ = ~new_n18478_ & new_n18480_;
  assign new_n18482_ = pi0627 & ~new_n18413_;
  assign new_n18483_ = ~new_n18481_ & new_n18482_;
  assign new_n18484_ = ~new_n18477_ & ~new_n18483_;
  assign new_n18485_ = pi0781 & ~new_n18484_;
  assign new_n18486_ = ~pi0781 & ~new_n18471_;
  assign new_n18487_ = ~new_n18485_ & ~new_n18486_;
  assign new_n18488_ = pi0619 & ~new_n18487_;
  assign new_n18489_ = ~pi0619 & new_n18395_;
  assign new_n18490_ = pi1159 & ~new_n18489_;
  assign new_n18491_ = ~new_n18488_ & new_n18490_;
  assign new_n18492_ = pi0648 & ~new_n18425_;
  assign new_n18493_ = ~new_n18491_ & new_n18492_;
  assign new_n18494_ = ~pi0619 & ~new_n18487_;
  assign new_n18495_ = pi0619 & new_n18395_;
  assign new_n18496_ = ~pi1159 & ~new_n18495_;
  assign new_n18497_ = ~new_n18494_ & new_n18496_;
  assign new_n18498_ = ~pi0648 & ~new_n18421_;
  assign new_n18499_ = ~new_n18497_ & new_n18498_;
  assign new_n18500_ = pi0789 & ~new_n18499_;
  assign new_n18501_ = ~new_n18493_ & new_n18500_;
  assign new_n18502_ = ~pi0789 & new_n18487_;
  assign new_n18503_ = new_n17969_ & ~new_n18502_;
  assign new_n18504_ = ~new_n18501_ & new_n18503_;
  assign new_n18505_ = ~new_n18440_ & ~new_n18504_;
  assign new_n18506_ = ~pi0628 & ~new_n18505_;
  assign new_n18507_ = ~pi0788 & ~new_n18428_;
  assign new_n18508_ = pi0788 & ~new_n18437_;
  assign new_n18509_ = ~new_n18507_ & ~new_n18508_;
  assign new_n18510_ = pi0628 & new_n18509_;
  assign new_n18511_ = ~pi1156 & ~new_n18510_;
  assign new_n18512_ = ~new_n18506_ & new_n18511_;
  assign new_n18513_ = ~new_n17980_ & new_n18396_;
  assign new_n18514_ = ~new_n17982_ & new_n18513_;
  assign new_n18515_ = pi1156 & ~new_n18514_;
  assign new_n18516_ = ~pi0629 & ~new_n18515_;
  assign new_n18517_ = ~new_n18512_ & new_n18516_;
  assign new_n18518_ = pi0628 & ~new_n18505_;
  assign new_n18519_ = ~pi0628 & new_n18509_;
  assign new_n18520_ = pi1156 & ~new_n18519_;
  assign new_n18521_ = ~new_n18518_ & new_n18520_;
  assign new_n18522_ = ~new_n17991_ & new_n18513_;
  assign new_n18523_ = ~pi1156 & ~new_n18522_;
  assign new_n18524_ = pi0629 & ~new_n18523_;
  assign new_n18525_ = ~new_n18521_ & new_n18524_;
  assign new_n18526_ = ~new_n18517_ & ~new_n18525_;
  assign new_n18527_ = pi0792 & ~new_n18526_;
  assign new_n18528_ = ~pi0792 & ~new_n18505_;
  assign new_n18529_ = ~new_n18527_ & ~new_n18528_;
  assign new_n18530_ = ~pi0647 & ~new_n18529_;
  assign new_n18531_ = ~new_n17762_ & new_n18509_;
  assign new_n18532_ = new_n17762_ & new_n18382_;
  assign new_n18533_ = ~new_n18531_ & ~new_n18532_;
  assign new_n18534_ = pi0647 & ~new_n18533_;
  assign new_n18535_ = ~pi1157 & ~new_n18534_;
  assign new_n18536_ = ~new_n18530_ & new_n18535_;
  assign new_n18537_ = ~new_n18011_ & new_n18513_;
  assign new_n18538_ = pi0647 & new_n18537_;
  assign new_n18539_ = ~pi0647 & new_n18382_;
  assign new_n18540_ = pi1157 & ~new_n18539_;
  assign new_n18541_ = ~new_n18538_ & new_n18540_;
  assign new_n18542_ = ~pi0630 & ~new_n18541_;
  assign new_n18543_ = ~new_n18536_ & new_n18542_;
  assign new_n18544_ = pi0647 & ~new_n18529_;
  assign new_n18545_ = ~pi0647 & ~new_n18533_;
  assign new_n18546_ = pi1157 & ~new_n18545_;
  assign new_n18547_ = ~new_n18544_ & new_n18546_;
  assign new_n18548_ = ~pi0647 & new_n18537_;
  assign new_n18549_ = pi0647 & new_n18382_;
  assign new_n18550_ = ~pi1157 & ~new_n18549_;
  assign new_n18551_ = ~new_n18548_ & new_n18550_;
  assign new_n18552_ = pi0630 & ~new_n18551_;
  assign new_n18553_ = ~new_n18547_ & new_n18552_;
  assign new_n18554_ = ~new_n18543_ & ~new_n18553_;
  assign new_n18555_ = pi0787 & ~new_n18554_;
  assign new_n18556_ = ~pi0787 & ~new_n18529_;
  assign new_n18557_ = ~new_n18555_ & ~new_n18556_;
  assign new_n18558_ = pi0644 & ~new_n18557_;
  assign new_n18559_ = ~pi0787 & ~new_n18537_;
  assign new_n18560_ = ~new_n18541_ & ~new_n18551_;
  assign new_n18561_ = pi0787 & ~new_n18560_;
  assign new_n18562_ = ~new_n18559_ & ~new_n18561_;
  assign new_n18563_ = ~pi0644 & new_n18562_;
  assign new_n18564_ = pi0715 & ~new_n18563_;
  assign new_n18565_ = ~new_n18558_ & new_n18564_;
  assign new_n18566_ = new_n17804_ & ~new_n18382_;
  assign new_n18567_ = ~new_n17804_ & new_n18533_;
  assign new_n18568_ = ~new_n18566_ & ~new_n18567_;
  assign new_n18569_ = pi0644 & new_n18568_;
  assign new_n18570_ = ~pi0644 & new_n18382_;
  assign new_n18571_ = ~pi0715 & ~new_n18570_;
  assign new_n18572_ = ~new_n18569_ & new_n18571_;
  assign new_n18573_ = pi1160 & ~new_n18572_;
  assign new_n18574_ = ~new_n18565_ & new_n18573_;
  assign new_n18575_ = ~pi0644 & ~new_n18557_;
  assign new_n18576_ = pi0644 & new_n18562_;
  assign new_n18577_ = ~pi0715 & ~new_n18576_;
  assign new_n18578_ = ~new_n18575_ & new_n18577_;
  assign new_n18579_ = ~pi0644 & new_n18568_;
  assign new_n18580_ = pi0644 & new_n18382_;
  assign new_n18581_ = pi0715 & ~new_n18580_;
  assign new_n18582_ = ~new_n18579_ & new_n18581_;
  assign new_n18583_ = ~pi1160 & ~new_n18582_;
  assign new_n18584_ = ~new_n18578_ & new_n18583_;
  assign new_n18585_ = ~new_n18574_ & ~new_n18584_;
  assign new_n18586_ = pi0790 & ~new_n18585_;
  assign new_n18587_ = ~pi0790 & ~new_n18557_;
  assign new_n18588_ = pi0832 & ~new_n18587_;
  assign new_n18589_ = ~new_n18586_ & new_n18588_;
  assign po0298 = ~new_n18381_ & ~new_n18589_;
  assign new_n18591_ = pi0142 & ~new_n3272_;
  assign new_n18592_ = pi0142 & ~new_n17224_;
  assign new_n18593_ = new_n17189_ & new_n18592_;
  assign new_n18594_ = ~pi0142 & ~new_n17208_;
  assign new_n18595_ = ~new_n17229_ & new_n18594_;
  assign new_n18596_ = ~new_n18593_ & ~new_n18595_;
  assign new_n18597_ = pi0743 & ~new_n18596_;
  assign new_n18598_ = ~pi0142 & new_n17164_;
  assign new_n18599_ = pi0142 & ~new_n17189_;
  assign new_n18600_ = ~new_n17208_ & new_n18599_;
  assign new_n18601_ = ~pi0743 & ~new_n18600_;
  assign new_n18602_ = ~new_n18598_ & new_n18601_;
  assign new_n18603_ = ~pi0299 & ~new_n18602_;
  assign new_n18604_ = ~new_n18597_ & new_n18603_;
  assign new_n18605_ = ~pi0142 & new_n17176_;
  assign new_n18606_ = pi0142 & ~new_n17198_;
  assign new_n18607_ = ~new_n17213_ & new_n18606_;
  assign new_n18608_ = ~pi0743 & ~new_n18607_;
  assign new_n18609_ = ~new_n18605_ & new_n18608_;
  assign new_n18610_ = ~pi0142 & ~new_n17213_;
  assign new_n18611_ = ~new_n17231_ & new_n18610_;
  assign new_n18612_ = pi0142 & new_n17221_;
  assign new_n18613_ = ~new_n17197_ & new_n18612_;
  assign new_n18614_ = ~new_n18611_ & ~new_n18613_;
  assign new_n18615_ = pi0743 & ~new_n18614_;
  assign new_n18616_ = pi0299 & ~new_n18615_;
  assign new_n18617_ = ~new_n18609_ & new_n18616_;
  assign new_n18618_ = ~new_n18604_ & ~new_n18617_;
  assign new_n18619_ = pi0735 & ~new_n18618_;
  assign new_n18620_ = pi0743 & ~new_n18594_;
  assign new_n18621_ = ~new_n18592_ & new_n18620_;
  assign new_n18622_ = pi0142 & ~pi0743;
  assign new_n18623_ = ~new_n17182_ & new_n18622_;
  assign new_n18624_ = ~pi0299 & ~new_n18623_;
  assign new_n18625_ = ~new_n18621_ & new_n18624_;
  assign new_n18626_ = pi0142 & ~new_n17193_;
  assign new_n18627_ = ~pi0743 & ~new_n18626_;
  assign new_n18628_ = ~new_n18610_ & ~new_n18627_;
  assign new_n18629_ = ~new_n18612_ & new_n18628_;
  assign new_n18630_ = pi0299 & ~new_n18629_;
  assign new_n18631_ = ~new_n18625_ & ~new_n18630_;
  assign new_n18632_ = ~pi0735 & new_n18631_;
  assign new_n18633_ = ~pi0039 & ~new_n18632_;
  assign new_n18634_ = ~new_n18619_ & new_n18633_;
  assign new_n18635_ = pi0142 & new_n17049_;
  assign new_n18636_ = ~pi0142 & new_n16988_;
  assign new_n18637_ = pi0743 & ~new_n18636_;
  assign new_n18638_ = ~new_n18635_ & new_n18637_;
  assign new_n18639_ = ~pi0142 & ~new_n16888_;
  assign new_n18640_ = pi0142 & new_n16716_;
  assign new_n18641_ = ~pi0743 & ~new_n18640_;
  assign new_n18642_ = ~new_n18639_ & new_n18641_;
  assign new_n18643_ = ~new_n18638_ & ~new_n18642_;
  assign new_n18644_ = pi0735 & ~new_n18643_;
  assign new_n18645_ = pi0142 & ~new_n17272_;
  assign new_n18646_ = ~pi0743 & ~new_n18645_;
  assign new_n18647_ = pi0142 & ~new_n17372_;
  assign new_n18648_ = pi0743 & new_n16984_;
  assign new_n18649_ = ~new_n18647_ & new_n18648_;
  assign new_n18650_ = ~new_n18646_ & ~new_n18649_;
  assign new_n18651_ = ~pi0735 & new_n18650_;
  assign new_n18652_ = ~new_n18644_ & ~new_n18651_;
  assign new_n18653_ = ~new_n6212_ & new_n18652_;
  assign new_n18654_ = pi0142 & ~new_n17055_;
  assign new_n18655_ = ~pi0142 & ~new_n16982_;
  assign new_n18656_ = pi0743 & ~new_n18655_;
  assign new_n18657_ = ~new_n18654_ & new_n18656_;
  assign new_n18658_ = pi0142 & new_n16698_;
  assign new_n18659_ = ~pi0142 & new_n16900_;
  assign new_n18660_ = ~pi0743 & ~new_n18659_;
  assign new_n18661_ = ~new_n18658_ & new_n18660_;
  assign new_n18662_ = ~new_n18657_ & ~new_n18661_;
  assign new_n18663_ = pi0735 & ~new_n18662_;
  assign new_n18664_ = pi0142 & ~new_n17292_;
  assign new_n18665_ = ~pi0743 & ~new_n18664_;
  assign new_n18666_ = pi0142 & new_n17367_;
  assign new_n18667_ = pi0743 & new_n16978_;
  assign new_n18668_ = ~new_n18666_ & new_n18667_;
  assign new_n18669_ = ~new_n18665_ & ~new_n18668_;
  assign new_n18670_ = ~pi0735 & new_n18669_;
  assign new_n18671_ = ~new_n18663_ & ~new_n18670_;
  assign new_n18672_ = new_n6212_ & new_n18671_;
  assign new_n18673_ = pi0215 & ~new_n18672_;
  assign new_n18674_ = ~new_n18653_ & new_n18673_;
  assign new_n18675_ = ~pi0142 & ~new_n16963_;
  assign new_n18676_ = pi0142 & new_n17030_;
  assign new_n18677_ = pi0743 & ~new_n18676_;
  assign new_n18678_ = ~new_n18675_ & new_n18677_;
  assign new_n18679_ = pi0142 & new_n16768_;
  assign new_n18680_ = ~pi0142 & new_n16861_;
  assign new_n18681_ = ~pi0743 & ~new_n18680_;
  assign new_n18682_ = ~new_n18679_ & new_n18681_;
  assign new_n18683_ = ~new_n18678_ & ~new_n18682_;
  assign new_n18684_ = pi0735 & ~new_n18683_;
  assign new_n18685_ = ~pi0142 & new_n17401_;
  assign new_n18686_ = pi0142 & new_n17355_;
  assign new_n18687_ = ~new_n18685_ & ~new_n18686_;
  assign new_n18688_ = pi0743 & ~new_n18687_;
  assign new_n18689_ = pi0142 & ~new_n17313_;
  assign new_n18690_ = ~pi0743 & ~new_n18689_;
  assign new_n18691_ = ~new_n18688_ & ~new_n18690_;
  assign new_n18692_ = ~pi0735 & new_n18691_;
  assign new_n18693_ = ~new_n18684_ & ~new_n18692_;
  assign new_n18694_ = new_n6212_ & ~new_n18693_;
  assign new_n18695_ = ~pi0142 & ~new_n16945_;
  assign new_n18696_ = pi0142 & new_n17017_;
  assign new_n18697_ = pi0743 & ~new_n18696_;
  assign new_n18698_ = ~new_n18695_ & new_n18697_;
  assign new_n18699_ = ~pi0142 & ~new_n16840_;
  assign new_n18700_ = pi0142 & new_n16786_;
  assign new_n18701_ = ~pi0743 & ~new_n18700_;
  assign new_n18702_ = ~new_n18699_ & new_n18701_;
  assign new_n18703_ = ~new_n18698_ & ~new_n18702_;
  assign new_n18704_ = pi0735 & ~new_n18703_;
  assign new_n18705_ = pi0142 & ~new_n17320_;
  assign new_n18706_ = ~pi0743 & ~new_n18705_;
  assign new_n18707_ = pi0142 & ~new_n17360_;
  assign new_n18708_ = pi0743 & ~new_n16942_;
  assign new_n18709_ = ~new_n18707_ & new_n18708_;
  assign new_n18710_ = ~new_n18706_ & ~new_n18709_;
  assign new_n18711_ = ~pi0735 & new_n18710_;
  assign new_n18712_ = ~new_n18704_ & ~new_n18711_;
  assign new_n18713_ = ~new_n6212_ & ~new_n18712_;
  assign new_n18714_ = ~new_n3467_ & ~new_n18713_;
  assign new_n18715_ = ~new_n18694_ & new_n18714_;
  assign new_n18716_ = pi0142 & ~new_n16636_;
  assign new_n18717_ = pi0743 & new_n16661_;
  assign new_n18718_ = ~new_n18716_ & ~new_n18717_;
  assign new_n18719_ = ~pi0735 & new_n18718_;
  assign new_n18720_ = pi0142 & ~new_n16647_;
  assign new_n18721_ = pi0743 & new_n16913_;
  assign new_n18722_ = new_n3100_ & new_n18721_;
  assign new_n18723_ = ~new_n18720_ & ~new_n18722_;
  assign new_n18724_ = ~new_n17247_ & new_n18723_;
  assign new_n18725_ = ~new_n16633_ & ~new_n18724_;
  assign new_n18726_ = pi0735 & ~new_n18725_;
  assign new_n18727_ = ~new_n18716_ & new_n18726_;
  assign new_n18728_ = ~new_n18719_ & ~new_n18727_;
  assign new_n18729_ = new_n3467_ & ~new_n18728_;
  assign new_n18730_ = ~pi0215 & ~new_n18729_;
  assign new_n18731_ = ~new_n18715_ & new_n18730_;
  assign new_n18732_ = ~new_n18674_ & ~new_n18731_;
  assign new_n18733_ = pi0299 & ~new_n18732_;
  assign new_n18734_ = ~new_n6238_ & new_n18652_;
  assign new_n18735_ = new_n6238_ & new_n18671_;
  assign new_n18736_ = pi0223 & ~new_n18735_;
  assign new_n18737_ = ~new_n18734_ & new_n18736_;
  assign new_n18738_ = new_n6238_ & ~new_n18693_;
  assign new_n18739_ = ~new_n6238_ & ~new_n18712_;
  assign new_n18740_ = ~new_n3057_ & ~new_n18739_;
  assign new_n18741_ = ~new_n18738_ & new_n18740_;
  assign new_n18742_ = new_n3057_ & ~new_n18728_;
  assign new_n18743_ = ~pi0223 & ~new_n18742_;
  assign new_n18744_ = ~new_n18741_ & new_n18743_;
  assign new_n18745_ = ~new_n18737_ & ~new_n18744_;
  assign new_n18746_ = ~pi0299 & ~new_n18745_;
  assign new_n18747_ = pi0039 & ~new_n18746_;
  assign new_n18748_ = ~new_n18733_ & new_n18747_;
  assign new_n18749_ = ~new_n18634_ & ~new_n18748_;
  assign new_n18750_ = ~pi0038 & ~new_n18749_;
  assign new_n18751_ = pi0039 & pi0142;
  assign new_n18752_ = pi0038 & ~new_n18751_;
  assign new_n18753_ = pi0735 & new_n17247_;
  assign new_n18754_ = new_n18723_ & ~new_n18753_;
  assign new_n18755_ = ~pi0039 & ~new_n18754_;
  assign new_n18756_ = new_n18752_ & ~new_n18755_;
  assign new_n18757_ = new_n3272_ & ~new_n18756_;
  assign new_n18758_ = ~new_n18750_ & new_n18757_;
  assign new_n18759_ = ~new_n18591_ & ~new_n18758_;
  assign new_n18760_ = pi0625 & new_n18759_;
  assign new_n18761_ = ~new_n6212_ & new_n18710_;
  assign new_n18762_ = new_n6212_ & new_n18691_;
  assign new_n18763_ = ~new_n18761_ & ~new_n18762_;
  assign new_n18764_ = ~new_n3467_ & ~new_n18763_;
  assign new_n18765_ = new_n3467_ & ~new_n18718_;
  assign new_n18766_ = ~pi0215 & ~new_n18765_;
  assign new_n18767_ = ~new_n18764_ & new_n18766_;
  assign new_n18768_ = ~new_n6212_ & new_n18650_;
  assign new_n18769_ = new_n6212_ & new_n18669_;
  assign new_n18770_ = pi0215 & ~new_n18769_;
  assign new_n18771_ = ~new_n18768_ & new_n18770_;
  assign new_n18772_ = ~new_n18767_ & ~new_n18771_;
  assign new_n18773_ = pi0299 & ~new_n18772_;
  assign new_n18774_ = new_n6238_ & new_n18691_;
  assign new_n18775_ = ~new_n6238_ & new_n18710_;
  assign new_n18776_ = ~new_n3057_ & ~new_n18775_;
  assign new_n18777_ = ~new_n18774_ & new_n18776_;
  assign new_n18778_ = new_n3057_ & new_n18718_;
  assign new_n18779_ = ~pi0223 & ~new_n18778_;
  assign new_n18780_ = ~new_n18777_ & new_n18779_;
  assign new_n18781_ = ~new_n6238_ & ~new_n18650_;
  assign new_n18782_ = new_n6238_ & ~new_n18669_;
  assign new_n18783_ = pi0223 & ~new_n18782_;
  assign new_n18784_ = ~new_n18781_ & new_n18783_;
  assign new_n18785_ = ~pi0299 & ~new_n18784_;
  assign new_n18786_ = ~new_n18780_ & new_n18785_;
  assign new_n18787_ = pi0039 & ~new_n18786_;
  assign new_n18788_ = ~new_n18773_ & new_n18787_;
  assign new_n18789_ = ~pi0039 & new_n18631_;
  assign new_n18790_ = ~pi0038 & ~new_n18789_;
  assign new_n18791_ = ~new_n18788_ & new_n18790_;
  assign new_n18792_ = ~pi0039 & ~new_n18723_;
  assign new_n18793_ = new_n18752_ & ~new_n18792_;
  assign new_n18794_ = new_n3272_ & ~new_n18793_;
  assign new_n18795_ = ~new_n18791_ & new_n18794_;
  assign new_n18796_ = ~new_n18591_ & ~new_n18795_;
  assign new_n18797_ = ~pi0625 & new_n18796_;
  assign new_n18798_ = pi1153 & ~new_n18797_;
  assign new_n18799_ = ~new_n18760_ & new_n18798_;
  assign new_n18800_ = ~pi0142 & ~new_n17458_;
  assign new_n18801_ = pi0142 & ~new_n17494_;
  assign new_n18802_ = ~new_n18800_ & ~new_n18801_;
  assign new_n18803_ = pi0735 & ~new_n18802_;
  assign new_n18804_ = ~pi0735 & ~new_n18689_;
  assign new_n18805_ = ~new_n18803_ & ~new_n18804_;
  assign new_n18806_ = new_n6238_ & new_n18805_;
  assign new_n18807_ = ~pi0142 & new_n17451_;
  assign new_n18808_ = pi0142 & new_n17500_;
  assign new_n18809_ = ~new_n18807_ & ~new_n18808_;
  assign new_n18810_ = pi0735 & ~new_n18809_;
  assign new_n18811_ = ~pi0735 & ~new_n18705_;
  assign new_n18812_ = ~new_n18810_ & ~new_n18811_;
  assign new_n18813_ = ~new_n6238_ & new_n18812_;
  assign new_n18814_ = ~new_n3057_ & ~new_n18813_;
  assign new_n18815_ = ~new_n18806_ & new_n18814_;
  assign new_n18816_ = pi0735 & new_n16915_;
  assign new_n18817_ = new_n16635_ & new_n18816_;
  assign new_n18818_ = ~new_n18716_ & ~new_n18817_;
  assign new_n18819_ = new_n3057_ & new_n18818_;
  assign new_n18820_ = ~pi0223 & ~new_n18819_;
  assign new_n18821_ = ~new_n18815_ & new_n18820_;
  assign new_n18822_ = ~pi0735 & ~new_n18645_;
  assign new_n18823_ = pi0142 & ~new_n17511_;
  assign new_n18824_ = ~pi0142 & new_n16986_;
  assign new_n18825_ = new_n16985_ & new_n18824_;
  assign new_n18826_ = pi0735 & ~new_n18825_;
  assign new_n18827_ = ~new_n18823_ & new_n18826_;
  assign new_n18828_ = ~new_n18822_ & ~new_n18827_;
  assign new_n18829_ = ~new_n6238_ & ~new_n18828_;
  assign new_n18830_ = ~pi0735 & ~new_n18664_;
  assign new_n18831_ = pi0142 & ~new_n17513_;
  assign new_n18832_ = pi0735 & ~new_n18824_;
  assign new_n18833_ = ~new_n18831_ & new_n18832_;
  assign new_n18834_ = ~new_n18830_ & ~new_n18833_;
  assign new_n18835_ = new_n6238_ & ~new_n18834_;
  assign new_n18836_ = pi0223 & ~new_n18835_;
  assign new_n18837_ = ~new_n18829_ & new_n18836_;
  assign new_n18838_ = ~pi0299 & ~new_n18837_;
  assign new_n18839_ = ~new_n18821_ & new_n18838_;
  assign new_n18840_ = new_n6212_ & new_n18805_;
  assign new_n18841_ = ~new_n6212_ & new_n18812_;
  assign new_n18842_ = ~new_n3467_ & ~new_n18841_;
  assign new_n18843_ = ~new_n18840_ & new_n18842_;
  assign new_n18844_ = new_n3467_ & new_n18818_;
  assign new_n18845_ = ~pi0215 & ~new_n18844_;
  assign new_n18846_ = ~new_n18843_ & new_n18845_;
  assign new_n18847_ = ~new_n6212_ & ~new_n18828_;
  assign new_n18848_ = new_n6212_ & ~new_n18834_;
  assign new_n18849_ = pi0215 & ~new_n18848_;
  assign new_n18850_ = ~new_n18847_ & new_n18849_;
  assign new_n18851_ = pi0299 & ~new_n18850_;
  assign new_n18852_ = ~new_n18846_ & new_n18851_;
  assign new_n18853_ = pi0039 & ~new_n18852_;
  assign new_n18854_ = ~new_n18839_ & new_n18853_;
  assign new_n18855_ = pi0142 & new_n17200_;
  assign new_n18856_ = ~pi0142 & ~new_n17233_;
  assign new_n18857_ = pi0735 & ~new_n18856_;
  assign new_n18858_ = ~new_n18855_ & new_n18857_;
  assign new_n18859_ = pi0142 & ~pi0735;
  assign new_n18860_ = ~new_n17260_ & new_n18859_;
  assign new_n18861_ = ~new_n18858_ & ~new_n18860_;
  assign new_n18862_ = ~pi0039 & ~new_n18861_;
  assign new_n18863_ = ~pi0038 & ~new_n18862_;
  assign new_n18864_ = ~new_n18854_ & new_n18863_;
  assign new_n18865_ = new_n3100_ & new_n18816_;
  assign new_n18866_ = ~new_n18720_ & ~new_n18865_;
  assign new_n18867_ = ~pi0039 & ~new_n18866_;
  assign new_n18868_ = new_n18752_ & ~new_n18867_;
  assign new_n18869_ = new_n3272_ & ~new_n18868_;
  assign new_n18870_ = ~new_n18864_ & new_n18869_;
  assign new_n18871_ = ~new_n18591_ & ~new_n18870_;
  assign new_n18872_ = ~pi0625 & new_n18871_;
  assign new_n18873_ = new_n3272_ & ~new_n17550_;
  assign new_n18874_ = pi0142 & ~new_n18873_;
  assign new_n18875_ = pi0039 & ~new_n17327_;
  assign new_n18876_ = pi0142 & ~new_n18106_;
  assign new_n18877_ = ~new_n18875_ & new_n18876_;
  assign new_n18878_ = ~new_n6212_ & ~new_n18645_;
  assign new_n18879_ = new_n6212_ & ~new_n18664_;
  assign new_n18880_ = pi0215 & ~new_n18879_;
  assign new_n18881_ = ~new_n18878_ & new_n18880_;
  assign new_n18882_ = ~new_n6212_ & ~new_n18705_;
  assign new_n18883_ = new_n6212_ & ~new_n18689_;
  assign new_n18884_ = ~new_n18882_ & ~new_n18883_;
  assign new_n18885_ = ~new_n3467_ & ~new_n18884_;
  assign new_n18886_ = new_n3467_ & ~new_n18716_;
  assign new_n18887_ = ~pi0215 & ~new_n18886_;
  assign new_n18888_ = ~new_n18885_ & new_n18887_;
  assign new_n18889_ = ~new_n18881_ & ~new_n18888_;
  assign new_n18890_ = pi0039 & pi0299;
  assign new_n18891_ = ~new_n18889_ & new_n18890_;
  assign new_n18892_ = ~new_n18877_ & ~new_n18891_;
  assign new_n18893_ = new_n14865_ & ~new_n18892_;
  assign new_n18894_ = ~new_n18874_ & ~new_n18893_;
  assign new_n18895_ = pi0625 & new_n18894_;
  assign new_n18896_ = ~pi1153 & ~new_n18895_;
  assign new_n18897_ = ~new_n18872_ & new_n18896_;
  assign new_n18898_ = pi0608 & ~new_n18897_;
  assign new_n18899_ = ~new_n18799_ & new_n18898_;
  assign new_n18900_ = ~pi0625 & new_n18759_;
  assign new_n18901_ = pi0625 & new_n18796_;
  assign new_n18902_ = ~pi1153 & ~new_n18901_;
  assign new_n18903_ = ~new_n18900_ & new_n18902_;
  assign new_n18904_ = pi0625 & new_n18871_;
  assign new_n18905_ = ~pi0625 & new_n18894_;
  assign new_n18906_ = pi1153 & ~new_n18905_;
  assign new_n18907_ = ~new_n18904_ & new_n18906_;
  assign new_n18908_ = ~pi0608 & ~new_n18907_;
  assign new_n18909_ = ~new_n18903_ & new_n18908_;
  assign new_n18910_ = ~new_n18899_ & ~new_n18909_;
  assign new_n18911_ = pi0778 & ~new_n18910_;
  assign new_n18912_ = ~pi0778 & new_n18759_;
  assign new_n18913_ = ~new_n18911_ & ~new_n18912_;
  assign new_n18914_ = ~pi0609 & ~new_n18913_;
  assign new_n18915_ = ~pi0778 & ~new_n18871_;
  assign new_n18916_ = ~new_n18897_ & ~new_n18907_;
  assign new_n18917_ = pi0778 & ~new_n18916_;
  assign new_n18918_ = ~new_n18915_ & ~new_n18917_;
  assign new_n18919_ = pi0609 & new_n18918_;
  assign new_n18920_ = ~pi1155 & ~new_n18919_;
  assign new_n18921_ = ~new_n18914_ & new_n18920_;
  assign new_n18922_ = ~new_n17591_ & ~new_n18894_;
  assign new_n18923_ = ~new_n17590_ & ~new_n18796_;
  assign new_n18924_ = pi0609 & new_n18923_;
  assign new_n18925_ = ~new_n18922_ & ~new_n18924_;
  assign new_n18926_ = pi1155 & ~new_n18925_;
  assign new_n18927_ = ~pi0660 & ~new_n18926_;
  assign new_n18928_ = ~new_n18921_ & new_n18927_;
  assign new_n18929_ = pi0609 & ~new_n18913_;
  assign new_n18930_ = ~pi0609 & new_n18918_;
  assign new_n18931_ = pi1155 & ~new_n18930_;
  assign new_n18932_ = ~new_n18929_ & new_n18931_;
  assign new_n18933_ = ~new_n17603_ & ~new_n18894_;
  assign new_n18934_ = ~pi0609 & new_n18923_;
  assign new_n18935_ = ~new_n18933_ & ~new_n18934_;
  assign new_n18936_ = ~pi1155 & ~new_n18935_;
  assign new_n18937_ = pi0660 & ~new_n18936_;
  assign new_n18938_ = ~new_n18932_ & new_n18937_;
  assign new_n18939_ = ~new_n18928_ & ~new_n18938_;
  assign new_n18940_ = pi0785 & ~new_n18939_;
  assign new_n18941_ = ~pi0785 & ~new_n18913_;
  assign new_n18942_ = ~new_n18940_ & ~new_n18941_;
  assign new_n18943_ = ~pi0618 & ~new_n18942_;
  assign new_n18944_ = ~new_n17618_ & new_n18918_;
  assign new_n18945_ = new_n17618_ & new_n18894_;
  assign new_n18946_ = ~new_n18944_ & ~new_n18945_;
  assign new_n18947_ = pi0618 & ~new_n18946_;
  assign new_n18948_ = ~pi1154 & ~new_n18947_;
  assign new_n18949_ = ~new_n18943_ & new_n18948_;
  assign new_n18950_ = new_n17590_ & ~new_n18894_;
  assign new_n18951_ = ~new_n18923_ & ~new_n18950_;
  assign new_n18952_ = ~pi0785 & ~new_n18951_;
  assign new_n18953_ = ~new_n18926_ & ~new_n18936_;
  assign new_n18954_ = pi0785 & ~new_n18953_;
  assign new_n18955_ = ~new_n18952_ & ~new_n18954_;
  assign new_n18956_ = pi0618 & new_n18955_;
  assign new_n18957_ = ~pi0618 & new_n18894_;
  assign new_n18958_ = pi1154 & ~new_n18957_;
  assign new_n18959_ = ~new_n18956_ & new_n18958_;
  assign new_n18960_ = ~pi0627 & ~new_n18959_;
  assign new_n18961_ = ~new_n18949_ & new_n18960_;
  assign new_n18962_ = pi0618 & ~new_n18942_;
  assign new_n18963_ = ~pi0618 & ~new_n18946_;
  assign new_n18964_ = pi1154 & ~new_n18963_;
  assign new_n18965_ = ~new_n18962_ & new_n18964_;
  assign new_n18966_ = ~pi0618 & new_n18955_;
  assign new_n18967_ = pi0618 & new_n18894_;
  assign new_n18968_ = ~pi1154 & ~new_n18967_;
  assign new_n18969_ = ~new_n18966_ & new_n18968_;
  assign new_n18970_ = pi0627 & ~new_n18969_;
  assign new_n18971_ = ~new_n18965_ & new_n18970_;
  assign new_n18972_ = ~new_n18961_ & ~new_n18971_;
  assign new_n18973_ = pi0781 & ~new_n18972_;
  assign new_n18974_ = ~pi0781 & ~new_n18942_;
  assign new_n18975_ = ~new_n18973_ & ~new_n18974_;
  assign new_n18976_ = ~pi0619 & ~new_n18975_;
  assign new_n18977_ = new_n17655_ & ~new_n18894_;
  assign new_n18978_ = ~new_n17655_ & new_n18946_;
  assign new_n18979_ = ~new_n18977_ & ~new_n18978_;
  assign new_n18980_ = pi0619 & new_n18979_;
  assign new_n18981_ = ~pi1159 & ~new_n18980_;
  assign new_n18982_ = ~new_n18976_ & new_n18981_;
  assign new_n18983_ = ~pi0781 & ~new_n18955_;
  assign new_n18984_ = ~new_n18959_ & ~new_n18969_;
  assign new_n18985_ = pi0781 & ~new_n18984_;
  assign new_n18986_ = ~new_n18983_ & ~new_n18985_;
  assign new_n18987_ = pi0619 & new_n18986_;
  assign new_n18988_ = ~pi0619 & new_n18894_;
  assign new_n18989_ = pi1159 & ~new_n18988_;
  assign new_n18990_ = ~new_n18987_ & new_n18989_;
  assign new_n18991_ = ~pi0648 & ~new_n18990_;
  assign new_n18992_ = ~new_n18982_ & new_n18991_;
  assign new_n18993_ = pi0619 & ~new_n18975_;
  assign new_n18994_ = ~pi0619 & new_n18979_;
  assign new_n18995_ = pi1159 & ~new_n18994_;
  assign new_n18996_ = ~new_n18993_ & new_n18995_;
  assign new_n18997_ = ~pi0619 & new_n18986_;
  assign new_n18998_ = pi0619 & new_n18894_;
  assign new_n18999_ = ~pi1159 & ~new_n18998_;
  assign new_n19000_ = ~new_n18997_ & new_n18999_;
  assign new_n19001_ = pi0648 & ~new_n19000_;
  assign new_n19002_ = ~new_n18996_ & new_n19001_;
  assign new_n19003_ = ~new_n18992_ & ~new_n19002_;
  assign new_n19004_ = pi0789 & ~new_n19003_;
  assign new_n19005_ = ~pi0789 & ~new_n18975_;
  assign new_n19006_ = ~new_n19004_ & ~new_n19005_;
  assign new_n19007_ = ~pi0788 & new_n19006_;
  assign new_n19008_ = ~pi0626 & new_n19006_;
  assign new_n19009_ = ~new_n17691_ & new_n18979_;
  assign new_n19010_ = new_n17691_ & new_n18894_;
  assign new_n19011_ = ~new_n19009_ & ~new_n19010_;
  assign new_n19012_ = pi0626 & new_n19011_;
  assign new_n19013_ = ~pi0641 & ~new_n19012_;
  assign new_n19014_ = ~new_n19008_ & new_n19013_;
  assign new_n19015_ = ~pi0789 & ~new_n18986_;
  assign new_n19016_ = ~new_n18990_ & ~new_n19000_;
  assign new_n19017_ = pi0789 & ~new_n19016_;
  assign new_n19018_ = ~new_n19015_ & ~new_n19017_;
  assign new_n19019_ = ~pi0626 & new_n19018_;
  assign new_n19020_ = pi0626 & new_n18894_;
  assign new_n19021_ = ~pi1158 & ~new_n19020_;
  assign new_n19022_ = ~new_n19019_ & new_n19021_;
  assign new_n19023_ = ~new_n17698_ & ~new_n19022_;
  assign new_n19024_ = ~new_n19014_ & ~new_n19023_;
  assign new_n19025_ = pi0626 & new_n19006_;
  assign new_n19026_ = ~pi0626 & new_n19011_;
  assign new_n19027_ = pi0641 & ~new_n19026_;
  assign new_n19028_ = ~new_n19025_ & new_n19027_;
  assign new_n19029_ = pi0626 & new_n19018_;
  assign new_n19030_ = ~pi0626 & new_n18894_;
  assign new_n19031_ = pi1158 & ~new_n19030_;
  assign new_n19032_ = ~new_n19029_ & new_n19031_;
  assign new_n19033_ = ~new_n17713_ & ~new_n19032_;
  assign new_n19034_ = ~new_n19028_ & ~new_n19033_;
  assign new_n19035_ = ~new_n19024_ & ~new_n19034_;
  assign new_n19036_ = pi0788 & ~new_n19035_;
  assign new_n19037_ = ~new_n19007_ & ~new_n19036_;
  assign new_n19038_ = ~pi0628 & new_n19037_;
  assign new_n19039_ = ~new_n19022_ & ~new_n19032_;
  assign new_n19040_ = pi0788 & ~new_n19039_;
  assign new_n19041_ = ~pi0788 & ~new_n19018_;
  assign new_n19042_ = ~new_n19040_ & ~new_n19041_;
  assign new_n19043_ = pi0628 & new_n19042_;
  assign new_n19044_ = ~pi1156 & ~new_n19043_;
  assign new_n19045_ = ~new_n19038_ & new_n19044_;
  assign new_n19046_ = ~new_n17734_ & ~new_n19011_;
  assign new_n19047_ = new_n17734_ & new_n18894_;
  assign new_n19048_ = ~new_n19046_ & ~new_n19047_;
  assign new_n19049_ = pi0628 & ~new_n19048_;
  assign new_n19050_ = ~pi0628 & new_n18894_;
  assign new_n19051_ = pi1156 & ~new_n19050_;
  assign new_n19052_ = ~new_n19049_ & new_n19051_;
  assign new_n19053_ = ~pi0629 & ~new_n19052_;
  assign new_n19054_ = ~new_n19045_ & new_n19053_;
  assign new_n19055_ = pi0628 & new_n19037_;
  assign new_n19056_ = ~pi0628 & new_n19042_;
  assign new_n19057_ = pi1156 & ~new_n19056_;
  assign new_n19058_ = ~new_n19055_ & new_n19057_;
  assign new_n19059_ = ~pi0628 & ~new_n19048_;
  assign new_n19060_ = pi0628 & new_n18894_;
  assign new_n19061_ = ~pi1156 & ~new_n19060_;
  assign new_n19062_ = ~new_n19059_ & new_n19061_;
  assign new_n19063_ = pi0629 & ~new_n19062_;
  assign new_n19064_ = ~new_n19058_ & new_n19063_;
  assign new_n19065_ = ~new_n19054_ & ~new_n19064_;
  assign new_n19066_ = pi0792 & ~new_n19065_;
  assign new_n19067_ = ~pi0792 & new_n19037_;
  assign new_n19068_ = ~new_n19066_ & ~new_n19067_;
  assign new_n19069_ = ~pi0647 & ~new_n19068_;
  assign new_n19070_ = ~new_n17762_ & new_n19042_;
  assign new_n19071_ = new_n17762_ & new_n18894_;
  assign new_n19072_ = ~new_n19070_ & ~new_n19071_;
  assign new_n19073_ = pi0647 & ~new_n19072_;
  assign new_n19074_ = ~pi1157 & ~new_n19073_;
  assign new_n19075_ = ~new_n19069_ & new_n19074_;
  assign new_n19076_ = ~pi0792 & new_n19048_;
  assign new_n19077_ = ~new_n19052_ & ~new_n19062_;
  assign new_n19078_ = pi0792 & ~new_n19077_;
  assign new_n19079_ = ~new_n19076_ & ~new_n19078_;
  assign new_n19080_ = pi0647 & new_n19079_;
  assign new_n19081_ = ~pi0647 & new_n18894_;
  assign new_n19082_ = pi1157 & ~new_n19081_;
  assign new_n19083_ = ~new_n19080_ & new_n19082_;
  assign new_n19084_ = ~pi0630 & ~new_n19083_;
  assign new_n19085_ = ~new_n19075_ & new_n19084_;
  assign new_n19086_ = pi0647 & ~new_n19068_;
  assign new_n19087_ = ~pi0647 & ~new_n19072_;
  assign new_n19088_ = pi1157 & ~new_n19087_;
  assign new_n19089_ = ~new_n19086_ & new_n19088_;
  assign new_n19090_ = ~pi0647 & new_n19079_;
  assign new_n19091_ = pi0647 & new_n18894_;
  assign new_n19092_ = ~pi1157 & ~new_n19091_;
  assign new_n19093_ = ~new_n19090_ & new_n19092_;
  assign new_n19094_ = pi0630 & ~new_n19093_;
  assign new_n19095_ = ~new_n19089_ & new_n19094_;
  assign new_n19096_ = ~new_n19085_ & ~new_n19095_;
  assign new_n19097_ = pi0787 & ~new_n19096_;
  assign new_n19098_ = ~pi0787 & ~new_n19068_;
  assign new_n19099_ = ~new_n19097_ & ~new_n19098_;
  assign new_n19100_ = ~pi0644 & ~new_n19099_;
  assign new_n19101_ = ~pi0787 & ~new_n19079_;
  assign new_n19102_ = ~new_n19083_ & ~new_n19093_;
  assign new_n19103_ = pi0787 & ~new_n19102_;
  assign new_n19104_ = ~new_n19101_ & ~new_n19103_;
  assign new_n19105_ = pi0644 & new_n19104_;
  assign new_n19106_ = ~pi0715 & ~new_n19105_;
  assign new_n19107_ = ~new_n19100_ & new_n19106_;
  assign new_n19108_ = new_n17804_ & ~new_n18894_;
  assign new_n19109_ = ~new_n17804_ & new_n19072_;
  assign new_n19110_ = ~new_n19108_ & ~new_n19109_;
  assign new_n19111_ = ~pi0644 & new_n19110_;
  assign new_n19112_ = pi0644 & new_n18894_;
  assign new_n19113_ = pi0715 & ~new_n19112_;
  assign new_n19114_ = ~new_n19111_ & new_n19113_;
  assign new_n19115_ = ~pi1160 & ~new_n19114_;
  assign new_n19116_ = ~new_n19107_ & new_n19115_;
  assign new_n19117_ = pi0644 & ~new_n19099_;
  assign new_n19118_ = ~pi0644 & new_n19104_;
  assign new_n19119_ = pi0715 & ~new_n19118_;
  assign new_n19120_ = ~new_n19117_ & new_n19119_;
  assign new_n19121_ = pi0644 & new_n19110_;
  assign new_n19122_ = ~pi0644 & new_n18894_;
  assign new_n19123_ = ~pi0715 & ~new_n19122_;
  assign new_n19124_ = ~new_n19121_ & new_n19123_;
  assign new_n19125_ = pi1160 & ~new_n19124_;
  assign new_n19126_ = ~new_n19120_ & new_n19125_;
  assign new_n19127_ = pi0790 & ~new_n19126_;
  assign new_n19128_ = ~new_n19116_ & new_n19127_;
  assign new_n19129_ = ~pi0790 & new_n19099_;
  assign new_n19130_ = new_n6305_ & ~new_n19129_;
  assign new_n19131_ = ~new_n19128_ & new_n19130_;
  assign new_n19132_ = ~pi0142 & ~new_n6305_;
  assign new_n19133_ = ~pi0057 & ~new_n19132_;
  assign new_n19134_ = ~new_n19131_ & new_n19133_;
  assign new_n19135_ = pi0057 & pi0142;
  assign new_n19136_ = ~pi0832 & ~new_n19135_;
  assign new_n19137_ = ~new_n19134_ & new_n19136_;
  assign new_n19138_ = ~new_n17590_ & new_n18721_;
  assign new_n19139_ = pi0609 & new_n19138_;
  assign new_n19140_ = pi0142 & ~new_n2754_;
  assign new_n19141_ = pi1155 & ~new_n19140_;
  assign new_n19142_ = ~new_n19139_ & new_n19141_;
  assign new_n19143_ = ~pi0609 & new_n19138_;
  assign new_n19144_ = ~pi1155 & ~new_n19140_;
  assign new_n19145_ = ~new_n19143_ & new_n19144_;
  assign new_n19146_ = ~new_n19142_ & ~new_n19145_;
  assign new_n19147_ = pi0785 & ~new_n19146_;
  assign new_n19148_ = ~pi0785 & ~new_n19140_;
  assign new_n19149_ = ~new_n19138_ & new_n19148_;
  assign new_n19150_ = ~new_n19147_ & ~new_n19149_;
  assign new_n19151_ = ~pi0781 & ~new_n19150_;
  assign new_n19152_ = pi0618 & new_n19150_;
  assign new_n19153_ = ~pi0618 & new_n19140_;
  assign new_n19154_ = pi1154 & ~new_n19153_;
  assign new_n19155_ = ~new_n19152_ & new_n19154_;
  assign new_n19156_ = ~pi0618 & new_n19150_;
  assign new_n19157_ = pi0618 & new_n19140_;
  assign new_n19158_ = ~pi1154 & ~new_n19157_;
  assign new_n19159_ = ~new_n19156_ & new_n19158_;
  assign new_n19160_ = ~new_n19155_ & ~new_n19159_;
  assign new_n19161_ = pi0781 & ~new_n19160_;
  assign new_n19162_ = ~new_n19151_ & ~new_n19161_;
  assign new_n19163_ = ~pi0789 & ~new_n19162_;
  assign new_n19164_ = pi0619 & new_n19162_;
  assign new_n19165_ = ~pi0619 & new_n19140_;
  assign new_n19166_ = pi1159 & ~new_n19165_;
  assign new_n19167_ = ~new_n19164_ & new_n19166_;
  assign new_n19168_ = ~pi0619 & new_n19162_;
  assign new_n19169_ = pi0619 & new_n19140_;
  assign new_n19170_ = ~pi1159 & ~new_n19169_;
  assign new_n19171_ = ~new_n19168_ & new_n19170_;
  assign new_n19172_ = ~new_n19167_ & ~new_n19171_;
  assign new_n19173_ = pi0789 & ~new_n19172_;
  assign new_n19174_ = ~new_n19163_ & ~new_n19173_;
  assign new_n19175_ = pi0626 & new_n19174_;
  assign new_n19176_ = ~pi0626 & new_n19140_;
  assign new_n19177_ = pi1158 & ~new_n19176_;
  assign new_n19178_ = ~new_n19175_ & new_n19177_;
  assign new_n19179_ = ~pi0626 & new_n19174_;
  assign new_n19180_ = pi0626 & new_n19140_;
  assign new_n19181_ = ~pi1158 & ~new_n19180_;
  assign new_n19182_ = ~new_n19179_ & new_n19181_;
  assign new_n19183_ = ~new_n19178_ & ~new_n19182_;
  assign new_n19184_ = ~new_n17733_ & new_n19183_;
  assign new_n19185_ = ~pi0625 & pi1153;
  assign new_n19186_ = pi0625 & ~pi1153;
  assign new_n19187_ = ~new_n19185_ & ~new_n19186_;
  assign new_n19188_ = pi0778 & ~new_n19187_;
  assign new_n19189_ = new_n18816_ & ~new_n19188_;
  assign new_n19190_ = ~new_n19140_ & ~new_n19189_;
  assign new_n19191_ = ~new_n17618_ & ~new_n19190_;
  assign new_n19192_ = ~new_n17655_ & new_n19191_;
  assign new_n19193_ = ~new_n19140_ & ~new_n19192_;
  assign new_n19194_ = new_n17691_ & ~new_n19140_;
  assign new_n19195_ = new_n17856_ & ~new_n19194_;
  assign new_n19196_ = ~new_n19193_ & new_n19195_;
  assign new_n19197_ = ~new_n19184_ & ~new_n19196_;
  assign new_n19198_ = pi0788 & ~new_n19197_;
  assign new_n19199_ = pi0735 & new_n16916_;
  assign new_n19200_ = pi0625 & new_n19199_;
  assign new_n19201_ = ~new_n18721_ & ~new_n19140_;
  assign new_n19202_ = ~new_n19199_ & new_n19201_;
  assign new_n19203_ = ~new_n19200_ & ~new_n19202_;
  assign new_n19204_ = ~pi1153 & ~new_n19203_;
  assign new_n19205_ = pi0625 & new_n18816_;
  assign new_n19206_ = pi1153 & ~new_n19140_;
  assign new_n19207_ = ~new_n19205_ & new_n19206_;
  assign new_n19208_ = ~pi0608 & ~new_n19207_;
  assign new_n19209_ = ~new_n19204_ & new_n19208_;
  assign new_n19210_ = ~new_n18721_ & ~new_n19200_;
  assign new_n19211_ = pi1153 & ~new_n19210_;
  assign new_n19212_ = ~pi0625 & ~pi1153;
  assign new_n19213_ = new_n18816_ & new_n19212_;
  assign new_n19214_ = ~new_n19140_ & ~new_n19213_;
  assign new_n19215_ = ~new_n19211_ & new_n19214_;
  assign new_n19216_ = pi0608 & ~new_n19215_;
  assign new_n19217_ = ~new_n19209_ & ~new_n19216_;
  assign new_n19218_ = pi0778 & ~new_n19217_;
  assign new_n19219_ = ~pi0778 & ~new_n19202_;
  assign new_n19220_ = ~new_n19218_ & ~new_n19219_;
  assign new_n19221_ = ~pi0609 & ~new_n19220_;
  assign new_n19222_ = pi0609 & ~new_n19190_;
  assign new_n19223_ = ~pi1155 & ~new_n19222_;
  assign new_n19224_ = ~new_n19221_ & new_n19223_;
  assign new_n19225_ = ~pi0660 & ~new_n19142_;
  assign new_n19226_ = ~new_n19224_ & new_n19225_;
  assign new_n19227_ = pi0609 & ~new_n19220_;
  assign new_n19228_ = ~pi0609 & ~new_n19190_;
  assign new_n19229_ = pi1155 & ~new_n19228_;
  assign new_n19230_ = ~new_n19227_ & new_n19229_;
  assign new_n19231_ = pi0660 & ~new_n19145_;
  assign new_n19232_ = ~new_n19230_ & new_n19231_;
  assign new_n19233_ = ~new_n19226_ & ~new_n19232_;
  assign new_n19234_ = pi0785 & ~new_n19233_;
  assign new_n19235_ = ~pi0785 & ~new_n19220_;
  assign new_n19236_ = ~new_n19234_ & ~new_n19235_;
  assign new_n19237_ = ~pi0618 & ~new_n19236_;
  assign new_n19238_ = ~new_n19140_ & ~new_n19191_;
  assign new_n19239_ = pi0618 & ~new_n19238_;
  assign new_n19240_ = ~pi1154 & ~new_n19239_;
  assign new_n19241_ = ~new_n19237_ & new_n19240_;
  assign new_n19242_ = ~pi0627 & ~new_n19155_;
  assign new_n19243_ = ~new_n19241_ & new_n19242_;
  assign new_n19244_ = pi0618 & ~new_n19236_;
  assign new_n19245_ = ~pi0618 & ~new_n19238_;
  assign new_n19246_ = pi1154 & ~new_n19245_;
  assign new_n19247_ = ~new_n19244_ & new_n19246_;
  assign new_n19248_ = pi0627 & ~new_n19159_;
  assign new_n19249_ = ~new_n19247_ & new_n19248_;
  assign new_n19250_ = ~new_n19243_ & ~new_n19249_;
  assign new_n19251_ = pi0781 & ~new_n19250_;
  assign new_n19252_ = ~pi0781 & ~new_n19236_;
  assign new_n19253_ = ~new_n19251_ & ~new_n19252_;
  assign new_n19254_ = pi0619 & ~new_n19253_;
  assign new_n19255_ = ~pi0619 & ~new_n19193_;
  assign new_n19256_ = pi1159 & ~new_n19255_;
  assign new_n19257_ = ~new_n19254_ & new_n19256_;
  assign new_n19258_ = pi0648 & ~new_n19171_;
  assign new_n19259_ = ~new_n19257_ & new_n19258_;
  assign new_n19260_ = ~pi0619 & ~new_n19253_;
  assign new_n19261_ = pi0619 & ~new_n19193_;
  assign new_n19262_ = ~pi1159 & ~new_n19261_;
  assign new_n19263_ = ~new_n19260_ & new_n19262_;
  assign new_n19264_ = ~pi0648 & ~new_n19167_;
  assign new_n19265_ = ~new_n19263_ & new_n19264_;
  assign new_n19266_ = pi0789 & ~new_n19265_;
  assign new_n19267_ = ~new_n19259_ & new_n19266_;
  assign new_n19268_ = ~pi0789 & new_n19253_;
  assign new_n19269_ = new_n17969_ & ~new_n19268_;
  assign new_n19270_ = ~new_n19267_ & new_n19269_;
  assign new_n19271_ = ~new_n19198_ & ~new_n19270_;
  assign new_n19272_ = ~pi0628 & new_n19271_;
  assign new_n19273_ = ~pi0788 & ~new_n19174_;
  assign new_n19274_ = pi0788 & ~new_n19183_;
  assign new_n19275_ = ~new_n19273_ & ~new_n19274_;
  assign new_n19276_ = pi0628 & ~new_n19275_;
  assign new_n19277_ = ~pi1156 & ~new_n19276_;
  assign new_n19278_ = ~new_n19272_ & new_n19277_;
  assign new_n19279_ = ~new_n17691_ & ~new_n17734_;
  assign new_n19280_ = ~new_n17618_ & ~new_n17655_;
  assign new_n19281_ = new_n19279_ & new_n19280_;
  assign new_n19282_ = ~new_n19190_ & new_n19281_;
  assign new_n19283_ = pi0628 & new_n19282_;
  assign new_n19284_ = ~new_n19140_ & ~new_n19283_;
  assign new_n19285_ = pi1156 & ~new_n19284_;
  assign new_n19286_ = ~pi0629 & ~new_n19285_;
  assign new_n19287_ = ~new_n19278_ & new_n19286_;
  assign new_n19288_ = pi0628 & new_n19271_;
  assign new_n19289_ = ~pi0628 & ~new_n19275_;
  assign new_n19290_ = pi1156 & ~new_n19289_;
  assign new_n19291_ = ~new_n19288_ & new_n19290_;
  assign new_n19292_ = ~pi0628 & new_n19282_;
  assign new_n19293_ = ~new_n19140_ & ~new_n19292_;
  assign new_n19294_ = ~pi1156 & ~new_n19293_;
  assign new_n19295_ = pi0629 & ~new_n19294_;
  assign new_n19296_ = ~new_n19291_ & new_n19295_;
  assign new_n19297_ = ~new_n19287_ & ~new_n19296_;
  assign new_n19298_ = pi0792 & ~new_n19297_;
  assign new_n19299_ = ~pi0792 & new_n19271_;
  assign new_n19300_ = ~new_n19298_ & ~new_n19299_;
  assign new_n19301_ = ~pi0647 & new_n19300_;
  assign new_n19302_ = ~new_n17762_ & new_n19275_;
  assign new_n19303_ = new_n17762_ & new_n19140_;
  assign new_n19304_ = ~new_n19302_ & ~new_n19303_;
  assign new_n19305_ = pi0647 & ~new_n19304_;
  assign new_n19306_ = ~pi1157 & ~new_n19305_;
  assign new_n19307_ = ~new_n19301_ & new_n19306_;
  assign new_n19308_ = ~pi0628 & ~pi1156;
  assign new_n19309_ = pi0628 & pi1156;
  assign new_n19310_ = pi0792 & ~new_n19309_;
  assign new_n19311_ = ~new_n19308_ & new_n19310_;
  assign new_n19312_ = new_n19282_ & ~new_n19311_;
  assign new_n19313_ = pi0647 & new_n19312_;
  assign new_n19314_ = pi1157 & ~new_n19140_;
  assign new_n19315_ = ~new_n19313_ & new_n19314_;
  assign new_n19316_ = ~pi0630 & ~new_n19315_;
  assign new_n19317_ = ~new_n19307_ & new_n19316_;
  assign new_n19318_ = pi0647 & new_n19300_;
  assign new_n19319_ = ~pi0647 & ~new_n19304_;
  assign new_n19320_ = pi1157 & ~new_n19319_;
  assign new_n19321_ = ~new_n19318_ & new_n19320_;
  assign new_n19322_ = ~pi0647 & new_n19312_;
  assign new_n19323_ = ~pi1157 & ~new_n19140_;
  assign new_n19324_ = ~new_n19322_ & new_n19323_;
  assign new_n19325_ = pi0630 & ~new_n19324_;
  assign new_n19326_ = ~new_n19321_ & new_n19325_;
  assign new_n19327_ = ~new_n19317_ & ~new_n19326_;
  assign new_n19328_ = pi0787 & ~new_n19327_;
  assign new_n19329_ = ~pi0787 & new_n19300_;
  assign new_n19330_ = ~new_n19328_ & ~new_n19329_;
  assign new_n19331_ = pi0644 & ~new_n19330_;
  assign new_n19332_ = ~pi0647 & pi1157;
  assign new_n19333_ = pi0647 & ~pi1157;
  assign new_n19334_ = ~new_n19332_ & ~new_n19333_;
  assign new_n19335_ = pi0787 & ~new_n19334_;
  assign new_n19336_ = new_n19312_ & ~new_n19335_;
  assign new_n19337_ = ~new_n19140_ & ~new_n19336_;
  assign new_n19338_ = ~pi0644 & ~new_n19337_;
  assign new_n19339_ = pi0715 & ~new_n19338_;
  assign new_n19340_ = ~new_n19331_ & new_n19339_;
  assign new_n19341_ = new_n17804_ & ~new_n19140_;
  assign new_n19342_ = ~new_n17804_ & new_n19304_;
  assign new_n19343_ = ~new_n19341_ & ~new_n19342_;
  assign new_n19344_ = pi0644 & new_n19343_;
  assign new_n19345_ = ~pi0644 & new_n19140_;
  assign new_n19346_ = ~pi0715 & ~new_n19345_;
  assign new_n19347_ = ~new_n19344_ & new_n19346_;
  assign new_n19348_ = pi1160 & ~new_n19347_;
  assign new_n19349_ = ~new_n19340_ & new_n19348_;
  assign new_n19350_ = ~pi0644 & ~new_n19330_;
  assign new_n19351_ = pi0644 & ~new_n19337_;
  assign new_n19352_ = ~pi0715 & ~new_n19351_;
  assign new_n19353_ = ~new_n19350_ & new_n19352_;
  assign new_n19354_ = ~pi0644 & new_n19343_;
  assign new_n19355_ = pi0644 & new_n19140_;
  assign new_n19356_ = pi0715 & ~new_n19355_;
  assign new_n19357_ = ~new_n19354_ & new_n19356_;
  assign new_n19358_ = ~pi1160 & ~new_n19357_;
  assign new_n19359_ = ~new_n19353_ & new_n19358_;
  assign new_n19360_ = ~new_n19349_ & ~new_n19359_;
  assign new_n19361_ = pi0790 & ~new_n19360_;
  assign new_n19362_ = ~pi0790 & ~new_n19330_;
  assign new_n19363_ = pi0832 & ~new_n19362_;
  assign new_n19364_ = ~new_n19361_ & new_n19363_;
  assign po0299 = ~new_n19137_ & ~new_n19364_;
  assign new_n19366_ = pi0143 & ~new_n3272_;
  assign new_n19367_ = ~pi0143 & ~new_n17551_;
  assign new_n19368_ = pi0774 & ~new_n19367_;
  assign new_n19369_ = new_n6132_ & new_n16913_;
  assign new_n19370_ = pi0038 & new_n19369_;
  assign new_n19371_ = ~pi0038 & new_n17426_;
  assign new_n19372_ = pi0143 & ~new_n19371_;
  assign new_n19373_ = ~pi0038 & ~new_n17393_;
  assign new_n19374_ = new_n6257_ & new_n16869_;
  assign new_n19375_ = pi0038 & ~new_n19374_;
  assign new_n19376_ = ~new_n19373_ & ~new_n19375_;
  assign new_n19377_ = ~pi0143 & ~pi0774;
  assign new_n19378_ = new_n19376_ & new_n19377_;
  assign new_n19379_ = ~new_n19372_ & ~new_n19378_;
  assign new_n19380_ = ~new_n19370_ & ~new_n19379_;
  assign new_n19381_ = ~new_n19368_ & ~new_n19380_;
  assign new_n19382_ = ~pi0687 & new_n19381_;
  assign new_n19383_ = ~new_n16790_ & new_n17431_;
  assign new_n19384_ = pi0038 & new_n19383_;
  assign new_n19385_ = pi0039 & ~new_n16810_;
  assign new_n19386_ = ~pi0039 & ~new_n17217_;
  assign new_n19387_ = ~new_n19385_ & ~new_n19386_;
  assign new_n19388_ = ~pi0038 & ~new_n19387_;
  assign new_n19389_ = ~new_n19384_ & ~new_n19388_;
  assign new_n19390_ = ~pi0143 & new_n19389_;
  assign new_n19391_ = ~pi0039 & ~new_n17178_;
  assign new_n19392_ = pi0039 & ~new_n16928_;
  assign new_n19393_ = ~new_n19391_ & ~new_n19392_;
  assign new_n19394_ = ~pi0038 & new_n19393_;
  assign new_n19395_ = pi0143 & new_n19394_;
  assign new_n19396_ = pi0038 & new_n18092_;
  assign new_n19397_ = pi0774 & ~new_n19396_;
  assign new_n19398_ = ~new_n19395_ & new_n19397_;
  assign new_n19399_ = ~new_n19390_ & new_n19398_;
  assign new_n19400_ = new_n6257_ & ~new_n16917_;
  assign new_n19401_ = pi0038 & ~new_n19400_;
  assign new_n19402_ = pi0039 & ~new_n17007_;
  assign new_n19403_ = ~new_n17233_ & new_n17397_;
  assign new_n19404_ = ~new_n19402_ & ~new_n19403_;
  assign new_n19405_ = ~pi0038 & ~new_n19404_;
  assign new_n19406_ = ~new_n19401_ & ~new_n19405_;
  assign new_n19407_ = pi0143 & new_n19406_;
  assign new_n19408_ = pi0039 & ~new_n17074_;
  assign new_n19409_ = ~pi0039 & ~new_n17227_;
  assign new_n19410_ = ~pi0038 & new_n19409_;
  assign new_n19411_ = ~pi0039 & new_n17035_;
  assign new_n19412_ = pi0038 & ~new_n19411_;
  assign new_n19413_ = ~new_n19410_ & ~new_n19412_;
  assign new_n19414_ = ~new_n19408_ & new_n19413_;
  assign new_n19415_ = ~pi0143 & ~new_n19414_;
  assign new_n19416_ = ~pi0774 & ~new_n19415_;
  assign new_n19417_ = ~new_n19407_ & new_n19416_;
  assign new_n19418_ = pi0687 & ~new_n19417_;
  assign new_n19419_ = ~new_n19399_ & new_n19418_;
  assign new_n19420_ = new_n3272_ & ~new_n19419_;
  assign new_n19421_ = ~new_n19382_ & new_n19420_;
  assign new_n19422_ = ~new_n19366_ & ~new_n19421_;
  assign new_n19423_ = ~pi0625 & new_n19422_;
  assign new_n19424_ = new_n3272_ & ~new_n19381_;
  assign new_n19425_ = ~new_n19366_ & ~new_n19424_;
  assign new_n19426_ = pi0625 & new_n19425_;
  assign new_n19427_ = ~pi1153 & ~new_n19426_;
  assign new_n19428_ = ~new_n19423_ & new_n19427_;
  assign new_n19429_ = ~pi0143 & new_n18124_;
  assign new_n19430_ = pi0143 & ~new_n18128_;
  assign new_n19431_ = ~pi0038 & ~new_n19430_;
  assign new_n19432_ = ~new_n19429_ & new_n19431_;
  assign new_n19433_ = ~pi0143 & ~new_n17431_;
  assign new_n19434_ = new_n17544_ & ~new_n19433_;
  assign new_n19435_ = pi0687 & ~new_n19434_;
  assign new_n19436_ = ~new_n19432_ & new_n19435_;
  assign new_n19437_ = ~pi0687 & new_n19367_;
  assign new_n19438_ = new_n3272_ & ~new_n19437_;
  assign new_n19439_ = ~new_n19436_ & new_n19438_;
  assign new_n19440_ = ~new_n19366_ & ~new_n19439_;
  assign new_n19441_ = pi0625 & new_n19440_;
  assign new_n19442_ = ~pi0143 & ~new_n17558_;
  assign new_n19443_ = ~pi0625 & new_n19442_;
  assign new_n19444_ = pi1153 & ~new_n19443_;
  assign new_n19445_ = ~new_n19441_ & new_n19444_;
  assign new_n19446_ = ~pi0608 & ~new_n19445_;
  assign new_n19447_ = ~new_n19428_ & new_n19446_;
  assign new_n19448_ = pi0625 & new_n19422_;
  assign new_n19449_ = ~pi0625 & new_n19425_;
  assign new_n19450_ = pi1153 & ~new_n19449_;
  assign new_n19451_ = ~new_n19448_ & new_n19450_;
  assign new_n19452_ = ~pi0625 & new_n19440_;
  assign new_n19453_ = pi0625 & new_n19442_;
  assign new_n19454_ = ~pi1153 & ~new_n19453_;
  assign new_n19455_ = ~new_n19452_ & new_n19454_;
  assign new_n19456_ = pi0608 & ~new_n19455_;
  assign new_n19457_ = ~new_n19451_ & new_n19456_;
  assign new_n19458_ = ~new_n19447_ & ~new_n19457_;
  assign new_n19459_ = pi0778 & ~new_n19458_;
  assign new_n19460_ = ~pi0778 & new_n19422_;
  assign new_n19461_ = ~new_n19459_ & ~new_n19460_;
  assign new_n19462_ = ~pi0609 & ~new_n19461_;
  assign new_n19463_ = ~pi0778 & ~new_n19440_;
  assign new_n19464_ = ~new_n19445_ & ~new_n19455_;
  assign new_n19465_ = pi0778 & ~new_n19464_;
  assign new_n19466_ = ~new_n19463_ & ~new_n19465_;
  assign new_n19467_ = pi0609 & new_n19466_;
  assign new_n19468_ = ~pi1155 & ~new_n19467_;
  assign new_n19469_ = ~new_n19462_ & new_n19468_;
  assign new_n19470_ = ~new_n17591_ & ~new_n19442_;
  assign new_n19471_ = ~new_n17590_ & ~new_n19425_;
  assign new_n19472_ = pi0609 & new_n19471_;
  assign new_n19473_ = ~new_n19470_ & ~new_n19472_;
  assign new_n19474_ = pi1155 & ~new_n19473_;
  assign new_n19475_ = ~pi0660 & ~new_n19474_;
  assign new_n19476_ = ~new_n19469_ & new_n19475_;
  assign new_n19477_ = pi0609 & ~new_n19461_;
  assign new_n19478_ = ~pi0609 & new_n19466_;
  assign new_n19479_ = pi1155 & ~new_n19478_;
  assign new_n19480_ = ~new_n19477_ & new_n19479_;
  assign new_n19481_ = ~new_n17603_ & ~new_n19442_;
  assign new_n19482_ = ~pi0609 & new_n19471_;
  assign new_n19483_ = ~new_n19481_ & ~new_n19482_;
  assign new_n19484_ = ~pi1155 & ~new_n19483_;
  assign new_n19485_ = pi0660 & ~new_n19484_;
  assign new_n19486_ = ~new_n19480_ & new_n19485_;
  assign new_n19487_ = ~new_n19476_ & ~new_n19486_;
  assign new_n19488_ = pi0785 & ~new_n19487_;
  assign new_n19489_ = ~pi0785 & ~new_n19461_;
  assign new_n19490_ = ~new_n19488_ & ~new_n19489_;
  assign new_n19491_ = ~pi0618 & ~new_n19490_;
  assign new_n19492_ = ~new_n17618_ & ~new_n19466_;
  assign new_n19493_ = new_n17618_ & ~new_n19442_;
  assign new_n19494_ = ~new_n19492_ & ~new_n19493_;
  assign new_n19495_ = pi0618 & new_n19494_;
  assign new_n19496_ = ~pi1154 & ~new_n19495_;
  assign new_n19497_ = ~new_n19491_ & new_n19496_;
  assign new_n19498_ = new_n17590_ & ~new_n19442_;
  assign new_n19499_ = ~new_n19471_ & ~new_n19498_;
  assign new_n19500_ = ~pi0785 & ~new_n19499_;
  assign new_n19501_ = ~new_n19474_ & ~new_n19484_;
  assign new_n19502_ = pi0785 & ~new_n19501_;
  assign new_n19503_ = ~new_n19500_ & ~new_n19502_;
  assign new_n19504_ = pi0618 & new_n19503_;
  assign new_n19505_ = ~pi0618 & new_n19442_;
  assign new_n19506_ = pi1154 & ~new_n19505_;
  assign new_n19507_ = ~new_n19504_ & new_n19506_;
  assign new_n19508_ = ~pi0627 & ~new_n19507_;
  assign new_n19509_ = ~new_n19497_ & new_n19508_;
  assign new_n19510_ = pi0618 & ~new_n19490_;
  assign new_n19511_ = ~pi0618 & new_n19494_;
  assign new_n19512_ = pi1154 & ~new_n19511_;
  assign new_n19513_ = ~new_n19510_ & new_n19512_;
  assign new_n19514_ = ~pi0618 & new_n19503_;
  assign new_n19515_ = pi0618 & new_n19442_;
  assign new_n19516_ = ~pi1154 & ~new_n19515_;
  assign new_n19517_ = ~new_n19514_ & new_n19516_;
  assign new_n19518_ = pi0627 & ~new_n19517_;
  assign new_n19519_ = ~new_n19513_ & new_n19518_;
  assign new_n19520_ = ~new_n19509_ & ~new_n19519_;
  assign new_n19521_ = pi0781 & ~new_n19520_;
  assign new_n19522_ = ~pi0781 & ~new_n19490_;
  assign new_n19523_ = ~new_n19521_ & ~new_n19522_;
  assign new_n19524_ = ~pi0619 & ~new_n19523_;
  assign new_n19525_ = ~new_n17655_ & new_n19494_;
  assign new_n19526_ = new_n17655_ & new_n19442_;
  assign new_n19527_ = ~new_n19525_ & ~new_n19526_;
  assign new_n19528_ = pi0619 & ~new_n19527_;
  assign new_n19529_ = ~pi1159 & ~new_n19528_;
  assign new_n19530_ = ~new_n19524_ & new_n19529_;
  assign new_n19531_ = ~pi0781 & ~new_n19503_;
  assign new_n19532_ = ~new_n19507_ & ~new_n19517_;
  assign new_n19533_ = pi0781 & ~new_n19532_;
  assign new_n19534_ = ~new_n19531_ & ~new_n19533_;
  assign new_n19535_ = pi0619 & new_n19534_;
  assign new_n19536_ = ~pi0619 & new_n19442_;
  assign new_n19537_ = pi1159 & ~new_n19536_;
  assign new_n19538_ = ~new_n19535_ & new_n19537_;
  assign new_n19539_ = ~pi0648 & ~new_n19538_;
  assign new_n19540_ = ~new_n19530_ & new_n19539_;
  assign new_n19541_ = pi0619 & ~new_n19523_;
  assign new_n19542_ = ~pi0619 & ~new_n19527_;
  assign new_n19543_ = pi1159 & ~new_n19542_;
  assign new_n19544_ = ~new_n19541_ & new_n19543_;
  assign new_n19545_ = ~pi0619 & new_n19534_;
  assign new_n19546_ = pi0619 & new_n19442_;
  assign new_n19547_ = ~pi1159 & ~new_n19546_;
  assign new_n19548_ = ~new_n19545_ & new_n19547_;
  assign new_n19549_ = pi0648 & ~new_n19548_;
  assign new_n19550_ = ~new_n19544_ & new_n19549_;
  assign new_n19551_ = ~new_n19540_ & ~new_n19550_;
  assign new_n19552_ = pi0789 & ~new_n19551_;
  assign new_n19553_ = ~pi0789 & ~new_n19523_;
  assign new_n19554_ = ~new_n19552_ & ~new_n19553_;
  assign new_n19555_ = ~pi0788 & new_n19554_;
  assign new_n19556_ = ~pi0626 & new_n19554_;
  assign new_n19557_ = new_n17691_ & ~new_n19442_;
  assign new_n19558_ = ~new_n17691_ & new_n19527_;
  assign new_n19559_ = ~new_n19557_ & ~new_n19558_;
  assign new_n19560_ = pi0626 & ~new_n19559_;
  assign new_n19561_ = ~pi0641 & ~new_n19560_;
  assign new_n19562_ = ~new_n19556_ & new_n19561_;
  assign new_n19563_ = ~pi0789 & ~new_n19534_;
  assign new_n19564_ = ~new_n19538_ & ~new_n19548_;
  assign new_n19565_ = pi0789 & ~new_n19564_;
  assign new_n19566_ = ~new_n19563_ & ~new_n19565_;
  assign new_n19567_ = ~pi0626 & new_n19566_;
  assign new_n19568_ = pi0626 & new_n19442_;
  assign new_n19569_ = ~pi1158 & ~new_n19568_;
  assign new_n19570_ = ~new_n19567_ & new_n19569_;
  assign new_n19571_ = ~new_n17698_ & ~new_n19570_;
  assign new_n19572_ = ~new_n19562_ & ~new_n19571_;
  assign new_n19573_ = pi0626 & new_n19554_;
  assign new_n19574_ = ~pi0626 & ~new_n19559_;
  assign new_n19575_ = pi0641 & ~new_n19574_;
  assign new_n19576_ = ~new_n19573_ & new_n19575_;
  assign new_n19577_ = pi0626 & new_n19566_;
  assign new_n19578_ = ~pi0626 & new_n19442_;
  assign new_n19579_ = pi1158 & ~new_n19578_;
  assign new_n19580_ = ~new_n19577_ & new_n19579_;
  assign new_n19581_ = ~new_n17713_ & ~new_n19580_;
  assign new_n19582_ = ~new_n19576_ & ~new_n19581_;
  assign new_n19583_ = ~new_n19572_ & ~new_n19582_;
  assign new_n19584_ = pi0788 & ~new_n19583_;
  assign new_n19585_ = ~new_n19555_ & ~new_n19584_;
  assign new_n19586_ = ~pi0628 & new_n19585_;
  assign new_n19587_ = ~new_n19570_ & ~new_n19580_;
  assign new_n19588_ = pi0788 & ~new_n19587_;
  assign new_n19589_ = ~pi0788 & ~new_n19566_;
  assign new_n19590_ = ~new_n19588_ & ~new_n19589_;
  assign new_n19591_ = pi0628 & new_n19590_;
  assign new_n19592_ = ~pi1156 & ~new_n19591_;
  assign new_n19593_ = ~new_n19586_ & new_n19592_;
  assign new_n19594_ = ~new_n17734_ & new_n19559_;
  assign new_n19595_ = new_n17734_ & new_n19442_;
  assign new_n19596_ = ~new_n19594_ & ~new_n19595_;
  assign new_n19597_ = pi0628 & ~new_n19596_;
  assign new_n19598_ = ~pi0628 & new_n19442_;
  assign new_n19599_ = pi1156 & ~new_n19598_;
  assign new_n19600_ = ~new_n19597_ & new_n19599_;
  assign new_n19601_ = ~pi0629 & ~new_n19600_;
  assign new_n19602_ = ~new_n19593_ & new_n19601_;
  assign new_n19603_ = pi0628 & new_n19585_;
  assign new_n19604_ = ~pi0628 & new_n19590_;
  assign new_n19605_ = pi1156 & ~new_n19604_;
  assign new_n19606_ = ~new_n19603_ & new_n19605_;
  assign new_n19607_ = ~pi0628 & ~new_n19596_;
  assign new_n19608_ = pi0628 & new_n19442_;
  assign new_n19609_ = ~pi1156 & ~new_n19608_;
  assign new_n19610_ = ~new_n19607_ & new_n19609_;
  assign new_n19611_ = pi0629 & ~new_n19610_;
  assign new_n19612_ = ~new_n19606_ & new_n19611_;
  assign new_n19613_ = ~new_n19602_ & ~new_n19612_;
  assign new_n19614_ = pi0792 & ~new_n19613_;
  assign new_n19615_ = ~pi0792 & new_n19585_;
  assign new_n19616_ = ~new_n19614_ & ~new_n19615_;
  assign new_n19617_ = ~pi0647 & ~new_n19616_;
  assign new_n19618_ = ~new_n17762_ & new_n19590_;
  assign new_n19619_ = new_n17762_ & new_n19442_;
  assign new_n19620_ = ~new_n19618_ & ~new_n19619_;
  assign new_n19621_ = pi0647 & ~new_n19620_;
  assign new_n19622_ = ~pi1157 & ~new_n19621_;
  assign new_n19623_ = ~new_n19617_ & new_n19622_;
  assign new_n19624_ = ~pi0792 & new_n19596_;
  assign new_n19625_ = ~new_n19600_ & ~new_n19610_;
  assign new_n19626_ = pi0792 & ~new_n19625_;
  assign new_n19627_ = ~new_n19624_ & ~new_n19626_;
  assign new_n19628_ = pi0647 & new_n19627_;
  assign new_n19629_ = ~pi0647 & new_n19442_;
  assign new_n19630_ = pi1157 & ~new_n19629_;
  assign new_n19631_ = ~new_n19628_ & new_n19630_;
  assign new_n19632_ = ~pi0630 & ~new_n19631_;
  assign new_n19633_ = ~new_n19623_ & new_n19632_;
  assign new_n19634_ = pi0647 & ~new_n19616_;
  assign new_n19635_ = ~pi0647 & ~new_n19620_;
  assign new_n19636_ = pi1157 & ~new_n19635_;
  assign new_n19637_ = ~new_n19634_ & new_n19636_;
  assign new_n19638_ = ~pi0647 & new_n19627_;
  assign new_n19639_ = pi0647 & new_n19442_;
  assign new_n19640_ = ~pi1157 & ~new_n19639_;
  assign new_n19641_ = ~new_n19638_ & new_n19640_;
  assign new_n19642_ = pi0630 & ~new_n19641_;
  assign new_n19643_ = ~new_n19637_ & new_n19642_;
  assign new_n19644_ = ~new_n19633_ & ~new_n19643_;
  assign new_n19645_ = pi0787 & ~new_n19644_;
  assign new_n19646_ = ~pi0787 & ~new_n19616_;
  assign new_n19647_ = ~new_n19645_ & ~new_n19646_;
  assign new_n19648_ = ~pi0644 & ~new_n19647_;
  assign new_n19649_ = ~pi0787 & ~new_n19627_;
  assign new_n19650_ = ~new_n19631_ & ~new_n19641_;
  assign new_n19651_ = pi0787 & ~new_n19650_;
  assign new_n19652_ = ~new_n19649_ & ~new_n19651_;
  assign new_n19653_ = pi0644 & new_n19652_;
  assign new_n19654_ = ~pi0715 & ~new_n19653_;
  assign new_n19655_ = ~new_n19648_ & new_n19654_;
  assign new_n19656_ = new_n17804_ & ~new_n19442_;
  assign new_n19657_ = ~new_n17804_ & new_n19620_;
  assign new_n19658_ = ~new_n19656_ & ~new_n19657_;
  assign new_n19659_ = ~pi0644 & new_n19658_;
  assign new_n19660_ = pi0644 & new_n19442_;
  assign new_n19661_ = pi0715 & ~new_n19660_;
  assign new_n19662_ = ~new_n19659_ & new_n19661_;
  assign new_n19663_ = ~pi1160 & ~new_n19662_;
  assign new_n19664_ = ~new_n19655_ & new_n19663_;
  assign new_n19665_ = pi0644 & ~new_n19647_;
  assign new_n19666_ = ~pi0644 & new_n19652_;
  assign new_n19667_ = pi0715 & ~new_n19666_;
  assign new_n19668_ = ~new_n19665_ & new_n19667_;
  assign new_n19669_ = pi0644 & new_n19658_;
  assign new_n19670_ = ~pi0644 & new_n19442_;
  assign new_n19671_ = ~pi0715 & ~new_n19670_;
  assign new_n19672_ = ~new_n19669_ & new_n19671_;
  assign new_n19673_ = pi1160 & ~new_n19672_;
  assign new_n19674_ = ~new_n19668_ & new_n19673_;
  assign new_n19675_ = pi0790 & ~new_n19674_;
  assign new_n19676_ = ~new_n19664_ & new_n19675_;
  assign new_n19677_ = ~pi0790 & new_n19647_;
  assign new_n19678_ = ~po1038 & ~new_n19677_;
  assign new_n19679_ = ~new_n19676_ & new_n19678_;
  assign new_n19680_ = ~pi0143 & po1038;
  assign new_n19681_ = ~pi0832 & ~new_n19680_;
  assign new_n19682_ = ~new_n19679_ & new_n19681_;
  assign new_n19683_ = ~pi0143 & ~new_n2754_;
  assign new_n19684_ = pi0687 & new_n16915_;
  assign new_n19685_ = ~new_n19683_ & ~new_n19684_;
  assign new_n19686_ = ~pi0778 & new_n19685_;
  assign new_n19687_ = ~pi0625 & new_n19684_;
  assign new_n19688_ = ~new_n19685_ & ~new_n19687_;
  assign new_n19689_ = pi1153 & ~new_n19688_;
  assign new_n19690_ = ~pi1153 & ~new_n19683_;
  assign new_n19691_ = ~new_n19687_ & new_n19690_;
  assign new_n19692_ = ~new_n19689_ & ~new_n19691_;
  assign new_n19693_ = pi0778 & ~new_n19692_;
  assign new_n19694_ = ~new_n19686_ & ~new_n19693_;
  assign new_n19695_ = ~new_n17844_ & new_n19694_;
  assign new_n19696_ = ~new_n17846_ & new_n19695_;
  assign new_n19697_ = ~new_n17848_ & new_n19696_;
  assign new_n19698_ = new_n17856_ & new_n19697_;
  assign new_n19699_ = ~pi0774 & new_n16913_;
  assign new_n19700_ = ~new_n19683_ & ~new_n19699_;
  assign new_n19701_ = ~new_n17858_ & ~new_n19700_;
  assign new_n19702_ = ~pi0785 & ~new_n19701_;
  assign new_n19703_ = ~new_n17863_ & ~new_n19700_;
  assign new_n19704_ = pi1155 & ~new_n19703_;
  assign new_n19705_ = ~new_n17866_ & new_n19701_;
  assign new_n19706_ = ~pi1155 & ~new_n19705_;
  assign new_n19707_ = ~new_n19704_ & ~new_n19706_;
  assign new_n19708_ = pi0785 & ~new_n19707_;
  assign new_n19709_ = ~new_n19702_ & ~new_n19708_;
  assign new_n19710_ = ~pi0781 & ~new_n19709_;
  assign new_n19711_ = ~new_n17873_ & new_n19709_;
  assign new_n19712_ = pi1154 & ~new_n19711_;
  assign new_n19713_ = ~new_n17876_ & new_n19709_;
  assign new_n19714_ = ~pi1154 & ~new_n19713_;
  assign new_n19715_ = ~new_n19712_ & ~new_n19714_;
  assign new_n19716_ = pi0781 & ~new_n19715_;
  assign new_n19717_ = ~new_n19710_ & ~new_n19716_;
  assign new_n19718_ = ~pi0789 & ~new_n19717_;
  assign new_n19719_ = pi0619 & new_n19717_;
  assign new_n19720_ = ~pi0619 & new_n19683_;
  assign new_n19721_ = pi1159 & ~new_n19720_;
  assign new_n19722_ = ~new_n19719_ & new_n19721_;
  assign new_n19723_ = ~pi0619 & new_n19717_;
  assign new_n19724_ = pi0619 & new_n19683_;
  assign new_n19725_ = ~pi1159 & ~new_n19724_;
  assign new_n19726_ = ~new_n19723_ & new_n19725_;
  assign new_n19727_ = ~new_n19722_ & ~new_n19726_;
  assign new_n19728_ = pi0789 & ~new_n19727_;
  assign new_n19729_ = ~new_n19718_ & ~new_n19728_;
  assign new_n19730_ = pi0626 & new_n19729_;
  assign new_n19731_ = ~pi0626 & new_n19683_;
  assign new_n19732_ = pi1158 & ~new_n19731_;
  assign new_n19733_ = ~new_n19730_ & new_n19732_;
  assign new_n19734_ = ~pi0626 & new_n19729_;
  assign new_n19735_ = pi0626 & new_n19683_;
  assign new_n19736_ = ~pi1158 & ~new_n19735_;
  assign new_n19737_ = ~new_n19734_ & new_n19736_;
  assign new_n19738_ = ~new_n19733_ & ~new_n19737_;
  assign new_n19739_ = ~new_n17733_ & new_n19738_;
  assign new_n19740_ = ~new_n19698_ & ~new_n19739_;
  assign new_n19741_ = pi0788 & ~new_n19740_;
  assign new_n19742_ = ~new_n16639_ & ~new_n19685_;
  assign new_n19743_ = pi0625 & new_n19742_;
  assign new_n19744_ = new_n19700_ & ~new_n19742_;
  assign new_n19745_ = ~new_n19743_ & ~new_n19744_;
  assign new_n19746_ = new_n19690_ & ~new_n19745_;
  assign new_n19747_ = ~pi0608 & ~new_n19689_;
  assign new_n19748_ = ~new_n19746_ & new_n19747_;
  assign new_n19749_ = pi1153 & new_n19700_;
  assign new_n19750_ = ~new_n19743_ & new_n19749_;
  assign new_n19751_ = pi0608 & ~new_n19691_;
  assign new_n19752_ = ~new_n19750_ & new_n19751_;
  assign new_n19753_ = ~new_n19748_ & ~new_n19752_;
  assign new_n19754_ = pi0778 & ~new_n19753_;
  assign new_n19755_ = ~pi0778 & ~new_n19744_;
  assign new_n19756_ = ~new_n19754_ & ~new_n19755_;
  assign new_n19757_ = ~pi0609 & ~new_n19756_;
  assign new_n19758_ = pi0609 & new_n19694_;
  assign new_n19759_ = ~pi1155 & ~new_n19758_;
  assign new_n19760_ = ~new_n19757_ & new_n19759_;
  assign new_n19761_ = ~pi0660 & ~new_n19704_;
  assign new_n19762_ = ~new_n19760_ & new_n19761_;
  assign new_n19763_ = pi0609 & ~new_n19756_;
  assign new_n19764_ = ~pi0609 & new_n19694_;
  assign new_n19765_ = pi1155 & ~new_n19764_;
  assign new_n19766_ = ~new_n19763_ & new_n19765_;
  assign new_n19767_ = pi0660 & ~new_n19706_;
  assign new_n19768_ = ~new_n19766_ & new_n19767_;
  assign new_n19769_ = ~new_n19762_ & ~new_n19768_;
  assign new_n19770_ = pi0785 & ~new_n19769_;
  assign new_n19771_ = ~pi0785 & ~new_n19756_;
  assign new_n19772_ = ~new_n19770_ & ~new_n19771_;
  assign new_n19773_ = ~pi0618 & ~new_n19772_;
  assign new_n19774_ = pi0618 & new_n19695_;
  assign new_n19775_ = ~pi1154 & ~new_n19774_;
  assign new_n19776_ = ~new_n19773_ & new_n19775_;
  assign new_n19777_ = ~pi0627 & ~new_n19712_;
  assign new_n19778_ = ~new_n19776_ & new_n19777_;
  assign new_n19779_ = pi0618 & ~new_n19772_;
  assign new_n19780_ = ~pi0618 & new_n19695_;
  assign new_n19781_ = pi1154 & ~new_n19780_;
  assign new_n19782_ = ~new_n19779_ & new_n19781_;
  assign new_n19783_ = pi0627 & ~new_n19714_;
  assign new_n19784_ = ~new_n19782_ & new_n19783_;
  assign new_n19785_ = ~new_n19778_ & ~new_n19784_;
  assign new_n19786_ = pi0781 & ~new_n19785_;
  assign new_n19787_ = ~pi0781 & ~new_n19772_;
  assign new_n19788_ = ~new_n19786_ & ~new_n19787_;
  assign new_n19789_ = pi0619 & ~new_n19788_;
  assign new_n19790_ = ~pi0619 & new_n19696_;
  assign new_n19791_ = pi1159 & ~new_n19790_;
  assign new_n19792_ = ~new_n19789_ & new_n19791_;
  assign new_n19793_ = pi0648 & ~new_n19726_;
  assign new_n19794_ = ~new_n19792_ & new_n19793_;
  assign new_n19795_ = ~pi0619 & ~new_n19788_;
  assign new_n19796_ = pi0619 & new_n19696_;
  assign new_n19797_ = ~pi1159 & ~new_n19796_;
  assign new_n19798_ = ~new_n19795_ & new_n19797_;
  assign new_n19799_ = ~pi0648 & ~new_n19722_;
  assign new_n19800_ = ~new_n19798_ & new_n19799_;
  assign new_n19801_ = pi0789 & ~new_n19800_;
  assign new_n19802_ = ~new_n19794_ & new_n19801_;
  assign new_n19803_ = ~pi0789 & new_n19788_;
  assign new_n19804_ = new_n17969_ & ~new_n19803_;
  assign new_n19805_ = ~new_n19802_ & new_n19804_;
  assign new_n19806_ = ~new_n19741_ & ~new_n19805_;
  assign new_n19807_ = ~pi0628 & ~new_n19806_;
  assign new_n19808_ = ~pi0788 & ~new_n19729_;
  assign new_n19809_ = pi0788 & ~new_n19738_;
  assign new_n19810_ = ~new_n19808_ & ~new_n19809_;
  assign new_n19811_ = pi0628 & new_n19810_;
  assign new_n19812_ = ~pi1156 & ~new_n19811_;
  assign new_n19813_ = ~new_n19807_ & new_n19812_;
  assign new_n19814_ = ~new_n17980_ & new_n19697_;
  assign new_n19815_ = ~new_n17982_ & new_n19814_;
  assign new_n19816_ = pi1156 & ~new_n19815_;
  assign new_n19817_ = ~pi0629 & ~new_n19816_;
  assign new_n19818_ = ~new_n19813_ & new_n19817_;
  assign new_n19819_ = pi0628 & ~new_n19806_;
  assign new_n19820_ = ~pi0628 & new_n19810_;
  assign new_n19821_ = pi1156 & ~new_n19820_;
  assign new_n19822_ = ~new_n19819_ & new_n19821_;
  assign new_n19823_ = ~new_n17991_ & new_n19814_;
  assign new_n19824_ = ~pi1156 & ~new_n19823_;
  assign new_n19825_ = pi0629 & ~new_n19824_;
  assign new_n19826_ = ~new_n19822_ & new_n19825_;
  assign new_n19827_ = ~new_n19818_ & ~new_n19826_;
  assign new_n19828_ = pi0792 & ~new_n19827_;
  assign new_n19829_ = ~pi0792 & ~new_n19806_;
  assign new_n19830_ = ~new_n19828_ & ~new_n19829_;
  assign new_n19831_ = ~pi0647 & ~new_n19830_;
  assign new_n19832_ = ~new_n17762_ & new_n19810_;
  assign new_n19833_ = new_n17762_ & new_n19683_;
  assign new_n19834_ = ~new_n19832_ & ~new_n19833_;
  assign new_n19835_ = pi0647 & ~new_n19834_;
  assign new_n19836_ = ~pi1157 & ~new_n19835_;
  assign new_n19837_ = ~new_n19831_ & new_n19836_;
  assign new_n19838_ = ~new_n18011_ & new_n19814_;
  assign new_n19839_ = pi0647 & new_n19838_;
  assign new_n19840_ = ~pi0647 & new_n19683_;
  assign new_n19841_ = pi1157 & ~new_n19840_;
  assign new_n19842_ = ~new_n19839_ & new_n19841_;
  assign new_n19843_ = ~pi0630 & ~new_n19842_;
  assign new_n19844_ = ~new_n19837_ & new_n19843_;
  assign new_n19845_ = pi0647 & ~new_n19830_;
  assign new_n19846_ = ~pi0647 & ~new_n19834_;
  assign new_n19847_ = pi1157 & ~new_n19846_;
  assign new_n19848_ = ~new_n19845_ & new_n19847_;
  assign new_n19849_ = ~pi0647 & new_n19838_;
  assign new_n19850_ = pi0647 & new_n19683_;
  assign new_n19851_ = ~pi1157 & ~new_n19850_;
  assign new_n19852_ = ~new_n19849_ & new_n19851_;
  assign new_n19853_ = pi0630 & ~new_n19852_;
  assign new_n19854_ = ~new_n19848_ & new_n19853_;
  assign new_n19855_ = ~new_n19844_ & ~new_n19854_;
  assign new_n19856_ = pi0787 & ~new_n19855_;
  assign new_n19857_ = ~pi0787 & ~new_n19830_;
  assign new_n19858_ = ~new_n19856_ & ~new_n19857_;
  assign new_n19859_ = pi0644 & ~new_n19858_;
  assign new_n19860_ = ~pi0787 & ~new_n19838_;
  assign new_n19861_ = ~new_n19842_ & ~new_n19852_;
  assign new_n19862_ = pi0787 & ~new_n19861_;
  assign new_n19863_ = ~new_n19860_ & ~new_n19862_;
  assign new_n19864_ = ~pi0644 & new_n19863_;
  assign new_n19865_ = pi0715 & ~new_n19864_;
  assign new_n19866_ = ~new_n19859_ & new_n19865_;
  assign new_n19867_ = new_n17804_ & ~new_n19683_;
  assign new_n19868_ = ~new_n17804_ & new_n19834_;
  assign new_n19869_ = ~new_n19867_ & ~new_n19868_;
  assign new_n19870_ = pi0644 & new_n19869_;
  assign new_n19871_ = ~pi0644 & new_n19683_;
  assign new_n19872_ = ~pi0715 & ~new_n19871_;
  assign new_n19873_ = ~new_n19870_ & new_n19872_;
  assign new_n19874_ = pi1160 & ~new_n19873_;
  assign new_n19875_ = ~new_n19866_ & new_n19874_;
  assign new_n19876_ = ~pi0644 & ~new_n19858_;
  assign new_n19877_ = pi0644 & new_n19863_;
  assign new_n19878_ = ~pi0715 & ~new_n19877_;
  assign new_n19879_ = ~new_n19876_ & new_n19878_;
  assign new_n19880_ = ~pi0644 & new_n19869_;
  assign new_n19881_ = pi0644 & new_n19683_;
  assign new_n19882_ = pi0715 & ~new_n19881_;
  assign new_n19883_ = ~new_n19880_ & new_n19882_;
  assign new_n19884_ = ~pi1160 & ~new_n19883_;
  assign new_n19885_ = ~new_n19879_ & new_n19884_;
  assign new_n19886_ = ~new_n19875_ & ~new_n19885_;
  assign new_n19887_ = pi0790 & ~new_n19886_;
  assign new_n19888_ = ~pi0790 & ~new_n19858_;
  assign new_n19889_ = pi0832 & ~new_n19888_;
  assign new_n19890_ = ~new_n19887_ & new_n19889_;
  assign po0300 = ~new_n19682_ & ~new_n19890_;
  assign new_n19892_ = pi0144 & ~new_n3272_;
  assign new_n19893_ = ~pi0758 & ~new_n17347_;
  assign new_n19894_ = pi0758 & new_n17391_;
  assign new_n19895_ = ~new_n19893_ & ~new_n19894_;
  assign new_n19896_ = pi0039 & ~new_n19895_;
  assign new_n19897_ = pi0758 & new_n17226_;
  assign new_n19898_ = ~pi0758 & new_n17260_;
  assign new_n19899_ = ~pi0039 & ~new_n19898_;
  assign new_n19900_ = ~new_n19897_ & new_n19899_;
  assign new_n19901_ = ~new_n19896_ & ~new_n19900_;
  assign new_n19902_ = pi0144 & ~new_n19901_;
  assign new_n19903_ = ~pi0144 & pi0758;
  assign new_n19904_ = new_n17426_ & new_n19903_;
  assign new_n19905_ = ~new_n19902_ & ~new_n19904_;
  assign new_n19906_ = ~pi0038 & ~new_n19905_;
  assign new_n19907_ = pi0758 & new_n16639_;
  assign new_n19908_ = new_n17431_ & ~new_n19907_;
  assign new_n19909_ = ~pi0144 & ~new_n17431_;
  assign new_n19910_ = pi0038 & ~new_n19909_;
  assign new_n19911_ = ~new_n19908_ & new_n19910_;
  assign new_n19912_ = ~new_n19906_ & ~new_n19911_;
  assign new_n19913_ = ~pi0736 & new_n19912_;
  assign new_n19914_ = pi0144 & ~new_n16810_;
  assign new_n19915_ = ~pi0144 & ~new_n16928_;
  assign new_n19916_ = ~pi0758 & ~new_n19915_;
  assign new_n19917_ = ~new_n19914_ & new_n19916_;
  assign new_n19918_ = ~pi0144 & ~new_n17007_;
  assign new_n19919_ = pi0144 & new_n17074_;
  assign new_n19920_ = pi0758 & ~new_n19919_;
  assign new_n19921_ = ~new_n19918_ & new_n19920_;
  assign new_n19922_ = pi0039 & ~new_n19921_;
  assign new_n19923_ = ~new_n19917_ & new_n19922_;
  assign new_n19924_ = pi0144 & ~new_n17217_;
  assign new_n19925_ = ~pi0144 & ~new_n17178_;
  assign new_n19926_ = ~pi0758 & ~new_n19925_;
  assign new_n19927_ = ~new_n19924_ & new_n19926_;
  assign new_n19928_ = pi0144 & new_n17227_;
  assign new_n19929_ = ~pi0144 & new_n17234_;
  assign new_n19930_ = pi0758 & ~new_n19929_;
  assign new_n19931_ = ~new_n19928_ & new_n19930_;
  assign new_n19932_ = ~pi0039 & ~new_n19931_;
  assign new_n19933_ = ~new_n19927_ & new_n19932_;
  assign new_n19934_ = ~pi0038 & ~new_n19933_;
  assign new_n19935_ = ~new_n19923_ & new_n19934_;
  assign new_n19936_ = pi0736 & ~new_n19396_;
  assign new_n19937_ = ~new_n19911_ & new_n19936_;
  assign new_n19938_ = ~new_n19935_ & new_n19937_;
  assign new_n19939_ = new_n3272_ & ~new_n19938_;
  assign new_n19940_ = ~new_n19913_ & new_n19939_;
  assign new_n19941_ = ~new_n19892_ & ~new_n19940_;
  assign new_n19942_ = ~pi0625 & new_n19941_;
  assign new_n19943_ = new_n3272_ & ~new_n19912_;
  assign new_n19944_ = ~new_n19892_ & ~new_n19943_;
  assign new_n19945_ = pi0625 & new_n19944_;
  assign new_n19946_ = ~pi1153 & ~new_n19945_;
  assign new_n19947_ = ~new_n19942_ & new_n19946_;
  assign new_n19948_ = pi0144 & ~new_n17558_;
  assign new_n19949_ = pi0736 & new_n3272_;
  assign new_n19950_ = ~new_n19948_ & ~new_n19949_;
  assign new_n19951_ = pi0144 & ~new_n18124_;
  assign new_n19952_ = ~pi0144 & new_n18128_;
  assign new_n19953_ = ~pi0038 & ~new_n19952_;
  assign new_n19954_ = ~new_n19951_ & new_n19953_;
  assign new_n19955_ = ~new_n16914_ & new_n17431_;
  assign new_n19956_ = pi0038 & ~new_n19955_;
  assign new_n19957_ = ~new_n19909_ & new_n19956_;
  assign new_n19958_ = new_n19949_ & ~new_n19957_;
  assign new_n19959_ = ~new_n19954_ & new_n19958_;
  assign new_n19960_ = ~new_n19950_ & ~new_n19959_;
  assign new_n19961_ = pi0625 & ~new_n19960_;
  assign new_n19962_ = ~pi0625 & ~new_n19948_;
  assign new_n19963_ = pi1153 & ~new_n19962_;
  assign new_n19964_ = ~new_n19961_ & new_n19963_;
  assign new_n19965_ = ~pi0608 & ~new_n19964_;
  assign new_n19966_ = ~new_n19947_ & new_n19965_;
  assign new_n19967_ = pi0625 & new_n19941_;
  assign new_n19968_ = ~pi0625 & new_n19944_;
  assign new_n19969_ = pi1153 & ~new_n19968_;
  assign new_n19970_ = ~new_n19967_ & new_n19969_;
  assign new_n19971_ = ~pi0625 & ~new_n19960_;
  assign new_n19972_ = pi0625 & ~new_n19948_;
  assign new_n19973_ = ~pi1153 & ~new_n19972_;
  assign new_n19974_ = ~new_n19971_ & new_n19973_;
  assign new_n19975_ = pi0608 & ~new_n19974_;
  assign new_n19976_ = ~new_n19970_ & new_n19975_;
  assign new_n19977_ = ~new_n19966_ & ~new_n19976_;
  assign new_n19978_ = pi0778 & ~new_n19977_;
  assign new_n19979_ = ~pi0778 & new_n19941_;
  assign new_n19980_ = ~new_n19978_ & ~new_n19979_;
  assign new_n19981_ = ~pi0609 & ~new_n19980_;
  assign new_n19982_ = ~pi0778 & new_n19960_;
  assign new_n19983_ = ~new_n19964_ & ~new_n19974_;
  assign new_n19984_ = pi0778 & ~new_n19983_;
  assign new_n19985_ = ~new_n19982_ & ~new_n19984_;
  assign new_n19986_ = pi0609 & new_n19985_;
  assign new_n19987_ = ~pi1155 & ~new_n19986_;
  assign new_n19988_ = ~new_n19981_ & new_n19987_;
  assign new_n19989_ = new_n17590_ & ~new_n19948_;
  assign new_n19990_ = ~new_n17590_ & new_n19944_;
  assign new_n19991_ = ~new_n19989_ & ~new_n19990_;
  assign new_n19992_ = pi0609 & ~new_n19991_;
  assign new_n19993_ = ~pi0609 & ~new_n19948_;
  assign new_n19994_ = pi1155 & ~new_n19993_;
  assign new_n19995_ = ~new_n19992_ & new_n19994_;
  assign new_n19996_ = ~pi0660 & ~new_n19995_;
  assign new_n19997_ = ~new_n19988_ & new_n19996_;
  assign new_n19998_ = pi0609 & ~new_n19980_;
  assign new_n19999_ = ~pi0609 & new_n19985_;
  assign new_n20000_ = pi1155 & ~new_n19999_;
  assign new_n20001_ = ~new_n19998_ & new_n20000_;
  assign new_n20002_ = ~pi0609 & ~new_n19991_;
  assign new_n20003_ = pi0609 & ~new_n19948_;
  assign new_n20004_ = ~pi1155 & ~new_n20003_;
  assign new_n20005_ = ~new_n20002_ & new_n20004_;
  assign new_n20006_ = pi0660 & ~new_n20005_;
  assign new_n20007_ = ~new_n20001_ & new_n20006_;
  assign new_n20008_ = ~new_n19997_ & ~new_n20007_;
  assign new_n20009_ = pi0785 & ~new_n20008_;
  assign new_n20010_ = ~pi0785 & ~new_n19980_;
  assign new_n20011_ = ~new_n20009_ & ~new_n20010_;
  assign new_n20012_ = ~pi0618 & ~new_n20011_;
  assign new_n20013_ = new_n17618_ & ~new_n19948_;
  assign new_n20014_ = ~new_n17618_ & new_n19985_;
  assign new_n20015_ = ~new_n20013_ & ~new_n20014_;
  assign new_n20016_ = pi0618 & ~new_n20015_;
  assign new_n20017_ = ~pi1154 & ~new_n20016_;
  assign new_n20018_ = ~new_n20012_ & new_n20017_;
  assign new_n20019_ = ~pi0785 & new_n19991_;
  assign new_n20020_ = ~new_n19995_ & ~new_n20005_;
  assign new_n20021_ = pi0785 & ~new_n20020_;
  assign new_n20022_ = ~new_n20019_ & ~new_n20021_;
  assign new_n20023_ = pi0618 & new_n20022_;
  assign new_n20024_ = ~pi0618 & ~new_n19948_;
  assign new_n20025_ = pi1154 & ~new_n20024_;
  assign new_n20026_ = ~new_n20023_ & new_n20025_;
  assign new_n20027_ = ~pi0627 & ~new_n20026_;
  assign new_n20028_ = ~new_n20018_ & new_n20027_;
  assign new_n20029_ = pi0618 & ~new_n20011_;
  assign new_n20030_ = ~pi0618 & ~new_n20015_;
  assign new_n20031_ = pi1154 & ~new_n20030_;
  assign new_n20032_ = ~new_n20029_ & new_n20031_;
  assign new_n20033_ = ~pi0618 & new_n20022_;
  assign new_n20034_ = pi0618 & ~new_n19948_;
  assign new_n20035_ = ~pi1154 & ~new_n20034_;
  assign new_n20036_ = ~new_n20033_ & new_n20035_;
  assign new_n20037_ = pi0627 & ~new_n20036_;
  assign new_n20038_ = ~new_n20032_ & new_n20037_;
  assign new_n20039_ = ~new_n20028_ & ~new_n20038_;
  assign new_n20040_ = pi0781 & ~new_n20039_;
  assign new_n20041_ = ~pi0781 & ~new_n20011_;
  assign new_n20042_ = ~new_n20040_ & ~new_n20041_;
  assign new_n20043_ = ~pi0619 & ~new_n20042_;
  assign new_n20044_ = ~new_n17655_ & new_n20015_;
  assign new_n20045_ = new_n17655_ & new_n19948_;
  assign new_n20046_ = ~new_n20044_ & ~new_n20045_;
  assign new_n20047_ = pi0619 & new_n20046_;
  assign new_n20048_ = ~pi1159 & ~new_n20047_;
  assign new_n20049_ = ~new_n20043_ & new_n20048_;
  assign new_n20050_ = ~pi0781 & ~new_n20022_;
  assign new_n20051_ = ~new_n20026_ & ~new_n20036_;
  assign new_n20052_ = pi0781 & ~new_n20051_;
  assign new_n20053_ = ~new_n20050_ & ~new_n20052_;
  assign new_n20054_ = pi0619 & new_n20053_;
  assign new_n20055_ = ~pi0619 & ~new_n19948_;
  assign new_n20056_ = pi1159 & ~new_n20055_;
  assign new_n20057_ = ~new_n20054_ & new_n20056_;
  assign new_n20058_ = ~pi0648 & ~new_n20057_;
  assign new_n20059_ = ~new_n20049_ & new_n20058_;
  assign new_n20060_ = pi0619 & ~new_n20042_;
  assign new_n20061_ = ~pi0619 & new_n20046_;
  assign new_n20062_ = pi1159 & ~new_n20061_;
  assign new_n20063_ = ~new_n20060_ & new_n20062_;
  assign new_n20064_ = ~pi0619 & new_n20053_;
  assign new_n20065_ = pi0619 & ~new_n19948_;
  assign new_n20066_ = ~pi1159 & ~new_n20065_;
  assign new_n20067_ = ~new_n20064_ & new_n20066_;
  assign new_n20068_ = pi0648 & ~new_n20067_;
  assign new_n20069_ = ~new_n20063_ & new_n20068_;
  assign new_n20070_ = ~new_n20059_ & ~new_n20069_;
  assign new_n20071_ = pi0789 & ~new_n20070_;
  assign new_n20072_ = ~pi0789 & ~new_n20042_;
  assign new_n20073_ = ~new_n20071_ & ~new_n20072_;
  assign new_n20074_ = ~pi0788 & new_n20073_;
  assign new_n20075_ = ~pi0626 & new_n20073_;
  assign new_n20076_ = new_n17691_ & ~new_n19948_;
  assign new_n20077_ = ~new_n17691_ & new_n20046_;
  assign new_n20078_ = ~new_n20076_ & ~new_n20077_;
  assign new_n20079_ = pi0626 & new_n20078_;
  assign new_n20080_ = ~pi0641 & ~new_n20079_;
  assign new_n20081_ = ~new_n20075_ & new_n20080_;
  assign new_n20082_ = ~pi0789 & ~new_n20053_;
  assign new_n20083_ = ~new_n20057_ & ~new_n20067_;
  assign new_n20084_ = pi0789 & ~new_n20083_;
  assign new_n20085_ = ~new_n20082_ & ~new_n20084_;
  assign new_n20086_ = ~pi0626 & new_n20085_;
  assign new_n20087_ = pi0626 & ~new_n19948_;
  assign new_n20088_ = ~pi1158 & ~new_n20087_;
  assign new_n20089_ = ~new_n20086_ & new_n20088_;
  assign new_n20090_ = ~new_n17698_ & ~new_n20089_;
  assign new_n20091_ = ~new_n20081_ & ~new_n20090_;
  assign new_n20092_ = pi0626 & new_n20073_;
  assign new_n20093_ = ~pi0626 & new_n20078_;
  assign new_n20094_ = pi0641 & ~new_n20093_;
  assign new_n20095_ = ~new_n20092_ & new_n20094_;
  assign new_n20096_ = pi0626 & new_n20085_;
  assign new_n20097_ = ~pi0626 & ~new_n19948_;
  assign new_n20098_ = pi1158 & ~new_n20097_;
  assign new_n20099_ = ~new_n20096_ & new_n20098_;
  assign new_n20100_ = ~new_n17713_ & ~new_n20099_;
  assign new_n20101_ = ~new_n20095_ & ~new_n20100_;
  assign new_n20102_ = ~new_n20091_ & ~new_n20101_;
  assign new_n20103_ = pi0788 & ~new_n20102_;
  assign new_n20104_ = ~new_n20074_ & ~new_n20103_;
  assign new_n20105_ = ~pi0628 & new_n20104_;
  assign new_n20106_ = ~new_n20089_ & ~new_n20099_;
  assign new_n20107_ = pi0788 & ~new_n20106_;
  assign new_n20108_ = ~pi0788 & ~new_n20085_;
  assign new_n20109_ = ~new_n20107_ & ~new_n20108_;
  assign new_n20110_ = pi0628 & new_n20109_;
  assign new_n20111_ = ~pi1156 & ~new_n20110_;
  assign new_n20112_ = ~new_n20105_ & new_n20111_;
  assign new_n20113_ = ~new_n17734_ & new_n20078_;
  assign new_n20114_ = new_n17734_ & new_n19948_;
  assign new_n20115_ = ~new_n20113_ & ~new_n20114_;
  assign new_n20116_ = pi0628 & new_n20115_;
  assign new_n20117_ = ~pi0628 & ~new_n19948_;
  assign new_n20118_ = pi1156 & ~new_n20117_;
  assign new_n20119_ = ~new_n20116_ & new_n20118_;
  assign new_n20120_ = ~pi0629 & ~new_n20119_;
  assign new_n20121_ = ~new_n20112_ & new_n20120_;
  assign new_n20122_ = pi0628 & new_n20104_;
  assign new_n20123_ = ~pi0628 & new_n20109_;
  assign new_n20124_ = pi1156 & ~new_n20123_;
  assign new_n20125_ = ~new_n20122_ & new_n20124_;
  assign new_n20126_ = ~pi0628 & new_n20115_;
  assign new_n20127_ = pi0628 & ~new_n19948_;
  assign new_n20128_ = ~pi1156 & ~new_n20127_;
  assign new_n20129_ = ~new_n20126_ & new_n20128_;
  assign new_n20130_ = pi0629 & ~new_n20129_;
  assign new_n20131_ = ~new_n20125_ & new_n20130_;
  assign new_n20132_ = ~new_n20121_ & ~new_n20131_;
  assign new_n20133_ = pi0792 & ~new_n20132_;
  assign new_n20134_ = ~pi0792 & new_n20104_;
  assign new_n20135_ = ~new_n20133_ & ~new_n20134_;
  assign new_n20136_ = ~pi0647 & ~new_n20135_;
  assign new_n20137_ = ~new_n17762_ & ~new_n20109_;
  assign new_n20138_ = new_n17762_ & new_n19948_;
  assign new_n20139_ = ~new_n20137_ & ~new_n20138_;
  assign new_n20140_ = pi0647 & new_n20139_;
  assign new_n20141_ = ~pi1157 & ~new_n20140_;
  assign new_n20142_ = ~new_n20136_ & new_n20141_;
  assign new_n20143_ = ~pi0792 & ~new_n20115_;
  assign new_n20144_ = ~new_n20119_ & ~new_n20129_;
  assign new_n20145_ = pi0792 & ~new_n20144_;
  assign new_n20146_ = ~new_n20143_ & ~new_n20145_;
  assign new_n20147_ = pi0647 & new_n20146_;
  assign new_n20148_ = ~pi0647 & ~new_n19948_;
  assign new_n20149_ = pi1157 & ~new_n20148_;
  assign new_n20150_ = ~new_n20147_ & new_n20149_;
  assign new_n20151_ = ~pi0630 & ~new_n20150_;
  assign new_n20152_ = ~new_n20142_ & new_n20151_;
  assign new_n20153_ = pi0647 & ~new_n20135_;
  assign new_n20154_ = ~pi0647 & new_n20139_;
  assign new_n20155_ = pi1157 & ~new_n20154_;
  assign new_n20156_ = ~new_n20153_ & new_n20155_;
  assign new_n20157_ = ~pi0647 & new_n20146_;
  assign new_n20158_ = pi0647 & ~new_n19948_;
  assign new_n20159_ = ~pi1157 & ~new_n20158_;
  assign new_n20160_ = ~new_n20157_ & new_n20159_;
  assign new_n20161_ = pi0630 & ~new_n20160_;
  assign new_n20162_ = ~new_n20156_ & new_n20161_;
  assign new_n20163_ = ~new_n20152_ & ~new_n20162_;
  assign new_n20164_ = pi0787 & ~new_n20163_;
  assign new_n20165_ = ~pi0787 & ~new_n20135_;
  assign new_n20166_ = ~new_n20164_ & ~new_n20165_;
  assign new_n20167_ = ~pi0644 & ~new_n20166_;
  assign new_n20168_ = ~pi0787 & ~new_n20146_;
  assign new_n20169_ = ~new_n20150_ & ~new_n20160_;
  assign new_n20170_ = pi0787 & ~new_n20169_;
  assign new_n20171_ = ~new_n20168_ & ~new_n20170_;
  assign new_n20172_ = pi0644 & new_n20171_;
  assign new_n20173_ = ~pi0715 & ~new_n20172_;
  assign new_n20174_ = ~new_n20167_ & new_n20173_;
  assign new_n20175_ = new_n17804_ & ~new_n19948_;
  assign new_n20176_ = ~new_n17804_ & new_n20139_;
  assign new_n20177_ = ~new_n20175_ & ~new_n20176_;
  assign new_n20178_ = ~pi0644 & ~new_n20177_;
  assign new_n20179_ = pi0644 & ~new_n19948_;
  assign new_n20180_ = pi0715 & ~new_n20179_;
  assign new_n20181_ = ~new_n20178_ & new_n20180_;
  assign new_n20182_ = ~pi1160 & ~new_n20181_;
  assign new_n20183_ = ~new_n20174_ & new_n20182_;
  assign new_n20184_ = pi0644 & ~new_n20166_;
  assign new_n20185_ = ~pi0644 & new_n20171_;
  assign new_n20186_ = pi0715 & ~new_n20185_;
  assign new_n20187_ = ~new_n20184_ & new_n20186_;
  assign new_n20188_ = pi0644 & ~new_n20177_;
  assign new_n20189_ = ~pi0644 & ~new_n19948_;
  assign new_n20190_ = ~pi0715 & ~new_n20189_;
  assign new_n20191_ = ~new_n20188_ & new_n20190_;
  assign new_n20192_ = pi1160 & ~new_n20191_;
  assign new_n20193_ = ~new_n20187_ & new_n20192_;
  assign new_n20194_ = pi0790 & ~new_n20193_;
  assign new_n20195_ = ~new_n20183_ & new_n20194_;
  assign new_n20196_ = ~pi0790 & new_n20166_;
  assign new_n20197_ = new_n6305_ & ~new_n20196_;
  assign new_n20198_ = ~new_n20195_ & new_n20197_;
  assign new_n20199_ = ~pi0144 & ~new_n6305_;
  assign new_n20200_ = ~pi0057 & ~new_n20199_;
  assign new_n20201_ = ~new_n20198_ & new_n20200_;
  assign new_n20202_ = pi0057 & pi0144;
  assign new_n20203_ = ~pi0832 & ~new_n20202_;
  assign new_n20204_ = ~new_n20201_ & new_n20203_;
  assign new_n20205_ = pi0144 & ~new_n2754_;
  assign new_n20206_ = pi0736 & new_n16915_;
  assign new_n20207_ = ~new_n20205_ & ~new_n20206_;
  assign new_n20208_ = ~pi0778 & new_n20207_;
  assign new_n20209_ = pi0625 & new_n20206_;
  assign new_n20210_ = ~new_n20207_ & ~new_n20209_;
  assign new_n20211_ = ~pi1153 & ~new_n20210_;
  assign new_n20212_ = pi1153 & ~new_n20205_;
  assign new_n20213_ = ~new_n20209_ & new_n20212_;
  assign new_n20214_ = ~new_n20211_ & ~new_n20213_;
  assign new_n20215_ = pi0778 & ~new_n20214_;
  assign new_n20216_ = ~new_n20208_ & ~new_n20215_;
  assign new_n20217_ = new_n19281_ & new_n20216_;
  assign new_n20218_ = ~pi0628 & new_n20217_;
  assign new_n20219_ = pi0629 & ~new_n20218_;
  assign new_n20220_ = pi0609 & pi1155;
  assign new_n20221_ = ~pi0609 & ~pi1155;
  assign new_n20222_ = pi0785 & ~new_n20221_;
  assign new_n20223_ = ~new_n20220_ & new_n20222_;
  assign new_n20224_ = pi0758 & new_n16913_;
  assign new_n20225_ = ~new_n20223_ & new_n20224_;
  assign new_n20226_ = pi0618 & pi1154;
  assign new_n20227_ = ~pi0618 & ~pi1154;
  assign new_n20228_ = pi0781 & ~new_n20227_;
  assign new_n20229_ = ~new_n20226_ & new_n20228_;
  assign new_n20230_ = ~pi0619 & pi1159;
  assign new_n20231_ = pi0619 & ~pi1159;
  assign new_n20232_ = ~new_n20230_ & ~new_n20231_;
  assign new_n20233_ = pi0789 & ~new_n20232_;
  assign new_n20234_ = ~new_n17590_ & ~new_n20233_;
  assign new_n20235_ = ~new_n20229_ & new_n20234_;
  assign new_n20236_ = new_n20225_ & new_n20235_;
  assign new_n20237_ = ~new_n17968_ & new_n20236_;
  assign new_n20238_ = pi0628 & ~new_n20237_;
  assign new_n20239_ = ~new_n20219_ & ~new_n20238_;
  assign new_n20240_ = ~pi1156 & ~new_n20239_;
  assign new_n20241_ = pi0628 & new_n20217_;
  assign new_n20242_ = ~pi0628 & ~new_n20237_;
  assign new_n20243_ = pi0629 & ~new_n20242_;
  assign new_n20244_ = pi1156 & ~new_n20243_;
  assign new_n20245_ = ~new_n20241_ & new_n20244_;
  assign new_n20246_ = ~new_n20240_ & ~new_n20245_;
  assign new_n20247_ = ~new_n20205_ & ~new_n20246_;
  assign new_n20248_ = pi0792 & new_n20247_;
  assign new_n20249_ = new_n17691_ & ~new_n20205_;
  assign new_n20250_ = ~new_n17618_ & new_n20216_;
  assign new_n20251_ = ~new_n17655_ & new_n20250_;
  assign new_n20252_ = ~new_n20205_ & ~new_n20251_;
  assign new_n20253_ = ~new_n20249_ & ~new_n20252_;
  assign new_n20254_ = new_n17851_ & new_n20253_;
  assign new_n20255_ = pi0626 & new_n20236_;
  assign new_n20256_ = ~new_n20205_ & ~new_n20255_;
  assign new_n20257_ = pi1158 & ~new_n20256_;
  assign new_n20258_ = ~pi0641 & ~new_n20257_;
  assign new_n20259_ = ~new_n20254_ & new_n20258_;
  assign new_n20260_ = new_n17850_ & new_n20253_;
  assign new_n20261_ = ~pi0626 & new_n20236_;
  assign new_n20262_ = ~new_n20205_ & ~new_n20261_;
  assign new_n20263_ = ~pi1158 & ~new_n20262_;
  assign new_n20264_ = pi0641 & ~new_n20263_;
  assign new_n20265_ = ~new_n20260_ & new_n20264_;
  assign new_n20266_ = pi0788 & ~new_n20265_;
  assign new_n20267_ = ~new_n20259_ & new_n20266_;
  assign new_n20268_ = ~new_n20205_ & ~new_n20224_;
  assign new_n20269_ = pi0736 & new_n16916_;
  assign new_n20270_ = new_n20268_ & ~new_n20269_;
  assign new_n20271_ = pi0625 & new_n20269_;
  assign new_n20272_ = ~new_n20270_ & ~new_n20271_;
  assign new_n20273_ = ~pi1153 & ~new_n20272_;
  assign new_n20274_ = ~pi0608 & ~new_n20213_;
  assign new_n20275_ = ~new_n20273_ & new_n20274_;
  assign new_n20276_ = pi1153 & new_n20268_;
  assign new_n20277_ = ~new_n20271_ & new_n20276_;
  assign new_n20278_ = pi0608 & ~new_n20211_;
  assign new_n20279_ = ~new_n20277_ & new_n20278_;
  assign new_n20280_ = ~new_n20275_ & ~new_n20279_;
  assign new_n20281_ = pi0778 & ~new_n20280_;
  assign new_n20282_ = ~pi0778 & ~new_n20270_;
  assign new_n20283_ = ~new_n20281_ & ~new_n20282_;
  assign new_n20284_ = ~pi0609 & ~new_n20283_;
  assign new_n20285_ = pi0609 & new_n20216_;
  assign new_n20286_ = ~pi1155 & ~new_n20285_;
  assign new_n20287_ = ~new_n20284_ & new_n20286_;
  assign new_n20288_ = new_n17591_ & new_n20224_;
  assign new_n20289_ = pi1155 & ~new_n20205_;
  assign new_n20290_ = ~new_n20288_ & new_n20289_;
  assign new_n20291_ = ~pi0660 & ~new_n20290_;
  assign new_n20292_ = ~new_n20287_ & new_n20291_;
  assign new_n20293_ = pi0609 & ~new_n20283_;
  assign new_n20294_ = ~pi0609 & new_n20216_;
  assign new_n20295_ = pi1155 & ~new_n20294_;
  assign new_n20296_ = ~new_n20293_ & new_n20295_;
  assign new_n20297_ = new_n17603_ & new_n20224_;
  assign new_n20298_ = ~pi1155 & ~new_n20205_;
  assign new_n20299_ = ~new_n20297_ & new_n20298_;
  assign new_n20300_ = pi0660 & ~new_n20299_;
  assign new_n20301_ = ~new_n20296_ & new_n20300_;
  assign new_n20302_ = ~new_n20292_ & ~new_n20301_;
  assign new_n20303_ = pi0785 & ~new_n20302_;
  assign new_n20304_ = ~pi0785 & ~new_n20283_;
  assign new_n20305_ = ~new_n20303_ & ~new_n20304_;
  assign new_n20306_ = ~pi0618 & ~new_n20305_;
  assign new_n20307_ = ~new_n20205_ & ~new_n20250_;
  assign new_n20308_ = pi0618 & ~new_n20307_;
  assign new_n20309_ = ~pi1154 & ~new_n20308_;
  assign new_n20310_ = ~new_n20306_ & new_n20309_;
  assign new_n20311_ = pi0618 & ~new_n17590_;
  assign new_n20312_ = new_n20225_ & new_n20311_;
  assign new_n20313_ = pi1154 & ~new_n20205_;
  assign new_n20314_ = ~new_n20312_ & new_n20313_;
  assign new_n20315_ = ~pi0627 & ~new_n20314_;
  assign new_n20316_ = ~new_n20310_ & new_n20315_;
  assign new_n20317_ = pi0618 & ~new_n20305_;
  assign new_n20318_ = ~pi0618 & ~new_n20307_;
  assign new_n20319_ = pi1154 & ~new_n20318_;
  assign new_n20320_ = ~new_n20317_ & new_n20319_;
  assign new_n20321_ = ~pi0618 & ~new_n17590_;
  assign new_n20322_ = new_n20225_ & new_n20321_;
  assign new_n20323_ = ~pi1154 & ~new_n20205_;
  assign new_n20324_ = ~new_n20322_ & new_n20323_;
  assign new_n20325_ = pi0627 & ~new_n20324_;
  assign new_n20326_ = ~new_n20320_ & new_n20325_;
  assign new_n20327_ = ~new_n20316_ & ~new_n20326_;
  assign new_n20328_ = pi0781 & ~new_n20327_;
  assign new_n20329_ = ~pi0781 & ~new_n20305_;
  assign new_n20330_ = ~new_n20328_ & ~new_n20329_;
  assign new_n20331_ = pi0619 & ~new_n20330_;
  assign new_n20332_ = ~pi0619 & ~new_n20252_;
  assign new_n20333_ = pi1159 & ~new_n20332_;
  assign new_n20334_ = ~new_n20331_ & new_n20333_;
  assign new_n20335_ = new_n20225_ & ~new_n20229_;
  assign new_n20336_ = ~pi0619 & ~new_n17590_;
  assign new_n20337_ = new_n20335_ & new_n20336_;
  assign new_n20338_ = ~pi1159 & ~new_n20205_;
  assign new_n20339_ = ~new_n20337_ & new_n20338_;
  assign new_n20340_ = pi0648 & ~new_n20339_;
  assign new_n20341_ = ~new_n20334_ & new_n20340_;
  assign new_n20342_ = ~pi0619 & ~new_n20330_;
  assign new_n20343_ = pi0619 & ~new_n20252_;
  assign new_n20344_ = ~pi1159 & ~new_n20343_;
  assign new_n20345_ = ~new_n20342_ & new_n20344_;
  assign new_n20346_ = pi0619 & ~new_n17590_;
  assign new_n20347_ = new_n20335_ & new_n20346_;
  assign new_n20348_ = pi1159 & ~new_n20205_;
  assign new_n20349_ = ~new_n20347_ & new_n20348_;
  assign new_n20350_ = ~pi0648 & ~new_n20349_;
  assign new_n20351_ = ~new_n20345_ & new_n20350_;
  assign new_n20352_ = pi0789 & ~new_n20351_;
  assign new_n20353_ = ~new_n20341_ & new_n20352_;
  assign new_n20354_ = ~pi0789 & new_n20330_;
  assign new_n20355_ = new_n17969_ & ~new_n20354_;
  assign new_n20356_ = ~new_n20353_ & new_n20355_;
  assign new_n20357_ = ~new_n20267_ & ~new_n20356_;
  assign new_n20358_ = ~new_n20248_ & ~new_n20357_;
  assign new_n20359_ = new_n17803_ & new_n19334_;
  assign new_n20360_ = pi0787 & ~new_n20359_;
  assign new_n20361_ = ~pi0629 & new_n19308_;
  assign new_n20362_ = pi0629 & new_n19309_;
  assign new_n20363_ = pi0792 & ~new_n20362_;
  assign new_n20364_ = ~new_n20361_ & new_n20363_;
  assign new_n20365_ = ~new_n20247_ & new_n20364_;
  assign new_n20366_ = ~new_n20360_ & ~new_n20365_;
  assign new_n20367_ = ~new_n20358_ & new_n20366_;
  assign new_n20368_ = ~new_n17762_ & new_n20237_;
  assign new_n20369_ = ~pi0630 & new_n20368_;
  assign new_n20370_ = pi0647 & ~new_n20369_;
  assign new_n20371_ = ~new_n19311_ & new_n20217_;
  assign new_n20372_ = pi0630 & ~new_n20371_;
  assign new_n20373_ = ~new_n20370_ & ~new_n20372_;
  assign new_n20374_ = ~pi1157 & ~new_n20373_;
  assign new_n20375_ = ~pi0630 & ~new_n20371_;
  assign new_n20376_ = pi0647 & ~new_n20375_;
  assign new_n20377_ = pi0630 & new_n20368_;
  assign new_n20378_ = pi1157 & ~new_n20377_;
  assign new_n20379_ = ~new_n20376_ & new_n20378_;
  assign new_n20380_ = ~new_n20374_ & ~new_n20379_;
  assign new_n20381_ = pi0787 & ~new_n20205_;
  assign new_n20382_ = ~new_n20380_ & new_n20381_;
  assign new_n20383_ = ~new_n20367_ & ~new_n20382_;
  assign new_n20384_ = pi0644 & new_n20383_;
  assign new_n20385_ = ~new_n19335_ & new_n20371_;
  assign new_n20386_ = ~new_n20205_ & ~new_n20385_;
  assign new_n20387_ = ~pi0644 & ~new_n20386_;
  assign new_n20388_ = pi0715 & ~new_n20387_;
  assign new_n20389_ = ~new_n20384_ & new_n20388_;
  assign new_n20390_ = ~new_n17804_ & new_n20368_;
  assign new_n20391_ = pi0644 & new_n20390_;
  assign new_n20392_ = ~pi0715 & ~new_n20205_;
  assign new_n20393_ = ~new_n20391_ & new_n20392_;
  assign new_n20394_ = pi1160 & ~new_n20393_;
  assign new_n20395_ = ~new_n20389_ & new_n20394_;
  assign new_n20396_ = ~pi0644 & new_n20383_;
  assign new_n20397_ = pi0644 & ~new_n20386_;
  assign new_n20398_ = ~pi0715 & ~new_n20397_;
  assign new_n20399_ = ~new_n20396_ & new_n20398_;
  assign new_n20400_ = ~pi0644 & new_n20390_;
  assign new_n20401_ = pi0715 & ~new_n20205_;
  assign new_n20402_ = ~new_n20400_ & new_n20401_;
  assign new_n20403_ = ~pi1160 & ~new_n20402_;
  assign new_n20404_ = ~new_n20399_ & new_n20403_;
  assign new_n20405_ = ~new_n20395_ & ~new_n20404_;
  assign new_n20406_ = pi0790 & ~new_n20405_;
  assign new_n20407_ = ~pi0790 & new_n20383_;
  assign new_n20408_ = pi0832 & ~new_n20407_;
  assign new_n20409_ = ~new_n20406_ & new_n20408_;
  assign po0301 = ~new_n20204_ & ~new_n20409_;
  assign new_n20411_ = ~pi0145 & ~new_n17558_;
  assign new_n20412_ = new_n17691_ & ~new_n20411_;
  assign new_n20413_ = ~pi0698 & new_n3272_;
  assign new_n20414_ = new_n20411_ & ~new_n20413_;
  assign new_n20415_ = pi0145 & ~new_n18128_;
  assign new_n20416_ = ~pi0038 & ~new_n20415_;
  assign new_n20417_ = new_n3272_ & ~new_n20416_;
  assign new_n20418_ = ~pi0145 & new_n18124_;
  assign new_n20419_ = ~new_n20417_ & ~new_n20418_;
  assign new_n20420_ = ~pi0145 & ~new_n17431_;
  assign new_n20421_ = new_n17544_ & ~new_n20420_;
  assign new_n20422_ = ~pi0698 & ~new_n20421_;
  assign new_n20423_ = ~new_n20419_ & new_n20422_;
  assign new_n20424_ = ~new_n20414_ & ~new_n20423_;
  assign new_n20425_ = ~pi0778 & new_n20424_;
  assign new_n20426_ = pi0625 & ~new_n20424_;
  assign new_n20427_ = ~pi0625 & new_n20411_;
  assign new_n20428_ = pi1153 & ~new_n20427_;
  assign new_n20429_ = ~new_n20426_ & new_n20428_;
  assign new_n20430_ = ~pi0625 & ~new_n20424_;
  assign new_n20431_ = pi0625 & new_n20411_;
  assign new_n20432_ = ~pi1153 & ~new_n20431_;
  assign new_n20433_ = ~new_n20430_ & new_n20432_;
  assign new_n20434_ = ~new_n20429_ & ~new_n20433_;
  assign new_n20435_ = pi0778 & ~new_n20434_;
  assign new_n20436_ = ~new_n20425_ & ~new_n20435_;
  assign new_n20437_ = ~new_n17618_ & ~new_n20436_;
  assign new_n20438_ = new_n17618_ & ~new_n20411_;
  assign new_n20439_ = ~new_n20437_ & ~new_n20438_;
  assign new_n20440_ = ~new_n17655_ & new_n20439_;
  assign new_n20441_ = new_n17655_ & new_n20411_;
  assign new_n20442_ = ~new_n20440_ & ~new_n20441_;
  assign new_n20443_ = ~new_n17691_ & new_n20442_;
  assign new_n20444_ = ~new_n20412_ & ~new_n20443_;
  assign new_n20445_ = ~new_n17734_ & new_n20444_;
  assign new_n20446_ = new_n17734_ & new_n20411_;
  assign new_n20447_ = ~new_n20445_ & ~new_n20446_;
  assign new_n20448_ = ~pi0792 & new_n20447_;
  assign new_n20449_ = pi0628 & ~new_n20447_;
  assign new_n20450_ = ~pi0628 & new_n20411_;
  assign new_n20451_ = pi1156 & ~new_n20450_;
  assign new_n20452_ = ~new_n20449_ & new_n20451_;
  assign new_n20453_ = ~pi0628 & ~new_n20447_;
  assign new_n20454_ = pi0628 & new_n20411_;
  assign new_n20455_ = ~pi1156 & ~new_n20454_;
  assign new_n20456_ = ~new_n20453_ & new_n20455_;
  assign new_n20457_ = ~new_n20452_ & ~new_n20456_;
  assign new_n20458_ = pi0792 & ~new_n20457_;
  assign new_n20459_ = ~new_n20448_ & ~new_n20458_;
  assign new_n20460_ = ~pi0647 & ~new_n20459_;
  assign new_n20461_ = pi0647 & ~new_n20411_;
  assign new_n20462_ = ~new_n20460_ & ~new_n20461_;
  assign new_n20463_ = ~pi1157 & new_n20462_;
  assign new_n20464_ = pi0647 & ~new_n20459_;
  assign new_n20465_ = ~pi0647 & ~new_n20411_;
  assign new_n20466_ = ~new_n20464_ & ~new_n20465_;
  assign new_n20467_ = pi1157 & new_n20466_;
  assign new_n20468_ = ~new_n20463_ & ~new_n20467_;
  assign new_n20469_ = pi0787 & ~new_n20468_;
  assign new_n20470_ = ~pi0787 & new_n20459_;
  assign new_n20471_ = ~new_n20469_ & ~new_n20470_;
  assign new_n20472_ = ~pi0644 & ~new_n20471_;
  assign new_n20473_ = pi0715 & ~new_n20472_;
  assign new_n20474_ = pi0145 & ~new_n3272_;
  assign new_n20475_ = ~pi0145 & ~new_n17349_;
  assign new_n20476_ = pi0767 & ~new_n20475_;
  assign new_n20477_ = pi0145 & ~new_n17426_;
  assign new_n20478_ = ~pi0145 & ~pi0767;
  assign new_n20479_ = new_n17393_ & new_n20478_;
  assign new_n20480_ = ~new_n20477_ & ~new_n20479_;
  assign new_n20481_ = ~new_n20476_ & new_n20480_;
  assign new_n20482_ = ~pi0038 & ~new_n20481_;
  assign new_n20483_ = ~pi0767 & new_n17433_;
  assign new_n20484_ = pi0038 & ~new_n20420_;
  assign new_n20485_ = ~new_n20483_ & new_n20484_;
  assign new_n20486_ = ~new_n20482_ & ~new_n20485_;
  assign new_n20487_ = new_n3272_ & ~new_n20486_;
  assign new_n20488_ = ~new_n20474_ & ~new_n20487_;
  assign new_n20489_ = ~new_n17590_ & ~new_n20488_;
  assign new_n20490_ = new_n17590_ & ~new_n20411_;
  assign new_n20491_ = ~new_n20489_ & ~new_n20490_;
  assign new_n20492_ = ~pi0785 & ~new_n20491_;
  assign new_n20493_ = ~new_n17591_ & ~new_n20411_;
  assign new_n20494_ = pi0609 & new_n20489_;
  assign new_n20495_ = ~new_n20493_ & ~new_n20494_;
  assign new_n20496_ = pi1155 & ~new_n20495_;
  assign new_n20497_ = ~new_n17603_ & ~new_n20411_;
  assign new_n20498_ = ~pi0609 & new_n20489_;
  assign new_n20499_ = ~new_n20497_ & ~new_n20498_;
  assign new_n20500_ = ~pi1155 & ~new_n20499_;
  assign new_n20501_ = ~new_n20496_ & ~new_n20500_;
  assign new_n20502_ = pi0785 & ~new_n20501_;
  assign new_n20503_ = ~new_n20492_ & ~new_n20502_;
  assign new_n20504_ = ~pi0781 & ~new_n20503_;
  assign new_n20505_ = pi0618 & new_n20503_;
  assign new_n20506_ = ~pi0618 & new_n20411_;
  assign new_n20507_ = pi1154 & ~new_n20506_;
  assign new_n20508_ = ~new_n20505_ & new_n20507_;
  assign new_n20509_ = ~pi0618 & new_n20503_;
  assign new_n20510_ = pi0618 & new_n20411_;
  assign new_n20511_ = ~pi1154 & ~new_n20510_;
  assign new_n20512_ = ~new_n20509_ & new_n20511_;
  assign new_n20513_ = ~new_n20508_ & ~new_n20512_;
  assign new_n20514_ = pi0781 & ~new_n20513_;
  assign new_n20515_ = ~new_n20504_ & ~new_n20514_;
  assign new_n20516_ = ~pi0789 & ~new_n20515_;
  assign new_n20517_ = pi0619 & new_n20515_;
  assign new_n20518_ = ~pi0619 & new_n20411_;
  assign new_n20519_ = pi1159 & ~new_n20518_;
  assign new_n20520_ = ~new_n20517_ & new_n20519_;
  assign new_n20521_ = ~pi0619 & new_n20515_;
  assign new_n20522_ = pi0619 & new_n20411_;
  assign new_n20523_ = ~pi1159 & ~new_n20522_;
  assign new_n20524_ = ~new_n20521_ & new_n20523_;
  assign new_n20525_ = ~new_n20520_ & ~new_n20524_;
  assign new_n20526_ = pi0789 & ~new_n20525_;
  assign new_n20527_ = ~new_n20516_ & ~new_n20526_;
  assign new_n20528_ = ~pi0788 & ~new_n20527_;
  assign new_n20529_ = pi0626 & new_n20527_;
  assign new_n20530_ = ~pi0626 & new_n20411_;
  assign new_n20531_ = pi1158 & ~new_n20530_;
  assign new_n20532_ = ~new_n20529_ & new_n20531_;
  assign new_n20533_ = ~pi0626 & new_n20527_;
  assign new_n20534_ = pi0626 & new_n20411_;
  assign new_n20535_ = ~pi1158 & ~new_n20534_;
  assign new_n20536_ = ~new_n20533_ & new_n20535_;
  assign new_n20537_ = ~new_n20532_ & ~new_n20536_;
  assign new_n20538_ = pi0788 & ~new_n20537_;
  assign new_n20539_ = ~new_n20528_ & ~new_n20538_;
  assign new_n20540_ = ~new_n17762_ & new_n20539_;
  assign new_n20541_ = new_n17762_ & new_n20411_;
  assign new_n20542_ = ~new_n20540_ & ~new_n20541_;
  assign new_n20543_ = ~new_n17804_ & ~new_n20542_;
  assign new_n20544_ = new_n17804_ & new_n20411_;
  assign new_n20545_ = ~new_n20543_ & ~new_n20544_;
  assign new_n20546_ = pi0644 & ~new_n20545_;
  assign new_n20547_ = ~pi0644 & new_n20411_;
  assign new_n20548_ = ~pi0715 & ~new_n20547_;
  assign new_n20549_ = ~new_n20546_ & new_n20548_;
  assign new_n20550_ = pi1160 & ~new_n20549_;
  assign new_n20551_ = ~new_n20473_ & new_n20550_;
  assign new_n20552_ = pi0630 & ~pi0647;
  assign new_n20553_ = pi1157 & new_n20552_;
  assign new_n20554_ = ~pi0630 & pi0647;
  assign new_n20555_ = ~pi1157 & new_n20554_;
  assign new_n20556_ = ~new_n20553_ & ~new_n20555_;
  assign new_n20557_ = new_n20542_ & ~new_n20556_;
  assign new_n20558_ = new_n17802_ & ~new_n20462_;
  assign new_n20559_ = new_n17801_ & ~new_n20466_;
  assign new_n20560_ = ~new_n20558_ & ~new_n20559_;
  assign new_n20561_ = ~new_n20557_ & new_n20560_;
  assign new_n20562_ = pi0787 & ~new_n20561_;
  assign new_n20563_ = ~pi0628 & pi0629;
  assign new_n20564_ = pi1156 & new_n20563_;
  assign new_n20565_ = pi0628 & ~pi0629;
  assign new_n20566_ = ~pi1156 & new_n20565_;
  assign new_n20567_ = ~new_n20564_ & ~new_n20566_;
  assign new_n20568_ = ~new_n20539_ & ~new_n20567_;
  assign new_n20569_ = ~pi0629 & new_n20452_;
  assign new_n20570_ = pi0629 & new_n20456_;
  assign new_n20571_ = ~new_n20569_ & ~new_n20570_;
  assign new_n20572_ = ~new_n20568_ & new_n20571_;
  assign new_n20573_ = pi0792 & ~new_n20572_;
  assign new_n20574_ = pi0698 & new_n20486_;
  assign new_n20575_ = ~pi0145 & new_n16810_;
  assign new_n20576_ = pi0145 & new_n16928_;
  assign new_n20577_ = pi0767 & ~new_n20576_;
  assign new_n20578_ = ~new_n20575_ & new_n20577_;
  assign new_n20579_ = pi0145 & new_n17007_;
  assign new_n20580_ = ~pi0145 & ~new_n17074_;
  assign new_n20581_ = ~pi0767 & ~new_n20580_;
  assign new_n20582_ = ~new_n20579_ & new_n20581_;
  assign new_n20583_ = pi0039 & ~new_n20582_;
  assign new_n20584_ = ~new_n20578_ & new_n20583_;
  assign new_n20585_ = ~pi0145 & ~new_n17217_;
  assign new_n20586_ = pi0145 & ~new_n17178_;
  assign new_n20587_ = pi0767 & ~new_n20586_;
  assign new_n20588_ = ~new_n20585_ & new_n20587_;
  assign new_n20589_ = ~pi0145 & new_n17227_;
  assign new_n20590_ = pi0145 & new_n17234_;
  assign new_n20591_ = ~pi0767 & ~new_n20590_;
  assign new_n20592_ = ~new_n20589_ & new_n20591_;
  assign new_n20593_ = ~new_n20588_ & ~new_n20592_;
  assign new_n20594_ = ~pi0039 & ~new_n20593_;
  assign new_n20595_ = ~pi0038 & ~new_n20594_;
  assign new_n20596_ = ~new_n20584_ & new_n20595_;
  assign new_n20597_ = ~pi0767 & ~new_n17035_;
  assign new_n20598_ = new_n19383_ & ~new_n20597_;
  assign new_n20599_ = ~pi0145 & ~new_n20598_;
  assign new_n20600_ = ~pi0767 & new_n16913_;
  assign new_n20601_ = ~new_n16916_ & ~new_n20600_;
  assign new_n20602_ = pi0145 & ~new_n20601_;
  assign new_n20603_ = new_n6257_ & new_n20602_;
  assign new_n20604_ = pi0038 & ~new_n20603_;
  assign new_n20605_ = ~new_n20599_ & new_n20604_;
  assign new_n20606_ = ~pi0698 & ~new_n20605_;
  assign new_n20607_ = ~new_n20596_ & new_n20606_;
  assign new_n20608_ = new_n3272_ & ~new_n20607_;
  assign new_n20609_ = ~new_n20574_ & new_n20608_;
  assign new_n20610_ = ~new_n20474_ & ~new_n20609_;
  assign new_n20611_ = ~pi0625 & new_n20610_;
  assign new_n20612_ = pi0625 & new_n20488_;
  assign new_n20613_ = ~pi1153 & ~new_n20612_;
  assign new_n20614_ = ~new_n20611_ & new_n20613_;
  assign new_n20615_ = ~pi0608 & ~new_n20429_;
  assign new_n20616_ = ~new_n20614_ & new_n20615_;
  assign new_n20617_ = pi0625 & new_n20610_;
  assign new_n20618_ = ~pi0625 & new_n20488_;
  assign new_n20619_ = pi1153 & ~new_n20618_;
  assign new_n20620_ = ~new_n20617_ & new_n20619_;
  assign new_n20621_ = pi0608 & ~new_n20433_;
  assign new_n20622_ = ~new_n20620_ & new_n20621_;
  assign new_n20623_ = ~new_n20616_ & ~new_n20622_;
  assign new_n20624_ = pi0778 & ~new_n20623_;
  assign new_n20625_ = ~pi0778 & new_n20610_;
  assign new_n20626_ = ~new_n20624_ & ~new_n20625_;
  assign new_n20627_ = ~pi0609 & ~new_n20626_;
  assign new_n20628_ = pi0609 & new_n20436_;
  assign new_n20629_ = ~pi1155 & ~new_n20628_;
  assign new_n20630_ = ~new_n20627_ & new_n20629_;
  assign new_n20631_ = ~pi0660 & ~new_n20496_;
  assign new_n20632_ = ~new_n20630_ & new_n20631_;
  assign new_n20633_ = pi0609 & ~new_n20626_;
  assign new_n20634_ = ~pi0609 & new_n20436_;
  assign new_n20635_ = pi1155 & ~new_n20634_;
  assign new_n20636_ = ~new_n20633_ & new_n20635_;
  assign new_n20637_ = pi0660 & ~new_n20500_;
  assign new_n20638_ = ~new_n20636_ & new_n20637_;
  assign new_n20639_ = ~new_n20632_ & ~new_n20638_;
  assign new_n20640_ = pi0785 & ~new_n20639_;
  assign new_n20641_ = ~pi0785 & ~new_n20626_;
  assign new_n20642_ = ~new_n20640_ & ~new_n20641_;
  assign new_n20643_ = ~pi0618 & ~new_n20642_;
  assign new_n20644_ = pi0618 & new_n20439_;
  assign new_n20645_ = ~pi1154 & ~new_n20644_;
  assign new_n20646_ = ~new_n20643_ & new_n20645_;
  assign new_n20647_ = ~pi0627 & ~new_n20508_;
  assign new_n20648_ = ~new_n20646_ & new_n20647_;
  assign new_n20649_ = pi0618 & ~new_n20642_;
  assign new_n20650_ = ~pi0618 & new_n20439_;
  assign new_n20651_ = pi1154 & ~new_n20650_;
  assign new_n20652_ = ~new_n20649_ & new_n20651_;
  assign new_n20653_ = pi0627 & ~new_n20512_;
  assign new_n20654_ = ~new_n20652_ & new_n20653_;
  assign new_n20655_ = ~new_n20648_ & ~new_n20654_;
  assign new_n20656_ = pi0781 & ~new_n20655_;
  assign new_n20657_ = ~pi0781 & ~new_n20642_;
  assign new_n20658_ = ~new_n20656_ & ~new_n20657_;
  assign new_n20659_ = pi0619 & ~new_n20658_;
  assign new_n20660_ = ~pi0619 & ~new_n20442_;
  assign new_n20661_ = pi1159 & ~new_n20660_;
  assign new_n20662_ = ~new_n20659_ & new_n20661_;
  assign new_n20663_ = pi0648 & ~new_n20524_;
  assign new_n20664_ = ~new_n20662_ & new_n20663_;
  assign new_n20665_ = ~pi0619 & ~new_n20658_;
  assign new_n20666_ = pi0619 & ~new_n20442_;
  assign new_n20667_ = ~pi1159 & ~new_n20666_;
  assign new_n20668_ = ~new_n20665_ & new_n20667_;
  assign new_n20669_ = ~pi0648 & ~new_n20520_;
  assign new_n20670_ = ~new_n20668_ & new_n20669_;
  assign new_n20671_ = pi0789 & ~new_n20670_;
  assign new_n20672_ = ~new_n20664_ & new_n20671_;
  assign new_n20673_ = ~pi0789 & new_n20658_;
  assign new_n20674_ = new_n17969_ & ~new_n20673_;
  assign new_n20675_ = ~new_n20672_ & new_n20674_;
  assign new_n20676_ = new_n17856_ & new_n20444_;
  assign new_n20677_ = ~new_n17733_ & new_n20537_;
  assign new_n20678_ = ~new_n20676_ & ~new_n20677_;
  assign new_n20679_ = pi0788 & ~new_n20678_;
  assign new_n20680_ = ~new_n20364_ & ~new_n20679_;
  assign new_n20681_ = ~new_n20675_ & new_n20680_;
  assign new_n20682_ = ~new_n20573_ & ~new_n20681_;
  assign new_n20683_ = ~new_n20360_ & ~new_n20682_;
  assign new_n20684_ = ~new_n20562_ & ~new_n20683_;
  assign new_n20685_ = ~pi0644 & new_n20684_;
  assign new_n20686_ = pi0644 & ~new_n20471_;
  assign new_n20687_ = ~pi0715 & ~new_n20686_;
  assign new_n20688_ = ~new_n20685_ & new_n20687_;
  assign new_n20689_ = ~pi0644 & ~new_n20545_;
  assign new_n20690_ = pi0644 & new_n20411_;
  assign new_n20691_ = pi0715 & ~new_n20690_;
  assign new_n20692_ = ~new_n20689_ & new_n20691_;
  assign new_n20693_ = ~pi1160 & ~new_n20692_;
  assign new_n20694_ = ~new_n20688_ & new_n20693_;
  assign new_n20695_ = ~new_n20551_ & ~new_n20694_;
  assign new_n20696_ = pi0790 & ~new_n20695_;
  assign new_n20697_ = pi0644 & new_n20550_;
  assign new_n20698_ = pi0790 & ~new_n20697_;
  assign new_n20699_ = new_n20684_ & ~new_n20698_;
  assign new_n20700_ = ~new_n20696_ & ~new_n20699_;
  assign new_n20701_ = ~po1038 & ~new_n20700_;
  assign new_n20702_ = ~pi0145 & po1038;
  assign new_n20703_ = ~pi0832 & ~new_n20702_;
  assign new_n20704_ = ~new_n20701_ & new_n20703_;
  assign new_n20705_ = ~pi0145 & ~new_n2754_;
  assign new_n20706_ = ~new_n20600_ & ~new_n20705_;
  assign new_n20707_ = ~new_n17858_ & ~new_n20706_;
  assign new_n20708_ = ~pi0785 & ~new_n20707_;
  assign new_n20709_ = ~new_n17863_ & ~new_n20706_;
  assign new_n20710_ = pi1155 & ~new_n20709_;
  assign new_n20711_ = ~new_n17866_ & new_n20707_;
  assign new_n20712_ = ~pi1155 & ~new_n20711_;
  assign new_n20713_ = ~new_n20710_ & ~new_n20712_;
  assign new_n20714_ = pi0785 & ~new_n20713_;
  assign new_n20715_ = ~new_n20708_ & ~new_n20714_;
  assign new_n20716_ = ~pi0781 & ~new_n20715_;
  assign new_n20717_ = ~new_n17873_ & new_n20715_;
  assign new_n20718_ = pi1154 & ~new_n20717_;
  assign new_n20719_ = ~new_n17876_ & new_n20715_;
  assign new_n20720_ = ~pi1154 & ~new_n20719_;
  assign new_n20721_ = ~new_n20718_ & ~new_n20720_;
  assign new_n20722_ = pi0781 & ~new_n20721_;
  assign new_n20723_ = ~new_n20716_ & ~new_n20722_;
  assign new_n20724_ = ~pi0789 & ~new_n20723_;
  assign new_n20725_ = pi0619 & new_n20723_;
  assign new_n20726_ = ~pi0619 & new_n20705_;
  assign new_n20727_ = pi1159 & ~new_n20726_;
  assign new_n20728_ = ~new_n20725_ & new_n20727_;
  assign new_n20729_ = ~pi0619 & new_n20723_;
  assign new_n20730_ = pi0619 & new_n20705_;
  assign new_n20731_ = ~pi1159 & ~new_n20730_;
  assign new_n20732_ = ~new_n20729_ & new_n20731_;
  assign new_n20733_ = ~new_n20728_ & ~new_n20732_;
  assign new_n20734_ = pi0789 & ~new_n20733_;
  assign new_n20735_ = ~new_n20724_ & ~new_n20734_;
  assign new_n20736_ = ~pi0788 & ~new_n20735_;
  assign new_n20737_ = pi0626 & new_n20735_;
  assign new_n20738_ = ~pi0626 & new_n20705_;
  assign new_n20739_ = pi1158 & ~new_n20738_;
  assign new_n20740_ = ~new_n20737_ & new_n20739_;
  assign new_n20741_ = ~pi0626 & new_n20735_;
  assign new_n20742_ = pi0626 & new_n20705_;
  assign new_n20743_ = ~pi1158 & ~new_n20742_;
  assign new_n20744_ = ~new_n20741_ & new_n20743_;
  assign new_n20745_ = ~new_n20740_ & ~new_n20744_;
  assign new_n20746_ = pi0788 & ~new_n20745_;
  assign new_n20747_ = ~new_n20736_ & ~new_n20746_;
  assign new_n20748_ = ~new_n17762_ & new_n20747_;
  assign new_n20749_ = new_n17762_ & new_n20705_;
  assign new_n20750_ = ~new_n20748_ & ~new_n20749_;
  assign new_n20751_ = ~new_n20556_ & new_n20750_;
  assign new_n20752_ = ~pi0698 & new_n16915_;
  assign new_n20753_ = ~new_n20705_ & ~new_n20752_;
  assign new_n20754_ = ~pi0778 & new_n20753_;
  assign new_n20755_ = ~pi0625 & new_n20752_;
  assign new_n20756_ = ~new_n20753_ & ~new_n20755_;
  assign new_n20757_ = pi1153 & ~new_n20756_;
  assign new_n20758_ = ~pi1153 & ~new_n20705_;
  assign new_n20759_ = ~new_n20755_ & new_n20758_;
  assign new_n20760_ = ~new_n20757_ & ~new_n20759_;
  assign new_n20761_ = pi0778 & ~new_n20760_;
  assign new_n20762_ = ~new_n20754_ & ~new_n20761_;
  assign new_n20763_ = ~new_n17844_ & new_n20762_;
  assign new_n20764_ = ~new_n17846_ & new_n20763_;
  assign new_n20765_ = ~new_n17848_ & new_n20764_;
  assign new_n20766_ = ~new_n17980_ & new_n20765_;
  assign new_n20767_ = ~new_n18011_ & new_n20766_;
  assign new_n20768_ = ~pi0647 & new_n20767_;
  assign new_n20769_ = pi0647 & new_n20705_;
  assign new_n20770_ = ~pi1157 & ~new_n20769_;
  assign new_n20771_ = ~new_n20768_ & new_n20770_;
  assign new_n20772_ = pi0630 & new_n20771_;
  assign new_n20773_ = pi0647 & ~new_n20767_;
  assign new_n20774_ = ~pi0647 & ~new_n20705_;
  assign new_n20775_ = ~new_n20773_ & ~new_n20774_;
  assign new_n20776_ = new_n17801_ & ~new_n20775_;
  assign new_n20777_ = ~new_n20772_ & ~new_n20776_;
  assign new_n20778_ = ~new_n20751_ & new_n20777_;
  assign new_n20779_ = pi0787 & ~new_n20778_;
  assign new_n20780_ = new_n17856_ & new_n20765_;
  assign new_n20781_ = ~new_n17733_ & new_n20745_;
  assign new_n20782_ = ~new_n20780_ & ~new_n20781_;
  assign new_n20783_ = pi0788 & ~new_n20782_;
  assign new_n20784_ = ~new_n16639_ & ~new_n20753_;
  assign new_n20785_ = pi0625 & new_n20784_;
  assign new_n20786_ = new_n20706_ & ~new_n20784_;
  assign new_n20787_ = ~new_n20785_ & ~new_n20786_;
  assign new_n20788_ = new_n20758_ & ~new_n20787_;
  assign new_n20789_ = ~pi0608 & ~new_n20757_;
  assign new_n20790_ = ~new_n20788_ & new_n20789_;
  assign new_n20791_ = pi1153 & new_n20706_;
  assign new_n20792_ = ~new_n20785_ & new_n20791_;
  assign new_n20793_ = pi0608 & ~new_n20759_;
  assign new_n20794_ = ~new_n20792_ & new_n20793_;
  assign new_n20795_ = ~new_n20790_ & ~new_n20794_;
  assign new_n20796_ = pi0778 & ~new_n20795_;
  assign new_n20797_ = ~pi0778 & ~new_n20786_;
  assign new_n20798_ = ~new_n20796_ & ~new_n20797_;
  assign new_n20799_ = ~pi0609 & ~new_n20798_;
  assign new_n20800_ = pi0609 & new_n20762_;
  assign new_n20801_ = ~pi1155 & ~new_n20800_;
  assign new_n20802_ = ~new_n20799_ & new_n20801_;
  assign new_n20803_ = ~pi0660 & ~new_n20710_;
  assign new_n20804_ = ~new_n20802_ & new_n20803_;
  assign new_n20805_ = pi0609 & ~new_n20798_;
  assign new_n20806_ = ~pi0609 & new_n20762_;
  assign new_n20807_ = pi1155 & ~new_n20806_;
  assign new_n20808_ = ~new_n20805_ & new_n20807_;
  assign new_n20809_ = pi0660 & ~new_n20712_;
  assign new_n20810_ = ~new_n20808_ & new_n20809_;
  assign new_n20811_ = ~new_n20804_ & ~new_n20810_;
  assign new_n20812_ = pi0785 & ~new_n20811_;
  assign new_n20813_ = ~pi0785 & ~new_n20798_;
  assign new_n20814_ = ~new_n20812_ & ~new_n20813_;
  assign new_n20815_ = ~pi0618 & ~new_n20814_;
  assign new_n20816_ = pi0618 & new_n20763_;
  assign new_n20817_ = ~pi1154 & ~new_n20816_;
  assign new_n20818_ = ~new_n20815_ & new_n20817_;
  assign new_n20819_ = ~pi0627 & ~new_n20718_;
  assign new_n20820_ = ~new_n20818_ & new_n20819_;
  assign new_n20821_ = pi0618 & ~new_n20814_;
  assign new_n20822_ = ~pi0618 & new_n20763_;
  assign new_n20823_ = pi1154 & ~new_n20822_;
  assign new_n20824_ = ~new_n20821_ & new_n20823_;
  assign new_n20825_ = pi0627 & ~new_n20720_;
  assign new_n20826_ = ~new_n20824_ & new_n20825_;
  assign new_n20827_ = ~new_n20820_ & ~new_n20826_;
  assign new_n20828_ = pi0781 & ~new_n20827_;
  assign new_n20829_ = ~pi0781 & ~new_n20814_;
  assign new_n20830_ = ~new_n20828_ & ~new_n20829_;
  assign new_n20831_ = pi0619 & ~new_n20830_;
  assign new_n20832_ = ~pi0619 & new_n20764_;
  assign new_n20833_ = pi1159 & ~new_n20832_;
  assign new_n20834_ = ~new_n20831_ & new_n20833_;
  assign new_n20835_ = pi0648 & ~new_n20732_;
  assign new_n20836_ = ~new_n20834_ & new_n20835_;
  assign new_n20837_ = ~pi0619 & ~new_n20830_;
  assign new_n20838_ = pi0619 & new_n20764_;
  assign new_n20839_ = ~pi1159 & ~new_n20838_;
  assign new_n20840_ = ~new_n20837_ & new_n20839_;
  assign new_n20841_ = ~pi0648 & ~new_n20728_;
  assign new_n20842_ = ~new_n20840_ & new_n20841_;
  assign new_n20843_ = pi0789 & ~new_n20842_;
  assign new_n20844_ = ~new_n20836_ & new_n20843_;
  assign new_n20845_ = ~pi0789 & new_n20830_;
  assign new_n20846_ = new_n17969_ & ~new_n20845_;
  assign new_n20847_ = ~new_n20844_ & new_n20846_;
  assign new_n20848_ = ~new_n20783_ & ~new_n20847_;
  assign new_n20849_ = ~new_n20364_ & ~new_n20848_;
  assign new_n20850_ = new_n18008_ & new_n20747_;
  assign new_n20851_ = pi1156 & ~new_n17982_;
  assign new_n20852_ = new_n20766_ & new_n20851_;
  assign new_n20853_ = ~new_n20850_ & ~new_n20852_;
  assign new_n20854_ = ~pi0629 & ~new_n20853_;
  assign new_n20855_ = ~pi1156 & ~new_n17991_;
  assign new_n20856_ = new_n20766_ & new_n20855_;
  assign new_n20857_ = new_n18007_ & new_n20747_;
  assign new_n20858_ = ~new_n20856_ & ~new_n20857_;
  assign new_n20859_ = pi0629 & ~new_n20858_;
  assign new_n20860_ = ~new_n20854_ & ~new_n20859_;
  assign new_n20861_ = pi0792 & ~new_n20860_;
  assign new_n20862_ = ~new_n20360_ & ~new_n20861_;
  assign new_n20863_ = ~new_n20849_ & new_n20862_;
  assign new_n20864_ = ~new_n20779_ & ~new_n20863_;
  assign new_n20865_ = pi0644 & new_n20864_;
  assign new_n20866_ = ~pi0787 & ~new_n20767_;
  assign new_n20867_ = pi1157 & ~new_n20775_;
  assign new_n20868_ = ~new_n20771_ & ~new_n20867_;
  assign new_n20869_ = pi0787 & ~new_n20868_;
  assign new_n20870_ = ~new_n20866_ & ~new_n20869_;
  assign new_n20871_ = ~pi0644 & new_n20870_;
  assign new_n20872_ = pi0715 & ~new_n20871_;
  assign new_n20873_ = ~new_n20865_ & new_n20872_;
  assign new_n20874_ = ~new_n17804_ & ~new_n20750_;
  assign new_n20875_ = new_n17804_ & new_n20705_;
  assign new_n20876_ = ~new_n20874_ & ~new_n20875_;
  assign new_n20877_ = pi0644 & ~new_n20876_;
  assign new_n20878_ = ~pi0644 & new_n20705_;
  assign new_n20879_ = ~pi0715 & ~new_n20878_;
  assign new_n20880_ = ~new_n20877_ & new_n20879_;
  assign new_n20881_ = pi1160 & ~new_n20880_;
  assign new_n20882_ = ~new_n20873_ & new_n20881_;
  assign new_n20883_ = ~pi0644 & new_n20864_;
  assign new_n20884_ = pi0644 & new_n20870_;
  assign new_n20885_ = ~pi0715 & ~new_n20884_;
  assign new_n20886_ = ~new_n20883_ & new_n20885_;
  assign new_n20887_ = ~pi0644 & ~new_n20876_;
  assign new_n20888_ = pi0644 & new_n20705_;
  assign new_n20889_ = pi0715 & ~new_n20888_;
  assign new_n20890_ = ~new_n20887_ & new_n20889_;
  assign new_n20891_ = ~pi1160 & ~new_n20890_;
  assign new_n20892_ = ~new_n20886_ & new_n20891_;
  assign new_n20893_ = ~new_n20882_ & ~new_n20892_;
  assign new_n20894_ = pi0790 & ~new_n20893_;
  assign new_n20895_ = ~pi0790 & new_n20864_;
  assign new_n20896_ = pi0832 & ~new_n20895_;
  assign new_n20897_ = ~new_n20894_ & new_n20896_;
  assign po0302 = ~new_n20704_ & ~new_n20897_;
  assign new_n20899_ = ~pi0907 & new_n6211_;
  assign new_n20900_ = pi0146 & ~new_n17320_;
  assign new_n20901_ = ~new_n20899_ & new_n20900_;
  assign new_n20902_ = pi0146 & ~new_n17313_;
  assign new_n20903_ = new_n20899_ & new_n20902_;
  assign new_n20904_ = pi0735 & pi0907;
  assign new_n20905_ = new_n17320_ & new_n20904_;
  assign new_n20906_ = ~pi0947 & ~new_n20905_;
  assign new_n20907_ = ~new_n20903_ & new_n20906_;
  assign new_n20908_ = pi0743 & new_n17320_;
  assign new_n20909_ = pi0947 & ~new_n20900_;
  assign new_n20910_ = ~new_n20908_ & new_n20909_;
  assign new_n20911_ = ~new_n20907_ & ~new_n20910_;
  assign new_n20912_ = ~new_n20901_ & ~new_n20911_;
  assign new_n20913_ = ~new_n3467_ & ~new_n20912_;
  assign new_n20914_ = pi0743 & pi0947;
  assign new_n20915_ = pi0907 & ~pi0947;
  assign new_n20916_ = pi0735 & new_n20915_;
  assign new_n20917_ = ~new_n20914_ & ~new_n20916_;
  assign new_n20918_ = new_n16636_ & ~new_n20917_;
  assign new_n20919_ = pi0146 & ~new_n16636_;
  assign new_n20920_ = ~new_n20918_ & ~new_n20919_;
  assign new_n20921_ = new_n3467_ & ~new_n20920_;
  assign new_n20922_ = ~pi0215 & ~new_n20921_;
  assign new_n20923_ = ~new_n20913_ & new_n20922_;
  assign new_n20924_ = pi0146 & new_n17343_;
  assign new_n20925_ = new_n17272_ & ~new_n20917_;
  assign new_n20926_ = pi0215 & ~new_n20925_;
  assign new_n20927_ = ~new_n20924_ & new_n20926_;
  assign new_n20928_ = ~new_n20923_ & ~new_n20927_;
  assign new_n20929_ = pi0299 & ~new_n20928_;
  assign new_n20930_ = new_n17320_ & ~new_n20917_;
  assign new_n20931_ = ~new_n6238_ & ~new_n20900_;
  assign new_n20932_ = ~new_n20930_ & new_n20931_;
  assign new_n20933_ = new_n17313_ & ~new_n20917_;
  assign new_n20934_ = new_n6238_ & ~new_n20902_;
  assign new_n20935_ = ~new_n20933_ & new_n20934_;
  assign new_n20936_ = ~new_n20932_ & ~new_n20935_;
  assign new_n20937_ = ~new_n3057_ & ~new_n20936_;
  assign new_n20938_ = new_n3057_ & new_n20920_;
  assign new_n20939_ = ~pi0223 & ~new_n20938_;
  assign new_n20940_ = ~new_n20937_ & new_n20939_;
  assign new_n20941_ = pi0146 & ~new_n17272_;
  assign new_n20942_ = ~new_n20925_ & ~new_n20941_;
  assign new_n20943_ = ~new_n6238_ & ~new_n20942_;
  assign new_n20944_ = new_n17292_ & new_n20917_;
  assign new_n20945_ = ~pi0146 & ~new_n17292_;
  assign new_n20946_ = new_n6238_ & ~new_n20945_;
  assign new_n20947_ = ~new_n20944_ & new_n20946_;
  assign new_n20948_ = ~new_n20943_ & ~new_n20947_;
  assign new_n20949_ = pi0223 & ~new_n20948_;
  assign new_n20950_ = ~pi0299 & ~new_n20949_;
  assign new_n20951_ = ~new_n20940_ & new_n20950_;
  assign new_n20952_ = ~new_n20929_ & ~new_n20951_;
  assign new_n20953_ = pi0039 & ~new_n20952_;
  assign new_n20954_ = new_n17182_ & new_n20917_;
  assign new_n20955_ = ~pi0146 & ~new_n17182_;
  assign new_n20956_ = ~pi0299 & ~new_n20955_;
  assign new_n20957_ = ~new_n20954_ & new_n20956_;
  assign new_n20958_ = new_n17193_ & new_n20917_;
  assign new_n20959_ = ~pi0146 & ~new_n17193_;
  assign new_n20960_ = pi0299 & ~new_n20959_;
  assign new_n20961_ = ~new_n20958_ & new_n20960_;
  assign new_n20962_ = ~pi0039 & ~new_n20961_;
  assign new_n20963_ = ~new_n20957_ & new_n20962_;
  assign new_n20964_ = ~pi0038 & ~new_n20963_;
  assign new_n20965_ = ~new_n20953_ & new_n20964_;
  assign new_n20966_ = ~pi0146 & ~new_n17431_;
  assign new_n20967_ = new_n2754_ & new_n20917_;
  assign new_n20968_ = new_n6257_ & new_n20967_;
  assign new_n20969_ = pi0038 & ~new_n20968_;
  assign new_n20970_ = ~new_n20966_ & new_n20969_;
  assign new_n20971_ = new_n10197_ & ~new_n20970_;
  assign new_n20972_ = ~new_n20965_ & new_n20971_;
  assign new_n20973_ = ~pi0146 & ~new_n10197_;
  assign new_n20974_ = ~pi0832 & ~new_n20973_;
  assign new_n20975_ = ~new_n20972_ & new_n20974_;
  assign new_n20976_ = ~pi0146 & ~new_n2754_;
  assign new_n20977_ = pi0832 & ~new_n20976_;
  assign new_n20978_ = ~new_n20967_ & new_n20977_;
  assign po0303 = new_n20975_ | new_n20978_;
  assign new_n20980_ = ~pi0770 & pi0947;
  assign new_n20981_ = pi0726 & new_n20915_;
  assign new_n20982_ = ~new_n20980_ & ~new_n20981_;
  assign new_n20983_ = new_n2754_ & ~new_n20982_;
  assign new_n20984_ = ~pi0147 & ~new_n2754_;
  assign new_n20985_ = pi0832 & ~new_n20984_;
  assign new_n20986_ = ~new_n20983_ & new_n20985_;
  assign new_n20987_ = ~pi0947 & new_n17260_;
  assign new_n20988_ = ~pi0039 & ~new_n20987_;
  assign new_n20989_ = ~pi0299 & new_n17326_;
  assign new_n20990_ = pi0947 & new_n20989_;
  assign new_n20991_ = ~pi0947 & new_n16865_;
  assign new_n20992_ = new_n17320_ & new_n20915_;
  assign new_n20993_ = ~new_n17331_ & ~new_n20992_;
  assign new_n20994_ = ~new_n3467_ & ~new_n20993_;
  assign new_n20995_ = ~pi0215 & ~new_n20994_;
  assign new_n20996_ = ~new_n20991_ & new_n20995_;
  assign new_n20997_ = pi0215 & ~new_n17342_;
  assign new_n20998_ = new_n17272_ & new_n20915_;
  assign new_n20999_ = new_n20997_ & ~new_n20998_;
  assign new_n21000_ = ~new_n20996_ & ~new_n20999_;
  assign new_n21001_ = pi0299 & ~new_n21000_;
  assign new_n21002_ = ~new_n17327_ & ~new_n21001_;
  assign new_n21003_ = ~new_n20990_ & new_n21002_;
  assign new_n21004_ = pi0039 & ~new_n21003_;
  assign new_n21005_ = ~new_n20988_ & ~new_n21004_;
  assign new_n21006_ = ~pi0038 & new_n21005_;
  assign new_n21007_ = pi0038 & ~pi0947;
  assign new_n21008_ = new_n17549_ & new_n21007_;
  assign new_n21009_ = ~new_n21006_ & ~new_n21008_;
  assign new_n21010_ = ~pi0770 & new_n21009_;
  assign new_n21011_ = pi0770 & ~new_n17551_;
  assign new_n21012_ = ~new_n21010_ & ~new_n21011_;
  assign new_n21013_ = ~pi0147 & ~new_n21012_;
  assign new_n21014_ = ~new_n17550_ & ~new_n21008_;
  assign new_n21015_ = pi0947 & new_n17260_;
  assign new_n21016_ = ~pi0039 & ~new_n21015_;
  assign new_n21017_ = pi0947 & new_n17326_;
  assign new_n21018_ = ~pi0299 & ~new_n21017_;
  assign new_n21019_ = pi0215 & pi0947;
  assign new_n21020_ = new_n17272_ & new_n21019_;
  assign new_n21021_ = pi0299 & ~new_n21020_;
  assign new_n21022_ = pi0947 & new_n17320_;
  assign new_n21023_ = ~new_n3467_ & ~new_n21022_;
  assign new_n21024_ = pi0947 & new_n16636_;
  assign new_n21025_ = new_n3467_ & ~new_n21024_;
  assign new_n21026_ = ~pi0215 & ~new_n21025_;
  assign new_n21027_ = ~new_n21023_ & new_n21026_;
  assign new_n21028_ = new_n21021_ & ~new_n21027_;
  assign new_n21029_ = ~new_n21018_ & ~new_n21028_;
  assign new_n21030_ = pi0039 & ~new_n21029_;
  assign new_n21031_ = ~new_n21016_ & ~new_n21030_;
  assign new_n21032_ = ~pi0038 & ~new_n21031_;
  assign new_n21033_ = new_n21014_ & ~new_n21032_;
  assign new_n21034_ = pi0147 & ~pi0770;
  assign new_n21035_ = new_n21033_ & new_n21034_;
  assign new_n21036_ = ~pi0726 & ~new_n21035_;
  assign new_n21037_ = ~new_n21013_ & new_n21036_;
  assign new_n21038_ = new_n16865_ & ~new_n20915_;
  assign new_n21039_ = ~new_n17331_ & ~new_n21022_;
  assign new_n21040_ = ~new_n3467_ & ~new_n21039_;
  assign new_n21041_ = ~pi0215 & ~new_n21040_;
  assign new_n21042_ = ~new_n21038_ & new_n21041_;
  assign new_n21043_ = ~new_n20997_ & ~new_n21042_;
  assign new_n21044_ = ~new_n21020_ & ~new_n21043_;
  assign new_n21045_ = pi0299 & ~new_n21044_;
  assign new_n21046_ = ~new_n20915_ & new_n20989_;
  assign new_n21047_ = ~new_n21045_ & ~new_n21046_;
  assign new_n21048_ = pi0039 & ~new_n21047_;
  assign new_n21049_ = new_n17260_ & ~new_n20915_;
  assign new_n21050_ = ~pi0039 & new_n21049_;
  assign new_n21051_ = ~new_n21048_ & ~new_n21050_;
  assign new_n21052_ = ~pi0147 & new_n21051_;
  assign new_n21053_ = pi0215 & ~new_n20998_;
  assign new_n21054_ = ~new_n3467_ & ~new_n20992_;
  assign new_n21055_ = pi0907 & new_n16636_;
  assign new_n21056_ = ~pi0947 & new_n21055_;
  assign new_n21057_ = new_n3467_ & ~new_n21056_;
  assign new_n21058_ = ~new_n21054_ & ~new_n21057_;
  assign new_n21059_ = ~pi0215 & ~new_n21058_;
  assign new_n21060_ = ~new_n21053_ & ~new_n21059_;
  assign new_n21061_ = pi0299 & ~new_n21060_;
  assign new_n21062_ = new_n17326_ & new_n20915_;
  assign new_n21063_ = ~pi0299 & ~new_n21062_;
  assign new_n21064_ = ~new_n21061_ & ~new_n21063_;
  assign new_n21065_ = pi0039 & ~new_n21064_;
  assign new_n21066_ = new_n17260_ & new_n20915_;
  assign new_n21067_ = ~pi0039 & ~new_n21066_;
  assign new_n21068_ = ~new_n21065_ & ~new_n21067_;
  assign new_n21069_ = pi0147 & new_n21068_;
  assign new_n21070_ = ~pi0038 & ~new_n21069_;
  assign new_n21071_ = ~new_n21052_ & new_n21070_;
  assign new_n21072_ = ~pi0147 & ~new_n17431_;
  assign new_n21073_ = new_n17431_ & new_n20915_;
  assign new_n21074_ = pi0038 & ~new_n21073_;
  assign new_n21075_ = ~new_n21072_ & new_n21074_;
  assign new_n21076_ = pi0770 & ~new_n21075_;
  assign new_n21077_ = ~new_n21071_ & new_n21076_;
  assign new_n21078_ = new_n3100_ & new_n16910_;
  assign new_n21079_ = ~new_n17323_ & ~new_n21078_;
  assign new_n21080_ = new_n6206_ & ~new_n21079_;
  assign new_n21081_ = ~pi0223 & ~new_n21080_;
  assign new_n21082_ = ~pi0947 & new_n17294_;
  assign new_n21083_ = pi0223 & ~new_n21082_;
  assign new_n21084_ = new_n17294_ & ~new_n20915_;
  assign new_n21085_ = pi0223 & ~new_n21084_;
  assign new_n21086_ = ~new_n21083_ & ~new_n21085_;
  assign new_n21087_ = ~new_n21081_ & new_n21086_;
  assign new_n21088_ = ~pi0299 & ~new_n21087_;
  assign new_n21089_ = pi0299 & pi0947;
  assign new_n21090_ = pi0299 & ~new_n21043_;
  assign new_n21091_ = ~new_n21089_ & ~new_n21090_;
  assign new_n21092_ = ~new_n21088_ & new_n21091_;
  assign new_n21093_ = pi0039 & new_n21092_;
  assign new_n21094_ = ~new_n6206_ & new_n17260_;
  assign new_n21095_ = ~pi0039 & ~new_n21094_;
  assign new_n21096_ = new_n17260_ & new_n21095_;
  assign new_n21097_ = ~new_n21093_ & ~new_n21096_;
  assign new_n21098_ = ~pi0147 & new_n21097_;
  assign new_n21099_ = ~new_n6206_ & new_n17326_;
  assign new_n21100_ = ~pi0299 & new_n21099_;
  assign new_n21101_ = ~new_n6206_ & new_n16636_;
  assign new_n21102_ = new_n3467_ & new_n21101_;
  assign new_n21103_ = ~pi0215 & ~new_n21102_;
  assign new_n21104_ = ~new_n17334_ & new_n21103_;
  assign new_n21105_ = pi0215 & ~new_n17338_;
  assign new_n21106_ = pi0299 & ~new_n21105_;
  assign new_n21107_ = ~new_n21104_ & new_n21106_;
  assign new_n21108_ = ~new_n21100_ & ~new_n21107_;
  assign new_n21109_ = pi0039 & new_n21108_;
  assign new_n21110_ = ~new_n21095_ & ~new_n21109_;
  assign new_n21111_ = pi0147 & new_n21110_;
  assign new_n21112_ = ~pi0038 & ~new_n21111_;
  assign new_n21113_ = ~new_n21098_ & new_n21112_;
  assign new_n21114_ = new_n6206_ & new_n17549_;
  assign new_n21115_ = ~pi0147 & ~new_n21114_;
  assign new_n21116_ = ~new_n6206_ & new_n17431_;
  assign new_n21117_ = pi0038 & ~new_n21116_;
  assign new_n21118_ = ~new_n21115_ & new_n21117_;
  assign new_n21119_ = ~pi0770 & ~new_n21118_;
  assign new_n21120_ = ~new_n21113_ & new_n21119_;
  assign new_n21121_ = pi0726 & ~new_n21120_;
  assign new_n21122_ = ~new_n21077_ & new_n21121_;
  assign new_n21123_ = new_n10197_ & ~new_n21122_;
  assign new_n21124_ = ~new_n21037_ & new_n21123_;
  assign new_n21125_ = ~pi0147 & ~new_n10197_;
  assign new_n21126_ = ~pi0832 & ~new_n21125_;
  assign new_n21127_ = ~new_n21124_ & new_n21126_;
  assign po0304 = ~new_n20986_ & ~new_n21127_;
  assign new_n21129_ = ~pi0148 & new_n21092_;
  assign new_n21130_ = pi0148 & new_n21108_;
  assign new_n21131_ = pi0749 & ~new_n21130_;
  assign new_n21132_ = ~new_n21129_ & new_n21131_;
  assign new_n21133_ = ~new_n9740_ & ~new_n21047_;
  assign new_n21134_ = ~new_n17327_ & ~new_n21061_;
  assign new_n21135_ = pi0148 & ~new_n21134_;
  assign new_n21136_ = ~pi0749 & ~new_n21135_;
  assign new_n21137_ = ~new_n21133_ & new_n21136_;
  assign new_n21138_ = pi0039 & ~new_n21137_;
  assign new_n21139_ = ~new_n21132_ & new_n21138_;
  assign new_n21140_ = ~pi0148 & ~new_n17260_;
  assign new_n21141_ = ~pi0039 & ~new_n21140_;
  assign new_n21142_ = ~pi0749 & pi0947;
  assign new_n21143_ = new_n21094_ & ~new_n21142_;
  assign new_n21144_ = new_n21141_ & ~new_n21143_;
  assign new_n21145_ = ~pi0038 & ~new_n21144_;
  assign new_n21146_ = ~new_n21139_ & new_n21145_;
  assign new_n21147_ = new_n21116_ & ~new_n21142_;
  assign new_n21148_ = ~pi0148 & ~new_n17431_;
  assign new_n21149_ = ~new_n21147_ & ~new_n21148_;
  assign new_n21150_ = pi0038 & ~new_n21149_;
  assign new_n21151_ = pi0706 & ~new_n21150_;
  assign new_n21152_ = ~new_n21146_ & new_n21151_;
  assign new_n21153_ = new_n3272_ & new_n6305_;
  assign new_n21154_ = ~pi0148 & ~new_n21000_;
  assign new_n21155_ = ~new_n21020_ & ~new_n21027_;
  assign new_n21156_ = pi0148 & ~new_n21155_;
  assign new_n21157_ = pi0299 & ~new_n21156_;
  assign new_n21158_ = ~new_n21154_ & new_n21157_;
  assign new_n21159_ = ~pi0148 & ~new_n17326_;
  assign new_n21160_ = new_n21018_ & ~new_n21159_;
  assign new_n21161_ = pi0749 & ~new_n21160_;
  assign new_n21162_ = ~new_n21158_ & new_n21161_;
  assign new_n21163_ = ~pi0148 & ~pi0749;
  assign new_n21164_ = ~new_n17347_ & new_n21163_;
  assign new_n21165_ = pi0039 & ~new_n21164_;
  assign new_n21166_ = ~new_n21162_ & new_n21165_;
  assign new_n21167_ = pi0749 & pi0947;
  assign new_n21168_ = new_n17260_ & new_n21167_;
  assign new_n21169_ = new_n21141_ & ~new_n21168_;
  assign new_n21170_ = ~pi0038 & ~new_n21169_;
  assign new_n21171_ = ~new_n21166_ & new_n21170_;
  assign new_n21172_ = pi0148 & ~new_n17549_;
  assign new_n21173_ = new_n17431_ & ~new_n21167_;
  assign new_n21174_ = pi0038 & ~new_n21173_;
  assign new_n21175_ = ~new_n21172_ & new_n21174_;
  assign new_n21176_ = ~pi0706 & ~new_n21175_;
  assign new_n21177_ = ~new_n21171_ & new_n21176_;
  assign new_n21178_ = new_n21153_ & ~new_n21177_;
  assign new_n21179_ = ~new_n21152_ & new_n21178_;
  assign new_n21180_ = ~pi0148 & ~new_n21153_;
  assign new_n21181_ = ~pi0057 & ~new_n21180_;
  assign new_n21182_ = ~new_n21179_ & new_n21181_;
  assign new_n21183_ = pi0057 & pi0148;
  assign new_n21184_ = ~pi0832 & ~new_n21183_;
  assign new_n21185_ = ~new_n21182_ & new_n21184_;
  assign new_n21186_ = pi0706 & new_n20915_;
  assign new_n21187_ = new_n2754_ & ~new_n21167_;
  assign new_n21188_ = ~new_n21186_ & new_n21187_;
  assign new_n21189_ = pi0148 & ~new_n2754_;
  assign new_n21190_ = pi0832 & ~new_n21189_;
  assign new_n21191_ = ~new_n21188_ & new_n21190_;
  assign po0305 = new_n21185_ | new_n21191_;
  assign new_n21193_ = ~pi0755 & pi0947;
  assign new_n21194_ = ~pi0725 & new_n20915_;
  assign new_n21195_ = ~new_n21193_ & ~new_n21194_;
  assign new_n21196_ = new_n2754_ & ~new_n21195_;
  assign new_n21197_ = ~pi0149 & ~new_n2754_;
  assign new_n21198_ = pi0832 & ~new_n21197_;
  assign new_n21199_ = ~new_n21196_ & new_n21198_;
  assign new_n21200_ = pi0149 & ~new_n17549_;
  assign new_n21201_ = new_n17431_ & ~new_n21193_;
  assign new_n21202_ = pi0038 & ~new_n21201_;
  assign new_n21203_ = ~new_n21200_ & new_n21202_;
  assign new_n21204_ = ~pi0149 & ~new_n21000_;
  assign new_n21205_ = ~new_n16145_ & ~new_n21028_;
  assign new_n21206_ = ~new_n21204_ & ~new_n21205_;
  assign new_n21207_ = ~pi0149 & ~new_n17326_;
  assign new_n21208_ = new_n21018_ & ~new_n21207_;
  assign new_n21209_ = ~pi0755 & ~new_n21208_;
  assign new_n21210_ = ~new_n21206_ & new_n21209_;
  assign new_n21211_ = ~pi0149 & pi0755;
  assign new_n21212_ = ~new_n17347_ & new_n21211_;
  assign new_n21213_ = pi0039 & ~new_n21212_;
  assign new_n21214_ = ~new_n21210_ & new_n21213_;
  assign new_n21215_ = new_n17260_ & new_n21193_;
  assign new_n21216_ = ~pi0149 & ~new_n17260_;
  assign new_n21217_ = ~pi0039 & ~new_n21216_;
  assign new_n21218_ = ~new_n21215_ & new_n21217_;
  assign new_n21219_ = ~pi0038 & ~new_n21218_;
  assign new_n21220_ = ~new_n21214_ & new_n21219_;
  assign new_n21221_ = ~new_n21203_ & ~new_n21220_;
  assign new_n21222_ = pi0725 & ~new_n21221_;
  assign new_n21223_ = ~new_n21066_ & new_n21218_;
  assign new_n21224_ = ~pi0149 & new_n21092_;
  assign new_n21225_ = pi0149 & new_n21108_;
  assign new_n21226_ = ~pi0755 & ~new_n21225_;
  assign new_n21227_ = ~new_n21224_ & new_n21226_;
  assign new_n21228_ = ~pi0149 & new_n21045_;
  assign new_n21229_ = pi0149 & ~new_n21134_;
  assign new_n21230_ = pi0755 & ~new_n21046_;
  assign new_n21231_ = ~new_n21229_ & new_n21230_;
  assign new_n21232_ = ~new_n21228_ & new_n21231_;
  assign new_n21233_ = pi0039 & ~new_n21232_;
  assign new_n21234_ = ~new_n21227_ & new_n21233_;
  assign new_n21235_ = ~new_n21223_ & ~new_n21234_;
  assign new_n21236_ = ~pi0038 & ~new_n21235_;
  assign new_n21237_ = ~new_n6206_ & new_n16647_;
  assign new_n21238_ = pi0755 & pi0947;
  assign new_n21239_ = ~pi0039 & ~new_n21238_;
  assign new_n21240_ = new_n21237_ & new_n21239_;
  assign new_n21241_ = ~pi0149 & ~new_n17431_;
  assign new_n21242_ = pi0038 & ~new_n21241_;
  assign new_n21243_ = ~new_n21240_ & new_n21242_;
  assign new_n21244_ = ~pi0725 & ~new_n21243_;
  assign new_n21245_ = ~new_n21236_ & new_n21244_;
  assign new_n21246_ = ~new_n21222_ & ~new_n21245_;
  assign new_n21247_ = new_n10197_ & ~new_n21246_;
  assign new_n21248_ = ~pi0149 & ~new_n10197_;
  assign new_n21249_ = ~pi0832 & ~new_n21248_;
  assign new_n21250_ = ~new_n21247_ & new_n21249_;
  assign po0306 = ~new_n21199_ & ~new_n21250_;
  assign new_n21252_ = ~pi0150 & new_n21003_;
  assign new_n21253_ = pi0150 & ~new_n21029_;
  assign new_n21254_ = ~pi0751 & ~new_n21253_;
  assign new_n21255_ = ~new_n21252_ & new_n21254_;
  assign new_n21256_ = ~pi0150 & pi0751;
  assign new_n21257_ = ~new_n17347_ & new_n21256_;
  assign new_n21258_ = ~new_n21255_ & ~new_n21257_;
  assign new_n21259_ = pi0039 & ~new_n21258_;
  assign new_n21260_ = pi0150 & ~new_n17260_;
  assign new_n21261_ = pi0751 & new_n17260_;
  assign new_n21262_ = ~new_n21260_ & ~new_n21261_;
  assign new_n21263_ = new_n20988_ & new_n21262_;
  assign new_n21264_ = ~pi0038 & ~new_n21263_;
  assign new_n21265_ = ~new_n21259_ & new_n21264_;
  assign new_n21266_ = pi0150 & ~new_n17549_;
  assign new_n21267_ = ~pi0751 & pi0947;
  assign new_n21268_ = new_n17431_ & ~new_n21267_;
  assign new_n21269_ = ~new_n21266_ & ~new_n21268_;
  assign new_n21270_ = pi0038 & ~new_n21269_;
  assign new_n21271_ = pi0701 & ~new_n21270_;
  assign new_n21272_ = ~new_n21265_ & new_n21271_;
  assign new_n21273_ = ~pi0150 & ~new_n21047_;
  assign new_n21274_ = pi0150 & ~new_n21064_;
  assign new_n21275_ = pi0751 & ~new_n21274_;
  assign new_n21276_ = ~new_n21273_ & new_n21275_;
  assign new_n21277_ = ~pi0150 & new_n21092_;
  assign new_n21278_ = pi0150 & new_n21108_;
  assign new_n21279_ = ~pi0751 & ~new_n21278_;
  assign new_n21280_ = ~new_n21277_ & new_n21279_;
  assign new_n21281_ = ~new_n21276_ & ~new_n21280_;
  assign new_n21282_ = pi0039 & ~new_n21281_;
  assign new_n21283_ = new_n21049_ & ~new_n21267_;
  assign new_n21284_ = ~pi0039 & ~new_n21260_;
  assign new_n21285_ = ~new_n21283_ & new_n21284_;
  assign new_n21286_ = ~pi0038 & ~new_n21285_;
  assign new_n21287_ = ~new_n21282_ & new_n21286_;
  assign new_n21288_ = pi0751 & pi0947;
  assign new_n21289_ = ~pi0039 & ~new_n21288_;
  assign new_n21290_ = new_n21237_ & new_n21289_;
  assign new_n21291_ = ~pi0150 & ~new_n17431_;
  assign new_n21292_ = pi0038 & ~new_n21291_;
  assign new_n21293_ = ~new_n21290_ & new_n21292_;
  assign new_n21294_ = ~pi0701 & ~new_n21293_;
  assign new_n21295_ = ~new_n21287_ & new_n21294_;
  assign new_n21296_ = ~new_n21272_ & ~new_n21295_;
  assign new_n21297_ = new_n10197_ & ~new_n21296_;
  assign new_n21298_ = ~pi0150 & ~new_n10197_;
  assign new_n21299_ = ~pi0832 & ~new_n21298_;
  assign new_n21300_ = ~new_n21297_ & new_n21299_;
  assign new_n21301_ = ~pi0701 & new_n20915_;
  assign new_n21302_ = ~new_n21267_ & ~new_n21301_;
  assign new_n21303_ = new_n2754_ & ~new_n21302_;
  assign new_n21304_ = ~pi0150 & ~new_n2754_;
  assign new_n21305_ = pi0832 & ~new_n21304_;
  assign new_n21306_ = ~new_n21303_ & new_n21305_;
  assign po0307 = ~new_n21300_ & ~new_n21306_;
  assign new_n21308_ = ~pi0745 & pi0947;
  assign new_n21309_ = ~pi0723 & new_n20915_;
  assign new_n21310_ = ~new_n21308_ & ~new_n21309_;
  assign new_n21311_ = new_n2754_ & ~new_n21310_;
  assign new_n21312_ = ~pi0151 & ~new_n2754_;
  assign new_n21313_ = pi0832 & ~new_n21312_;
  assign new_n21314_ = ~new_n21311_ & new_n21313_;
  assign new_n21315_ = ~pi0151 & ~new_n17260_;
  assign new_n21316_ = ~pi0745 & new_n21015_;
  assign new_n21317_ = ~new_n21315_ & ~new_n21316_;
  assign new_n21318_ = new_n21067_ & new_n21317_;
  assign new_n21319_ = ~new_n17342_ & ~new_n20998_;
  assign new_n21320_ = ~pi0151 & new_n21319_;
  assign new_n21321_ = ~new_n17338_ & ~new_n21320_;
  assign new_n21322_ = pi0215 & ~new_n21321_;
  assign new_n21323_ = pi0151 & ~new_n3467_;
  assign new_n21324_ = ~new_n17333_ & new_n21323_;
  assign new_n21325_ = ~new_n17332_ & ~new_n21324_;
  assign new_n21326_ = ~pi0151 & ~new_n16636_;
  assign new_n21327_ = new_n21057_ & ~new_n21326_;
  assign new_n21328_ = ~new_n21101_ & new_n21327_;
  assign new_n21329_ = ~pi0215 & ~new_n21328_;
  assign new_n21330_ = new_n21325_ & new_n21329_;
  assign new_n21331_ = ~new_n21322_ & ~new_n21330_;
  assign new_n21332_ = pi0299 & ~new_n21331_;
  assign new_n21333_ = pi0151 & ~new_n21099_;
  assign new_n21334_ = new_n21088_ & ~new_n21333_;
  assign new_n21335_ = ~new_n21332_ & ~new_n21334_;
  assign new_n21336_ = ~pi0745 & ~new_n21335_;
  assign new_n21337_ = new_n21325_ & ~new_n21327_;
  assign new_n21338_ = new_n21041_ & new_n21337_;
  assign new_n21339_ = ~new_n21322_ & ~new_n21338_;
  assign new_n21340_ = ~new_n21020_ & ~new_n21339_;
  assign new_n21341_ = pi0299 & ~new_n21340_;
  assign new_n21342_ = ~pi0151 & ~new_n17326_;
  assign new_n21343_ = new_n21063_ & ~new_n21342_;
  assign new_n21344_ = pi0745 & ~new_n21343_;
  assign new_n21345_ = ~new_n21341_ & new_n21344_;
  assign new_n21346_ = pi0039 & ~new_n21345_;
  assign new_n21347_ = ~new_n21336_ & new_n21346_;
  assign new_n21348_ = ~new_n21318_ & ~new_n21347_;
  assign new_n21349_ = ~pi0038 & ~new_n21348_;
  assign new_n21350_ = pi0745 & pi0947;
  assign new_n21351_ = ~pi0039 & ~new_n21350_;
  assign new_n21352_ = new_n21237_ & new_n21351_;
  assign new_n21353_ = ~pi0151 & ~new_n17431_;
  assign new_n21354_ = pi0038 & ~new_n21353_;
  assign new_n21355_ = ~new_n21352_ & new_n21354_;
  assign new_n21356_ = ~pi0723 & ~new_n21355_;
  assign new_n21357_ = ~new_n21349_ & new_n21356_;
  assign new_n21358_ = ~pi0745 & ~new_n17327_;
  assign new_n21359_ = ~pi0151 & ~new_n17347_;
  assign new_n21360_ = ~new_n21358_ & new_n21359_;
  assign new_n21361_ = new_n21025_ & ~new_n21326_;
  assign new_n21362_ = new_n21325_ & ~new_n21361_;
  assign new_n21363_ = new_n20995_ & new_n21362_;
  assign new_n21364_ = new_n21053_ & ~new_n21321_;
  assign new_n21365_ = pi0299 & ~new_n21364_;
  assign new_n21366_ = ~new_n21363_ & new_n21365_;
  assign new_n21367_ = ~pi0745 & ~new_n21018_;
  assign new_n21368_ = ~new_n21366_ & new_n21367_;
  assign new_n21369_ = ~new_n21360_ & ~new_n21368_;
  assign new_n21370_ = pi0039 & ~new_n21369_;
  assign new_n21371_ = ~pi0039 & ~new_n21317_;
  assign new_n21372_ = ~pi0038 & ~new_n21371_;
  assign new_n21373_ = ~new_n21370_ & new_n21372_;
  assign new_n21374_ = pi0151 & ~new_n17549_;
  assign new_n21375_ = new_n17431_ & ~new_n21308_;
  assign new_n21376_ = ~new_n21374_ & ~new_n21375_;
  assign new_n21377_ = pi0038 & ~new_n21376_;
  assign new_n21378_ = pi0723 & ~new_n21377_;
  assign new_n21379_ = ~new_n21373_ & new_n21378_;
  assign new_n21380_ = ~new_n21357_ & ~new_n21379_;
  assign new_n21381_ = new_n10197_ & ~new_n21380_;
  assign new_n21382_ = ~pi0151 & ~new_n10197_;
  assign new_n21383_ = ~pi0832 & ~new_n21382_;
  assign new_n21384_ = ~new_n21381_ & new_n21383_;
  assign po0308 = ~new_n21314_ & ~new_n21384_;
  assign new_n21386_ = ~pi0152 & ~new_n17322_;
  assign new_n21387_ = ~pi0947 & new_n17322_;
  assign new_n21388_ = ~new_n3057_ & ~new_n21387_;
  assign new_n21389_ = ~new_n21386_ & new_n21388_;
  assign new_n21390_ = ~new_n6206_ & new_n17322_;
  assign new_n21391_ = ~new_n3057_ & ~new_n21390_;
  assign new_n21392_ = ~new_n21389_ & new_n21391_;
  assign new_n21393_ = pi0152 & ~new_n16636_;
  assign new_n21394_ = ~new_n21101_ & ~new_n21393_;
  assign new_n21395_ = new_n3057_ & new_n21394_;
  assign new_n21396_ = ~pi0223 & ~new_n21395_;
  assign new_n21397_ = ~new_n21392_ & new_n21396_;
  assign new_n21398_ = ~pi0152 & ~new_n17294_;
  assign new_n21399_ = new_n21085_ & ~new_n21398_;
  assign new_n21400_ = new_n21083_ & ~new_n21398_;
  assign new_n21401_ = ~pi0299 & ~new_n21400_;
  assign new_n21402_ = ~new_n21399_ & new_n21401_;
  assign new_n21403_ = ~new_n21397_ & new_n21402_;
  assign new_n21404_ = new_n3467_ & new_n21394_;
  assign new_n21405_ = ~pi0215 & ~new_n21404_;
  assign new_n21406_ = pi0152 & new_n21039_;
  assign new_n21407_ = new_n21054_ & ~new_n21406_;
  assign new_n21408_ = ~new_n17333_ & new_n21407_;
  assign new_n21409_ = new_n21405_ & ~new_n21408_;
  assign new_n21410_ = ~pi0152 & ~new_n17338_;
  assign new_n21411_ = new_n20997_ & ~new_n21410_;
  assign new_n21412_ = pi0299 & ~new_n21411_;
  assign new_n21413_ = ~new_n21409_ & new_n21412_;
  assign new_n21414_ = pi0759 & ~new_n21413_;
  assign new_n21415_ = ~new_n21403_ & new_n21414_;
  assign new_n21416_ = ~new_n21056_ & ~new_n21393_;
  assign new_n21417_ = new_n3057_ & ~new_n21416_;
  assign new_n21418_ = new_n17322_ & ~new_n20915_;
  assign new_n21419_ = ~new_n3057_ & ~new_n21418_;
  assign new_n21420_ = ~new_n21386_ & new_n21419_;
  assign new_n21421_ = ~new_n21417_ & ~new_n21420_;
  assign new_n21422_ = ~pi0223 & ~new_n21421_;
  assign new_n21423_ = ~pi0299 & ~new_n21399_;
  assign new_n21424_ = ~new_n21422_ & new_n21423_;
  assign new_n21425_ = ~new_n21038_ & new_n21405_;
  assign new_n21426_ = ~new_n21407_ & new_n21425_;
  assign new_n21427_ = ~new_n20915_ & ~new_n21105_;
  assign new_n21428_ = new_n21411_ & ~new_n21427_;
  assign new_n21429_ = pi0299 & ~new_n21428_;
  assign new_n21430_ = ~new_n21426_ & new_n21429_;
  assign new_n21431_ = ~pi0759 & ~new_n21430_;
  assign new_n21432_ = ~new_n21424_ & new_n21431_;
  assign new_n21433_ = pi0039 & ~new_n21432_;
  assign new_n21434_ = ~new_n21415_ & new_n21433_;
  assign new_n21435_ = pi0152 & ~new_n17260_;
  assign new_n21436_ = pi0759 & pi0947;
  assign new_n21437_ = ~pi0039 & ~new_n21436_;
  assign new_n21438_ = ~new_n17261_ & ~new_n21437_;
  assign new_n21439_ = ~new_n21435_ & ~new_n21438_;
  assign new_n21440_ = ~new_n21066_ & new_n21439_;
  assign new_n21441_ = ~pi0038 & ~new_n21440_;
  assign new_n21442_ = ~new_n21434_ & new_n21441_;
  assign new_n21443_ = new_n16647_ & ~new_n20915_;
  assign new_n21444_ = new_n21437_ & new_n21443_;
  assign new_n21445_ = ~pi0152 & ~new_n17431_;
  assign new_n21446_ = pi0038 & ~new_n21445_;
  assign new_n21447_ = ~new_n21444_ & new_n21446_;
  assign new_n21448_ = pi0696 & ~new_n21447_;
  assign new_n21449_ = ~new_n21442_ & new_n21448_;
  assign new_n21450_ = ~new_n20994_ & ~new_n21407_;
  assign new_n21451_ = ~new_n21022_ & ~new_n21450_;
  assign new_n21452_ = ~new_n21024_ & ~new_n21393_;
  assign new_n21453_ = new_n3467_ & new_n21452_;
  assign new_n21454_ = ~pi0215 & ~new_n21453_;
  assign new_n21455_ = ~new_n21451_ & new_n21454_;
  assign new_n21456_ = pi0152 & new_n20999_;
  assign new_n21457_ = new_n21021_ & ~new_n21456_;
  assign new_n21458_ = ~new_n21455_ & new_n21457_;
  assign new_n21459_ = new_n3057_ & ~new_n21452_;
  assign new_n21460_ = ~new_n21389_ & ~new_n21459_;
  assign new_n21461_ = ~pi0223 & ~new_n21460_;
  assign new_n21462_ = new_n21401_ & ~new_n21461_;
  assign new_n21463_ = pi0759 & ~new_n21462_;
  assign new_n21464_ = ~new_n21458_ & new_n21463_;
  assign new_n21465_ = ~pi0759 & ~new_n17347_;
  assign new_n21466_ = pi0152 & new_n21465_;
  assign new_n21467_ = pi0039 & ~new_n21466_;
  assign new_n21468_ = ~new_n21464_ & new_n21467_;
  assign new_n21469_ = ~pi0038 & ~new_n21439_;
  assign new_n21470_ = ~new_n21468_ & new_n21469_;
  assign new_n21471_ = ~pi0152 & ~new_n17549_;
  assign new_n21472_ = new_n17431_ & ~new_n21436_;
  assign new_n21473_ = pi0038 & ~new_n21472_;
  assign new_n21474_ = ~new_n21471_ & new_n21473_;
  assign new_n21475_ = ~pi0696 & ~new_n21474_;
  assign new_n21476_ = ~new_n21470_ & new_n21475_;
  assign new_n21477_ = ~new_n21449_ & ~new_n21476_;
  assign new_n21478_ = new_n10197_ & ~new_n21477_;
  assign new_n21479_ = ~pi0152 & ~new_n10197_;
  assign new_n21480_ = ~pi0832 & ~new_n21479_;
  assign new_n21481_ = ~new_n21478_ & new_n21480_;
  assign new_n21482_ = pi0696 & new_n20915_;
  assign new_n21483_ = new_n2754_ & ~new_n21436_;
  assign new_n21484_ = ~new_n21482_ & new_n21483_;
  assign new_n21485_ = ~pi0152 & ~new_n2754_;
  assign new_n21486_ = pi0832 & ~new_n21485_;
  assign new_n21487_ = ~new_n21484_ & new_n21486_;
  assign po0309 = new_n21481_ | new_n21487_;
  assign new_n21489_ = pi0766 & pi0947;
  assign new_n21490_ = new_n2754_ & ~new_n21489_;
  assign new_n21491_ = pi0700 & new_n20915_;
  assign new_n21492_ = new_n21490_ & ~new_n21491_;
  assign new_n21493_ = pi0153 & ~new_n2754_;
  assign new_n21494_ = pi0832 & ~new_n21493_;
  assign new_n21495_ = ~new_n21492_ & new_n21494_;
  assign new_n21496_ = ~pi0153 & ~new_n17260_;
  assign new_n21497_ = ~pi0766 & new_n18106_;
  assign new_n21498_ = ~new_n21016_ & ~new_n21497_;
  assign new_n21499_ = ~new_n21496_ & ~new_n21498_;
  assign new_n21500_ = ~new_n21066_ & new_n21499_;
  assign new_n21501_ = pi0153 & ~new_n17338_;
  assign new_n21502_ = new_n20997_ & ~new_n21501_;
  assign new_n21503_ = pi0153 & ~new_n3467_;
  assign new_n21504_ = ~new_n17333_ & new_n21503_;
  assign new_n21505_ = ~new_n17332_ & ~new_n21504_;
  assign new_n21506_ = ~pi0153 & ~new_n16636_;
  assign new_n21507_ = new_n21025_ & ~new_n21506_;
  assign new_n21508_ = ~new_n21055_ & new_n21507_;
  assign new_n21509_ = ~pi0215 & ~new_n21508_;
  assign new_n21510_ = new_n21505_ & new_n21509_;
  assign new_n21511_ = ~new_n21502_ & ~new_n21510_;
  assign new_n21512_ = pi0299 & ~new_n21511_;
  assign new_n21513_ = pi0153 & ~new_n21099_;
  assign new_n21514_ = new_n21088_ & ~new_n21513_;
  assign new_n21515_ = ~new_n21512_ & ~new_n21514_;
  assign new_n21516_ = pi0766 & ~new_n21515_;
  assign new_n21517_ = new_n21057_ & ~new_n21506_;
  assign new_n21518_ = ~new_n21040_ & ~new_n21517_;
  assign new_n21519_ = new_n21505_ & new_n21518_;
  assign new_n21520_ = ~pi0215 & ~new_n21519_;
  assign new_n21521_ = new_n21105_ & ~new_n21502_;
  assign new_n21522_ = ~new_n21020_ & ~new_n21521_;
  assign new_n21523_ = ~new_n21520_ & new_n21522_;
  assign new_n21524_ = pi0299 & ~new_n21523_;
  assign new_n21525_ = ~pi0153 & ~new_n17326_;
  assign new_n21526_ = new_n21063_ & ~new_n21525_;
  assign new_n21527_ = ~pi0766 & ~new_n21526_;
  assign new_n21528_ = ~new_n21524_ & new_n21527_;
  assign new_n21529_ = pi0039 & ~new_n21528_;
  assign new_n21530_ = ~new_n21516_ & new_n21529_;
  assign new_n21531_ = ~new_n21500_ & ~new_n21530_;
  assign new_n21532_ = ~pi0038 & ~new_n21531_;
  assign new_n21533_ = ~pi0766 & pi0947;
  assign new_n21534_ = ~pi0039 & ~new_n21533_;
  assign new_n21535_ = new_n21237_ & new_n21534_;
  assign new_n21536_ = ~pi0153 & ~new_n17431_;
  assign new_n21537_ = pi0038 & ~new_n21536_;
  assign new_n21538_ = ~new_n21535_ & new_n21537_;
  assign new_n21539_ = ~new_n21532_ & ~new_n21538_;
  assign new_n21540_ = pi0700 & ~new_n21539_;
  assign new_n21541_ = new_n21018_ & ~new_n21525_;
  assign new_n21542_ = new_n21505_ & ~new_n21507_;
  assign new_n21543_ = new_n20995_ & new_n21542_;
  assign new_n21544_ = new_n20999_ & ~new_n21501_;
  assign new_n21545_ = pi0299 & ~new_n21544_;
  assign new_n21546_ = ~new_n21543_ & new_n21545_;
  assign new_n21547_ = pi0766 & ~new_n21546_;
  assign new_n21548_ = ~new_n21541_ & new_n21547_;
  assign new_n21549_ = ~pi0153 & ~pi0766;
  assign new_n21550_ = ~new_n17347_ & new_n21549_;
  assign new_n21551_ = pi0039 & ~new_n21550_;
  assign new_n21552_ = ~new_n21548_ & new_n21551_;
  assign new_n21553_ = ~pi0038 & ~new_n21499_;
  assign new_n21554_ = ~new_n21552_ & new_n21553_;
  assign new_n21555_ = pi0153 & ~new_n17549_;
  assign new_n21556_ = new_n6257_ & new_n21490_;
  assign new_n21557_ = pi0038 & ~new_n21556_;
  assign new_n21558_ = ~new_n21555_ & new_n21557_;
  assign new_n21559_ = ~pi0700 & ~new_n21558_;
  assign new_n21560_ = ~new_n21554_ & new_n21559_;
  assign new_n21561_ = new_n21153_ & ~new_n21560_;
  assign new_n21562_ = ~new_n21540_ & new_n21561_;
  assign new_n21563_ = ~pi0153 & ~new_n21153_;
  assign new_n21564_ = ~pi0057 & ~new_n21563_;
  assign new_n21565_ = ~new_n21562_ & new_n21564_;
  assign new_n21566_ = pi0057 & pi0153;
  assign new_n21567_ = ~pi0832 & ~new_n21566_;
  assign new_n21568_ = ~new_n21565_ & new_n21567_;
  assign po0310 = new_n21495_ | new_n21568_;
  assign new_n21570_ = ~pi0742 & pi0947;
  assign new_n21571_ = ~pi0704 & new_n20915_;
  assign new_n21572_ = ~new_n21570_ & ~new_n21571_;
  assign new_n21573_ = new_n2754_ & ~new_n21572_;
  assign new_n21574_ = ~pi0154 & ~new_n2754_;
  assign new_n21575_ = pi0832 & ~new_n21574_;
  assign new_n21576_ = ~new_n21573_ & new_n21575_;
  assign new_n21577_ = ~pi0154 & ~new_n17260_;
  assign new_n21578_ = new_n21067_ & ~new_n21577_;
  assign new_n21579_ = ~new_n21094_ & new_n21578_;
  assign new_n21580_ = ~pi0154 & ~new_n21092_;
  assign new_n21581_ = pi0154 & ~new_n21108_;
  assign new_n21582_ = pi0039 & ~new_n21581_;
  assign new_n21583_ = ~new_n21580_ & new_n21582_;
  assign new_n21584_ = ~new_n21579_ & ~new_n21583_;
  assign new_n21585_ = ~pi0038 & ~new_n21584_;
  assign new_n21586_ = ~pi0154 & ~new_n17431_;
  assign new_n21587_ = new_n21117_ & ~new_n21586_;
  assign new_n21588_ = ~pi0742 & ~new_n21587_;
  assign new_n21589_ = ~new_n21585_ & new_n21588_;
  assign new_n21590_ = ~pi0154 & new_n21047_;
  assign new_n21591_ = pi0154 & new_n21064_;
  assign new_n21592_ = pi0039 & ~new_n21591_;
  assign new_n21593_ = ~new_n21590_ & new_n21592_;
  assign new_n21594_ = ~new_n21578_ & ~new_n21593_;
  assign new_n21595_ = ~pi0038 & ~new_n21594_;
  assign new_n21596_ = new_n21074_ & ~new_n21586_;
  assign new_n21597_ = pi0742 & ~new_n21596_;
  assign new_n21598_ = ~new_n21595_ & new_n21597_;
  assign new_n21599_ = ~pi0704 & ~new_n21598_;
  assign new_n21600_ = ~new_n21589_ & new_n21599_;
  assign new_n21601_ = new_n21016_ & ~new_n21577_;
  assign new_n21602_ = ~pi0154 & ~new_n21003_;
  assign new_n21603_ = pi0154 & new_n21029_;
  assign new_n21604_ = pi0039 & ~new_n21603_;
  assign new_n21605_ = ~new_n21602_ & new_n21604_;
  assign new_n21606_ = ~new_n21601_ & ~new_n21605_;
  assign new_n21607_ = ~pi0038 & ~new_n21606_;
  assign new_n21608_ = ~pi0154 & ~new_n17549_;
  assign new_n21609_ = ~new_n21014_ & ~new_n21608_;
  assign new_n21610_ = ~pi0742 & ~new_n21609_;
  assign new_n21611_ = ~new_n21607_ & new_n21610_;
  assign new_n21612_ = ~pi0154 & pi0742;
  assign new_n21613_ = ~new_n17551_ & new_n21612_;
  assign new_n21614_ = pi0704 & ~new_n21613_;
  assign new_n21615_ = ~new_n21611_ & new_n21614_;
  assign new_n21616_ = new_n10197_ & ~new_n21615_;
  assign new_n21617_ = ~new_n21600_ & new_n21616_;
  assign new_n21618_ = ~pi0154 & ~new_n10197_;
  assign new_n21619_ = ~pi0832 & ~new_n21618_;
  assign new_n21620_ = ~new_n21617_ & new_n21619_;
  assign po0311 = ~new_n21576_ & ~new_n21620_;
  assign new_n21622_ = ~pi0038 & ~new_n21068_;
  assign new_n21623_ = ~new_n21074_ & ~new_n21622_;
  assign new_n21624_ = pi0757 & new_n21623_;
  assign new_n21625_ = ~pi0038 & ~new_n21110_;
  assign new_n21626_ = ~new_n21117_ & ~new_n21625_;
  assign new_n21627_ = ~pi0757 & new_n21626_;
  assign new_n21628_ = ~pi0686 & ~new_n21627_;
  assign new_n21629_ = ~new_n21624_ & new_n21628_;
  assign new_n21630_ = ~pi0757 & new_n21033_;
  assign new_n21631_ = pi0686 & ~new_n21630_;
  assign new_n21632_ = new_n10197_ & ~new_n21631_;
  assign new_n21633_ = ~new_n21629_ & new_n21632_;
  assign new_n21634_ = pi0155 & ~new_n21633_;
  assign new_n21635_ = ~pi0038 & ~new_n21051_;
  assign new_n21636_ = new_n17431_ & new_n21074_;
  assign new_n21637_ = ~new_n21635_ & ~new_n21636_;
  assign new_n21638_ = pi0757 & new_n21637_;
  assign new_n21639_ = ~pi0038 & ~new_n21097_;
  assign new_n21640_ = pi0038 & new_n21114_;
  assign new_n21641_ = ~new_n21639_ & ~new_n21640_;
  assign new_n21642_ = ~pi0757 & new_n21641_;
  assign new_n21643_ = ~pi0686 & ~new_n21642_;
  assign new_n21644_ = ~new_n21638_ & new_n21643_;
  assign new_n21645_ = ~pi0757 & new_n21009_;
  assign new_n21646_ = pi0757 & ~new_n17551_;
  assign new_n21647_ = pi0686 & ~new_n21646_;
  assign new_n21648_ = ~new_n21645_ & new_n21647_;
  assign new_n21649_ = ~new_n21644_ & ~new_n21648_;
  assign new_n21650_ = ~pi0155 & new_n10197_;
  assign new_n21651_ = ~new_n21649_ & new_n21650_;
  assign new_n21652_ = ~new_n21634_ & ~new_n21651_;
  assign new_n21653_ = ~pi0832 & ~new_n21652_;
  assign new_n21654_ = ~pi0757 & pi0947;
  assign new_n21655_ = ~pi0686 & new_n20915_;
  assign new_n21656_ = ~new_n21654_ & ~new_n21655_;
  assign new_n21657_ = new_n2754_ & ~new_n21656_;
  assign new_n21658_ = ~pi0155 & ~new_n2754_;
  assign new_n21659_ = pi0832 & ~new_n21658_;
  assign new_n21660_ = ~new_n21657_ & new_n21659_;
  assign po0312 = ~new_n21653_ & ~new_n21660_;
  assign new_n21662_ = ~pi0741 & pi0947;
  assign new_n21663_ = ~pi0724 & new_n20915_;
  assign new_n21664_ = ~new_n21662_ & ~new_n21663_;
  assign new_n21665_ = new_n2754_ & ~new_n21664_;
  assign new_n21666_ = ~pi0156 & ~new_n2754_;
  assign new_n21667_ = pi0832 & ~new_n21666_;
  assign new_n21668_ = ~new_n21665_ & new_n21667_;
  assign new_n21669_ = pi0741 & ~new_n21637_;
  assign new_n21670_ = ~pi0741 & ~new_n21641_;
  assign new_n21671_ = ~pi0724 & ~new_n21670_;
  assign new_n21672_ = ~new_n21669_ & new_n21671_;
  assign new_n21673_ = ~pi0741 & ~new_n21009_;
  assign new_n21674_ = pi0741 & new_n17551_;
  assign new_n21675_ = pi0724 & ~new_n21674_;
  assign new_n21676_ = ~new_n21673_ & new_n21675_;
  assign new_n21677_ = new_n10197_ & ~new_n21676_;
  assign new_n21678_ = ~new_n21672_ & new_n21677_;
  assign new_n21679_ = ~pi0156 & ~new_n21678_;
  assign new_n21680_ = pi0741 & ~new_n21623_;
  assign new_n21681_ = ~pi0741 & ~new_n21626_;
  assign new_n21682_ = ~pi0724 & ~new_n21681_;
  assign new_n21683_ = ~new_n21680_ & new_n21682_;
  assign new_n21684_ = pi0724 & ~pi0741;
  assign new_n21685_ = new_n21033_ & new_n21684_;
  assign new_n21686_ = ~new_n21683_ & ~new_n21685_;
  assign new_n21687_ = pi0156 & new_n10197_;
  assign new_n21688_ = ~new_n21686_ & new_n21687_;
  assign new_n21689_ = ~pi0832 & ~new_n21688_;
  assign new_n21690_ = ~new_n21679_ & new_n21689_;
  assign po0313 = ~new_n21668_ & ~new_n21690_;
  assign new_n21692_ = ~pi0760 & pi0947;
  assign new_n21693_ = ~pi0688 & new_n20915_;
  assign new_n21694_ = ~new_n21692_ & ~new_n21693_;
  assign new_n21695_ = new_n2754_ & ~new_n21694_;
  assign new_n21696_ = ~pi0157 & ~new_n2754_;
  assign new_n21697_ = pi0832 & ~new_n21696_;
  assign new_n21698_ = ~new_n21695_ & new_n21697_;
  assign new_n21699_ = pi0157 & ~new_n17549_;
  assign new_n21700_ = new_n17431_ & ~new_n21692_;
  assign new_n21701_ = pi0038 & ~new_n21700_;
  assign new_n21702_ = ~new_n21699_ & new_n21701_;
  assign new_n21703_ = ~pi0157 & ~new_n21000_;
  assign new_n21704_ = ~new_n13815_ & ~new_n21028_;
  assign new_n21705_ = ~new_n21703_ & ~new_n21704_;
  assign new_n21706_ = ~pi0157 & ~new_n17326_;
  assign new_n21707_ = new_n21018_ & ~new_n21706_;
  assign new_n21708_ = ~pi0760 & ~new_n21707_;
  assign new_n21709_ = ~new_n21705_ & new_n21708_;
  assign new_n21710_ = ~pi0157 & pi0760;
  assign new_n21711_ = ~new_n17347_ & new_n21710_;
  assign new_n21712_ = pi0039 & ~new_n21711_;
  assign new_n21713_ = ~new_n21709_ & new_n21712_;
  assign new_n21714_ = new_n17260_ & new_n21692_;
  assign new_n21715_ = ~pi0157 & ~new_n17260_;
  assign new_n21716_ = ~pi0039 & ~new_n21715_;
  assign new_n21717_ = ~new_n21714_ & new_n21716_;
  assign new_n21718_ = ~pi0038 & ~new_n21717_;
  assign new_n21719_ = ~new_n21713_ & new_n21718_;
  assign new_n21720_ = ~new_n21702_ & ~new_n21719_;
  assign new_n21721_ = pi0688 & ~new_n21720_;
  assign new_n21722_ = ~new_n21066_ & new_n21717_;
  assign new_n21723_ = ~pi0760 & new_n21092_;
  assign new_n21724_ = pi0760 & ~new_n21047_;
  assign new_n21725_ = ~pi0157 & ~new_n21724_;
  assign new_n21726_ = ~new_n21723_ & new_n21725_;
  assign new_n21727_ = pi0760 & ~new_n21064_;
  assign new_n21728_ = ~pi0760 & new_n21108_;
  assign new_n21729_ = pi0157 & ~new_n21728_;
  assign new_n21730_ = ~new_n21727_ & new_n21729_;
  assign new_n21731_ = pi0039 & ~new_n21730_;
  assign new_n21732_ = ~new_n21726_ & new_n21731_;
  assign new_n21733_ = ~new_n21722_ & ~new_n21732_;
  assign new_n21734_ = ~pi0038 & ~new_n21733_;
  assign new_n21735_ = pi0760 & pi0947;
  assign new_n21736_ = ~pi0039 & ~new_n21735_;
  assign new_n21737_ = new_n21237_ & new_n21736_;
  assign new_n21738_ = ~pi0157 & ~new_n17431_;
  assign new_n21739_ = pi0038 & ~new_n21738_;
  assign new_n21740_ = ~new_n21737_ & new_n21739_;
  assign new_n21741_ = ~pi0688 & ~new_n21740_;
  assign new_n21742_ = ~new_n21734_ & new_n21741_;
  assign new_n21743_ = ~new_n21721_ & ~new_n21742_;
  assign new_n21744_ = new_n10197_ & ~new_n21743_;
  assign new_n21745_ = ~pi0157 & ~new_n10197_;
  assign new_n21746_ = ~pi0832 & ~new_n21745_;
  assign new_n21747_ = ~new_n21744_ & new_n21746_;
  assign po0314 = ~new_n21698_ & ~new_n21747_;
  assign new_n21749_ = ~pi0158 & new_n21003_;
  assign new_n21750_ = pi0158 & ~new_n21029_;
  assign new_n21751_ = ~pi0753 & ~new_n21750_;
  assign new_n21752_ = ~new_n21749_ & new_n21751_;
  assign new_n21753_ = ~pi0158 & pi0753;
  assign new_n21754_ = ~new_n17347_ & new_n21753_;
  assign new_n21755_ = ~new_n21752_ & ~new_n21754_;
  assign new_n21756_ = pi0039 & ~new_n21755_;
  assign new_n21757_ = pi0158 & ~new_n17260_;
  assign new_n21758_ = pi0753 & new_n17260_;
  assign new_n21759_ = ~new_n21757_ & ~new_n21758_;
  assign new_n21760_ = new_n20988_ & new_n21759_;
  assign new_n21761_ = ~pi0038 & ~new_n21760_;
  assign new_n21762_ = ~new_n21756_ & new_n21761_;
  assign new_n21763_ = pi0158 & ~new_n17549_;
  assign new_n21764_ = ~pi0753 & pi0947;
  assign new_n21765_ = new_n17431_ & ~new_n21764_;
  assign new_n21766_ = ~new_n21763_ & ~new_n21765_;
  assign new_n21767_ = pi0038 & ~new_n21766_;
  assign new_n21768_ = pi0702 & ~new_n21767_;
  assign new_n21769_ = ~new_n21762_ & new_n21768_;
  assign new_n21770_ = ~pi0158 & ~new_n21047_;
  assign new_n21771_ = pi0158 & ~new_n21064_;
  assign new_n21772_ = pi0753 & ~new_n21771_;
  assign new_n21773_ = ~new_n21770_ & new_n21772_;
  assign new_n21774_ = ~pi0158 & new_n21092_;
  assign new_n21775_ = pi0158 & new_n21108_;
  assign new_n21776_ = ~pi0753 & ~new_n21775_;
  assign new_n21777_ = ~new_n21774_ & new_n21776_;
  assign new_n21778_ = ~new_n21773_ & ~new_n21777_;
  assign new_n21779_ = pi0039 & ~new_n21778_;
  assign new_n21780_ = new_n21049_ & ~new_n21764_;
  assign new_n21781_ = ~pi0039 & ~new_n21757_;
  assign new_n21782_ = ~new_n21780_ & new_n21781_;
  assign new_n21783_ = ~pi0038 & ~new_n21782_;
  assign new_n21784_ = ~new_n21779_ & new_n21783_;
  assign new_n21785_ = pi0753 & pi0947;
  assign new_n21786_ = ~pi0039 & ~new_n21785_;
  assign new_n21787_ = new_n21237_ & new_n21786_;
  assign new_n21788_ = ~pi0158 & ~new_n17431_;
  assign new_n21789_ = pi0038 & ~new_n21788_;
  assign new_n21790_ = ~new_n21787_ & new_n21789_;
  assign new_n21791_ = ~pi0702 & ~new_n21790_;
  assign new_n21792_ = ~new_n21784_ & new_n21791_;
  assign new_n21793_ = ~new_n21769_ & ~new_n21792_;
  assign new_n21794_ = new_n10197_ & ~new_n21793_;
  assign new_n21795_ = ~pi0158 & ~new_n10197_;
  assign new_n21796_ = ~pi0832 & ~new_n21795_;
  assign new_n21797_ = ~new_n21794_ & new_n21796_;
  assign new_n21798_ = ~pi0702 & new_n20915_;
  assign new_n21799_ = ~new_n21764_ & ~new_n21798_;
  assign new_n21800_ = new_n2754_ & ~new_n21799_;
  assign new_n21801_ = ~pi0158 & ~new_n2754_;
  assign new_n21802_ = pi0832 & ~new_n21801_;
  assign new_n21803_ = ~new_n21800_ & new_n21802_;
  assign po0315 = ~new_n21797_ & ~new_n21803_;
  assign new_n21805_ = ~pi0159 & new_n21003_;
  assign new_n21806_ = pi0159 & ~new_n21029_;
  assign new_n21807_ = ~pi0754 & ~new_n21806_;
  assign new_n21808_ = ~new_n21805_ & new_n21807_;
  assign new_n21809_ = ~pi0159 & pi0754;
  assign new_n21810_ = ~new_n17347_ & new_n21809_;
  assign new_n21811_ = ~new_n21808_ & ~new_n21810_;
  assign new_n21812_ = pi0039 & ~new_n21811_;
  assign new_n21813_ = pi0159 & ~new_n17260_;
  assign new_n21814_ = pi0754 & new_n17260_;
  assign new_n21815_ = ~new_n21813_ & ~new_n21814_;
  assign new_n21816_ = new_n20988_ & new_n21815_;
  assign new_n21817_ = ~pi0038 & ~new_n21816_;
  assign new_n21818_ = ~new_n21812_ & new_n21817_;
  assign new_n21819_ = pi0159 & ~new_n17549_;
  assign new_n21820_ = ~pi0754 & pi0947;
  assign new_n21821_ = new_n17431_ & ~new_n21820_;
  assign new_n21822_ = ~new_n21819_ & ~new_n21821_;
  assign new_n21823_ = pi0038 & ~new_n21822_;
  assign new_n21824_ = pi0709 & ~new_n21823_;
  assign new_n21825_ = ~new_n21818_ & new_n21824_;
  assign new_n21826_ = ~pi0159 & ~new_n21047_;
  assign new_n21827_ = pi0159 & ~new_n21064_;
  assign new_n21828_ = pi0754 & ~new_n21827_;
  assign new_n21829_ = ~new_n21826_ & new_n21828_;
  assign new_n21830_ = ~pi0159 & new_n21092_;
  assign new_n21831_ = pi0159 & new_n21108_;
  assign new_n21832_ = ~pi0754 & ~new_n21831_;
  assign new_n21833_ = ~new_n21830_ & new_n21832_;
  assign new_n21834_ = ~new_n21829_ & ~new_n21833_;
  assign new_n21835_ = pi0039 & ~new_n21834_;
  assign new_n21836_ = new_n21049_ & ~new_n21820_;
  assign new_n21837_ = ~pi0039 & ~new_n21813_;
  assign new_n21838_ = ~new_n21836_ & new_n21837_;
  assign new_n21839_ = ~pi0038 & ~new_n21838_;
  assign new_n21840_ = ~new_n21835_ & new_n21839_;
  assign new_n21841_ = pi0754 & pi0947;
  assign new_n21842_ = ~pi0039 & ~new_n21841_;
  assign new_n21843_ = new_n21237_ & new_n21842_;
  assign new_n21844_ = ~pi0159 & ~new_n17431_;
  assign new_n21845_ = pi0038 & ~new_n21844_;
  assign new_n21846_ = ~new_n21843_ & new_n21845_;
  assign new_n21847_ = ~pi0709 & ~new_n21846_;
  assign new_n21848_ = ~new_n21840_ & new_n21847_;
  assign new_n21849_ = ~new_n21825_ & ~new_n21848_;
  assign new_n21850_ = new_n10197_ & ~new_n21849_;
  assign new_n21851_ = ~pi0159 & ~new_n10197_;
  assign new_n21852_ = ~pi0832 & ~new_n21851_;
  assign new_n21853_ = ~new_n21850_ & new_n21852_;
  assign new_n21854_ = ~pi0709 & new_n20915_;
  assign new_n21855_ = ~new_n21820_ & ~new_n21854_;
  assign new_n21856_ = new_n2754_ & ~new_n21855_;
  assign new_n21857_ = ~pi0159 & ~new_n2754_;
  assign new_n21858_ = pi0832 & ~new_n21857_;
  assign new_n21859_ = ~new_n21856_ & new_n21858_;
  assign po0316 = ~new_n21853_ & ~new_n21859_;
  assign new_n21861_ = ~pi0756 & pi0947;
  assign new_n21862_ = ~pi0734 & new_n20915_;
  assign new_n21863_ = ~new_n21861_ & ~new_n21862_;
  assign new_n21864_ = new_n2754_ & ~new_n21863_;
  assign new_n21865_ = ~pi0160 & ~new_n2754_;
  assign new_n21866_ = pi0832 & ~new_n21865_;
  assign new_n21867_ = ~new_n21864_ & new_n21866_;
  assign new_n21868_ = pi0160 & ~new_n17549_;
  assign new_n21869_ = new_n17431_ & ~new_n21861_;
  assign new_n21870_ = pi0038 & ~new_n21869_;
  assign new_n21871_ = ~new_n21868_ & new_n21870_;
  assign new_n21872_ = ~pi0160 & ~new_n21000_;
  assign new_n21873_ = pi0160 & ~new_n21155_;
  assign new_n21874_ = pi0299 & ~new_n21873_;
  assign new_n21875_ = ~new_n21872_ & new_n21874_;
  assign new_n21876_ = ~pi0160 & ~new_n17326_;
  assign new_n21877_ = new_n21018_ & ~new_n21876_;
  assign new_n21878_ = ~pi0756 & ~new_n21877_;
  assign new_n21879_ = ~new_n21875_ & new_n21878_;
  assign new_n21880_ = ~pi0160 & pi0756;
  assign new_n21881_ = ~new_n17347_ & new_n21880_;
  assign new_n21882_ = pi0039 & ~new_n21881_;
  assign new_n21883_ = ~new_n21879_ & new_n21882_;
  assign new_n21884_ = new_n17260_ & new_n21861_;
  assign new_n21885_ = ~pi0160 & ~new_n17260_;
  assign new_n21886_ = ~pi0039 & ~new_n21885_;
  assign new_n21887_ = ~new_n21884_ & new_n21886_;
  assign new_n21888_ = ~pi0038 & ~new_n21887_;
  assign new_n21889_ = ~new_n21883_ & new_n21888_;
  assign new_n21890_ = ~new_n21871_ & ~new_n21889_;
  assign new_n21891_ = pi0734 & ~new_n21890_;
  assign new_n21892_ = ~new_n21066_ & new_n21887_;
  assign new_n21893_ = ~pi0160 & new_n21092_;
  assign new_n21894_ = pi0160 & new_n21108_;
  assign new_n21895_ = ~pi0756 & ~new_n21894_;
  assign new_n21896_ = ~new_n21893_ & new_n21895_;
  assign new_n21897_ = ~pi0160 & new_n21045_;
  assign new_n21898_ = pi0160 & ~new_n21134_;
  assign new_n21899_ = pi0756 & ~new_n21046_;
  assign new_n21900_ = ~new_n21898_ & new_n21899_;
  assign new_n21901_ = ~new_n21897_ & new_n21900_;
  assign new_n21902_ = pi0039 & ~new_n21901_;
  assign new_n21903_ = ~new_n21896_ & new_n21902_;
  assign new_n21904_ = ~new_n21892_ & ~new_n21903_;
  assign new_n21905_ = ~pi0038 & ~new_n21904_;
  assign new_n21906_ = pi0756 & pi0947;
  assign new_n21907_ = ~pi0039 & ~new_n21906_;
  assign new_n21908_ = new_n21237_ & new_n21907_;
  assign new_n21909_ = ~pi0160 & ~new_n17431_;
  assign new_n21910_ = pi0038 & ~new_n21909_;
  assign new_n21911_ = ~new_n21908_ & new_n21910_;
  assign new_n21912_ = ~pi0734 & ~new_n21911_;
  assign new_n21913_ = ~new_n21905_ & new_n21912_;
  assign new_n21914_ = ~new_n21891_ & ~new_n21913_;
  assign new_n21915_ = new_n10197_ & ~new_n21914_;
  assign new_n21916_ = ~pi0160 & ~new_n10197_;
  assign new_n21917_ = ~pi0832 & ~new_n21916_;
  assign new_n21918_ = ~new_n21915_ & new_n21917_;
  assign po0317 = ~new_n21867_ & ~new_n21918_;
  assign new_n21920_ = ~pi0161 & ~new_n17322_;
  assign new_n21921_ = new_n21388_ & ~new_n21920_;
  assign new_n21922_ = new_n21391_ & ~new_n21921_;
  assign new_n21923_ = pi0161 & ~new_n16636_;
  assign new_n21924_ = ~new_n21101_ & ~new_n21923_;
  assign new_n21925_ = new_n3057_ & new_n21924_;
  assign new_n21926_ = ~pi0223 & ~new_n21925_;
  assign new_n21927_ = ~new_n21922_ & new_n21926_;
  assign new_n21928_ = ~pi0161 & ~new_n17294_;
  assign new_n21929_ = new_n21085_ & ~new_n21928_;
  assign new_n21930_ = new_n21083_ & ~new_n21928_;
  assign new_n21931_ = ~pi0299 & ~new_n21930_;
  assign new_n21932_ = ~new_n21929_ & new_n21931_;
  assign new_n21933_ = ~new_n21927_ & new_n21932_;
  assign new_n21934_ = new_n3467_ & new_n21924_;
  assign new_n21935_ = ~pi0215 & ~new_n21934_;
  assign new_n21936_ = pi0161 & new_n21039_;
  assign new_n21937_ = new_n21054_ & ~new_n21936_;
  assign new_n21938_ = ~new_n17333_ & new_n21937_;
  assign new_n21939_ = new_n21935_ & ~new_n21938_;
  assign new_n21940_ = ~pi0161 & ~new_n17338_;
  assign new_n21941_ = new_n20997_ & ~new_n21940_;
  assign new_n21942_ = pi0299 & ~new_n21941_;
  assign new_n21943_ = ~new_n21939_ & new_n21942_;
  assign new_n21944_ = pi0758 & ~new_n21943_;
  assign new_n21945_ = ~new_n21933_ & new_n21944_;
  assign new_n21946_ = ~new_n21056_ & ~new_n21923_;
  assign new_n21947_ = new_n3057_ & ~new_n21946_;
  assign new_n21948_ = new_n21419_ & ~new_n21920_;
  assign new_n21949_ = ~new_n21947_ & ~new_n21948_;
  assign new_n21950_ = ~pi0223 & ~new_n21949_;
  assign new_n21951_ = ~pi0299 & ~new_n21929_;
  assign new_n21952_ = ~new_n21950_ & new_n21951_;
  assign new_n21953_ = ~new_n21038_ & new_n21935_;
  assign new_n21954_ = ~new_n21937_ & new_n21953_;
  assign new_n21955_ = ~new_n21427_ & new_n21941_;
  assign new_n21956_ = pi0299 & ~new_n21955_;
  assign new_n21957_ = ~new_n21954_ & new_n21956_;
  assign new_n21958_ = ~pi0758 & ~new_n21957_;
  assign new_n21959_ = ~new_n21952_ & new_n21958_;
  assign new_n21960_ = pi0039 & ~new_n21959_;
  assign new_n21961_ = ~new_n21945_ & new_n21960_;
  assign new_n21962_ = pi0161 & ~new_n17260_;
  assign new_n21963_ = pi0758 & pi0947;
  assign new_n21964_ = new_n17260_ & new_n21963_;
  assign new_n21965_ = ~pi0039 & ~new_n21964_;
  assign new_n21966_ = ~new_n21962_ & new_n21965_;
  assign new_n21967_ = ~new_n21066_ & new_n21966_;
  assign new_n21968_ = ~pi0038 & ~new_n21967_;
  assign new_n21969_ = ~new_n21961_ & new_n21968_;
  assign new_n21970_ = ~pi0039 & ~new_n21963_;
  assign new_n21971_ = new_n21443_ & new_n21970_;
  assign new_n21972_ = ~pi0161 & ~new_n17431_;
  assign new_n21973_ = pi0038 & ~new_n21972_;
  assign new_n21974_ = ~new_n21971_ & new_n21973_;
  assign new_n21975_ = pi0736 & ~new_n21974_;
  assign new_n21976_ = ~new_n21969_ & new_n21975_;
  assign new_n21977_ = ~new_n20994_ & ~new_n21937_;
  assign new_n21978_ = ~new_n21022_ & ~new_n21977_;
  assign new_n21979_ = ~new_n21024_ & ~new_n21923_;
  assign new_n21980_ = new_n3467_ & new_n21979_;
  assign new_n21981_ = ~pi0215 & ~new_n21980_;
  assign new_n21982_ = ~new_n21978_ & new_n21981_;
  assign new_n21983_ = pi0161 & new_n20999_;
  assign new_n21984_ = new_n21021_ & ~new_n21983_;
  assign new_n21985_ = ~new_n21982_ & new_n21984_;
  assign new_n21986_ = new_n3057_ & ~new_n21979_;
  assign new_n21987_ = ~new_n21921_ & ~new_n21986_;
  assign new_n21988_ = ~pi0223 & ~new_n21987_;
  assign new_n21989_ = new_n21931_ & ~new_n21988_;
  assign new_n21990_ = pi0758 & ~new_n21989_;
  assign new_n21991_ = ~new_n21985_ & new_n21990_;
  assign new_n21992_ = pi0161 & new_n19893_;
  assign new_n21993_ = pi0039 & ~new_n21992_;
  assign new_n21994_ = ~new_n21991_ & new_n21993_;
  assign new_n21995_ = ~pi0038 & ~new_n21966_;
  assign new_n21996_ = ~new_n21994_ & new_n21995_;
  assign new_n21997_ = ~pi0161 & ~new_n17549_;
  assign new_n21998_ = new_n17431_ & ~new_n21963_;
  assign new_n21999_ = pi0038 & ~new_n21998_;
  assign new_n22000_ = ~new_n21997_ & new_n21999_;
  assign new_n22001_ = ~pi0736 & ~new_n22000_;
  assign new_n22002_ = ~new_n21996_ & new_n22001_;
  assign new_n22003_ = ~new_n21976_ & ~new_n22002_;
  assign new_n22004_ = new_n10197_ & ~new_n22003_;
  assign new_n22005_ = ~pi0161 & ~new_n10197_;
  assign new_n22006_ = ~pi0832 & ~new_n22005_;
  assign new_n22007_ = ~new_n22004_ & new_n22006_;
  assign new_n22008_ = pi0736 & new_n20915_;
  assign new_n22009_ = new_n2754_ & ~new_n21963_;
  assign new_n22010_ = ~new_n22008_ & new_n22009_;
  assign new_n22011_ = ~pi0161 & ~new_n2754_;
  assign new_n22012_ = pi0832 & ~new_n22011_;
  assign new_n22013_ = ~new_n22010_ & new_n22012_;
  assign po0318 = new_n22007_ | new_n22013_;
  assign new_n22015_ = pi0162 & ~new_n17549_;
  assign new_n22016_ = ~pi0761 & pi0947;
  assign new_n22017_ = new_n17431_ & ~new_n22016_;
  assign new_n22018_ = pi0038 & ~new_n22017_;
  assign new_n22019_ = ~new_n22015_ & new_n22018_;
  assign new_n22020_ = ~pi0761 & new_n21002_;
  assign new_n22021_ = pi0761 & new_n17347_;
  assign new_n22022_ = ~pi0162 & ~new_n22021_;
  assign new_n22023_ = ~new_n22020_ & new_n22022_;
  assign new_n22024_ = new_n15128_ & ~new_n21155_;
  assign new_n22025_ = ~new_n20990_ & ~new_n22024_;
  assign new_n22026_ = ~pi0761 & ~new_n22025_;
  assign new_n22027_ = pi0039 & ~new_n22026_;
  assign new_n22028_ = ~new_n22023_ & new_n22027_;
  assign new_n22029_ = new_n17260_ & new_n22016_;
  assign new_n22030_ = ~pi0162 & ~new_n17260_;
  assign new_n22031_ = ~pi0039 & ~new_n22030_;
  assign new_n22032_ = ~new_n22029_ & new_n22031_;
  assign new_n22033_ = ~pi0038 & ~new_n22032_;
  assign new_n22034_ = ~new_n22028_ & new_n22033_;
  assign new_n22035_ = ~new_n22019_ & ~new_n22034_;
  assign new_n22036_ = pi0738 & ~new_n22035_;
  assign new_n22037_ = ~new_n21066_ & new_n22032_;
  assign new_n22038_ = ~pi0162 & new_n21092_;
  assign new_n22039_ = pi0162 & new_n21108_;
  assign new_n22040_ = ~pi0761 & ~new_n22039_;
  assign new_n22041_ = ~new_n22038_ & new_n22040_;
  assign new_n22042_ = ~new_n15128_ & ~new_n21047_;
  assign new_n22043_ = pi0162 & ~new_n21134_;
  assign new_n22044_ = pi0761 & ~new_n22043_;
  assign new_n22045_ = ~new_n22042_ & new_n22044_;
  assign new_n22046_ = pi0039 & ~new_n22045_;
  assign new_n22047_ = ~new_n22041_ & new_n22046_;
  assign new_n22048_ = ~new_n22037_ & ~new_n22047_;
  assign new_n22049_ = ~pi0038 & ~new_n22048_;
  assign new_n22050_ = pi0761 & pi0947;
  assign new_n22051_ = ~pi0039 & ~new_n22050_;
  assign new_n22052_ = new_n21237_ & new_n22051_;
  assign new_n22053_ = ~pi0162 & ~new_n17431_;
  assign new_n22054_ = pi0038 & ~new_n22053_;
  assign new_n22055_ = ~new_n22052_ & new_n22054_;
  assign new_n22056_ = ~pi0738 & ~new_n22055_;
  assign new_n22057_ = ~new_n22049_ & new_n22056_;
  assign new_n22058_ = ~new_n22036_ & ~new_n22057_;
  assign new_n22059_ = new_n10197_ & ~new_n22058_;
  assign new_n22060_ = ~pi0162 & ~new_n10197_;
  assign new_n22061_ = ~pi0832 & ~new_n22060_;
  assign new_n22062_ = ~new_n22059_ & new_n22061_;
  assign new_n22063_ = ~pi0738 & new_n20915_;
  assign new_n22064_ = ~new_n22016_ & ~new_n22063_;
  assign new_n22065_ = new_n2754_ & ~new_n22064_;
  assign new_n22066_ = ~pi0162 & ~new_n2754_;
  assign new_n22067_ = pi0832 & ~new_n22066_;
  assign new_n22068_ = ~new_n22065_ & new_n22067_;
  assign po0319 = ~new_n22062_ & ~new_n22068_;
  assign new_n22070_ = ~pi0777 & pi0947;
  assign new_n22071_ = ~pi0737 & new_n20915_;
  assign new_n22072_ = ~new_n22070_ & ~new_n22071_;
  assign new_n22073_ = new_n2754_ & ~new_n22072_;
  assign new_n22074_ = ~pi0163 & ~new_n2754_;
  assign new_n22075_ = pi0832 & ~new_n22074_;
  assign new_n22076_ = ~new_n22073_ & new_n22075_;
  assign new_n22077_ = pi0163 & ~new_n17549_;
  assign new_n22078_ = new_n17431_ & ~new_n22070_;
  assign new_n22079_ = pi0038 & ~new_n22078_;
  assign new_n22080_ = ~new_n22077_ & new_n22079_;
  assign new_n22081_ = ~pi0163 & ~new_n21000_;
  assign new_n22082_ = ~new_n14735_ & ~new_n21028_;
  assign new_n22083_ = ~new_n22081_ & ~new_n22082_;
  assign new_n22084_ = ~pi0163 & ~new_n17326_;
  assign new_n22085_ = new_n21018_ & ~new_n22084_;
  assign new_n22086_ = ~pi0777 & ~new_n22085_;
  assign new_n22087_ = ~new_n22083_ & new_n22086_;
  assign new_n22088_ = ~pi0163 & pi0777;
  assign new_n22089_ = ~new_n17347_ & new_n22088_;
  assign new_n22090_ = pi0039 & ~new_n22089_;
  assign new_n22091_ = ~new_n22087_ & new_n22090_;
  assign new_n22092_ = new_n17260_ & new_n22070_;
  assign new_n22093_ = ~pi0163 & ~new_n17260_;
  assign new_n22094_ = ~pi0039 & ~new_n22093_;
  assign new_n22095_ = ~new_n22092_ & new_n22094_;
  assign new_n22096_ = ~pi0038 & ~new_n22095_;
  assign new_n22097_ = ~new_n22091_ & new_n22096_;
  assign new_n22098_ = ~new_n22080_ & ~new_n22097_;
  assign new_n22099_ = pi0737 & ~new_n22098_;
  assign new_n22100_ = ~new_n21066_ & new_n22095_;
  assign new_n22101_ = ~pi0163 & new_n21092_;
  assign new_n22102_ = pi0163 & new_n21108_;
  assign new_n22103_ = ~pi0777 & ~new_n22102_;
  assign new_n22104_ = ~new_n22101_ & new_n22103_;
  assign new_n22105_ = ~pi0163 & new_n21045_;
  assign new_n22106_ = pi0163 & ~new_n21134_;
  assign new_n22107_ = pi0777 & ~new_n21046_;
  assign new_n22108_ = ~new_n22106_ & new_n22107_;
  assign new_n22109_ = ~new_n22105_ & new_n22108_;
  assign new_n22110_ = pi0039 & ~new_n22109_;
  assign new_n22111_ = ~new_n22104_ & new_n22110_;
  assign new_n22112_ = ~new_n22100_ & ~new_n22111_;
  assign new_n22113_ = ~pi0038 & ~new_n22112_;
  assign new_n22114_ = pi0777 & pi0947;
  assign new_n22115_ = ~pi0039 & ~new_n22114_;
  assign new_n22116_ = new_n21237_ & new_n22115_;
  assign new_n22117_ = ~pi0163 & ~new_n17431_;
  assign new_n22118_ = pi0038 & ~new_n22117_;
  assign new_n22119_ = ~new_n22116_ & new_n22118_;
  assign new_n22120_ = ~pi0737 & ~new_n22119_;
  assign new_n22121_ = ~new_n22113_ & new_n22120_;
  assign new_n22122_ = ~new_n22099_ & ~new_n22121_;
  assign new_n22123_ = new_n10197_ & ~new_n22122_;
  assign new_n22124_ = ~pi0163 & ~new_n10197_;
  assign new_n22125_ = ~pi0832 & ~new_n22124_;
  assign new_n22126_ = ~new_n22123_ & new_n22125_;
  assign po0320 = ~new_n22076_ & ~new_n22126_;
  assign new_n22128_ = ~pi0752 & pi0947;
  assign new_n22129_ = pi0703 & new_n20915_;
  assign new_n22130_ = ~new_n22128_ & ~new_n22129_;
  assign new_n22131_ = new_n2754_ & ~new_n22130_;
  assign new_n22132_ = ~pi0164 & ~new_n2754_;
  assign new_n22133_ = pi0832 & ~new_n22132_;
  assign new_n22134_ = ~new_n22131_ & new_n22133_;
  assign new_n22135_ = ~pi0164 & new_n21097_;
  assign new_n22136_ = pi0164 & new_n21110_;
  assign new_n22137_ = ~pi0038 & ~new_n22136_;
  assign new_n22138_ = ~new_n22135_ & new_n22137_;
  assign new_n22139_ = ~pi0164 & ~new_n21114_;
  assign new_n22140_ = new_n21117_ & ~new_n22139_;
  assign new_n22141_ = ~pi0752 & ~new_n22140_;
  assign new_n22142_ = ~new_n22138_ & new_n22141_;
  assign new_n22143_ = ~pi0164 & new_n21051_;
  assign new_n22144_ = pi0164 & new_n21068_;
  assign new_n22145_ = ~pi0038 & ~new_n22144_;
  assign new_n22146_ = ~new_n22143_ & new_n22145_;
  assign new_n22147_ = ~pi0164 & ~new_n17431_;
  assign new_n22148_ = new_n21074_ & ~new_n22147_;
  assign new_n22149_ = pi0752 & ~new_n22148_;
  assign new_n22150_ = ~new_n22146_ & new_n22149_;
  assign new_n22151_ = ~new_n22142_ & ~new_n22150_;
  assign new_n22152_ = pi0703 & ~new_n22151_;
  assign new_n22153_ = pi0164 & ~new_n21008_;
  assign new_n22154_ = ~pi0752 & ~new_n22153_;
  assign new_n22155_ = ~new_n21009_ & new_n22154_;
  assign new_n22156_ = ~pi0752 & new_n21033_;
  assign new_n22157_ = pi0164 & ~new_n22156_;
  assign new_n22158_ = pi0752 & new_n17551_;
  assign new_n22159_ = ~pi0703 & ~new_n22158_;
  assign new_n22160_ = ~new_n22157_ & new_n22159_;
  assign new_n22161_ = ~new_n22155_ & new_n22160_;
  assign new_n22162_ = ~new_n22152_ & ~new_n22161_;
  assign new_n22163_ = new_n10197_ & ~new_n22162_;
  assign new_n22164_ = ~pi0164 & ~new_n10197_;
  assign new_n22165_ = ~pi0832 & ~new_n22164_;
  assign new_n22166_ = ~new_n22163_ & new_n22165_;
  assign po0321 = ~new_n22134_ & ~new_n22166_;
  assign new_n22168_ = ~pi0774 & pi0947;
  assign new_n22169_ = pi0687 & new_n20915_;
  assign new_n22170_ = ~new_n22168_ & ~new_n22169_;
  assign new_n22171_ = new_n2754_ & ~new_n22170_;
  assign new_n22172_ = ~pi0165 & ~new_n2754_;
  assign new_n22173_ = pi0832 & ~new_n22172_;
  assign new_n22174_ = ~new_n22171_ & new_n22173_;
  assign new_n22175_ = ~pi0165 & new_n21097_;
  assign new_n22176_ = pi0165 & new_n21110_;
  assign new_n22177_ = ~pi0038 & ~new_n22176_;
  assign new_n22178_ = ~new_n22175_ & new_n22177_;
  assign new_n22179_ = ~pi0165 & ~new_n21114_;
  assign new_n22180_ = new_n21117_ & ~new_n22179_;
  assign new_n22181_ = ~pi0774 & ~new_n22180_;
  assign new_n22182_ = ~new_n22178_ & new_n22181_;
  assign new_n22183_ = ~pi0165 & new_n21051_;
  assign new_n22184_ = pi0165 & new_n21068_;
  assign new_n22185_ = ~pi0038 & ~new_n22184_;
  assign new_n22186_ = ~new_n22183_ & new_n22185_;
  assign new_n22187_ = ~pi0165 & ~new_n17431_;
  assign new_n22188_ = new_n21074_ & ~new_n22187_;
  assign new_n22189_ = pi0774 & ~new_n22188_;
  assign new_n22190_ = ~new_n22186_ & new_n22189_;
  assign new_n22191_ = ~new_n22182_ & ~new_n22190_;
  assign new_n22192_ = pi0687 & ~new_n22191_;
  assign new_n22193_ = pi0165 & ~new_n21008_;
  assign new_n22194_ = ~pi0774 & ~new_n22193_;
  assign new_n22195_ = ~new_n21009_ & new_n22194_;
  assign new_n22196_ = ~pi0774 & new_n21033_;
  assign new_n22197_ = pi0165 & ~new_n22196_;
  assign new_n22198_ = pi0774 & new_n17551_;
  assign new_n22199_ = ~pi0687 & ~new_n22198_;
  assign new_n22200_ = ~new_n22197_ & new_n22199_;
  assign new_n22201_ = ~new_n22195_ & new_n22200_;
  assign new_n22202_ = ~new_n22192_ & ~new_n22201_;
  assign new_n22203_ = new_n10197_ & ~new_n22202_;
  assign new_n22204_ = ~pi0165 & ~new_n10197_;
  assign new_n22205_ = ~pi0832 & ~new_n22204_;
  assign new_n22206_ = ~new_n22203_ & new_n22205_;
  assign po0322 = ~new_n22174_ & ~new_n22206_;
  assign new_n22208_ = pi0166 & new_n21039_;
  assign new_n22209_ = new_n21054_ & ~new_n22208_;
  assign new_n22210_ = ~new_n20994_ & ~new_n22209_;
  assign new_n22211_ = ~new_n21022_ & ~new_n22210_;
  assign new_n22212_ = pi0166 & ~new_n16636_;
  assign new_n22213_ = ~new_n21024_ & ~new_n22212_;
  assign new_n22214_ = new_n3467_ & new_n22213_;
  assign new_n22215_ = ~pi0215 & ~new_n22214_;
  assign new_n22216_ = ~new_n22211_ & new_n22215_;
  assign new_n22217_ = pi0166 & new_n20999_;
  assign new_n22218_ = new_n21021_ & ~new_n22217_;
  assign new_n22219_ = ~new_n22216_ & new_n22218_;
  assign new_n22220_ = ~pi0166 & ~new_n17294_;
  assign new_n22221_ = new_n21083_ & ~new_n22220_;
  assign new_n22222_ = ~pi0299 & ~new_n22221_;
  assign new_n22223_ = new_n3057_ & ~new_n22213_;
  assign new_n22224_ = ~pi0166 & ~new_n17322_;
  assign new_n22225_ = new_n21388_ & ~new_n22224_;
  assign new_n22226_ = ~new_n22223_ & ~new_n22225_;
  assign new_n22227_ = ~pi0223 & ~new_n22226_;
  assign new_n22228_ = new_n22222_ & ~new_n22227_;
  assign new_n22229_ = pi0772 & ~new_n22228_;
  assign new_n22230_ = ~new_n22219_ & new_n22229_;
  assign new_n22231_ = ~pi0772 & ~new_n17347_;
  assign new_n22232_ = pi0166 & new_n22231_;
  assign new_n22233_ = pi0039 & ~new_n22232_;
  assign new_n22234_ = ~new_n22230_ & new_n22233_;
  assign new_n22235_ = pi0166 & ~new_n17260_;
  assign new_n22236_ = pi0772 & pi0947;
  assign new_n22237_ = ~pi0039 & ~new_n22236_;
  assign new_n22238_ = ~new_n17261_ & ~new_n22237_;
  assign new_n22239_ = ~new_n22235_ & ~new_n22238_;
  assign new_n22240_ = ~pi0038 & ~new_n22239_;
  assign new_n22241_ = ~new_n22234_ & new_n22240_;
  assign new_n22242_ = ~pi0166 & ~new_n17549_;
  assign new_n22243_ = new_n17431_ & ~new_n22236_;
  assign new_n22244_ = pi0038 & ~new_n22243_;
  assign new_n22245_ = ~new_n22242_ & new_n22244_;
  assign new_n22246_ = ~pi0727 & ~new_n22245_;
  assign new_n22247_ = ~new_n22241_ & new_n22246_;
  assign new_n22248_ = ~new_n21101_ & ~new_n22212_;
  assign new_n22249_ = new_n3467_ & new_n22248_;
  assign new_n22250_ = ~pi0215 & ~new_n22249_;
  assign new_n22251_ = ~new_n21038_ & new_n22250_;
  assign new_n22252_ = ~new_n22209_ & new_n22251_;
  assign new_n22253_ = ~pi0166 & ~new_n17338_;
  assign new_n22254_ = new_n20997_ & ~new_n22253_;
  assign new_n22255_ = ~new_n21427_ & new_n22254_;
  assign new_n22256_ = pi0299 & ~new_n22255_;
  assign new_n22257_ = ~new_n22252_ & new_n22256_;
  assign new_n22258_ = ~new_n21418_ & ~new_n22224_;
  assign new_n22259_ = ~new_n3057_ & ~new_n22258_;
  assign new_n22260_ = new_n3057_ & new_n22248_;
  assign new_n22261_ = ~pi0223 & ~new_n22260_;
  assign new_n22262_ = new_n3057_ & new_n21024_;
  assign new_n22263_ = new_n22261_ & ~new_n22262_;
  assign new_n22264_ = ~new_n22259_ & new_n22263_;
  assign new_n22265_ = ~new_n6206_ & new_n17294_;
  assign new_n22266_ = ~pi0166 & ~new_n22265_;
  assign new_n22267_ = new_n21085_ & ~new_n22266_;
  assign new_n22268_ = ~pi0299 & ~new_n22267_;
  assign new_n22269_ = ~new_n22264_ & new_n22268_;
  assign new_n22270_ = ~pi0772 & ~new_n22269_;
  assign new_n22271_ = ~new_n22257_ & new_n22270_;
  assign new_n22272_ = ~new_n17333_ & new_n22209_;
  assign new_n22273_ = new_n22250_ & ~new_n22272_;
  assign new_n22274_ = pi0299 & ~new_n22254_;
  assign new_n22275_ = ~new_n22273_ & new_n22274_;
  assign new_n22276_ = new_n21391_ & ~new_n22258_;
  assign new_n22277_ = new_n22261_ & ~new_n22276_;
  assign new_n22278_ = new_n22222_ & ~new_n22267_;
  assign new_n22279_ = ~new_n22277_ & new_n22278_;
  assign new_n22280_ = pi0772 & ~new_n22279_;
  assign new_n22281_ = ~new_n22275_ & new_n22280_;
  assign new_n22282_ = pi0039 & ~new_n22281_;
  assign new_n22283_ = ~new_n22271_ & new_n22282_;
  assign new_n22284_ = ~new_n21066_ & new_n22239_;
  assign new_n22285_ = ~pi0038 & ~new_n22284_;
  assign new_n22286_ = ~new_n22283_ & new_n22285_;
  assign new_n22287_ = ~pi0166 & ~new_n17431_;
  assign new_n22288_ = new_n21443_ & new_n22237_;
  assign new_n22289_ = pi0038 & ~new_n22288_;
  assign new_n22290_ = ~new_n22287_ & new_n22289_;
  assign new_n22291_ = pi0727 & ~new_n22290_;
  assign new_n22292_ = ~new_n22286_ & new_n22291_;
  assign new_n22293_ = ~new_n22247_ & ~new_n22292_;
  assign new_n22294_ = new_n10197_ & ~new_n22293_;
  assign new_n22295_ = ~pi0166 & ~new_n10197_;
  assign new_n22296_ = ~pi0832 & ~new_n22295_;
  assign new_n22297_ = ~new_n22294_ & new_n22296_;
  assign new_n22298_ = pi0727 & new_n20915_;
  assign new_n22299_ = new_n2754_ & ~new_n22236_;
  assign new_n22300_ = ~new_n22298_ & new_n22299_;
  assign new_n22301_ = ~pi0166 & ~new_n2754_;
  assign new_n22302_ = pi0832 & ~new_n22301_;
  assign new_n22303_ = ~new_n22300_ & new_n22302_;
  assign po0323 = new_n22297_ | new_n22303_;
  assign new_n22305_ = ~pi0768 & pi0947;
  assign new_n22306_ = pi0705 & new_n20915_;
  assign new_n22307_ = ~new_n22305_ & ~new_n22306_;
  assign new_n22308_ = new_n2754_ & ~new_n22307_;
  assign new_n22309_ = ~pi0167 & ~new_n2754_;
  assign new_n22310_ = pi0832 & ~new_n22309_;
  assign new_n22311_ = ~new_n22308_ & new_n22310_;
  assign new_n22312_ = ~pi0167 & new_n21097_;
  assign new_n22313_ = pi0167 & new_n21110_;
  assign new_n22314_ = ~pi0038 & ~new_n22313_;
  assign new_n22315_ = ~new_n22312_ & new_n22314_;
  assign new_n22316_ = ~pi0167 & ~new_n21114_;
  assign new_n22317_ = new_n21117_ & ~new_n22316_;
  assign new_n22318_ = ~pi0768 & ~new_n22317_;
  assign new_n22319_ = ~new_n22315_ & new_n22318_;
  assign new_n22320_ = ~pi0167 & new_n21051_;
  assign new_n22321_ = pi0167 & new_n21068_;
  assign new_n22322_ = ~pi0038 & ~new_n22321_;
  assign new_n22323_ = ~new_n22320_ & new_n22322_;
  assign new_n22324_ = ~pi0167 & ~new_n17431_;
  assign new_n22325_ = new_n21074_ & ~new_n22324_;
  assign new_n22326_ = pi0768 & ~new_n22325_;
  assign new_n22327_ = ~new_n22323_ & new_n22326_;
  assign new_n22328_ = pi0705 & ~new_n22327_;
  assign new_n22329_ = ~new_n22319_ & new_n22328_;
  assign new_n22330_ = ~pi0167 & ~new_n21005_;
  assign new_n22331_ = pi0167 & new_n21031_;
  assign new_n22332_ = ~pi0038 & ~new_n22331_;
  assign new_n22333_ = ~new_n22330_ & new_n22332_;
  assign new_n22334_ = ~pi0167 & ~new_n17549_;
  assign new_n22335_ = ~new_n21014_ & ~new_n22334_;
  assign new_n22336_ = ~pi0768 & ~new_n22335_;
  assign new_n22337_ = ~new_n22333_ & new_n22336_;
  assign new_n22338_ = pi0768 & ~new_n17551_;
  assign new_n22339_ = ~pi0167 & new_n22338_;
  assign new_n22340_ = ~pi0705 & ~new_n22339_;
  assign new_n22341_ = ~new_n22337_ & new_n22340_;
  assign new_n22342_ = new_n10197_ & ~new_n22341_;
  assign new_n22343_ = ~new_n22329_ & new_n22342_;
  assign new_n22344_ = ~pi0167 & ~new_n10197_;
  assign new_n22345_ = ~pi0832 & ~new_n22344_;
  assign new_n22346_ = ~new_n22343_ & new_n22345_;
  assign po0324 = ~new_n22311_ & ~new_n22346_;
  assign new_n22348_ = pi0763 & pi0947;
  assign new_n22349_ = new_n2754_ & ~new_n22348_;
  assign new_n22350_ = pi0699 & new_n20915_;
  assign new_n22351_ = new_n22349_ & ~new_n22350_;
  assign new_n22352_ = pi0168 & ~new_n2754_;
  assign new_n22353_ = pi0832 & ~new_n22352_;
  assign new_n22354_ = ~new_n22351_ & new_n22353_;
  assign new_n22355_ = ~pi0168 & ~new_n17260_;
  assign new_n22356_ = ~pi0763 & new_n18106_;
  assign new_n22357_ = ~new_n21016_ & ~new_n22356_;
  assign new_n22358_ = ~new_n22355_ & ~new_n22357_;
  assign new_n22359_ = ~new_n21066_ & new_n22358_;
  assign new_n22360_ = pi0168 & ~new_n17338_;
  assign new_n22361_ = new_n20997_ & ~new_n22360_;
  assign new_n22362_ = pi0168 & ~new_n3467_;
  assign new_n22363_ = ~new_n17333_ & new_n22362_;
  assign new_n22364_ = ~new_n17332_ & ~new_n22363_;
  assign new_n22365_ = ~pi0168 & ~new_n16636_;
  assign new_n22366_ = new_n21025_ & ~new_n22365_;
  assign new_n22367_ = ~new_n21055_ & new_n22366_;
  assign new_n22368_ = ~pi0215 & ~new_n22367_;
  assign new_n22369_ = new_n22364_ & new_n22368_;
  assign new_n22370_ = ~new_n22361_ & ~new_n22369_;
  assign new_n22371_ = pi0299 & ~new_n22370_;
  assign new_n22372_ = pi0168 & ~new_n21099_;
  assign new_n22373_ = new_n21088_ & ~new_n22372_;
  assign new_n22374_ = ~new_n22371_ & ~new_n22373_;
  assign new_n22375_ = pi0763 & ~new_n22374_;
  assign new_n22376_ = new_n21057_ & ~new_n22365_;
  assign new_n22377_ = ~new_n21040_ & ~new_n22376_;
  assign new_n22378_ = new_n22364_ & new_n22377_;
  assign new_n22379_ = ~pi0215 & ~new_n22378_;
  assign new_n22380_ = new_n21105_ & ~new_n22361_;
  assign new_n22381_ = ~new_n21020_ & ~new_n22380_;
  assign new_n22382_ = ~new_n22379_ & new_n22381_;
  assign new_n22383_ = pi0299 & ~new_n22382_;
  assign new_n22384_ = ~pi0168 & ~new_n17326_;
  assign new_n22385_ = new_n21063_ & ~new_n22384_;
  assign new_n22386_ = ~pi0763 & ~new_n22385_;
  assign new_n22387_ = ~new_n22383_ & new_n22386_;
  assign new_n22388_ = pi0039 & ~new_n22387_;
  assign new_n22389_ = ~new_n22375_ & new_n22388_;
  assign new_n22390_ = ~new_n22359_ & ~new_n22389_;
  assign new_n22391_ = ~pi0038 & ~new_n22390_;
  assign new_n22392_ = ~pi0763 & pi0947;
  assign new_n22393_ = ~pi0039 & ~new_n22392_;
  assign new_n22394_ = new_n21237_ & new_n22393_;
  assign new_n22395_ = ~pi0168 & ~new_n17431_;
  assign new_n22396_ = pi0038 & ~new_n22395_;
  assign new_n22397_ = ~new_n22394_ & new_n22396_;
  assign new_n22398_ = ~new_n22391_ & ~new_n22397_;
  assign new_n22399_ = pi0699 & ~new_n22398_;
  assign new_n22400_ = new_n21018_ & ~new_n22384_;
  assign new_n22401_ = new_n22364_ & ~new_n22366_;
  assign new_n22402_ = new_n20995_ & new_n22401_;
  assign new_n22403_ = new_n20999_ & ~new_n22360_;
  assign new_n22404_ = pi0299 & ~new_n22403_;
  assign new_n22405_ = ~new_n22402_ & new_n22404_;
  assign new_n22406_ = pi0763 & ~new_n22405_;
  assign new_n22407_ = ~new_n22400_ & new_n22406_;
  assign new_n22408_ = ~pi0168 & ~pi0763;
  assign new_n22409_ = ~new_n17347_ & new_n22408_;
  assign new_n22410_ = pi0039 & ~new_n22409_;
  assign new_n22411_ = ~new_n22407_ & new_n22410_;
  assign new_n22412_ = ~pi0038 & ~new_n22358_;
  assign new_n22413_ = ~new_n22411_ & new_n22412_;
  assign new_n22414_ = pi0168 & ~new_n17549_;
  assign new_n22415_ = new_n6257_ & new_n22349_;
  assign new_n22416_ = pi0038 & ~new_n22415_;
  assign new_n22417_ = ~new_n22414_ & new_n22416_;
  assign new_n22418_ = ~pi0699 & ~new_n22417_;
  assign new_n22419_ = ~new_n22413_ & new_n22418_;
  assign new_n22420_ = new_n21153_ & ~new_n22419_;
  assign new_n22421_ = ~new_n22399_ & new_n22420_;
  assign new_n22422_ = ~pi0168 & ~new_n21153_;
  assign new_n22423_ = ~pi0057 & ~new_n22422_;
  assign new_n22424_ = ~new_n22421_ & new_n22423_;
  assign new_n22425_ = pi0057 & pi0168;
  assign new_n22426_ = ~pi0832 & ~new_n22425_;
  assign new_n22427_ = ~new_n22424_ & new_n22426_;
  assign po0325 = new_n22354_ | new_n22427_;
  assign new_n22429_ = pi0746 & pi0947;
  assign new_n22430_ = new_n2754_ & ~new_n22429_;
  assign new_n22431_ = pi0729 & new_n20915_;
  assign new_n22432_ = new_n22430_ & ~new_n22431_;
  assign new_n22433_ = pi0169 & ~new_n2754_;
  assign new_n22434_ = pi0832 & ~new_n22433_;
  assign new_n22435_ = ~new_n22432_ & new_n22434_;
  assign new_n22436_ = ~pi0169 & ~new_n17260_;
  assign new_n22437_ = ~pi0746 & new_n18106_;
  assign new_n22438_ = ~new_n21016_ & ~new_n22437_;
  assign new_n22439_ = ~new_n22436_ & ~new_n22438_;
  assign new_n22440_ = ~new_n21066_ & new_n22439_;
  assign new_n22441_ = pi0169 & ~new_n17338_;
  assign new_n22442_ = new_n20997_ & ~new_n22441_;
  assign new_n22443_ = pi0169 & ~new_n3467_;
  assign new_n22444_ = ~new_n17333_ & new_n22443_;
  assign new_n22445_ = ~new_n17332_ & ~new_n22444_;
  assign new_n22446_ = ~pi0169 & ~new_n16636_;
  assign new_n22447_ = new_n21025_ & ~new_n22446_;
  assign new_n22448_ = ~new_n21055_ & new_n22447_;
  assign new_n22449_ = ~pi0215 & ~new_n22448_;
  assign new_n22450_ = new_n22445_ & new_n22449_;
  assign new_n22451_ = ~new_n22442_ & ~new_n22450_;
  assign new_n22452_ = pi0299 & ~new_n22451_;
  assign new_n22453_ = pi0169 & ~new_n21099_;
  assign new_n22454_ = new_n21088_ & ~new_n22453_;
  assign new_n22455_ = ~new_n22452_ & ~new_n22454_;
  assign new_n22456_ = pi0746 & ~new_n22455_;
  assign new_n22457_ = new_n21057_ & ~new_n22446_;
  assign new_n22458_ = ~new_n21040_ & ~new_n22457_;
  assign new_n22459_ = new_n22445_ & new_n22458_;
  assign new_n22460_ = ~pi0215 & ~new_n22459_;
  assign new_n22461_ = new_n21105_ & ~new_n22442_;
  assign new_n22462_ = ~new_n21020_ & ~new_n22461_;
  assign new_n22463_ = ~new_n22460_ & new_n22462_;
  assign new_n22464_ = pi0299 & ~new_n22463_;
  assign new_n22465_ = ~pi0169 & ~new_n17326_;
  assign new_n22466_ = new_n21063_ & ~new_n22465_;
  assign new_n22467_ = ~pi0746 & ~new_n22466_;
  assign new_n22468_ = ~new_n22464_ & new_n22467_;
  assign new_n22469_ = pi0039 & ~new_n22468_;
  assign new_n22470_ = ~new_n22456_ & new_n22469_;
  assign new_n22471_ = ~new_n22440_ & ~new_n22470_;
  assign new_n22472_ = ~pi0038 & ~new_n22471_;
  assign new_n22473_ = ~pi0746 & pi0947;
  assign new_n22474_ = ~pi0039 & ~new_n22473_;
  assign new_n22475_ = new_n21237_ & new_n22474_;
  assign new_n22476_ = ~pi0169 & ~new_n17431_;
  assign new_n22477_ = pi0038 & ~new_n22476_;
  assign new_n22478_ = ~new_n22475_ & new_n22477_;
  assign new_n22479_ = ~new_n22472_ & ~new_n22478_;
  assign new_n22480_ = pi0729 & ~new_n22479_;
  assign new_n22481_ = new_n21018_ & ~new_n22465_;
  assign new_n22482_ = new_n22445_ & ~new_n22447_;
  assign new_n22483_ = new_n20995_ & new_n22482_;
  assign new_n22484_ = new_n20999_ & ~new_n22441_;
  assign new_n22485_ = pi0299 & ~new_n22484_;
  assign new_n22486_ = ~new_n22483_ & new_n22485_;
  assign new_n22487_ = pi0746 & ~new_n22486_;
  assign new_n22488_ = ~new_n22481_ & new_n22487_;
  assign new_n22489_ = ~pi0169 & ~pi0746;
  assign new_n22490_ = ~new_n17347_ & new_n22489_;
  assign new_n22491_ = pi0039 & ~new_n22490_;
  assign new_n22492_ = ~new_n22488_ & new_n22491_;
  assign new_n22493_ = ~pi0038 & ~new_n22439_;
  assign new_n22494_ = ~new_n22492_ & new_n22493_;
  assign new_n22495_ = pi0169 & ~new_n17549_;
  assign new_n22496_ = new_n6257_ & new_n22430_;
  assign new_n22497_ = pi0038 & ~new_n22496_;
  assign new_n22498_ = ~new_n22495_ & new_n22497_;
  assign new_n22499_ = ~pi0729 & ~new_n22498_;
  assign new_n22500_ = ~new_n22494_ & new_n22499_;
  assign new_n22501_ = new_n21153_ & ~new_n22500_;
  assign new_n22502_ = ~new_n22480_ & new_n22501_;
  assign new_n22503_ = ~pi0169 & ~new_n21153_;
  assign new_n22504_ = ~pi0057 & ~new_n22503_;
  assign new_n22505_ = ~new_n22502_ & new_n22504_;
  assign new_n22506_ = pi0057 & pi0169;
  assign new_n22507_ = ~pi0832 & ~new_n22506_;
  assign new_n22508_ = ~new_n22505_ & new_n22507_;
  assign po0326 = new_n22435_ | new_n22508_;
  assign new_n22510_ = pi0730 & new_n20915_;
  assign new_n22511_ = pi0748 & pi0947;
  assign new_n22512_ = new_n2754_ & ~new_n22511_;
  assign new_n22513_ = ~new_n22510_ & new_n22512_;
  assign new_n22514_ = pi0170 & ~new_n2754_;
  assign new_n22515_ = pi0832 & ~new_n22514_;
  assign new_n22516_ = ~new_n22513_ & new_n22515_;
  assign new_n22517_ = pi0170 & ~new_n3467_;
  assign new_n22518_ = ~new_n17333_ & new_n22517_;
  assign new_n22519_ = ~new_n17332_ & ~new_n22518_;
  assign new_n22520_ = ~pi0170 & ~new_n16636_;
  assign new_n22521_ = new_n21057_ & ~new_n22520_;
  assign new_n22522_ = ~new_n21040_ & ~new_n22521_;
  assign new_n22523_ = new_n22519_ & new_n22522_;
  assign new_n22524_ = ~pi0215 & ~new_n22523_;
  assign new_n22525_ = pi0170 & ~new_n17338_;
  assign new_n22526_ = new_n20997_ & ~new_n22525_;
  assign new_n22527_ = new_n21105_ & ~new_n22526_;
  assign new_n22528_ = ~new_n21020_ & ~new_n22527_;
  assign new_n22529_ = ~new_n22524_ & new_n22528_;
  assign new_n22530_ = pi0299 & ~new_n22529_;
  assign new_n22531_ = ~pi0170 & ~new_n17326_;
  assign new_n22532_ = ~pi0299 & ~new_n22531_;
  assign new_n22533_ = ~new_n21062_ & new_n22532_;
  assign new_n22534_ = ~new_n22530_ & ~new_n22533_;
  assign new_n22535_ = pi0039 & ~new_n22534_;
  assign new_n22536_ = ~pi0170 & ~new_n17260_;
  assign new_n22537_ = new_n21067_ & ~new_n22536_;
  assign new_n22538_ = ~new_n22535_ & ~new_n22537_;
  assign new_n22539_ = ~pi0038 & ~new_n22538_;
  assign new_n22540_ = ~pi0170 & ~new_n17431_;
  assign new_n22541_ = new_n21074_ & ~new_n22540_;
  assign new_n22542_ = ~pi0748 & ~new_n22541_;
  assign new_n22543_ = ~new_n22539_ & new_n22542_;
  assign new_n22544_ = new_n21095_ & ~new_n22536_;
  assign new_n22545_ = pi0170 & ~new_n21099_;
  assign new_n22546_ = new_n21088_ & ~new_n22545_;
  assign new_n22547_ = new_n21025_ & ~new_n22520_;
  assign new_n22548_ = ~new_n21055_ & new_n22547_;
  assign new_n22549_ = ~pi0215 & ~new_n22548_;
  assign new_n22550_ = new_n22519_ & new_n22549_;
  assign new_n22551_ = ~new_n22526_ & ~new_n22550_;
  assign new_n22552_ = pi0299 & ~new_n22551_;
  assign new_n22553_ = pi0039 & ~new_n22552_;
  assign new_n22554_ = ~new_n22546_ & new_n22553_;
  assign new_n22555_ = ~new_n22544_ & ~new_n22554_;
  assign new_n22556_ = ~pi0038 & ~new_n22555_;
  assign new_n22557_ = new_n21117_ & ~new_n22540_;
  assign new_n22558_ = pi0748 & ~new_n22557_;
  assign new_n22559_ = ~new_n22556_ & new_n22558_;
  assign new_n22560_ = pi0730 & ~new_n22559_;
  assign new_n22561_ = ~new_n22543_ & new_n22560_;
  assign new_n22562_ = new_n21016_ & ~new_n22536_;
  assign new_n22563_ = new_n22519_ & ~new_n22547_;
  assign new_n22564_ = new_n20995_ & new_n22563_;
  assign new_n22565_ = new_n20999_ & ~new_n22525_;
  assign new_n22566_ = pi0299 & ~new_n22565_;
  assign new_n22567_ = ~new_n22564_ & new_n22566_;
  assign new_n22568_ = ~new_n21017_ & new_n22532_;
  assign new_n22569_ = ~new_n22567_ & ~new_n22568_;
  assign new_n22570_ = pi0039 & ~new_n22569_;
  assign new_n22571_ = ~new_n22562_ & ~new_n22570_;
  assign new_n22572_ = ~pi0038 & ~new_n22571_;
  assign new_n22573_ = ~pi0170 & ~new_n17549_;
  assign new_n22574_ = ~new_n21014_ & ~new_n22573_;
  assign new_n22575_ = pi0748 & ~new_n22574_;
  assign new_n22576_ = ~new_n22572_ & new_n22575_;
  assign new_n22577_ = ~pi0170 & ~pi0748;
  assign new_n22578_ = ~new_n17551_ & new_n22577_;
  assign new_n22579_ = ~pi0730 & ~new_n22578_;
  assign new_n22580_ = ~new_n22576_ & new_n22579_;
  assign new_n22581_ = new_n21153_ & ~new_n22580_;
  assign new_n22582_ = ~new_n22561_ & new_n22581_;
  assign new_n22583_ = ~pi0170 & ~new_n21153_;
  assign new_n22584_ = ~pi0057 & ~new_n22583_;
  assign new_n22585_ = ~new_n22582_ & new_n22584_;
  assign new_n22586_ = pi0057 & pi0170;
  assign new_n22587_ = ~pi0832 & ~new_n22586_;
  assign new_n22588_ = ~new_n22585_ & new_n22587_;
  assign po0327 = new_n22516_ | new_n22588_;
  assign new_n22590_ = pi0764 & pi0947;
  assign new_n22591_ = new_n2754_ & ~new_n22590_;
  assign new_n22592_ = pi0691 & new_n20915_;
  assign new_n22593_ = new_n22591_ & ~new_n22592_;
  assign new_n22594_ = pi0171 & ~new_n2754_;
  assign new_n22595_ = pi0832 & ~new_n22594_;
  assign new_n22596_ = ~new_n22593_ & new_n22595_;
  assign new_n22597_ = ~pi0171 & ~new_n17260_;
  assign new_n22598_ = ~pi0764 & new_n18106_;
  assign new_n22599_ = ~new_n21016_ & ~new_n22598_;
  assign new_n22600_ = ~new_n22597_ & ~new_n22599_;
  assign new_n22601_ = ~new_n21066_ & new_n22600_;
  assign new_n22602_ = pi0171 & ~new_n17338_;
  assign new_n22603_ = new_n20997_ & ~new_n22602_;
  assign new_n22604_ = pi0171 & ~new_n3467_;
  assign new_n22605_ = ~new_n17333_ & new_n22604_;
  assign new_n22606_ = ~new_n17332_ & ~new_n22605_;
  assign new_n22607_ = ~pi0171 & ~new_n16636_;
  assign new_n22608_ = new_n21025_ & ~new_n22607_;
  assign new_n22609_ = ~new_n21055_ & new_n22608_;
  assign new_n22610_ = ~pi0215 & ~new_n22609_;
  assign new_n22611_ = new_n22606_ & new_n22610_;
  assign new_n22612_ = ~new_n22603_ & ~new_n22611_;
  assign new_n22613_ = pi0299 & ~new_n22612_;
  assign new_n22614_ = pi0171 & ~new_n21099_;
  assign new_n22615_ = new_n21088_ & ~new_n22614_;
  assign new_n22616_ = ~new_n22613_ & ~new_n22615_;
  assign new_n22617_ = pi0764 & ~new_n22616_;
  assign new_n22618_ = new_n21057_ & ~new_n22607_;
  assign new_n22619_ = ~new_n21040_ & ~new_n22618_;
  assign new_n22620_ = new_n22606_ & new_n22619_;
  assign new_n22621_ = ~pi0215 & ~new_n22620_;
  assign new_n22622_ = new_n21105_ & ~new_n22603_;
  assign new_n22623_ = ~new_n21020_ & ~new_n22622_;
  assign new_n22624_ = ~new_n22621_ & new_n22623_;
  assign new_n22625_ = pi0299 & ~new_n22624_;
  assign new_n22626_ = ~pi0171 & ~new_n17326_;
  assign new_n22627_ = new_n21063_ & ~new_n22626_;
  assign new_n22628_ = ~pi0764 & ~new_n22627_;
  assign new_n22629_ = ~new_n22625_ & new_n22628_;
  assign new_n22630_ = pi0039 & ~new_n22629_;
  assign new_n22631_ = ~new_n22617_ & new_n22630_;
  assign new_n22632_ = ~new_n22601_ & ~new_n22631_;
  assign new_n22633_ = ~pi0038 & ~new_n22632_;
  assign new_n22634_ = ~pi0764 & pi0947;
  assign new_n22635_ = ~pi0039 & ~new_n22634_;
  assign new_n22636_ = new_n21237_ & new_n22635_;
  assign new_n22637_ = ~pi0171 & ~new_n17431_;
  assign new_n22638_ = pi0038 & ~new_n22637_;
  assign new_n22639_ = ~new_n22636_ & new_n22638_;
  assign new_n22640_ = ~new_n22633_ & ~new_n22639_;
  assign new_n22641_ = pi0691 & ~new_n22640_;
  assign new_n22642_ = new_n21018_ & ~new_n22626_;
  assign new_n22643_ = new_n22606_ & ~new_n22608_;
  assign new_n22644_ = new_n20995_ & new_n22643_;
  assign new_n22645_ = new_n20999_ & ~new_n22602_;
  assign new_n22646_ = pi0299 & ~new_n22645_;
  assign new_n22647_ = ~new_n22644_ & new_n22646_;
  assign new_n22648_ = pi0764 & ~new_n22647_;
  assign new_n22649_ = ~new_n22642_ & new_n22648_;
  assign new_n22650_ = ~pi0171 & ~pi0764;
  assign new_n22651_ = ~new_n17347_ & new_n22650_;
  assign new_n22652_ = pi0039 & ~new_n22651_;
  assign new_n22653_ = ~new_n22649_ & new_n22652_;
  assign new_n22654_ = ~pi0038 & ~new_n22600_;
  assign new_n22655_ = ~new_n22653_ & new_n22654_;
  assign new_n22656_ = pi0171 & ~new_n17549_;
  assign new_n22657_ = new_n6257_ & new_n22591_;
  assign new_n22658_ = pi0038 & ~new_n22657_;
  assign new_n22659_ = ~new_n22656_ & new_n22658_;
  assign new_n22660_ = ~pi0691 & ~new_n22659_;
  assign new_n22661_ = ~new_n22655_ & new_n22660_;
  assign new_n22662_ = new_n21153_ & ~new_n22661_;
  assign new_n22663_ = ~new_n22641_ & new_n22662_;
  assign new_n22664_ = ~pi0171 & ~new_n21153_;
  assign new_n22665_ = ~pi0057 & ~new_n22664_;
  assign new_n22666_ = ~new_n22663_ & new_n22665_;
  assign new_n22667_ = pi0057 & pi0171;
  assign new_n22668_ = ~pi0832 & ~new_n22667_;
  assign new_n22669_ = ~new_n22666_ & new_n22668_;
  assign po0328 = new_n22596_ | new_n22669_;
  assign new_n22671_ = pi0739 & pi0947;
  assign new_n22672_ = new_n2754_ & ~new_n22671_;
  assign new_n22673_ = pi0690 & new_n20915_;
  assign new_n22674_ = new_n22672_ & ~new_n22673_;
  assign new_n22675_ = pi0172 & ~new_n2754_;
  assign new_n22676_ = pi0832 & ~new_n22675_;
  assign new_n22677_ = ~new_n22674_ & new_n22676_;
  assign new_n22678_ = new_n17260_ & new_n22671_;
  assign new_n22679_ = ~pi0172 & ~new_n17260_;
  assign new_n22680_ = ~pi0039 & ~new_n22679_;
  assign new_n22681_ = ~new_n22678_ & new_n22680_;
  assign new_n22682_ = ~new_n21066_ & new_n22681_;
  assign new_n22683_ = pi0172 & ~new_n17338_;
  assign new_n22684_ = new_n20997_ & ~new_n22683_;
  assign new_n22685_ = pi0172 & ~new_n3467_;
  assign new_n22686_ = ~new_n17333_ & new_n22685_;
  assign new_n22687_ = ~new_n17332_ & ~new_n22686_;
  assign new_n22688_ = ~pi0172 & ~new_n16636_;
  assign new_n22689_ = new_n21025_ & ~new_n22688_;
  assign new_n22690_ = ~new_n21055_ & new_n22689_;
  assign new_n22691_ = ~pi0215 & ~new_n22690_;
  assign new_n22692_ = new_n22687_ & new_n22691_;
  assign new_n22693_ = ~new_n22684_ & ~new_n22692_;
  assign new_n22694_ = pi0299 & ~new_n22693_;
  assign new_n22695_ = pi0172 & ~new_n21099_;
  assign new_n22696_ = new_n21088_ & ~new_n22695_;
  assign new_n22697_ = ~new_n22694_ & ~new_n22696_;
  assign new_n22698_ = pi0739 & ~new_n22697_;
  assign new_n22699_ = new_n21057_ & ~new_n22688_;
  assign new_n22700_ = ~new_n21040_ & ~new_n22699_;
  assign new_n22701_ = new_n22687_ & new_n22700_;
  assign new_n22702_ = ~pi0215 & ~new_n22701_;
  assign new_n22703_ = new_n21105_ & ~new_n22684_;
  assign new_n22704_ = ~new_n21020_ & ~new_n22703_;
  assign new_n22705_ = ~new_n22702_ & new_n22704_;
  assign new_n22706_ = pi0299 & ~new_n22705_;
  assign new_n22707_ = ~pi0172 & ~new_n17326_;
  assign new_n22708_ = new_n21063_ & ~new_n22707_;
  assign new_n22709_ = ~pi0739 & ~new_n22708_;
  assign new_n22710_ = ~new_n22706_ & new_n22709_;
  assign new_n22711_ = pi0039 & ~new_n22710_;
  assign new_n22712_ = ~new_n22698_ & new_n22711_;
  assign new_n22713_ = ~new_n22682_ & ~new_n22712_;
  assign new_n22714_ = ~pi0038 & ~new_n22713_;
  assign new_n22715_ = ~pi0739 & pi0947;
  assign new_n22716_ = ~pi0039 & ~new_n22715_;
  assign new_n22717_ = new_n21237_ & new_n22716_;
  assign new_n22718_ = ~pi0172 & ~new_n17431_;
  assign new_n22719_ = pi0038 & ~new_n22718_;
  assign new_n22720_ = ~new_n22717_ & new_n22719_;
  assign new_n22721_ = ~new_n22714_ & ~new_n22720_;
  assign new_n22722_ = pi0690 & ~new_n22721_;
  assign new_n22723_ = new_n21018_ & ~new_n22707_;
  assign new_n22724_ = new_n22687_ & ~new_n22689_;
  assign new_n22725_ = new_n20995_ & new_n22724_;
  assign new_n22726_ = new_n20999_ & ~new_n22683_;
  assign new_n22727_ = pi0299 & ~new_n22726_;
  assign new_n22728_ = ~new_n22725_ & new_n22727_;
  assign new_n22729_ = pi0739 & ~new_n22728_;
  assign new_n22730_ = ~new_n22723_ & new_n22729_;
  assign new_n22731_ = ~pi0172 & ~pi0739;
  assign new_n22732_ = ~new_n17347_ & new_n22731_;
  assign new_n22733_ = pi0039 & ~new_n22732_;
  assign new_n22734_ = ~new_n22730_ & new_n22733_;
  assign new_n22735_ = ~pi0038 & ~new_n22681_;
  assign new_n22736_ = ~new_n22734_ & new_n22735_;
  assign new_n22737_ = pi0172 & ~new_n17549_;
  assign new_n22738_ = new_n6257_ & new_n22672_;
  assign new_n22739_ = pi0038 & ~new_n22738_;
  assign new_n22740_ = ~new_n22737_ & new_n22739_;
  assign new_n22741_ = ~pi0690 & ~new_n22740_;
  assign new_n22742_ = ~new_n22736_ & new_n22741_;
  assign new_n22743_ = new_n21153_ & ~new_n22742_;
  assign new_n22744_ = ~new_n22722_ & new_n22743_;
  assign new_n22745_ = ~pi0172 & ~new_n21153_;
  assign new_n22746_ = ~pi0057 & ~new_n22745_;
  assign new_n22747_ = ~new_n22744_ & new_n22746_;
  assign new_n22748_ = pi0057 & pi0172;
  assign new_n22749_ = ~pi0832 & ~new_n22748_;
  assign new_n22750_ = ~new_n22747_ & new_n22749_;
  assign po0329 = new_n22677_ | new_n22750_;
  assign new_n22752_ = ~pi0173 & ~new_n17558_;
  assign new_n22753_ = new_n17691_ & ~new_n22752_;
  assign new_n22754_ = ~pi0723 & new_n3272_;
  assign new_n22755_ = new_n22752_ & ~new_n22754_;
  assign new_n22756_ = pi0173 & ~new_n18128_;
  assign new_n22757_ = ~pi0038 & ~new_n22756_;
  assign new_n22758_ = new_n3272_ & ~new_n22757_;
  assign new_n22759_ = ~pi0173 & new_n18124_;
  assign new_n22760_ = ~new_n22758_ & ~new_n22759_;
  assign new_n22761_ = ~pi0173 & ~new_n17431_;
  assign new_n22762_ = new_n17544_ & ~new_n22761_;
  assign new_n22763_ = ~pi0723 & ~new_n22762_;
  assign new_n22764_ = ~new_n22760_ & new_n22763_;
  assign new_n22765_ = ~new_n22755_ & ~new_n22764_;
  assign new_n22766_ = ~pi0778 & new_n22765_;
  assign new_n22767_ = pi0625 & ~new_n22765_;
  assign new_n22768_ = ~pi0625 & new_n22752_;
  assign new_n22769_ = pi1153 & ~new_n22768_;
  assign new_n22770_ = ~new_n22767_ & new_n22769_;
  assign new_n22771_ = ~pi0625 & ~new_n22765_;
  assign new_n22772_ = pi0625 & new_n22752_;
  assign new_n22773_ = ~pi1153 & ~new_n22772_;
  assign new_n22774_ = ~new_n22771_ & new_n22773_;
  assign new_n22775_ = ~new_n22770_ & ~new_n22774_;
  assign new_n22776_ = pi0778 & ~new_n22775_;
  assign new_n22777_ = ~new_n22766_ & ~new_n22776_;
  assign new_n22778_ = ~new_n17618_ & ~new_n22777_;
  assign new_n22779_ = new_n17618_ & ~new_n22752_;
  assign new_n22780_ = ~new_n22778_ & ~new_n22779_;
  assign new_n22781_ = ~new_n17655_ & new_n22780_;
  assign new_n22782_ = new_n17655_ & new_n22752_;
  assign new_n22783_ = ~new_n22781_ & ~new_n22782_;
  assign new_n22784_ = ~new_n17691_ & new_n22783_;
  assign new_n22785_ = ~new_n22753_ & ~new_n22784_;
  assign new_n22786_ = ~new_n17734_ & new_n22785_;
  assign new_n22787_ = new_n17734_ & new_n22752_;
  assign new_n22788_ = ~new_n22786_ & ~new_n22787_;
  assign new_n22789_ = ~pi0792 & new_n22788_;
  assign new_n22790_ = pi0628 & ~new_n22788_;
  assign new_n22791_ = ~pi0628 & new_n22752_;
  assign new_n22792_ = pi1156 & ~new_n22791_;
  assign new_n22793_ = ~new_n22790_ & new_n22792_;
  assign new_n22794_ = ~pi0628 & ~new_n22788_;
  assign new_n22795_ = pi0628 & new_n22752_;
  assign new_n22796_ = ~pi1156 & ~new_n22795_;
  assign new_n22797_ = ~new_n22794_ & new_n22796_;
  assign new_n22798_ = ~new_n22793_ & ~new_n22797_;
  assign new_n22799_ = pi0792 & ~new_n22798_;
  assign new_n22800_ = ~new_n22789_ & ~new_n22799_;
  assign new_n22801_ = ~pi0647 & ~new_n22800_;
  assign new_n22802_ = pi0647 & ~new_n22752_;
  assign new_n22803_ = ~new_n22801_ & ~new_n22802_;
  assign new_n22804_ = ~pi1157 & new_n22803_;
  assign new_n22805_ = pi0647 & ~new_n22800_;
  assign new_n22806_ = ~pi0647 & ~new_n22752_;
  assign new_n22807_ = ~new_n22805_ & ~new_n22806_;
  assign new_n22808_ = pi1157 & new_n22807_;
  assign new_n22809_ = ~new_n22804_ & ~new_n22808_;
  assign new_n22810_ = pi0787 & ~new_n22809_;
  assign new_n22811_ = ~pi0787 & new_n22800_;
  assign new_n22812_ = ~new_n22810_ & ~new_n22811_;
  assign new_n22813_ = ~pi0644 & ~new_n22812_;
  assign new_n22814_ = pi0715 & ~new_n22813_;
  assign new_n22815_ = pi0173 & ~new_n3272_;
  assign new_n22816_ = ~pi0173 & ~new_n17349_;
  assign new_n22817_ = pi0745 & ~new_n22816_;
  assign new_n22818_ = pi0173 & ~new_n17426_;
  assign new_n22819_ = ~pi0173 & ~pi0745;
  assign new_n22820_ = new_n17393_ & new_n22819_;
  assign new_n22821_ = ~new_n22818_ & ~new_n22820_;
  assign new_n22822_ = ~new_n22817_ & new_n22821_;
  assign new_n22823_ = ~pi0038 & ~new_n22822_;
  assign new_n22824_ = ~pi0745 & new_n17433_;
  assign new_n22825_ = pi0038 & ~new_n22761_;
  assign new_n22826_ = ~new_n22824_ & new_n22825_;
  assign new_n22827_ = ~new_n22823_ & ~new_n22826_;
  assign new_n22828_ = new_n3272_ & ~new_n22827_;
  assign new_n22829_ = ~new_n22815_ & ~new_n22828_;
  assign new_n22830_ = ~new_n17590_ & ~new_n22829_;
  assign new_n22831_ = new_n17590_ & ~new_n22752_;
  assign new_n22832_ = ~new_n22830_ & ~new_n22831_;
  assign new_n22833_ = ~pi0785 & ~new_n22832_;
  assign new_n22834_ = ~new_n17591_ & ~new_n22752_;
  assign new_n22835_ = pi0609 & new_n22830_;
  assign new_n22836_ = ~new_n22834_ & ~new_n22835_;
  assign new_n22837_ = pi1155 & ~new_n22836_;
  assign new_n22838_ = ~new_n17603_ & ~new_n22752_;
  assign new_n22839_ = ~pi0609 & new_n22830_;
  assign new_n22840_ = ~new_n22838_ & ~new_n22839_;
  assign new_n22841_ = ~pi1155 & ~new_n22840_;
  assign new_n22842_ = ~new_n22837_ & ~new_n22841_;
  assign new_n22843_ = pi0785 & ~new_n22842_;
  assign new_n22844_ = ~new_n22833_ & ~new_n22843_;
  assign new_n22845_ = ~pi0781 & ~new_n22844_;
  assign new_n22846_ = pi0618 & new_n22844_;
  assign new_n22847_ = ~pi0618 & new_n22752_;
  assign new_n22848_ = pi1154 & ~new_n22847_;
  assign new_n22849_ = ~new_n22846_ & new_n22848_;
  assign new_n22850_ = ~pi0618 & new_n22844_;
  assign new_n22851_ = pi0618 & new_n22752_;
  assign new_n22852_ = ~pi1154 & ~new_n22851_;
  assign new_n22853_ = ~new_n22850_ & new_n22852_;
  assign new_n22854_ = ~new_n22849_ & ~new_n22853_;
  assign new_n22855_ = pi0781 & ~new_n22854_;
  assign new_n22856_ = ~new_n22845_ & ~new_n22855_;
  assign new_n22857_ = ~pi0789 & ~new_n22856_;
  assign new_n22858_ = pi0619 & new_n22856_;
  assign new_n22859_ = ~pi0619 & new_n22752_;
  assign new_n22860_ = pi1159 & ~new_n22859_;
  assign new_n22861_ = ~new_n22858_ & new_n22860_;
  assign new_n22862_ = ~pi0619 & new_n22856_;
  assign new_n22863_ = pi0619 & new_n22752_;
  assign new_n22864_ = ~pi1159 & ~new_n22863_;
  assign new_n22865_ = ~new_n22862_ & new_n22864_;
  assign new_n22866_ = ~new_n22861_ & ~new_n22865_;
  assign new_n22867_ = pi0789 & ~new_n22866_;
  assign new_n22868_ = ~new_n22857_ & ~new_n22867_;
  assign new_n22869_ = ~pi0788 & ~new_n22868_;
  assign new_n22870_ = pi0626 & new_n22868_;
  assign new_n22871_ = ~pi0626 & new_n22752_;
  assign new_n22872_ = pi1158 & ~new_n22871_;
  assign new_n22873_ = ~new_n22870_ & new_n22872_;
  assign new_n22874_ = ~pi0626 & new_n22868_;
  assign new_n22875_ = pi0626 & new_n22752_;
  assign new_n22876_ = ~pi1158 & ~new_n22875_;
  assign new_n22877_ = ~new_n22874_ & new_n22876_;
  assign new_n22878_ = ~new_n22873_ & ~new_n22877_;
  assign new_n22879_ = pi0788 & ~new_n22878_;
  assign new_n22880_ = ~new_n22869_ & ~new_n22879_;
  assign new_n22881_ = ~new_n17762_ & new_n22880_;
  assign new_n22882_ = new_n17762_ & new_n22752_;
  assign new_n22883_ = ~new_n22881_ & ~new_n22882_;
  assign new_n22884_ = ~new_n17804_ & ~new_n22883_;
  assign new_n22885_ = new_n17804_ & new_n22752_;
  assign new_n22886_ = ~new_n22884_ & ~new_n22885_;
  assign new_n22887_ = pi0644 & ~new_n22886_;
  assign new_n22888_ = ~pi0644 & new_n22752_;
  assign new_n22889_ = ~pi0715 & ~new_n22888_;
  assign new_n22890_ = ~new_n22887_ & new_n22889_;
  assign new_n22891_ = pi1160 & ~new_n22890_;
  assign new_n22892_ = ~new_n22814_ & new_n22891_;
  assign new_n22893_ = ~new_n20556_ & new_n22883_;
  assign new_n22894_ = new_n17802_ & ~new_n22803_;
  assign new_n22895_ = new_n17801_ & ~new_n22807_;
  assign new_n22896_ = ~new_n22894_ & ~new_n22895_;
  assign new_n22897_ = ~new_n22893_ & new_n22896_;
  assign new_n22898_ = pi0787 & ~new_n22897_;
  assign new_n22899_ = ~new_n20567_ & ~new_n22880_;
  assign new_n22900_ = ~pi0629 & new_n22793_;
  assign new_n22901_ = pi0629 & new_n22797_;
  assign new_n22902_ = ~new_n22900_ & ~new_n22901_;
  assign new_n22903_ = ~new_n22899_ & new_n22902_;
  assign new_n22904_ = pi0792 & ~new_n22903_;
  assign new_n22905_ = pi0723 & new_n22827_;
  assign new_n22906_ = ~pi0173 & new_n16810_;
  assign new_n22907_ = pi0173 & new_n16928_;
  assign new_n22908_ = pi0745 & ~new_n22907_;
  assign new_n22909_ = ~new_n22906_ & new_n22908_;
  assign new_n22910_ = pi0173 & new_n17007_;
  assign new_n22911_ = ~pi0173 & ~new_n17074_;
  assign new_n22912_ = ~pi0745 & ~new_n22911_;
  assign new_n22913_ = ~new_n22910_ & new_n22912_;
  assign new_n22914_ = pi0039 & ~new_n22913_;
  assign new_n22915_ = ~new_n22909_ & new_n22914_;
  assign new_n22916_ = ~pi0173 & ~new_n17217_;
  assign new_n22917_ = pi0173 & ~new_n17178_;
  assign new_n22918_ = pi0745 & ~new_n22917_;
  assign new_n22919_ = ~new_n22916_ & new_n22918_;
  assign new_n22920_ = ~pi0173 & new_n17227_;
  assign new_n22921_ = pi0173 & new_n17234_;
  assign new_n22922_ = ~pi0745 & ~new_n22921_;
  assign new_n22923_ = ~new_n22920_ & new_n22922_;
  assign new_n22924_ = ~new_n22919_ & ~new_n22923_;
  assign new_n22925_ = ~pi0039 & ~new_n22924_;
  assign new_n22926_ = ~pi0038 & ~new_n22925_;
  assign new_n22927_ = ~new_n22915_ & new_n22926_;
  assign new_n22928_ = ~pi0745 & ~new_n17035_;
  assign new_n22929_ = new_n19383_ & ~new_n22928_;
  assign new_n22930_ = ~pi0173 & ~new_n22929_;
  assign new_n22931_ = ~pi0745 & new_n16913_;
  assign new_n22932_ = ~new_n16916_ & ~new_n22931_;
  assign new_n22933_ = pi0173 & ~new_n22932_;
  assign new_n22934_ = new_n6257_ & new_n22933_;
  assign new_n22935_ = pi0038 & ~new_n22934_;
  assign new_n22936_ = ~new_n22930_ & new_n22935_;
  assign new_n22937_ = ~pi0723 & ~new_n22936_;
  assign new_n22938_ = ~new_n22927_ & new_n22937_;
  assign new_n22939_ = new_n3272_ & ~new_n22938_;
  assign new_n22940_ = ~new_n22905_ & new_n22939_;
  assign new_n22941_ = ~new_n22815_ & ~new_n22940_;
  assign new_n22942_ = ~pi0625 & new_n22941_;
  assign new_n22943_ = pi0625 & new_n22829_;
  assign new_n22944_ = ~pi1153 & ~new_n22943_;
  assign new_n22945_ = ~new_n22942_ & new_n22944_;
  assign new_n22946_ = ~pi0608 & ~new_n22770_;
  assign new_n22947_ = ~new_n22945_ & new_n22946_;
  assign new_n22948_ = pi0625 & new_n22941_;
  assign new_n22949_ = ~pi0625 & new_n22829_;
  assign new_n22950_ = pi1153 & ~new_n22949_;
  assign new_n22951_ = ~new_n22948_ & new_n22950_;
  assign new_n22952_ = pi0608 & ~new_n22774_;
  assign new_n22953_ = ~new_n22951_ & new_n22952_;
  assign new_n22954_ = ~new_n22947_ & ~new_n22953_;
  assign new_n22955_ = pi0778 & ~new_n22954_;
  assign new_n22956_ = ~pi0778 & new_n22941_;
  assign new_n22957_ = ~new_n22955_ & ~new_n22956_;
  assign new_n22958_ = ~pi0609 & ~new_n22957_;
  assign new_n22959_ = pi0609 & new_n22777_;
  assign new_n22960_ = ~pi1155 & ~new_n22959_;
  assign new_n22961_ = ~new_n22958_ & new_n22960_;
  assign new_n22962_ = ~pi0660 & ~new_n22837_;
  assign new_n22963_ = ~new_n22961_ & new_n22962_;
  assign new_n22964_ = pi0609 & ~new_n22957_;
  assign new_n22965_ = ~pi0609 & new_n22777_;
  assign new_n22966_ = pi1155 & ~new_n22965_;
  assign new_n22967_ = ~new_n22964_ & new_n22966_;
  assign new_n22968_ = pi0660 & ~new_n22841_;
  assign new_n22969_ = ~new_n22967_ & new_n22968_;
  assign new_n22970_ = ~new_n22963_ & ~new_n22969_;
  assign new_n22971_ = pi0785 & ~new_n22970_;
  assign new_n22972_ = ~pi0785 & ~new_n22957_;
  assign new_n22973_ = ~new_n22971_ & ~new_n22972_;
  assign new_n22974_ = ~pi0618 & ~new_n22973_;
  assign new_n22975_ = pi0618 & new_n22780_;
  assign new_n22976_ = ~pi1154 & ~new_n22975_;
  assign new_n22977_ = ~new_n22974_ & new_n22976_;
  assign new_n22978_ = ~pi0627 & ~new_n22849_;
  assign new_n22979_ = ~new_n22977_ & new_n22978_;
  assign new_n22980_ = pi0618 & ~new_n22973_;
  assign new_n22981_ = ~pi0618 & new_n22780_;
  assign new_n22982_ = pi1154 & ~new_n22981_;
  assign new_n22983_ = ~new_n22980_ & new_n22982_;
  assign new_n22984_ = pi0627 & ~new_n22853_;
  assign new_n22985_ = ~new_n22983_ & new_n22984_;
  assign new_n22986_ = ~new_n22979_ & ~new_n22985_;
  assign new_n22987_ = pi0781 & ~new_n22986_;
  assign new_n22988_ = ~pi0781 & ~new_n22973_;
  assign new_n22989_ = ~new_n22987_ & ~new_n22988_;
  assign new_n22990_ = pi0619 & ~new_n22989_;
  assign new_n22991_ = ~pi0619 & ~new_n22783_;
  assign new_n22992_ = pi1159 & ~new_n22991_;
  assign new_n22993_ = ~new_n22990_ & new_n22992_;
  assign new_n22994_ = pi0648 & ~new_n22865_;
  assign new_n22995_ = ~new_n22993_ & new_n22994_;
  assign new_n22996_ = ~pi0619 & ~new_n22989_;
  assign new_n22997_ = pi0619 & ~new_n22783_;
  assign new_n22998_ = ~pi1159 & ~new_n22997_;
  assign new_n22999_ = ~new_n22996_ & new_n22998_;
  assign new_n23000_ = ~pi0648 & ~new_n22861_;
  assign new_n23001_ = ~new_n22999_ & new_n23000_;
  assign new_n23002_ = pi0789 & ~new_n23001_;
  assign new_n23003_ = ~new_n22995_ & new_n23002_;
  assign new_n23004_ = ~pi0789 & new_n22989_;
  assign new_n23005_ = new_n17969_ & ~new_n23004_;
  assign new_n23006_ = ~new_n23003_ & new_n23005_;
  assign new_n23007_ = new_n17856_ & new_n22785_;
  assign new_n23008_ = ~new_n17733_ & new_n22878_;
  assign new_n23009_ = ~new_n23007_ & ~new_n23008_;
  assign new_n23010_ = pi0788 & ~new_n23009_;
  assign new_n23011_ = ~new_n20364_ & ~new_n23010_;
  assign new_n23012_ = ~new_n23006_ & new_n23011_;
  assign new_n23013_ = ~new_n22904_ & ~new_n23012_;
  assign new_n23014_ = ~new_n20360_ & ~new_n23013_;
  assign new_n23015_ = ~new_n22898_ & ~new_n23014_;
  assign new_n23016_ = ~pi0644 & new_n23015_;
  assign new_n23017_ = pi0644 & ~new_n22812_;
  assign new_n23018_ = ~pi0715 & ~new_n23017_;
  assign new_n23019_ = ~new_n23016_ & new_n23018_;
  assign new_n23020_ = ~pi0644 & ~new_n22886_;
  assign new_n23021_ = pi0644 & new_n22752_;
  assign new_n23022_ = pi0715 & ~new_n23021_;
  assign new_n23023_ = ~new_n23020_ & new_n23022_;
  assign new_n23024_ = ~pi1160 & ~new_n23023_;
  assign new_n23025_ = ~new_n23019_ & new_n23024_;
  assign new_n23026_ = ~new_n22892_ & ~new_n23025_;
  assign new_n23027_ = pi0790 & ~new_n23026_;
  assign new_n23028_ = pi0644 & new_n22891_;
  assign new_n23029_ = pi0790 & ~new_n23028_;
  assign new_n23030_ = new_n23015_ & ~new_n23029_;
  assign new_n23031_ = ~new_n23027_ & ~new_n23030_;
  assign new_n23032_ = ~po1038 & ~new_n23031_;
  assign new_n23033_ = ~pi0173 & po1038;
  assign new_n23034_ = ~pi0832 & ~new_n23033_;
  assign new_n23035_ = ~new_n23032_ & new_n23034_;
  assign new_n23036_ = ~pi0173 & ~new_n2754_;
  assign new_n23037_ = ~new_n22931_ & ~new_n23036_;
  assign new_n23038_ = ~new_n17858_ & ~new_n23037_;
  assign new_n23039_ = ~pi0785 & ~new_n23038_;
  assign new_n23040_ = new_n17603_ & new_n22931_;
  assign new_n23041_ = new_n23038_ & ~new_n23040_;
  assign new_n23042_ = pi1155 & ~new_n23041_;
  assign new_n23043_ = ~pi1155 & ~new_n23036_;
  assign new_n23044_ = ~new_n23040_ & new_n23043_;
  assign new_n23045_ = ~new_n23042_ & ~new_n23044_;
  assign new_n23046_ = pi0785 & ~new_n23045_;
  assign new_n23047_ = ~new_n23039_ & ~new_n23046_;
  assign new_n23048_ = ~pi0781 & ~new_n23047_;
  assign new_n23049_ = ~new_n17873_ & new_n23047_;
  assign new_n23050_ = pi1154 & ~new_n23049_;
  assign new_n23051_ = ~new_n17876_ & new_n23047_;
  assign new_n23052_ = ~pi1154 & ~new_n23051_;
  assign new_n23053_ = ~new_n23050_ & ~new_n23052_;
  assign new_n23054_ = pi0781 & ~new_n23053_;
  assign new_n23055_ = ~new_n23048_ & ~new_n23054_;
  assign new_n23056_ = ~pi0789 & ~new_n23055_;
  assign new_n23057_ = ~pi0619 & new_n2754_;
  assign new_n23058_ = new_n23055_ & ~new_n23057_;
  assign new_n23059_ = pi1159 & ~new_n23058_;
  assign new_n23060_ = pi0619 & new_n2754_;
  assign new_n23061_ = new_n23055_ & ~new_n23060_;
  assign new_n23062_ = ~pi1159 & ~new_n23061_;
  assign new_n23063_ = ~new_n23059_ & ~new_n23062_;
  assign new_n23064_ = pi0789 & ~new_n23063_;
  assign new_n23065_ = ~new_n23056_ & ~new_n23064_;
  assign new_n23066_ = ~pi0788 & ~new_n23065_;
  assign new_n23067_ = pi0626 & new_n23065_;
  assign new_n23068_ = ~pi0626 & new_n23036_;
  assign new_n23069_ = pi1158 & ~new_n23068_;
  assign new_n23070_ = ~new_n23067_ & new_n23069_;
  assign new_n23071_ = ~pi0626 & new_n23065_;
  assign new_n23072_ = pi0626 & new_n23036_;
  assign new_n23073_ = ~pi1158 & ~new_n23072_;
  assign new_n23074_ = ~new_n23071_ & new_n23073_;
  assign new_n23075_ = ~new_n23070_ & ~new_n23074_;
  assign new_n23076_ = pi0788 & ~new_n23075_;
  assign new_n23077_ = ~new_n23066_ & ~new_n23076_;
  assign new_n23078_ = ~new_n17762_ & new_n23077_;
  assign new_n23079_ = new_n17762_ & new_n23036_;
  assign new_n23080_ = ~new_n23078_ & ~new_n23079_;
  assign new_n23081_ = ~new_n20556_ & new_n23080_;
  assign new_n23082_ = ~pi0723 & new_n16915_;
  assign new_n23083_ = ~new_n23036_ & ~new_n23082_;
  assign new_n23084_ = ~pi0778 & ~new_n23083_;
  assign new_n23085_ = ~pi0625 & new_n23082_;
  assign new_n23086_ = ~new_n23083_ & ~new_n23085_;
  assign new_n23087_ = pi1153 & ~new_n23086_;
  assign new_n23088_ = ~pi1153 & ~new_n23036_;
  assign new_n23089_ = ~new_n23085_ & new_n23088_;
  assign new_n23090_ = pi0778 & ~new_n23089_;
  assign new_n23091_ = ~new_n23087_ & new_n23090_;
  assign new_n23092_ = ~new_n23084_ & ~new_n23091_;
  assign new_n23093_ = ~new_n17844_ & ~new_n23092_;
  assign new_n23094_ = ~new_n17846_ & new_n23093_;
  assign new_n23095_ = ~new_n17848_ & new_n23094_;
  assign new_n23096_ = ~new_n17980_ & new_n23095_;
  assign new_n23097_ = ~new_n18011_ & new_n23096_;
  assign new_n23098_ = ~pi0647 & new_n23097_;
  assign new_n23099_ = pi0647 & new_n23036_;
  assign new_n23100_ = ~pi1157 & ~new_n23099_;
  assign new_n23101_ = ~new_n23098_ & new_n23100_;
  assign new_n23102_ = pi0630 & new_n23101_;
  assign new_n23103_ = pi0647 & ~new_n23097_;
  assign new_n23104_ = ~pi0647 & ~new_n23036_;
  assign new_n23105_ = ~new_n23103_ & ~new_n23104_;
  assign new_n23106_ = new_n17801_ & ~new_n23105_;
  assign new_n23107_ = ~new_n23102_ & ~new_n23106_;
  assign new_n23108_ = ~new_n23081_ & new_n23107_;
  assign new_n23109_ = pi0787 & ~new_n23108_;
  assign new_n23110_ = new_n17856_ & new_n23095_;
  assign new_n23111_ = ~new_n17733_ & new_n23075_;
  assign new_n23112_ = ~new_n23110_ & ~new_n23111_;
  assign new_n23113_ = pi0788 & ~new_n23112_;
  assign new_n23114_ = ~new_n16639_ & ~new_n23083_;
  assign new_n23115_ = pi0625 & new_n23114_;
  assign new_n23116_ = new_n23037_ & ~new_n23114_;
  assign new_n23117_ = ~new_n23115_ & ~new_n23116_;
  assign new_n23118_ = new_n23088_ & ~new_n23117_;
  assign new_n23119_ = ~pi0608 & ~new_n23087_;
  assign new_n23120_ = ~new_n23118_ & new_n23119_;
  assign new_n23121_ = pi1153 & new_n23037_;
  assign new_n23122_ = ~new_n23115_ & new_n23121_;
  assign new_n23123_ = pi0608 & ~new_n23089_;
  assign new_n23124_ = ~new_n23122_ & new_n23123_;
  assign new_n23125_ = ~new_n23120_ & ~new_n23124_;
  assign new_n23126_ = pi0778 & ~new_n23125_;
  assign new_n23127_ = ~pi0778 & ~new_n23116_;
  assign new_n23128_ = ~new_n23126_ & ~new_n23127_;
  assign new_n23129_ = ~pi0609 & ~new_n23128_;
  assign new_n23130_ = pi0609 & ~new_n23092_;
  assign new_n23131_ = ~pi1155 & ~new_n23130_;
  assign new_n23132_ = ~new_n23129_ & new_n23131_;
  assign new_n23133_ = ~pi0660 & ~new_n23042_;
  assign new_n23134_ = ~new_n23132_ & new_n23133_;
  assign new_n23135_ = pi0609 & ~new_n23128_;
  assign new_n23136_ = ~pi0609 & ~new_n23092_;
  assign new_n23137_ = pi1155 & ~new_n23136_;
  assign new_n23138_ = ~new_n23135_ & new_n23137_;
  assign new_n23139_ = pi0660 & ~new_n23044_;
  assign new_n23140_ = ~new_n23138_ & new_n23139_;
  assign new_n23141_ = ~new_n23134_ & ~new_n23140_;
  assign new_n23142_ = pi0785 & ~new_n23141_;
  assign new_n23143_ = ~pi0785 & ~new_n23128_;
  assign new_n23144_ = ~new_n23142_ & ~new_n23143_;
  assign new_n23145_ = ~pi0618 & ~new_n23144_;
  assign new_n23146_ = pi0618 & new_n23093_;
  assign new_n23147_ = ~pi1154 & ~new_n23146_;
  assign new_n23148_ = ~new_n23145_ & new_n23147_;
  assign new_n23149_ = ~pi0627 & ~new_n23050_;
  assign new_n23150_ = ~new_n23148_ & new_n23149_;
  assign new_n23151_ = pi0618 & ~new_n23144_;
  assign new_n23152_ = ~pi0618 & new_n23093_;
  assign new_n23153_ = pi1154 & ~new_n23152_;
  assign new_n23154_ = ~new_n23151_ & new_n23153_;
  assign new_n23155_ = pi0627 & ~new_n23052_;
  assign new_n23156_ = ~new_n23154_ & new_n23155_;
  assign new_n23157_ = ~new_n23150_ & ~new_n23156_;
  assign new_n23158_ = pi0781 & ~new_n23157_;
  assign new_n23159_ = ~pi0781 & ~new_n23144_;
  assign new_n23160_ = ~new_n23158_ & ~new_n23159_;
  assign new_n23161_ = pi0619 & ~new_n23160_;
  assign new_n23162_ = ~pi0619 & new_n23094_;
  assign new_n23163_ = pi1159 & ~new_n23162_;
  assign new_n23164_ = ~new_n23161_ & new_n23163_;
  assign new_n23165_ = pi0648 & ~new_n23062_;
  assign new_n23166_ = ~new_n23164_ & new_n23165_;
  assign new_n23167_ = ~pi0619 & ~new_n23160_;
  assign new_n23168_ = pi0619 & new_n23094_;
  assign new_n23169_ = ~pi1159 & ~new_n23168_;
  assign new_n23170_ = ~new_n23167_ & new_n23169_;
  assign new_n23171_ = ~pi0648 & ~new_n23059_;
  assign new_n23172_ = ~new_n23170_ & new_n23171_;
  assign new_n23173_ = pi0789 & ~new_n23172_;
  assign new_n23174_ = ~new_n23166_ & new_n23173_;
  assign new_n23175_ = ~pi0789 & new_n23160_;
  assign new_n23176_ = new_n17969_ & ~new_n23175_;
  assign new_n23177_ = ~new_n23174_ & new_n23176_;
  assign new_n23178_ = ~new_n23113_ & ~new_n23177_;
  assign new_n23179_ = ~new_n20364_ & ~new_n23178_;
  assign new_n23180_ = new_n18008_ & new_n23077_;
  assign new_n23181_ = new_n20851_ & new_n23096_;
  assign new_n23182_ = ~new_n23180_ & ~new_n23181_;
  assign new_n23183_ = ~pi0629 & ~new_n23182_;
  assign new_n23184_ = new_n20855_ & new_n23096_;
  assign new_n23185_ = new_n18007_ & new_n23077_;
  assign new_n23186_ = ~new_n23184_ & ~new_n23185_;
  assign new_n23187_ = pi0629 & ~new_n23186_;
  assign new_n23188_ = ~new_n23183_ & ~new_n23187_;
  assign new_n23189_ = pi0792 & ~new_n23188_;
  assign new_n23190_ = ~new_n20360_ & ~new_n23189_;
  assign new_n23191_ = ~new_n23179_ & new_n23190_;
  assign new_n23192_ = ~new_n23109_ & ~new_n23191_;
  assign new_n23193_ = pi0644 & new_n23192_;
  assign new_n23194_ = ~pi0787 & ~new_n23097_;
  assign new_n23195_ = pi1157 & ~new_n23105_;
  assign new_n23196_ = ~new_n23101_ & ~new_n23195_;
  assign new_n23197_ = pi0787 & ~new_n23196_;
  assign new_n23198_ = ~new_n23194_ & ~new_n23197_;
  assign new_n23199_ = ~pi0644 & new_n23198_;
  assign new_n23200_ = pi0715 & ~new_n23199_;
  assign new_n23201_ = ~new_n23193_ & new_n23200_;
  assign new_n23202_ = ~new_n17804_ & ~new_n23080_;
  assign new_n23203_ = new_n17804_ & new_n23036_;
  assign new_n23204_ = ~new_n23202_ & ~new_n23203_;
  assign new_n23205_ = pi0644 & ~new_n23204_;
  assign new_n23206_ = ~pi0644 & new_n23036_;
  assign new_n23207_ = ~pi0715 & ~new_n23206_;
  assign new_n23208_ = ~new_n23205_ & new_n23207_;
  assign new_n23209_ = pi1160 & ~new_n23208_;
  assign new_n23210_ = ~new_n23201_ & new_n23209_;
  assign new_n23211_ = ~pi0644 & new_n23192_;
  assign new_n23212_ = pi0644 & new_n23198_;
  assign new_n23213_ = ~pi0715 & ~new_n23212_;
  assign new_n23214_ = ~new_n23211_ & new_n23213_;
  assign new_n23215_ = ~pi0644 & ~new_n23204_;
  assign new_n23216_ = pi0644 & new_n23036_;
  assign new_n23217_ = pi0715 & ~new_n23216_;
  assign new_n23218_ = ~new_n23215_ & new_n23217_;
  assign new_n23219_ = ~pi1160 & ~new_n23218_;
  assign new_n23220_ = ~new_n23214_ & new_n23219_;
  assign new_n23221_ = ~new_n23210_ & ~new_n23220_;
  assign new_n23222_ = pi0790 & ~new_n23221_;
  assign new_n23223_ = ~pi0790 & new_n23192_;
  assign new_n23224_ = pi0832 & ~new_n23223_;
  assign new_n23225_ = ~new_n23222_ & new_n23224_;
  assign po0330 = ~new_n23035_ & ~new_n23225_;
  assign new_n23227_ = pi0174 & ~new_n3272_;
  assign new_n23228_ = pi0759 & new_n17391_;
  assign new_n23229_ = ~new_n21465_ & ~new_n23228_;
  assign new_n23230_ = pi0039 & ~new_n23229_;
  assign new_n23231_ = pi0759 & new_n17226_;
  assign new_n23232_ = ~pi0759 & new_n17260_;
  assign new_n23233_ = ~pi0039 & ~new_n23232_;
  assign new_n23234_ = ~new_n23231_ & new_n23233_;
  assign new_n23235_ = ~new_n23230_ & ~new_n23234_;
  assign new_n23236_ = pi0174 & ~new_n23235_;
  assign new_n23237_ = ~pi0174 & pi0759;
  assign new_n23238_ = new_n17426_ & new_n23237_;
  assign new_n23239_ = ~new_n23236_ & ~new_n23238_;
  assign new_n23240_ = ~pi0038 & ~new_n23239_;
  assign new_n23241_ = pi0759 & new_n16639_;
  assign new_n23242_ = new_n17431_ & ~new_n23241_;
  assign new_n23243_ = ~pi0174 & ~new_n17431_;
  assign new_n23244_ = pi0038 & ~new_n23243_;
  assign new_n23245_ = ~new_n23242_ & new_n23244_;
  assign new_n23246_ = ~new_n23240_ & ~new_n23245_;
  assign new_n23247_ = ~pi0696 & new_n23246_;
  assign new_n23248_ = pi0174 & ~new_n16810_;
  assign new_n23249_ = ~pi0174 & ~new_n16928_;
  assign new_n23250_ = ~pi0759 & ~new_n23249_;
  assign new_n23251_ = ~new_n23248_ & new_n23250_;
  assign new_n23252_ = ~pi0174 & ~new_n17007_;
  assign new_n23253_ = pi0174 & new_n17074_;
  assign new_n23254_ = pi0759 & ~new_n23253_;
  assign new_n23255_ = ~new_n23252_ & new_n23254_;
  assign new_n23256_ = pi0039 & ~new_n23255_;
  assign new_n23257_ = ~new_n23251_ & new_n23256_;
  assign new_n23258_ = pi0174 & ~new_n17217_;
  assign new_n23259_ = ~pi0174 & ~new_n17178_;
  assign new_n23260_ = ~pi0759 & ~new_n23259_;
  assign new_n23261_ = ~new_n23258_ & new_n23260_;
  assign new_n23262_ = pi0174 & new_n17227_;
  assign new_n23263_ = ~pi0174 & new_n17234_;
  assign new_n23264_ = pi0759 & ~new_n23263_;
  assign new_n23265_ = ~new_n23262_ & new_n23264_;
  assign new_n23266_ = ~pi0039 & ~new_n23265_;
  assign new_n23267_ = ~new_n23261_ & new_n23266_;
  assign new_n23268_ = ~pi0038 & ~new_n23267_;
  assign new_n23269_ = ~new_n23257_ & new_n23268_;
  assign new_n23270_ = pi0696 & ~new_n19396_;
  assign new_n23271_ = ~new_n23245_ & new_n23270_;
  assign new_n23272_ = ~new_n23269_ & new_n23271_;
  assign new_n23273_ = new_n3272_ & ~new_n23272_;
  assign new_n23274_ = ~new_n23247_ & new_n23273_;
  assign new_n23275_ = ~new_n23227_ & ~new_n23274_;
  assign new_n23276_ = ~pi0625 & new_n23275_;
  assign new_n23277_ = new_n3272_ & ~new_n23246_;
  assign new_n23278_ = ~new_n23227_ & ~new_n23277_;
  assign new_n23279_ = pi0625 & new_n23278_;
  assign new_n23280_ = ~pi1153 & ~new_n23279_;
  assign new_n23281_ = ~new_n23276_ & new_n23280_;
  assign new_n23282_ = pi0174 & ~new_n17558_;
  assign new_n23283_ = pi0696 & new_n3272_;
  assign new_n23284_ = ~new_n23282_ & ~new_n23283_;
  assign new_n23285_ = pi0174 & ~new_n18124_;
  assign new_n23286_ = ~pi0174 & new_n18128_;
  assign new_n23287_ = ~pi0038 & ~new_n23286_;
  assign new_n23288_ = ~new_n23285_ & new_n23287_;
  assign new_n23289_ = new_n19956_ & ~new_n23243_;
  assign new_n23290_ = new_n23283_ & ~new_n23289_;
  assign new_n23291_ = ~new_n23288_ & new_n23290_;
  assign new_n23292_ = ~new_n23284_ & ~new_n23291_;
  assign new_n23293_ = pi0625 & ~new_n23292_;
  assign new_n23294_ = ~pi0625 & ~new_n23282_;
  assign new_n23295_ = pi1153 & ~new_n23294_;
  assign new_n23296_ = ~new_n23293_ & new_n23295_;
  assign new_n23297_ = ~pi0608 & ~new_n23296_;
  assign new_n23298_ = ~new_n23281_ & new_n23297_;
  assign new_n23299_ = pi0625 & new_n23275_;
  assign new_n23300_ = ~pi0625 & new_n23278_;
  assign new_n23301_ = pi1153 & ~new_n23300_;
  assign new_n23302_ = ~new_n23299_ & new_n23301_;
  assign new_n23303_ = ~pi0625 & ~new_n23292_;
  assign new_n23304_ = pi0625 & ~new_n23282_;
  assign new_n23305_ = ~pi1153 & ~new_n23304_;
  assign new_n23306_ = ~new_n23303_ & new_n23305_;
  assign new_n23307_ = pi0608 & ~new_n23306_;
  assign new_n23308_ = ~new_n23302_ & new_n23307_;
  assign new_n23309_ = ~new_n23298_ & ~new_n23308_;
  assign new_n23310_ = pi0778 & ~new_n23309_;
  assign new_n23311_ = ~pi0778 & new_n23275_;
  assign new_n23312_ = ~new_n23310_ & ~new_n23311_;
  assign new_n23313_ = ~pi0609 & ~new_n23312_;
  assign new_n23314_ = ~pi0778 & new_n23292_;
  assign new_n23315_ = ~new_n23296_ & ~new_n23306_;
  assign new_n23316_ = pi0778 & ~new_n23315_;
  assign new_n23317_ = ~new_n23314_ & ~new_n23316_;
  assign new_n23318_ = pi0609 & new_n23317_;
  assign new_n23319_ = ~pi1155 & ~new_n23318_;
  assign new_n23320_ = ~new_n23313_ & new_n23319_;
  assign new_n23321_ = new_n17590_ & ~new_n23282_;
  assign new_n23322_ = ~new_n17590_ & new_n23278_;
  assign new_n23323_ = ~new_n23321_ & ~new_n23322_;
  assign new_n23324_ = pi0609 & ~new_n23323_;
  assign new_n23325_ = ~pi0609 & ~new_n23282_;
  assign new_n23326_ = pi1155 & ~new_n23325_;
  assign new_n23327_ = ~new_n23324_ & new_n23326_;
  assign new_n23328_ = ~pi0660 & ~new_n23327_;
  assign new_n23329_ = ~new_n23320_ & new_n23328_;
  assign new_n23330_ = pi0609 & ~new_n23312_;
  assign new_n23331_ = ~pi0609 & new_n23317_;
  assign new_n23332_ = pi1155 & ~new_n23331_;
  assign new_n23333_ = ~new_n23330_ & new_n23332_;
  assign new_n23334_ = ~pi0609 & ~new_n23323_;
  assign new_n23335_ = pi0609 & ~new_n23282_;
  assign new_n23336_ = ~pi1155 & ~new_n23335_;
  assign new_n23337_ = ~new_n23334_ & new_n23336_;
  assign new_n23338_ = pi0660 & ~new_n23337_;
  assign new_n23339_ = ~new_n23333_ & new_n23338_;
  assign new_n23340_ = ~new_n23329_ & ~new_n23339_;
  assign new_n23341_ = pi0785 & ~new_n23340_;
  assign new_n23342_ = ~pi0785 & ~new_n23312_;
  assign new_n23343_ = ~new_n23341_ & ~new_n23342_;
  assign new_n23344_ = ~pi0618 & ~new_n23343_;
  assign new_n23345_ = new_n17618_ & ~new_n23282_;
  assign new_n23346_ = ~new_n17618_ & new_n23317_;
  assign new_n23347_ = ~new_n23345_ & ~new_n23346_;
  assign new_n23348_ = pi0618 & ~new_n23347_;
  assign new_n23349_ = ~pi1154 & ~new_n23348_;
  assign new_n23350_ = ~new_n23344_ & new_n23349_;
  assign new_n23351_ = ~pi0785 & new_n23323_;
  assign new_n23352_ = ~new_n23327_ & ~new_n23337_;
  assign new_n23353_ = pi0785 & ~new_n23352_;
  assign new_n23354_ = ~new_n23351_ & ~new_n23353_;
  assign new_n23355_ = pi0618 & new_n23354_;
  assign new_n23356_ = ~pi0618 & ~new_n23282_;
  assign new_n23357_ = pi1154 & ~new_n23356_;
  assign new_n23358_ = ~new_n23355_ & new_n23357_;
  assign new_n23359_ = ~pi0627 & ~new_n23358_;
  assign new_n23360_ = ~new_n23350_ & new_n23359_;
  assign new_n23361_ = pi0618 & ~new_n23343_;
  assign new_n23362_ = ~pi0618 & ~new_n23347_;
  assign new_n23363_ = pi1154 & ~new_n23362_;
  assign new_n23364_ = ~new_n23361_ & new_n23363_;
  assign new_n23365_ = ~pi0618 & new_n23354_;
  assign new_n23366_ = pi0618 & ~new_n23282_;
  assign new_n23367_ = ~pi1154 & ~new_n23366_;
  assign new_n23368_ = ~new_n23365_ & new_n23367_;
  assign new_n23369_ = pi0627 & ~new_n23368_;
  assign new_n23370_ = ~new_n23364_ & new_n23369_;
  assign new_n23371_ = ~new_n23360_ & ~new_n23370_;
  assign new_n23372_ = pi0781 & ~new_n23371_;
  assign new_n23373_ = ~pi0781 & ~new_n23343_;
  assign new_n23374_ = ~new_n23372_ & ~new_n23373_;
  assign new_n23375_ = ~pi0619 & ~new_n23374_;
  assign new_n23376_ = ~new_n17655_ & new_n23347_;
  assign new_n23377_ = new_n17655_ & new_n23282_;
  assign new_n23378_ = ~new_n23376_ & ~new_n23377_;
  assign new_n23379_ = pi0619 & new_n23378_;
  assign new_n23380_ = ~pi1159 & ~new_n23379_;
  assign new_n23381_ = ~new_n23375_ & new_n23380_;
  assign new_n23382_ = ~pi0781 & ~new_n23354_;
  assign new_n23383_ = ~new_n23358_ & ~new_n23368_;
  assign new_n23384_ = pi0781 & ~new_n23383_;
  assign new_n23385_ = ~new_n23382_ & ~new_n23384_;
  assign new_n23386_ = pi0619 & new_n23385_;
  assign new_n23387_ = ~pi0619 & ~new_n23282_;
  assign new_n23388_ = pi1159 & ~new_n23387_;
  assign new_n23389_ = ~new_n23386_ & new_n23388_;
  assign new_n23390_ = ~pi0648 & ~new_n23389_;
  assign new_n23391_ = ~new_n23381_ & new_n23390_;
  assign new_n23392_ = pi0619 & ~new_n23374_;
  assign new_n23393_ = ~pi0619 & new_n23378_;
  assign new_n23394_ = pi1159 & ~new_n23393_;
  assign new_n23395_ = ~new_n23392_ & new_n23394_;
  assign new_n23396_ = ~pi0619 & new_n23385_;
  assign new_n23397_ = pi0619 & ~new_n23282_;
  assign new_n23398_ = ~pi1159 & ~new_n23397_;
  assign new_n23399_ = ~new_n23396_ & new_n23398_;
  assign new_n23400_ = pi0648 & ~new_n23399_;
  assign new_n23401_ = ~new_n23395_ & new_n23400_;
  assign new_n23402_ = ~new_n23391_ & ~new_n23401_;
  assign new_n23403_ = pi0789 & ~new_n23402_;
  assign new_n23404_ = ~pi0789 & ~new_n23374_;
  assign new_n23405_ = ~new_n23403_ & ~new_n23404_;
  assign new_n23406_ = ~pi0788 & new_n23405_;
  assign new_n23407_ = ~pi0626 & new_n23405_;
  assign new_n23408_ = new_n17691_ & ~new_n23282_;
  assign new_n23409_ = ~new_n17691_ & new_n23378_;
  assign new_n23410_ = ~new_n23408_ & ~new_n23409_;
  assign new_n23411_ = pi0626 & new_n23410_;
  assign new_n23412_ = ~pi0641 & ~new_n23411_;
  assign new_n23413_ = ~new_n23407_ & new_n23412_;
  assign new_n23414_ = ~pi0789 & ~new_n23385_;
  assign new_n23415_ = ~new_n23389_ & ~new_n23399_;
  assign new_n23416_ = pi0789 & ~new_n23415_;
  assign new_n23417_ = ~new_n23414_ & ~new_n23416_;
  assign new_n23418_ = ~pi0626 & ~new_n23417_;
  assign new_n23419_ = pi0626 & new_n23282_;
  assign new_n23420_ = pi0641 & ~new_n23419_;
  assign new_n23421_ = ~new_n23418_ & new_n23420_;
  assign new_n23422_ = ~pi1158 & ~new_n23421_;
  assign new_n23423_ = ~new_n23413_ & new_n23422_;
  assign new_n23424_ = pi0626 & new_n23405_;
  assign new_n23425_ = ~pi0626 & new_n23410_;
  assign new_n23426_ = pi0641 & ~new_n23425_;
  assign new_n23427_ = ~new_n23424_ & new_n23426_;
  assign new_n23428_ = pi0626 & ~new_n23417_;
  assign new_n23429_ = ~pi0626 & new_n23282_;
  assign new_n23430_ = ~pi0641 & ~new_n23429_;
  assign new_n23431_ = ~new_n23428_ & new_n23430_;
  assign new_n23432_ = pi1158 & ~new_n23431_;
  assign new_n23433_ = ~new_n23427_ & new_n23432_;
  assign new_n23434_ = ~new_n23423_ & ~new_n23433_;
  assign new_n23435_ = pi0788 & ~new_n23434_;
  assign new_n23436_ = ~new_n23406_ & ~new_n23435_;
  assign new_n23437_ = ~pi0628 & new_n23436_;
  assign new_n23438_ = ~new_n17968_ & ~new_n23417_;
  assign new_n23439_ = new_n17968_ & new_n23282_;
  assign new_n23440_ = ~new_n23438_ & ~new_n23439_;
  assign new_n23441_ = pi0628 & new_n23440_;
  assign new_n23442_ = ~pi1156 & ~new_n23441_;
  assign new_n23443_ = ~new_n23437_ & new_n23442_;
  assign new_n23444_ = ~new_n17734_ & new_n23410_;
  assign new_n23445_ = new_n17734_ & new_n23282_;
  assign new_n23446_ = ~new_n23444_ & ~new_n23445_;
  assign new_n23447_ = pi0628 & new_n23446_;
  assign new_n23448_ = ~pi0628 & ~new_n23282_;
  assign new_n23449_ = pi1156 & ~new_n23448_;
  assign new_n23450_ = ~new_n23447_ & new_n23449_;
  assign new_n23451_ = ~pi0629 & ~new_n23450_;
  assign new_n23452_ = ~new_n23443_ & new_n23451_;
  assign new_n23453_ = pi0628 & new_n23436_;
  assign new_n23454_ = ~pi0628 & new_n23440_;
  assign new_n23455_ = pi1156 & ~new_n23454_;
  assign new_n23456_ = ~new_n23453_ & new_n23455_;
  assign new_n23457_ = ~pi0628 & new_n23446_;
  assign new_n23458_ = pi0628 & ~new_n23282_;
  assign new_n23459_ = ~pi1156 & ~new_n23458_;
  assign new_n23460_ = ~new_n23457_ & new_n23459_;
  assign new_n23461_ = pi0629 & ~new_n23460_;
  assign new_n23462_ = ~new_n23456_ & new_n23461_;
  assign new_n23463_ = ~new_n23452_ & ~new_n23462_;
  assign new_n23464_ = pi0792 & ~new_n23463_;
  assign new_n23465_ = ~pi0792 & new_n23436_;
  assign new_n23466_ = ~new_n23464_ & ~new_n23465_;
  assign new_n23467_ = ~pi0647 & ~new_n23466_;
  assign new_n23468_ = ~new_n17762_ & ~new_n23440_;
  assign new_n23469_ = new_n17762_ & new_n23282_;
  assign new_n23470_ = ~new_n23468_ & ~new_n23469_;
  assign new_n23471_ = pi0647 & new_n23470_;
  assign new_n23472_ = ~pi1157 & ~new_n23471_;
  assign new_n23473_ = ~new_n23467_ & new_n23472_;
  assign new_n23474_ = ~pi0792 & ~new_n23446_;
  assign new_n23475_ = ~new_n23450_ & ~new_n23460_;
  assign new_n23476_ = pi0792 & ~new_n23475_;
  assign new_n23477_ = ~new_n23474_ & ~new_n23476_;
  assign new_n23478_ = pi0647 & new_n23477_;
  assign new_n23479_ = ~pi0647 & ~new_n23282_;
  assign new_n23480_ = pi1157 & ~new_n23479_;
  assign new_n23481_ = ~new_n23478_ & new_n23480_;
  assign new_n23482_ = ~pi0630 & ~new_n23481_;
  assign new_n23483_ = ~new_n23473_ & new_n23482_;
  assign new_n23484_ = pi0647 & ~new_n23466_;
  assign new_n23485_ = ~pi0647 & new_n23470_;
  assign new_n23486_ = pi1157 & ~new_n23485_;
  assign new_n23487_ = ~new_n23484_ & new_n23486_;
  assign new_n23488_ = ~pi0647 & new_n23477_;
  assign new_n23489_ = pi0647 & ~new_n23282_;
  assign new_n23490_ = ~pi1157 & ~new_n23489_;
  assign new_n23491_ = ~new_n23488_ & new_n23490_;
  assign new_n23492_ = pi0630 & ~new_n23491_;
  assign new_n23493_ = ~new_n23487_ & new_n23492_;
  assign new_n23494_ = ~new_n23483_ & ~new_n23493_;
  assign new_n23495_ = pi0787 & ~new_n23494_;
  assign new_n23496_ = ~pi0787 & ~new_n23466_;
  assign new_n23497_ = ~new_n23495_ & ~new_n23496_;
  assign new_n23498_ = ~pi0644 & ~new_n23497_;
  assign new_n23499_ = ~pi0787 & ~new_n23477_;
  assign new_n23500_ = ~new_n23481_ & ~new_n23491_;
  assign new_n23501_ = pi0787 & ~new_n23500_;
  assign new_n23502_ = ~new_n23499_ & ~new_n23501_;
  assign new_n23503_ = pi0644 & new_n23502_;
  assign new_n23504_ = ~pi0715 & ~new_n23503_;
  assign new_n23505_ = ~new_n23498_ & new_n23504_;
  assign new_n23506_ = new_n17804_ & ~new_n23282_;
  assign new_n23507_ = ~new_n17804_ & new_n23470_;
  assign new_n23508_ = ~new_n23506_ & ~new_n23507_;
  assign new_n23509_ = ~pi0644 & ~new_n23508_;
  assign new_n23510_ = pi0644 & ~new_n23282_;
  assign new_n23511_ = pi0715 & ~new_n23510_;
  assign new_n23512_ = ~new_n23509_ & new_n23511_;
  assign new_n23513_ = ~pi1160 & ~new_n23512_;
  assign new_n23514_ = ~new_n23505_ & new_n23513_;
  assign new_n23515_ = pi0644 & ~new_n23497_;
  assign new_n23516_ = ~pi0644 & new_n23502_;
  assign new_n23517_ = pi0715 & ~new_n23516_;
  assign new_n23518_ = ~new_n23515_ & new_n23517_;
  assign new_n23519_ = pi0644 & ~new_n23508_;
  assign new_n23520_ = ~pi0644 & ~new_n23282_;
  assign new_n23521_ = ~pi0715 & ~new_n23520_;
  assign new_n23522_ = ~new_n23519_ & new_n23521_;
  assign new_n23523_ = pi1160 & ~new_n23522_;
  assign new_n23524_ = ~new_n23518_ & new_n23523_;
  assign new_n23525_ = pi0790 & ~new_n23524_;
  assign new_n23526_ = ~new_n23514_ & new_n23525_;
  assign new_n23527_ = ~pi0790 & new_n23497_;
  assign new_n23528_ = new_n6305_ & ~new_n23527_;
  assign new_n23529_ = ~new_n23526_ & new_n23528_;
  assign new_n23530_ = ~pi0174 & ~new_n6305_;
  assign new_n23531_ = ~pi0057 & ~new_n23530_;
  assign new_n23532_ = ~new_n23529_ & new_n23531_;
  assign new_n23533_ = pi0057 & pi0174;
  assign new_n23534_ = ~pi0832 & ~new_n23533_;
  assign new_n23535_ = ~new_n23532_ & new_n23534_;
  assign new_n23536_ = pi0174 & ~new_n2754_;
  assign new_n23537_ = pi0759 & new_n16913_;
  assign new_n23538_ = ~new_n23536_ & ~new_n23537_;
  assign new_n23539_ = pi0696 & new_n16916_;
  assign new_n23540_ = new_n23538_ & ~new_n23539_;
  assign new_n23541_ = pi0625 & new_n23539_;
  assign new_n23542_ = ~new_n23540_ & ~new_n23541_;
  assign new_n23543_ = ~pi1153 & ~new_n23542_;
  assign new_n23544_ = pi0696 & new_n16915_;
  assign new_n23545_ = pi0625 & new_n23544_;
  assign new_n23546_ = pi1153 & ~new_n23536_;
  assign new_n23547_ = ~new_n23545_ & new_n23546_;
  assign new_n23548_ = ~pi0608 & ~new_n23547_;
  assign new_n23549_ = ~new_n23543_ & new_n23548_;
  assign new_n23550_ = pi1153 & new_n23538_;
  assign new_n23551_ = ~new_n23541_ & new_n23550_;
  assign new_n23552_ = ~new_n23536_ & ~new_n23544_;
  assign new_n23553_ = ~new_n23545_ & ~new_n23552_;
  assign new_n23554_ = ~pi1153 & ~new_n23553_;
  assign new_n23555_ = pi0608 & ~new_n23554_;
  assign new_n23556_ = ~new_n23551_ & new_n23555_;
  assign new_n23557_ = ~new_n23549_ & ~new_n23556_;
  assign new_n23558_ = pi0778 & ~new_n23557_;
  assign new_n23559_ = ~pi0778 & ~new_n23540_;
  assign new_n23560_ = ~new_n23558_ & ~new_n23559_;
  assign new_n23561_ = ~pi0609 & ~new_n23560_;
  assign new_n23562_ = ~pi0778 & new_n23552_;
  assign new_n23563_ = ~new_n23547_ & ~new_n23554_;
  assign new_n23564_ = pi0778 & ~new_n23563_;
  assign new_n23565_ = ~new_n23562_ & ~new_n23564_;
  assign new_n23566_ = pi0609 & new_n23565_;
  assign new_n23567_ = ~pi1155 & ~new_n23566_;
  assign new_n23568_ = ~new_n23561_ & new_n23567_;
  assign new_n23569_ = new_n17591_ & new_n23537_;
  assign new_n23570_ = pi1155 & ~new_n23536_;
  assign new_n23571_ = ~new_n23569_ & new_n23570_;
  assign new_n23572_ = ~pi0660 & ~new_n23571_;
  assign new_n23573_ = ~new_n23568_ & new_n23572_;
  assign new_n23574_ = pi0609 & ~new_n23560_;
  assign new_n23575_ = ~pi0609 & new_n23565_;
  assign new_n23576_ = pi1155 & ~new_n23575_;
  assign new_n23577_ = ~new_n23574_ & new_n23576_;
  assign new_n23578_ = new_n17603_ & new_n23537_;
  assign new_n23579_ = ~pi1155 & ~new_n23536_;
  assign new_n23580_ = ~new_n23578_ & new_n23579_;
  assign new_n23581_ = pi0660 & ~new_n23580_;
  assign new_n23582_ = ~new_n23577_ & new_n23581_;
  assign new_n23583_ = ~new_n23573_ & ~new_n23582_;
  assign new_n23584_ = pi0785 & ~new_n23583_;
  assign new_n23585_ = ~pi0785 & ~new_n23560_;
  assign new_n23586_ = ~new_n23584_ & ~new_n23585_;
  assign new_n23587_ = ~pi0618 & ~new_n23586_;
  assign new_n23588_ = ~new_n17618_ & new_n23565_;
  assign new_n23589_ = ~new_n23536_ & ~new_n23588_;
  assign new_n23590_ = pi0618 & ~new_n23589_;
  assign new_n23591_ = ~pi1154 & ~new_n23590_;
  assign new_n23592_ = ~new_n23587_ & new_n23591_;
  assign new_n23593_ = ~new_n20223_ & new_n23537_;
  assign new_n23594_ = new_n20311_ & new_n23593_;
  assign new_n23595_ = pi1154 & ~new_n23536_;
  assign new_n23596_ = ~new_n23594_ & new_n23595_;
  assign new_n23597_ = ~pi0627 & ~new_n23596_;
  assign new_n23598_ = ~new_n23592_ & new_n23597_;
  assign new_n23599_ = pi0618 & ~new_n23586_;
  assign new_n23600_ = ~pi0618 & ~new_n23589_;
  assign new_n23601_ = pi1154 & ~new_n23600_;
  assign new_n23602_ = ~new_n23599_ & new_n23601_;
  assign new_n23603_ = new_n20321_ & new_n23593_;
  assign new_n23604_ = ~pi1154 & ~new_n23536_;
  assign new_n23605_ = ~new_n23603_ & new_n23604_;
  assign new_n23606_ = pi0627 & ~new_n23605_;
  assign new_n23607_ = ~new_n23602_ & new_n23606_;
  assign new_n23608_ = ~new_n23598_ & ~new_n23607_;
  assign new_n23609_ = pi0781 & ~new_n23608_;
  assign new_n23610_ = ~pi0781 & ~new_n23586_;
  assign new_n23611_ = pi0648 & new_n20230_;
  assign new_n23612_ = ~pi0648 & new_n20231_;
  assign new_n23613_ = ~new_n23611_ & ~new_n23612_;
  assign new_n23614_ = new_n17690_ & new_n23613_;
  assign new_n23615_ = pi0789 & ~new_n23614_;
  assign new_n23616_ = ~new_n23610_ & ~new_n23615_;
  assign new_n23617_ = ~new_n23609_ & new_n23616_;
  assign new_n23618_ = new_n19280_ & new_n23565_;
  assign new_n23619_ = ~new_n23613_ & ~new_n23618_;
  assign new_n23620_ = ~new_n20229_ & new_n23593_;
  assign new_n23621_ = new_n20336_ & new_n23620_;
  assign new_n23622_ = new_n17689_ & ~new_n23621_;
  assign new_n23623_ = new_n20346_ & new_n23620_;
  assign new_n23624_ = new_n17688_ & ~new_n23623_;
  assign new_n23625_ = ~new_n23622_ & ~new_n23624_;
  assign new_n23626_ = ~new_n23619_ & new_n23625_;
  assign new_n23627_ = pi0789 & ~new_n23536_;
  assign new_n23628_ = ~new_n23626_ & new_n23627_;
  assign new_n23629_ = new_n17969_ & ~new_n23628_;
  assign new_n23630_ = ~new_n23617_ & new_n23629_;
  assign new_n23631_ = ~new_n17691_ & new_n23618_;
  assign new_n23632_ = ~new_n23536_ & ~new_n23631_;
  assign new_n23633_ = new_n17851_ & ~new_n23632_;
  assign new_n23634_ = new_n20235_ & new_n23593_;
  assign new_n23635_ = pi0626 & new_n23634_;
  assign new_n23636_ = ~new_n23536_ & ~new_n23635_;
  assign new_n23637_ = pi1158 & ~new_n23636_;
  assign new_n23638_ = ~pi0641 & ~new_n23637_;
  assign new_n23639_ = ~new_n23633_ & new_n23638_;
  assign new_n23640_ = new_n17850_ & ~new_n23632_;
  assign new_n23641_ = ~pi0626 & new_n23634_;
  assign new_n23642_ = ~new_n23536_ & ~new_n23641_;
  assign new_n23643_ = ~pi1158 & ~new_n23642_;
  assign new_n23644_ = pi0641 & ~new_n23643_;
  assign new_n23645_ = ~new_n23640_ & new_n23644_;
  assign new_n23646_ = pi0788 & ~new_n23645_;
  assign new_n23647_ = ~new_n23639_ & new_n23646_;
  assign new_n23648_ = ~new_n20364_ & ~new_n23647_;
  assign new_n23649_ = ~new_n23630_ & new_n23648_;
  assign new_n23650_ = ~new_n17968_ & new_n23634_;
  assign new_n23651_ = ~pi0629 & new_n23650_;
  assign new_n23652_ = pi0628 & ~new_n23651_;
  assign new_n23653_ = new_n19281_ & new_n23565_;
  assign new_n23654_ = pi0629 & ~new_n23653_;
  assign new_n23655_ = ~new_n23652_ & ~new_n23654_;
  assign new_n23656_ = ~pi1156 & ~new_n23655_;
  assign new_n23657_ = pi0628 & new_n23653_;
  assign new_n23658_ = ~pi0628 & ~new_n23650_;
  assign new_n23659_ = pi0629 & ~new_n23658_;
  assign new_n23660_ = pi1156 & ~new_n23659_;
  assign new_n23661_ = ~new_n23657_ & new_n23660_;
  assign new_n23662_ = ~new_n23656_ & ~new_n23661_;
  assign new_n23663_ = pi0792 & ~new_n23536_;
  assign new_n23664_ = ~new_n23662_ & new_n23663_;
  assign new_n23665_ = ~new_n23649_ & ~new_n23664_;
  assign new_n23666_ = ~new_n20360_ & ~new_n23665_;
  assign new_n23667_ = ~new_n17762_ & new_n23650_;
  assign new_n23668_ = ~pi0630 & new_n23667_;
  assign new_n23669_ = pi0647 & ~new_n23668_;
  assign new_n23670_ = ~new_n19311_ & new_n23653_;
  assign new_n23671_ = pi0630 & ~new_n23670_;
  assign new_n23672_ = ~new_n23669_ & ~new_n23671_;
  assign new_n23673_ = ~pi1157 & ~new_n23672_;
  assign new_n23674_ = ~pi0630 & ~new_n23670_;
  assign new_n23675_ = pi0647 & ~new_n23674_;
  assign new_n23676_ = pi0630 & new_n23667_;
  assign new_n23677_ = pi1157 & ~new_n23676_;
  assign new_n23678_ = ~new_n23675_ & new_n23677_;
  assign new_n23679_ = ~new_n23673_ & ~new_n23678_;
  assign new_n23680_ = pi0787 & ~new_n23536_;
  assign new_n23681_ = ~new_n23679_ & new_n23680_;
  assign new_n23682_ = ~new_n23666_ & ~new_n23681_;
  assign new_n23683_ = pi0644 & new_n23682_;
  assign new_n23684_ = ~new_n19335_ & new_n23670_;
  assign new_n23685_ = ~new_n23536_ & ~new_n23684_;
  assign new_n23686_ = ~pi0644 & ~new_n23685_;
  assign new_n23687_ = pi0715 & ~new_n23686_;
  assign new_n23688_ = ~new_n23683_ & new_n23687_;
  assign new_n23689_ = ~new_n17762_ & ~new_n17804_;
  assign new_n23690_ = new_n23650_ & new_n23689_;
  assign new_n23691_ = pi0644 & new_n23690_;
  assign new_n23692_ = ~pi0715 & ~new_n23536_;
  assign new_n23693_ = ~new_n23691_ & new_n23692_;
  assign new_n23694_ = pi1160 & ~new_n23693_;
  assign new_n23695_ = ~new_n23688_ & new_n23694_;
  assign new_n23696_ = ~pi0644 & new_n23682_;
  assign new_n23697_ = pi0644 & ~new_n23685_;
  assign new_n23698_ = ~pi0715 & ~new_n23697_;
  assign new_n23699_ = ~new_n23696_ & new_n23698_;
  assign new_n23700_ = ~pi0644 & new_n23690_;
  assign new_n23701_ = pi0715 & ~new_n23536_;
  assign new_n23702_ = ~new_n23700_ & new_n23701_;
  assign new_n23703_ = ~pi1160 & ~new_n23702_;
  assign new_n23704_ = ~new_n23699_ & new_n23703_;
  assign new_n23705_ = ~new_n23695_ & ~new_n23704_;
  assign new_n23706_ = pi0790 & ~new_n23705_;
  assign new_n23707_ = ~pi0790 & new_n23682_;
  assign new_n23708_ = pi0832 & ~new_n23707_;
  assign new_n23709_ = ~new_n23706_ & new_n23708_;
  assign po0331 = ~new_n23535_ & ~new_n23709_;
  assign new_n23711_ = ~pi0175 & ~new_n2754_;
  assign new_n23712_ = pi0766 & new_n16913_;
  assign new_n23713_ = ~new_n23711_ & ~new_n23712_;
  assign new_n23714_ = ~new_n17858_ & ~new_n23713_;
  assign new_n23715_ = ~pi0785 & ~new_n23714_;
  assign new_n23716_ = new_n17603_ & new_n23712_;
  assign new_n23717_ = new_n23714_ & ~new_n23716_;
  assign new_n23718_ = pi1155 & ~new_n23717_;
  assign new_n23719_ = ~pi1155 & ~new_n23711_;
  assign new_n23720_ = ~new_n23716_ & new_n23719_;
  assign new_n23721_ = ~new_n23718_ & ~new_n23720_;
  assign new_n23722_ = pi0785 & ~new_n23721_;
  assign new_n23723_ = ~new_n23715_ & ~new_n23722_;
  assign new_n23724_ = ~pi0781 & ~new_n23723_;
  assign new_n23725_ = ~new_n17873_ & new_n23723_;
  assign new_n23726_ = pi1154 & ~new_n23725_;
  assign new_n23727_ = ~new_n17876_ & new_n23723_;
  assign new_n23728_ = ~pi1154 & ~new_n23727_;
  assign new_n23729_ = ~new_n23726_ & ~new_n23728_;
  assign new_n23730_ = pi0781 & ~new_n23729_;
  assign new_n23731_ = ~new_n23724_ & ~new_n23730_;
  assign new_n23732_ = ~pi0789 & ~new_n23731_;
  assign new_n23733_ = ~new_n23057_ & new_n23731_;
  assign new_n23734_ = pi1159 & ~new_n23733_;
  assign new_n23735_ = ~new_n23060_ & new_n23731_;
  assign new_n23736_ = ~pi1159 & ~new_n23735_;
  assign new_n23737_ = ~new_n23734_ & ~new_n23736_;
  assign new_n23738_ = pi0789 & ~new_n23737_;
  assign new_n23739_ = ~new_n23732_ & ~new_n23738_;
  assign new_n23740_ = ~new_n17968_ & new_n23739_;
  assign new_n23741_ = new_n17968_ & new_n23711_;
  assign new_n23742_ = ~new_n23740_ & ~new_n23741_;
  assign new_n23743_ = ~new_n17762_ & ~new_n23742_;
  assign new_n23744_ = new_n17762_ & new_n23711_;
  assign new_n23745_ = ~new_n23743_ & ~new_n23744_;
  assign new_n23746_ = ~new_n20556_ & new_n23745_;
  assign new_n23747_ = pi0700 & new_n16915_;
  assign new_n23748_ = ~new_n23711_ & ~new_n23747_;
  assign new_n23749_ = ~pi0778 & ~new_n23748_;
  assign new_n23750_ = ~pi0625 & new_n23747_;
  assign new_n23751_ = ~new_n23748_ & ~new_n23750_;
  assign new_n23752_ = pi1153 & ~new_n23751_;
  assign new_n23753_ = ~pi1153 & ~new_n23711_;
  assign new_n23754_ = ~new_n23750_ & new_n23753_;
  assign new_n23755_ = pi0778 & ~new_n23754_;
  assign new_n23756_ = ~new_n23752_ & new_n23755_;
  assign new_n23757_ = ~new_n23749_ & ~new_n23756_;
  assign new_n23758_ = ~new_n17844_ & ~new_n23757_;
  assign new_n23759_ = ~new_n17846_ & new_n23758_;
  assign new_n23760_ = ~new_n17848_ & new_n23759_;
  assign new_n23761_ = ~new_n17980_ & new_n23760_;
  assign new_n23762_ = ~new_n18011_ & new_n23761_;
  assign new_n23763_ = ~pi0647 & new_n23762_;
  assign new_n23764_ = pi0647 & new_n23711_;
  assign new_n23765_ = ~pi1157 & ~new_n23764_;
  assign new_n23766_ = ~new_n23763_ & new_n23765_;
  assign new_n23767_ = pi0630 & new_n23766_;
  assign new_n23768_ = pi0647 & ~new_n23762_;
  assign new_n23769_ = ~pi0647 & ~new_n23711_;
  assign new_n23770_ = ~new_n23768_ & ~new_n23769_;
  assign new_n23771_ = new_n17801_ & ~new_n23770_;
  assign new_n23772_ = ~new_n23767_ & ~new_n23771_;
  assign new_n23773_ = ~new_n23746_ & new_n23772_;
  assign new_n23774_ = pi0787 & ~new_n23773_;
  assign new_n23775_ = pi0626 & ~new_n23739_;
  assign new_n23776_ = ~pi0626 & ~new_n23711_;
  assign new_n23777_ = new_n17731_ & ~new_n23776_;
  assign new_n23778_ = ~new_n23775_ & new_n23777_;
  assign new_n23779_ = new_n17856_ & new_n23760_;
  assign new_n23780_ = ~pi0626 & ~new_n23739_;
  assign new_n23781_ = pi0626 & ~new_n23711_;
  assign new_n23782_ = new_n17732_ & ~new_n23781_;
  assign new_n23783_ = ~new_n23780_ & new_n23782_;
  assign new_n23784_ = ~new_n23779_ & ~new_n23783_;
  assign new_n23785_ = ~new_n23778_ & new_n23784_;
  assign new_n23786_ = pi0788 & ~new_n23785_;
  assign new_n23787_ = ~new_n16639_ & ~new_n23748_;
  assign new_n23788_ = pi0625 & new_n23787_;
  assign new_n23789_ = new_n23713_ & ~new_n23787_;
  assign new_n23790_ = ~new_n23788_ & ~new_n23789_;
  assign new_n23791_ = new_n23753_ & ~new_n23790_;
  assign new_n23792_ = ~pi0608 & ~new_n23752_;
  assign new_n23793_ = ~new_n23791_ & new_n23792_;
  assign new_n23794_ = pi1153 & new_n23713_;
  assign new_n23795_ = ~new_n23788_ & new_n23794_;
  assign new_n23796_ = pi0608 & ~new_n23754_;
  assign new_n23797_ = ~new_n23795_ & new_n23796_;
  assign new_n23798_ = ~new_n23793_ & ~new_n23797_;
  assign new_n23799_ = pi0778 & ~new_n23798_;
  assign new_n23800_ = ~pi0778 & ~new_n23789_;
  assign new_n23801_ = ~new_n23799_ & ~new_n23800_;
  assign new_n23802_ = ~pi0609 & ~new_n23801_;
  assign new_n23803_ = pi0609 & ~new_n23757_;
  assign new_n23804_ = ~pi1155 & ~new_n23803_;
  assign new_n23805_ = ~new_n23802_ & new_n23804_;
  assign new_n23806_ = ~pi0660 & ~new_n23718_;
  assign new_n23807_ = ~new_n23805_ & new_n23806_;
  assign new_n23808_ = pi0609 & ~new_n23801_;
  assign new_n23809_ = ~pi0609 & ~new_n23757_;
  assign new_n23810_ = pi1155 & ~new_n23809_;
  assign new_n23811_ = ~new_n23808_ & new_n23810_;
  assign new_n23812_ = pi0660 & ~new_n23720_;
  assign new_n23813_ = ~new_n23811_ & new_n23812_;
  assign new_n23814_ = ~new_n23807_ & ~new_n23813_;
  assign new_n23815_ = pi0785 & ~new_n23814_;
  assign new_n23816_ = ~pi0785 & ~new_n23801_;
  assign new_n23817_ = ~new_n23815_ & ~new_n23816_;
  assign new_n23818_ = ~pi0618 & ~new_n23817_;
  assign new_n23819_ = pi0618 & new_n23758_;
  assign new_n23820_ = ~pi1154 & ~new_n23819_;
  assign new_n23821_ = ~new_n23818_ & new_n23820_;
  assign new_n23822_ = ~pi0627 & ~new_n23726_;
  assign new_n23823_ = ~new_n23821_ & new_n23822_;
  assign new_n23824_ = pi0618 & ~new_n23817_;
  assign new_n23825_ = ~pi0618 & new_n23758_;
  assign new_n23826_ = pi1154 & ~new_n23825_;
  assign new_n23827_ = ~new_n23824_ & new_n23826_;
  assign new_n23828_ = pi0627 & ~new_n23728_;
  assign new_n23829_ = ~new_n23827_ & new_n23828_;
  assign new_n23830_ = ~new_n23823_ & ~new_n23829_;
  assign new_n23831_ = pi0781 & ~new_n23830_;
  assign new_n23832_ = ~pi0781 & ~new_n23817_;
  assign new_n23833_ = ~new_n23831_ & ~new_n23832_;
  assign new_n23834_ = pi0619 & ~new_n23833_;
  assign new_n23835_ = ~pi0619 & new_n23759_;
  assign new_n23836_ = pi1159 & ~new_n23835_;
  assign new_n23837_ = ~new_n23834_ & new_n23836_;
  assign new_n23838_ = pi0648 & ~new_n23736_;
  assign new_n23839_ = ~new_n23837_ & new_n23838_;
  assign new_n23840_ = ~pi0619 & ~new_n23833_;
  assign new_n23841_ = pi0619 & new_n23759_;
  assign new_n23842_ = ~pi1159 & ~new_n23841_;
  assign new_n23843_ = ~new_n23840_ & new_n23842_;
  assign new_n23844_ = ~pi0648 & ~new_n23734_;
  assign new_n23845_ = ~new_n23843_ & new_n23844_;
  assign new_n23846_ = pi0789 & ~new_n23845_;
  assign new_n23847_ = ~new_n23839_ & new_n23846_;
  assign new_n23848_ = ~pi0789 & new_n23833_;
  assign new_n23849_ = new_n17969_ & ~new_n23848_;
  assign new_n23850_ = ~new_n23847_ & new_n23849_;
  assign new_n23851_ = ~new_n23786_ & ~new_n23850_;
  assign new_n23852_ = ~new_n20364_ & ~new_n23851_;
  assign new_n23853_ = new_n18008_ & ~new_n23742_;
  assign new_n23854_ = new_n20851_ & new_n23761_;
  assign new_n23855_ = ~new_n23853_ & ~new_n23854_;
  assign new_n23856_ = ~pi0629 & ~new_n23855_;
  assign new_n23857_ = new_n20855_ & new_n23761_;
  assign new_n23858_ = new_n18007_ & ~new_n23742_;
  assign new_n23859_ = ~new_n23857_ & ~new_n23858_;
  assign new_n23860_ = pi0629 & ~new_n23859_;
  assign new_n23861_ = ~new_n23856_ & ~new_n23860_;
  assign new_n23862_ = pi0792 & ~new_n23861_;
  assign new_n23863_ = ~new_n20360_ & ~new_n23862_;
  assign new_n23864_ = ~new_n23852_ & new_n23863_;
  assign new_n23865_ = ~new_n23774_ & ~new_n23864_;
  assign new_n23866_ = pi0644 & new_n23865_;
  assign new_n23867_ = ~pi0787 & ~new_n23762_;
  assign new_n23868_ = pi1157 & ~new_n23770_;
  assign new_n23869_ = ~new_n23766_ & ~new_n23868_;
  assign new_n23870_ = pi0787 & ~new_n23869_;
  assign new_n23871_ = ~new_n23867_ & ~new_n23870_;
  assign new_n23872_ = ~pi0644 & new_n23871_;
  assign new_n23873_ = pi0715 & ~new_n23872_;
  assign new_n23874_ = ~new_n23866_ & new_n23873_;
  assign new_n23875_ = ~new_n17804_ & ~new_n23745_;
  assign new_n23876_ = new_n17804_ & new_n23711_;
  assign new_n23877_ = ~new_n23875_ & ~new_n23876_;
  assign new_n23878_ = pi0644 & ~new_n23877_;
  assign new_n23879_ = ~pi0644 & new_n23711_;
  assign new_n23880_ = ~pi0715 & ~new_n23879_;
  assign new_n23881_ = ~new_n23878_ & new_n23880_;
  assign new_n23882_ = pi1160 & ~new_n23881_;
  assign new_n23883_ = ~new_n23874_ & new_n23882_;
  assign new_n23884_ = ~pi0644 & new_n23865_;
  assign new_n23885_ = pi0644 & new_n23871_;
  assign new_n23886_ = ~pi0715 & ~new_n23885_;
  assign new_n23887_ = ~new_n23884_ & new_n23886_;
  assign new_n23888_ = ~pi0644 & ~new_n23877_;
  assign new_n23889_ = pi0644 & new_n23711_;
  assign new_n23890_ = pi0715 & ~new_n23889_;
  assign new_n23891_ = ~new_n23888_ & new_n23890_;
  assign new_n23892_ = ~pi1160 & ~new_n23891_;
  assign new_n23893_ = ~new_n23887_ & new_n23892_;
  assign new_n23894_ = ~new_n23883_ & ~new_n23893_;
  assign new_n23895_ = pi0790 & ~new_n23894_;
  assign new_n23896_ = ~pi0790 & new_n23865_;
  assign new_n23897_ = pi0832 & ~new_n23896_;
  assign new_n23898_ = ~new_n23895_ & new_n23897_;
  assign new_n23899_ = ~pi0175 & ~new_n17558_;
  assign new_n23900_ = new_n17691_ & ~new_n23899_;
  assign new_n23901_ = pi0175 & ~new_n3272_;
  assign new_n23902_ = ~pi0175 & new_n18124_;
  assign new_n23903_ = pi0175 & ~new_n18128_;
  assign new_n23904_ = ~pi0038 & ~new_n23903_;
  assign new_n23905_ = ~new_n23902_ & new_n23904_;
  assign new_n23906_ = ~pi0175 & ~new_n17431_;
  assign new_n23907_ = new_n17544_ & ~new_n23906_;
  assign new_n23908_ = pi0700 & ~new_n23907_;
  assign new_n23909_ = ~new_n23905_ & new_n23908_;
  assign new_n23910_ = ~pi0175 & ~pi0700;
  assign new_n23911_ = ~new_n17551_ & new_n23910_;
  assign new_n23912_ = new_n3272_ & ~new_n23911_;
  assign new_n23913_ = ~new_n23909_ & new_n23912_;
  assign new_n23914_ = ~new_n23901_ & ~new_n23913_;
  assign new_n23915_ = ~pi0778 & ~new_n23914_;
  assign new_n23916_ = pi0625 & new_n23914_;
  assign new_n23917_ = ~pi0625 & new_n23899_;
  assign new_n23918_ = pi1153 & ~new_n23917_;
  assign new_n23919_ = ~new_n23916_ & new_n23918_;
  assign new_n23920_ = ~pi0625 & new_n23914_;
  assign new_n23921_ = pi0625 & new_n23899_;
  assign new_n23922_ = ~pi1153 & ~new_n23921_;
  assign new_n23923_ = ~new_n23920_ & new_n23922_;
  assign new_n23924_ = ~new_n23919_ & ~new_n23923_;
  assign new_n23925_ = pi0778 & ~new_n23924_;
  assign new_n23926_ = ~new_n23915_ & ~new_n23925_;
  assign new_n23927_ = ~new_n17618_ & ~new_n23926_;
  assign new_n23928_ = new_n17618_ & ~new_n23899_;
  assign new_n23929_ = ~new_n23927_ & ~new_n23928_;
  assign new_n23930_ = ~new_n17655_ & new_n23929_;
  assign new_n23931_ = new_n17655_ & new_n23899_;
  assign new_n23932_ = ~new_n23930_ & ~new_n23931_;
  assign new_n23933_ = ~new_n17691_ & new_n23932_;
  assign new_n23934_ = ~new_n23900_ & ~new_n23933_;
  assign new_n23935_ = ~new_n17734_ & new_n23934_;
  assign new_n23936_ = new_n17734_ & new_n23899_;
  assign new_n23937_ = ~new_n23935_ & ~new_n23936_;
  assign new_n23938_ = ~pi0628 & ~new_n23937_;
  assign new_n23939_ = pi0628 & new_n23899_;
  assign new_n23940_ = ~new_n23938_ & ~new_n23939_;
  assign new_n23941_ = ~pi1156 & ~new_n23940_;
  assign new_n23942_ = pi0628 & ~new_n23937_;
  assign new_n23943_ = ~pi0628 & new_n23899_;
  assign new_n23944_ = ~new_n23942_ & ~new_n23943_;
  assign new_n23945_ = pi1156 & ~new_n23944_;
  assign new_n23946_ = ~new_n23941_ & ~new_n23945_;
  assign new_n23947_ = pi0792 & ~new_n23946_;
  assign new_n23948_ = ~pi0792 & ~new_n23937_;
  assign new_n23949_ = ~new_n23947_ & ~new_n23948_;
  assign new_n23950_ = ~pi0647 & ~new_n23949_;
  assign new_n23951_ = pi0647 & new_n23899_;
  assign new_n23952_ = ~new_n23950_ & ~new_n23951_;
  assign new_n23953_ = ~pi1157 & ~new_n23952_;
  assign new_n23954_ = pi0647 & ~new_n23949_;
  assign new_n23955_ = ~pi0647 & new_n23899_;
  assign new_n23956_ = ~new_n23954_ & ~new_n23955_;
  assign new_n23957_ = pi1157 & ~new_n23956_;
  assign new_n23958_ = ~new_n23953_ & ~new_n23957_;
  assign new_n23959_ = pi0787 & ~new_n23958_;
  assign new_n23960_ = ~pi0787 & ~new_n23949_;
  assign new_n23961_ = ~new_n23959_ & ~new_n23960_;
  assign new_n23962_ = ~pi0644 & ~new_n23961_;
  assign new_n23963_ = pi0715 & ~new_n23962_;
  assign new_n23964_ = ~pi0766 & new_n17347_;
  assign new_n23965_ = pi0175 & new_n17424_;
  assign new_n23966_ = ~new_n23964_ & ~new_n23965_;
  assign new_n23967_ = pi0039 & ~new_n23966_;
  assign new_n23968_ = ~pi0175 & pi0766;
  assign new_n23969_ = new_n17393_ & new_n23968_;
  assign new_n23970_ = pi0766 & ~new_n17397_;
  assign new_n23971_ = pi0175 & ~new_n23970_;
  assign new_n23972_ = ~new_n21497_ & ~new_n23971_;
  assign new_n23973_ = ~new_n23969_ & new_n23972_;
  assign new_n23974_ = ~new_n23967_ & new_n23973_;
  assign new_n23975_ = ~pi0038 & ~new_n23974_;
  assign new_n23976_ = pi0766 & new_n17433_;
  assign new_n23977_ = pi0038 & ~new_n23906_;
  assign new_n23978_ = ~new_n23976_ & new_n23977_;
  assign new_n23979_ = ~new_n23975_ & ~new_n23978_;
  assign new_n23980_ = new_n3272_ & ~new_n23979_;
  assign new_n23981_ = ~new_n23901_ & ~new_n23980_;
  assign new_n23982_ = ~new_n17590_ & ~new_n23981_;
  assign new_n23983_ = new_n17590_ & ~new_n23899_;
  assign new_n23984_ = ~new_n23982_ & ~new_n23983_;
  assign new_n23985_ = ~pi0785 & ~new_n23984_;
  assign new_n23986_ = ~new_n17591_ & ~new_n23899_;
  assign new_n23987_ = pi0609 & new_n23982_;
  assign new_n23988_ = ~new_n23986_ & ~new_n23987_;
  assign new_n23989_ = pi1155 & ~new_n23988_;
  assign new_n23990_ = ~new_n17603_ & ~new_n23899_;
  assign new_n23991_ = ~pi0609 & new_n23982_;
  assign new_n23992_ = ~new_n23990_ & ~new_n23991_;
  assign new_n23993_ = ~pi1155 & ~new_n23992_;
  assign new_n23994_ = ~new_n23989_ & ~new_n23993_;
  assign new_n23995_ = pi0785 & ~new_n23994_;
  assign new_n23996_ = ~new_n23985_ & ~new_n23995_;
  assign new_n23997_ = ~pi0781 & ~new_n23996_;
  assign new_n23998_ = pi0618 & new_n23996_;
  assign new_n23999_ = ~pi0618 & new_n23899_;
  assign new_n24000_ = pi1154 & ~new_n23999_;
  assign new_n24001_ = ~new_n23998_ & new_n24000_;
  assign new_n24002_ = ~pi0618 & new_n23996_;
  assign new_n24003_ = pi0618 & new_n23899_;
  assign new_n24004_ = ~pi1154 & ~new_n24003_;
  assign new_n24005_ = ~new_n24002_ & new_n24004_;
  assign new_n24006_ = ~new_n24001_ & ~new_n24005_;
  assign new_n24007_ = pi0781 & ~new_n24006_;
  assign new_n24008_ = ~new_n23997_ & ~new_n24007_;
  assign new_n24009_ = ~pi0789 & ~new_n24008_;
  assign new_n24010_ = pi0619 & new_n24008_;
  assign new_n24011_ = ~pi0619 & new_n23899_;
  assign new_n24012_ = pi1159 & ~new_n24011_;
  assign new_n24013_ = ~new_n24010_ & new_n24012_;
  assign new_n24014_ = ~pi0619 & new_n24008_;
  assign new_n24015_ = pi0619 & new_n23899_;
  assign new_n24016_ = ~pi1159 & ~new_n24015_;
  assign new_n24017_ = ~new_n24014_ & new_n24016_;
  assign new_n24018_ = ~new_n24013_ & ~new_n24017_;
  assign new_n24019_ = pi0789 & ~new_n24018_;
  assign new_n24020_ = ~new_n24009_ & ~new_n24019_;
  assign new_n24021_ = ~new_n17968_ & new_n24020_;
  assign new_n24022_ = new_n17968_ & new_n23899_;
  assign new_n24023_ = ~new_n24021_ & ~new_n24022_;
  assign new_n24024_ = ~new_n17762_ & ~new_n24023_;
  assign new_n24025_ = new_n17762_ & new_n23899_;
  assign new_n24026_ = ~new_n24024_ & ~new_n24025_;
  assign new_n24027_ = ~new_n17804_ & ~new_n24026_;
  assign new_n24028_ = new_n17804_ & new_n23899_;
  assign new_n24029_ = ~new_n24027_ & ~new_n24028_;
  assign new_n24030_ = pi0644 & ~new_n24029_;
  assign new_n24031_ = ~pi0644 & new_n23899_;
  assign new_n24032_ = ~pi0715 & ~new_n24031_;
  assign new_n24033_ = ~new_n24030_ & new_n24032_;
  assign new_n24034_ = pi1160 & ~new_n24033_;
  assign new_n24035_ = ~new_n23963_ & new_n24034_;
  assign new_n24036_ = pi0644 & ~new_n23961_;
  assign new_n24037_ = ~pi0715 & ~new_n24036_;
  assign new_n24038_ = ~pi0644 & ~new_n24029_;
  assign new_n24039_ = pi0644 & new_n23899_;
  assign new_n24040_ = pi0715 & ~new_n24039_;
  assign new_n24041_ = ~new_n24038_ & new_n24040_;
  assign new_n24042_ = ~pi1160 & ~new_n24041_;
  assign new_n24043_ = ~new_n24037_ & new_n24042_;
  assign new_n24044_ = ~new_n24035_ & ~new_n24043_;
  assign new_n24045_ = pi0790 & ~new_n24044_;
  assign new_n24046_ = pi0644 & new_n24034_;
  assign new_n24047_ = ~pi0644 & new_n24042_;
  assign new_n24048_ = pi0790 & ~new_n24047_;
  assign new_n24049_ = ~new_n24046_ & new_n24048_;
  assign new_n24050_ = ~new_n20567_ & new_n24023_;
  assign new_n24051_ = new_n17760_ & new_n23940_;
  assign new_n24052_ = new_n17759_ & new_n23944_;
  assign new_n24053_ = ~new_n24051_ & ~new_n24052_;
  assign new_n24054_ = ~new_n24050_ & new_n24053_;
  assign new_n24055_ = pi0792 & ~new_n24054_;
  assign new_n24056_ = ~pi0700 & new_n23979_;
  assign new_n24057_ = ~pi0175 & new_n16810_;
  assign new_n24058_ = pi0175 & new_n16928_;
  assign new_n24059_ = ~pi0766 & ~new_n24058_;
  assign new_n24060_ = ~new_n24057_ & new_n24059_;
  assign new_n24061_ = pi0175 & new_n17007_;
  assign new_n24062_ = ~pi0175 & ~new_n17074_;
  assign new_n24063_ = pi0766 & ~new_n24062_;
  assign new_n24064_ = ~new_n24061_ & new_n24063_;
  assign new_n24065_ = pi0039 & ~new_n24064_;
  assign new_n24066_ = ~new_n24060_ & new_n24065_;
  assign new_n24067_ = pi0175 & new_n17178_;
  assign new_n24068_ = ~pi0175 & new_n17217_;
  assign new_n24069_ = ~pi0766 & ~new_n24068_;
  assign new_n24070_ = ~new_n24067_ & new_n24069_;
  assign new_n24071_ = ~pi0175 & ~new_n17227_;
  assign new_n24072_ = pi0175 & ~new_n17234_;
  assign new_n24073_ = pi0766 & ~new_n24072_;
  assign new_n24074_ = ~new_n24071_ & new_n24073_;
  assign new_n24075_ = ~pi0039 & ~new_n24074_;
  assign new_n24076_ = ~new_n24070_ & new_n24075_;
  assign new_n24077_ = ~pi0038 & ~new_n24076_;
  assign new_n24078_ = ~new_n24066_ & new_n24077_;
  assign new_n24079_ = ~new_n16640_ & new_n16647_;
  assign new_n24080_ = ~pi0766 & new_n24079_;
  assign new_n24081_ = ~new_n17035_ & ~new_n24080_;
  assign new_n24082_ = ~pi0039 & ~new_n24081_;
  assign new_n24083_ = ~pi0175 & ~new_n24082_;
  assign new_n24084_ = ~new_n16916_ & ~new_n23712_;
  assign new_n24085_ = pi0175 & ~new_n24084_;
  assign new_n24086_ = new_n6257_ & new_n24085_;
  assign new_n24087_ = pi0038 & ~new_n24086_;
  assign new_n24088_ = ~new_n24083_ & new_n24087_;
  assign new_n24089_ = pi0700 & ~new_n24088_;
  assign new_n24090_ = ~new_n24078_ & new_n24089_;
  assign new_n24091_ = new_n3272_ & ~new_n24090_;
  assign new_n24092_ = ~new_n24056_ & new_n24091_;
  assign new_n24093_ = ~new_n23901_ & ~new_n24092_;
  assign new_n24094_ = ~pi0625 & new_n24093_;
  assign new_n24095_ = pi0625 & new_n23981_;
  assign new_n24096_ = ~pi1153 & ~new_n24095_;
  assign new_n24097_ = ~new_n24094_ & new_n24096_;
  assign new_n24098_ = ~pi0608 & ~new_n23919_;
  assign new_n24099_ = ~new_n24097_ & new_n24098_;
  assign new_n24100_ = pi0625 & new_n24093_;
  assign new_n24101_ = ~pi0625 & new_n23981_;
  assign new_n24102_ = pi1153 & ~new_n24101_;
  assign new_n24103_ = ~new_n24100_ & new_n24102_;
  assign new_n24104_ = pi0608 & ~new_n23923_;
  assign new_n24105_ = ~new_n24103_ & new_n24104_;
  assign new_n24106_ = ~new_n24099_ & ~new_n24105_;
  assign new_n24107_ = pi0778 & ~new_n24106_;
  assign new_n24108_ = ~pi0778 & new_n24093_;
  assign new_n24109_ = ~new_n24107_ & ~new_n24108_;
  assign new_n24110_ = ~pi0609 & ~new_n24109_;
  assign new_n24111_ = pi0609 & new_n23926_;
  assign new_n24112_ = ~pi1155 & ~new_n24111_;
  assign new_n24113_ = ~new_n24110_ & new_n24112_;
  assign new_n24114_ = ~pi0660 & ~new_n23989_;
  assign new_n24115_ = ~new_n24113_ & new_n24114_;
  assign new_n24116_ = pi0609 & ~new_n24109_;
  assign new_n24117_ = ~pi0609 & new_n23926_;
  assign new_n24118_ = pi1155 & ~new_n24117_;
  assign new_n24119_ = ~new_n24116_ & new_n24118_;
  assign new_n24120_ = pi0660 & ~new_n23993_;
  assign new_n24121_ = ~new_n24119_ & new_n24120_;
  assign new_n24122_ = ~new_n24115_ & ~new_n24121_;
  assign new_n24123_ = pi0785 & ~new_n24122_;
  assign new_n24124_ = ~pi0785 & ~new_n24109_;
  assign new_n24125_ = ~new_n24123_ & ~new_n24124_;
  assign new_n24126_ = ~pi0618 & ~new_n24125_;
  assign new_n24127_ = pi0618 & new_n23929_;
  assign new_n24128_ = ~pi1154 & ~new_n24127_;
  assign new_n24129_ = ~new_n24126_ & new_n24128_;
  assign new_n24130_ = ~pi0627 & ~new_n24001_;
  assign new_n24131_ = ~new_n24129_ & new_n24130_;
  assign new_n24132_ = pi0618 & ~new_n24125_;
  assign new_n24133_ = ~pi0618 & new_n23929_;
  assign new_n24134_ = pi1154 & ~new_n24133_;
  assign new_n24135_ = ~new_n24132_ & new_n24134_;
  assign new_n24136_ = pi0627 & ~new_n24005_;
  assign new_n24137_ = ~new_n24135_ & new_n24136_;
  assign new_n24138_ = ~new_n24131_ & ~new_n24137_;
  assign new_n24139_ = pi0781 & ~new_n24138_;
  assign new_n24140_ = ~pi0781 & ~new_n24125_;
  assign new_n24141_ = ~new_n24139_ & ~new_n24140_;
  assign new_n24142_ = pi0619 & ~new_n24141_;
  assign new_n24143_ = ~pi0619 & ~new_n23932_;
  assign new_n24144_ = pi1159 & ~new_n24143_;
  assign new_n24145_ = ~new_n24142_ & new_n24144_;
  assign new_n24146_ = pi0648 & ~new_n24017_;
  assign new_n24147_ = ~new_n24145_ & new_n24146_;
  assign new_n24148_ = ~pi0619 & ~new_n24141_;
  assign new_n24149_ = pi0619 & ~new_n23932_;
  assign new_n24150_ = ~pi1159 & ~new_n24149_;
  assign new_n24151_ = ~new_n24148_ & new_n24150_;
  assign new_n24152_ = ~pi0648 & ~new_n24013_;
  assign new_n24153_ = ~new_n24151_ & new_n24152_;
  assign new_n24154_ = pi0789 & ~new_n24153_;
  assign new_n24155_ = ~new_n24147_ & new_n24154_;
  assign new_n24156_ = ~pi0789 & new_n24141_;
  assign new_n24157_ = new_n17969_ & ~new_n24156_;
  assign new_n24158_ = ~new_n24155_ & new_n24157_;
  assign new_n24159_ = pi0626 & ~new_n24020_;
  assign new_n24160_ = ~pi0626 & ~new_n23899_;
  assign new_n24161_ = new_n17731_ & ~new_n24160_;
  assign new_n24162_ = ~new_n24159_ & new_n24161_;
  assign new_n24163_ = new_n17856_ & new_n23934_;
  assign new_n24164_ = ~pi0626 & ~new_n24020_;
  assign new_n24165_ = pi0626 & ~new_n23899_;
  assign new_n24166_ = new_n17732_ & ~new_n24165_;
  assign new_n24167_ = ~new_n24164_ & new_n24166_;
  assign new_n24168_ = ~new_n24163_ & ~new_n24167_;
  assign new_n24169_ = ~new_n24162_ & new_n24168_;
  assign new_n24170_ = pi0788 & ~new_n24169_;
  assign new_n24171_ = ~new_n20364_ & ~new_n24170_;
  assign new_n24172_ = ~new_n24158_ & new_n24171_;
  assign new_n24173_ = ~new_n24055_ & ~new_n24172_;
  assign new_n24174_ = ~new_n20360_ & ~new_n24173_;
  assign new_n24175_ = new_n17801_ & new_n23956_;
  assign new_n24176_ = new_n17802_ & new_n23952_;
  assign new_n24177_ = ~new_n20556_ & new_n24026_;
  assign new_n24178_ = ~new_n24176_ & ~new_n24177_;
  assign new_n24179_ = ~new_n24175_ & new_n24178_;
  assign new_n24180_ = pi0787 & ~new_n24179_;
  assign new_n24181_ = ~new_n24174_ & ~new_n24180_;
  assign new_n24182_ = ~new_n24049_ & new_n24181_;
  assign new_n24183_ = ~new_n24045_ & ~new_n24182_;
  assign new_n24184_ = ~po1038 & ~new_n24183_;
  assign new_n24185_ = ~pi0175 & po1038;
  assign new_n24186_ = ~pi0832 & ~new_n24185_;
  assign new_n24187_ = ~new_n24184_ & new_n24186_;
  assign po0332 = ~new_n23898_ & ~new_n24187_;
  assign new_n24189_ = ~pi0176 & ~new_n2754_;
  assign new_n24190_ = ~pi0742 & new_n16913_;
  assign new_n24191_ = ~new_n24189_ & ~new_n24190_;
  assign new_n24192_ = ~new_n17858_ & ~new_n24191_;
  assign new_n24193_ = ~pi0785 & ~new_n24192_;
  assign new_n24194_ = ~new_n17863_ & ~new_n24191_;
  assign new_n24195_ = pi1155 & ~new_n24194_;
  assign new_n24196_ = ~new_n17866_ & new_n24192_;
  assign new_n24197_ = ~pi1155 & ~new_n24196_;
  assign new_n24198_ = ~new_n24195_ & ~new_n24197_;
  assign new_n24199_ = pi0785 & ~new_n24198_;
  assign new_n24200_ = ~new_n24193_ & ~new_n24199_;
  assign new_n24201_ = ~pi0781 & ~new_n24200_;
  assign new_n24202_ = ~new_n17873_ & new_n24200_;
  assign new_n24203_ = pi1154 & ~new_n24202_;
  assign new_n24204_ = ~new_n17876_ & new_n24200_;
  assign new_n24205_ = ~pi1154 & ~new_n24204_;
  assign new_n24206_ = ~new_n24203_ & ~new_n24205_;
  assign new_n24207_ = pi0781 & ~new_n24206_;
  assign new_n24208_ = ~new_n24201_ & ~new_n24207_;
  assign new_n24209_ = ~pi0789 & ~new_n24208_;
  assign new_n24210_ = pi0619 & new_n24208_;
  assign new_n24211_ = ~pi0619 & new_n24189_;
  assign new_n24212_ = pi1159 & ~new_n24211_;
  assign new_n24213_ = ~new_n24210_ & new_n24212_;
  assign new_n24214_ = ~pi0619 & new_n24208_;
  assign new_n24215_ = pi0619 & new_n24189_;
  assign new_n24216_ = ~pi1159 & ~new_n24215_;
  assign new_n24217_ = ~new_n24214_ & new_n24216_;
  assign new_n24218_ = ~new_n24213_ & ~new_n24217_;
  assign new_n24219_ = pi0789 & ~new_n24218_;
  assign new_n24220_ = ~new_n24209_ & ~new_n24219_;
  assign new_n24221_ = ~new_n17968_ & new_n24220_;
  assign new_n24222_ = new_n17968_ & new_n24189_;
  assign new_n24223_ = ~new_n24221_ & ~new_n24222_;
  assign new_n24224_ = ~new_n17762_ & ~new_n24223_;
  assign new_n24225_ = new_n17762_ & new_n24189_;
  assign new_n24226_ = ~new_n24224_ & ~new_n24225_;
  assign new_n24227_ = ~new_n20556_ & new_n24226_;
  assign new_n24228_ = ~pi0704 & new_n16915_;
  assign new_n24229_ = ~new_n24189_ & ~new_n24228_;
  assign new_n24230_ = ~pi0778 & new_n24229_;
  assign new_n24231_ = ~pi0625 & new_n24228_;
  assign new_n24232_ = ~new_n24229_ & ~new_n24231_;
  assign new_n24233_ = pi1153 & ~new_n24232_;
  assign new_n24234_ = ~pi1153 & ~new_n24189_;
  assign new_n24235_ = ~new_n24231_ & new_n24234_;
  assign new_n24236_ = ~new_n24233_ & ~new_n24235_;
  assign new_n24237_ = pi0778 & ~new_n24236_;
  assign new_n24238_ = ~new_n24230_ & ~new_n24237_;
  assign new_n24239_ = ~new_n17844_ & new_n24238_;
  assign new_n24240_ = ~new_n17846_ & new_n24239_;
  assign new_n24241_ = ~new_n17848_ & new_n24240_;
  assign new_n24242_ = ~new_n17980_ & new_n24241_;
  assign new_n24243_ = ~new_n18011_ & new_n24242_;
  assign new_n24244_ = ~pi0647 & new_n24243_;
  assign new_n24245_ = pi0647 & new_n24189_;
  assign new_n24246_ = ~pi1157 & ~new_n24245_;
  assign new_n24247_ = ~new_n24244_ & new_n24246_;
  assign new_n24248_ = pi0630 & new_n24247_;
  assign new_n24249_ = pi0647 & ~new_n24243_;
  assign new_n24250_ = ~pi0647 & ~new_n24189_;
  assign new_n24251_ = ~new_n24249_ & ~new_n24250_;
  assign new_n24252_ = new_n17801_ & ~new_n24251_;
  assign new_n24253_ = ~new_n24248_ & ~new_n24252_;
  assign new_n24254_ = ~new_n24227_ & new_n24253_;
  assign new_n24255_ = pi0787 & ~new_n24254_;
  assign new_n24256_ = pi0626 & ~new_n24220_;
  assign new_n24257_ = ~pi0626 & ~new_n24189_;
  assign new_n24258_ = new_n17731_ & ~new_n24257_;
  assign new_n24259_ = ~new_n24256_ & new_n24258_;
  assign new_n24260_ = new_n17856_ & new_n24241_;
  assign new_n24261_ = ~pi0626 & ~new_n24220_;
  assign new_n24262_ = pi0626 & ~new_n24189_;
  assign new_n24263_ = new_n17732_ & ~new_n24262_;
  assign new_n24264_ = ~new_n24261_ & new_n24263_;
  assign new_n24265_ = ~new_n24260_ & ~new_n24264_;
  assign new_n24266_ = ~new_n24259_ & new_n24265_;
  assign new_n24267_ = pi0788 & ~new_n24266_;
  assign new_n24268_ = ~new_n16639_ & ~new_n24229_;
  assign new_n24269_ = pi0625 & new_n24268_;
  assign new_n24270_ = new_n24191_ & ~new_n24268_;
  assign new_n24271_ = ~new_n24269_ & ~new_n24270_;
  assign new_n24272_ = new_n24234_ & ~new_n24271_;
  assign new_n24273_ = ~pi0608 & ~new_n24233_;
  assign new_n24274_ = ~new_n24272_ & new_n24273_;
  assign new_n24275_ = pi1153 & new_n24191_;
  assign new_n24276_ = ~new_n24269_ & new_n24275_;
  assign new_n24277_ = pi0608 & ~new_n24235_;
  assign new_n24278_ = ~new_n24276_ & new_n24277_;
  assign new_n24279_ = ~new_n24274_ & ~new_n24278_;
  assign new_n24280_ = pi0778 & ~new_n24279_;
  assign new_n24281_ = ~pi0778 & ~new_n24270_;
  assign new_n24282_ = ~new_n24280_ & ~new_n24281_;
  assign new_n24283_ = ~pi0609 & ~new_n24282_;
  assign new_n24284_ = pi0609 & new_n24238_;
  assign new_n24285_ = ~pi1155 & ~new_n24284_;
  assign new_n24286_ = ~new_n24283_ & new_n24285_;
  assign new_n24287_ = ~pi0660 & ~new_n24195_;
  assign new_n24288_ = ~new_n24286_ & new_n24287_;
  assign new_n24289_ = pi0609 & ~new_n24282_;
  assign new_n24290_ = ~pi0609 & new_n24238_;
  assign new_n24291_ = pi1155 & ~new_n24290_;
  assign new_n24292_ = ~new_n24289_ & new_n24291_;
  assign new_n24293_ = pi0660 & ~new_n24197_;
  assign new_n24294_ = ~new_n24292_ & new_n24293_;
  assign new_n24295_ = ~new_n24288_ & ~new_n24294_;
  assign new_n24296_ = pi0785 & ~new_n24295_;
  assign new_n24297_ = ~pi0785 & ~new_n24282_;
  assign new_n24298_ = ~new_n24296_ & ~new_n24297_;
  assign new_n24299_ = ~pi0618 & ~new_n24298_;
  assign new_n24300_ = pi0618 & new_n24239_;
  assign new_n24301_ = ~pi1154 & ~new_n24300_;
  assign new_n24302_ = ~new_n24299_ & new_n24301_;
  assign new_n24303_ = ~pi0627 & ~new_n24203_;
  assign new_n24304_ = ~new_n24302_ & new_n24303_;
  assign new_n24305_ = pi0618 & ~new_n24298_;
  assign new_n24306_ = ~pi0618 & new_n24239_;
  assign new_n24307_ = pi1154 & ~new_n24306_;
  assign new_n24308_ = ~new_n24305_ & new_n24307_;
  assign new_n24309_ = pi0627 & ~new_n24205_;
  assign new_n24310_ = ~new_n24308_ & new_n24309_;
  assign new_n24311_ = ~new_n24304_ & ~new_n24310_;
  assign new_n24312_ = pi0781 & ~new_n24311_;
  assign new_n24313_ = ~pi0781 & ~new_n24298_;
  assign new_n24314_ = ~new_n24312_ & ~new_n24313_;
  assign new_n24315_ = pi0619 & ~new_n24314_;
  assign new_n24316_ = ~pi0619 & new_n24240_;
  assign new_n24317_ = pi1159 & ~new_n24316_;
  assign new_n24318_ = ~new_n24315_ & new_n24317_;
  assign new_n24319_ = pi0648 & ~new_n24217_;
  assign new_n24320_ = ~new_n24318_ & new_n24319_;
  assign new_n24321_ = ~pi0619 & ~new_n24314_;
  assign new_n24322_ = pi0619 & new_n24240_;
  assign new_n24323_ = ~pi1159 & ~new_n24322_;
  assign new_n24324_ = ~new_n24321_ & new_n24323_;
  assign new_n24325_ = ~pi0648 & ~new_n24213_;
  assign new_n24326_ = ~new_n24324_ & new_n24325_;
  assign new_n24327_ = pi0789 & ~new_n24326_;
  assign new_n24328_ = ~new_n24320_ & new_n24327_;
  assign new_n24329_ = ~pi0789 & new_n24314_;
  assign new_n24330_ = new_n17969_ & ~new_n24329_;
  assign new_n24331_ = ~new_n24328_ & new_n24330_;
  assign new_n24332_ = ~new_n24267_ & ~new_n24331_;
  assign new_n24333_ = ~new_n20364_ & ~new_n24332_;
  assign new_n24334_ = new_n18008_ & ~new_n24223_;
  assign new_n24335_ = new_n20851_ & new_n24242_;
  assign new_n24336_ = ~new_n24334_ & ~new_n24335_;
  assign new_n24337_ = ~pi0629 & ~new_n24336_;
  assign new_n24338_ = new_n20855_ & new_n24242_;
  assign new_n24339_ = new_n18007_ & ~new_n24223_;
  assign new_n24340_ = ~new_n24338_ & ~new_n24339_;
  assign new_n24341_ = pi0629 & ~new_n24340_;
  assign new_n24342_ = ~new_n24337_ & ~new_n24341_;
  assign new_n24343_ = pi0792 & ~new_n24342_;
  assign new_n24344_ = ~new_n20360_ & ~new_n24343_;
  assign new_n24345_ = ~new_n24333_ & new_n24344_;
  assign new_n24346_ = ~new_n24255_ & ~new_n24345_;
  assign new_n24347_ = pi0644 & new_n24346_;
  assign new_n24348_ = ~pi0787 & ~new_n24243_;
  assign new_n24349_ = pi1157 & ~new_n24251_;
  assign new_n24350_ = ~new_n24247_ & ~new_n24349_;
  assign new_n24351_ = pi0787 & ~new_n24350_;
  assign new_n24352_ = ~new_n24348_ & ~new_n24351_;
  assign new_n24353_ = ~pi0644 & new_n24352_;
  assign new_n24354_ = pi0715 & ~new_n24353_;
  assign new_n24355_ = ~new_n24347_ & new_n24354_;
  assign new_n24356_ = ~new_n17804_ & ~new_n24226_;
  assign new_n24357_ = new_n17804_ & new_n24189_;
  assign new_n24358_ = ~new_n24356_ & ~new_n24357_;
  assign new_n24359_ = pi0644 & ~new_n24358_;
  assign new_n24360_ = ~pi0644 & new_n24189_;
  assign new_n24361_ = ~pi0715 & ~new_n24360_;
  assign new_n24362_ = ~new_n24359_ & new_n24361_;
  assign new_n24363_ = pi1160 & ~new_n24362_;
  assign new_n24364_ = ~new_n24355_ & new_n24363_;
  assign new_n24365_ = ~pi0644 & new_n24346_;
  assign new_n24366_ = pi0644 & new_n24352_;
  assign new_n24367_ = ~pi0715 & ~new_n24366_;
  assign new_n24368_ = ~new_n24365_ & new_n24367_;
  assign new_n24369_ = ~pi0644 & ~new_n24358_;
  assign new_n24370_ = pi0644 & new_n24189_;
  assign new_n24371_ = pi0715 & ~new_n24370_;
  assign new_n24372_ = ~new_n24369_ & new_n24371_;
  assign new_n24373_ = ~pi1160 & ~new_n24372_;
  assign new_n24374_ = ~new_n24368_ & new_n24373_;
  assign new_n24375_ = ~new_n24364_ & ~new_n24374_;
  assign new_n24376_ = pi0790 & ~new_n24375_;
  assign new_n24377_ = ~pi0790 & new_n24346_;
  assign new_n24378_ = pi0832 & ~new_n24377_;
  assign new_n24379_ = ~new_n24376_ & new_n24378_;
  assign new_n24380_ = ~pi0176 & ~new_n17558_;
  assign new_n24381_ = new_n17691_ & ~new_n24380_;
  assign new_n24382_ = ~pi0038 & new_n18128_;
  assign new_n24383_ = new_n3272_ & ~new_n17544_;
  assign new_n24384_ = ~new_n24382_ & new_n24383_;
  assign new_n24385_ = pi0176 & ~new_n24384_;
  assign new_n24386_ = ~pi0038 & new_n18124_;
  assign new_n24387_ = ~new_n19956_ & ~new_n24386_;
  assign new_n24388_ = ~pi0176 & new_n24387_;
  assign new_n24389_ = ~pi0704 & ~new_n24388_;
  assign new_n24390_ = ~pi0176 & ~new_n17551_;
  assign new_n24391_ = pi0704 & new_n24390_;
  assign new_n24392_ = new_n3272_ & ~new_n24391_;
  assign new_n24393_ = ~new_n24389_ & new_n24392_;
  assign new_n24394_ = ~new_n24385_ & ~new_n24393_;
  assign new_n24395_ = ~pi0778 & ~new_n24394_;
  assign new_n24396_ = pi0625 & new_n24394_;
  assign new_n24397_ = ~pi0625 & new_n24380_;
  assign new_n24398_ = pi1153 & ~new_n24397_;
  assign new_n24399_ = ~new_n24396_ & new_n24398_;
  assign new_n24400_ = ~pi0625 & new_n24394_;
  assign new_n24401_ = pi0625 & new_n24380_;
  assign new_n24402_ = ~pi1153 & ~new_n24401_;
  assign new_n24403_ = ~new_n24400_ & new_n24402_;
  assign new_n24404_ = ~new_n24399_ & ~new_n24403_;
  assign new_n24405_ = pi0778 & ~new_n24404_;
  assign new_n24406_ = ~new_n24395_ & ~new_n24405_;
  assign new_n24407_ = ~new_n17618_ & ~new_n24406_;
  assign new_n24408_ = new_n17618_ & ~new_n24380_;
  assign new_n24409_ = ~new_n24407_ & ~new_n24408_;
  assign new_n24410_ = ~new_n17655_ & new_n24409_;
  assign new_n24411_ = new_n17655_ & new_n24380_;
  assign new_n24412_ = ~new_n24410_ & ~new_n24411_;
  assign new_n24413_ = ~new_n17691_ & new_n24412_;
  assign new_n24414_ = ~new_n24381_ & ~new_n24413_;
  assign new_n24415_ = ~new_n17734_ & new_n24414_;
  assign new_n24416_ = new_n17734_ & new_n24380_;
  assign new_n24417_ = ~new_n24415_ & ~new_n24416_;
  assign new_n24418_ = ~pi0628 & ~new_n24417_;
  assign new_n24419_ = pi0628 & new_n24380_;
  assign new_n24420_ = ~new_n24418_ & ~new_n24419_;
  assign new_n24421_ = ~pi1156 & ~new_n24420_;
  assign new_n24422_ = pi0628 & ~new_n24417_;
  assign new_n24423_ = ~pi0628 & new_n24380_;
  assign new_n24424_ = ~new_n24422_ & ~new_n24423_;
  assign new_n24425_ = pi1156 & ~new_n24424_;
  assign new_n24426_ = ~new_n24421_ & ~new_n24425_;
  assign new_n24427_ = pi0792 & ~new_n24426_;
  assign new_n24428_ = ~pi0792 & ~new_n24417_;
  assign new_n24429_ = ~new_n24427_ & ~new_n24428_;
  assign new_n24430_ = ~pi0647 & ~new_n24429_;
  assign new_n24431_ = pi0647 & new_n24380_;
  assign new_n24432_ = ~new_n24430_ & ~new_n24431_;
  assign new_n24433_ = ~pi1157 & ~new_n24432_;
  assign new_n24434_ = pi0647 & ~new_n24429_;
  assign new_n24435_ = ~pi0647 & new_n24380_;
  assign new_n24436_ = ~new_n24434_ & ~new_n24435_;
  assign new_n24437_ = pi1157 & ~new_n24436_;
  assign new_n24438_ = ~new_n24433_ & ~new_n24437_;
  assign new_n24439_ = pi0787 & ~new_n24438_;
  assign new_n24440_ = ~pi0787 & ~new_n24429_;
  assign new_n24441_ = ~new_n24439_ & ~new_n24440_;
  assign new_n24442_ = ~pi0644 & ~new_n24441_;
  assign new_n24443_ = pi0715 & ~new_n24442_;
  assign new_n24444_ = pi0176 & ~new_n3272_;
  assign new_n24445_ = ~pi0176 & new_n19376_;
  assign new_n24446_ = ~new_n19370_ & ~new_n19371_;
  assign new_n24447_ = pi0176 & new_n24446_;
  assign new_n24448_ = ~new_n24445_ & ~new_n24447_;
  assign new_n24449_ = ~pi0742 & ~new_n24448_;
  assign new_n24450_ = pi0742 & ~new_n24390_;
  assign new_n24451_ = ~new_n24449_ & ~new_n24450_;
  assign new_n24452_ = new_n3272_ & ~new_n24451_;
  assign new_n24453_ = ~new_n24444_ & ~new_n24452_;
  assign new_n24454_ = ~new_n17590_ & ~new_n24453_;
  assign new_n24455_ = new_n17590_ & ~new_n24380_;
  assign new_n24456_ = ~new_n24454_ & ~new_n24455_;
  assign new_n24457_ = ~pi0785 & ~new_n24456_;
  assign new_n24458_ = ~new_n17591_ & ~new_n24380_;
  assign new_n24459_ = pi0609 & new_n24454_;
  assign new_n24460_ = ~new_n24458_ & ~new_n24459_;
  assign new_n24461_ = pi1155 & ~new_n24460_;
  assign new_n24462_ = ~new_n17603_ & ~new_n24380_;
  assign new_n24463_ = ~pi0609 & new_n24454_;
  assign new_n24464_ = ~new_n24462_ & ~new_n24463_;
  assign new_n24465_ = ~pi1155 & ~new_n24464_;
  assign new_n24466_ = ~new_n24461_ & ~new_n24465_;
  assign new_n24467_ = pi0785 & ~new_n24466_;
  assign new_n24468_ = ~new_n24457_ & ~new_n24467_;
  assign new_n24469_ = ~pi0781 & ~new_n24468_;
  assign new_n24470_ = pi0618 & new_n24468_;
  assign new_n24471_ = ~pi0618 & new_n24380_;
  assign new_n24472_ = pi1154 & ~new_n24471_;
  assign new_n24473_ = ~new_n24470_ & new_n24472_;
  assign new_n24474_ = ~pi0618 & new_n24468_;
  assign new_n24475_ = pi0618 & new_n24380_;
  assign new_n24476_ = ~pi1154 & ~new_n24475_;
  assign new_n24477_ = ~new_n24474_ & new_n24476_;
  assign new_n24478_ = ~new_n24473_ & ~new_n24477_;
  assign new_n24479_ = pi0781 & ~new_n24478_;
  assign new_n24480_ = ~new_n24469_ & ~new_n24479_;
  assign new_n24481_ = ~pi0789 & ~new_n24480_;
  assign new_n24482_ = pi0619 & new_n24480_;
  assign new_n24483_ = ~pi0619 & new_n24380_;
  assign new_n24484_ = pi1159 & ~new_n24483_;
  assign new_n24485_ = ~new_n24482_ & new_n24484_;
  assign new_n24486_ = ~pi0619 & new_n24480_;
  assign new_n24487_ = pi0619 & new_n24380_;
  assign new_n24488_ = ~pi1159 & ~new_n24487_;
  assign new_n24489_ = ~new_n24486_ & new_n24488_;
  assign new_n24490_ = ~new_n24485_ & ~new_n24489_;
  assign new_n24491_ = pi0789 & ~new_n24490_;
  assign new_n24492_ = ~new_n24481_ & ~new_n24491_;
  assign new_n24493_ = ~new_n17968_ & new_n24492_;
  assign new_n24494_ = new_n17968_ & new_n24380_;
  assign new_n24495_ = ~new_n24493_ & ~new_n24494_;
  assign new_n24496_ = ~new_n17762_ & ~new_n24495_;
  assign new_n24497_ = new_n17762_ & new_n24380_;
  assign new_n24498_ = ~new_n24496_ & ~new_n24497_;
  assign new_n24499_ = ~new_n17804_ & ~new_n24498_;
  assign new_n24500_ = new_n17804_ & new_n24380_;
  assign new_n24501_ = ~new_n24499_ & ~new_n24500_;
  assign new_n24502_ = pi0644 & ~new_n24501_;
  assign new_n24503_ = ~pi0644 & new_n24380_;
  assign new_n24504_ = ~pi0715 & ~new_n24503_;
  assign new_n24505_ = ~new_n24502_ & new_n24504_;
  assign new_n24506_ = pi1160 & ~new_n24505_;
  assign new_n24507_ = ~new_n24443_ & new_n24506_;
  assign new_n24508_ = pi0644 & ~new_n24441_;
  assign new_n24509_ = ~pi0715 & ~new_n24508_;
  assign new_n24510_ = ~pi0644 & ~new_n24501_;
  assign new_n24511_ = pi0644 & new_n24380_;
  assign new_n24512_ = pi0715 & ~new_n24511_;
  assign new_n24513_ = ~new_n24510_ & new_n24512_;
  assign new_n24514_ = ~pi1160 & ~new_n24513_;
  assign new_n24515_ = ~new_n24509_ & new_n24514_;
  assign new_n24516_ = ~new_n24507_ & ~new_n24515_;
  assign new_n24517_ = pi0790 & ~new_n24516_;
  assign new_n24518_ = pi0644 & new_n24506_;
  assign new_n24519_ = ~pi0644 & new_n24514_;
  assign new_n24520_ = pi0790 & ~new_n24519_;
  assign new_n24521_ = ~new_n24518_ & new_n24520_;
  assign new_n24522_ = new_n17801_ & new_n24436_;
  assign new_n24523_ = new_n17802_ & new_n24432_;
  assign new_n24524_ = ~new_n20556_ & new_n24498_;
  assign new_n24525_ = ~new_n24523_ & ~new_n24524_;
  assign new_n24526_ = ~new_n24522_ & new_n24525_;
  assign new_n24527_ = pi0787 & ~new_n24526_;
  assign new_n24528_ = ~new_n20567_ & new_n24495_;
  assign new_n24529_ = new_n17760_ & new_n24420_;
  assign new_n24530_ = new_n17759_ & new_n24424_;
  assign new_n24531_ = ~new_n24529_ & ~new_n24530_;
  assign new_n24532_ = ~new_n24528_ & new_n24531_;
  assign new_n24533_ = pi0792 & ~new_n24532_;
  assign new_n24534_ = pi0626 & ~new_n24492_;
  assign new_n24535_ = ~pi0626 & ~new_n24380_;
  assign new_n24536_ = new_n17731_ & ~new_n24535_;
  assign new_n24537_ = ~new_n24534_ & new_n24536_;
  assign new_n24538_ = new_n17856_ & new_n24414_;
  assign new_n24539_ = ~pi0626 & ~new_n24492_;
  assign new_n24540_ = pi0626 & ~new_n24380_;
  assign new_n24541_ = new_n17732_ & ~new_n24540_;
  assign new_n24542_ = ~new_n24539_ & new_n24541_;
  assign new_n24543_ = ~new_n24538_ & ~new_n24542_;
  assign new_n24544_ = ~new_n24537_ & new_n24543_;
  assign new_n24545_ = pi0788 & ~new_n24544_;
  assign new_n24546_ = pi0704 & new_n24451_;
  assign new_n24547_ = ~pi0176 & new_n19389_;
  assign new_n24548_ = ~new_n19394_ & ~new_n19396_;
  assign new_n24549_ = pi0176 & ~new_n24548_;
  assign new_n24550_ = pi0742 & ~new_n24549_;
  assign new_n24551_ = ~new_n24547_ & new_n24550_;
  assign new_n24552_ = pi0176 & new_n19406_;
  assign new_n24553_ = ~pi0176 & ~new_n19414_;
  assign new_n24554_ = ~pi0742 & ~new_n24553_;
  assign new_n24555_ = ~new_n24552_ & new_n24554_;
  assign new_n24556_ = ~pi0704 & ~new_n24555_;
  assign new_n24557_ = ~new_n24551_ & new_n24556_;
  assign new_n24558_ = new_n3272_ & ~new_n24557_;
  assign new_n24559_ = ~new_n24546_ & new_n24558_;
  assign new_n24560_ = ~new_n24444_ & ~new_n24559_;
  assign new_n24561_ = ~pi0625 & new_n24560_;
  assign new_n24562_ = pi0625 & new_n24453_;
  assign new_n24563_ = ~pi1153 & ~new_n24562_;
  assign new_n24564_ = ~new_n24561_ & new_n24563_;
  assign new_n24565_ = ~pi0608 & ~new_n24399_;
  assign new_n24566_ = ~new_n24564_ & new_n24565_;
  assign new_n24567_ = pi0625 & new_n24560_;
  assign new_n24568_ = ~pi0625 & new_n24453_;
  assign new_n24569_ = pi1153 & ~new_n24568_;
  assign new_n24570_ = ~new_n24567_ & new_n24569_;
  assign new_n24571_ = pi0608 & ~new_n24403_;
  assign new_n24572_ = ~new_n24570_ & new_n24571_;
  assign new_n24573_ = ~new_n24566_ & ~new_n24572_;
  assign new_n24574_ = pi0778 & ~new_n24573_;
  assign new_n24575_ = ~pi0778 & new_n24560_;
  assign new_n24576_ = ~new_n24574_ & ~new_n24575_;
  assign new_n24577_ = ~pi0609 & ~new_n24576_;
  assign new_n24578_ = pi0609 & new_n24406_;
  assign new_n24579_ = ~pi1155 & ~new_n24578_;
  assign new_n24580_ = ~new_n24577_ & new_n24579_;
  assign new_n24581_ = ~pi0660 & ~new_n24461_;
  assign new_n24582_ = ~new_n24580_ & new_n24581_;
  assign new_n24583_ = pi0609 & ~new_n24576_;
  assign new_n24584_ = ~pi0609 & new_n24406_;
  assign new_n24585_ = pi1155 & ~new_n24584_;
  assign new_n24586_ = ~new_n24583_ & new_n24585_;
  assign new_n24587_ = pi0660 & ~new_n24465_;
  assign new_n24588_ = ~new_n24586_ & new_n24587_;
  assign new_n24589_ = ~new_n24582_ & ~new_n24588_;
  assign new_n24590_ = pi0785 & ~new_n24589_;
  assign new_n24591_ = ~pi0785 & ~new_n24576_;
  assign new_n24592_ = ~new_n24590_ & ~new_n24591_;
  assign new_n24593_ = ~pi0618 & ~new_n24592_;
  assign new_n24594_ = pi0618 & new_n24409_;
  assign new_n24595_ = ~pi1154 & ~new_n24594_;
  assign new_n24596_ = ~new_n24593_ & new_n24595_;
  assign new_n24597_ = ~pi0627 & ~new_n24473_;
  assign new_n24598_ = ~new_n24596_ & new_n24597_;
  assign new_n24599_ = pi0618 & ~new_n24592_;
  assign new_n24600_ = ~pi0618 & new_n24409_;
  assign new_n24601_ = pi1154 & ~new_n24600_;
  assign new_n24602_ = ~new_n24599_ & new_n24601_;
  assign new_n24603_ = pi0627 & ~new_n24477_;
  assign new_n24604_ = ~new_n24602_ & new_n24603_;
  assign new_n24605_ = ~new_n24598_ & ~new_n24604_;
  assign new_n24606_ = pi0781 & ~new_n24605_;
  assign new_n24607_ = ~pi0781 & ~new_n24592_;
  assign new_n24608_ = ~new_n24606_ & ~new_n24607_;
  assign new_n24609_ = pi0619 & ~new_n24608_;
  assign new_n24610_ = ~pi0619 & ~new_n24412_;
  assign new_n24611_ = pi1159 & ~new_n24610_;
  assign new_n24612_ = ~new_n24609_ & new_n24611_;
  assign new_n24613_ = pi0648 & ~new_n24489_;
  assign new_n24614_ = ~new_n24612_ & new_n24613_;
  assign new_n24615_ = ~pi0619 & ~new_n24608_;
  assign new_n24616_ = pi0619 & ~new_n24412_;
  assign new_n24617_ = ~pi1159 & ~new_n24616_;
  assign new_n24618_ = ~new_n24615_ & new_n24617_;
  assign new_n24619_ = ~pi0648 & ~new_n24485_;
  assign new_n24620_ = ~new_n24618_ & new_n24619_;
  assign new_n24621_ = pi0789 & ~new_n24620_;
  assign new_n24622_ = ~new_n24614_ & new_n24621_;
  assign new_n24623_ = ~pi0789 & new_n24608_;
  assign new_n24624_ = new_n17969_ & ~new_n24623_;
  assign new_n24625_ = ~new_n24622_ & new_n24624_;
  assign new_n24626_ = ~new_n24545_ & ~new_n24625_;
  assign new_n24627_ = ~new_n24533_ & ~new_n24626_;
  assign new_n24628_ = new_n20364_ & new_n24532_;
  assign new_n24629_ = ~new_n20360_ & ~new_n24628_;
  assign new_n24630_ = ~new_n24627_ & new_n24629_;
  assign new_n24631_ = ~new_n24527_ & ~new_n24630_;
  assign new_n24632_ = ~new_n24521_ & new_n24631_;
  assign new_n24633_ = ~new_n24517_ & ~new_n24632_;
  assign new_n24634_ = ~po1038 & ~new_n24633_;
  assign new_n24635_ = ~pi0176 & po1038;
  assign new_n24636_ = ~pi0832 & ~new_n24635_;
  assign new_n24637_ = ~new_n24634_ & new_n24636_;
  assign po0333 = ~new_n24379_ & ~new_n24637_;
  assign new_n24639_ = pi0177 & ~new_n3272_;
  assign new_n24640_ = ~pi0757 & ~new_n19376_;
  assign new_n24641_ = ~new_n21646_ & ~new_n24640_;
  assign new_n24642_ = ~pi0177 & ~new_n24641_;
  assign new_n24643_ = ~pi0177 & ~new_n19370_;
  assign new_n24644_ = ~pi0757 & ~new_n24643_;
  assign new_n24645_ = ~new_n24446_ & new_n24644_;
  assign new_n24646_ = ~new_n24642_ & ~new_n24645_;
  assign new_n24647_ = pi0686 & ~new_n24646_;
  assign new_n24648_ = ~pi0177 & new_n19387_;
  assign new_n24649_ = pi0177 & new_n19393_;
  assign new_n24650_ = ~pi0038 & ~new_n24649_;
  assign new_n24651_ = ~new_n24648_ & new_n24650_;
  assign new_n24652_ = ~pi0177 & ~new_n17431_;
  assign new_n24653_ = new_n18093_ & ~new_n24652_;
  assign new_n24654_ = pi0757 & ~new_n24653_;
  assign new_n24655_ = ~new_n24651_ & new_n24654_;
  assign new_n24656_ = pi0177 & new_n19404_;
  assign new_n24657_ = ~new_n19408_ & ~new_n19409_;
  assign new_n24658_ = ~pi0177 & ~new_n24657_;
  assign new_n24659_ = ~pi0038 & ~new_n24658_;
  assign new_n24660_ = ~new_n24656_ & new_n24659_;
  assign new_n24661_ = ~pi0177 & ~new_n19411_;
  assign new_n24662_ = pi0177 & new_n19400_;
  assign new_n24663_ = pi0038 & ~new_n24662_;
  assign new_n24664_ = ~new_n24661_ & new_n24663_;
  assign new_n24665_ = ~pi0757 & ~new_n24664_;
  assign new_n24666_ = ~new_n24660_ & new_n24665_;
  assign new_n24667_ = ~new_n24655_ & ~new_n24666_;
  assign new_n24668_ = ~pi0686 & ~new_n24667_;
  assign new_n24669_ = new_n3272_ & ~new_n24668_;
  assign new_n24670_ = ~new_n24647_ & new_n24669_;
  assign new_n24671_ = ~new_n24639_ & ~new_n24670_;
  assign new_n24672_ = ~pi0625 & new_n24671_;
  assign new_n24673_ = new_n3272_ & new_n24646_;
  assign new_n24674_ = ~new_n24639_ & ~new_n24673_;
  assign new_n24675_ = pi0625 & new_n24674_;
  assign new_n24676_ = ~pi1153 & ~new_n24675_;
  assign new_n24677_ = ~new_n24672_ & new_n24676_;
  assign new_n24678_ = ~pi0177 & new_n18124_;
  assign new_n24679_ = pi0177 & ~new_n18128_;
  assign new_n24680_ = ~pi0038 & ~new_n24679_;
  assign new_n24681_ = ~new_n24678_ & new_n24680_;
  assign new_n24682_ = new_n17544_ & ~new_n24652_;
  assign new_n24683_ = ~pi0686 & ~new_n24682_;
  assign new_n24684_ = ~new_n24681_ & new_n24683_;
  assign new_n24685_ = ~pi0177 & pi0686;
  assign new_n24686_ = ~new_n17551_ & new_n24685_;
  assign new_n24687_ = new_n3272_ & ~new_n24686_;
  assign new_n24688_ = ~new_n24684_ & new_n24687_;
  assign new_n24689_ = ~new_n24639_ & ~new_n24688_;
  assign new_n24690_ = pi0625 & new_n24689_;
  assign new_n24691_ = ~pi0177 & ~new_n17558_;
  assign new_n24692_ = ~pi0625 & new_n24691_;
  assign new_n24693_ = pi1153 & ~new_n24692_;
  assign new_n24694_ = ~new_n24690_ & new_n24693_;
  assign new_n24695_ = ~pi0608 & ~new_n24694_;
  assign new_n24696_ = ~new_n24677_ & new_n24695_;
  assign new_n24697_ = pi0625 & new_n24671_;
  assign new_n24698_ = ~pi0625 & new_n24674_;
  assign new_n24699_ = pi1153 & ~new_n24698_;
  assign new_n24700_ = ~new_n24697_ & new_n24699_;
  assign new_n24701_ = ~pi0625 & new_n24689_;
  assign new_n24702_ = pi0625 & new_n24691_;
  assign new_n24703_ = ~pi1153 & ~new_n24702_;
  assign new_n24704_ = ~new_n24701_ & new_n24703_;
  assign new_n24705_ = pi0608 & ~new_n24704_;
  assign new_n24706_ = ~new_n24700_ & new_n24705_;
  assign new_n24707_ = ~new_n24696_ & ~new_n24706_;
  assign new_n24708_ = pi0778 & ~new_n24707_;
  assign new_n24709_ = ~pi0778 & new_n24671_;
  assign new_n24710_ = ~new_n24708_ & ~new_n24709_;
  assign new_n24711_ = ~pi0609 & ~new_n24710_;
  assign new_n24712_ = ~pi0778 & ~new_n24689_;
  assign new_n24713_ = ~new_n24694_ & ~new_n24704_;
  assign new_n24714_ = pi0778 & ~new_n24713_;
  assign new_n24715_ = ~new_n24712_ & ~new_n24714_;
  assign new_n24716_ = pi0609 & new_n24715_;
  assign new_n24717_ = ~pi1155 & ~new_n24716_;
  assign new_n24718_ = ~new_n24711_ & new_n24717_;
  assign new_n24719_ = ~new_n17591_ & ~new_n24691_;
  assign new_n24720_ = ~new_n17590_ & ~new_n24674_;
  assign new_n24721_ = pi0609 & new_n24720_;
  assign new_n24722_ = ~new_n24719_ & ~new_n24721_;
  assign new_n24723_ = pi1155 & ~new_n24722_;
  assign new_n24724_ = ~pi0660 & ~new_n24723_;
  assign new_n24725_ = ~new_n24718_ & new_n24724_;
  assign new_n24726_ = pi0609 & ~new_n24710_;
  assign new_n24727_ = ~pi0609 & new_n24715_;
  assign new_n24728_ = pi1155 & ~new_n24727_;
  assign new_n24729_ = ~new_n24726_ & new_n24728_;
  assign new_n24730_ = ~new_n17603_ & ~new_n24691_;
  assign new_n24731_ = ~pi0609 & new_n24720_;
  assign new_n24732_ = ~new_n24730_ & ~new_n24731_;
  assign new_n24733_ = ~pi1155 & ~new_n24732_;
  assign new_n24734_ = pi0660 & ~new_n24733_;
  assign new_n24735_ = ~new_n24729_ & new_n24734_;
  assign new_n24736_ = ~new_n24725_ & ~new_n24735_;
  assign new_n24737_ = pi0785 & ~new_n24736_;
  assign new_n24738_ = ~pi0785 & ~new_n24710_;
  assign new_n24739_ = ~new_n24737_ & ~new_n24738_;
  assign new_n24740_ = ~pi0618 & ~new_n24739_;
  assign new_n24741_ = ~new_n17618_ & ~new_n24715_;
  assign new_n24742_ = new_n17618_ & ~new_n24691_;
  assign new_n24743_ = ~new_n24741_ & ~new_n24742_;
  assign new_n24744_ = pi0618 & new_n24743_;
  assign new_n24745_ = ~pi1154 & ~new_n24744_;
  assign new_n24746_ = ~new_n24740_ & new_n24745_;
  assign new_n24747_ = new_n17590_ & ~new_n24691_;
  assign new_n24748_ = ~new_n24720_ & ~new_n24747_;
  assign new_n24749_ = ~pi0785 & ~new_n24748_;
  assign new_n24750_ = ~new_n24723_ & ~new_n24733_;
  assign new_n24751_ = pi0785 & ~new_n24750_;
  assign new_n24752_ = ~new_n24749_ & ~new_n24751_;
  assign new_n24753_ = pi0618 & new_n24752_;
  assign new_n24754_ = ~pi0618 & new_n24691_;
  assign new_n24755_ = pi1154 & ~new_n24754_;
  assign new_n24756_ = ~new_n24753_ & new_n24755_;
  assign new_n24757_ = ~pi0627 & ~new_n24756_;
  assign new_n24758_ = ~new_n24746_ & new_n24757_;
  assign new_n24759_ = pi0618 & ~new_n24739_;
  assign new_n24760_ = ~pi0618 & new_n24743_;
  assign new_n24761_ = pi1154 & ~new_n24760_;
  assign new_n24762_ = ~new_n24759_ & new_n24761_;
  assign new_n24763_ = ~pi0618 & new_n24752_;
  assign new_n24764_ = pi0618 & new_n24691_;
  assign new_n24765_ = ~pi1154 & ~new_n24764_;
  assign new_n24766_ = ~new_n24763_ & new_n24765_;
  assign new_n24767_ = pi0627 & ~new_n24766_;
  assign new_n24768_ = ~new_n24762_ & new_n24767_;
  assign new_n24769_ = ~new_n24758_ & ~new_n24768_;
  assign new_n24770_ = pi0781 & ~new_n24769_;
  assign new_n24771_ = ~pi0781 & ~new_n24739_;
  assign new_n24772_ = ~new_n24770_ & ~new_n24771_;
  assign new_n24773_ = ~pi0619 & ~new_n24772_;
  assign new_n24774_ = ~new_n17655_ & new_n24743_;
  assign new_n24775_ = new_n17655_ & new_n24691_;
  assign new_n24776_ = ~new_n24774_ & ~new_n24775_;
  assign new_n24777_ = pi0619 & ~new_n24776_;
  assign new_n24778_ = ~pi1159 & ~new_n24777_;
  assign new_n24779_ = ~new_n24773_ & new_n24778_;
  assign new_n24780_ = ~pi0781 & ~new_n24752_;
  assign new_n24781_ = ~new_n24756_ & ~new_n24766_;
  assign new_n24782_ = pi0781 & ~new_n24781_;
  assign new_n24783_ = ~new_n24780_ & ~new_n24782_;
  assign new_n24784_ = pi0619 & new_n24783_;
  assign new_n24785_ = ~pi0619 & new_n24691_;
  assign new_n24786_ = pi1159 & ~new_n24785_;
  assign new_n24787_ = ~new_n24784_ & new_n24786_;
  assign new_n24788_ = ~pi0648 & ~new_n24787_;
  assign new_n24789_ = ~new_n24779_ & new_n24788_;
  assign new_n24790_ = pi0619 & ~new_n24772_;
  assign new_n24791_ = ~pi0619 & ~new_n24776_;
  assign new_n24792_ = pi1159 & ~new_n24791_;
  assign new_n24793_ = ~new_n24790_ & new_n24792_;
  assign new_n24794_ = ~pi0619 & new_n24783_;
  assign new_n24795_ = pi0619 & new_n24691_;
  assign new_n24796_ = ~pi1159 & ~new_n24795_;
  assign new_n24797_ = ~new_n24794_ & new_n24796_;
  assign new_n24798_ = pi0648 & ~new_n24797_;
  assign new_n24799_ = ~new_n24793_ & new_n24798_;
  assign new_n24800_ = ~new_n24789_ & ~new_n24799_;
  assign new_n24801_ = pi0789 & ~new_n24800_;
  assign new_n24802_ = ~pi0789 & ~new_n24772_;
  assign new_n24803_ = ~new_n24801_ & ~new_n24802_;
  assign new_n24804_ = ~pi0788 & new_n24803_;
  assign new_n24805_ = ~pi0626 & new_n24803_;
  assign new_n24806_ = new_n17691_ & ~new_n24691_;
  assign new_n24807_ = ~new_n17691_ & new_n24776_;
  assign new_n24808_ = ~new_n24806_ & ~new_n24807_;
  assign new_n24809_ = pi0626 & ~new_n24808_;
  assign new_n24810_ = ~pi0641 & ~new_n24809_;
  assign new_n24811_ = ~new_n24805_ & new_n24810_;
  assign new_n24812_ = ~pi0789 & ~new_n24783_;
  assign new_n24813_ = ~new_n24787_ & ~new_n24797_;
  assign new_n24814_ = pi0789 & ~new_n24813_;
  assign new_n24815_ = ~new_n24812_ & ~new_n24814_;
  assign new_n24816_ = ~pi0626 & ~new_n24815_;
  assign new_n24817_ = pi0626 & ~new_n24691_;
  assign new_n24818_ = pi0641 & ~new_n24817_;
  assign new_n24819_ = ~new_n24816_ & new_n24818_;
  assign new_n24820_ = ~pi1158 & ~new_n24819_;
  assign new_n24821_ = ~new_n24811_ & new_n24820_;
  assign new_n24822_ = pi0626 & new_n24803_;
  assign new_n24823_ = ~pi0626 & ~new_n24808_;
  assign new_n24824_ = pi0641 & ~new_n24823_;
  assign new_n24825_ = ~new_n24822_ & new_n24824_;
  assign new_n24826_ = pi0626 & ~new_n24815_;
  assign new_n24827_ = ~pi0626 & ~new_n24691_;
  assign new_n24828_ = ~pi0641 & ~new_n24827_;
  assign new_n24829_ = ~new_n24826_ & new_n24828_;
  assign new_n24830_ = pi1158 & ~new_n24829_;
  assign new_n24831_ = ~new_n24825_ & new_n24830_;
  assign new_n24832_ = ~new_n24821_ & ~new_n24831_;
  assign new_n24833_ = pi0788 & ~new_n24832_;
  assign new_n24834_ = ~new_n24804_ & ~new_n24833_;
  assign new_n24835_ = ~pi0628 & new_n24834_;
  assign new_n24836_ = ~new_n17968_ & new_n24815_;
  assign new_n24837_ = new_n17968_ & new_n24691_;
  assign new_n24838_ = ~new_n24836_ & ~new_n24837_;
  assign new_n24839_ = pi0628 & ~new_n24838_;
  assign new_n24840_ = ~pi1156 & ~new_n24839_;
  assign new_n24841_ = ~new_n24835_ & new_n24840_;
  assign new_n24842_ = ~new_n17734_ & new_n24808_;
  assign new_n24843_ = new_n17734_ & new_n24691_;
  assign new_n24844_ = ~new_n24842_ & ~new_n24843_;
  assign new_n24845_ = pi0628 & ~new_n24844_;
  assign new_n24846_ = ~pi0628 & new_n24691_;
  assign new_n24847_ = pi1156 & ~new_n24846_;
  assign new_n24848_ = ~new_n24845_ & new_n24847_;
  assign new_n24849_ = ~pi0629 & ~new_n24848_;
  assign new_n24850_ = ~new_n24841_ & new_n24849_;
  assign new_n24851_ = pi0628 & new_n24834_;
  assign new_n24852_ = ~pi0628 & ~new_n24838_;
  assign new_n24853_ = pi1156 & ~new_n24852_;
  assign new_n24854_ = ~new_n24851_ & new_n24853_;
  assign new_n24855_ = ~pi0628 & ~new_n24844_;
  assign new_n24856_ = pi0628 & new_n24691_;
  assign new_n24857_ = ~pi1156 & ~new_n24856_;
  assign new_n24858_ = ~new_n24855_ & new_n24857_;
  assign new_n24859_ = pi0629 & ~new_n24858_;
  assign new_n24860_ = ~new_n24854_ & new_n24859_;
  assign new_n24861_ = ~new_n24850_ & ~new_n24860_;
  assign new_n24862_ = pi0792 & ~new_n24861_;
  assign new_n24863_ = ~pi0792 & new_n24834_;
  assign new_n24864_ = ~new_n24862_ & ~new_n24863_;
  assign new_n24865_ = ~pi0647 & ~new_n24864_;
  assign new_n24866_ = ~new_n17762_ & ~new_n24838_;
  assign new_n24867_ = new_n17762_ & new_n24691_;
  assign new_n24868_ = ~new_n24866_ & ~new_n24867_;
  assign new_n24869_ = pi0647 & ~new_n24868_;
  assign new_n24870_ = ~pi1157 & ~new_n24869_;
  assign new_n24871_ = ~new_n24865_ & new_n24870_;
  assign new_n24872_ = ~pi0792 & new_n24844_;
  assign new_n24873_ = ~new_n24848_ & ~new_n24858_;
  assign new_n24874_ = pi0792 & ~new_n24873_;
  assign new_n24875_ = ~new_n24872_ & ~new_n24874_;
  assign new_n24876_ = pi0647 & new_n24875_;
  assign new_n24877_ = ~pi0647 & new_n24691_;
  assign new_n24878_ = pi1157 & ~new_n24877_;
  assign new_n24879_ = ~new_n24876_ & new_n24878_;
  assign new_n24880_ = ~pi0630 & ~new_n24879_;
  assign new_n24881_ = ~new_n24871_ & new_n24880_;
  assign new_n24882_ = pi0647 & ~new_n24864_;
  assign new_n24883_ = ~pi0647 & ~new_n24868_;
  assign new_n24884_ = pi1157 & ~new_n24883_;
  assign new_n24885_ = ~new_n24882_ & new_n24884_;
  assign new_n24886_ = ~pi0647 & new_n24875_;
  assign new_n24887_ = pi0647 & new_n24691_;
  assign new_n24888_ = ~pi1157 & ~new_n24887_;
  assign new_n24889_ = ~new_n24886_ & new_n24888_;
  assign new_n24890_ = pi0630 & ~new_n24889_;
  assign new_n24891_ = ~new_n24885_ & new_n24890_;
  assign new_n24892_ = ~new_n24881_ & ~new_n24891_;
  assign new_n24893_ = pi0787 & ~new_n24892_;
  assign new_n24894_ = ~pi0787 & ~new_n24864_;
  assign new_n24895_ = ~new_n24893_ & ~new_n24894_;
  assign new_n24896_ = ~pi0644 & ~new_n24895_;
  assign new_n24897_ = ~pi0787 & ~new_n24875_;
  assign new_n24898_ = ~new_n24879_ & ~new_n24889_;
  assign new_n24899_ = pi0787 & ~new_n24898_;
  assign new_n24900_ = ~new_n24897_ & ~new_n24899_;
  assign new_n24901_ = pi0644 & new_n24900_;
  assign new_n24902_ = ~pi0715 & ~new_n24901_;
  assign new_n24903_ = ~new_n24896_ & new_n24902_;
  assign new_n24904_ = new_n17804_ & ~new_n24691_;
  assign new_n24905_ = ~new_n17804_ & new_n24868_;
  assign new_n24906_ = ~new_n24904_ & ~new_n24905_;
  assign new_n24907_ = ~pi0644 & new_n24906_;
  assign new_n24908_ = pi0644 & new_n24691_;
  assign new_n24909_ = pi0715 & ~new_n24908_;
  assign new_n24910_ = ~new_n24907_ & new_n24909_;
  assign new_n24911_ = ~pi1160 & ~new_n24910_;
  assign new_n24912_ = ~new_n24903_ & new_n24911_;
  assign new_n24913_ = pi0644 & ~new_n24895_;
  assign new_n24914_ = ~pi0644 & new_n24900_;
  assign new_n24915_ = pi0715 & ~new_n24914_;
  assign new_n24916_ = ~new_n24913_ & new_n24915_;
  assign new_n24917_ = pi0644 & new_n24906_;
  assign new_n24918_ = ~pi0644 & new_n24691_;
  assign new_n24919_ = ~pi0715 & ~new_n24918_;
  assign new_n24920_ = ~new_n24917_ & new_n24919_;
  assign new_n24921_ = pi1160 & ~new_n24920_;
  assign new_n24922_ = ~new_n24916_ & new_n24921_;
  assign new_n24923_ = pi0790 & ~new_n24922_;
  assign new_n24924_ = ~new_n24912_ & new_n24923_;
  assign new_n24925_ = ~pi0790 & new_n24895_;
  assign new_n24926_ = ~po1038 & ~new_n24925_;
  assign new_n24927_ = ~new_n24924_ & new_n24926_;
  assign new_n24928_ = ~pi0177 & po1038;
  assign new_n24929_ = ~pi0832 & ~new_n24928_;
  assign new_n24930_ = ~new_n24927_ & new_n24929_;
  assign new_n24931_ = ~pi0177 & ~new_n2754_;
  assign new_n24932_ = ~pi0757 & new_n16913_;
  assign new_n24933_ = ~new_n24931_ & ~new_n24932_;
  assign new_n24934_ = ~new_n17858_ & ~new_n24933_;
  assign new_n24935_ = ~pi0785 & ~new_n24934_;
  assign new_n24936_ = ~new_n17863_ & ~new_n24933_;
  assign new_n24937_ = pi1155 & ~new_n24936_;
  assign new_n24938_ = ~new_n17866_ & new_n24934_;
  assign new_n24939_ = ~pi1155 & ~new_n24938_;
  assign new_n24940_ = ~new_n24937_ & ~new_n24939_;
  assign new_n24941_ = pi0785 & ~new_n24940_;
  assign new_n24942_ = ~new_n24935_ & ~new_n24941_;
  assign new_n24943_ = ~pi0781 & ~new_n24942_;
  assign new_n24944_ = ~new_n17873_ & new_n24942_;
  assign new_n24945_ = pi1154 & ~new_n24944_;
  assign new_n24946_ = ~new_n17876_ & new_n24942_;
  assign new_n24947_ = ~pi1154 & ~new_n24946_;
  assign new_n24948_ = ~new_n24945_ & ~new_n24947_;
  assign new_n24949_ = pi0781 & ~new_n24948_;
  assign new_n24950_ = ~new_n24943_ & ~new_n24949_;
  assign new_n24951_ = ~pi0789 & ~new_n24950_;
  assign new_n24952_ = pi0619 & new_n24950_;
  assign new_n24953_ = ~pi0619 & new_n24931_;
  assign new_n24954_ = pi1159 & ~new_n24953_;
  assign new_n24955_ = ~new_n24952_ & new_n24954_;
  assign new_n24956_ = ~pi0619 & new_n24950_;
  assign new_n24957_ = pi0619 & new_n24931_;
  assign new_n24958_ = ~pi1159 & ~new_n24957_;
  assign new_n24959_ = ~new_n24956_ & new_n24958_;
  assign new_n24960_ = ~new_n24955_ & ~new_n24959_;
  assign new_n24961_ = pi0789 & ~new_n24960_;
  assign new_n24962_ = ~new_n24951_ & ~new_n24961_;
  assign new_n24963_ = ~new_n17968_ & new_n24962_;
  assign new_n24964_ = new_n17968_ & new_n24931_;
  assign new_n24965_ = ~new_n24963_ & ~new_n24964_;
  assign new_n24966_ = ~new_n17762_ & ~new_n24965_;
  assign new_n24967_ = new_n17762_ & new_n24931_;
  assign new_n24968_ = ~new_n24966_ & ~new_n24967_;
  assign new_n24969_ = ~new_n20556_ & new_n24968_;
  assign new_n24970_ = ~pi0686 & new_n16915_;
  assign new_n24971_ = ~new_n24931_ & ~new_n24970_;
  assign new_n24972_ = ~pi0778 & new_n24971_;
  assign new_n24973_ = ~pi0625 & new_n24970_;
  assign new_n24974_ = ~new_n24971_ & ~new_n24973_;
  assign new_n24975_ = pi1153 & ~new_n24974_;
  assign new_n24976_ = ~pi1153 & ~new_n24931_;
  assign new_n24977_ = ~new_n24973_ & new_n24976_;
  assign new_n24978_ = ~new_n24975_ & ~new_n24977_;
  assign new_n24979_ = pi0778 & ~new_n24978_;
  assign new_n24980_ = ~new_n24972_ & ~new_n24979_;
  assign new_n24981_ = ~new_n17844_ & new_n24980_;
  assign new_n24982_ = ~new_n17846_ & new_n24981_;
  assign new_n24983_ = ~new_n17848_ & new_n24982_;
  assign new_n24984_ = ~new_n17980_ & new_n24983_;
  assign new_n24985_ = ~new_n18011_ & new_n24984_;
  assign new_n24986_ = ~pi0647 & new_n24985_;
  assign new_n24987_ = pi0647 & new_n24931_;
  assign new_n24988_ = ~pi1157 & ~new_n24987_;
  assign new_n24989_ = ~new_n24986_ & new_n24988_;
  assign new_n24990_ = pi0630 & new_n24989_;
  assign new_n24991_ = pi0647 & ~new_n24985_;
  assign new_n24992_ = ~pi0647 & ~new_n24931_;
  assign new_n24993_ = ~new_n24991_ & ~new_n24992_;
  assign new_n24994_ = new_n17801_ & ~new_n24993_;
  assign new_n24995_ = ~new_n24990_ & ~new_n24994_;
  assign new_n24996_ = ~new_n24969_ & new_n24995_;
  assign new_n24997_ = pi0787 & ~new_n24996_;
  assign new_n24998_ = pi0626 & ~new_n24962_;
  assign new_n24999_ = ~pi0626 & ~new_n24931_;
  assign new_n25000_ = new_n17731_ & ~new_n24999_;
  assign new_n25001_ = ~new_n24998_ & new_n25000_;
  assign new_n25002_ = new_n17856_ & new_n24983_;
  assign new_n25003_ = ~pi0626 & ~new_n24962_;
  assign new_n25004_ = pi0626 & ~new_n24931_;
  assign new_n25005_ = new_n17732_ & ~new_n25004_;
  assign new_n25006_ = ~new_n25003_ & new_n25005_;
  assign new_n25007_ = ~new_n25002_ & ~new_n25006_;
  assign new_n25008_ = ~new_n25001_ & new_n25007_;
  assign new_n25009_ = pi0788 & ~new_n25008_;
  assign new_n25010_ = ~new_n16639_ & ~new_n24971_;
  assign new_n25011_ = pi0625 & new_n25010_;
  assign new_n25012_ = new_n24933_ & ~new_n25010_;
  assign new_n25013_ = ~new_n25011_ & ~new_n25012_;
  assign new_n25014_ = new_n24976_ & ~new_n25013_;
  assign new_n25015_ = ~pi0608 & ~new_n24975_;
  assign new_n25016_ = ~new_n25014_ & new_n25015_;
  assign new_n25017_ = pi1153 & new_n24933_;
  assign new_n25018_ = ~new_n25011_ & new_n25017_;
  assign new_n25019_ = pi0608 & ~new_n24977_;
  assign new_n25020_ = ~new_n25018_ & new_n25019_;
  assign new_n25021_ = ~new_n25016_ & ~new_n25020_;
  assign new_n25022_ = pi0778 & ~new_n25021_;
  assign new_n25023_ = ~pi0778 & ~new_n25012_;
  assign new_n25024_ = ~new_n25022_ & ~new_n25023_;
  assign new_n25025_ = ~pi0609 & ~new_n25024_;
  assign new_n25026_ = pi0609 & new_n24980_;
  assign new_n25027_ = ~pi1155 & ~new_n25026_;
  assign new_n25028_ = ~new_n25025_ & new_n25027_;
  assign new_n25029_ = ~pi0660 & ~new_n24937_;
  assign new_n25030_ = ~new_n25028_ & new_n25029_;
  assign new_n25031_ = pi0609 & ~new_n25024_;
  assign new_n25032_ = ~pi0609 & new_n24980_;
  assign new_n25033_ = pi1155 & ~new_n25032_;
  assign new_n25034_ = ~new_n25031_ & new_n25033_;
  assign new_n25035_ = pi0660 & ~new_n24939_;
  assign new_n25036_ = ~new_n25034_ & new_n25035_;
  assign new_n25037_ = ~new_n25030_ & ~new_n25036_;
  assign new_n25038_ = pi0785 & ~new_n25037_;
  assign new_n25039_ = ~pi0785 & ~new_n25024_;
  assign new_n25040_ = ~new_n25038_ & ~new_n25039_;
  assign new_n25041_ = ~pi0618 & ~new_n25040_;
  assign new_n25042_ = pi0618 & new_n24981_;
  assign new_n25043_ = ~pi1154 & ~new_n25042_;
  assign new_n25044_ = ~new_n25041_ & new_n25043_;
  assign new_n25045_ = ~pi0627 & ~new_n24945_;
  assign new_n25046_ = ~new_n25044_ & new_n25045_;
  assign new_n25047_ = pi0618 & ~new_n25040_;
  assign new_n25048_ = ~pi0618 & new_n24981_;
  assign new_n25049_ = pi1154 & ~new_n25048_;
  assign new_n25050_ = ~new_n25047_ & new_n25049_;
  assign new_n25051_ = pi0627 & ~new_n24947_;
  assign new_n25052_ = ~new_n25050_ & new_n25051_;
  assign new_n25053_ = ~new_n25046_ & ~new_n25052_;
  assign new_n25054_ = pi0781 & ~new_n25053_;
  assign new_n25055_ = ~pi0781 & ~new_n25040_;
  assign new_n25056_ = ~new_n25054_ & ~new_n25055_;
  assign new_n25057_ = pi0619 & ~new_n25056_;
  assign new_n25058_ = ~pi0619 & new_n24982_;
  assign new_n25059_ = pi1159 & ~new_n25058_;
  assign new_n25060_ = ~new_n25057_ & new_n25059_;
  assign new_n25061_ = pi0648 & ~new_n24959_;
  assign new_n25062_ = ~new_n25060_ & new_n25061_;
  assign new_n25063_ = ~pi0619 & ~new_n25056_;
  assign new_n25064_ = pi0619 & new_n24982_;
  assign new_n25065_ = ~pi1159 & ~new_n25064_;
  assign new_n25066_ = ~new_n25063_ & new_n25065_;
  assign new_n25067_ = ~pi0648 & ~new_n24955_;
  assign new_n25068_ = ~new_n25066_ & new_n25067_;
  assign new_n25069_ = pi0789 & ~new_n25068_;
  assign new_n25070_ = ~new_n25062_ & new_n25069_;
  assign new_n25071_ = ~pi0789 & new_n25056_;
  assign new_n25072_ = new_n17969_ & ~new_n25071_;
  assign new_n25073_ = ~new_n25070_ & new_n25072_;
  assign new_n25074_ = ~new_n25009_ & ~new_n25073_;
  assign new_n25075_ = ~new_n20364_ & ~new_n25074_;
  assign new_n25076_ = new_n18008_ & ~new_n24965_;
  assign new_n25077_ = new_n20851_ & new_n24984_;
  assign new_n25078_ = ~new_n25076_ & ~new_n25077_;
  assign new_n25079_ = ~pi0629 & ~new_n25078_;
  assign new_n25080_ = new_n20855_ & new_n24984_;
  assign new_n25081_ = new_n18007_ & ~new_n24965_;
  assign new_n25082_ = ~new_n25080_ & ~new_n25081_;
  assign new_n25083_ = pi0629 & ~new_n25082_;
  assign new_n25084_ = ~new_n25079_ & ~new_n25083_;
  assign new_n25085_ = pi0792 & ~new_n25084_;
  assign new_n25086_ = ~new_n20360_ & ~new_n25085_;
  assign new_n25087_ = ~new_n25075_ & new_n25086_;
  assign new_n25088_ = ~new_n24997_ & ~new_n25087_;
  assign new_n25089_ = pi0644 & new_n25088_;
  assign new_n25090_ = ~pi0787 & ~new_n24985_;
  assign new_n25091_ = pi1157 & ~new_n24993_;
  assign new_n25092_ = ~new_n24989_ & ~new_n25091_;
  assign new_n25093_ = pi0787 & ~new_n25092_;
  assign new_n25094_ = ~new_n25090_ & ~new_n25093_;
  assign new_n25095_ = ~pi0644 & new_n25094_;
  assign new_n25096_ = pi0715 & ~new_n25095_;
  assign new_n25097_ = ~new_n25089_ & new_n25096_;
  assign new_n25098_ = ~new_n17804_ & ~new_n24968_;
  assign new_n25099_ = new_n17804_ & new_n24931_;
  assign new_n25100_ = ~new_n25098_ & ~new_n25099_;
  assign new_n25101_ = pi0644 & ~new_n25100_;
  assign new_n25102_ = ~pi0644 & new_n24931_;
  assign new_n25103_ = ~pi0715 & ~new_n25102_;
  assign new_n25104_ = ~new_n25101_ & new_n25103_;
  assign new_n25105_ = pi1160 & ~new_n25104_;
  assign new_n25106_ = ~new_n25097_ & new_n25105_;
  assign new_n25107_ = ~pi0644 & new_n25088_;
  assign new_n25108_ = pi0644 & new_n25094_;
  assign new_n25109_ = ~pi0715 & ~new_n25108_;
  assign new_n25110_ = ~new_n25107_ & new_n25109_;
  assign new_n25111_ = ~pi0644 & ~new_n25100_;
  assign new_n25112_ = pi0644 & new_n24931_;
  assign new_n25113_ = pi0715 & ~new_n25112_;
  assign new_n25114_ = ~new_n25111_ & new_n25113_;
  assign new_n25115_ = ~pi1160 & ~new_n25114_;
  assign new_n25116_ = ~new_n25110_ & new_n25115_;
  assign new_n25117_ = ~new_n25106_ & ~new_n25116_;
  assign new_n25118_ = pi0790 & ~new_n25117_;
  assign new_n25119_ = ~pi0790 & new_n25088_;
  assign new_n25120_ = pi0832 & ~new_n25119_;
  assign new_n25121_ = ~new_n25118_ & new_n25120_;
  assign po0334 = ~new_n24930_ & ~new_n25121_;
  assign new_n25123_ = ~pi0178 & ~new_n2754_;
  assign new_n25124_ = ~pi0760 & new_n16913_;
  assign new_n25125_ = ~new_n25123_ & ~new_n25124_;
  assign new_n25126_ = ~new_n17858_ & ~new_n25125_;
  assign new_n25127_ = ~pi0785 & ~new_n25126_;
  assign new_n25128_ = new_n17603_ & new_n25124_;
  assign new_n25129_ = new_n25126_ & ~new_n25128_;
  assign new_n25130_ = pi1155 & ~new_n25129_;
  assign new_n25131_ = ~pi1155 & ~new_n25123_;
  assign new_n25132_ = ~new_n25128_ & new_n25131_;
  assign new_n25133_ = ~new_n25130_ & ~new_n25132_;
  assign new_n25134_ = pi0785 & ~new_n25133_;
  assign new_n25135_ = ~new_n25127_ & ~new_n25134_;
  assign new_n25136_ = ~pi0781 & ~new_n25135_;
  assign new_n25137_ = ~new_n17873_ & new_n25135_;
  assign new_n25138_ = pi1154 & ~new_n25137_;
  assign new_n25139_ = ~new_n17876_ & new_n25135_;
  assign new_n25140_ = ~pi1154 & ~new_n25139_;
  assign new_n25141_ = ~new_n25138_ & ~new_n25140_;
  assign new_n25142_ = pi0781 & ~new_n25141_;
  assign new_n25143_ = ~new_n25136_ & ~new_n25142_;
  assign new_n25144_ = ~pi0789 & ~new_n25143_;
  assign new_n25145_ = ~new_n23057_ & new_n25143_;
  assign new_n25146_ = pi1159 & ~new_n25145_;
  assign new_n25147_ = ~new_n23060_ & new_n25143_;
  assign new_n25148_ = ~pi1159 & ~new_n25147_;
  assign new_n25149_ = ~new_n25146_ & ~new_n25148_;
  assign new_n25150_ = pi0789 & ~new_n25149_;
  assign new_n25151_ = ~new_n25144_ & ~new_n25150_;
  assign new_n25152_ = ~new_n17968_ & new_n25151_;
  assign new_n25153_ = new_n17968_ & new_n25123_;
  assign new_n25154_ = ~new_n25152_ & ~new_n25153_;
  assign new_n25155_ = ~new_n17762_ & ~new_n25154_;
  assign new_n25156_ = new_n17762_ & new_n25123_;
  assign new_n25157_ = ~new_n25155_ & ~new_n25156_;
  assign new_n25158_ = ~new_n20556_ & new_n25157_;
  assign new_n25159_ = ~pi0688 & new_n16915_;
  assign new_n25160_ = ~new_n25123_ & ~new_n25159_;
  assign new_n25161_ = ~pi0778 & ~new_n25160_;
  assign new_n25162_ = ~pi0625 & new_n25159_;
  assign new_n25163_ = ~new_n25160_ & ~new_n25162_;
  assign new_n25164_ = pi1153 & ~new_n25163_;
  assign new_n25165_ = ~pi1153 & ~new_n25123_;
  assign new_n25166_ = ~new_n25162_ & new_n25165_;
  assign new_n25167_ = pi0778 & ~new_n25166_;
  assign new_n25168_ = ~new_n25164_ & new_n25167_;
  assign new_n25169_ = ~new_n25161_ & ~new_n25168_;
  assign new_n25170_ = ~new_n17844_ & ~new_n25169_;
  assign new_n25171_ = ~new_n17846_ & new_n25170_;
  assign new_n25172_ = ~new_n17848_ & new_n25171_;
  assign new_n25173_ = ~new_n17980_ & new_n25172_;
  assign new_n25174_ = ~new_n18011_ & new_n25173_;
  assign new_n25175_ = ~pi0647 & new_n25174_;
  assign new_n25176_ = pi0647 & new_n25123_;
  assign new_n25177_ = ~pi1157 & ~new_n25176_;
  assign new_n25178_ = ~new_n25175_ & new_n25177_;
  assign new_n25179_ = pi0630 & new_n25178_;
  assign new_n25180_ = pi0647 & ~new_n25174_;
  assign new_n25181_ = ~pi0647 & ~new_n25123_;
  assign new_n25182_ = ~new_n25180_ & ~new_n25181_;
  assign new_n25183_ = new_n17801_ & ~new_n25182_;
  assign new_n25184_ = ~new_n25179_ & ~new_n25183_;
  assign new_n25185_ = ~new_n25158_ & new_n25184_;
  assign new_n25186_ = pi0787 & ~new_n25185_;
  assign new_n25187_ = pi0626 & ~new_n25151_;
  assign new_n25188_ = ~pi0626 & ~new_n25123_;
  assign new_n25189_ = new_n17731_ & ~new_n25188_;
  assign new_n25190_ = ~new_n25187_ & new_n25189_;
  assign new_n25191_ = new_n17856_ & new_n25172_;
  assign new_n25192_ = ~pi0626 & ~new_n25151_;
  assign new_n25193_ = pi0626 & ~new_n25123_;
  assign new_n25194_ = new_n17732_ & ~new_n25193_;
  assign new_n25195_ = ~new_n25192_ & new_n25194_;
  assign new_n25196_ = ~new_n25191_ & ~new_n25195_;
  assign new_n25197_ = ~new_n25190_ & new_n25196_;
  assign new_n25198_ = pi0788 & ~new_n25197_;
  assign new_n25199_ = ~new_n16639_ & ~new_n25160_;
  assign new_n25200_ = pi0625 & new_n25199_;
  assign new_n25201_ = new_n25125_ & ~new_n25199_;
  assign new_n25202_ = ~new_n25200_ & ~new_n25201_;
  assign new_n25203_ = new_n25165_ & ~new_n25202_;
  assign new_n25204_ = ~pi0608 & ~new_n25164_;
  assign new_n25205_ = ~new_n25203_ & new_n25204_;
  assign new_n25206_ = pi1153 & new_n25125_;
  assign new_n25207_ = ~new_n25200_ & new_n25206_;
  assign new_n25208_ = pi0608 & ~new_n25166_;
  assign new_n25209_ = ~new_n25207_ & new_n25208_;
  assign new_n25210_ = ~new_n25205_ & ~new_n25209_;
  assign new_n25211_ = pi0778 & ~new_n25210_;
  assign new_n25212_ = ~pi0778 & ~new_n25201_;
  assign new_n25213_ = ~new_n25211_ & ~new_n25212_;
  assign new_n25214_ = ~pi0609 & ~new_n25213_;
  assign new_n25215_ = pi0609 & ~new_n25169_;
  assign new_n25216_ = ~pi1155 & ~new_n25215_;
  assign new_n25217_ = ~new_n25214_ & new_n25216_;
  assign new_n25218_ = ~pi0660 & ~new_n25130_;
  assign new_n25219_ = ~new_n25217_ & new_n25218_;
  assign new_n25220_ = pi0609 & ~new_n25213_;
  assign new_n25221_ = ~pi0609 & ~new_n25169_;
  assign new_n25222_ = pi1155 & ~new_n25221_;
  assign new_n25223_ = ~new_n25220_ & new_n25222_;
  assign new_n25224_ = pi0660 & ~new_n25132_;
  assign new_n25225_ = ~new_n25223_ & new_n25224_;
  assign new_n25226_ = ~new_n25219_ & ~new_n25225_;
  assign new_n25227_ = pi0785 & ~new_n25226_;
  assign new_n25228_ = ~pi0785 & ~new_n25213_;
  assign new_n25229_ = ~new_n25227_ & ~new_n25228_;
  assign new_n25230_ = ~pi0618 & ~new_n25229_;
  assign new_n25231_ = pi0618 & new_n25170_;
  assign new_n25232_ = ~pi1154 & ~new_n25231_;
  assign new_n25233_ = ~new_n25230_ & new_n25232_;
  assign new_n25234_ = ~pi0627 & ~new_n25138_;
  assign new_n25235_ = ~new_n25233_ & new_n25234_;
  assign new_n25236_ = pi0618 & ~new_n25229_;
  assign new_n25237_ = ~pi0618 & new_n25170_;
  assign new_n25238_ = pi1154 & ~new_n25237_;
  assign new_n25239_ = ~new_n25236_ & new_n25238_;
  assign new_n25240_ = pi0627 & ~new_n25140_;
  assign new_n25241_ = ~new_n25239_ & new_n25240_;
  assign new_n25242_ = ~new_n25235_ & ~new_n25241_;
  assign new_n25243_ = pi0781 & ~new_n25242_;
  assign new_n25244_ = ~pi0781 & ~new_n25229_;
  assign new_n25245_ = ~new_n25243_ & ~new_n25244_;
  assign new_n25246_ = pi0619 & ~new_n25245_;
  assign new_n25247_ = ~pi0619 & new_n25171_;
  assign new_n25248_ = pi1159 & ~new_n25247_;
  assign new_n25249_ = ~new_n25246_ & new_n25248_;
  assign new_n25250_ = pi0648 & ~new_n25148_;
  assign new_n25251_ = ~new_n25249_ & new_n25250_;
  assign new_n25252_ = ~pi0619 & ~new_n25245_;
  assign new_n25253_ = pi0619 & new_n25171_;
  assign new_n25254_ = ~pi1159 & ~new_n25253_;
  assign new_n25255_ = ~new_n25252_ & new_n25254_;
  assign new_n25256_ = ~pi0648 & ~new_n25146_;
  assign new_n25257_ = ~new_n25255_ & new_n25256_;
  assign new_n25258_ = pi0789 & ~new_n25257_;
  assign new_n25259_ = ~new_n25251_ & new_n25258_;
  assign new_n25260_ = ~pi0789 & new_n25245_;
  assign new_n25261_ = new_n17969_ & ~new_n25260_;
  assign new_n25262_ = ~new_n25259_ & new_n25261_;
  assign new_n25263_ = ~new_n25198_ & ~new_n25262_;
  assign new_n25264_ = ~new_n20364_ & ~new_n25263_;
  assign new_n25265_ = new_n18008_ & ~new_n25154_;
  assign new_n25266_ = new_n20851_ & new_n25173_;
  assign new_n25267_ = ~new_n25265_ & ~new_n25266_;
  assign new_n25268_ = ~pi0629 & ~new_n25267_;
  assign new_n25269_ = new_n20855_ & new_n25173_;
  assign new_n25270_ = new_n18007_ & ~new_n25154_;
  assign new_n25271_ = ~new_n25269_ & ~new_n25270_;
  assign new_n25272_ = pi0629 & ~new_n25271_;
  assign new_n25273_ = ~new_n25268_ & ~new_n25272_;
  assign new_n25274_ = pi0792 & ~new_n25273_;
  assign new_n25275_ = ~new_n20360_ & ~new_n25274_;
  assign new_n25276_ = ~new_n25264_ & new_n25275_;
  assign new_n25277_ = ~new_n25186_ & ~new_n25276_;
  assign new_n25278_ = pi0644 & new_n25277_;
  assign new_n25279_ = ~pi0787 & ~new_n25174_;
  assign new_n25280_ = pi1157 & ~new_n25182_;
  assign new_n25281_ = ~new_n25178_ & ~new_n25280_;
  assign new_n25282_ = pi0787 & ~new_n25281_;
  assign new_n25283_ = ~new_n25279_ & ~new_n25282_;
  assign new_n25284_ = ~pi0644 & new_n25283_;
  assign new_n25285_ = pi0715 & ~new_n25284_;
  assign new_n25286_ = ~new_n25278_ & new_n25285_;
  assign new_n25287_ = ~new_n17804_ & ~new_n25157_;
  assign new_n25288_ = new_n17804_ & new_n25123_;
  assign new_n25289_ = ~new_n25287_ & ~new_n25288_;
  assign new_n25290_ = pi0644 & ~new_n25289_;
  assign new_n25291_ = ~pi0644 & new_n25123_;
  assign new_n25292_ = ~pi0715 & ~new_n25291_;
  assign new_n25293_ = ~new_n25290_ & new_n25292_;
  assign new_n25294_ = pi1160 & ~new_n25293_;
  assign new_n25295_ = ~new_n25286_ & new_n25294_;
  assign new_n25296_ = ~pi0644 & new_n25277_;
  assign new_n25297_ = pi0644 & new_n25283_;
  assign new_n25298_ = ~pi0715 & ~new_n25297_;
  assign new_n25299_ = ~new_n25296_ & new_n25298_;
  assign new_n25300_ = ~pi0644 & ~new_n25289_;
  assign new_n25301_ = pi0644 & new_n25123_;
  assign new_n25302_ = pi0715 & ~new_n25301_;
  assign new_n25303_ = ~new_n25300_ & new_n25302_;
  assign new_n25304_ = ~pi1160 & ~new_n25303_;
  assign new_n25305_ = ~new_n25299_ & new_n25304_;
  assign new_n25306_ = ~new_n25295_ & ~new_n25305_;
  assign new_n25307_ = pi0790 & ~new_n25306_;
  assign new_n25308_ = ~pi0790 & new_n25277_;
  assign new_n25309_ = pi0832 & ~new_n25308_;
  assign new_n25310_ = ~new_n25307_ & new_n25309_;
  assign new_n25311_ = ~pi0178 & ~new_n17558_;
  assign new_n25312_ = new_n17691_ & ~new_n25311_;
  assign new_n25313_ = ~pi0688 & new_n3272_;
  assign new_n25314_ = new_n25311_ & ~new_n25313_;
  assign new_n25315_ = pi0178 & ~new_n18128_;
  assign new_n25316_ = ~pi0038 & ~new_n25315_;
  assign new_n25317_ = new_n3272_ & ~new_n25316_;
  assign new_n25318_ = ~pi0178 & new_n18124_;
  assign new_n25319_ = ~new_n25317_ & ~new_n25318_;
  assign new_n25320_ = ~pi0178 & ~new_n17431_;
  assign new_n25321_ = new_n17544_ & ~new_n25320_;
  assign new_n25322_ = ~pi0688 & ~new_n25321_;
  assign new_n25323_ = ~new_n25319_ & new_n25322_;
  assign new_n25324_ = ~new_n25314_ & ~new_n25323_;
  assign new_n25325_ = ~pi0778 & new_n25324_;
  assign new_n25326_ = pi0625 & ~new_n25324_;
  assign new_n25327_ = ~pi0625 & new_n25311_;
  assign new_n25328_ = pi1153 & ~new_n25327_;
  assign new_n25329_ = ~new_n25326_ & new_n25328_;
  assign new_n25330_ = ~pi0625 & ~new_n25324_;
  assign new_n25331_ = pi0625 & new_n25311_;
  assign new_n25332_ = ~pi1153 & ~new_n25331_;
  assign new_n25333_ = ~new_n25330_ & new_n25332_;
  assign new_n25334_ = ~new_n25329_ & ~new_n25333_;
  assign new_n25335_ = pi0778 & ~new_n25334_;
  assign new_n25336_ = ~new_n25325_ & ~new_n25335_;
  assign new_n25337_ = ~new_n17618_ & ~new_n25336_;
  assign new_n25338_ = new_n17618_ & ~new_n25311_;
  assign new_n25339_ = ~new_n25337_ & ~new_n25338_;
  assign new_n25340_ = ~new_n17655_ & new_n25339_;
  assign new_n25341_ = new_n17655_ & new_n25311_;
  assign new_n25342_ = ~new_n25340_ & ~new_n25341_;
  assign new_n25343_ = ~new_n17691_ & new_n25342_;
  assign new_n25344_ = ~new_n25312_ & ~new_n25343_;
  assign new_n25345_ = ~new_n17734_ & new_n25344_;
  assign new_n25346_ = new_n17734_ & new_n25311_;
  assign new_n25347_ = ~new_n25345_ & ~new_n25346_;
  assign new_n25348_ = ~pi0792 & new_n25347_;
  assign new_n25349_ = pi0628 & ~new_n25347_;
  assign new_n25350_ = ~pi0628 & new_n25311_;
  assign new_n25351_ = pi1156 & ~new_n25350_;
  assign new_n25352_ = ~new_n25349_ & new_n25351_;
  assign new_n25353_ = ~pi0628 & ~new_n25347_;
  assign new_n25354_ = pi0628 & new_n25311_;
  assign new_n25355_ = ~pi1156 & ~new_n25354_;
  assign new_n25356_ = ~new_n25353_ & new_n25355_;
  assign new_n25357_ = ~new_n25352_ & ~new_n25356_;
  assign new_n25358_ = pi0792 & ~new_n25357_;
  assign new_n25359_ = ~new_n25348_ & ~new_n25358_;
  assign new_n25360_ = ~pi0647 & ~new_n25359_;
  assign new_n25361_ = pi0647 & ~new_n25311_;
  assign new_n25362_ = ~new_n25360_ & ~new_n25361_;
  assign new_n25363_ = ~pi1157 & new_n25362_;
  assign new_n25364_ = pi0647 & ~new_n25359_;
  assign new_n25365_ = ~pi0647 & ~new_n25311_;
  assign new_n25366_ = ~new_n25364_ & ~new_n25365_;
  assign new_n25367_ = pi1157 & new_n25366_;
  assign new_n25368_ = ~new_n25363_ & ~new_n25367_;
  assign new_n25369_ = pi0787 & ~new_n25368_;
  assign new_n25370_ = ~pi0787 & new_n25359_;
  assign new_n25371_ = ~new_n25369_ & ~new_n25370_;
  assign new_n25372_ = ~pi0644 & ~new_n25371_;
  assign new_n25373_ = pi0715 & ~new_n25372_;
  assign new_n25374_ = pi0178 & ~new_n3272_;
  assign new_n25375_ = ~pi0760 & new_n17433_;
  assign new_n25376_ = ~new_n25320_ & ~new_n25375_;
  assign new_n25377_ = pi0038 & ~new_n25376_;
  assign new_n25378_ = ~pi0178 & new_n17393_;
  assign new_n25379_ = pi0178 & ~new_n17426_;
  assign new_n25380_ = ~pi0760 & ~new_n25379_;
  assign new_n25381_ = ~new_n25378_ & new_n25380_;
  assign new_n25382_ = ~pi0178 & pi0760;
  assign new_n25383_ = ~new_n17349_ & new_n25382_;
  assign new_n25384_ = ~new_n25381_ & ~new_n25383_;
  assign new_n25385_ = ~pi0038 & ~new_n25384_;
  assign new_n25386_ = ~new_n25377_ & ~new_n25385_;
  assign new_n25387_ = new_n3272_ & new_n25386_;
  assign new_n25388_ = ~new_n25374_ & ~new_n25387_;
  assign new_n25389_ = ~new_n17590_ & ~new_n25388_;
  assign new_n25390_ = new_n17590_ & ~new_n25311_;
  assign new_n25391_ = ~new_n25389_ & ~new_n25390_;
  assign new_n25392_ = ~pi0785 & ~new_n25391_;
  assign new_n25393_ = ~new_n17591_ & ~new_n25311_;
  assign new_n25394_ = pi0609 & new_n25389_;
  assign new_n25395_ = ~new_n25393_ & ~new_n25394_;
  assign new_n25396_ = pi1155 & ~new_n25395_;
  assign new_n25397_ = ~new_n17603_ & ~new_n25311_;
  assign new_n25398_ = ~pi0609 & new_n25389_;
  assign new_n25399_ = ~new_n25397_ & ~new_n25398_;
  assign new_n25400_ = ~pi1155 & ~new_n25399_;
  assign new_n25401_ = ~new_n25396_ & ~new_n25400_;
  assign new_n25402_ = pi0785 & ~new_n25401_;
  assign new_n25403_ = ~new_n25392_ & ~new_n25402_;
  assign new_n25404_ = ~pi0781 & ~new_n25403_;
  assign new_n25405_ = pi0618 & new_n25403_;
  assign new_n25406_ = ~pi0618 & new_n25311_;
  assign new_n25407_ = pi1154 & ~new_n25406_;
  assign new_n25408_ = ~new_n25405_ & new_n25407_;
  assign new_n25409_ = ~pi0618 & new_n25403_;
  assign new_n25410_ = pi0618 & new_n25311_;
  assign new_n25411_ = ~pi1154 & ~new_n25410_;
  assign new_n25412_ = ~new_n25409_ & new_n25411_;
  assign new_n25413_ = ~new_n25408_ & ~new_n25412_;
  assign new_n25414_ = pi0781 & ~new_n25413_;
  assign new_n25415_ = ~new_n25404_ & ~new_n25414_;
  assign new_n25416_ = ~pi0789 & ~new_n25415_;
  assign new_n25417_ = pi0619 & new_n25415_;
  assign new_n25418_ = ~pi0619 & new_n25311_;
  assign new_n25419_ = pi1159 & ~new_n25418_;
  assign new_n25420_ = ~new_n25417_ & new_n25419_;
  assign new_n25421_ = ~pi0619 & new_n25415_;
  assign new_n25422_ = pi0619 & new_n25311_;
  assign new_n25423_ = ~pi1159 & ~new_n25422_;
  assign new_n25424_ = ~new_n25421_ & new_n25423_;
  assign new_n25425_ = ~new_n25420_ & ~new_n25424_;
  assign new_n25426_ = pi0789 & ~new_n25425_;
  assign new_n25427_ = ~new_n25416_ & ~new_n25426_;
  assign new_n25428_ = ~new_n17968_ & new_n25427_;
  assign new_n25429_ = new_n17968_ & new_n25311_;
  assign new_n25430_ = ~new_n25428_ & ~new_n25429_;
  assign new_n25431_ = ~new_n17762_ & ~new_n25430_;
  assign new_n25432_ = new_n17762_ & new_n25311_;
  assign new_n25433_ = ~new_n25431_ & ~new_n25432_;
  assign new_n25434_ = ~new_n17804_ & ~new_n25433_;
  assign new_n25435_ = new_n17804_ & new_n25311_;
  assign new_n25436_ = ~new_n25434_ & ~new_n25435_;
  assign new_n25437_ = pi0644 & ~new_n25436_;
  assign new_n25438_ = ~pi0644 & new_n25311_;
  assign new_n25439_ = ~pi0715 & ~new_n25438_;
  assign new_n25440_ = ~new_n25437_ & new_n25439_;
  assign new_n25441_ = pi1160 & ~new_n25440_;
  assign new_n25442_ = ~new_n25373_ & new_n25441_;
  assign new_n25443_ = pi0644 & ~new_n25371_;
  assign new_n25444_ = ~pi0715 & ~new_n25443_;
  assign new_n25445_ = ~pi0644 & ~new_n25436_;
  assign new_n25446_ = pi0644 & new_n25311_;
  assign new_n25447_ = pi0715 & ~new_n25446_;
  assign new_n25448_ = ~new_n25445_ & new_n25447_;
  assign new_n25449_ = ~pi1160 & ~new_n25448_;
  assign new_n25450_ = ~new_n25444_ & new_n25449_;
  assign new_n25451_ = ~new_n25442_ & ~new_n25450_;
  assign new_n25452_ = pi0790 & ~new_n25451_;
  assign new_n25453_ = pi0644 & new_n25441_;
  assign new_n25454_ = ~pi0644 & new_n25449_;
  assign new_n25455_ = pi0790 & ~new_n25454_;
  assign new_n25456_ = ~new_n25453_ & new_n25455_;
  assign new_n25457_ = ~new_n20567_ & new_n25430_;
  assign new_n25458_ = ~pi0629 & new_n25352_;
  assign new_n25459_ = pi0629 & new_n25356_;
  assign new_n25460_ = ~new_n25458_ & ~new_n25459_;
  assign new_n25461_ = ~new_n25457_ & new_n25460_;
  assign new_n25462_ = pi0792 & ~new_n25461_;
  assign new_n25463_ = pi0688 & ~new_n25386_;
  assign new_n25464_ = ~pi0178 & new_n16810_;
  assign new_n25465_ = pi0178 & new_n16928_;
  assign new_n25466_ = pi0760 & ~new_n25465_;
  assign new_n25467_ = ~new_n25464_ & new_n25466_;
  assign new_n25468_ = pi0178 & new_n17007_;
  assign new_n25469_ = ~pi0178 & ~new_n17074_;
  assign new_n25470_ = ~pi0760 & ~new_n25469_;
  assign new_n25471_ = ~new_n25468_ & new_n25470_;
  assign new_n25472_ = pi0039 & ~new_n25471_;
  assign new_n25473_ = ~new_n25467_ & new_n25472_;
  assign new_n25474_ = ~pi0178 & ~new_n17217_;
  assign new_n25475_ = pi0178 & ~new_n17178_;
  assign new_n25476_ = pi0760 & ~new_n25475_;
  assign new_n25477_ = ~new_n25474_ & new_n25476_;
  assign new_n25478_ = ~pi0178 & new_n17227_;
  assign new_n25479_ = pi0178 & new_n17234_;
  assign new_n25480_ = ~pi0760 & ~new_n25479_;
  assign new_n25481_ = ~new_n25478_ & new_n25480_;
  assign new_n25482_ = ~new_n25477_ & ~new_n25481_;
  assign new_n25483_ = ~pi0039 & ~new_n25482_;
  assign new_n25484_ = ~pi0038 & ~new_n25483_;
  assign new_n25485_ = ~new_n25473_ & new_n25484_;
  assign new_n25486_ = ~pi0760 & ~new_n17035_;
  assign new_n25487_ = new_n19383_ & ~new_n25486_;
  assign new_n25488_ = ~pi0178 & ~new_n25487_;
  assign new_n25489_ = ~new_n16916_ & ~new_n25124_;
  assign new_n25490_ = pi0178 & ~new_n25489_;
  assign new_n25491_ = new_n6257_ & new_n25490_;
  assign new_n25492_ = pi0038 & ~new_n25491_;
  assign new_n25493_ = ~new_n25488_ & new_n25492_;
  assign new_n25494_ = ~pi0688 & ~new_n25493_;
  assign new_n25495_ = ~new_n25485_ & new_n25494_;
  assign new_n25496_ = new_n3272_ & ~new_n25495_;
  assign new_n25497_ = ~new_n25463_ & new_n25496_;
  assign new_n25498_ = ~new_n25374_ & ~new_n25497_;
  assign new_n25499_ = ~pi0625 & new_n25498_;
  assign new_n25500_ = pi0625 & new_n25388_;
  assign new_n25501_ = ~pi1153 & ~new_n25500_;
  assign new_n25502_ = ~new_n25499_ & new_n25501_;
  assign new_n25503_ = ~pi0608 & ~new_n25329_;
  assign new_n25504_ = ~new_n25502_ & new_n25503_;
  assign new_n25505_ = pi0625 & new_n25498_;
  assign new_n25506_ = ~pi0625 & new_n25388_;
  assign new_n25507_ = pi1153 & ~new_n25506_;
  assign new_n25508_ = ~new_n25505_ & new_n25507_;
  assign new_n25509_ = pi0608 & ~new_n25333_;
  assign new_n25510_ = ~new_n25508_ & new_n25509_;
  assign new_n25511_ = ~new_n25504_ & ~new_n25510_;
  assign new_n25512_ = pi0778 & ~new_n25511_;
  assign new_n25513_ = ~pi0778 & new_n25498_;
  assign new_n25514_ = ~new_n25512_ & ~new_n25513_;
  assign new_n25515_ = ~pi0609 & ~new_n25514_;
  assign new_n25516_ = pi0609 & new_n25336_;
  assign new_n25517_ = ~pi1155 & ~new_n25516_;
  assign new_n25518_ = ~new_n25515_ & new_n25517_;
  assign new_n25519_ = ~pi0660 & ~new_n25396_;
  assign new_n25520_ = ~new_n25518_ & new_n25519_;
  assign new_n25521_ = pi0609 & ~new_n25514_;
  assign new_n25522_ = ~pi0609 & new_n25336_;
  assign new_n25523_ = pi1155 & ~new_n25522_;
  assign new_n25524_ = ~new_n25521_ & new_n25523_;
  assign new_n25525_ = pi0660 & ~new_n25400_;
  assign new_n25526_ = ~new_n25524_ & new_n25525_;
  assign new_n25527_ = ~new_n25520_ & ~new_n25526_;
  assign new_n25528_ = pi0785 & ~new_n25527_;
  assign new_n25529_ = ~pi0785 & ~new_n25514_;
  assign new_n25530_ = ~new_n25528_ & ~new_n25529_;
  assign new_n25531_ = ~pi0618 & ~new_n25530_;
  assign new_n25532_ = pi0618 & new_n25339_;
  assign new_n25533_ = ~pi1154 & ~new_n25532_;
  assign new_n25534_ = ~new_n25531_ & new_n25533_;
  assign new_n25535_ = ~pi0627 & ~new_n25408_;
  assign new_n25536_ = ~new_n25534_ & new_n25535_;
  assign new_n25537_ = pi0618 & ~new_n25530_;
  assign new_n25538_ = ~pi0618 & new_n25339_;
  assign new_n25539_ = pi1154 & ~new_n25538_;
  assign new_n25540_ = ~new_n25537_ & new_n25539_;
  assign new_n25541_ = pi0627 & ~new_n25412_;
  assign new_n25542_ = ~new_n25540_ & new_n25541_;
  assign new_n25543_ = ~new_n25536_ & ~new_n25542_;
  assign new_n25544_ = pi0781 & ~new_n25543_;
  assign new_n25545_ = ~pi0781 & ~new_n25530_;
  assign new_n25546_ = ~new_n25544_ & ~new_n25545_;
  assign new_n25547_ = pi0619 & ~new_n25546_;
  assign new_n25548_ = ~pi0619 & ~new_n25342_;
  assign new_n25549_ = pi1159 & ~new_n25548_;
  assign new_n25550_ = ~new_n25547_ & new_n25549_;
  assign new_n25551_ = pi0648 & ~new_n25424_;
  assign new_n25552_ = ~new_n25550_ & new_n25551_;
  assign new_n25553_ = ~pi0619 & ~new_n25546_;
  assign new_n25554_ = pi0619 & ~new_n25342_;
  assign new_n25555_ = ~pi1159 & ~new_n25554_;
  assign new_n25556_ = ~new_n25553_ & new_n25555_;
  assign new_n25557_ = ~pi0648 & ~new_n25420_;
  assign new_n25558_ = ~new_n25556_ & new_n25557_;
  assign new_n25559_ = pi0789 & ~new_n25558_;
  assign new_n25560_ = ~new_n25552_ & new_n25559_;
  assign new_n25561_ = ~pi0789 & new_n25546_;
  assign new_n25562_ = new_n17969_ & ~new_n25561_;
  assign new_n25563_ = ~new_n25560_ & new_n25562_;
  assign new_n25564_ = pi0626 & ~new_n25427_;
  assign new_n25565_ = ~pi0626 & ~new_n25311_;
  assign new_n25566_ = new_n17731_ & ~new_n25565_;
  assign new_n25567_ = ~new_n25564_ & new_n25566_;
  assign new_n25568_ = new_n17856_ & new_n25344_;
  assign new_n25569_ = ~pi0626 & ~new_n25427_;
  assign new_n25570_ = pi0626 & ~new_n25311_;
  assign new_n25571_ = new_n17732_ & ~new_n25570_;
  assign new_n25572_ = ~new_n25569_ & new_n25571_;
  assign new_n25573_ = ~new_n25568_ & ~new_n25572_;
  assign new_n25574_ = ~new_n25567_ & new_n25573_;
  assign new_n25575_ = pi0788 & ~new_n25574_;
  assign new_n25576_ = ~new_n20364_ & ~new_n25575_;
  assign new_n25577_ = ~new_n25563_ & new_n25576_;
  assign new_n25578_ = ~new_n25462_ & ~new_n25577_;
  assign new_n25579_ = ~new_n20360_ & ~new_n25578_;
  assign new_n25580_ = ~new_n20556_ & new_n25433_;
  assign new_n25581_ = new_n17802_ & ~new_n25362_;
  assign new_n25582_ = new_n17801_ & ~new_n25366_;
  assign new_n25583_ = ~new_n25581_ & ~new_n25582_;
  assign new_n25584_ = ~new_n25580_ & new_n25583_;
  assign new_n25585_ = pi0787 & ~new_n25584_;
  assign new_n25586_ = ~new_n25579_ & ~new_n25585_;
  assign new_n25587_ = ~new_n25456_ & new_n25586_;
  assign new_n25588_ = ~new_n25452_ & ~new_n25587_;
  assign new_n25589_ = ~po1038 & ~new_n25588_;
  assign new_n25590_ = ~pi0178 & po1038;
  assign new_n25591_ = ~pi0832 & ~new_n25590_;
  assign new_n25592_ = ~new_n25589_ & new_n25591_;
  assign po0335 = ~new_n25310_ & ~new_n25592_;
  assign new_n25594_ = pi0179 & ~new_n3272_;
  assign new_n25595_ = ~pi0179 & ~new_n17431_;
  assign new_n25596_ = new_n18093_ & ~new_n25595_;
  assign new_n25597_ = ~pi0179 & new_n16810_;
  assign new_n25598_ = pi0179 & new_n16928_;
  assign new_n25599_ = pi0039 & ~new_n25598_;
  assign new_n25600_ = ~new_n25597_ & new_n25599_;
  assign new_n25601_ = pi0179 & new_n17178_;
  assign new_n25602_ = ~pi0179 & new_n17217_;
  assign new_n25603_ = ~pi0039 & ~new_n25602_;
  assign new_n25604_ = ~new_n25601_ & new_n25603_;
  assign new_n25605_ = ~new_n25600_ & ~new_n25604_;
  assign new_n25606_ = ~pi0038 & ~new_n25605_;
  assign new_n25607_ = ~new_n25596_ & ~new_n25606_;
  assign new_n25608_ = pi0741 & ~new_n25607_;
  assign new_n25609_ = pi0179 & new_n19406_;
  assign new_n25610_ = ~pi0179 & ~new_n19414_;
  assign new_n25611_ = ~pi0741 & ~new_n25610_;
  assign new_n25612_ = ~new_n25609_ & new_n25611_;
  assign new_n25613_ = ~pi0724 & ~new_n25612_;
  assign new_n25614_ = ~new_n25608_ & new_n25613_;
  assign new_n25615_ = ~pi0741 & ~new_n24446_;
  assign new_n25616_ = pi0179 & ~new_n25615_;
  assign new_n25617_ = ~pi0179 & ~pi0741;
  assign new_n25618_ = ~new_n19370_ & new_n25617_;
  assign new_n25619_ = new_n19376_ & new_n25618_;
  assign new_n25620_ = ~new_n25616_ & ~new_n25619_;
  assign new_n25621_ = ~new_n21674_ & new_n25620_;
  assign new_n25622_ = pi0724 & new_n25621_;
  assign new_n25623_ = new_n3272_ & ~new_n25622_;
  assign new_n25624_ = ~new_n25614_ & new_n25623_;
  assign new_n25625_ = ~new_n25594_ & ~new_n25624_;
  assign new_n25626_ = ~pi0625 & new_n25625_;
  assign new_n25627_ = new_n3272_ & ~new_n25621_;
  assign new_n25628_ = ~new_n25594_ & ~new_n25627_;
  assign new_n25629_ = pi0625 & new_n25628_;
  assign new_n25630_ = ~pi1153 & ~new_n25629_;
  assign new_n25631_ = ~new_n25626_ & new_n25630_;
  assign new_n25632_ = ~pi0179 & ~new_n17558_;
  assign new_n25633_ = ~pi0724 & new_n3272_;
  assign new_n25634_ = new_n25632_ & ~new_n25633_;
  assign new_n25635_ = ~pi0179 & new_n18124_;
  assign new_n25636_ = pi0179 & ~new_n18128_;
  assign new_n25637_ = ~pi0038 & ~new_n25636_;
  assign new_n25638_ = new_n3272_ & ~new_n25637_;
  assign new_n25639_ = ~new_n25635_ & ~new_n25638_;
  assign new_n25640_ = new_n17544_ & ~new_n25595_;
  assign new_n25641_ = ~pi0724 & ~new_n25640_;
  assign new_n25642_ = ~new_n25639_ & new_n25641_;
  assign new_n25643_ = ~new_n25634_ & ~new_n25642_;
  assign new_n25644_ = pi0625 & ~new_n25643_;
  assign new_n25645_ = ~pi0625 & new_n25632_;
  assign new_n25646_ = pi1153 & ~new_n25645_;
  assign new_n25647_ = ~new_n25644_ & new_n25646_;
  assign new_n25648_ = ~pi0608 & ~new_n25647_;
  assign new_n25649_ = ~new_n25631_ & new_n25648_;
  assign new_n25650_ = pi0625 & new_n25625_;
  assign new_n25651_ = ~pi0625 & new_n25628_;
  assign new_n25652_ = pi1153 & ~new_n25651_;
  assign new_n25653_ = ~new_n25650_ & new_n25652_;
  assign new_n25654_ = ~pi0625 & ~new_n25643_;
  assign new_n25655_ = pi0625 & new_n25632_;
  assign new_n25656_ = ~pi1153 & ~new_n25655_;
  assign new_n25657_ = ~new_n25654_ & new_n25656_;
  assign new_n25658_ = pi0608 & ~new_n25657_;
  assign new_n25659_ = ~new_n25653_ & new_n25658_;
  assign new_n25660_ = ~new_n25649_ & ~new_n25659_;
  assign new_n25661_ = pi0778 & ~new_n25660_;
  assign new_n25662_ = ~pi0778 & new_n25625_;
  assign new_n25663_ = ~new_n25661_ & ~new_n25662_;
  assign new_n25664_ = ~pi0609 & ~new_n25663_;
  assign new_n25665_ = ~pi0778 & new_n25643_;
  assign new_n25666_ = ~new_n25647_ & ~new_n25657_;
  assign new_n25667_ = pi0778 & ~new_n25666_;
  assign new_n25668_ = ~new_n25665_ & ~new_n25667_;
  assign new_n25669_ = pi0609 & new_n25668_;
  assign new_n25670_ = ~pi1155 & ~new_n25669_;
  assign new_n25671_ = ~new_n25664_ & new_n25670_;
  assign new_n25672_ = ~new_n17591_ & ~new_n25632_;
  assign new_n25673_ = ~new_n17590_ & ~new_n25628_;
  assign new_n25674_ = pi0609 & new_n25673_;
  assign new_n25675_ = ~new_n25672_ & ~new_n25674_;
  assign new_n25676_ = pi1155 & ~new_n25675_;
  assign new_n25677_ = ~pi0660 & ~new_n25676_;
  assign new_n25678_ = ~new_n25671_ & new_n25677_;
  assign new_n25679_ = pi0609 & ~new_n25663_;
  assign new_n25680_ = ~pi0609 & new_n25668_;
  assign new_n25681_ = pi1155 & ~new_n25680_;
  assign new_n25682_ = ~new_n25679_ & new_n25681_;
  assign new_n25683_ = ~new_n17603_ & ~new_n25632_;
  assign new_n25684_ = ~pi0609 & new_n25673_;
  assign new_n25685_ = ~new_n25683_ & ~new_n25684_;
  assign new_n25686_ = ~pi1155 & ~new_n25685_;
  assign new_n25687_ = pi0660 & ~new_n25686_;
  assign new_n25688_ = ~new_n25682_ & new_n25687_;
  assign new_n25689_ = ~new_n25678_ & ~new_n25688_;
  assign new_n25690_ = pi0785 & ~new_n25689_;
  assign new_n25691_ = ~pi0785 & ~new_n25663_;
  assign new_n25692_ = ~new_n25690_ & ~new_n25691_;
  assign new_n25693_ = ~pi0618 & ~new_n25692_;
  assign new_n25694_ = ~new_n17618_ & ~new_n25668_;
  assign new_n25695_ = new_n17618_ & ~new_n25632_;
  assign new_n25696_ = ~new_n25694_ & ~new_n25695_;
  assign new_n25697_ = pi0618 & new_n25696_;
  assign new_n25698_ = ~pi1154 & ~new_n25697_;
  assign new_n25699_ = ~new_n25693_ & new_n25698_;
  assign new_n25700_ = new_n17590_ & ~new_n25632_;
  assign new_n25701_ = ~new_n25673_ & ~new_n25700_;
  assign new_n25702_ = ~pi0785 & ~new_n25701_;
  assign new_n25703_ = ~new_n25676_ & ~new_n25686_;
  assign new_n25704_ = pi0785 & ~new_n25703_;
  assign new_n25705_ = ~new_n25702_ & ~new_n25704_;
  assign new_n25706_ = pi0618 & new_n25705_;
  assign new_n25707_ = ~pi0618 & new_n25632_;
  assign new_n25708_ = pi1154 & ~new_n25707_;
  assign new_n25709_ = ~new_n25706_ & new_n25708_;
  assign new_n25710_ = ~pi0627 & ~new_n25709_;
  assign new_n25711_ = ~new_n25699_ & new_n25710_;
  assign new_n25712_ = pi0618 & ~new_n25692_;
  assign new_n25713_ = ~pi0618 & new_n25696_;
  assign new_n25714_ = pi1154 & ~new_n25713_;
  assign new_n25715_ = ~new_n25712_ & new_n25714_;
  assign new_n25716_ = ~pi0618 & new_n25705_;
  assign new_n25717_ = pi0618 & new_n25632_;
  assign new_n25718_ = ~pi1154 & ~new_n25717_;
  assign new_n25719_ = ~new_n25716_ & new_n25718_;
  assign new_n25720_ = pi0627 & ~new_n25719_;
  assign new_n25721_ = ~new_n25715_ & new_n25720_;
  assign new_n25722_ = ~new_n25711_ & ~new_n25721_;
  assign new_n25723_ = pi0781 & ~new_n25722_;
  assign new_n25724_ = ~pi0781 & ~new_n25692_;
  assign new_n25725_ = ~new_n25723_ & ~new_n25724_;
  assign new_n25726_ = ~pi0619 & ~new_n25725_;
  assign new_n25727_ = ~new_n17655_ & new_n25696_;
  assign new_n25728_ = new_n17655_ & new_n25632_;
  assign new_n25729_ = ~new_n25727_ & ~new_n25728_;
  assign new_n25730_ = pi0619 & ~new_n25729_;
  assign new_n25731_ = ~pi1159 & ~new_n25730_;
  assign new_n25732_ = ~new_n25726_ & new_n25731_;
  assign new_n25733_ = ~pi0781 & ~new_n25705_;
  assign new_n25734_ = ~new_n25709_ & ~new_n25719_;
  assign new_n25735_ = pi0781 & ~new_n25734_;
  assign new_n25736_ = ~new_n25733_ & ~new_n25735_;
  assign new_n25737_ = pi0619 & new_n25736_;
  assign new_n25738_ = ~pi0619 & new_n25632_;
  assign new_n25739_ = pi1159 & ~new_n25738_;
  assign new_n25740_ = ~new_n25737_ & new_n25739_;
  assign new_n25741_ = ~pi0648 & ~new_n25740_;
  assign new_n25742_ = ~new_n25732_ & new_n25741_;
  assign new_n25743_ = pi0619 & ~new_n25725_;
  assign new_n25744_ = ~pi0619 & ~new_n25729_;
  assign new_n25745_ = pi1159 & ~new_n25744_;
  assign new_n25746_ = ~new_n25743_ & new_n25745_;
  assign new_n25747_ = ~pi0619 & new_n25736_;
  assign new_n25748_ = pi0619 & new_n25632_;
  assign new_n25749_ = ~pi1159 & ~new_n25748_;
  assign new_n25750_ = ~new_n25747_ & new_n25749_;
  assign new_n25751_ = pi0648 & ~new_n25750_;
  assign new_n25752_ = ~new_n25746_ & new_n25751_;
  assign new_n25753_ = ~new_n25742_ & ~new_n25752_;
  assign new_n25754_ = pi0789 & ~new_n25753_;
  assign new_n25755_ = ~pi0789 & ~new_n25725_;
  assign new_n25756_ = ~new_n25754_ & ~new_n25755_;
  assign new_n25757_ = ~pi0788 & new_n25756_;
  assign new_n25758_ = ~pi0626 & new_n25756_;
  assign new_n25759_ = new_n17691_ & ~new_n25632_;
  assign new_n25760_ = ~new_n17691_ & new_n25729_;
  assign new_n25761_ = ~new_n25759_ & ~new_n25760_;
  assign new_n25762_ = pi0626 & ~new_n25761_;
  assign new_n25763_ = ~pi0641 & ~new_n25762_;
  assign new_n25764_ = ~new_n25758_ & new_n25763_;
  assign new_n25765_ = ~pi0789 & ~new_n25736_;
  assign new_n25766_ = ~new_n25740_ & ~new_n25750_;
  assign new_n25767_ = pi0789 & ~new_n25766_;
  assign new_n25768_ = ~new_n25765_ & ~new_n25767_;
  assign new_n25769_ = ~pi0626 & ~new_n25768_;
  assign new_n25770_ = pi0626 & ~new_n25632_;
  assign new_n25771_ = pi0641 & ~new_n25770_;
  assign new_n25772_ = ~new_n25769_ & new_n25771_;
  assign new_n25773_ = ~pi1158 & ~new_n25772_;
  assign new_n25774_ = ~new_n25764_ & new_n25773_;
  assign new_n25775_ = pi0626 & new_n25756_;
  assign new_n25776_ = ~pi0626 & ~new_n25761_;
  assign new_n25777_ = pi0641 & ~new_n25776_;
  assign new_n25778_ = ~new_n25775_ & new_n25777_;
  assign new_n25779_ = pi0626 & ~new_n25768_;
  assign new_n25780_ = ~pi0626 & ~new_n25632_;
  assign new_n25781_ = ~pi0641 & ~new_n25780_;
  assign new_n25782_ = ~new_n25779_ & new_n25781_;
  assign new_n25783_ = pi1158 & ~new_n25782_;
  assign new_n25784_ = ~new_n25778_ & new_n25783_;
  assign new_n25785_ = ~new_n25774_ & ~new_n25784_;
  assign new_n25786_ = pi0788 & ~new_n25785_;
  assign new_n25787_ = ~new_n25757_ & ~new_n25786_;
  assign new_n25788_ = ~pi0628 & new_n25787_;
  assign new_n25789_ = ~new_n17968_ & new_n25768_;
  assign new_n25790_ = new_n17968_ & new_n25632_;
  assign new_n25791_ = ~new_n25789_ & ~new_n25790_;
  assign new_n25792_ = pi0628 & ~new_n25791_;
  assign new_n25793_ = ~pi1156 & ~new_n25792_;
  assign new_n25794_ = ~new_n25788_ & new_n25793_;
  assign new_n25795_ = ~new_n17734_ & new_n25761_;
  assign new_n25796_ = new_n17734_ & new_n25632_;
  assign new_n25797_ = ~new_n25795_ & ~new_n25796_;
  assign new_n25798_ = pi0628 & ~new_n25797_;
  assign new_n25799_ = ~pi0628 & new_n25632_;
  assign new_n25800_ = pi1156 & ~new_n25799_;
  assign new_n25801_ = ~new_n25798_ & new_n25800_;
  assign new_n25802_ = ~pi0629 & ~new_n25801_;
  assign new_n25803_ = ~new_n25794_ & new_n25802_;
  assign new_n25804_ = pi0628 & new_n25787_;
  assign new_n25805_ = ~pi0628 & ~new_n25791_;
  assign new_n25806_ = pi1156 & ~new_n25805_;
  assign new_n25807_ = ~new_n25804_ & new_n25806_;
  assign new_n25808_ = ~pi0628 & ~new_n25797_;
  assign new_n25809_ = pi0628 & new_n25632_;
  assign new_n25810_ = ~pi1156 & ~new_n25809_;
  assign new_n25811_ = ~new_n25808_ & new_n25810_;
  assign new_n25812_ = pi0629 & ~new_n25811_;
  assign new_n25813_ = ~new_n25807_ & new_n25812_;
  assign new_n25814_ = ~new_n25803_ & ~new_n25813_;
  assign new_n25815_ = pi0792 & ~new_n25814_;
  assign new_n25816_ = ~pi0792 & new_n25787_;
  assign new_n25817_ = ~new_n25815_ & ~new_n25816_;
  assign new_n25818_ = ~pi0647 & ~new_n25817_;
  assign new_n25819_ = ~new_n17762_ & ~new_n25791_;
  assign new_n25820_ = new_n17762_ & new_n25632_;
  assign new_n25821_ = ~new_n25819_ & ~new_n25820_;
  assign new_n25822_ = pi0647 & ~new_n25821_;
  assign new_n25823_ = ~pi1157 & ~new_n25822_;
  assign new_n25824_ = ~new_n25818_ & new_n25823_;
  assign new_n25825_ = ~pi0792 & new_n25797_;
  assign new_n25826_ = ~new_n25801_ & ~new_n25811_;
  assign new_n25827_ = pi0792 & ~new_n25826_;
  assign new_n25828_ = ~new_n25825_ & ~new_n25827_;
  assign new_n25829_ = pi0647 & new_n25828_;
  assign new_n25830_ = ~pi0647 & new_n25632_;
  assign new_n25831_ = pi1157 & ~new_n25830_;
  assign new_n25832_ = ~new_n25829_ & new_n25831_;
  assign new_n25833_ = ~pi0630 & ~new_n25832_;
  assign new_n25834_ = ~new_n25824_ & new_n25833_;
  assign new_n25835_ = pi0647 & ~new_n25817_;
  assign new_n25836_ = ~pi0647 & ~new_n25821_;
  assign new_n25837_ = pi1157 & ~new_n25836_;
  assign new_n25838_ = ~new_n25835_ & new_n25837_;
  assign new_n25839_ = ~pi0647 & new_n25828_;
  assign new_n25840_ = pi0647 & new_n25632_;
  assign new_n25841_ = ~pi1157 & ~new_n25840_;
  assign new_n25842_ = ~new_n25839_ & new_n25841_;
  assign new_n25843_ = pi0630 & ~new_n25842_;
  assign new_n25844_ = ~new_n25838_ & new_n25843_;
  assign new_n25845_ = ~new_n25834_ & ~new_n25844_;
  assign new_n25846_ = pi0787 & ~new_n25845_;
  assign new_n25847_ = ~pi0787 & ~new_n25817_;
  assign new_n25848_ = ~new_n25846_ & ~new_n25847_;
  assign new_n25849_ = ~pi0644 & ~new_n25848_;
  assign new_n25850_ = ~pi0787 & ~new_n25828_;
  assign new_n25851_ = ~new_n25832_ & ~new_n25842_;
  assign new_n25852_ = pi0787 & ~new_n25851_;
  assign new_n25853_ = ~new_n25850_ & ~new_n25852_;
  assign new_n25854_ = pi0644 & new_n25853_;
  assign new_n25855_ = ~pi0715 & ~new_n25854_;
  assign new_n25856_ = ~new_n25849_ & new_n25855_;
  assign new_n25857_ = new_n17804_ & ~new_n25632_;
  assign new_n25858_ = ~new_n17804_ & new_n25821_;
  assign new_n25859_ = ~new_n25857_ & ~new_n25858_;
  assign new_n25860_ = ~pi0644 & new_n25859_;
  assign new_n25861_ = pi0644 & new_n25632_;
  assign new_n25862_ = pi0715 & ~new_n25861_;
  assign new_n25863_ = ~new_n25860_ & new_n25862_;
  assign new_n25864_ = ~pi1160 & ~new_n25863_;
  assign new_n25865_ = ~new_n25856_ & new_n25864_;
  assign new_n25866_ = pi0644 & ~new_n25848_;
  assign new_n25867_ = ~pi0644 & new_n25853_;
  assign new_n25868_ = pi0715 & ~new_n25867_;
  assign new_n25869_ = ~new_n25866_ & new_n25868_;
  assign new_n25870_ = pi0644 & new_n25859_;
  assign new_n25871_ = ~pi0644 & new_n25632_;
  assign new_n25872_ = ~pi0715 & ~new_n25871_;
  assign new_n25873_ = ~new_n25870_ & new_n25872_;
  assign new_n25874_ = pi1160 & ~new_n25873_;
  assign new_n25875_ = ~new_n25869_ & new_n25874_;
  assign new_n25876_ = pi0790 & ~new_n25875_;
  assign new_n25877_ = ~new_n25865_ & new_n25876_;
  assign new_n25878_ = ~pi0790 & new_n25848_;
  assign new_n25879_ = ~po1038 & ~new_n25878_;
  assign new_n25880_ = ~new_n25877_ & new_n25879_;
  assign new_n25881_ = ~pi0179 & po1038;
  assign new_n25882_ = ~pi0832 & ~new_n25881_;
  assign new_n25883_ = ~new_n25880_ & new_n25882_;
  assign new_n25884_ = ~pi0179 & ~new_n2754_;
  assign new_n25885_ = ~pi0741 & new_n16913_;
  assign new_n25886_ = ~new_n25884_ & ~new_n25885_;
  assign new_n25887_ = ~new_n17858_ & ~new_n25886_;
  assign new_n25888_ = ~pi0785 & ~new_n25887_;
  assign new_n25889_ = ~new_n17863_ & ~new_n25886_;
  assign new_n25890_ = pi1155 & ~new_n25889_;
  assign new_n25891_ = ~new_n17866_ & new_n25887_;
  assign new_n25892_ = ~pi1155 & ~new_n25891_;
  assign new_n25893_ = ~new_n25890_ & ~new_n25892_;
  assign new_n25894_ = pi0785 & ~new_n25893_;
  assign new_n25895_ = ~new_n25888_ & ~new_n25894_;
  assign new_n25896_ = ~pi0781 & ~new_n25895_;
  assign new_n25897_ = ~new_n17873_ & new_n25895_;
  assign new_n25898_ = pi1154 & ~new_n25897_;
  assign new_n25899_ = ~new_n17876_ & new_n25895_;
  assign new_n25900_ = ~pi1154 & ~new_n25899_;
  assign new_n25901_ = ~new_n25898_ & ~new_n25900_;
  assign new_n25902_ = pi0781 & ~new_n25901_;
  assign new_n25903_ = ~new_n25896_ & ~new_n25902_;
  assign new_n25904_ = ~pi0789 & ~new_n25903_;
  assign new_n25905_ = pi0619 & new_n25903_;
  assign new_n25906_ = ~pi0619 & new_n25884_;
  assign new_n25907_ = pi1159 & ~new_n25906_;
  assign new_n25908_ = ~new_n25905_ & new_n25907_;
  assign new_n25909_ = ~pi0619 & new_n25903_;
  assign new_n25910_ = pi0619 & new_n25884_;
  assign new_n25911_ = ~pi1159 & ~new_n25910_;
  assign new_n25912_ = ~new_n25909_ & new_n25911_;
  assign new_n25913_ = ~new_n25908_ & ~new_n25912_;
  assign new_n25914_ = pi0789 & ~new_n25913_;
  assign new_n25915_ = ~new_n25904_ & ~new_n25914_;
  assign new_n25916_ = ~new_n17968_ & new_n25915_;
  assign new_n25917_ = new_n17968_ & new_n25884_;
  assign new_n25918_ = ~new_n25916_ & ~new_n25917_;
  assign new_n25919_ = ~new_n17762_ & ~new_n25918_;
  assign new_n25920_ = new_n17762_ & new_n25884_;
  assign new_n25921_ = ~new_n25919_ & ~new_n25920_;
  assign new_n25922_ = ~new_n20556_ & new_n25921_;
  assign new_n25923_ = ~pi0724 & new_n16915_;
  assign new_n25924_ = ~new_n25884_ & ~new_n25923_;
  assign new_n25925_ = ~pi0778 & new_n25924_;
  assign new_n25926_ = ~pi0625 & new_n25923_;
  assign new_n25927_ = ~new_n25924_ & ~new_n25926_;
  assign new_n25928_ = pi1153 & ~new_n25927_;
  assign new_n25929_ = ~pi1153 & ~new_n25884_;
  assign new_n25930_ = ~new_n25926_ & new_n25929_;
  assign new_n25931_ = ~new_n25928_ & ~new_n25930_;
  assign new_n25932_ = pi0778 & ~new_n25931_;
  assign new_n25933_ = ~new_n25925_ & ~new_n25932_;
  assign new_n25934_ = ~new_n17844_ & new_n25933_;
  assign new_n25935_ = ~new_n17846_ & new_n25934_;
  assign new_n25936_ = ~new_n17848_ & new_n25935_;
  assign new_n25937_ = ~new_n17980_ & new_n25936_;
  assign new_n25938_ = ~new_n18011_ & new_n25937_;
  assign new_n25939_ = ~pi0647 & new_n25938_;
  assign new_n25940_ = pi0647 & new_n25884_;
  assign new_n25941_ = ~pi1157 & ~new_n25940_;
  assign new_n25942_ = ~new_n25939_ & new_n25941_;
  assign new_n25943_ = pi0630 & new_n25942_;
  assign new_n25944_ = pi0647 & ~new_n25938_;
  assign new_n25945_ = ~pi0647 & ~new_n25884_;
  assign new_n25946_ = ~new_n25944_ & ~new_n25945_;
  assign new_n25947_ = new_n17801_ & ~new_n25946_;
  assign new_n25948_ = ~new_n25943_ & ~new_n25947_;
  assign new_n25949_ = ~new_n25922_ & new_n25948_;
  assign new_n25950_ = pi0787 & ~new_n25949_;
  assign new_n25951_ = pi0626 & ~new_n25915_;
  assign new_n25952_ = ~pi0626 & ~new_n25884_;
  assign new_n25953_ = new_n17731_ & ~new_n25952_;
  assign new_n25954_ = ~new_n25951_ & new_n25953_;
  assign new_n25955_ = new_n17856_ & new_n25936_;
  assign new_n25956_ = ~pi0626 & ~new_n25915_;
  assign new_n25957_ = pi0626 & ~new_n25884_;
  assign new_n25958_ = new_n17732_ & ~new_n25957_;
  assign new_n25959_ = ~new_n25956_ & new_n25958_;
  assign new_n25960_ = ~new_n25955_ & ~new_n25959_;
  assign new_n25961_ = ~new_n25954_ & new_n25960_;
  assign new_n25962_ = pi0788 & ~new_n25961_;
  assign new_n25963_ = ~new_n16639_ & ~new_n25924_;
  assign new_n25964_ = pi0625 & new_n25963_;
  assign new_n25965_ = new_n25886_ & ~new_n25963_;
  assign new_n25966_ = ~new_n25964_ & ~new_n25965_;
  assign new_n25967_ = new_n25929_ & ~new_n25966_;
  assign new_n25968_ = ~pi0608 & ~new_n25928_;
  assign new_n25969_ = ~new_n25967_ & new_n25968_;
  assign new_n25970_ = pi1153 & new_n25886_;
  assign new_n25971_ = ~new_n25964_ & new_n25970_;
  assign new_n25972_ = pi0608 & ~new_n25930_;
  assign new_n25973_ = ~new_n25971_ & new_n25972_;
  assign new_n25974_ = ~new_n25969_ & ~new_n25973_;
  assign new_n25975_ = pi0778 & ~new_n25974_;
  assign new_n25976_ = ~pi0778 & ~new_n25965_;
  assign new_n25977_ = ~new_n25975_ & ~new_n25976_;
  assign new_n25978_ = ~pi0609 & ~new_n25977_;
  assign new_n25979_ = pi0609 & new_n25933_;
  assign new_n25980_ = ~pi1155 & ~new_n25979_;
  assign new_n25981_ = ~new_n25978_ & new_n25980_;
  assign new_n25982_ = ~pi0660 & ~new_n25890_;
  assign new_n25983_ = ~new_n25981_ & new_n25982_;
  assign new_n25984_ = pi0609 & ~new_n25977_;
  assign new_n25985_ = ~pi0609 & new_n25933_;
  assign new_n25986_ = pi1155 & ~new_n25985_;
  assign new_n25987_ = ~new_n25984_ & new_n25986_;
  assign new_n25988_ = pi0660 & ~new_n25892_;
  assign new_n25989_ = ~new_n25987_ & new_n25988_;
  assign new_n25990_ = ~new_n25983_ & ~new_n25989_;
  assign new_n25991_ = pi0785 & ~new_n25990_;
  assign new_n25992_ = ~pi0785 & ~new_n25977_;
  assign new_n25993_ = ~new_n25991_ & ~new_n25992_;
  assign new_n25994_ = ~pi0618 & ~new_n25993_;
  assign new_n25995_ = pi0618 & new_n25934_;
  assign new_n25996_ = ~pi1154 & ~new_n25995_;
  assign new_n25997_ = ~new_n25994_ & new_n25996_;
  assign new_n25998_ = ~pi0627 & ~new_n25898_;
  assign new_n25999_ = ~new_n25997_ & new_n25998_;
  assign new_n26000_ = pi0618 & ~new_n25993_;
  assign new_n26001_ = ~pi0618 & new_n25934_;
  assign new_n26002_ = pi1154 & ~new_n26001_;
  assign new_n26003_ = ~new_n26000_ & new_n26002_;
  assign new_n26004_ = pi0627 & ~new_n25900_;
  assign new_n26005_ = ~new_n26003_ & new_n26004_;
  assign new_n26006_ = ~new_n25999_ & ~new_n26005_;
  assign new_n26007_ = pi0781 & ~new_n26006_;
  assign new_n26008_ = ~pi0781 & ~new_n25993_;
  assign new_n26009_ = ~new_n26007_ & ~new_n26008_;
  assign new_n26010_ = pi0619 & ~new_n26009_;
  assign new_n26011_ = ~pi0619 & new_n25935_;
  assign new_n26012_ = pi1159 & ~new_n26011_;
  assign new_n26013_ = ~new_n26010_ & new_n26012_;
  assign new_n26014_ = pi0648 & ~new_n25912_;
  assign new_n26015_ = ~new_n26013_ & new_n26014_;
  assign new_n26016_ = ~pi0619 & ~new_n26009_;
  assign new_n26017_ = pi0619 & new_n25935_;
  assign new_n26018_ = ~pi1159 & ~new_n26017_;
  assign new_n26019_ = ~new_n26016_ & new_n26018_;
  assign new_n26020_ = ~pi0648 & ~new_n25908_;
  assign new_n26021_ = ~new_n26019_ & new_n26020_;
  assign new_n26022_ = pi0789 & ~new_n26021_;
  assign new_n26023_ = ~new_n26015_ & new_n26022_;
  assign new_n26024_ = ~pi0789 & new_n26009_;
  assign new_n26025_ = new_n17969_ & ~new_n26024_;
  assign new_n26026_ = ~new_n26023_ & new_n26025_;
  assign new_n26027_ = ~new_n25962_ & ~new_n26026_;
  assign new_n26028_ = ~new_n20364_ & ~new_n26027_;
  assign new_n26029_ = new_n18008_ & ~new_n25918_;
  assign new_n26030_ = new_n20851_ & new_n25937_;
  assign new_n26031_ = ~new_n26029_ & ~new_n26030_;
  assign new_n26032_ = ~pi0629 & ~new_n26031_;
  assign new_n26033_ = new_n20855_ & new_n25937_;
  assign new_n26034_ = new_n18007_ & ~new_n25918_;
  assign new_n26035_ = ~new_n26033_ & ~new_n26034_;
  assign new_n26036_ = pi0629 & ~new_n26035_;
  assign new_n26037_ = ~new_n26032_ & ~new_n26036_;
  assign new_n26038_ = pi0792 & ~new_n26037_;
  assign new_n26039_ = ~new_n20360_ & ~new_n26038_;
  assign new_n26040_ = ~new_n26028_ & new_n26039_;
  assign new_n26041_ = ~new_n25950_ & ~new_n26040_;
  assign new_n26042_ = pi0644 & new_n26041_;
  assign new_n26043_ = ~pi0787 & ~new_n25938_;
  assign new_n26044_ = pi1157 & ~new_n25946_;
  assign new_n26045_ = ~new_n25942_ & ~new_n26044_;
  assign new_n26046_ = pi0787 & ~new_n26045_;
  assign new_n26047_ = ~new_n26043_ & ~new_n26046_;
  assign new_n26048_ = ~pi0644 & new_n26047_;
  assign new_n26049_ = pi0715 & ~new_n26048_;
  assign new_n26050_ = ~new_n26042_ & new_n26049_;
  assign new_n26051_ = ~new_n17804_ & ~new_n25921_;
  assign new_n26052_ = new_n17804_ & new_n25884_;
  assign new_n26053_ = ~new_n26051_ & ~new_n26052_;
  assign new_n26054_ = pi0644 & ~new_n26053_;
  assign new_n26055_ = ~pi0644 & new_n25884_;
  assign new_n26056_ = ~pi0715 & ~new_n26055_;
  assign new_n26057_ = ~new_n26054_ & new_n26056_;
  assign new_n26058_ = pi1160 & ~new_n26057_;
  assign new_n26059_ = ~new_n26050_ & new_n26058_;
  assign new_n26060_ = ~pi0644 & new_n26041_;
  assign new_n26061_ = pi0644 & new_n26047_;
  assign new_n26062_ = ~pi0715 & ~new_n26061_;
  assign new_n26063_ = ~new_n26060_ & new_n26062_;
  assign new_n26064_ = ~pi0644 & ~new_n26053_;
  assign new_n26065_ = pi0644 & new_n25884_;
  assign new_n26066_ = pi0715 & ~new_n26065_;
  assign new_n26067_ = ~new_n26064_ & new_n26066_;
  assign new_n26068_ = ~pi1160 & ~new_n26067_;
  assign new_n26069_ = ~new_n26063_ & new_n26068_;
  assign new_n26070_ = ~new_n26059_ & ~new_n26069_;
  assign new_n26071_ = pi0790 & ~new_n26070_;
  assign new_n26072_ = ~pi0790 & new_n26041_;
  assign new_n26073_ = pi0832 & ~new_n26072_;
  assign new_n26074_ = ~new_n26071_ & new_n26073_;
  assign po0336 = ~new_n25883_ & ~new_n26074_;
  assign new_n26076_ = ~pi0180 & ~new_n2754_;
  assign new_n26077_ = ~pi0753 & new_n16913_;
  assign new_n26078_ = ~new_n26076_ & ~new_n26077_;
  assign new_n26079_ = ~new_n17858_ & ~new_n26078_;
  assign new_n26080_ = ~pi0785 & ~new_n26079_;
  assign new_n26081_ = new_n17603_ & new_n26077_;
  assign new_n26082_ = new_n26079_ & ~new_n26081_;
  assign new_n26083_ = pi1155 & ~new_n26082_;
  assign new_n26084_ = ~pi1155 & ~new_n26076_;
  assign new_n26085_ = ~new_n26081_ & new_n26084_;
  assign new_n26086_ = ~new_n26083_ & ~new_n26085_;
  assign new_n26087_ = pi0785 & ~new_n26086_;
  assign new_n26088_ = ~new_n26080_ & ~new_n26087_;
  assign new_n26089_ = ~pi0781 & ~new_n26088_;
  assign new_n26090_ = ~new_n17873_ & new_n26088_;
  assign new_n26091_ = pi1154 & ~new_n26090_;
  assign new_n26092_ = ~new_n17876_ & new_n26088_;
  assign new_n26093_ = ~pi1154 & ~new_n26092_;
  assign new_n26094_ = ~new_n26091_ & ~new_n26093_;
  assign new_n26095_ = pi0781 & ~new_n26094_;
  assign new_n26096_ = ~new_n26089_ & ~new_n26095_;
  assign new_n26097_ = ~pi0789 & ~new_n26096_;
  assign new_n26098_ = ~new_n23057_ & new_n26096_;
  assign new_n26099_ = pi1159 & ~new_n26098_;
  assign new_n26100_ = ~new_n23060_ & new_n26096_;
  assign new_n26101_ = ~pi1159 & ~new_n26100_;
  assign new_n26102_ = ~new_n26099_ & ~new_n26101_;
  assign new_n26103_ = pi0789 & ~new_n26102_;
  assign new_n26104_ = ~new_n26097_ & ~new_n26103_;
  assign new_n26105_ = ~new_n17968_ & new_n26104_;
  assign new_n26106_ = new_n17968_ & new_n26076_;
  assign new_n26107_ = ~new_n26105_ & ~new_n26106_;
  assign new_n26108_ = ~new_n17762_ & ~new_n26107_;
  assign new_n26109_ = new_n17762_ & new_n26076_;
  assign new_n26110_ = ~new_n26108_ & ~new_n26109_;
  assign new_n26111_ = ~new_n20556_ & new_n26110_;
  assign new_n26112_ = ~pi0702 & new_n16915_;
  assign new_n26113_ = ~new_n26076_ & ~new_n26112_;
  assign new_n26114_ = ~pi0778 & ~new_n26113_;
  assign new_n26115_ = ~pi0625 & new_n26112_;
  assign new_n26116_ = ~new_n26113_ & ~new_n26115_;
  assign new_n26117_ = pi1153 & ~new_n26116_;
  assign new_n26118_ = ~pi1153 & ~new_n26076_;
  assign new_n26119_ = ~new_n26115_ & new_n26118_;
  assign new_n26120_ = pi0778 & ~new_n26119_;
  assign new_n26121_ = ~new_n26117_ & new_n26120_;
  assign new_n26122_ = ~new_n26114_ & ~new_n26121_;
  assign new_n26123_ = ~new_n17844_ & ~new_n26122_;
  assign new_n26124_ = ~new_n17846_ & new_n26123_;
  assign new_n26125_ = ~new_n17848_ & new_n26124_;
  assign new_n26126_ = ~new_n17980_ & new_n26125_;
  assign new_n26127_ = ~new_n18011_ & new_n26126_;
  assign new_n26128_ = ~pi0647 & new_n26127_;
  assign new_n26129_ = pi0647 & new_n26076_;
  assign new_n26130_ = ~pi1157 & ~new_n26129_;
  assign new_n26131_ = ~new_n26128_ & new_n26130_;
  assign new_n26132_ = pi0630 & new_n26131_;
  assign new_n26133_ = pi0647 & ~new_n26127_;
  assign new_n26134_ = ~pi0647 & ~new_n26076_;
  assign new_n26135_ = ~new_n26133_ & ~new_n26134_;
  assign new_n26136_ = new_n17801_ & ~new_n26135_;
  assign new_n26137_ = ~new_n26132_ & ~new_n26136_;
  assign new_n26138_ = ~new_n26111_ & new_n26137_;
  assign new_n26139_ = pi0787 & ~new_n26138_;
  assign new_n26140_ = pi0626 & ~new_n26104_;
  assign new_n26141_ = ~pi0626 & ~new_n26076_;
  assign new_n26142_ = new_n17731_ & ~new_n26141_;
  assign new_n26143_ = ~new_n26140_ & new_n26142_;
  assign new_n26144_ = new_n17856_ & new_n26125_;
  assign new_n26145_ = ~pi0626 & ~new_n26104_;
  assign new_n26146_ = pi0626 & ~new_n26076_;
  assign new_n26147_ = new_n17732_ & ~new_n26146_;
  assign new_n26148_ = ~new_n26145_ & new_n26147_;
  assign new_n26149_ = ~new_n26144_ & ~new_n26148_;
  assign new_n26150_ = ~new_n26143_ & new_n26149_;
  assign new_n26151_ = pi0788 & ~new_n26150_;
  assign new_n26152_ = ~new_n16639_ & ~new_n26113_;
  assign new_n26153_ = pi0625 & new_n26152_;
  assign new_n26154_ = new_n26078_ & ~new_n26152_;
  assign new_n26155_ = ~new_n26153_ & ~new_n26154_;
  assign new_n26156_ = new_n26118_ & ~new_n26155_;
  assign new_n26157_ = ~pi0608 & ~new_n26117_;
  assign new_n26158_ = ~new_n26156_ & new_n26157_;
  assign new_n26159_ = pi1153 & new_n26078_;
  assign new_n26160_ = ~new_n26153_ & new_n26159_;
  assign new_n26161_ = pi0608 & ~new_n26119_;
  assign new_n26162_ = ~new_n26160_ & new_n26161_;
  assign new_n26163_ = ~new_n26158_ & ~new_n26162_;
  assign new_n26164_ = pi0778 & ~new_n26163_;
  assign new_n26165_ = ~pi0778 & ~new_n26154_;
  assign new_n26166_ = ~new_n26164_ & ~new_n26165_;
  assign new_n26167_ = ~pi0609 & ~new_n26166_;
  assign new_n26168_ = pi0609 & ~new_n26122_;
  assign new_n26169_ = ~pi1155 & ~new_n26168_;
  assign new_n26170_ = ~new_n26167_ & new_n26169_;
  assign new_n26171_ = ~pi0660 & ~new_n26083_;
  assign new_n26172_ = ~new_n26170_ & new_n26171_;
  assign new_n26173_ = pi0609 & ~new_n26166_;
  assign new_n26174_ = ~pi0609 & ~new_n26122_;
  assign new_n26175_ = pi1155 & ~new_n26174_;
  assign new_n26176_ = ~new_n26173_ & new_n26175_;
  assign new_n26177_ = pi0660 & ~new_n26085_;
  assign new_n26178_ = ~new_n26176_ & new_n26177_;
  assign new_n26179_ = ~new_n26172_ & ~new_n26178_;
  assign new_n26180_ = pi0785 & ~new_n26179_;
  assign new_n26181_ = ~pi0785 & ~new_n26166_;
  assign new_n26182_ = ~new_n26180_ & ~new_n26181_;
  assign new_n26183_ = ~pi0618 & ~new_n26182_;
  assign new_n26184_ = pi0618 & new_n26123_;
  assign new_n26185_ = ~pi1154 & ~new_n26184_;
  assign new_n26186_ = ~new_n26183_ & new_n26185_;
  assign new_n26187_ = ~pi0627 & ~new_n26091_;
  assign new_n26188_ = ~new_n26186_ & new_n26187_;
  assign new_n26189_ = pi0618 & ~new_n26182_;
  assign new_n26190_ = ~pi0618 & new_n26123_;
  assign new_n26191_ = pi1154 & ~new_n26190_;
  assign new_n26192_ = ~new_n26189_ & new_n26191_;
  assign new_n26193_ = pi0627 & ~new_n26093_;
  assign new_n26194_ = ~new_n26192_ & new_n26193_;
  assign new_n26195_ = ~new_n26188_ & ~new_n26194_;
  assign new_n26196_ = pi0781 & ~new_n26195_;
  assign new_n26197_ = ~pi0781 & ~new_n26182_;
  assign new_n26198_ = ~new_n26196_ & ~new_n26197_;
  assign new_n26199_ = pi0619 & ~new_n26198_;
  assign new_n26200_ = ~pi0619 & new_n26124_;
  assign new_n26201_ = pi1159 & ~new_n26200_;
  assign new_n26202_ = ~new_n26199_ & new_n26201_;
  assign new_n26203_ = pi0648 & ~new_n26101_;
  assign new_n26204_ = ~new_n26202_ & new_n26203_;
  assign new_n26205_ = ~pi0619 & ~new_n26198_;
  assign new_n26206_ = pi0619 & new_n26124_;
  assign new_n26207_ = ~pi1159 & ~new_n26206_;
  assign new_n26208_ = ~new_n26205_ & new_n26207_;
  assign new_n26209_ = ~pi0648 & ~new_n26099_;
  assign new_n26210_ = ~new_n26208_ & new_n26209_;
  assign new_n26211_ = pi0789 & ~new_n26210_;
  assign new_n26212_ = ~new_n26204_ & new_n26211_;
  assign new_n26213_ = ~pi0789 & new_n26198_;
  assign new_n26214_ = new_n17969_ & ~new_n26213_;
  assign new_n26215_ = ~new_n26212_ & new_n26214_;
  assign new_n26216_ = ~new_n26151_ & ~new_n26215_;
  assign new_n26217_ = ~new_n20364_ & ~new_n26216_;
  assign new_n26218_ = new_n18008_ & ~new_n26107_;
  assign new_n26219_ = new_n20851_ & new_n26126_;
  assign new_n26220_ = ~new_n26218_ & ~new_n26219_;
  assign new_n26221_ = ~pi0629 & ~new_n26220_;
  assign new_n26222_ = new_n20855_ & new_n26126_;
  assign new_n26223_ = new_n18007_ & ~new_n26107_;
  assign new_n26224_ = ~new_n26222_ & ~new_n26223_;
  assign new_n26225_ = pi0629 & ~new_n26224_;
  assign new_n26226_ = ~new_n26221_ & ~new_n26225_;
  assign new_n26227_ = pi0792 & ~new_n26226_;
  assign new_n26228_ = ~new_n20360_ & ~new_n26227_;
  assign new_n26229_ = ~new_n26217_ & new_n26228_;
  assign new_n26230_ = ~new_n26139_ & ~new_n26229_;
  assign new_n26231_ = pi0644 & new_n26230_;
  assign new_n26232_ = ~pi0787 & ~new_n26127_;
  assign new_n26233_ = pi1157 & ~new_n26135_;
  assign new_n26234_ = ~new_n26131_ & ~new_n26233_;
  assign new_n26235_ = pi0787 & ~new_n26234_;
  assign new_n26236_ = ~new_n26232_ & ~new_n26235_;
  assign new_n26237_ = ~pi0644 & new_n26236_;
  assign new_n26238_ = pi0715 & ~new_n26237_;
  assign new_n26239_ = ~new_n26231_ & new_n26238_;
  assign new_n26240_ = ~new_n17804_ & ~new_n26110_;
  assign new_n26241_ = new_n17804_ & new_n26076_;
  assign new_n26242_ = ~new_n26240_ & ~new_n26241_;
  assign new_n26243_ = pi0644 & ~new_n26242_;
  assign new_n26244_ = ~pi0644 & new_n26076_;
  assign new_n26245_ = ~pi0715 & ~new_n26244_;
  assign new_n26246_ = ~new_n26243_ & new_n26245_;
  assign new_n26247_ = pi1160 & ~new_n26246_;
  assign new_n26248_ = ~new_n26239_ & new_n26247_;
  assign new_n26249_ = ~pi0644 & new_n26230_;
  assign new_n26250_ = pi0644 & new_n26236_;
  assign new_n26251_ = ~pi0715 & ~new_n26250_;
  assign new_n26252_ = ~new_n26249_ & new_n26251_;
  assign new_n26253_ = ~pi0644 & ~new_n26242_;
  assign new_n26254_ = pi0644 & new_n26076_;
  assign new_n26255_ = pi0715 & ~new_n26254_;
  assign new_n26256_ = ~new_n26253_ & new_n26255_;
  assign new_n26257_ = ~pi1160 & ~new_n26256_;
  assign new_n26258_ = ~new_n26252_ & new_n26257_;
  assign new_n26259_ = ~new_n26248_ & ~new_n26258_;
  assign new_n26260_ = pi0790 & ~new_n26259_;
  assign new_n26261_ = ~pi0790 & new_n26230_;
  assign new_n26262_ = pi0832 & ~new_n26261_;
  assign new_n26263_ = ~new_n26260_ & new_n26262_;
  assign new_n26264_ = ~pi0180 & ~new_n17558_;
  assign new_n26265_ = new_n17691_ & ~new_n26264_;
  assign new_n26266_ = ~pi0702 & new_n3272_;
  assign new_n26267_ = new_n26264_ & ~new_n26266_;
  assign new_n26268_ = pi0180 & ~new_n18128_;
  assign new_n26269_ = ~pi0038 & ~new_n26268_;
  assign new_n26270_ = new_n3272_ & ~new_n26269_;
  assign new_n26271_ = ~pi0180 & new_n18124_;
  assign new_n26272_ = ~new_n26270_ & ~new_n26271_;
  assign new_n26273_ = ~pi0180 & ~new_n17431_;
  assign new_n26274_ = new_n17544_ & ~new_n26273_;
  assign new_n26275_ = ~pi0702 & ~new_n26274_;
  assign new_n26276_ = ~new_n26272_ & new_n26275_;
  assign new_n26277_ = ~new_n26267_ & ~new_n26276_;
  assign new_n26278_ = ~pi0778 & new_n26277_;
  assign new_n26279_ = pi0625 & ~new_n26277_;
  assign new_n26280_ = ~pi0625 & new_n26264_;
  assign new_n26281_ = pi1153 & ~new_n26280_;
  assign new_n26282_ = ~new_n26279_ & new_n26281_;
  assign new_n26283_ = ~pi0625 & ~new_n26277_;
  assign new_n26284_ = pi0625 & new_n26264_;
  assign new_n26285_ = ~pi1153 & ~new_n26284_;
  assign new_n26286_ = ~new_n26283_ & new_n26285_;
  assign new_n26287_ = ~new_n26282_ & ~new_n26286_;
  assign new_n26288_ = pi0778 & ~new_n26287_;
  assign new_n26289_ = ~new_n26278_ & ~new_n26288_;
  assign new_n26290_ = ~new_n17618_ & ~new_n26289_;
  assign new_n26291_ = new_n17618_ & ~new_n26264_;
  assign new_n26292_ = ~new_n26290_ & ~new_n26291_;
  assign new_n26293_ = ~new_n17655_ & new_n26292_;
  assign new_n26294_ = new_n17655_ & new_n26264_;
  assign new_n26295_ = ~new_n26293_ & ~new_n26294_;
  assign new_n26296_ = ~new_n17691_ & new_n26295_;
  assign new_n26297_ = ~new_n26265_ & ~new_n26296_;
  assign new_n26298_ = ~new_n17734_ & new_n26297_;
  assign new_n26299_ = new_n17734_ & new_n26264_;
  assign new_n26300_ = ~new_n26298_ & ~new_n26299_;
  assign new_n26301_ = ~pi0792 & new_n26300_;
  assign new_n26302_ = pi0628 & ~new_n26300_;
  assign new_n26303_ = ~pi0628 & new_n26264_;
  assign new_n26304_ = pi1156 & ~new_n26303_;
  assign new_n26305_ = ~new_n26302_ & new_n26304_;
  assign new_n26306_ = ~pi0628 & ~new_n26300_;
  assign new_n26307_ = pi0628 & new_n26264_;
  assign new_n26308_ = ~pi1156 & ~new_n26307_;
  assign new_n26309_ = ~new_n26306_ & new_n26308_;
  assign new_n26310_ = ~new_n26305_ & ~new_n26309_;
  assign new_n26311_ = pi0792 & ~new_n26310_;
  assign new_n26312_ = ~new_n26301_ & ~new_n26311_;
  assign new_n26313_ = ~pi0647 & ~new_n26312_;
  assign new_n26314_ = pi0647 & ~new_n26264_;
  assign new_n26315_ = ~new_n26313_ & ~new_n26314_;
  assign new_n26316_ = ~pi1157 & new_n26315_;
  assign new_n26317_ = pi0647 & ~new_n26312_;
  assign new_n26318_ = ~pi0647 & ~new_n26264_;
  assign new_n26319_ = ~new_n26317_ & ~new_n26318_;
  assign new_n26320_ = pi1157 & new_n26319_;
  assign new_n26321_ = ~new_n26316_ & ~new_n26320_;
  assign new_n26322_ = pi0787 & ~new_n26321_;
  assign new_n26323_ = ~pi0787 & new_n26312_;
  assign new_n26324_ = ~new_n26322_ & ~new_n26323_;
  assign new_n26325_ = ~pi0644 & ~new_n26324_;
  assign new_n26326_ = pi0715 & ~new_n26325_;
  assign new_n26327_ = pi0180 & ~new_n3272_;
  assign new_n26328_ = pi0753 & new_n17347_;
  assign new_n26329_ = pi0180 & new_n17424_;
  assign new_n26330_ = ~new_n26328_ & ~new_n26329_;
  assign new_n26331_ = pi0039 & ~new_n26330_;
  assign new_n26332_ = ~pi0180 & ~pi0753;
  assign new_n26333_ = new_n17393_ & new_n26332_;
  assign new_n26334_ = pi0180 & pi0753;
  assign new_n26335_ = pi0180 & ~new_n17215_;
  assign new_n26336_ = ~new_n21758_ & ~new_n26335_;
  assign new_n26337_ = ~pi0039 & ~new_n26336_;
  assign new_n26338_ = ~new_n26334_ & ~new_n26337_;
  assign new_n26339_ = ~new_n26333_ & new_n26338_;
  assign new_n26340_ = ~new_n26331_ & new_n26339_;
  assign new_n26341_ = ~pi0038 & ~new_n26340_;
  assign new_n26342_ = ~pi0753 & new_n17433_;
  assign new_n26343_ = pi0038 & ~new_n26273_;
  assign new_n26344_ = ~new_n26342_ & new_n26343_;
  assign new_n26345_ = ~new_n26341_ & ~new_n26344_;
  assign new_n26346_ = new_n3272_ & ~new_n26345_;
  assign new_n26347_ = ~new_n26327_ & ~new_n26346_;
  assign new_n26348_ = ~new_n17590_ & ~new_n26347_;
  assign new_n26349_ = new_n17590_ & ~new_n26264_;
  assign new_n26350_ = ~new_n26348_ & ~new_n26349_;
  assign new_n26351_ = ~pi0785 & ~new_n26350_;
  assign new_n26352_ = ~new_n17591_ & ~new_n26264_;
  assign new_n26353_ = pi0609 & new_n26348_;
  assign new_n26354_ = ~new_n26352_ & ~new_n26353_;
  assign new_n26355_ = pi1155 & ~new_n26354_;
  assign new_n26356_ = ~new_n17603_ & ~new_n26264_;
  assign new_n26357_ = ~pi0609 & new_n26348_;
  assign new_n26358_ = ~new_n26356_ & ~new_n26357_;
  assign new_n26359_ = ~pi1155 & ~new_n26358_;
  assign new_n26360_ = ~new_n26355_ & ~new_n26359_;
  assign new_n26361_ = pi0785 & ~new_n26360_;
  assign new_n26362_ = ~new_n26351_ & ~new_n26361_;
  assign new_n26363_ = ~pi0781 & ~new_n26362_;
  assign new_n26364_ = pi0618 & new_n26362_;
  assign new_n26365_ = ~pi0618 & new_n26264_;
  assign new_n26366_ = pi1154 & ~new_n26365_;
  assign new_n26367_ = ~new_n26364_ & new_n26366_;
  assign new_n26368_ = ~pi0618 & new_n26362_;
  assign new_n26369_ = pi0618 & new_n26264_;
  assign new_n26370_ = ~pi1154 & ~new_n26369_;
  assign new_n26371_ = ~new_n26368_ & new_n26370_;
  assign new_n26372_ = ~new_n26367_ & ~new_n26371_;
  assign new_n26373_ = pi0781 & ~new_n26372_;
  assign new_n26374_ = ~new_n26363_ & ~new_n26373_;
  assign new_n26375_ = ~pi0789 & ~new_n26374_;
  assign new_n26376_ = pi0619 & new_n26374_;
  assign new_n26377_ = ~pi0619 & new_n26264_;
  assign new_n26378_ = pi1159 & ~new_n26377_;
  assign new_n26379_ = ~new_n26376_ & new_n26378_;
  assign new_n26380_ = ~pi0619 & new_n26374_;
  assign new_n26381_ = pi0619 & new_n26264_;
  assign new_n26382_ = ~pi1159 & ~new_n26381_;
  assign new_n26383_ = ~new_n26380_ & new_n26382_;
  assign new_n26384_ = ~new_n26379_ & ~new_n26383_;
  assign new_n26385_ = pi0789 & ~new_n26384_;
  assign new_n26386_ = ~new_n26375_ & ~new_n26385_;
  assign new_n26387_ = ~new_n17968_ & new_n26386_;
  assign new_n26388_ = new_n17968_ & new_n26264_;
  assign new_n26389_ = ~new_n26387_ & ~new_n26388_;
  assign new_n26390_ = ~new_n17762_ & ~new_n26389_;
  assign new_n26391_ = new_n17762_ & new_n26264_;
  assign new_n26392_ = ~new_n26390_ & ~new_n26391_;
  assign new_n26393_ = ~new_n17804_ & ~new_n26392_;
  assign new_n26394_ = new_n17804_ & new_n26264_;
  assign new_n26395_ = ~new_n26393_ & ~new_n26394_;
  assign new_n26396_ = pi0644 & ~new_n26395_;
  assign new_n26397_ = ~pi0644 & new_n26264_;
  assign new_n26398_ = ~pi0715 & ~new_n26397_;
  assign new_n26399_ = ~new_n26396_ & new_n26398_;
  assign new_n26400_ = pi1160 & ~new_n26399_;
  assign new_n26401_ = ~new_n26326_ & new_n26400_;
  assign new_n26402_ = pi0644 & ~new_n26324_;
  assign new_n26403_ = ~pi0715 & ~new_n26402_;
  assign new_n26404_ = ~pi0644 & ~new_n26395_;
  assign new_n26405_ = pi0644 & new_n26264_;
  assign new_n26406_ = pi0715 & ~new_n26405_;
  assign new_n26407_ = ~new_n26404_ & new_n26406_;
  assign new_n26408_ = ~pi1160 & ~new_n26407_;
  assign new_n26409_ = ~new_n26403_ & new_n26408_;
  assign new_n26410_ = ~new_n26401_ & ~new_n26409_;
  assign new_n26411_ = pi0790 & ~new_n26410_;
  assign new_n26412_ = pi0644 & new_n26400_;
  assign new_n26413_ = ~pi0644 & new_n26408_;
  assign new_n26414_ = pi0790 & ~new_n26413_;
  assign new_n26415_ = ~new_n26412_ & new_n26414_;
  assign new_n26416_ = ~new_n20567_ & new_n26389_;
  assign new_n26417_ = ~pi0629 & new_n26305_;
  assign new_n26418_ = pi0629 & new_n26309_;
  assign new_n26419_ = ~new_n26417_ & ~new_n26418_;
  assign new_n26420_ = ~new_n26416_ & new_n26419_;
  assign new_n26421_ = pi0792 & ~new_n26420_;
  assign new_n26422_ = pi0702 & new_n26345_;
  assign new_n26423_ = ~pi0180 & new_n16810_;
  assign new_n26424_ = pi0180 & new_n16928_;
  assign new_n26425_ = pi0753 & ~new_n26424_;
  assign new_n26426_ = ~new_n26423_ & new_n26425_;
  assign new_n26427_ = pi0180 & new_n17007_;
  assign new_n26428_ = ~pi0180 & ~new_n17074_;
  assign new_n26429_ = ~pi0753 & ~new_n26428_;
  assign new_n26430_ = ~new_n26427_ & new_n26429_;
  assign new_n26431_ = pi0039 & ~new_n26430_;
  assign new_n26432_ = ~new_n26426_ & new_n26431_;
  assign new_n26433_ = ~pi0180 & ~new_n17217_;
  assign new_n26434_ = pi0180 & ~new_n17178_;
  assign new_n26435_ = pi0753 & ~new_n26434_;
  assign new_n26436_ = ~new_n26433_ & new_n26435_;
  assign new_n26437_ = ~pi0180 & new_n17227_;
  assign new_n26438_ = pi0180 & new_n17234_;
  assign new_n26439_ = ~pi0753 & ~new_n26438_;
  assign new_n26440_ = ~new_n26437_ & new_n26439_;
  assign new_n26441_ = ~new_n26436_ & ~new_n26440_;
  assign new_n26442_ = ~pi0039 & ~new_n26441_;
  assign new_n26443_ = ~pi0038 & ~new_n26442_;
  assign new_n26444_ = ~new_n26432_ & new_n26443_;
  assign new_n26445_ = ~pi0753 & ~new_n17035_;
  assign new_n26446_ = new_n19383_ & ~new_n26445_;
  assign new_n26447_ = ~pi0180 & ~new_n26446_;
  assign new_n26448_ = ~new_n16916_ & ~new_n26077_;
  assign new_n26449_ = pi0180 & ~new_n26448_;
  assign new_n26450_ = new_n6257_ & new_n26449_;
  assign new_n26451_ = pi0038 & ~new_n26450_;
  assign new_n26452_ = ~new_n26447_ & new_n26451_;
  assign new_n26453_ = ~pi0702 & ~new_n26452_;
  assign new_n26454_ = ~new_n26444_ & new_n26453_;
  assign new_n26455_ = new_n3272_ & ~new_n26454_;
  assign new_n26456_ = ~new_n26422_ & new_n26455_;
  assign new_n26457_ = ~new_n26327_ & ~new_n26456_;
  assign new_n26458_ = ~pi0625 & new_n26457_;
  assign new_n26459_ = pi0625 & new_n26347_;
  assign new_n26460_ = ~pi1153 & ~new_n26459_;
  assign new_n26461_ = ~new_n26458_ & new_n26460_;
  assign new_n26462_ = ~pi0608 & ~new_n26282_;
  assign new_n26463_ = ~new_n26461_ & new_n26462_;
  assign new_n26464_ = pi0625 & new_n26457_;
  assign new_n26465_ = ~pi0625 & new_n26347_;
  assign new_n26466_ = pi1153 & ~new_n26465_;
  assign new_n26467_ = ~new_n26464_ & new_n26466_;
  assign new_n26468_ = pi0608 & ~new_n26286_;
  assign new_n26469_ = ~new_n26467_ & new_n26468_;
  assign new_n26470_ = ~new_n26463_ & ~new_n26469_;
  assign new_n26471_ = pi0778 & ~new_n26470_;
  assign new_n26472_ = ~pi0778 & new_n26457_;
  assign new_n26473_ = ~new_n26471_ & ~new_n26472_;
  assign new_n26474_ = ~pi0609 & ~new_n26473_;
  assign new_n26475_ = pi0609 & new_n26289_;
  assign new_n26476_ = ~pi1155 & ~new_n26475_;
  assign new_n26477_ = ~new_n26474_ & new_n26476_;
  assign new_n26478_ = ~pi0660 & ~new_n26355_;
  assign new_n26479_ = ~new_n26477_ & new_n26478_;
  assign new_n26480_ = pi0609 & ~new_n26473_;
  assign new_n26481_ = ~pi0609 & new_n26289_;
  assign new_n26482_ = pi1155 & ~new_n26481_;
  assign new_n26483_ = ~new_n26480_ & new_n26482_;
  assign new_n26484_ = pi0660 & ~new_n26359_;
  assign new_n26485_ = ~new_n26483_ & new_n26484_;
  assign new_n26486_ = ~new_n26479_ & ~new_n26485_;
  assign new_n26487_ = pi0785 & ~new_n26486_;
  assign new_n26488_ = ~pi0785 & ~new_n26473_;
  assign new_n26489_ = ~new_n26487_ & ~new_n26488_;
  assign new_n26490_ = ~pi0618 & ~new_n26489_;
  assign new_n26491_ = pi0618 & new_n26292_;
  assign new_n26492_ = ~pi1154 & ~new_n26491_;
  assign new_n26493_ = ~new_n26490_ & new_n26492_;
  assign new_n26494_ = ~pi0627 & ~new_n26367_;
  assign new_n26495_ = ~new_n26493_ & new_n26494_;
  assign new_n26496_ = pi0618 & ~new_n26489_;
  assign new_n26497_ = ~pi0618 & new_n26292_;
  assign new_n26498_ = pi1154 & ~new_n26497_;
  assign new_n26499_ = ~new_n26496_ & new_n26498_;
  assign new_n26500_ = pi0627 & ~new_n26371_;
  assign new_n26501_ = ~new_n26499_ & new_n26500_;
  assign new_n26502_ = ~new_n26495_ & ~new_n26501_;
  assign new_n26503_ = pi0781 & ~new_n26502_;
  assign new_n26504_ = ~pi0781 & ~new_n26489_;
  assign new_n26505_ = ~new_n26503_ & ~new_n26504_;
  assign new_n26506_ = pi0619 & ~new_n26505_;
  assign new_n26507_ = ~pi0619 & ~new_n26295_;
  assign new_n26508_ = pi1159 & ~new_n26507_;
  assign new_n26509_ = ~new_n26506_ & new_n26508_;
  assign new_n26510_ = pi0648 & ~new_n26383_;
  assign new_n26511_ = ~new_n26509_ & new_n26510_;
  assign new_n26512_ = ~pi0619 & ~new_n26505_;
  assign new_n26513_ = pi0619 & ~new_n26295_;
  assign new_n26514_ = ~pi1159 & ~new_n26513_;
  assign new_n26515_ = ~new_n26512_ & new_n26514_;
  assign new_n26516_ = ~pi0648 & ~new_n26379_;
  assign new_n26517_ = ~new_n26515_ & new_n26516_;
  assign new_n26518_ = pi0789 & ~new_n26517_;
  assign new_n26519_ = ~new_n26511_ & new_n26518_;
  assign new_n26520_ = ~pi0789 & new_n26505_;
  assign new_n26521_ = new_n17969_ & ~new_n26520_;
  assign new_n26522_ = ~new_n26519_ & new_n26521_;
  assign new_n26523_ = pi0626 & ~new_n26386_;
  assign new_n26524_ = ~pi0626 & ~new_n26264_;
  assign new_n26525_ = new_n17731_ & ~new_n26524_;
  assign new_n26526_ = ~new_n26523_ & new_n26525_;
  assign new_n26527_ = new_n17856_ & new_n26297_;
  assign new_n26528_ = ~pi0626 & ~new_n26386_;
  assign new_n26529_ = pi0626 & ~new_n26264_;
  assign new_n26530_ = new_n17732_ & ~new_n26529_;
  assign new_n26531_ = ~new_n26528_ & new_n26530_;
  assign new_n26532_ = ~new_n26527_ & ~new_n26531_;
  assign new_n26533_ = ~new_n26526_ & new_n26532_;
  assign new_n26534_ = pi0788 & ~new_n26533_;
  assign new_n26535_ = ~new_n20364_ & ~new_n26534_;
  assign new_n26536_ = ~new_n26522_ & new_n26535_;
  assign new_n26537_ = ~new_n26421_ & ~new_n26536_;
  assign new_n26538_ = ~new_n20360_ & ~new_n26537_;
  assign new_n26539_ = ~new_n20556_ & new_n26392_;
  assign new_n26540_ = new_n17802_ & ~new_n26315_;
  assign new_n26541_ = new_n17801_ & ~new_n26319_;
  assign new_n26542_ = ~new_n26540_ & ~new_n26541_;
  assign new_n26543_ = ~new_n26539_ & new_n26542_;
  assign new_n26544_ = pi0787 & ~new_n26543_;
  assign new_n26545_ = ~new_n26538_ & ~new_n26544_;
  assign new_n26546_ = ~new_n26415_ & new_n26545_;
  assign new_n26547_ = ~new_n26411_ & ~new_n26546_;
  assign new_n26548_ = ~po1038 & ~new_n26547_;
  assign new_n26549_ = ~pi0180 & po1038;
  assign new_n26550_ = ~pi0832 & ~new_n26549_;
  assign new_n26551_ = ~new_n26548_ & new_n26550_;
  assign po0337 = ~new_n26263_ & ~new_n26551_;
  assign new_n26553_ = ~pi0181 & ~new_n2754_;
  assign new_n26554_ = ~pi0754 & new_n16913_;
  assign new_n26555_ = ~new_n26553_ & ~new_n26554_;
  assign new_n26556_ = ~new_n17858_ & ~new_n26555_;
  assign new_n26557_ = ~pi0785 & ~new_n26556_;
  assign new_n26558_ = new_n17603_ & new_n26554_;
  assign new_n26559_ = new_n26556_ & ~new_n26558_;
  assign new_n26560_ = pi1155 & ~new_n26559_;
  assign new_n26561_ = ~pi1155 & ~new_n26553_;
  assign new_n26562_ = ~new_n26558_ & new_n26561_;
  assign new_n26563_ = ~new_n26560_ & ~new_n26562_;
  assign new_n26564_ = pi0785 & ~new_n26563_;
  assign new_n26565_ = ~new_n26557_ & ~new_n26564_;
  assign new_n26566_ = ~pi0781 & ~new_n26565_;
  assign new_n26567_ = ~new_n17873_ & new_n26565_;
  assign new_n26568_ = pi1154 & ~new_n26567_;
  assign new_n26569_ = ~new_n17876_ & new_n26565_;
  assign new_n26570_ = ~pi1154 & ~new_n26569_;
  assign new_n26571_ = ~new_n26568_ & ~new_n26570_;
  assign new_n26572_ = pi0781 & ~new_n26571_;
  assign new_n26573_ = ~new_n26566_ & ~new_n26572_;
  assign new_n26574_ = ~pi0789 & ~new_n26573_;
  assign new_n26575_ = ~new_n23057_ & new_n26573_;
  assign new_n26576_ = pi1159 & ~new_n26575_;
  assign new_n26577_ = ~new_n23060_ & new_n26573_;
  assign new_n26578_ = ~pi1159 & ~new_n26577_;
  assign new_n26579_ = ~new_n26576_ & ~new_n26578_;
  assign new_n26580_ = pi0789 & ~new_n26579_;
  assign new_n26581_ = ~new_n26574_ & ~new_n26580_;
  assign new_n26582_ = ~new_n17968_ & new_n26581_;
  assign new_n26583_ = new_n17968_ & new_n26553_;
  assign new_n26584_ = ~new_n26582_ & ~new_n26583_;
  assign new_n26585_ = ~new_n17762_ & ~new_n26584_;
  assign new_n26586_ = new_n17762_ & new_n26553_;
  assign new_n26587_ = ~new_n26585_ & ~new_n26586_;
  assign new_n26588_ = ~new_n20556_ & new_n26587_;
  assign new_n26589_ = ~pi0709 & new_n16915_;
  assign new_n26590_ = ~new_n26553_ & ~new_n26589_;
  assign new_n26591_ = ~pi0778 & ~new_n26590_;
  assign new_n26592_ = ~pi0625 & new_n26589_;
  assign new_n26593_ = ~new_n26590_ & ~new_n26592_;
  assign new_n26594_ = pi1153 & ~new_n26593_;
  assign new_n26595_ = ~pi1153 & ~new_n26553_;
  assign new_n26596_ = ~new_n26592_ & new_n26595_;
  assign new_n26597_ = pi0778 & ~new_n26596_;
  assign new_n26598_ = ~new_n26594_ & new_n26597_;
  assign new_n26599_ = ~new_n26591_ & ~new_n26598_;
  assign new_n26600_ = ~new_n17844_ & ~new_n26599_;
  assign new_n26601_ = ~new_n17846_ & new_n26600_;
  assign new_n26602_ = ~new_n17848_ & new_n26601_;
  assign new_n26603_ = ~new_n17980_ & new_n26602_;
  assign new_n26604_ = ~new_n18011_ & new_n26603_;
  assign new_n26605_ = ~pi0647 & new_n26604_;
  assign new_n26606_ = pi0647 & new_n26553_;
  assign new_n26607_ = ~pi1157 & ~new_n26606_;
  assign new_n26608_ = ~new_n26605_ & new_n26607_;
  assign new_n26609_ = pi0630 & new_n26608_;
  assign new_n26610_ = pi0647 & ~new_n26604_;
  assign new_n26611_ = ~pi0647 & ~new_n26553_;
  assign new_n26612_ = ~new_n26610_ & ~new_n26611_;
  assign new_n26613_ = new_n17801_ & ~new_n26612_;
  assign new_n26614_ = ~new_n26609_ & ~new_n26613_;
  assign new_n26615_ = ~new_n26588_ & new_n26614_;
  assign new_n26616_ = pi0787 & ~new_n26615_;
  assign new_n26617_ = pi0626 & ~new_n26581_;
  assign new_n26618_ = ~pi0626 & ~new_n26553_;
  assign new_n26619_ = new_n17731_ & ~new_n26618_;
  assign new_n26620_ = ~new_n26617_ & new_n26619_;
  assign new_n26621_ = new_n17856_ & new_n26602_;
  assign new_n26622_ = ~pi0626 & ~new_n26581_;
  assign new_n26623_ = pi0626 & ~new_n26553_;
  assign new_n26624_ = new_n17732_ & ~new_n26623_;
  assign new_n26625_ = ~new_n26622_ & new_n26624_;
  assign new_n26626_ = ~new_n26621_ & ~new_n26625_;
  assign new_n26627_ = ~new_n26620_ & new_n26626_;
  assign new_n26628_ = pi0788 & ~new_n26627_;
  assign new_n26629_ = ~new_n16639_ & ~new_n26590_;
  assign new_n26630_ = pi0625 & new_n26629_;
  assign new_n26631_ = new_n26555_ & ~new_n26629_;
  assign new_n26632_ = ~new_n26630_ & ~new_n26631_;
  assign new_n26633_ = new_n26595_ & ~new_n26632_;
  assign new_n26634_ = ~pi0608 & ~new_n26594_;
  assign new_n26635_ = ~new_n26633_ & new_n26634_;
  assign new_n26636_ = pi1153 & new_n26555_;
  assign new_n26637_ = ~new_n26630_ & new_n26636_;
  assign new_n26638_ = pi0608 & ~new_n26596_;
  assign new_n26639_ = ~new_n26637_ & new_n26638_;
  assign new_n26640_ = ~new_n26635_ & ~new_n26639_;
  assign new_n26641_ = pi0778 & ~new_n26640_;
  assign new_n26642_ = ~pi0778 & ~new_n26631_;
  assign new_n26643_ = ~new_n26641_ & ~new_n26642_;
  assign new_n26644_ = ~pi0609 & ~new_n26643_;
  assign new_n26645_ = pi0609 & ~new_n26599_;
  assign new_n26646_ = ~pi1155 & ~new_n26645_;
  assign new_n26647_ = ~new_n26644_ & new_n26646_;
  assign new_n26648_ = ~pi0660 & ~new_n26560_;
  assign new_n26649_ = ~new_n26647_ & new_n26648_;
  assign new_n26650_ = pi0609 & ~new_n26643_;
  assign new_n26651_ = ~pi0609 & ~new_n26599_;
  assign new_n26652_ = pi1155 & ~new_n26651_;
  assign new_n26653_ = ~new_n26650_ & new_n26652_;
  assign new_n26654_ = pi0660 & ~new_n26562_;
  assign new_n26655_ = ~new_n26653_ & new_n26654_;
  assign new_n26656_ = ~new_n26649_ & ~new_n26655_;
  assign new_n26657_ = pi0785 & ~new_n26656_;
  assign new_n26658_ = ~pi0785 & ~new_n26643_;
  assign new_n26659_ = ~new_n26657_ & ~new_n26658_;
  assign new_n26660_ = ~pi0618 & ~new_n26659_;
  assign new_n26661_ = pi0618 & new_n26600_;
  assign new_n26662_ = ~pi1154 & ~new_n26661_;
  assign new_n26663_ = ~new_n26660_ & new_n26662_;
  assign new_n26664_ = ~pi0627 & ~new_n26568_;
  assign new_n26665_ = ~new_n26663_ & new_n26664_;
  assign new_n26666_ = pi0618 & ~new_n26659_;
  assign new_n26667_ = ~pi0618 & new_n26600_;
  assign new_n26668_ = pi1154 & ~new_n26667_;
  assign new_n26669_ = ~new_n26666_ & new_n26668_;
  assign new_n26670_ = pi0627 & ~new_n26570_;
  assign new_n26671_ = ~new_n26669_ & new_n26670_;
  assign new_n26672_ = ~new_n26665_ & ~new_n26671_;
  assign new_n26673_ = pi0781 & ~new_n26672_;
  assign new_n26674_ = ~pi0781 & ~new_n26659_;
  assign new_n26675_ = ~new_n26673_ & ~new_n26674_;
  assign new_n26676_ = pi0619 & ~new_n26675_;
  assign new_n26677_ = ~pi0619 & new_n26601_;
  assign new_n26678_ = pi1159 & ~new_n26677_;
  assign new_n26679_ = ~new_n26676_ & new_n26678_;
  assign new_n26680_ = pi0648 & ~new_n26578_;
  assign new_n26681_ = ~new_n26679_ & new_n26680_;
  assign new_n26682_ = ~pi0619 & ~new_n26675_;
  assign new_n26683_ = pi0619 & new_n26601_;
  assign new_n26684_ = ~pi1159 & ~new_n26683_;
  assign new_n26685_ = ~new_n26682_ & new_n26684_;
  assign new_n26686_ = ~pi0648 & ~new_n26576_;
  assign new_n26687_ = ~new_n26685_ & new_n26686_;
  assign new_n26688_ = pi0789 & ~new_n26687_;
  assign new_n26689_ = ~new_n26681_ & new_n26688_;
  assign new_n26690_ = ~pi0789 & new_n26675_;
  assign new_n26691_ = new_n17969_ & ~new_n26690_;
  assign new_n26692_ = ~new_n26689_ & new_n26691_;
  assign new_n26693_ = ~new_n26628_ & ~new_n26692_;
  assign new_n26694_ = ~new_n20364_ & ~new_n26693_;
  assign new_n26695_ = new_n18008_ & ~new_n26584_;
  assign new_n26696_ = new_n20851_ & new_n26603_;
  assign new_n26697_ = ~new_n26695_ & ~new_n26696_;
  assign new_n26698_ = ~pi0629 & ~new_n26697_;
  assign new_n26699_ = new_n20855_ & new_n26603_;
  assign new_n26700_ = new_n18007_ & ~new_n26584_;
  assign new_n26701_ = ~new_n26699_ & ~new_n26700_;
  assign new_n26702_ = pi0629 & ~new_n26701_;
  assign new_n26703_ = ~new_n26698_ & ~new_n26702_;
  assign new_n26704_ = pi0792 & ~new_n26703_;
  assign new_n26705_ = ~new_n20360_ & ~new_n26704_;
  assign new_n26706_ = ~new_n26694_ & new_n26705_;
  assign new_n26707_ = ~new_n26616_ & ~new_n26706_;
  assign new_n26708_ = pi0644 & new_n26707_;
  assign new_n26709_ = ~pi0787 & ~new_n26604_;
  assign new_n26710_ = pi1157 & ~new_n26612_;
  assign new_n26711_ = ~new_n26608_ & ~new_n26710_;
  assign new_n26712_ = pi0787 & ~new_n26711_;
  assign new_n26713_ = ~new_n26709_ & ~new_n26712_;
  assign new_n26714_ = ~pi0644 & new_n26713_;
  assign new_n26715_ = pi0715 & ~new_n26714_;
  assign new_n26716_ = ~new_n26708_ & new_n26715_;
  assign new_n26717_ = ~new_n17804_ & ~new_n26587_;
  assign new_n26718_ = new_n17804_ & new_n26553_;
  assign new_n26719_ = ~new_n26717_ & ~new_n26718_;
  assign new_n26720_ = pi0644 & ~new_n26719_;
  assign new_n26721_ = ~pi0644 & new_n26553_;
  assign new_n26722_ = ~pi0715 & ~new_n26721_;
  assign new_n26723_ = ~new_n26720_ & new_n26722_;
  assign new_n26724_ = pi1160 & ~new_n26723_;
  assign new_n26725_ = ~new_n26716_ & new_n26724_;
  assign new_n26726_ = ~pi0644 & new_n26707_;
  assign new_n26727_ = pi0644 & new_n26713_;
  assign new_n26728_ = ~pi0715 & ~new_n26727_;
  assign new_n26729_ = ~new_n26726_ & new_n26728_;
  assign new_n26730_ = ~pi0644 & ~new_n26719_;
  assign new_n26731_ = pi0644 & new_n26553_;
  assign new_n26732_ = pi0715 & ~new_n26731_;
  assign new_n26733_ = ~new_n26730_ & new_n26732_;
  assign new_n26734_ = ~pi1160 & ~new_n26733_;
  assign new_n26735_ = ~new_n26729_ & new_n26734_;
  assign new_n26736_ = ~new_n26725_ & ~new_n26735_;
  assign new_n26737_ = pi0790 & ~new_n26736_;
  assign new_n26738_ = ~pi0790 & new_n26707_;
  assign new_n26739_ = pi0832 & ~new_n26738_;
  assign new_n26740_ = ~new_n26737_ & new_n26739_;
  assign new_n26741_ = ~pi0181 & ~new_n17558_;
  assign new_n26742_ = new_n17691_ & ~new_n26741_;
  assign new_n26743_ = ~pi0709 & new_n3272_;
  assign new_n26744_ = new_n26741_ & ~new_n26743_;
  assign new_n26745_ = pi0181 & ~new_n18128_;
  assign new_n26746_ = ~pi0038 & ~new_n26745_;
  assign new_n26747_ = new_n3272_ & ~new_n26746_;
  assign new_n26748_ = ~pi0181 & new_n18124_;
  assign new_n26749_ = ~new_n26747_ & ~new_n26748_;
  assign new_n26750_ = ~pi0181 & ~new_n17431_;
  assign new_n26751_ = new_n17544_ & ~new_n26750_;
  assign new_n26752_ = ~pi0709 & ~new_n26751_;
  assign new_n26753_ = ~new_n26749_ & new_n26752_;
  assign new_n26754_ = ~new_n26744_ & ~new_n26753_;
  assign new_n26755_ = ~pi0778 & new_n26754_;
  assign new_n26756_ = pi0625 & ~new_n26754_;
  assign new_n26757_ = ~pi0625 & new_n26741_;
  assign new_n26758_ = pi1153 & ~new_n26757_;
  assign new_n26759_ = ~new_n26756_ & new_n26758_;
  assign new_n26760_ = ~pi0625 & ~new_n26754_;
  assign new_n26761_ = pi0625 & new_n26741_;
  assign new_n26762_ = ~pi1153 & ~new_n26761_;
  assign new_n26763_ = ~new_n26760_ & new_n26762_;
  assign new_n26764_ = ~new_n26759_ & ~new_n26763_;
  assign new_n26765_ = pi0778 & ~new_n26764_;
  assign new_n26766_ = ~new_n26755_ & ~new_n26765_;
  assign new_n26767_ = ~new_n17618_ & ~new_n26766_;
  assign new_n26768_ = new_n17618_ & ~new_n26741_;
  assign new_n26769_ = ~new_n26767_ & ~new_n26768_;
  assign new_n26770_ = ~new_n17655_ & new_n26769_;
  assign new_n26771_ = new_n17655_ & new_n26741_;
  assign new_n26772_ = ~new_n26770_ & ~new_n26771_;
  assign new_n26773_ = ~new_n17691_ & new_n26772_;
  assign new_n26774_ = ~new_n26742_ & ~new_n26773_;
  assign new_n26775_ = ~new_n17734_ & new_n26774_;
  assign new_n26776_ = new_n17734_ & new_n26741_;
  assign new_n26777_ = ~new_n26775_ & ~new_n26776_;
  assign new_n26778_ = ~pi0792 & new_n26777_;
  assign new_n26779_ = pi0628 & ~new_n26777_;
  assign new_n26780_ = ~pi0628 & new_n26741_;
  assign new_n26781_ = pi1156 & ~new_n26780_;
  assign new_n26782_ = ~new_n26779_ & new_n26781_;
  assign new_n26783_ = ~pi0628 & ~new_n26777_;
  assign new_n26784_ = pi0628 & new_n26741_;
  assign new_n26785_ = ~pi1156 & ~new_n26784_;
  assign new_n26786_ = ~new_n26783_ & new_n26785_;
  assign new_n26787_ = ~new_n26782_ & ~new_n26786_;
  assign new_n26788_ = pi0792 & ~new_n26787_;
  assign new_n26789_ = ~new_n26778_ & ~new_n26788_;
  assign new_n26790_ = ~pi0647 & ~new_n26789_;
  assign new_n26791_ = pi0647 & ~new_n26741_;
  assign new_n26792_ = ~new_n26790_ & ~new_n26791_;
  assign new_n26793_ = ~pi1157 & new_n26792_;
  assign new_n26794_ = pi0647 & ~new_n26789_;
  assign new_n26795_ = ~pi0647 & ~new_n26741_;
  assign new_n26796_ = ~new_n26794_ & ~new_n26795_;
  assign new_n26797_ = pi1157 & new_n26796_;
  assign new_n26798_ = ~new_n26793_ & ~new_n26797_;
  assign new_n26799_ = pi0787 & ~new_n26798_;
  assign new_n26800_ = ~pi0787 & new_n26789_;
  assign new_n26801_ = ~new_n26799_ & ~new_n26800_;
  assign new_n26802_ = ~pi0644 & ~new_n26801_;
  assign new_n26803_ = pi0715 & ~new_n26802_;
  assign new_n26804_ = pi0181 & ~new_n3272_;
  assign new_n26805_ = pi0754 & new_n17347_;
  assign new_n26806_ = pi0181 & new_n17424_;
  assign new_n26807_ = ~new_n26805_ & ~new_n26806_;
  assign new_n26808_ = pi0039 & ~new_n26807_;
  assign new_n26809_ = ~pi0181 & ~pi0754;
  assign new_n26810_ = new_n17393_ & new_n26809_;
  assign new_n26811_ = pi0181 & pi0754;
  assign new_n26812_ = pi0181 & ~new_n17215_;
  assign new_n26813_ = ~new_n21814_ & ~new_n26812_;
  assign new_n26814_ = ~pi0039 & ~new_n26813_;
  assign new_n26815_ = ~new_n26811_ & ~new_n26814_;
  assign new_n26816_ = ~new_n26810_ & new_n26815_;
  assign new_n26817_ = ~new_n26808_ & new_n26816_;
  assign new_n26818_ = ~pi0038 & ~new_n26817_;
  assign new_n26819_ = ~pi0754 & new_n17433_;
  assign new_n26820_ = pi0038 & ~new_n26750_;
  assign new_n26821_ = ~new_n26819_ & new_n26820_;
  assign new_n26822_ = ~new_n26818_ & ~new_n26821_;
  assign new_n26823_ = new_n3272_ & ~new_n26822_;
  assign new_n26824_ = ~new_n26804_ & ~new_n26823_;
  assign new_n26825_ = ~new_n17590_ & ~new_n26824_;
  assign new_n26826_ = new_n17590_ & ~new_n26741_;
  assign new_n26827_ = ~new_n26825_ & ~new_n26826_;
  assign new_n26828_ = ~pi0785 & ~new_n26827_;
  assign new_n26829_ = ~new_n17591_ & ~new_n26741_;
  assign new_n26830_ = pi0609 & new_n26825_;
  assign new_n26831_ = ~new_n26829_ & ~new_n26830_;
  assign new_n26832_ = pi1155 & ~new_n26831_;
  assign new_n26833_ = ~new_n17603_ & ~new_n26741_;
  assign new_n26834_ = ~pi0609 & new_n26825_;
  assign new_n26835_ = ~new_n26833_ & ~new_n26834_;
  assign new_n26836_ = ~pi1155 & ~new_n26835_;
  assign new_n26837_ = ~new_n26832_ & ~new_n26836_;
  assign new_n26838_ = pi0785 & ~new_n26837_;
  assign new_n26839_ = ~new_n26828_ & ~new_n26838_;
  assign new_n26840_ = ~pi0781 & ~new_n26839_;
  assign new_n26841_ = pi0618 & new_n26839_;
  assign new_n26842_ = ~pi0618 & new_n26741_;
  assign new_n26843_ = pi1154 & ~new_n26842_;
  assign new_n26844_ = ~new_n26841_ & new_n26843_;
  assign new_n26845_ = ~pi0618 & new_n26839_;
  assign new_n26846_ = pi0618 & new_n26741_;
  assign new_n26847_ = ~pi1154 & ~new_n26846_;
  assign new_n26848_ = ~new_n26845_ & new_n26847_;
  assign new_n26849_ = ~new_n26844_ & ~new_n26848_;
  assign new_n26850_ = pi0781 & ~new_n26849_;
  assign new_n26851_ = ~new_n26840_ & ~new_n26850_;
  assign new_n26852_ = ~pi0789 & ~new_n26851_;
  assign new_n26853_ = pi0619 & new_n26851_;
  assign new_n26854_ = ~pi0619 & new_n26741_;
  assign new_n26855_ = pi1159 & ~new_n26854_;
  assign new_n26856_ = ~new_n26853_ & new_n26855_;
  assign new_n26857_ = ~pi0619 & new_n26851_;
  assign new_n26858_ = pi0619 & new_n26741_;
  assign new_n26859_ = ~pi1159 & ~new_n26858_;
  assign new_n26860_ = ~new_n26857_ & new_n26859_;
  assign new_n26861_ = ~new_n26856_ & ~new_n26860_;
  assign new_n26862_ = pi0789 & ~new_n26861_;
  assign new_n26863_ = ~new_n26852_ & ~new_n26862_;
  assign new_n26864_ = ~new_n17968_ & new_n26863_;
  assign new_n26865_ = new_n17968_ & new_n26741_;
  assign new_n26866_ = ~new_n26864_ & ~new_n26865_;
  assign new_n26867_ = ~new_n17762_ & ~new_n26866_;
  assign new_n26868_ = new_n17762_ & new_n26741_;
  assign new_n26869_ = ~new_n26867_ & ~new_n26868_;
  assign new_n26870_ = ~new_n17804_ & ~new_n26869_;
  assign new_n26871_ = new_n17804_ & new_n26741_;
  assign new_n26872_ = ~new_n26870_ & ~new_n26871_;
  assign new_n26873_ = pi0644 & ~new_n26872_;
  assign new_n26874_ = ~pi0644 & new_n26741_;
  assign new_n26875_ = ~pi0715 & ~new_n26874_;
  assign new_n26876_ = ~new_n26873_ & new_n26875_;
  assign new_n26877_ = pi1160 & ~new_n26876_;
  assign new_n26878_ = ~new_n26803_ & new_n26877_;
  assign new_n26879_ = pi0644 & ~new_n26801_;
  assign new_n26880_ = ~pi0715 & ~new_n26879_;
  assign new_n26881_ = ~pi0644 & ~new_n26872_;
  assign new_n26882_ = pi0644 & new_n26741_;
  assign new_n26883_ = pi0715 & ~new_n26882_;
  assign new_n26884_ = ~new_n26881_ & new_n26883_;
  assign new_n26885_ = ~pi1160 & ~new_n26884_;
  assign new_n26886_ = ~new_n26880_ & new_n26885_;
  assign new_n26887_ = ~new_n26878_ & ~new_n26886_;
  assign new_n26888_ = pi0790 & ~new_n26887_;
  assign new_n26889_ = pi0644 & new_n26877_;
  assign new_n26890_ = ~pi0644 & new_n26885_;
  assign new_n26891_ = pi0790 & ~new_n26890_;
  assign new_n26892_ = ~new_n26889_ & new_n26891_;
  assign new_n26893_ = ~new_n20567_ & new_n26866_;
  assign new_n26894_ = ~pi0629 & new_n26782_;
  assign new_n26895_ = pi0629 & new_n26786_;
  assign new_n26896_ = ~new_n26894_ & ~new_n26895_;
  assign new_n26897_ = ~new_n26893_ & new_n26896_;
  assign new_n26898_ = pi0792 & ~new_n26897_;
  assign new_n26899_ = pi0709 & new_n26822_;
  assign new_n26900_ = ~pi0181 & new_n16810_;
  assign new_n26901_ = pi0181 & new_n16928_;
  assign new_n26902_ = pi0754 & ~new_n26901_;
  assign new_n26903_ = ~new_n26900_ & new_n26902_;
  assign new_n26904_ = pi0181 & new_n17007_;
  assign new_n26905_ = ~pi0181 & ~new_n17074_;
  assign new_n26906_ = ~pi0754 & ~new_n26905_;
  assign new_n26907_ = ~new_n26904_ & new_n26906_;
  assign new_n26908_ = pi0039 & ~new_n26907_;
  assign new_n26909_ = ~new_n26903_ & new_n26908_;
  assign new_n26910_ = ~pi0181 & ~new_n17217_;
  assign new_n26911_ = pi0181 & ~new_n17178_;
  assign new_n26912_ = pi0754 & ~new_n26911_;
  assign new_n26913_ = ~new_n26910_ & new_n26912_;
  assign new_n26914_ = ~pi0181 & new_n17227_;
  assign new_n26915_ = pi0181 & new_n17234_;
  assign new_n26916_ = ~pi0754 & ~new_n26915_;
  assign new_n26917_ = ~new_n26914_ & new_n26916_;
  assign new_n26918_ = ~new_n26913_ & ~new_n26917_;
  assign new_n26919_ = ~pi0039 & ~new_n26918_;
  assign new_n26920_ = ~pi0038 & ~new_n26919_;
  assign new_n26921_ = ~new_n26909_ & new_n26920_;
  assign new_n26922_ = ~pi0754 & ~new_n17035_;
  assign new_n26923_ = new_n19383_ & ~new_n26922_;
  assign new_n26924_ = ~pi0181 & ~new_n26923_;
  assign new_n26925_ = ~new_n16916_ & ~new_n26554_;
  assign new_n26926_ = pi0181 & ~new_n26925_;
  assign new_n26927_ = new_n6257_ & new_n26926_;
  assign new_n26928_ = pi0038 & ~new_n26927_;
  assign new_n26929_ = ~new_n26924_ & new_n26928_;
  assign new_n26930_ = ~pi0709 & ~new_n26929_;
  assign new_n26931_ = ~new_n26921_ & new_n26930_;
  assign new_n26932_ = new_n3272_ & ~new_n26931_;
  assign new_n26933_ = ~new_n26899_ & new_n26932_;
  assign new_n26934_ = ~new_n26804_ & ~new_n26933_;
  assign new_n26935_ = ~pi0625 & new_n26934_;
  assign new_n26936_ = pi0625 & new_n26824_;
  assign new_n26937_ = ~pi1153 & ~new_n26936_;
  assign new_n26938_ = ~new_n26935_ & new_n26937_;
  assign new_n26939_ = ~pi0608 & ~new_n26759_;
  assign new_n26940_ = ~new_n26938_ & new_n26939_;
  assign new_n26941_ = pi0625 & new_n26934_;
  assign new_n26942_ = ~pi0625 & new_n26824_;
  assign new_n26943_ = pi1153 & ~new_n26942_;
  assign new_n26944_ = ~new_n26941_ & new_n26943_;
  assign new_n26945_ = pi0608 & ~new_n26763_;
  assign new_n26946_ = ~new_n26944_ & new_n26945_;
  assign new_n26947_ = ~new_n26940_ & ~new_n26946_;
  assign new_n26948_ = pi0778 & ~new_n26947_;
  assign new_n26949_ = ~pi0778 & new_n26934_;
  assign new_n26950_ = ~new_n26948_ & ~new_n26949_;
  assign new_n26951_ = ~pi0609 & ~new_n26950_;
  assign new_n26952_ = pi0609 & new_n26766_;
  assign new_n26953_ = ~pi1155 & ~new_n26952_;
  assign new_n26954_ = ~new_n26951_ & new_n26953_;
  assign new_n26955_ = ~pi0660 & ~new_n26832_;
  assign new_n26956_ = ~new_n26954_ & new_n26955_;
  assign new_n26957_ = pi0609 & ~new_n26950_;
  assign new_n26958_ = ~pi0609 & new_n26766_;
  assign new_n26959_ = pi1155 & ~new_n26958_;
  assign new_n26960_ = ~new_n26957_ & new_n26959_;
  assign new_n26961_ = pi0660 & ~new_n26836_;
  assign new_n26962_ = ~new_n26960_ & new_n26961_;
  assign new_n26963_ = ~new_n26956_ & ~new_n26962_;
  assign new_n26964_ = pi0785 & ~new_n26963_;
  assign new_n26965_ = ~pi0785 & ~new_n26950_;
  assign new_n26966_ = ~new_n26964_ & ~new_n26965_;
  assign new_n26967_ = ~pi0618 & ~new_n26966_;
  assign new_n26968_ = pi0618 & new_n26769_;
  assign new_n26969_ = ~pi1154 & ~new_n26968_;
  assign new_n26970_ = ~new_n26967_ & new_n26969_;
  assign new_n26971_ = ~pi0627 & ~new_n26844_;
  assign new_n26972_ = ~new_n26970_ & new_n26971_;
  assign new_n26973_ = pi0618 & ~new_n26966_;
  assign new_n26974_ = ~pi0618 & new_n26769_;
  assign new_n26975_ = pi1154 & ~new_n26974_;
  assign new_n26976_ = ~new_n26973_ & new_n26975_;
  assign new_n26977_ = pi0627 & ~new_n26848_;
  assign new_n26978_ = ~new_n26976_ & new_n26977_;
  assign new_n26979_ = ~new_n26972_ & ~new_n26978_;
  assign new_n26980_ = pi0781 & ~new_n26979_;
  assign new_n26981_ = ~pi0781 & ~new_n26966_;
  assign new_n26982_ = ~new_n26980_ & ~new_n26981_;
  assign new_n26983_ = pi0619 & ~new_n26982_;
  assign new_n26984_ = ~pi0619 & ~new_n26772_;
  assign new_n26985_ = pi1159 & ~new_n26984_;
  assign new_n26986_ = ~new_n26983_ & new_n26985_;
  assign new_n26987_ = pi0648 & ~new_n26860_;
  assign new_n26988_ = ~new_n26986_ & new_n26987_;
  assign new_n26989_ = ~pi0619 & ~new_n26982_;
  assign new_n26990_ = pi0619 & ~new_n26772_;
  assign new_n26991_ = ~pi1159 & ~new_n26990_;
  assign new_n26992_ = ~new_n26989_ & new_n26991_;
  assign new_n26993_ = ~pi0648 & ~new_n26856_;
  assign new_n26994_ = ~new_n26992_ & new_n26993_;
  assign new_n26995_ = pi0789 & ~new_n26994_;
  assign new_n26996_ = ~new_n26988_ & new_n26995_;
  assign new_n26997_ = ~pi0789 & new_n26982_;
  assign new_n26998_ = new_n17969_ & ~new_n26997_;
  assign new_n26999_ = ~new_n26996_ & new_n26998_;
  assign new_n27000_ = pi0626 & ~new_n26863_;
  assign new_n27001_ = ~pi0626 & ~new_n26741_;
  assign new_n27002_ = new_n17731_ & ~new_n27001_;
  assign new_n27003_ = ~new_n27000_ & new_n27002_;
  assign new_n27004_ = new_n17856_ & new_n26774_;
  assign new_n27005_ = ~pi0626 & ~new_n26863_;
  assign new_n27006_ = pi0626 & ~new_n26741_;
  assign new_n27007_ = new_n17732_ & ~new_n27006_;
  assign new_n27008_ = ~new_n27005_ & new_n27007_;
  assign new_n27009_ = ~new_n27004_ & ~new_n27008_;
  assign new_n27010_ = ~new_n27003_ & new_n27009_;
  assign new_n27011_ = pi0788 & ~new_n27010_;
  assign new_n27012_ = ~new_n20364_ & ~new_n27011_;
  assign new_n27013_ = ~new_n26999_ & new_n27012_;
  assign new_n27014_ = ~new_n26898_ & ~new_n27013_;
  assign new_n27015_ = ~new_n20360_ & ~new_n27014_;
  assign new_n27016_ = ~new_n20556_ & new_n26869_;
  assign new_n27017_ = new_n17802_ & ~new_n26792_;
  assign new_n27018_ = new_n17801_ & ~new_n26796_;
  assign new_n27019_ = ~new_n27017_ & ~new_n27018_;
  assign new_n27020_ = ~new_n27016_ & new_n27019_;
  assign new_n27021_ = pi0787 & ~new_n27020_;
  assign new_n27022_ = ~new_n27015_ & ~new_n27021_;
  assign new_n27023_ = ~new_n26892_ & new_n27022_;
  assign new_n27024_ = ~new_n26888_ & ~new_n27023_;
  assign new_n27025_ = ~po1038 & ~new_n27024_;
  assign new_n27026_ = ~pi0181 & po1038;
  assign new_n27027_ = ~pi0832 & ~new_n27026_;
  assign new_n27028_ = ~new_n27025_ & new_n27027_;
  assign po0338 = ~new_n26740_ & ~new_n27028_;
  assign new_n27030_ = ~pi0182 & ~new_n2754_;
  assign new_n27031_ = ~pi0756 & new_n16913_;
  assign new_n27032_ = ~new_n27030_ & ~new_n27031_;
  assign new_n27033_ = ~new_n17858_ & ~new_n27032_;
  assign new_n27034_ = ~pi0785 & ~new_n27033_;
  assign new_n27035_ = new_n17603_ & new_n27031_;
  assign new_n27036_ = new_n27033_ & ~new_n27035_;
  assign new_n27037_ = pi1155 & ~new_n27036_;
  assign new_n27038_ = ~pi1155 & ~new_n27030_;
  assign new_n27039_ = ~new_n27035_ & new_n27038_;
  assign new_n27040_ = ~new_n27037_ & ~new_n27039_;
  assign new_n27041_ = pi0785 & ~new_n27040_;
  assign new_n27042_ = ~new_n27034_ & ~new_n27041_;
  assign new_n27043_ = ~pi0781 & ~new_n27042_;
  assign new_n27044_ = ~new_n17873_ & new_n27042_;
  assign new_n27045_ = pi1154 & ~new_n27044_;
  assign new_n27046_ = ~new_n17876_ & new_n27042_;
  assign new_n27047_ = ~pi1154 & ~new_n27046_;
  assign new_n27048_ = ~new_n27045_ & ~new_n27047_;
  assign new_n27049_ = pi0781 & ~new_n27048_;
  assign new_n27050_ = ~new_n27043_ & ~new_n27049_;
  assign new_n27051_ = ~pi0789 & ~new_n27050_;
  assign new_n27052_ = ~new_n23057_ & new_n27050_;
  assign new_n27053_ = pi1159 & ~new_n27052_;
  assign new_n27054_ = ~new_n23060_ & new_n27050_;
  assign new_n27055_ = ~pi1159 & ~new_n27054_;
  assign new_n27056_ = ~new_n27053_ & ~new_n27055_;
  assign new_n27057_ = pi0789 & ~new_n27056_;
  assign new_n27058_ = ~new_n27051_ & ~new_n27057_;
  assign new_n27059_ = ~new_n17968_ & new_n27058_;
  assign new_n27060_ = new_n17968_ & new_n27030_;
  assign new_n27061_ = ~new_n27059_ & ~new_n27060_;
  assign new_n27062_ = ~new_n17762_ & ~new_n27061_;
  assign new_n27063_ = new_n17762_ & new_n27030_;
  assign new_n27064_ = ~new_n27062_ & ~new_n27063_;
  assign new_n27065_ = ~new_n20556_ & new_n27064_;
  assign new_n27066_ = ~pi0734 & new_n16915_;
  assign new_n27067_ = ~new_n27030_ & ~new_n27066_;
  assign new_n27068_ = ~pi0778 & ~new_n27067_;
  assign new_n27069_ = ~pi0625 & new_n27066_;
  assign new_n27070_ = ~new_n27067_ & ~new_n27069_;
  assign new_n27071_ = pi1153 & ~new_n27070_;
  assign new_n27072_ = ~pi1153 & ~new_n27030_;
  assign new_n27073_ = ~new_n27069_ & new_n27072_;
  assign new_n27074_ = pi0778 & ~new_n27073_;
  assign new_n27075_ = ~new_n27071_ & new_n27074_;
  assign new_n27076_ = ~new_n27068_ & ~new_n27075_;
  assign new_n27077_ = ~new_n17844_ & ~new_n27076_;
  assign new_n27078_ = ~new_n17846_ & new_n27077_;
  assign new_n27079_ = ~new_n17848_ & new_n27078_;
  assign new_n27080_ = ~new_n17980_ & new_n27079_;
  assign new_n27081_ = ~new_n18011_ & new_n27080_;
  assign new_n27082_ = ~pi0647 & new_n27081_;
  assign new_n27083_ = pi0647 & new_n27030_;
  assign new_n27084_ = ~pi1157 & ~new_n27083_;
  assign new_n27085_ = ~new_n27082_ & new_n27084_;
  assign new_n27086_ = pi0630 & new_n27085_;
  assign new_n27087_ = pi0647 & ~new_n27081_;
  assign new_n27088_ = ~pi0647 & ~new_n27030_;
  assign new_n27089_ = ~new_n27087_ & ~new_n27088_;
  assign new_n27090_ = new_n17801_ & ~new_n27089_;
  assign new_n27091_ = ~new_n27086_ & ~new_n27090_;
  assign new_n27092_ = ~new_n27065_ & new_n27091_;
  assign new_n27093_ = pi0787 & ~new_n27092_;
  assign new_n27094_ = pi0626 & ~new_n27058_;
  assign new_n27095_ = ~pi0626 & ~new_n27030_;
  assign new_n27096_ = new_n17731_ & ~new_n27095_;
  assign new_n27097_ = ~new_n27094_ & new_n27096_;
  assign new_n27098_ = new_n17856_ & new_n27079_;
  assign new_n27099_ = ~pi0626 & ~new_n27058_;
  assign new_n27100_ = pi0626 & ~new_n27030_;
  assign new_n27101_ = new_n17732_ & ~new_n27100_;
  assign new_n27102_ = ~new_n27099_ & new_n27101_;
  assign new_n27103_ = ~new_n27098_ & ~new_n27102_;
  assign new_n27104_ = ~new_n27097_ & new_n27103_;
  assign new_n27105_ = pi0788 & ~new_n27104_;
  assign new_n27106_ = ~new_n16639_ & ~new_n27067_;
  assign new_n27107_ = pi0625 & new_n27106_;
  assign new_n27108_ = new_n27032_ & ~new_n27106_;
  assign new_n27109_ = ~new_n27107_ & ~new_n27108_;
  assign new_n27110_ = new_n27072_ & ~new_n27109_;
  assign new_n27111_ = ~pi0608 & ~new_n27071_;
  assign new_n27112_ = ~new_n27110_ & new_n27111_;
  assign new_n27113_ = pi1153 & new_n27032_;
  assign new_n27114_ = ~new_n27107_ & new_n27113_;
  assign new_n27115_ = pi0608 & ~new_n27073_;
  assign new_n27116_ = ~new_n27114_ & new_n27115_;
  assign new_n27117_ = ~new_n27112_ & ~new_n27116_;
  assign new_n27118_ = pi0778 & ~new_n27117_;
  assign new_n27119_ = ~pi0778 & ~new_n27108_;
  assign new_n27120_ = ~new_n27118_ & ~new_n27119_;
  assign new_n27121_ = ~pi0609 & ~new_n27120_;
  assign new_n27122_ = pi0609 & ~new_n27076_;
  assign new_n27123_ = ~pi1155 & ~new_n27122_;
  assign new_n27124_ = ~new_n27121_ & new_n27123_;
  assign new_n27125_ = ~pi0660 & ~new_n27037_;
  assign new_n27126_ = ~new_n27124_ & new_n27125_;
  assign new_n27127_ = pi0609 & ~new_n27120_;
  assign new_n27128_ = ~pi0609 & ~new_n27076_;
  assign new_n27129_ = pi1155 & ~new_n27128_;
  assign new_n27130_ = ~new_n27127_ & new_n27129_;
  assign new_n27131_ = pi0660 & ~new_n27039_;
  assign new_n27132_ = ~new_n27130_ & new_n27131_;
  assign new_n27133_ = ~new_n27126_ & ~new_n27132_;
  assign new_n27134_ = pi0785 & ~new_n27133_;
  assign new_n27135_ = ~pi0785 & ~new_n27120_;
  assign new_n27136_ = ~new_n27134_ & ~new_n27135_;
  assign new_n27137_ = ~pi0618 & ~new_n27136_;
  assign new_n27138_ = pi0618 & new_n27077_;
  assign new_n27139_ = ~pi1154 & ~new_n27138_;
  assign new_n27140_ = ~new_n27137_ & new_n27139_;
  assign new_n27141_ = ~pi0627 & ~new_n27045_;
  assign new_n27142_ = ~new_n27140_ & new_n27141_;
  assign new_n27143_ = pi0618 & ~new_n27136_;
  assign new_n27144_ = ~pi0618 & new_n27077_;
  assign new_n27145_ = pi1154 & ~new_n27144_;
  assign new_n27146_ = ~new_n27143_ & new_n27145_;
  assign new_n27147_ = pi0627 & ~new_n27047_;
  assign new_n27148_ = ~new_n27146_ & new_n27147_;
  assign new_n27149_ = ~new_n27142_ & ~new_n27148_;
  assign new_n27150_ = pi0781 & ~new_n27149_;
  assign new_n27151_ = ~pi0781 & ~new_n27136_;
  assign new_n27152_ = ~new_n27150_ & ~new_n27151_;
  assign new_n27153_ = pi0619 & ~new_n27152_;
  assign new_n27154_ = ~pi0619 & new_n27078_;
  assign new_n27155_ = pi1159 & ~new_n27154_;
  assign new_n27156_ = ~new_n27153_ & new_n27155_;
  assign new_n27157_ = pi0648 & ~new_n27055_;
  assign new_n27158_ = ~new_n27156_ & new_n27157_;
  assign new_n27159_ = ~pi0619 & ~new_n27152_;
  assign new_n27160_ = pi0619 & new_n27078_;
  assign new_n27161_ = ~pi1159 & ~new_n27160_;
  assign new_n27162_ = ~new_n27159_ & new_n27161_;
  assign new_n27163_ = ~pi0648 & ~new_n27053_;
  assign new_n27164_ = ~new_n27162_ & new_n27163_;
  assign new_n27165_ = pi0789 & ~new_n27164_;
  assign new_n27166_ = ~new_n27158_ & new_n27165_;
  assign new_n27167_ = ~pi0789 & new_n27152_;
  assign new_n27168_ = new_n17969_ & ~new_n27167_;
  assign new_n27169_ = ~new_n27166_ & new_n27168_;
  assign new_n27170_ = ~new_n27105_ & ~new_n27169_;
  assign new_n27171_ = ~new_n20364_ & ~new_n27170_;
  assign new_n27172_ = new_n18008_ & ~new_n27061_;
  assign new_n27173_ = new_n20851_ & new_n27080_;
  assign new_n27174_ = ~new_n27172_ & ~new_n27173_;
  assign new_n27175_ = ~pi0629 & ~new_n27174_;
  assign new_n27176_ = new_n20855_ & new_n27080_;
  assign new_n27177_ = new_n18007_ & ~new_n27061_;
  assign new_n27178_ = ~new_n27176_ & ~new_n27177_;
  assign new_n27179_ = pi0629 & ~new_n27178_;
  assign new_n27180_ = ~new_n27175_ & ~new_n27179_;
  assign new_n27181_ = pi0792 & ~new_n27180_;
  assign new_n27182_ = ~new_n20360_ & ~new_n27181_;
  assign new_n27183_ = ~new_n27171_ & new_n27182_;
  assign new_n27184_ = ~new_n27093_ & ~new_n27183_;
  assign new_n27185_ = pi0644 & new_n27184_;
  assign new_n27186_ = ~pi0787 & ~new_n27081_;
  assign new_n27187_ = pi1157 & ~new_n27089_;
  assign new_n27188_ = ~new_n27085_ & ~new_n27187_;
  assign new_n27189_ = pi0787 & ~new_n27188_;
  assign new_n27190_ = ~new_n27186_ & ~new_n27189_;
  assign new_n27191_ = ~pi0644 & new_n27190_;
  assign new_n27192_ = pi0715 & ~new_n27191_;
  assign new_n27193_ = ~new_n27185_ & new_n27192_;
  assign new_n27194_ = ~new_n17804_ & ~new_n27064_;
  assign new_n27195_ = new_n17804_ & new_n27030_;
  assign new_n27196_ = ~new_n27194_ & ~new_n27195_;
  assign new_n27197_ = pi0644 & ~new_n27196_;
  assign new_n27198_ = ~pi0644 & new_n27030_;
  assign new_n27199_ = ~pi0715 & ~new_n27198_;
  assign new_n27200_ = ~new_n27197_ & new_n27199_;
  assign new_n27201_ = pi1160 & ~new_n27200_;
  assign new_n27202_ = ~new_n27193_ & new_n27201_;
  assign new_n27203_ = ~pi0644 & new_n27184_;
  assign new_n27204_ = pi0644 & new_n27190_;
  assign new_n27205_ = ~pi0715 & ~new_n27204_;
  assign new_n27206_ = ~new_n27203_ & new_n27205_;
  assign new_n27207_ = ~pi0644 & ~new_n27196_;
  assign new_n27208_ = pi0644 & new_n27030_;
  assign new_n27209_ = pi0715 & ~new_n27208_;
  assign new_n27210_ = ~new_n27207_ & new_n27209_;
  assign new_n27211_ = ~pi1160 & ~new_n27210_;
  assign new_n27212_ = ~new_n27206_ & new_n27211_;
  assign new_n27213_ = ~new_n27202_ & ~new_n27212_;
  assign new_n27214_ = pi0790 & ~new_n27213_;
  assign new_n27215_ = ~pi0790 & new_n27184_;
  assign new_n27216_ = pi0832 & ~new_n27215_;
  assign new_n27217_ = ~new_n27214_ & new_n27216_;
  assign new_n27218_ = ~pi0182 & ~new_n17558_;
  assign new_n27219_ = new_n17691_ & ~new_n27218_;
  assign new_n27220_ = ~pi0734 & new_n3272_;
  assign new_n27221_ = new_n27218_ & ~new_n27220_;
  assign new_n27222_ = pi0182 & ~new_n18128_;
  assign new_n27223_ = ~pi0038 & ~new_n27222_;
  assign new_n27224_ = new_n3272_ & ~new_n27223_;
  assign new_n27225_ = ~pi0182 & new_n18124_;
  assign new_n27226_ = ~new_n27224_ & ~new_n27225_;
  assign new_n27227_ = ~pi0182 & ~new_n17431_;
  assign new_n27228_ = new_n17544_ & ~new_n27227_;
  assign new_n27229_ = ~pi0734 & ~new_n27228_;
  assign new_n27230_ = ~new_n27226_ & new_n27229_;
  assign new_n27231_ = ~new_n27221_ & ~new_n27230_;
  assign new_n27232_ = ~pi0778 & new_n27231_;
  assign new_n27233_ = pi0625 & ~new_n27231_;
  assign new_n27234_ = ~pi0625 & new_n27218_;
  assign new_n27235_ = pi1153 & ~new_n27234_;
  assign new_n27236_ = ~new_n27233_ & new_n27235_;
  assign new_n27237_ = ~pi0625 & ~new_n27231_;
  assign new_n27238_ = pi0625 & new_n27218_;
  assign new_n27239_ = ~pi1153 & ~new_n27238_;
  assign new_n27240_ = ~new_n27237_ & new_n27239_;
  assign new_n27241_ = ~new_n27236_ & ~new_n27240_;
  assign new_n27242_ = pi0778 & ~new_n27241_;
  assign new_n27243_ = ~new_n27232_ & ~new_n27242_;
  assign new_n27244_ = ~new_n17618_ & ~new_n27243_;
  assign new_n27245_ = new_n17618_ & ~new_n27218_;
  assign new_n27246_ = ~new_n27244_ & ~new_n27245_;
  assign new_n27247_ = ~new_n17655_ & new_n27246_;
  assign new_n27248_ = new_n17655_ & new_n27218_;
  assign new_n27249_ = ~new_n27247_ & ~new_n27248_;
  assign new_n27250_ = ~new_n17691_ & new_n27249_;
  assign new_n27251_ = ~new_n27219_ & ~new_n27250_;
  assign new_n27252_ = ~new_n17734_ & new_n27251_;
  assign new_n27253_ = new_n17734_ & new_n27218_;
  assign new_n27254_ = ~new_n27252_ & ~new_n27253_;
  assign new_n27255_ = ~pi0792 & new_n27254_;
  assign new_n27256_ = pi0628 & ~new_n27254_;
  assign new_n27257_ = ~pi0628 & new_n27218_;
  assign new_n27258_ = pi1156 & ~new_n27257_;
  assign new_n27259_ = ~new_n27256_ & new_n27258_;
  assign new_n27260_ = ~pi0628 & ~new_n27254_;
  assign new_n27261_ = pi0628 & new_n27218_;
  assign new_n27262_ = ~pi1156 & ~new_n27261_;
  assign new_n27263_ = ~new_n27260_ & new_n27262_;
  assign new_n27264_ = ~new_n27259_ & ~new_n27263_;
  assign new_n27265_ = pi0792 & ~new_n27264_;
  assign new_n27266_ = ~new_n27255_ & ~new_n27265_;
  assign new_n27267_ = ~pi0647 & ~new_n27266_;
  assign new_n27268_ = pi0647 & ~new_n27218_;
  assign new_n27269_ = ~new_n27267_ & ~new_n27268_;
  assign new_n27270_ = ~pi1157 & new_n27269_;
  assign new_n27271_ = pi0647 & ~new_n27266_;
  assign new_n27272_ = ~pi0647 & ~new_n27218_;
  assign new_n27273_ = ~new_n27271_ & ~new_n27272_;
  assign new_n27274_ = pi1157 & new_n27273_;
  assign new_n27275_ = ~new_n27270_ & ~new_n27274_;
  assign new_n27276_ = pi0787 & ~new_n27275_;
  assign new_n27277_ = ~pi0787 & new_n27266_;
  assign new_n27278_ = ~new_n27276_ & ~new_n27277_;
  assign new_n27279_ = ~pi0644 & ~new_n27278_;
  assign new_n27280_ = pi0715 & ~new_n27279_;
  assign new_n27281_ = pi0182 & ~new_n3272_;
  assign new_n27282_ = ~pi0756 & new_n17433_;
  assign new_n27283_ = ~new_n27227_ & ~new_n27282_;
  assign new_n27284_ = pi0038 & ~new_n27283_;
  assign new_n27285_ = ~pi0182 & new_n17393_;
  assign new_n27286_ = pi0182 & ~new_n17426_;
  assign new_n27287_ = ~pi0756 & ~new_n27286_;
  assign new_n27288_ = ~new_n27285_ & new_n27287_;
  assign new_n27289_ = ~pi0182 & pi0756;
  assign new_n27290_ = ~new_n17349_ & new_n27289_;
  assign new_n27291_ = ~new_n27288_ & ~new_n27290_;
  assign new_n27292_ = ~pi0038 & ~new_n27291_;
  assign new_n27293_ = ~new_n27284_ & ~new_n27292_;
  assign new_n27294_ = new_n3272_ & new_n27293_;
  assign new_n27295_ = ~new_n27281_ & ~new_n27294_;
  assign new_n27296_ = ~new_n17590_ & ~new_n27295_;
  assign new_n27297_ = new_n17590_ & ~new_n27218_;
  assign new_n27298_ = ~new_n27296_ & ~new_n27297_;
  assign new_n27299_ = ~pi0785 & ~new_n27298_;
  assign new_n27300_ = ~new_n17591_ & ~new_n27218_;
  assign new_n27301_ = pi0609 & new_n27296_;
  assign new_n27302_ = ~new_n27300_ & ~new_n27301_;
  assign new_n27303_ = pi1155 & ~new_n27302_;
  assign new_n27304_ = ~new_n17603_ & ~new_n27218_;
  assign new_n27305_ = ~pi0609 & new_n27296_;
  assign new_n27306_ = ~new_n27304_ & ~new_n27305_;
  assign new_n27307_ = ~pi1155 & ~new_n27306_;
  assign new_n27308_ = ~new_n27303_ & ~new_n27307_;
  assign new_n27309_ = pi0785 & ~new_n27308_;
  assign new_n27310_ = ~new_n27299_ & ~new_n27309_;
  assign new_n27311_ = ~pi0781 & ~new_n27310_;
  assign new_n27312_ = pi0618 & new_n27310_;
  assign new_n27313_ = ~pi0618 & new_n27218_;
  assign new_n27314_ = pi1154 & ~new_n27313_;
  assign new_n27315_ = ~new_n27312_ & new_n27314_;
  assign new_n27316_ = ~pi0618 & new_n27310_;
  assign new_n27317_ = pi0618 & new_n27218_;
  assign new_n27318_ = ~pi1154 & ~new_n27317_;
  assign new_n27319_ = ~new_n27316_ & new_n27318_;
  assign new_n27320_ = ~new_n27315_ & ~new_n27319_;
  assign new_n27321_ = pi0781 & ~new_n27320_;
  assign new_n27322_ = ~new_n27311_ & ~new_n27321_;
  assign new_n27323_ = ~pi0789 & ~new_n27322_;
  assign new_n27324_ = pi0619 & new_n27322_;
  assign new_n27325_ = ~pi0619 & new_n27218_;
  assign new_n27326_ = pi1159 & ~new_n27325_;
  assign new_n27327_ = ~new_n27324_ & new_n27326_;
  assign new_n27328_ = ~pi0619 & new_n27322_;
  assign new_n27329_ = pi0619 & new_n27218_;
  assign new_n27330_ = ~pi1159 & ~new_n27329_;
  assign new_n27331_ = ~new_n27328_ & new_n27330_;
  assign new_n27332_ = ~new_n27327_ & ~new_n27331_;
  assign new_n27333_ = pi0789 & ~new_n27332_;
  assign new_n27334_ = ~new_n27323_ & ~new_n27333_;
  assign new_n27335_ = ~new_n17968_ & new_n27334_;
  assign new_n27336_ = new_n17968_ & new_n27218_;
  assign new_n27337_ = ~new_n27335_ & ~new_n27336_;
  assign new_n27338_ = ~new_n17762_ & ~new_n27337_;
  assign new_n27339_ = new_n17762_ & new_n27218_;
  assign new_n27340_ = ~new_n27338_ & ~new_n27339_;
  assign new_n27341_ = ~new_n17804_ & ~new_n27340_;
  assign new_n27342_ = new_n17804_ & new_n27218_;
  assign new_n27343_ = ~new_n27341_ & ~new_n27342_;
  assign new_n27344_ = pi0644 & ~new_n27343_;
  assign new_n27345_ = ~pi0644 & new_n27218_;
  assign new_n27346_ = ~pi0715 & ~new_n27345_;
  assign new_n27347_ = ~new_n27344_ & new_n27346_;
  assign new_n27348_ = pi1160 & ~new_n27347_;
  assign new_n27349_ = ~new_n27280_ & new_n27348_;
  assign new_n27350_ = pi0644 & ~new_n27278_;
  assign new_n27351_ = ~pi0715 & ~new_n27350_;
  assign new_n27352_ = ~pi0644 & ~new_n27343_;
  assign new_n27353_ = pi0644 & new_n27218_;
  assign new_n27354_ = pi0715 & ~new_n27353_;
  assign new_n27355_ = ~new_n27352_ & new_n27354_;
  assign new_n27356_ = ~pi1160 & ~new_n27355_;
  assign new_n27357_ = ~new_n27351_ & new_n27356_;
  assign new_n27358_ = ~new_n27349_ & ~new_n27357_;
  assign new_n27359_ = pi0790 & ~new_n27358_;
  assign new_n27360_ = pi0644 & new_n27348_;
  assign new_n27361_ = ~pi0644 & new_n27356_;
  assign new_n27362_ = pi0790 & ~new_n27361_;
  assign new_n27363_ = ~new_n27360_ & new_n27362_;
  assign new_n27364_ = ~new_n20567_ & new_n27337_;
  assign new_n27365_ = ~pi0629 & new_n27259_;
  assign new_n27366_ = pi0629 & new_n27263_;
  assign new_n27367_ = ~new_n27365_ & ~new_n27366_;
  assign new_n27368_ = ~new_n27364_ & new_n27367_;
  assign new_n27369_ = pi0792 & ~new_n27368_;
  assign new_n27370_ = pi0734 & ~new_n27293_;
  assign new_n27371_ = ~pi0182 & new_n16810_;
  assign new_n27372_ = pi0182 & new_n16928_;
  assign new_n27373_ = pi0756 & ~new_n27372_;
  assign new_n27374_ = ~new_n27371_ & new_n27373_;
  assign new_n27375_ = pi0182 & new_n17007_;
  assign new_n27376_ = ~pi0182 & ~new_n17074_;
  assign new_n27377_ = ~pi0756 & ~new_n27376_;
  assign new_n27378_ = ~new_n27375_ & new_n27377_;
  assign new_n27379_ = pi0039 & ~new_n27378_;
  assign new_n27380_ = ~new_n27374_ & new_n27379_;
  assign new_n27381_ = ~pi0182 & ~new_n17217_;
  assign new_n27382_ = pi0182 & ~new_n17178_;
  assign new_n27383_ = pi0756 & ~new_n27382_;
  assign new_n27384_ = ~new_n27381_ & new_n27383_;
  assign new_n27385_ = ~pi0182 & new_n17227_;
  assign new_n27386_ = pi0182 & new_n17234_;
  assign new_n27387_ = ~pi0756 & ~new_n27386_;
  assign new_n27388_ = ~new_n27385_ & new_n27387_;
  assign new_n27389_ = ~new_n27384_ & ~new_n27388_;
  assign new_n27390_ = ~pi0039 & ~new_n27389_;
  assign new_n27391_ = ~pi0038 & ~new_n27390_;
  assign new_n27392_ = ~new_n27380_ & new_n27391_;
  assign new_n27393_ = ~pi0756 & ~new_n17035_;
  assign new_n27394_ = new_n19383_ & ~new_n27393_;
  assign new_n27395_ = ~pi0182 & ~new_n27394_;
  assign new_n27396_ = ~new_n16916_ & ~new_n27031_;
  assign new_n27397_ = pi0182 & ~new_n27396_;
  assign new_n27398_ = new_n6257_ & new_n27397_;
  assign new_n27399_ = pi0038 & ~new_n27398_;
  assign new_n27400_ = ~new_n27395_ & new_n27399_;
  assign new_n27401_ = ~pi0734 & ~new_n27400_;
  assign new_n27402_ = ~new_n27392_ & new_n27401_;
  assign new_n27403_ = new_n3272_ & ~new_n27402_;
  assign new_n27404_ = ~new_n27370_ & new_n27403_;
  assign new_n27405_ = ~new_n27281_ & ~new_n27404_;
  assign new_n27406_ = ~pi0625 & new_n27405_;
  assign new_n27407_ = pi0625 & new_n27295_;
  assign new_n27408_ = ~pi1153 & ~new_n27407_;
  assign new_n27409_ = ~new_n27406_ & new_n27408_;
  assign new_n27410_ = ~pi0608 & ~new_n27236_;
  assign new_n27411_ = ~new_n27409_ & new_n27410_;
  assign new_n27412_ = pi0625 & new_n27405_;
  assign new_n27413_ = ~pi0625 & new_n27295_;
  assign new_n27414_ = pi1153 & ~new_n27413_;
  assign new_n27415_ = ~new_n27412_ & new_n27414_;
  assign new_n27416_ = pi0608 & ~new_n27240_;
  assign new_n27417_ = ~new_n27415_ & new_n27416_;
  assign new_n27418_ = ~new_n27411_ & ~new_n27417_;
  assign new_n27419_ = pi0778 & ~new_n27418_;
  assign new_n27420_ = ~pi0778 & new_n27405_;
  assign new_n27421_ = ~new_n27419_ & ~new_n27420_;
  assign new_n27422_ = ~pi0609 & ~new_n27421_;
  assign new_n27423_ = pi0609 & new_n27243_;
  assign new_n27424_ = ~pi1155 & ~new_n27423_;
  assign new_n27425_ = ~new_n27422_ & new_n27424_;
  assign new_n27426_ = ~pi0660 & ~new_n27303_;
  assign new_n27427_ = ~new_n27425_ & new_n27426_;
  assign new_n27428_ = pi0609 & ~new_n27421_;
  assign new_n27429_ = ~pi0609 & new_n27243_;
  assign new_n27430_ = pi1155 & ~new_n27429_;
  assign new_n27431_ = ~new_n27428_ & new_n27430_;
  assign new_n27432_ = pi0660 & ~new_n27307_;
  assign new_n27433_ = ~new_n27431_ & new_n27432_;
  assign new_n27434_ = ~new_n27427_ & ~new_n27433_;
  assign new_n27435_ = pi0785 & ~new_n27434_;
  assign new_n27436_ = ~pi0785 & ~new_n27421_;
  assign new_n27437_ = ~new_n27435_ & ~new_n27436_;
  assign new_n27438_ = ~pi0618 & ~new_n27437_;
  assign new_n27439_ = pi0618 & new_n27246_;
  assign new_n27440_ = ~pi1154 & ~new_n27439_;
  assign new_n27441_ = ~new_n27438_ & new_n27440_;
  assign new_n27442_ = ~pi0627 & ~new_n27315_;
  assign new_n27443_ = ~new_n27441_ & new_n27442_;
  assign new_n27444_ = pi0618 & ~new_n27437_;
  assign new_n27445_ = ~pi0618 & new_n27246_;
  assign new_n27446_ = pi1154 & ~new_n27445_;
  assign new_n27447_ = ~new_n27444_ & new_n27446_;
  assign new_n27448_ = pi0627 & ~new_n27319_;
  assign new_n27449_ = ~new_n27447_ & new_n27448_;
  assign new_n27450_ = ~new_n27443_ & ~new_n27449_;
  assign new_n27451_ = pi0781 & ~new_n27450_;
  assign new_n27452_ = ~pi0781 & ~new_n27437_;
  assign new_n27453_ = ~new_n27451_ & ~new_n27452_;
  assign new_n27454_ = pi0619 & ~new_n27453_;
  assign new_n27455_ = ~pi0619 & ~new_n27249_;
  assign new_n27456_ = pi1159 & ~new_n27455_;
  assign new_n27457_ = ~new_n27454_ & new_n27456_;
  assign new_n27458_ = pi0648 & ~new_n27331_;
  assign new_n27459_ = ~new_n27457_ & new_n27458_;
  assign new_n27460_ = ~pi0619 & ~new_n27453_;
  assign new_n27461_ = pi0619 & ~new_n27249_;
  assign new_n27462_ = ~pi1159 & ~new_n27461_;
  assign new_n27463_ = ~new_n27460_ & new_n27462_;
  assign new_n27464_ = ~pi0648 & ~new_n27327_;
  assign new_n27465_ = ~new_n27463_ & new_n27464_;
  assign new_n27466_ = pi0789 & ~new_n27465_;
  assign new_n27467_ = ~new_n27459_ & new_n27466_;
  assign new_n27468_ = ~pi0789 & new_n27453_;
  assign new_n27469_ = new_n17969_ & ~new_n27468_;
  assign new_n27470_ = ~new_n27467_ & new_n27469_;
  assign new_n27471_ = pi0626 & ~new_n27334_;
  assign new_n27472_ = ~pi0626 & ~new_n27218_;
  assign new_n27473_ = new_n17731_ & ~new_n27472_;
  assign new_n27474_ = ~new_n27471_ & new_n27473_;
  assign new_n27475_ = new_n17856_ & new_n27251_;
  assign new_n27476_ = ~pi0626 & ~new_n27334_;
  assign new_n27477_ = pi0626 & ~new_n27218_;
  assign new_n27478_ = new_n17732_ & ~new_n27477_;
  assign new_n27479_ = ~new_n27476_ & new_n27478_;
  assign new_n27480_ = ~new_n27475_ & ~new_n27479_;
  assign new_n27481_ = ~new_n27474_ & new_n27480_;
  assign new_n27482_ = pi0788 & ~new_n27481_;
  assign new_n27483_ = ~new_n20364_ & ~new_n27482_;
  assign new_n27484_ = ~new_n27470_ & new_n27483_;
  assign new_n27485_ = ~new_n27369_ & ~new_n27484_;
  assign new_n27486_ = ~new_n20360_ & ~new_n27485_;
  assign new_n27487_ = ~new_n20556_ & new_n27340_;
  assign new_n27488_ = new_n17802_ & ~new_n27269_;
  assign new_n27489_ = new_n17801_ & ~new_n27273_;
  assign new_n27490_ = ~new_n27488_ & ~new_n27489_;
  assign new_n27491_ = ~new_n27487_ & new_n27490_;
  assign new_n27492_ = pi0787 & ~new_n27491_;
  assign new_n27493_ = ~new_n27486_ & ~new_n27492_;
  assign new_n27494_ = ~new_n27363_ & new_n27493_;
  assign new_n27495_ = ~new_n27359_ & ~new_n27494_;
  assign new_n27496_ = ~po1038 & ~new_n27495_;
  assign new_n27497_ = ~pi0182 & po1038;
  assign new_n27498_ = ~pi0832 & ~new_n27497_;
  assign new_n27499_ = ~new_n27496_ & new_n27498_;
  assign po0339 = ~new_n27217_ & ~new_n27499_;
  assign new_n27501_ = ~pi0183 & ~new_n2754_;
  assign new_n27502_ = ~pi0755 & new_n16913_;
  assign new_n27503_ = ~new_n27501_ & ~new_n27502_;
  assign new_n27504_ = ~new_n17858_ & ~new_n27503_;
  assign new_n27505_ = ~pi0785 & ~new_n27504_;
  assign new_n27506_ = new_n17603_ & new_n27502_;
  assign new_n27507_ = new_n27504_ & ~new_n27506_;
  assign new_n27508_ = pi1155 & ~new_n27507_;
  assign new_n27509_ = ~pi1155 & ~new_n27501_;
  assign new_n27510_ = ~new_n27506_ & new_n27509_;
  assign new_n27511_ = ~new_n27508_ & ~new_n27510_;
  assign new_n27512_ = pi0785 & ~new_n27511_;
  assign new_n27513_ = ~new_n27505_ & ~new_n27512_;
  assign new_n27514_ = ~pi0781 & ~new_n27513_;
  assign new_n27515_ = ~new_n17873_ & new_n27513_;
  assign new_n27516_ = pi1154 & ~new_n27515_;
  assign new_n27517_ = ~new_n17876_ & new_n27513_;
  assign new_n27518_ = ~pi1154 & ~new_n27517_;
  assign new_n27519_ = ~new_n27516_ & ~new_n27518_;
  assign new_n27520_ = pi0781 & ~new_n27519_;
  assign new_n27521_ = ~new_n27514_ & ~new_n27520_;
  assign new_n27522_ = ~pi0789 & ~new_n27521_;
  assign new_n27523_ = ~new_n23057_ & new_n27521_;
  assign new_n27524_ = pi1159 & ~new_n27523_;
  assign new_n27525_ = ~new_n23060_ & new_n27521_;
  assign new_n27526_ = ~pi1159 & ~new_n27525_;
  assign new_n27527_ = ~new_n27524_ & ~new_n27526_;
  assign new_n27528_ = pi0789 & ~new_n27527_;
  assign new_n27529_ = ~new_n27522_ & ~new_n27528_;
  assign new_n27530_ = ~new_n17968_ & new_n27529_;
  assign new_n27531_ = new_n17968_ & new_n27501_;
  assign new_n27532_ = ~new_n27530_ & ~new_n27531_;
  assign new_n27533_ = ~new_n17762_ & ~new_n27532_;
  assign new_n27534_ = new_n17762_ & new_n27501_;
  assign new_n27535_ = ~new_n27533_ & ~new_n27534_;
  assign new_n27536_ = ~new_n20556_ & new_n27535_;
  assign new_n27537_ = ~pi0725 & new_n16915_;
  assign new_n27538_ = ~new_n27501_ & ~new_n27537_;
  assign new_n27539_ = ~pi0778 & ~new_n27538_;
  assign new_n27540_ = ~pi0625 & new_n27537_;
  assign new_n27541_ = ~new_n27538_ & ~new_n27540_;
  assign new_n27542_ = pi1153 & ~new_n27541_;
  assign new_n27543_ = ~pi1153 & ~new_n27501_;
  assign new_n27544_ = ~new_n27540_ & new_n27543_;
  assign new_n27545_ = pi0778 & ~new_n27544_;
  assign new_n27546_ = ~new_n27542_ & new_n27545_;
  assign new_n27547_ = ~new_n27539_ & ~new_n27546_;
  assign new_n27548_ = ~new_n17844_ & ~new_n27547_;
  assign new_n27549_ = ~new_n17846_ & new_n27548_;
  assign new_n27550_ = ~new_n17848_ & new_n27549_;
  assign new_n27551_ = ~new_n17980_ & new_n27550_;
  assign new_n27552_ = ~new_n18011_ & new_n27551_;
  assign new_n27553_ = ~pi0647 & new_n27552_;
  assign new_n27554_ = pi0647 & new_n27501_;
  assign new_n27555_ = ~pi1157 & ~new_n27554_;
  assign new_n27556_ = ~new_n27553_ & new_n27555_;
  assign new_n27557_ = pi0630 & new_n27556_;
  assign new_n27558_ = pi0647 & ~new_n27552_;
  assign new_n27559_ = ~pi0647 & ~new_n27501_;
  assign new_n27560_ = ~new_n27558_ & ~new_n27559_;
  assign new_n27561_ = new_n17801_ & ~new_n27560_;
  assign new_n27562_ = ~new_n27557_ & ~new_n27561_;
  assign new_n27563_ = ~new_n27536_ & new_n27562_;
  assign new_n27564_ = pi0787 & ~new_n27563_;
  assign new_n27565_ = pi0626 & ~new_n27529_;
  assign new_n27566_ = ~pi0626 & ~new_n27501_;
  assign new_n27567_ = new_n17731_ & ~new_n27566_;
  assign new_n27568_ = ~new_n27565_ & new_n27567_;
  assign new_n27569_ = new_n17856_ & new_n27550_;
  assign new_n27570_ = ~pi0626 & ~new_n27529_;
  assign new_n27571_ = pi0626 & ~new_n27501_;
  assign new_n27572_ = new_n17732_ & ~new_n27571_;
  assign new_n27573_ = ~new_n27570_ & new_n27572_;
  assign new_n27574_ = ~new_n27569_ & ~new_n27573_;
  assign new_n27575_ = ~new_n27568_ & new_n27574_;
  assign new_n27576_ = pi0788 & ~new_n27575_;
  assign new_n27577_ = ~new_n16639_ & ~new_n27538_;
  assign new_n27578_ = pi0625 & new_n27577_;
  assign new_n27579_ = new_n27503_ & ~new_n27577_;
  assign new_n27580_ = ~new_n27578_ & ~new_n27579_;
  assign new_n27581_ = new_n27543_ & ~new_n27580_;
  assign new_n27582_ = ~pi0608 & ~new_n27542_;
  assign new_n27583_ = ~new_n27581_ & new_n27582_;
  assign new_n27584_ = pi1153 & new_n27503_;
  assign new_n27585_ = ~new_n27578_ & new_n27584_;
  assign new_n27586_ = pi0608 & ~new_n27544_;
  assign new_n27587_ = ~new_n27585_ & new_n27586_;
  assign new_n27588_ = ~new_n27583_ & ~new_n27587_;
  assign new_n27589_ = pi0778 & ~new_n27588_;
  assign new_n27590_ = ~pi0778 & ~new_n27579_;
  assign new_n27591_ = ~new_n27589_ & ~new_n27590_;
  assign new_n27592_ = ~pi0609 & ~new_n27591_;
  assign new_n27593_ = pi0609 & ~new_n27547_;
  assign new_n27594_ = ~pi1155 & ~new_n27593_;
  assign new_n27595_ = ~new_n27592_ & new_n27594_;
  assign new_n27596_ = ~pi0660 & ~new_n27508_;
  assign new_n27597_ = ~new_n27595_ & new_n27596_;
  assign new_n27598_ = pi0609 & ~new_n27591_;
  assign new_n27599_ = ~pi0609 & ~new_n27547_;
  assign new_n27600_ = pi1155 & ~new_n27599_;
  assign new_n27601_ = ~new_n27598_ & new_n27600_;
  assign new_n27602_ = pi0660 & ~new_n27510_;
  assign new_n27603_ = ~new_n27601_ & new_n27602_;
  assign new_n27604_ = ~new_n27597_ & ~new_n27603_;
  assign new_n27605_ = pi0785 & ~new_n27604_;
  assign new_n27606_ = ~pi0785 & ~new_n27591_;
  assign new_n27607_ = ~new_n27605_ & ~new_n27606_;
  assign new_n27608_ = ~pi0618 & ~new_n27607_;
  assign new_n27609_ = pi0618 & new_n27548_;
  assign new_n27610_ = ~pi1154 & ~new_n27609_;
  assign new_n27611_ = ~new_n27608_ & new_n27610_;
  assign new_n27612_ = ~pi0627 & ~new_n27516_;
  assign new_n27613_ = ~new_n27611_ & new_n27612_;
  assign new_n27614_ = pi0618 & ~new_n27607_;
  assign new_n27615_ = ~pi0618 & new_n27548_;
  assign new_n27616_ = pi1154 & ~new_n27615_;
  assign new_n27617_ = ~new_n27614_ & new_n27616_;
  assign new_n27618_ = pi0627 & ~new_n27518_;
  assign new_n27619_ = ~new_n27617_ & new_n27618_;
  assign new_n27620_ = ~new_n27613_ & ~new_n27619_;
  assign new_n27621_ = pi0781 & ~new_n27620_;
  assign new_n27622_ = ~pi0781 & ~new_n27607_;
  assign new_n27623_ = ~new_n27621_ & ~new_n27622_;
  assign new_n27624_ = pi0619 & ~new_n27623_;
  assign new_n27625_ = ~pi0619 & new_n27549_;
  assign new_n27626_ = pi1159 & ~new_n27625_;
  assign new_n27627_ = ~new_n27624_ & new_n27626_;
  assign new_n27628_ = pi0648 & ~new_n27526_;
  assign new_n27629_ = ~new_n27627_ & new_n27628_;
  assign new_n27630_ = ~pi0619 & ~new_n27623_;
  assign new_n27631_ = pi0619 & new_n27549_;
  assign new_n27632_ = ~pi1159 & ~new_n27631_;
  assign new_n27633_ = ~new_n27630_ & new_n27632_;
  assign new_n27634_ = ~pi0648 & ~new_n27524_;
  assign new_n27635_ = ~new_n27633_ & new_n27634_;
  assign new_n27636_ = pi0789 & ~new_n27635_;
  assign new_n27637_ = ~new_n27629_ & new_n27636_;
  assign new_n27638_ = ~pi0789 & new_n27623_;
  assign new_n27639_ = new_n17969_ & ~new_n27638_;
  assign new_n27640_ = ~new_n27637_ & new_n27639_;
  assign new_n27641_ = ~new_n27576_ & ~new_n27640_;
  assign new_n27642_ = ~new_n20364_ & ~new_n27641_;
  assign new_n27643_ = new_n18008_ & ~new_n27532_;
  assign new_n27644_ = new_n20851_ & new_n27551_;
  assign new_n27645_ = ~new_n27643_ & ~new_n27644_;
  assign new_n27646_ = ~pi0629 & ~new_n27645_;
  assign new_n27647_ = new_n20855_ & new_n27551_;
  assign new_n27648_ = new_n18007_ & ~new_n27532_;
  assign new_n27649_ = ~new_n27647_ & ~new_n27648_;
  assign new_n27650_ = pi0629 & ~new_n27649_;
  assign new_n27651_ = ~new_n27646_ & ~new_n27650_;
  assign new_n27652_ = pi0792 & ~new_n27651_;
  assign new_n27653_ = ~new_n20360_ & ~new_n27652_;
  assign new_n27654_ = ~new_n27642_ & new_n27653_;
  assign new_n27655_ = ~new_n27564_ & ~new_n27654_;
  assign new_n27656_ = pi0644 & new_n27655_;
  assign new_n27657_ = ~pi0787 & ~new_n27552_;
  assign new_n27658_ = pi1157 & ~new_n27560_;
  assign new_n27659_ = ~new_n27556_ & ~new_n27658_;
  assign new_n27660_ = pi0787 & ~new_n27659_;
  assign new_n27661_ = ~new_n27657_ & ~new_n27660_;
  assign new_n27662_ = ~pi0644 & new_n27661_;
  assign new_n27663_ = pi0715 & ~new_n27662_;
  assign new_n27664_ = ~new_n27656_ & new_n27663_;
  assign new_n27665_ = ~new_n17804_ & ~new_n27535_;
  assign new_n27666_ = new_n17804_ & new_n27501_;
  assign new_n27667_ = ~new_n27665_ & ~new_n27666_;
  assign new_n27668_ = pi0644 & ~new_n27667_;
  assign new_n27669_ = ~pi0644 & new_n27501_;
  assign new_n27670_ = ~pi0715 & ~new_n27669_;
  assign new_n27671_ = ~new_n27668_ & new_n27670_;
  assign new_n27672_ = pi1160 & ~new_n27671_;
  assign new_n27673_ = ~new_n27664_ & new_n27672_;
  assign new_n27674_ = ~pi0644 & new_n27655_;
  assign new_n27675_ = pi0644 & new_n27661_;
  assign new_n27676_ = ~pi0715 & ~new_n27675_;
  assign new_n27677_ = ~new_n27674_ & new_n27676_;
  assign new_n27678_ = ~pi0644 & ~new_n27667_;
  assign new_n27679_ = pi0644 & new_n27501_;
  assign new_n27680_ = pi0715 & ~new_n27679_;
  assign new_n27681_ = ~new_n27678_ & new_n27680_;
  assign new_n27682_ = ~pi1160 & ~new_n27681_;
  assign new_n27683_ = ~new_n27677_ & new_n27682_;
  assign new_n27684_ = ~new_n27673_ & ~new_n27683_;
  assign new_n27685_ = pi0790 & ~new_n27684_;
  assign new_n27686_ = ~pi0790 & new_n27655_;
  assign new_n27687_ = pi0832 & ~new_n27686_;
  assign new_n27688_ = ~new_n27685_ & new_n27687_;
  assign new_n27689_ = ~pi0183 & ~new_n17558_;
  assign new_n27690_ = new_n17691_ & ~new_n27689_;
  assign new_n27691_ = ~pi0725 & new_n3272_;
  assign new_n27692_ = new_n27689_ & ~new_n27691_;
  assign new_n27693_ = pi0183 & ~new_n18128_;
  assign new_n27694_ = ~pi0038 & ~new_n27693_;
  assign new_n27695_ = new_n3272_ & ~new_n27694_;
  assign new_n27696_ = ~pi0183 & new_n18124_;
  assign new_n27697_ = ~new_n27695_ & ~new_n27696_;
  assign new_n27698_ = ~pi0183 & ~new_n17431_;
  assign new_n27699_ = new_n17544_ & ~new_n27698_;
  assign new_n27700_ = ~pi0725 & ~new_n27699_;
  assign new_n27701_ = ~new_n27697_ & new_n27700_;
  assign new_n27702_ = ~new_n27692_ & ~new_n27701_;
  assign new_n27703_ = ~pi0778 & new_n27702_;
  assign new_n27704_ = pi0625 & ~new_n27702_;
  assign new_n27705_ = ~pi0625 & new_n27689_;
  assign new_n27706_ = pi1153 & ~new_n27705_;
  assign new_n27707_ = ~new_n27704_ & new_n27706_;
  assign new_n27708_ = ~pi0625 & ~new_n27702_;
  assign new_n27709_ = pi0625 & new_n27689_;
  assign new_n27710_ = ~pi1153 & ~new_n27709_;
  assign new_n27711_ = ~new_n27708_ & new_n27710_;
  assign new_n27712_ = ~new_n27707_ & ~new_n27711_;
  assign new_n27713_ = pi0778 & ~new_n27712_;
  assign new_n27714_ = ~new_n27703_ & ~new_n27713_;
  assign new_n27715_ = ~new_n17618_ & ~new_n27714_;
  assign new_n27716_ = new_n17618_ & ~new_n27689_;
  assign new_n27717_ = ~new_n27715_ & ~new_n27716_;
  assign new_n27718_ = ~new_n17655_ & new_n27717_;
  assign new_n27719_ = new_n17655_ & new_n27689_;
  assign new_n27720_ = ~new_n27718_ & ~new_n27719_;
  assign new_n27721_ = ~new_n17691_ & new_n27720_;
  assign new_n27722_ = ~new_n27690_ & ~new_n27721_;
  assign new_n27723_ = ~new_n17734_ & new_n27722_;
  assign new_n27724_ = new_n17734_ & new_n27689_;
  assign new_n27725_ = ~new_n27723_ & ~new_n27724_;
  assign new_n27726_ = ~pi0792 & new_n27725_;
  assign new_n27727_ = pi0628 & ~new_n27725_;
  assign new_n27728_ = ~pi0628 & new_n27689_;
  assign new_n27729_ = pi1156 & ~new_n27728_;
  assign new_n27730_ = ~new_n27727_ & new_n27729_;
  assign new_n27731_ = ~pi0628 & ~new_n27725_;
  assign new_n27732_ = pi0628 & new_n27689_;
  assign new_n27733_ = ~pi1156 & ~new_n27732_;
  assign new_n27734_ = ~new_n27731_ & new_n27733_;
  assign new_n27735_ = ~new_n27730_ & ~new_n27734_;
  assign new_n27736_ = pi0792 & ~new_n27735_;
  assign new_n27737_ = ~new_n27726_ & ~new_n27736_;
  assign new_n27738_ = ~pi0647 & ~new_n27737_;
  assign new_n27739_ = pi0647 & ~new_n27689_;
  assign new_n27740_ = ~new_n27738_ & ~new_n27739_;
  assign new_n27741_ = ~pi1157 & new_n27740_;
  assign new_n27742_ = pi0647 & ~new_n27737_;
  assign new_n27743_ = ~pi0647 & ~new_n27689_;
  assign new_n27744_ = ~new_n27742_ & ~new_n27743_;
  assign new_n27745_ = pi1157 & new_n27744_;
  assign new_n27746_ = ~new_n27741_ & ~new_n27745_;
  assign new_n27747_ = pi0787 & ~new_n27746_;
  assign new_n27748_ = ~pi0787 & new_n27737_;
  assign new_n27749_ = ~new_n27747_ & ~new_n27748_;
  assign new_n27750_ = ~pi0644 & ~new_n27749_;
  assign new_n27751_ = pi0715 & ~new_n27750_;
  assign new_n27752_ = pi0183 & ~new_n3272_;
  assign new_n27753_ = ~pi0755 & new_n17433_;
  assign new_n27754_ = ~new_n27698_ & ~new_n27753_;
  assign new_n27755_ = pi0038 & ~new_n27754_;
  assign new_n27756_ = ~pi0183 & new_n17393_;
  assign new_n27757_ = pi0183 & ~new_n17426_;
  assign new_n27758_ = ~pi0755 & ~new_n27757_;
  assign new_n27759_ = ~new_n27756_ & new_n27758_;
  assign new_n27760_ = ~pi0183 & pi0755;
  assign new_n27761_ = ~new_n17349_ & new_n27760_;
  assign new_n27762_ = ~new_n27759_ & ~new_n27761_;
  assign new_n27763_ = ~pi0038 & ~new_n27762_;
  assign new_n27764_ = ~new_n27755_ & ~new_n27763_;
  assign new_n27765_ = new_n3272_ & new_n27764_;
  assign new_n27766_ = ~new_n27752_ & ~new_n27765_;
  assign new_n27767_ = ~new_n17590_ & ~new_n27766_;
  assign new_n27768_ = new_n17590_ & ~new_n27689_;
  assign new_n27769_ = ~new_n27767_ & ~new_n27768_;
  assign new_n27770_ = ~pi0785 & ~new_n27769_;
  assign new_n27771_ = ~new_n17591_ & ~new_n27689_;
  assign new_n27772_ = pi0609 & new_n27767_;
  assign new_n27773_ = ~new_n27771_ & ~new_n27772_;
  assign new_n27774_ = pi1155 & ~new_n27773_;
  assign new_n27775_ = ~new_n17603_ & ~new_n27689_;
  assign new_n27776_ = ~pi0609 & new_n27767_;
  assign new_n27777_ = ~new_n27775_ & ~new_n27776_;
  assign new_n27778_ = ~pi1155 & ~new_n27777_;
  assign new_n27779_ = ~new_n27774_ & ~new_n27778_;
  assign new_n27780_ = pi0785 & ~new_n27779_;
  assign new_n27781_ = ~new_n27770_ & ~new_n27780_;
  assign new_n27782_ = ~pi0781 & ~new_n27781_;
  assign new_n27783_ = pi0618 & new_n27781_;
  assign new_n27784_ = ~pi0618 & new_n27689_;
  assign new_n27785_ = pi1154 & ~new_n27784_;
  assign new_n27786_ = ~new_n27783_ & new_n27785_;
  assign new_n27787_ = ~pi0618 & new_n27781_;
  assign new_n27788_ = pi0618 & new_n27689_;
  assign new_n27789_ = ~pi1154 & ~new_n27788_;
  assign new_n27790_ = ~new_n27787_ & new_n27789_;
  assign new_n27791_ = ~new_n27786_ & ~new_n27790_;
  assign new_n27792_ = pi0781 & ~new_n27791_;
  assign new_n27793_ = ~new_n27782_ & ~new_n27792_;
  assign new_n27794_ = ~pi0789 & ~new_n27793_;
  assign new_n27795_ = pi0619 & new_n27793_;
  assign new_n27796_ = ~pi0619 & new_n27689_;
  assign new_n27797_ = pi1159 & ~new_n27796_;
  assign new_n27798_ = ~new_n27795_ & new_n27797_;
  assign new_n27799_ = ~pi0619 & new_n27793_;
  assign new_n27800_ = pi0619 & new_n27689_;
  assign new_n27801_ = ~pi1159 & ~new_n27800_;
  assign new_n27802_ = ~new_n27799_ & new_n27801_;
  assign new_n27803_ = ~new_n27798_ & ~new_n27802_;
  assign new_n27804_ = pi0789 & ~new_n27803_;
  assign new_n27805_ = ~new_n27794_ & ~new_n27804_;
  assign new_n27806_ = ~new_n17968_ & new_n27805_;
  assign new_n27807_ = new_n17968_ & new_n27689_;
  assign new_n27808_ = ~new_n27806_ & ~new_n27807_;
  assign new_n27809_ = ~new_n17762_ & ~new_n27808_;
  assign new_n27810_ = new_n17762_ & new_n27689_;
  assign new_n27811_ = ~new_n27809_ & ~new_n27810_;
  assign new_n27812_ = ~new_n17804_ & ~new_n27811_;
  assign new_n27813_ = new_n17804_ & new_n27689_;
  assign new_n27814_ = ~new_n27812_ & ~new_n27813_;
  assign new_n27815_ = pi0644 & ~new_n27814_;
  assign new_n27816_ = ~pi0644 & new_n27689_;
  assign new_n27817_ = ~pi0715 & ~new_n27816_;
  assign new_n27818_ = ~new_n27815_ & new_n27817_;
  assign new_n27819_ = pi1160 & ~new_n27818_;
  assign new_n27820_ = ~new_n27751_ & new_n27819_;
  assign new_n27821_ = pi0644 & ~new_n27749_;
  assign new_n27822_ = ~pi0715 & ~new_n27821_;
  assign new_n27823_ = ~pi0644 & ~new_n27814_;
  assign new_n27824_ = pi0644 & new_n27689_;
  assign new_n27825_ = pi0715 & ~new_n27824_;
  assign new_n27826_ = ~new_n27823_ & new_n27825_;
  assign new_n27827_ = ~pi1160 & ~new_n27826_;
  assign new_n27828_ = ~new_n27822_ & new_n27827_;
  assign new_n27829_ = ~new_n27820_ & ~new_n27828_;
  assign new_n27830_ = pi0790 & ~new_n27829_;
  assign new_n27831_ = pi0644 & new_n27819_;
  assign new_n27832_ = ~pi0644 & new_n27827_;
  assign new_n27833_ = pi0790 & ~new_n27832_;
  assign new_n27834_ = ~new_n27831_ & new_n27833_;
  assign new_n27835_ = ~new_n20567_ & new_n27808_;
  assign new_n27836_ = ~pi0629 & new_n27730_;
  assign new_n27837_ = pi0629 & new_n27734_;
  assign new_n27838_ = ~new_n27836_ & ~new_n27837_;
  assign new_n27839_ = ~new_n27835_ & new_n27838_;
  assign new_n27840_ = pi0792 & ~new_n27839_;
  assign new_n27841_ = pi0725 & ~new_n27764_;
  assign new_n27842_ = ~pi0183 & new_n16810_;
  assign new_n27843_ = pi0183 & new_n16928_;
  assign new_n27844_ = pi0755 & ~new_n27843_;
  assign new_n27845_ = ~new_n27842_ & new_n27844_;
  assign new_n27846_ = pi0183 & new_n17007_;
  assign new_n27847_ = ~pi0183 & ~new_n17074_;
  assign new_n27848_ = ~pi0755 & ~new_n27847_;
  assign new_n27849_ = ~new_n27846_ & new_n27848_;
  assign new_n27850_ = pi0039 & ~new_n27849_;
  assign new_n27851_ = ~new_n27845_ & new_n27850_;
  assign new_n27852_ = ~pi0183 & ~new_n17217_;
  assign new_n27853_ = pi0183 & ~new_n17178_;
  assign new_n27854_ = pi0755 & ~new_n27853_;
  assign new_n27855_ = ~new_n27852_ & new_n27854_;
  assign new_n27856_ = ~pi0183 & new_n17227_;
  assign new_n27857_ = pi0183 & new_n17234_;
  assign new_n27858_ = ~pi0755 & ~new_n27857_;
  assign new_n27859_ = ~new_n27856_ & new_n27858_;
  assign new_n27860_ = ~new_n27855_ & ~new_n27859_;
  assign new_n27861_ = ~pi0039 & ~new_n27860_;
  assign new_n27862_ = ~pi0038 & ~new_n27861_;
  assign new_n27863_ = ~new_n27851_ & new_n27862_;
  assign new_n27864_ = ~pi0755 & ~new_n17035_;
  assign new_n27865_ = new_n19383_ & ~new_n27864_;
  assign new_n27866_ = ~pi0183 & ~new_n27865_;
  assign new_n27867_ = ~new_n16916_ & ~new_n27502_;
  assign new_n27868_ = pi0183 & ~new_n27867_;
  assign new_n27869_ = new_n6257_ & new_n27868_;
  assign new_n27870_ = pi0038 & ~new_n27869_;
  assign new_n27871_ = ~new_n27866_ & new_n27870_;
  assign new_n27872_ = ~pi0725 & ~new_n27871_;
  assign new_n27873_ = ~new_n27863_ & new_n27872_;
  assign new_n27874_ = new_n3272_ & ~new_n27873_;
  assign new_n27875_ = ~new_n27841_ & new_n27874_;
  assign new_n27876_ = ~new_n27752_ & ~new_n27875_;
  assign new_n27877_ = ~pi0625 & new_n27876_;
  assign new_n27878_ = pi0625 & new_n27766_;
  assign new_n27879_ = ~pi1153 & ~new_n27878_;
  assign new_n27880_ = ~new_n27877_ & new_n27879_;
  assign new_n27881_ = ~pi0608 & ~new_n27707_;
  assign new_n27882_ = ~new_n27880_ & new_n27881_;
  assign new_n27883_ = pi0625 & new_n27876_;
  assign new_n27884_ = ~pi0625 & new_n27766_;
  assign new_n27885_ = pi1153 & ~new_n27884_;
  assign new_n27886_ = ~new_n27883_ & new_n27885_;
  assign new_n27887_ = pi0608 & ~new_n27711_;
  assign new_n27888_ = ~new_n27886_ & new_n27887_;
  assign new_n27889_ = ~new_n27882_ & ~new_n27888_;
  assign new_n27890_ = pi0778 & ~new_n27889_;
  assign new_n27891_ = ~pi0778 & new_n27876_;
  assign new_n27892_ = ~new_n27890_ & ~new_n27891_;
  assign new_n27893_ = ~pi0609 & ~new_n27892_;
  assign new_n27894_ = pi0609 & new_n27714_;
  assign new_n27895_ = ~pi1155 & ~new_n27894_;
  assign new_n27896_ = ~new_n27893_ & new_n27895_;
  assign new_n27897_ = ~pi0660 & ~new_n27774_;
  assign new_n27898_ = ~new_n27896_ & new_n27897_;
  assign new_n27899_ = pi0609 & ~new_n27892_;
  assign new_n27900_ = ~pi0609 & new_n27714_;
  assign new_n27901_ = pi1155 & ~new_n27900_;
  assign new_n27902_ = ~new_n27899_ & new_n27901_;
  assign new_n27903_ = pi0660 & ~new_n27778_;
  assign new_n27904_ = ~new_n27902_ & new_n27903_;
  assign new_n27905_ = ~new_n27898_ & ~new_n27904_;
  assign new_n27906_ = pi0785 & ~new_n27905_;
  assign new_n27907_ = ~pi0785 & ~new_n27892_;
  assign new_n27908_ = ~new_n27906_ & ~new_n27907_;
  assign new_n27909_ = ~pi0618 & ~new_n27908_;
  assign new_n27910_ = pi0618 & new_n27717_;
  assign new_n27911_ = ~pi1154 & ~new_n27910_;
  assign new_n27912_ = ~new_n27909_ & new_n27911_;
  assign new_n27913_ = ~pi0627 & ~new_n27786_;
  assign new_n27914_ = ~new_n27912_ & new_n27913_;
  assign new_n27915_ = pi0618 & ~new_n27908_;
  assign new_n27916_ = ~pi0618 & new_n27717_;
  assign new_n27917_ = pi1154 & ~new_n27916_;
  assign new_n27918_ = ~new_n27915_ & new_n27917_;
  assign new_n27919_ = pi0627 & ~new_n27790_;
  assign new_n27920_ = ~new_n27918_ & new_n27919_;
  assign new_n27921_ = ~new_n27914_ & ~new_n27920_;
  assign new_n27922_ = pi0781 & ~new_n27921_;
  assign new_n27923_ = ~pi0781 & ~new_n27908_;
  assign new_n27924_ = ~new_n27922_ & ~new_n27923_;
  assign new_n27925_ = pi0619 & ~new_n27924_;
  assign new_n27926_ = ~pi0619 & ~new_n27720_;
  assign new_n27927_ = pi1159 & ~new_n27926_;
  assign new_n27928_ = ~new_n27925_ & new_n27927_;
  assign new_n27929_ = pi0648 & ~new_n27802_;
  assign new_n27930_ = ~new_n27928_ & new_n27929_;
  assign new_n27931_ = ~pi0619 & ~new_n27924_;
  assign new_n27932_ = pi0619 & ~new_n27720_;
  assign new_n27933_ = ~pi1159 & ~new_n27932_;
  assign new_n27934_ = ~new_n27931_ & new_n27933_;
  assign new_n27935_ = ~pi0648 & ~new_n27798_;
  assign new_n27936_ = ~new_n27934_ & new_n27935_;
  assign new_n27937_ = pi0789 & ~new_n27936_;
  assign new_n27938_ = ~new_n27930_ & new_n27937_;
  assign new_n27939_ = ~pi0789 & new_n27924_;
  assign new_n27940_ = new_n17969_ & ~new_n27939_;
  assign new_n27941_ = ~new_n27938_ & new_n27940_;
  assign new_n27942_ = pi0626 & ~new_n27805_;
  assign new_n27943_ = ~pi0626 & ~new_n27689_;
  assign new_n27944_ = new_n17731_ & ~new_n27943_;
  assign new_n27945_ = ~new_n27942_ & new_n27944_;
  assign new_n27946_ = new_n17856_ & new_n27722_;
  assign new_n27947_ = ~pi0626 & ~new_n27805_;
  assign new_n27948_ = pi0626 & ~new_n27689_;
  assign new_n27949_ = new_n17732_ & ~new_n27948_;
  assign new_n27950_ = ~new_n27947_ & new_n27949_;
  assign new_n27951_ = ~new_n27946_ & ~new_n27950_;
  assign new_n27952_ = ~new_n27945_ & new_n27951_;
  assign new_n27953_ = pi0788 & ~new_n27952_;
  assign new_n27954_ = ~new_n20364_ & ~new_n27953_;
  assign new_n27955_ = ~new_n27941_ & new_n27954_;
  assign new_n27956_ = ~new_n27840_ & ~new_n27955_;
  assign new_n27957_ = ~new_n20360_ & ~new_n27956_;
  assign new_n27958_ = ~new_n20556_ & new_n27811_;
  assign new_n27959_ = new_n17802_ & ~new_n27740_;
  assign new_n27960_ = new_n17801_ & ~new_n27744_;
  assign new_n27961_ = ~new_n27959_ & ~new_n27960_;
  assign new_n27962_ = ~new_n27958_ & new_n27961_;
  assign new_n27963_ = pi0787 & ~new_n27962_;
  assign new_n27964_ = ~new_n27957_ & ~new_n27963_;
  assign new_n27965_ = ~new_n27834_ & new_n27964_;
  assign new_n27966_ = ~new_n27830_ & ~new_n27965_;
  assign new_n27967_ = ~po1038 & ~new_n27966_;
  assign new_n27968_ = ~pi0183 & po1038;
  assign new_n27969_ = ~pi0832 & ~new_n27968_;
  assign new_n27970_ = ~new_n27967_ & new_n27969_;
  assign po0340 = ~new_n27688_ & ~new_n27970_;
  assign new_n27972_ = ~pi0184 & ~new_n2754_;
  assign new_n27973_ = ~pi0777 & new_n16913_;
  assign new_n27974_ = ~new_n27972_ & ~new_n27973_;
  assign new_n27975_ = ~new_n17858_ & ~new_n27974_;
  assign new_n27976_ = ~pi0785 & ~new_n27975_;
  assign new_n27977_ = new_n17603_ & new_n27973_;
  assign new_n27978_ = new_n27975_ & ~new_n27977_;
  assign new_n27979_ = pi1155 & ~new_n27978_;
  assign new_n27980_ = ~pi1155 & ~new_n27972_;
  assign new_n27981_ = ~new_n27977_ & new_n27980_;
  assign new_n27982_ = ~new_n27979_ & ~new_n27981_;
  assign new_n27983_ = pi0785 & ~new_n27982_;
  assign new_n27984_ = ~new_n27976_ & ~new_n27983_;
  assign new_n27985_ = ~pi0781 & ~new_n27984_;
  assign new_n27986_ = ~new_n17873_ & new_n27984_;
  assign new_n27987_ = pi1154 & ~new_n27986_;
  assign new_n27988_ = ~new_n17876_ & new_n27984_;
  assign new_n27989_ = ~pi1154 & ~new_n27988_;
  assign new_n27990_ = ~new_n27987_ & ~new_n27989_;
  assign new_n27991_ = pi0781 & ~new_n27990_;
  assign new_n27992_ = ~new_n27985_ & ~new_n27991_;
  assign new_n27993_ = ~pi0789 & ~new_n27992_;
  assign new_n27994_ = ~new_n23057_ & new_n27992_;
  assign new_n27995_ = pi1159 & ~new_n27994_;
  assign new_n27996_ = ~new_n23060_ & new_n27992_;
  assign new_n27997_ = ~pi1159 & ~new_n27996_;
  assign new_n27998_ = ~new_n27995_ & ~new_n27997_;
  assign new_n27999_ = pi0789 & ~new_n27998_;
  assign new_n28000_ = ~new_n27993_ & ~new_n27999_;
  assign new_n28001_ = ~new_n17968_ & new_n28000_;
  assign new_n28002_ = new_n17968_ & new_n27972_;
  assign new_n28003_ = ~new_n28001_ & ~new_n28002_;
  assign new_n28004_ = ~new_n17762_ & ~new_n28003_;
  assign new_n28005_ = new_n17762_ & new_n27972_;
  assign new_n28006_ = ~new_n28004_ & ~new_n28005_;
  assign new_n28007_ = ~new_n20556_ & new_n28006_;
  assign new_n28008_ = ~pi0737 & new_n16915_;
  assign new_n28009_ = ~new_n27972_ & ~new_n28008_;
  assign new_n28010_ = ~pi0778 & ~new_n28009_;
  assign new_n28011_ = ~pi0625 & new_n28008_;
  assign new_n28012_ = ~new_n28009_ & ~new_n28011_;
  assign new_n28013_ = pi1153 & ~new_n28012_;
  assign new_n28014_ = ~pi1153 & ~new_n27972_;
  assign new_n28015_ = ~new_n28011_ & new_n28014_;
  assign new_n28016_ = pi0778 & ~new_n28015_;
  assign new_n28017_ = ~new_n28013_ & new_n28016_;
  assign new_n28018_ = ~new_n28010_ & ~new_n28017_;
  assign new_n28019_ = ~new_n17844_ & ~new_n28018_;
  assign new_n28020_ = ~new_n17846_ & new_n28019_;
  assign new_n28021_ = ~new_n17848_ & new_n28020_;
  assign new_n28022_ = ~new_n17980_ & new_n28021_;
  assign new_n28023_ = ~new_n18011_ & new_n28022_;
  assign new_n28024_ = ~pi0647 & new_n28023_;
  assign new_n28025_ = pi0647 & new_n27972_;
  assign new_n28026_ = ~pi1157 & ~new_n28025_;
  assign new_n28027_ = ~new_n28024_ & new_n28026_;
  assign new_n28028_ = pi0630 & new_n28027_;
  assign new_n28029_ = pi0647 & ~new_n28023_;
  assign new_n28030_ = ~pi0647 & ~new_n27972_;
  assign new_n28031_ = ~new_n28029_ & ~new_n28030_;
  assign new_n28032_ = new_n17801_ & ~new_n28031_;
  assign new_n28033_ = ~new_n28028_ & ~new_n28032_;
  assign new_n28034_ = ~new_n28007_ & new_n28033_;
  assign new_n28035_ = pi0787 & ~new_n28034_;
  assign new_n28036_ = pi0626 & ~new_n28000_;
  assign new_n28037_ = ~pi0626 & ~new_n27972_;
  assign new_n28038_ = new_n17731_ & ~new_n28037_;
  assign new_n28039_ = ~new_n28036_ & new_n28038_;
  assign new_n28040_ = new_n17856_ & new_n28021_;
  assign new_n28041_ = ~pi0626 & ~new_n28000_;
  assign new_n28042_ = pi0626 & ~new_n27972_;
  assign new_n28043_ = new_n17732_ & ~new_n28042_;
  assign new_n28044_ = ~new_n28041_ & new_n28043_;
  assign new_n28045_ = ~new_n28040_ & ~new_n28044_;
  assign new_n28046_ = ~new_n28039_ & new_n28045_;
  assign new_n28047_ = pi0788 & ~new_n28046_;
  assign new_n28048_ = ~new_n16639_ & ~new_n28009_;
  assign new_n28049_ = pi0625 & new_n28048_;
  assign new_n28050_ = new_n27974_ & ~new_n28048_;
  assign new_n28051_ = ~new_n28049_ & ~new_n28050_;
  assign new_n28052_ = new_n28014_ & ~new_n28051_;
  assign new_n28053_ = ~pi0608 & ~new_n28013_;
  assign new_n28054_ = ~new_n28052_ & new_n28053_;
  assign new_n28055_ = pi1153 & new_n27974_;
  assign new_n28056_ = ~new_n28049_ & new_n28055_;
  assign new_n28057_ = pi0608 & ~new_n28015_;
  assign new_n28058_ = ~new_n28056_ & new_n28057_;
  assign new_n28059_ = ~new_n28054_ & ~new_n28058_;
  assign new_n28060_ = pi0778 & ~new_n28059_;
  assign new_n28061_ = ~pi0778 & ~new_n28050_;
  assign new_n28062_ = ~new_n28060_ & ~new_n28061_;
  assign new_n28063_ = ~pi0609 & ~new_n28062_;
  assign new_n28064_ = pi0609 & ~new_n28018_;
  assign new_n28065_ = ~pi1155 & ~new_n28064_;
  assign new_n28066_ = ~new_n28063_ & new_n28065_;
  assign new_n28067_ = ~pi0660 & ~new_n27979_;
  assign new_n28068_ = ~new_n28066_ & new_n28067_;
  assign new_n28069_ = pi0609 & ~new_n28062_;
  assign new_n28070_ = ~pi0609 & ~new_n28018_;
  assign new_n28071_ = pi1155 & ~new_n28070_;
  assign new_n28072_ = ~new_n28069_ & new_n28071_;
  assign new_n28073_ = pi0660 & ~new_n27981_;
  assign new_n28074_ = ~new_n28072_ & new_n28073_;
  assign new_n28075_ = ~new_n28068_ & ~new_n28074_;
  assign new_n28076_ = pi0785 & ~new_n28075_;
  assign new_n28077_ = ~pi0785 & ~new_n28062_;
  assign new_n28078_ = ~new_n28076_ & ~new_n28077_;
  assign new_n28079_ = ~pi0618 & ~new_n28078_;
  assign new_n28080_ = pi0618 & new_n28019_;
  assign new_n28081_ = ~pi1154 & ~new_n28080_;
  assign new_n28082_ = ~new_n28079_ & new_n28081_;
  assign new_n28083_ = ~pi0627 & ~new_n27987_;
  assign new_n28084_ = ~new_n28082_ & new_n28083_;
  assign new_n28085_ = pi0618 & ~new_n28078_;
  assign new_n28086_ = ~pi0618 & new_n28019_;
  assign new_n28087_ = pi1154 & ~new_n28086_;
  assign new_n28088_ = ~new_n28085_ & new_n28087_;
  assign new_n28089_ = pi0627 & ~new_n27989_;
  assign new_n28090_ = ~new_n28088_ & new_n28089_;
  assign new_n28091_ = ~new_n28084_ & ~new_n28090_;
  assign new_n28092_ = pi0781 & ~new_n28091_;
  assign new_n28093_ = ~pi0781 & ~new_n28078_;
  assign new_n28094_ = ~new_n28092_ & ~new_n28093_;
  assign new_n28095_ = pi0619 & ~new_n28094_;
  assign new_n28096_ = ~pi0619 & new_n28020_;
  assign new_n28097_ = pi1159 & ~new_n28096_;
  assign new_n28098_ = ~new_n28095_ & new_n28097_;
  assign new_n28099_ = pi0648 & ~new_n27997_;
  assign new_n28100_ = ~new_n28098_ & new_n28099_;
  assign new_n28101_ = ~pi0619 & ~new_n28094_;
  assign new_n28102_ = pi0619 & new_n28020_;
  assign new_n28103_ = ~pi1159 & ~new_n28102_;
  assign new_n28104_ = ~new_n28101_ & new_n28103_;
  assign new_n28105_ = ~pi0648 & ~new_n27995_;
  assign new_n28106_ = ~new_n28104_ & new_n28105_;
  assign new_n28107_ = pi0789 & ~new_n28106_;
  assign new_n28108_ = ~new_n28100_ & new_n28107_;
  assign new_n28109_ = ~pi0789 & new_n28094_;
  assign new_n28110_ = new_n17969_ & ~new_n28109_;
  assign new_n28111_ = ~new_n28108_ & new_n28110_;
  assign new_n28112_ = ~new_n28047_ & ~new_n28111_;
  assign new_n28113_ = ~new_n20364_ & ~new_n28112_;
  assign new_n28114_ = new_n18008_ & ~new_n28003_;
  assign new_n28115_ = new_n20851_ & new_n28022_;
  assign new_n28116_ = ~new_n28114_ & ~new_n28115_;
  assign new_n28117_ = ~pi0629 & ~new_n28116_;
  assign new_n28118_ = new_n20855_ & new_n28022_;
  assign new_n28119_ = new_n18007_ & ~new_n28003_;
  assign new_n28120_ = ~new_n28118_ & ~new_n28119_;
  assign new_n28121_ = pi0629 & ~new_n28120_;
  assign new_n28122_ = ~new_n28117_ & ~new_n28121_;
  assign new_n28123_ = pi0792 & ~new_n28122_;
  assign new_n28124_ = ~new_n20360_ & ~new_n28123_;
  assign new_n28125_ = ~new_n28113_ & new_n28124_;
  assign new_n28126_ = ~new_n28035_ & ~new_n28125_;
  assign new_n28127_ = pi0644 & new_n28126_;
  assign new_n28128_ = ~pi0787 & ~new_n28023_;
  assign new_n28129_ = pi1157 & ~new_n28031_;
  assign new_n28130_ = ~new_n28027_ & ~new_n28129_;
  assign new_n28131_ = pi0787 & ~new_n28130_;
  assign new_n28132_ = ~new_n28128_ & ~new_n28131_;
  assign new_n28133_ = ~pi0644 & new_n28132_;
  assign new_n28134_ = pi0715 & ~new_n28133_;
  assign new_n28135_ = ~new_n28127_ & new_n28134_;
  assign new_n28136_ = ~new_n17804_ & ~new_n28006_;
  assign new_n28137_ = new_n17804_ & new_n27972_;
  assign new_n28138_ = ~new_n28136_ & ~new_n28137_;
  assign new_n28139_ = pi0644 & ~new_n28138_;
  assign new_n28140_ = ~pi0644 & new_n27972_;
  assign new_n28141_ = ~pi0715 & ~new_n28140_;
  assign new_n28142_ = ~new_n28139_ & new_n28141_;
  assign new_n28143_ = pi1160 & ~new_n28142_;
  assign new_n28144_ = ~new_n28135_ & new_n28143_;
  assign new_n28145_ = ~pi0644 & new_n28126_;
  assign new_n28146_ = pi0644 & new_n28132_;
  assign new_n28147_ = ~pi0715 & ~new_n28146_;
  assign new_n28148_ = ~new_n28145_ & new_n28147_;
  assign new_n28149_ = ~pi0644 & ~new_n28138_;
  assign new_n28150_ = pi0644 & new_n27972_;
  assign new_n28151_ = pi0715 & ~new_n28150_;
  assign new_n28152_ = ~new_n28149_ & new_n28151_;
  assign new_n28153_ = ~pi1160 & ~new_n28152_;
  assign new_n28154_ = ~new_n28148_ & new_n28153_;
  assign new_n28155_ = ~new_n28144_ & ~new_n28154_;
  assign new_n28156_ = pi0790 & ~new_n28155_;
  assign new_n28157_ = ~pi0790 & new_n28126_;
  assign new_n28158_ = pi0832 & ~new_n28157_;
  assign new_n28159_ = ~new_n28156_ & new_n28158_;
  assign new_n28160_ = ~pi0184 & ~new_n17558_;
  assign new_n28161_ = new_n17691_ & ~new_n28160_;
  assign new_n28162_ = ~pi0737 & new_n3272_;
  assign new_n28163_ = new_n28160_ & ~new_n28162_;
  assign new_n28164_ = pi0184 & ~new_n18128_;
  assign new_n28165_ = ~pi0038 & ~new_n28164_;
  assign new_n28166_ = new_n3272_ & ~new_n28165_;
  assign new_n28167_ = ~pi0184 & new_n18124_;
  assign new_n28168_ = ~new_n28166_ & ~new_n28167_;
  assign new_n28169_ = ~pi0184 & ~new_n17431_;
  assign new_n28170_ = new_n17544_ & ~new_n28169_;
  assign new_n28171_ = ~pi0737 & ~new_n28170_;
  assign new_n28172_ = ~new_n28168_ & new_n28171_;
  assign new_n28173_ = ~new_n28163_ & ~new_n28172_;
  assign new_n28174_ = ~pi0778 & new_n28173_;
  assign new_n28175_ = pi0625 & ~new_n28173_;
  assign new_n28176_ = ~pi0625 & new_n28160_;
  assign new_n28177_ = pi1153 & ~new_n28176_;
  assign new_n28178_ = ~new_n28175_ & new_n28177_;
  assign new_n28179_ = ~pi0625 & ~new_n28173_;
  assign new_n28180_ = pi0625 & new_n28160_;
  assign new_n28181_ = ~pi1153 & ~new_n28180_;
  assign new_n28182_ = ~new_n28179_ & new_n28181_;
  assign new_n28183_ = ~new_n28178_ & ~new_n28182_;
  assign new_n28184_ = pi0778 & ~new_n28183_;
  assign new_n28185_ = ~new_n28174_ & ~new_n28184_;
  assign new_n28186_ = ~new_n17618_ & ~new_n28185_;
  assign new_n28187_ = new_n17618_ & ~new_n28160_;
  assign new_n28188_ = ~new_n28186_ & ~new_n28187_;
  assign new_n28189_ = ~new_n17655_ & new_n28188_;
  assign new_n28190_ = new_n17655_ & new_n28160_;
  assign new_n28191_ = ~new_n28189_ & ~new_n28190_;
  assign new_n28192_ = ~new_n17691_ & new_n28191_;
  assign new_n28193_ = ~new_n28161_ & ~new_n28192_;
  assign new_n28194_ = ~new_n17734_ & new_n28193_;
  assign new_n28195_ = new_n17734_ & new_n28160_;
  assign new_n28196_ = ~new_n28194_ & ~new_n28195_;
  assign new_n28197_ = ~pi0792 & new_n28196_;
  assign new_n28198_ = pi0628 & ~new_n28196_;
  assign new_n28199_ = ~pi0628 & new_n28160_;
  assign new_n28200_ = pi1156 & ~new_n28199_;
  assign new_n28201_ = ~new_n28198_ & new_n28200_;
  assign new_n28202_ = ~pi0628 & ~new_n28196_;
  assign new_n28203_ = pi0628 & new_n28160_;
  assign new_n28204_ = ~pi1156 & ~new_n28203_;
  assign new_n28205_ = ~new_n28202_ & new_n28204_;
  assign new_n28206_ = ~new_n28201_ & ~new_n28205_;
  assign new_n28207_ = pi0792 & ~new_n28206_;
  assign new_n28208_ = ~new_n28197_ & ~new_n28207_;
  assign new_n28209_ = ~pi0647 & ~new_n28208_;
  assign new_n28210_ = pi0647 & ~new_n28160_;
  assign new_n28211_ = ~new_n28209_ & ~new_n28210_;
  assign new_n28212_ = ~pi1157 & new_n28211_;
  assign new_n28213_ = pi0647 & ~new_n28208_;
  assign new_n28214_ = ~pi0647 & ~new_n28160_;
  assign new_n28215_ = ~new_n28213_ & ~new_n28214_;
  assign new_n28216_ = pi1157 & new_n28215_;
  assign new_n28217_ = ~new_n28212_ & ~new_n28216_;
  assign new_n28218_ = pi0787 & ~new_n28217_;
  assign new_n28219_ = ~pi0787 & new_n28208_;
  assign new_n28220_ = ~new_n28218_ & ~new_n28219_;
  assign new_n28221_ = ~pi0644 & ~new_n28220_;
  assign new_n28222_ = pi0715 & ~new_n28221_;
  assign new_n28223_ = pi0184 & ~new_n3272_;
  assign new_n28224_ = ~pi0777 & new_n17433_;
  assign new_n28225_ = ~new_n28169_ & ~new_n28224_;
  assign new_n28226_ = pi0038 & ~new_n28225_;
  assign new_n28227_ = ~pi0184 & new_n17393_;
  assign new_n28228_ = pi0184 & ~new_n17426_;
  assign new_n28229_ = ~pi0777 & ~new_n28228_;
  assign new_n28230_ = ~new_n28227_ & new_n28229_;
  assign new_n28231_ = ~pi0184 & pi0777;
  assign new_n28232_ = ~new_n17349_ & new_n28231_;
  assign new_n28233_ = ~new_n28230_ & ~new_n28232_;
  assign new_n28234_ = ~pi0038 & ~new_n28233_;
  assign new_n28235_ = ~new_n28226_ & ~new_n28234_;
  assign new_n28236_ = new_n3272_ & new_n28235_;
  assign new_n28237_ = ~new_n28223_ & ~new_n28236_;
  assign new_n28238_ = ~new_n17590_ & ~new_n28237_;
  assign new_n28239_ = new_n17590_ & ~new_n28160_;
  assign new_n28240_ = ~new_n28238_ & ~new_n28239_;
  assign new_n28241_ = ~pi0785 & ~new_n28240_;
  assign new_n28242_ = ~new_n17591_ & ~new_n28160_;
  assign new_n28243_ = pi0609 & new_n28238_;
  assign new_n28244_ = ~new_n28242_ & ~new_n28243_;
  assign new_n28245_ = pi1155 & ~new_n28244_;
  assign new_n28246_ = ~new_n17603_ & ~new_n28160_;
  assign new_n28247_ = ~pi0609 & new_n28238_;
  assign new_n28248_ = ~new_n28246_ & ~new_n28247_;
  assign new_n28249_ = ~pi1155 & ~new_n28248_;
  assign new_n28250_ = ~new_n28245_ & ~new_n28249_;
  assign new_n28251_ = pi0785 & ~new_n28250_;
  assign new_n28252_ = ~new_n28241_ & ~new_n28251_;
  assign new_n28253_ = ~pi0781 & ~new_n28252_;
  assign new_n28254_ = pi0618 & new_n28252_;
  assign new_n28255_ = ~pi0618 & new_n28160_;
  assign new_n28256_ = pi1154 & ~new_n28255_;
  assign new_n28257_ = ~new_n28254_ & new_n28256_;
  assign new_n28258_ = ~pi0618 & new_n28252_;
  assign new_n28259_ = pi0618 & new_n28160_;
  assign new_n28260_ = ~pi1154 & ~new_n28259_;
  assign new_n28261_ = ~new_n28258_ & new_n28260_;
  assign new_n28262_ = ~new_n28257_ & ~new_n28261_;
  assign new_n28263_ = pi0781 & ~new_n28262_;
  assign new_n28264_ = ~new_n28253_ & ~new_n28263_;
  assign new_n28265_ = ~pi0789 & ~new_n28264_;
  assign new_n28266_ = pi0619 & new_n28264_;
  assign new_n28267_ = ~pi0619 & new_n28160_;
  assign new_n28268_ = pi1159 & ~new_n28267_;
  assign new_n28269_ = ~new_n28266_ & new_n28268_;
  assign new_n28270_ = ~pi0619 & new_n28264_;
  assign new_n28271_ = pi0619 & new_n28160_;
  assign new_n28272_ = ~pi1159 & ~new_n28271_;
  assign new_n28273_ = ~new_n28270_ & new_n28272_;
  assign new_n28274_ = ~new_n28269_ & ~new_n28273_;
  assign new_n28275_ = pi0789 & ~new_n28274_;
  assign new_n28276_ = ~new_n28265_ & ~new_n28275_;
  assign new_n28277_ = ~new_n17968_ & new_n28276_;
  assign new_n28278_ = new_n17968_ & new_n28160_;
  assign new_n28279_ = ~new_n28277_ & ~new_n28278_;
  assign new_n28280_ = ~new_n17762_ & ~new_n28279_;
  assign new_n28281_ = new_n17762_ & new_n28160_;
  assign new_n28282_ = ~new_n28280_ & ~new_n28281_;
  assign new_n28283_ = ~new_n17804_ & ~new_n28282_;
  assign new_n28284_ = new_n17804_ & new_n28160_;
  assign new_n28285_ = ~new_n28283_ & ~new_n28284_;
  assign new_n28286_ = pi0644 & ~new_n28285_;
  assign new_n28287_ = ~pi0644 & new_n28160_;
  assign new_n28288_ = ~pi0715 & ~new_n28287_;
  assign new_n28289_ = ~new_n28286_ & new_n28288_;
  assign new_n28290_ = pi1160 & ~new_n28289_;
  assign new_n28291_ = ~new_n28222_ & new_n28290_;
  assign new_n28292_ = pi0644 & ~new_n28220_;
  assign new_n28293_ = ~pi0715 & ~new_n28292_;
  assign new_n28294_ = ~pi0644 & ~new_n28285_;
  assign new_n28295_ = pi0644 & new_n28160_;
  assign new_n28296_ = pi0715 & ~new_n28295_;
  assign new_n28297_ = ~new_n28294_ & new_n28296_;
  assign new_n28298_ = ~pi1160 & ~new_n28297_;
  assign new_n28299_ = ~new_n28293_ & new_n28298_;
  assign new_n28300_ = ~new_n28291_ & ~new_n28299_;
  assign new_n28301_ = pi0790 & ~new_n28300_;
  assign new_n28302_ = pi0644 & new_n28290_;
  assign new_n28303_ = ~pi0644 & new_n28298_;
  assign new_n28304_ = pi0790 & ~new_n28303_;
  assign new_n28305_ = ~new_n28302_ & new_n28304_;
  assign new_n28306_ = ~new_n20567_ & new_n28279_;
  assign new_n28307_ = ~pi0629 & new_n28201_;
  assign new_n28308_ = pi0629 & new_n28205_;
  assign new_n28309_ = ~new_n28307_ & ~new_n28308_;
  assign new_n28310_ = ~new_n28306_ & new_n28309_;
  assign new_n28311_ = pi0792 & ~new_n28310_;
  assign new_n28312_ = pi0737 & ~new_n28235_;
  assign new_n28313_ = ~pi0184 & new_n16810_;
  assign new_n28314_ = pi0184 & new_n16928_;
  assign new_n28315_ = pi0777 & ~new_n28314_;
  assign new_n28316_ = ~new_n28313_ & new_n28315_;
  assign new_n28317_ = pi0184 & new_n17007_;
  assign new_n28318_ = ~pi0184 & ~new_n17074_;
  assign new_n28319_ = ~pi0777 & ~new_n28318_;
  assign new_n28320_ = ~new_n28317_ & new_n28319_;
  assign new_n28321_ = pi0039 & ~new_n28320_;
  assign new_n28322_ = ~new_n28316_ & new_n28321_;
  assign new_n28323_ = ~pi0184 & ~new_n17217_;
  assign new_n28324_ = pi0184 & ~new_n17178_;
  assign new_n28325_ = pi0777 & ~new_n28324_;
  assign new_n28326_ = ~new_n28323_ & new_n28325_;
  assign new_n28327_ = ~pi0184 & new_n17227_;
  assign new_n28328_ = pi0184 & new_n17234_;
  assign new_n28329_ = ~pi0777 & ~new_n28328_;
  assign new_n28330_ = ~new_n28327_ & new_n28329_;
  assign new_n28331_ = ~new_n28326_ & ~new_n28330_;
  assign new_n28332_ = ~pi0039 & ~new_n28331_;
  assign new_n28333_ = ~pi0038 & ~new_n28332_;
  assign new_n28334_ = ~new_n28322_ & new_n28333_;
  assign new_n28335_ = ~pi0777 & ~new_n17035_;
  assign new_n28336_ = new_n19383_ & ~new_n28335_;
  assign new_n28337_ = ~pi0184 & ~new_n28336_;
  assign new_n28338_ = ~new_n16916_ & ~new_n27973_;
  assign new_n28339_ = pi0184 & ~new_n28338_;
  assign new_n28340_ = new_n6257_ & new_n28339_;
  assign new_n28341_ = pi0038 & ~new_n28340_;
  assign new_n28342_ = ~new_n28337_ & new_n28341_;
  assign new_n28343_ = ~pi0737 & ~new_n28342_;
  assign new_n28344_ = ~new_n28334_ & new_n28343_;
  assign new_n28345_ = new_n3272_ & ~new_n28344_;
  assign new_n28346_ = ~new_n28312_ & new_n28345_;
  assign new_n28347_ = ~new_n28223_ & ~new_n28346_;
  assign new_n28348_ = ~pi0625 & new_n28347_;
  assign new_n28349_ = pi0625 & new_n28237_;
  assign new_n28350_ = ~pi1153 & ~new_n28349_;
  assign new_n28351_ = ~new_n28348_ & new_n28350_;
  assign new_n28352_ = ~pi0608 & ~new_n28178_;
  assign new_n28353_ = ~new_n28351_ & new_n28352_;
  assign new_n28354_ = pi0625 & new_n28347_;
  assign new_n28355_ = ~pi0625 & new_n28237_;
  assign new_n28356_ = pi1153 & ~new_n28355_;
  assign new_n28357_ = ~new_n28354_ & new_n28356_;
  assign new_n28358_ = pi0608 & ~new_n28182_;
  assign new_n28359_ = ~new_n28357_ & new_n28358_;
  assign new_n28360_ = ~new_n28353_ & ~new_n28359_;
  assign new_n28361_ = pi0778 & ~new_n28360_;
  assign new_n28362_ = ~pi0778 & new_n28347_;
  assign new_n28363_ = ~new_n28361_ & ~new_n28362_;
  assign new_n28364_ = ~pi0609 & ~new_n28363_;
  assign new_n28365_ = pi0609 & new_n28185_;
  assign new_n28366_ = ~pi1155 & ~new_n28365_;
  assign new_n28367_ = ~new_n28364_ & new_n28366_;
  assign new_n28368_ = ~pi0660 & ~new_n28245_;
  assign new_n28369_ = ~new_n28367_ & new_n28368_;
  assign new_n28370_ = pi0609 & ~new_n28363_;
  assign new_n28371_ = ~pi0609 & new_n28185_;
  assign new_n28372_ = pi1155 & ~new_n28371_;
  assign new_n28373_ = ~new_n28370_ & new_n28372_;
  assign new_n28374_ = pi0660 & ~new_n28249_;
  assign new_n28375_ = ~new_n28373_ & new_n28374_;
  assign new_n28376_ = ~new_n28369_ & ~new_n28375_;
  assign new_n28377_ = pi0785 & ~new_n28376_;
  assign new_n28378_ = ~pi0785 & ~new_n28363_;
  assign new_n28379_ = ~new_n28377_ & ~new_n28378_;
  assign new_n28380_ = ~pi0618 & ~new_n28379_;
  assign new_n28381_ = pi0618 & new_n28188_;
  assign new_n28382_ = ~pi1154 & ~new_n28381_;
  assign new_n28383_ = ~new_n28380_ & new_n28382_;
  assign new_n28384_ = ~pi0627 & ~new_n28257_;
  assign new_n28385_ = ~new_n28383_ & new_n28384_;
  assign new_n28386_ = pi0618 & ~new_n28379_;
  assign new_n28387_ = ~pi0618 & new_n28188_;
  assign new_n28388_ = pi1154 & ~new_n28387_;
  assign new_n28389_ = ~new_n28386_ & new_n28388_;
  assign new_n28390_ = pi0627 & ~new_n28261_;
  assign new_n28391_ = ~new_n28389_ & new_n28390_;
  assign new_n28392_ = ~new_n28385_ & ~new_n28391_;
  assign new_n28393_ = pi0781 & ~new_n28392_;
  assign new_n28394_ = ~pi0781 & ~new_n28379_;
  assign new_n28395_ = ~new_n28393_ & ~new_n28394_;
  assign new_n28396_ = pi0619 & ~new_n28395_;
  assign new_n28397_ = ~pi0619 & ~new_n28191_;
  assign new_n28398_ = pi1159 & ~new_n28397_;
  assign new_n28399_ = ~new_n28396_ & new_n28398_;
  assign new_n28400_ = pi0648 & ~new_n28273_;
  assign new_n28401_ = ~new_n28399_ & new_n28400_;
  assign new_n28402_ = ~pi0619 & ~new_n28395_;
  assign new_n28403_ = pi0619 & ~new_n28191_;
  assign new_n28404_ = ~pi1159 & ~new_n28403_;
  assign new_n28405_ = ~new_n28402_ & new_n28404_;
  assign new_n28406_ = ~pi0648 & ~new_n28269_;
  assign new_n28407_ = ~new_n28405_ & new_n28406_;
  assign new_n28408_ = pi0789 & ~new_n28407_;
  assign new_n28409_ = ~new_n28401_ & new_n28408_;
  assign new_n28410_ = ~pi0789 & new_n28395_;
  assign new_n28411_ = new_n17969_ & ~new_n28410_;
  assign new_n28412_ = ~new_n28409_ & new_n28411_;
  assign new_n28413_ = pi0626 & ~new_n28276_;
  assign new_n28414_ = ~pi0626 & ~new_n28160_;
  assign new_n28415_ = new_n17731_ & ~new_n28414_;
  assign new_n28416_ = ~new_n28413_ & new_n28415_;
  assign new_n28417_ = new_n17856_ & new_n28193_;
  assign new_n28418_ = ~pi0626 & ~new_n28276_;
  assign new_n28419_ = pi0626 & ~new_n28160_;
  assign new_n28420_ = new_n17732_ & ~new_n28419_;
  assign new_n28421_ = ~new_n28418_ & new_n28420_;
  assign new_n28422_ = ~new_n28417_ & ~new_n28421_;
  assign new_n28423_ = ~new_n28416_ & new_n28422_;
  assign new_n28424_ = pi0788 & ~new_n28423_;
  assign new_n28425_ = ~new_n20364_ & ~new_n28424_;
  assign new_n28426_ = ~new_n28412_ & new_n28425_;
  assign new_n28427_ = ~new_n28311_ & ~new_n28426_;
  assign new_n28428_ = ~new_n20360_ & ~new_n28427_;
  assign new_n28429_ = ~new_n20556_ & new_n28282_;
  assign new_n28430_ = new_n17802_ & ~new_n28211_;
  assign new_n28431_ = new_n17801_ & ~new_n28215_;
  assign new_n28432_ = ~new_n28430_ & ~new_n28431_;
  assign new_n28433_ = ~new_n28429_ & new_n28432_;
  assign new_n28434_ = pi0787 & ~new_n28433_;
  assign new_n28435_ = ~new_n28428_ & ~new_n28434_;
  assign new_n28436_ = ~new_n28305_ & new_n28435_;
  assign new_n28437_ = ~new_n28301_ & ~new_n28436_;
  assign new_n28438_ = ~po1038 & ~new_n28437_;
  assign new_n28439_ = ~pi0184 & po1038;
  assign new_n28440_ = ~pi0832 & ~new_n28439_;
  assign new_n28441_ = ~new_n28438_ & new_n28440_;
  assign po0341 = ~new_n28159_ & ~new_n28441_;
  assign new_n28443_ = ~pi0185 & ~new_n2754_;
  assign new_n28444_ = ~pi0751 & new_n16913_;
  assign new_n28445_ = ~new_n28443_ & ~new_n28444_;
  assign new_n28446_ = ~new_n17858_ & ~new_n28445_;
  assign new_n28447_ = ~pi0785 & ~new_n28446_;
  assign new_n28448_ = new_n17603_ & new_n28444_;
  assign new_n28449_ = new_n28446_ & ~new_n28448_;
  assign new_n28450_ = pi1155 & ~new_n28449_;
  assign new_n28451_ = ~pi1155 & ~new_n28443_;
  assign new_n28452_ = ~new_n28448_ & new_n28451_;
  assign new_n28453_ = ~new_n28450_ & ~new_n28452_;
  assign new_n28454_ = pi0785 & ~new_n28453_;
  assign new_n28455_ = ~new_n28447_ & ~new_n28454_;
  assign new_n28456_ = ~pi0781 & ~new_n28455_;
  assign new_n28457_ = ~new_n17873_ & new_n28455_;
  assign new_n28458_ = pi1154 & ~new_n28457_;
  assign new_n28459_ = ~new_n17876_ & new_n28455_;
  assign new_n28460_ = ~pi1154 & ~new_n28459_;
  assign new_n28461_ = ~new_n28458_ & ~new_n28460_;
  assign new_n28462_ = pi0781 & ~new_n28461_;
  assign new_n28463_ = ~new_n28456_ & ~new_n28462_;
  assign new_n28464_ = ~pi0789 & ~new_n28463_;
  assign new_n28465_ = ~new_n23057_ & new_n28463_;
  assign new_n28466_ = pi1159 & ~new_n28465_;
  assign new_n28467_ = ~new_n23060_ & new_n28463_;
  assign new_n28468_ = ~pi1159 & ~new_n28467_;
  assign new_n28469_ = ~new_n28466_ & ~new_n28468_;
  assign new_n28470_ = pi0789 & ~new_n28469_;
  assign new_n28471_ = ~new_n28464_ & ~new_n28470_;
  assign new_n28472_ = ~new_n17968_ & new_n28471_;
  assign new_n28473_ = new_n17968_ & new_n28443_;
  assign new_n28474_ = ~new_n28472_ & ~new_n28473_;
  assign new_n28475_ = ~new_n17762_ & ~new_n28474_;
  assign new_n28476_ = new_n17762_ & new_n28443_;
  assign new_n28477_ = ~new_n28475_ & ~new_n28476_;
  assign new_n28478_ = ~new_n20556_ & new_n28477_;
  assign new_n28479_ = ~pi0701 & new_n16915_;
  assign new_n28480_ = ~new_n28443_ & ~new_n28479_;
  assign new_n28481_ = ~pi0778 & ~new_n28480_;
  assign new_n28482_ = ~pi0625 & new_n28479_;
  assign new_n28483_ = ~new_n28480_ & ~new_n28482_;
  assign new_n28484_ = pi1153 & ~new_n28483_;
  assign new_n28485_ = ~pi1153 & ~new_n28443_;
  assign new_n28486_ = ~new_n28482_ & new_n28485_;
  assign new_n28487_ = pi0778 & ~new_n28486_;
  assign new_n28488_ = ~new_n28484_ & new_n28487_;
  assign new_n28489_ = ~new_n28481_ & ~new_n28488_;
  assign new_n28490_ = ~new_n17844_ & ~new_n28489_;
  assign new_n28491_ = ~new_n17846_ & new_n28490_;
  assign new_n28492_ = ~new_n17848_ & new_n28491_;
  assign new_n28493_ = ~new_n17980_ & new_n28492_;
  assign new_n28494_ = ~new_n18011_ & new_n28493_;
  assign new_n28495_ = ~pi0647 & new_n28494_;
  assign new_n28496_ = pi0647 & new_n28443_;
  assign new_n28497_ = ~pi1157 & ~new_n28496_;
  assign new_n28498_ = ~new_n28495_ & new_n28497_;
  assign new_n28499_ = pi0630 & new_n28498_;
  assign new_n28500_ = pi0647 & ~new_n28494_;
  assign new_n28501_ = ~pi0647 & ~new_n28443_;
  assign new_n28502_ = ~new_n28500_ & ~new_n28501_;
  assign new_n28503_ = new_n17801_ & ~new_n28502_;
  assign new_n28504_ = ~new_n28499_ & ~new_n28503_;
  assign new_n28505_ = ~new_n28478_ & new_n28504_;
  assign new_n28506_ = pi0787 & ~new_n28505_;
  assign new_n28507_ = pi0626 & ~new_n28471_;
  assign new_n28508_ = ~pi0626 & ~new_n28443_;
  assign new_n28509_ = new_n17731_ & ~new_n28508_;
  assign new_n28510_ = ~new_n28507_ & new_n28509_;
  assign new_n28511_ = new_n17856_ & new_n28492_;
  assign new_n28512_ = ~pi0626 & ~new_n28471_;
  assign new_n28513_ = pi0626 & ~new_n28443_;
  assign new_n28514_ = new_n17732_ & ~new_n28513_;
  assign new_n28515_ = ~new_n28512_ & new_n28514_;
  assign new_n28516_ = ~new_n28511_ & ~new_n28515_;
  assign new_n28517_ = ~new_n28510_ & new_n28516_;
  assign new_n28518_ = pi0788 & ~new_n28517_;
  assign new_n28519_ = ~new_n16639_ & ~new_n28480_;
  assign new_n28520_ = pi0625 & new_n28519_;
  assign new_n28521_ = new_n28445_ & ~new_n28519_;
  assign new_n28522_ = ~new_n28520_ & ~new_n28521_;
  assign new_n28523_ = new_n28485_ & ~new_n28522_;
  assign new_n28524_ = ~pi0608 & ~new_n28484_;
  assign new_n28525_ = ~new_n28523_ & new_n28524_;
  assign new_n28526_ = pi1153 & new_n28445_;
  assign new_n28527_ = ~new_n28520_ & new_n28526_;
  assign new_n28528_ = pi0608 & ~new_n28486_;
  assign new_n28529_ = ~new_n28527_ & new_n28528_;
  assign new_n28530_ = ~new_n28525_ & ~new_n28529_;
  assign new_n28531_ = pi0778 & ~new_n28530_;
  assign new_n28532_ = ~pi0778 & ~new_n28521_;
  assign new_n28533_ = ~new_n28531_ & ~new_n28532_;
  assign new_n28534_ = ~pi0609 & ~new_n28533_;
  assign new_n28535_ = pi0609 & ~new_n28489_;
  assign new_n28536_ = ~pi1155 & ~new_n28535_;
  assign new_n28537_ = ~new_n28534_ & new_n28536_;
  assign new_n28538_ = ~pi0660 & ~new_n28450_;
  assign new_n28539_ = ~new_n28537_ & new_n28538_;
  assign new_n28540_ = pi0609 & ~new_n28533_;
  assign new_n28541_ = ~pi0609 & ~new_n28489_;
  assign new_n28542_ = pi1155 & ~new_n28541_;
  assign new_n28543_ = ~new_n28540_ & new_n28542_;
  assign new_n28544_ = pi0660 & ~new_n28452_;
  assign new_n28545_ = ~new_n28543_ & new_n28544_;
  assign new_n28546_ = ~new_n28539_ & ~new_n28545_;
  assign new_n28547_ = pi0785 & ~new_n28546_;
  assign new_n28548_ = ~pi0785 & ~new_n28533_;
  assign new_n28549_ = ~new_n28547_ & ~new_n28548_;
  assign new_n28550_ = ~pi0618 & ~new_n28549_;
  assign new_n28551_ = pi0618 & new_n28490_;
  assign new_n28552_ = ~pi1154 & ~new_n28551_;
  assign new_n28553_ = ~new_n28550_ & new_n28552_;
  assign new_n28554_ = ~pi0627 & ~new_n28458_;
  assign new_n28555_ = ~new_n28553_ & new_n28554_;
  assign new_n28556_ = pi0618 & ~new_n28549_;
  assign new_n28557_ = ~pi0618 & new_n28490_;
  assign new_n28558_ = pi1154 & ~new_n28557_;
  assign new_n28559_ = ~new_n28556_ & new_n28558_;
  assign new_n28560_ = pi0627 & ~new_n28460_;
  assign new_n28561_ = ~new_n28559_ & new_n28560_;
  assign new_n28562_ = ~new_n28555_ & ~new_n28561_;
  assign new_n28563_ = pi0781 & ~new_n28562_;
  assign new_n28564_ = ~pi0781 & ~new_n28549_;
  assign new_n28565_ = ~new_n28563_ & ~new_n28564_;
  assign new_n28566_ = pi0619 & ~new_n28565_;
  assign new_n28567_ = ~pi0619 & new_n28491_;
  assign new_n28568_ = pi1159 & ~new_n28567_;
  assign new_n28569_ = ~new_n28566_ & new_n28568_;
  assign new_n28570_ = pi0648 & ~new_n28468_;
  assign new_n28571_ = ~new_n28569_ & new_n28570_;
  assign new_n28572_ = ~pi0619 & ~new_n28565_;
  assign new_n28573_ = pi0619 & new_n28491_;
  assign new_n28574_ = ~pi1159 & ~new_n28573_;
  assign new_n28575_ = ~new_n28572_ & new_n28574_;
  assign new_n28576_ = ~pi0648 & ~new_n28466_;
  assign new_n28577_ = ~new_n28575_ & new_n28576_;
  assign new_n28578_ = pi0789 & ~new_n28577_;
  assign new_n28579_ = ~new_n28571_ & new_n28578_;
  assign new_n28580_ = ~pi0789 & new_n28565_;
  assign new_n28581_ = new_n17969_ & ~new_n28580_;
  assign new_n28582_ = ~new_n28579_ & new_n28581_;
  assign new_n28583_ = ~new_n28518_ & ~new_n28582_;
  assign new_n28584_ = ~new_n20364_ & ~new_n28583_;
  assign new_n28585_ = new_n18008_ & ~new_n28474_;
  assign new_n28586_ = new_n20851_ & new_n28493_;
  assign new_n28587_ = ~new_n28585_ & ~new_n28586_;
  assign new_n28588_ = ~pi0629 & ~new_n28587_;
  assign new_n28589_ = new_n20855_ & new_n28493_;
  assign new_n28590_ = new_n18007_ & ~new_n28474_;
  assign new_n28591_ = ~new_n28589_ & ~new_n28590_;
  assign new_n28592_ = pi0629 & ~new_n28591_;
  assign new_n28593_ = ~new_n28588_ & ~new_n28592_;
  assign new_n28594_ = pi0792 & ~new_n28593_;
  assign new_n28595_ = ~new_n20360_ & ~new_n28594_;
  assign new_n28596_ = ~new_n28584_ & new_n28595_;
  assign new_n28597_ = ~new_n28506_ & ~new_n28596_;
  assign new_n28598_ = pi0644 & new_n28597_;
  assign new_n28599_ = ~pi0787 & ~new_n28494_;
  assign new_n28600_ = pi1157 & ~new_n28502_;
  assign new_n28601_ = ~new_n28498_ & ~new_n28600_;
  assign new_n28602_ = pi0787 & ~new_n28601_;
  assign new_n28603_ = ~new_n28599_ & ~new_n28602_;
  assign new_n28604_ = ~pi0644 & new_n28603_;
  assign new_n28605_ = pi0715 & ~new_n28604_;
  assign new_n28606_ = ~new_n28598_ & new_n28605_;
  assign new_n28607_ = ~new_n17804_ & ~new_n28477_;
  assign new_n28608_ = new_n17804_ & new_n28443_;
  assign new_n28609_ = ~new_n28607_ & ~new_n28608_;
  assign new_n28610_ = pi0644 & ~new_n28609_;
  assign new_n28611_ = ~pi0644 & new_n28443_;
  assign new_n28612_ = ~pi0715 & ~new_n28611_;
  assign new_n28613_ = ~new_n28610_ & new_n28612_;
  assign new_n28614_ = pi1160 & ~new_n28613_;
  assign new_n28615_ = ~new_n28606_ & new_n28614_;
  assign new_n28616_ = ~pi0644 & new_n28597_;
  assign new_n28617_ = pi0644 & new_n28603_;
  assign new_n28618_ = ~pi0715 & ~new_n28617_;
  assign new_n28619_ = ~new_n28616_ & new_n28618_;
  assign new_n28620_ = ~pi0644 & ~new_n28609_;
  assign new_n28621_ = pi0644 & new_n28443_;
  assign new_n28622_ = pi0715 & ~new_n28621_;
  assign new_n28623_ = ~new_n28620_ & new_n28622_;
  assign new_n28624_ = ~pi1160 & ~new_n28623_;
  assign new_n28625_ = ~new_n28619_ & new_n28624_;
  assign new_n28626_ = ~new_n28615_ & ~new_n28625_;
  assign new_n28627_ = pi0790 & ~new_n28626_;
  assign new_n28628_ = ~pi0790 & new_n28597_;
  assign new_n28629_ = pi0832 & ~new_n28628_;
  assign new_n28630_ = ~new_n28627_ & new_n28629_;
  assign new_n28631_ = ~pi0185 & ~new_n17558_;
  assign new_n28632_ = new_n17691_ & ~new_n28631_;
  assign new_n28633_ = ~pi0701 & new_n3272_;
  assign new_n28634_ = new_n28631_ & ~new_n28633_;
  assign new_n28635_ = pi0185 & ~new_n18128_;
  assign new_n28636_ = ~pi0038 & ~new_n28635_;
  assign new_n28637_ = new_n3272_ & ~new_n28636_;
  assign new_n28638_ = ~pi0185 & new_n18124_;
  assign new_n28639_ = ~new_n28637_ & ~new_n28638_;
  assign new_n28640_ = ~pi0185 & ~new_n17431_;
  assign new_n28641_ = new_n17544_ & ~new_n28640_;
  assign new_n28642_ = ~pi0701 & ~new_n28641_;
  assign new_n28643_ = ~new_n28639_ & new_n28642_;
  assign new_n28644_ = ~new_n28634_ & ~new_n28643_;
  assign new_n28645_ = ~pi0778 & new_n28644_;
  assign new_n28646_ = pi0625 & ~new_n28644_;
  assign new_n28647_ = ~pi0625 & new_n28631_;
  assign new_n28648_ = pi1153 & ~new_n28647_;
  assign new_n28649_ = ~new_n28646_ & new_n28648_;
  assign new_n28650_ = ~pi0625 & ~new_n28644_;
  assign new_n28651_ = pi0625 & new_n28631_;
  assign new_n28652_ = ~pi1153 & ~new_n28651_;
  assign new_n28653_ = ~new_n28650_ & new_n28652_;
  assign new_n28654_ = ~new_n28649_ & ~new_n28653_;
  assign new_n28655_ = pi0778 & ~new_n28654_;
  assign new_n28656_ = ~new_n28645_ & ~new_n28655_;
  assign new_n28657_ = ~new_n17618_ & ~new_n28656_;
  assign new_n28658_ = new_n17618_ & ~new_n28631_;
  assign new_n28659_ = ~new_n28657_ & ~new_n28658_;
  assign new_n28660_ = ~new_n17655_ & new_n28659_;
  assign new_n28661_ = new_n17655_ & new_n28631_;
  assign new_n28662_ = ~new_n28660_ & ~new_n28661_;
  assign new_n28663_ = ~new_n17691_ & new_n28662_;
  assign new_n28664_ = ~new_n28632_ & ~new_n28663_;
  assign new_n28665_ = ~new_n17734_ & new_n28664_;
  assign new_n28666_ = new_n17734_ & new_n28631_;
  assign new_n28667_ = ~new_n28665_ & ~new_n28666_;
  assign new_n28668_ = ~pi0792 & new_n28667_;
  assign new_n28669_ = pi0628 & ~new_n28667_;
  assign new_n28670_ = ~pi0628 & new_n28631_;
  assign new_n28671_ = pi1156 & ~new_n28670_;
  assign new_n28672_ = ~new_n28669_ & new_n28671_;
  assign new_n28673_ = ~pi0628 & ~new_n28667_;
  assign new_n28674_ = pi0628 & new_n28631_;
  assign new_n28675_ = ~pi1156 & ~new_n28674_;
  assign new_n28676_ = ~new_n28673_ & new_n28675_;
  assign new_n28677_ = ~new_n28672_ & ~new_n28676_;
  assign new_n28678_ = pi0792 & ~new_n28677_;
  assign new_n28679_ = ~new_n28668_ & ~new_n28678_;
  assign new_n28680_ = ~pi0647 & ~new_n28679_;
  assign new_n28681_ = pi0647 & ~new_n28631_;
  assign new_n28682_ = ~new_n28680_ & ~new_n28681_;
  assign new_n28683_ = ~pi1157 & new_n28682_;
  assign new_n28684_ = pi0647 & ~new_n28679_;
  assign new_n28685_ = ~pi0647 & ~new_n28631_;
  assign new_n28686_ = ~new_n28684_ & ~new_n28685_;
  assign new_n28687_ = pi1157 & new_n28686_;
  assign new_n28688_ = ~new_n28683_ & ~new_n28687_;
  assign new_n28689_ = pi0787 & ~new_n28688_;
  assign new_n28690_ = ~pi0787 & new_n28679_;
  assign new_n28691_ = ~new_n28689_ & ~new_n28690_;
  assign new_n28692_ = ~pi0644 & ~new_n28691_;
  assign new_n28693_ = pi0715 & ~new_n28692_;
  assign new_n28694_ = pi0185 & ~new_n3272_;
  assign new_n28695_ = pi0751 & new_n17347_;
  assign new_n28696_ = pi0185 & new_n17424_;
  assign new_n28697_ = ~new_n28695_ & ~new_n28696_;
  assign new_n28698_ = pi0039 & ~new_n28697_;
  assign new_n28699_ = ~pi0185 & ~pi0751;
  assign new_n28700_ = new_n17393_ & new_n28699_;
  assign new_n28701_ = pi0185 & pi0751;
  assign new_n28702_ = pi0185 & ~new_n17215_;
  assign new_n28703_ = ~new_n21261_ & ~new_n28702_;
  assign new_n28704_ = ~pi0039 & ~new_n28703_;
  assign new_n28705_ = ~new_n28701_ & ~new_n28704_;
  assign new_n28706_ = ~new_n28700_ & new_n28705_;
  assign new_n28707_ = ~new_n28698_ & new_n28706_;
  assign new_n28708_ = ~pi0038 & ~new_n28707_;
  assign new_n28709_ = ~pi0751 & new_n17433_;
  assign new_n28710_ = pi0038 & ~new_n28640_;
  assign new_n28711_ = ~new_n28709_ & new_n28710_;
  assign new_n28712_ = ~new_n28708_ & ~new_n28711_;
  assign new_n28713_ = new_n3272_ & ~new_n28712_;
  assign new_n28714_ = ~new_n28694_ & ~new_n28713_;
  assign new_n28715_ = ~new_n17590_ & ~new_n28714_;
  assign new_n28716_ = new_n17590_ & ~new_n28631_;
  assign new_n28717_ = ~new_n28715_ & ~new_n28716_;
  assign new_n28718_ = ~pi0785 & ~new_n28717_;
  assign new_n28719_ = ~new_n17591_ & ~new_n28631_;
  assign new_n28720_ = pi0609 & new_n28715_;
  assign new_n28721_ = ~new_n28719_ & ~new_n28720_;
  assign new_n28722_ = pi1155 & ~new_n28721_;
  assign new_n28723_ = ~new_n17603_ & ~new_n28631_;
  assign new_n28724_ = ~pi0609 & new_n28715_;
  assign new_n28725_ = ~new_n28723_ & ~new_n28724_;
  assign new_n28726_ = ~pi1155 & ~new_n28725_;
  assign new_n28727_ = ~new_n28722_ & ~new_n28726_;
  assign new_n28728_ = pi0785 & ~new_n28727_;
  assign new_n28729_ = ~new_n28718_ & ~new_n28728_;
  assign new_n28730_ = ~pi0781 & ~new_n28729_;
  assign new_n28731_ = pi0618 & new_n28729_;
  assign new_n28732_ = ~pi0618 & new_n28631_;
  assign new_n28733_ = pi1154 & ~new_n28732_;
  assign new_n28734_ = ~new_n28731_ & new_n28733_;
  assign new_n28735_ = ~pi0618 & new_n28729_;
  assign new_n28736_ = pi0618 & new_n28631_;
  assign new_n28737_ = ~pi1154 & ~new_n28736_;
  assign new_n28738_ = ~new_n28735_ & new_n28737_;
  assign new_n28739_ = ~new_n28734_ & ~new_n28738_;
  assign new_n28740_ = pi0781 & ~new_n28739_;
  assign new_n28741_ = ~new_n28730_ & ~new_n28740_;
  assign new_n28742_ = ~pi0789 & ~new_n28741_;
  assign new_n28743_ = pi0619 & new_n28741_;
  assign new_n28744_ = ~pi0619 & new_n28631_;
  assign new_n28745_ = pi1159 & ~new_n28744_;
  assign new_n28746_ = ~new_n28743_ & new_n28745_;
  assign new_n28747_ = ~pi0619 & new_n28741_;
  assign new_n28748_ = pi0619 & new_n28631_;
  assign new_n28749_ = ~pi1159 & ~new_n28748_;
  assign new_n28750_ = ~new_n28747_ & new_n28749_;
  assign new_n28751_ = ~new_n28746_ & ~new_n28750_;
  assign new_n28752_ = pi0789 & ~new_n28751_;
  assign new_n28753_ = ~new_n28742_ & ~new_n28752_;
  assign new_n28754_ = ~new_n17968_ & new_n28753_;
  assign new_n28755_ = new_n17968_ & new_n28631_;
  assign new_n28756_ = ~new_n28754_ & ~new_n28755_;
  assign new_n28757_ = ~new_n17762_ & ~new_n28756_;
  assign new_n28758_ = new_n17762_ & new_n28631_;
  assign new_n28759_ = ~new_n28757_ & ~new_n28758_;
  assign new_n28760_ = ~new_n17804_ & ~new_n28759_;
  assign new_n28761_ = new_n17804_ & new_n28631_;
  assign new_n28762_ = ~new_n28760_ & ~new_n28761_;
  assign new_n28763_ = pi0644 & ~new_n28762_;
  assign new_n28764_ = ~pi0644 & new_n28631_;
  assign new_n28765_ = ~pi0715 & ~new_n28764_;
  assign new_n28766_ = ~new_n28763_ & new_n28765_;
  assign new_n28767_ = pi1160 & ~new_n28766_;
  assign new_n28768_ = ~new_n28693_ & new_n28767_;
  assign new_n28769_ = pi0644 & ~new_n28691_;
  assign new_n28770_ = ~pi0715 & ~new_n28769_;
  assign new_n28771_ = ~pi0644 & ~new_n28762_;
  assign new_n28772_ = pi0644 & new_n28631_;
  assign new_n28773_ = pi0715 & ~new_n28772_;
  assign new_n28774_ = ~new_n28771_ & new_n28773_;
  assign new_n28775_ = ~pi1160 & ~new_n28774_;
  assign new_n28776_ = ~new_n28770_ & new_n28775_;
  assign new_n28777_ = ~new_n28768_ & ~new_n28776_;
  assign new_n28778_ = pi0790 & ~new_n28777_;
  assign new_n28779_ = pi0644 & new_n28767_;
  assign new_n28780_ = ~pi0644 & new_n28775_;
  assign new_n28781_ = pi0790 & ~new_n28780_;
  assign new_n28782_ = ~new_n28779_ & new_n28781_;
  assign new_n28783_ = ~new_n20567_ & new_n28756_;
  assign new_n28784_ = ~pi0629 & new_n28672_;
  assign new_n28785_ = pi0629 & new_n28676_;
  assign new_n28786_ = ~new_n28784_ & ~new_n28785_;
  assign new_n28787_ = ~new_n28783_ & new_n28786_;
  assign new_n28788_ = pi0792 & ~new_n28787_;
  assign new_n28789_ = pi0701 & new_n28712_;
  assign new_n28790_ = ~pi0185 & new_n16810_;
  assign new_n28791_ = pi0185 & new_n16928_;
  assign new_n28792_ = pi0751 & ~new_n28791_;
  assign new_n28793_ = ~new_n28790_ & new_n28792_;
  assign new_n28794_ = pi0185 & new_n17007_;
  assign new_n28795_ = ~pi0185 & ~new_n17074_;
  assign new_n28796_ = ~pi0751 & ~new_n28795_;
  assign new_n28797_ = ~new_n28794_ & new_n28796_;
  assign new_n28798_ = pi0039 & ~new_n28797_;
  assign new_n28799_ = ~new_n28793_ & new_n28798_;
  assign new_n28800_ = ~pi0185 & ~new_n17217_;
  assign new_n28801_ = pi0185 & ~new_n17178_;
  assign new_n28802_ = pi0751 & ~new_n28801_;
  assign new_n28803_ = ~new_n28800_ & new_n28802_;
  assign new_n28804_ = ~pi0185 & new_n17227_;
  assign new_n28805_ = pi0185 & new_n17234_;
  assign new_n28806_ = ~pi0751 & ~new_n28805_;
  assign new_n28807_ = ~new_n28804_ & new_n28806_;
  assign new_n28808_ = ~new_n28803_ & ~new_n28807_;
  assign new_n28809_ = ~pi0039 & ~new_n28808_;
  assign new_n28810_ = ~pi0038 & ~new_n28809_;
  assign new_n28811_ = ~new_n28799_ & new_n28810_;
  assign new_n28812_ = ~pi0751 & ~new_n17035_;
  assign new_n28813_ = new_n19383_ & ~new_n28812_;
  assign new_n28814_ = ~pi0185 & ~new_n28813_;
  assign new_n28815_ = ~new_n16916_ & ~new_n28444_;
  assign new_n28816_ = pi0185 & ~new_n28815_;
  assign new_n28817_ = new_n6257_ & new_n28816_;
  assign new_n28818_ = pi0038 & ~new_n28817_;
  assign new_n28819_ = ~new_n28814_ & new_n28818_;
  assign new_n28820_ = ~pi0701 & ~new_n28819_;
  assign new_n28821_ = ~new_n28811_ & new_n28820_;
  assign new_n28822_ = new_n3272_ & ~new_n28821_;
  assign new_n28823_ = ~new_n28789_ & new_n28822_;
  assign new_n28824_ = ~new_n28694_ & ~new_n28823_;
  assign new_n28825_ = ~pi0625 & new_n28824_;
  assign new_n28826_ = pi0625 & new_n28714_;
  assign new_n28827_ = ~pi1153 & ~new_n28826_;
  assign new_n28828_ = ~new_n28825_ & new_n28827_;
  assign new_n28829_ = ~pi0608 & ~new_n28649_;
  assign new_n28830_ = ~new_n28828_ & new_n28829_;
  assign new_n28831_ = pi0625 & new_n28824_;
  assign new_n28832_ = ~pi0625 & new_n28714_;
  assign new_n28833_ = pi1153 & ~new_n28832_;
  assign new_n28834_ = ~new_n28831_ & new_n28833_;
  assign new_n28835_ = pi0608 & ~new_n28653_;
  assign new_n28836_ = ~new_n28834_ & new_n28835_;
  assign new_n28837_ = ~new_n28830_ & ~new_n28836_;
  assign new_n28838_ = pi0778 & ~new_n28837_;
  assign new_n28839_ = ~pi0778 & new_n28824_;
  assign new_n28840_ = ~new_n28838_ & ~new_n28839_;
  assign new_n28841_ = ~pi0609 & ~new_n28840_;
  assign new_n28842_ = pi0609 & new_n28656_;
  assign new_n28843_ = ~pi1155 & ~new_n28842_;
  assign new_n28844_ = ~new_n28841_ & new_n28843_;
  assign new_n28845_ = ~pi0660 & ~new_n28722_;
  assign new_n28846_ = ~new_n28844_ & new_n28845_;
  assign new_n28847_ = pi0609 & ~new_n28840_;
  assign new_n28848_ = ~pi0609 & new_n28656_;
  assign new_n28849_ = pi1155 & ~new_n28848_;
  assign new_n28850_ = ~new_n28847_ & new_n28849_;
  assign new_n28851_ = pi0660 & ~new_n28726_;
  assign new_n28852_ = ~new_n28850_ & new_n28851_;
  assign new_n28853_ = ~new_n28846_ & ~new_n28852_;
  assign new_n28854_ = pi0785 & ~new_n28853_;
  assign new_n28855_ = ~pi0785 & ~new_n28840_;
  assign new_n28856_ = ~new_n28854_ & ~new_n28855_;
  assign new_n28857_ = ~pi0618 & ~new_n28856_;
  assign new_n28858_ = pi0618 & new_n28659_;
  assign new_n28859_ = ~pi1154 & ~new_n28858_;
  assign new_n28860_ = ~new_n28857_ & new_n28859_;
  assign new_n28861_ = ~pi0627 & ~new_n28734_;
  assign new_n28862_ = ~new_n28860_ & new_n28861_;
  assign new_n28863_ = pi0618 & ~new_n28856_;
  assign new_n28864_ = ~pi0618 & new_n28659_;
  assign new_n28865_ = pi1154 & ~new_n28864_;
  assign new_n28866_ = ~new_n28863_ & new_n28865_;
  assign new_n28867_ = pi0627 & ~new_n28738_;
  assign new_n28868_ = ~new_n28866_ & new_n28867_;
  assign new_n28869_ = ~new_n28862_ & ~new_n28868_;
  assign new_n28870_ = pi0781 & ~new_n28869_;
  assign new_n28871_ = ~pi0781 & ~new_n28856_;
  assign new_n28872_ = ~new_n28870_ & ~new_n28871_;
  assign new_n28873_ = pi0619 & ~new_n28872_;
  assign new_n28874_ = ~pi0619 & ~new_n28662_;
  assign new_n28875_ = pi1159 & ~new_n28874_;
  assign new_n28876_ = ~new_n28873_ & new_n28875_;
  assign new_n28877_ = pi0648 & ~new_n28750_;
  assign new_n28878_ = ~new_n28876_ & new_n28877_;
  assign new_n28879_ = ~pi0619 & ~new_n28872_;
  assign new_n28880_ = pi0619 & ~new_n28662_;
  assign new_n28881_ = ~pi1159 & ~new_n28880_;
  assign new_n28882_ = ~new_n28879_ & new_n28881_;
  assign new_n28883_ = ~pi0648 & ~new_n28746_;
  assign new_n28884_ = ~new_n28882_ & new_n28883_;
  assign new_n28885_ = pi0789 & ~new_n28884_;
  assign new_n28886_ = ~new_n28878_ & new_n28885_;
  assign new_n28887_ = ~pi0789 & new_n28872_;
  assign new_n28888_ = new_n17969_ & ~new_n28887_;
  assign new_n28889_ = ~new_n28886_ & new_n28888_;
  assign new_n28890_ = pi0626 & ~new_n28753_;
  assign new_n28891_ = ~pi0626 & ~new_n28631_;
  assign new_n28892_ = new_n17731_ & ~new_n28891_;
  assign new_n28893_ = ~new_n28890_ & new_n28892_;
  assign new_n28894_ = new_n17856_ & new_n28664_;
  assign new_n28895_ = ~pi0626 & ~new_n28753_;
  assign new_n28896_ = pi0626 & ~new_n28631_;
  assign new_n28897_ = new_n17732_ & ~new_n28896_;
  assign new_n28898_ = ~new_n28895_ & new_n28897_;
  assign new_n28899_ = ~new_n28894_ & ~new_n28898_;
  assign new_n28900_ = ~new_n28893_ & new_n28899_;
  assign new_n28901_ = pi0788 & ~new_n28900_;
  assign new_n28902_ = ~new_n20364_ & ~new_n28901_;
  assign new_n28903_ = ~new_n28889_ & new_n28902_;
  assign new_n28904_ = ~new_n28788_ & ~new_n28903_;
  assign new_n28905_ = ~new_n20360_ & ~new_n28904_;
  assign new_n28906_ = ~new_n20556_ & new_n28759_;
  assign new_n28907_ = new_n17802_ & ~new_n28682_;
  assign new_n28908_ = new_n17801_ & ~new_n28686_;
  assign new_n28909_ = ~new_n28907_ & ~new_n28908_;
  assign new_n28910_ = ~new_n28906_ & new_n28909_;
  assign new_n28911_ = pi0787 & ~new_n28910_;
  assign new_n28912_ = ~new_n28905_ & ~new_n28911_;
  assign new_n28913_ = ~new_n28782_ & new_n28912_;
  assign new_n28914_ = ~new_n28778_ & ~new_n28913_;
  assign new_n28915_ = ~po1038 & ~new_n28914_;
  assign new_n28916_ = ~pi0185 & po1038;
  assign new_n28917_ = ~pi0832 & ~new_n28916_;
  assign new_n28918_ = ~new_n28915_ & new_n28917_;
  assign po0342 = ~new_n28630_ & ~new_n28918_;
  assign new_n28920_ = pi0186 & ~new_n3272_;
  assign new_n28921_ = ~pi0186 & ~new_n17551_;
  assign new_n28922_ = pi0752 & ~new_n28921_;
  assign new_n28923_ = pi0186 & ~new_n19371_;
  assign new_n28924_ = ~pi0186 & ~pi0752;
  assign new_n28925_ = new_n19376_ & new_n28924_;
  assign new_n28926_ = ~new_n28923_ & ~new_n28925_;
  assign new_n28927_ = ~new_n19370_ & ~new_n28926_;
  assign new_n28928_ = ~new_n28922_ & ~new_n28927_;
  assign new_n28929_ = ~pi0703 & new_n28928_;
  assign new_n28930_ = ~pi0186 & new_n19389_;
  assign new_n28931_ = pi0186 & new_n19394_;
  assign new_n28932_ = pi0752 & ~new_n19396_;
  assign new_n28933_ = ~new_n28931_ & new_n28932_;
  assign new_n28934_ = ~new_n28930_ & new_n28933_;
  assign new_n28935_ = pi0186 & new_n19406_;
  assign new_n28936_ = ~pi0186 & ~new_n19414_;
  assign new_n28937_ = ~pi0752 & ~new_n28936_;
  assign new_n28938_ = ~new_n28935_ & new_n28937_;
  assign new_n28939_ = pi0703 & ~new_n28938_;
  assign new_n28940_ = ~new_n28934_ & new_n28939_;
  assign new_n28941_ = new_n3272_ & ~new_n28940_;
  assign new_n28942_ = ~new_n28929_ & new_n28941_;
  assign new_n28943_ = ~new_n28920_ & ~new_n28942_;
  assign new_n28944_ = ~pi0625 & new_n28943_;
  assign new_n28945_ = new_n3272_ & ~new_n28928_;
  assign new_n28946_ = ~new_n28920_ & ~new_n28945_;
  assign new_n28947_ = pi0625 & new_n28946_;
  assign new_n28948_ = ~pi1153 & ~new_n28947_;
  assign new_n28949_ = ~new_n28944_ & new_n28948_;
  assign new_n28950_ = ~pi0186 & new_n18124_;
  assign new_n28951_ = pi0186 & ~new_n18128_;
  assign new_n28952_ = ~pi0038 & ~new_n28951_;
  assign new_n28953_ = ~new_n28950_ & new_n28952_;
  assign new_n28954_ = ~pi0186 & ~new_n17431_;
  assign new_n28955_ = new_n17544_ & ~new_n28954_;
  assign new_n28956_ = pi0703 & ~new_n28955_;
  assign new_n28957_ = ~new_n28953_ & new_n28956_;
  assign new_n28958_ = ~pi0703 & new_n28921_;
  assign new_n28959_ = new_n3272_ & ~new_n28958_;
  assign new_n28960_ = ~new_n28957_ & new_n28959_;
  assign new_n28961_ = ~new_n28920_ & ~new_n28960_;
  assign new_n28962_ = pi0625 & new_n28961_;
  assign new_n28963_ = ~pi0186 & ~new_n17558_;
  assign new_n28964_ = ~pi0625 & new_n28963_;
  assign new_n28965_ = pi1153 & ~new_n28964_;
  assign new_n28966_ = ~new_n28962_ & new_n28965_;
  assign new_n28967_ = ~pi0608 & ~new_n28966_;
  assign new_n28968_ = ~new_n28949_ & new_n28967_;
  assign new_n28969_ = pi0625 & new_n28943_;
  assign new_n28970_ = ~pi0625 & new_n28946_;
  assign new_n28971_ = pi1153 & ~new_n28970_;
  assign new_n28972_ = ~new_n28969_ & new_n28971_;
  assign new_n28973_ = ~pi0625 & new_n28961_;
  assign new_n28974_ = pi0625 & new_n28963_;
  assign new_n28975_ = ~pi1153 & ~new_n28974_;
  assign new_n28976_ = ~new_n28973_ & new_n28975_;
  assign new_n28977_ = pi0608 & ~new_n28976_;
  assign new_n28978_ = ~new_n28972_ & new_n28977_;
  assign new_n28979_ = ~new_n28968_ & ~new_n28978_;
  assign new_n28980_ = pi0778 & ~new_n28979_;
  assign new_n28981_ = ~pi0778 & new_n28943_;
  assign new_n28982_ = ~new_n28980_ & ~new_n28981_;
  assign new_n28983_ = ~pi0609 & ~new_n28982_;
  assign new_n28984_ = ~pi0778 & ~new_n28961_;
  assign new_n28985_ = ~new_n28966_ & ~new_n28976_;
  assign new_n28986_ = pi0778 & ~new_n28985_;
  assign new_n28987_ = ~new_n28984_ & ~new_n28986_;
  assign new_n28988_ = pi0609 & new_n28987_;
  assign new_n28989_ = ~pi1155 & ~new_n28988_;
  assign new_n28990_ = ~new_n28983_ & new_n28989_;
  assign new_n28991_ = ~new_n17591_ & ~new_n28963_;
  assign new_n28992_ = ~new_n17590_ & ~new_n28946_;
  assign new_n28993_ = pi0609 & new_n28992_;
  assign new_n28994_ = ~new_n28991_ & ~new_n28993_;
  assign new_n28995_ = pi1155 & ~new_n28994_;
  assign new_n28996_ = ~pi0660 & ~new_n28995_;
  assign new_n28997_ = ~new_n28990_ & new_n28996_;
  assign new_n28998_ = pi0609 & ~new_n28982_;
  assign new_n28999_ = ~pi0609 & new_n28987_;
  assign new_n29000_ = pi1155 & ~new_n28999_;
  assign new_n29001_ = ~new_n28998_ & new_n29000_;
  assign new_n29002_ = ~new_n17603_ & ~new_n28963_;
  assign new_n29003_ = ~pi0609 & new_n28992_;
  assign new_n29004_ = ~new_n29002_ & ~new_n29003_;
  assign new_n29005_ = ~pi1155 & ~new_n29004_;
  assign new_n29006_ = pi0660 & ~new_n29005_;
  assign new_n29007_ = ~new_n29001_ & new_n29006_;
  assign new_n29008_ = ~new_n28997_ & ~new_n29007_;
  assign new_n29009_ = pi0785 & ~new_n29008_;
  assign new_n29010_ = ~pi0785 & ~new_n28982_;
  assign new_n29011_ = ~new_n29009_ & ~new_n29010_;
  assign new_n29012_ = ~pi0618 & ~new_n29011_;
  assign new_n29013_ = ~new_n17618_ & ~new_n28987_;
  assign new_n29014_ = new_n17618_ & ~new_n28963_;
  assign new_n29015_ = ~new_n29013_ & ~new_n29014_;
  assign new_n29016_ = pi0618 & new_n29015_;
  assign new_n29017_ = ~pi1154 & ~new_n29016_;
  assign new_n29018_ = ~new_n29012_ & new_n29017_;
  assign new_n29019_ = new_n17590_ & ~new_n28963_;
  assign new_n29020_ = ~new_n28992_ & ~new_n29019_;
  assign new_n29021_ = ~pi0785 & ~new_n29020_;
  assign new_n29022_ = ~new_n28995_ & ~new_n29005_;
  assign new_n29023_ = pi0785 & ~new_n29022_;
  assign new_n29024_ = ~new_n29021_ & ~new_n29023_;
  assign new_n29025_ = pi0618 & new_n29024_;
  assign new_n29026_ = ~pi0618 & new_n28963_;
  assign new_n29027_ = pi1154 & ~new_n29026_;
  assign new_n29028_ = ~new_n29025_ & new_n29027_;
  assign new_n29029_ = ~pi0627 & ~new_n29028_;
  assign new_n29030_ = ~new_n29018_ & new_n29029_;
  assign new_n29031_ = pi0618 & ~new_n29011_;
  assign new_n29032_ = ~pi0618 & new_n29015_;
  assign new_n29033_ = pi1154 & ~new_n29032_;
  assign new_n29034_ = ~new_n29031_ & new_n29033_;
  assign new_n29035_ = ~pi0618 & new_n29024_;
  assign new_n29036_ = pi0618 & new_n28963_;
  assign new_n29037_ = ~pi1154 & ~new_n29036_;
  assign new_n29038_ = ~new_n29035_ & new_n29037_;
  assign new_n29039_ = pi0627 & ~new_n29038_;
  assign new_n29040_ = ~new_n29034_ & new_n29039_;
  assign new_n29041_ = ~new_n29030_ & ~new_n29040_;
  assign new_n29042_ = pi0781 & ~new_n29041_;
  assign new_n29043_ = ~pi0781 & ~new_n29011_;
  assign new_n29044_ = ~new_n29042_ & ~new_n29043_;
  assign new_n29045_ = ~pi0619 & ~new_n29044_;
  assign new_n29046_ = ~new_n17655_ & new_n29015_;
  assign new_n29047_ = new_n17655_ & new_n28963_;
  assign new_n29048_ = ~new_n29046_ & ~new_n29047_;
  assign new_n29049_ = pi0619 & ~new_n29048_;
  assign new_n29050_ = ~pi1159 & ~new_n29049_;
  assign new_n29051_ = ~new_n29045_ & new_n29050_;
  assign new_n29052_ = ~pi0781 & ~new_n29024_;
  assign new_n29053_ = ~new_n29028_ & ~new_n29038_;
  assign new_n29054_ = pi0781 & ~new_n29053_;
  assign new_n29055_ = ~new_n29052_ & ~new_n29054_;
  assign new_n29056_ = pi0619 & new_n29055_;
  assign new_n29057_ = ~pi0619 & new_n28963_;
  assign new_n29058_ = pi1159 & ~new_n29057_;
  assign new_n29059_ = ~new_n29056_ & new_n29058_;
  assign new_n29060_ = ~pi0648 & ~new_n29059_;
  assign new_n29061_ = ~new_n29051_ & new_n29060_;
  assign new_n29062_ = pi0619 & ~new_n29044_;
  assign new_n29063_ = ~pi0619 & ~new_n29048_;
  assign new_n29064_ = pi1159 & ~new_n29063_;
  assign new_n29065_ = ~new_n29062_ & new_n29064_;
  assign new_n29066_ = ~pi0619 & new_n29055_;
  assign new_n29067_ = pi0619 & new_n28963_;
  assign new_n29068_ = ~pi1159 & ~new_n29067_;
  assign new_n29069_ = ~new_n29066_ & new_n29068_;
  assign new_n29070_ = pi0648 & ~new_n29069_;
  assign new_n29071_ = ~new_n29065_ & new_n29070_;
  assign new_n29072_ = ~new_n29061_ & ~new_n29071_;
  assign new_n29073_ = pi0789 & ~new_n29072_;
  assign new_n29074_ = ~pi0789 & ~new_n29044_;
  assign new_n29075_ = ~new_n29073_ & ~new_n29074_;
  assign new_n29076_ = ~pi0788 & new_n29075_;
  assign new_n29077_ = ~pi0626 & new_n29075_;
  assign new_n29078_ = new_n17691_ & ~new_n28963_;
  assign new_n29079_ = ~new_n17691_ & new_n29048_;
  assign new_n29080_ = ~new_n29078_ & ~new_n29079_;
  assign new_n29081_ = pi0626 & ~new_n29080_;
  assign new_n29082_ = ~pi0641 & ~new_n29081_;
  assign new_n29083_ = ~new_n29077_ & new_n29082_;
  assign new_n29084_ = ~pi0789 & ~new_n29055_;
  assign new_n29085_ = ~new_n29059_ & ~new_n29069_;
  assign new_n29086_ = pi0789 & ~new_n29085_;
  assign new_n29087_ = ~new_n29084_ & ~new_n29086_;
  assign new_n29088_ = ~pi0626 & ~new_n29087_;
  assign new_n29089_ = pi0626 & ~new_n28963_;
  assign new_n29090_ = pi0641 & ~new_n29089_;
  assign new_n29091_ = ~new_n29088_ & new_n29090_;
  assign new_n29092_ = ~pi1158 & ~new_n29091_;
  assign new_n29093_ = ~new_n29083_ & new_n29092_;
  assign new_n29094_ = pi0626 & new_n29075_;
  assign new_n29095_ = ~pi0626 & ~new_n29080_;
  assign new_n29096_ = pi0641 & ~new_n29095_;
  assign new_n29097_ = ~new_n29094_ & new_n29096_;
  assign new_n29098_ = pi0626 & ~new_n29087_;
  assign new_n29099_ = ~pi0626 & ~new_n28963_;
  assign new_n29100_ = ~pi0641 & ~new_n29099_;
  assign new_n29101_ = ~new_n29098_ & new_n29100_;
  assign new_n29102_ = pi1158 & ~new_n29101_;
  assign new_n29103_ = ~new_n29097_ & new_n29102_;
  assign new_n29104_ = ~new_n29093_ & ~new_n29103_;
  assign new_n29105_ = pi0788 & ~new_n29104_;
  assign new_n29106_ = ~new_n29076_ & ~new_n29105_;
  assign new_n29107_ = ~pi0628 & new_n29106_;
  assign new_n29108_ = ~new_n17968_ & new_n29087_;
  assign new_n29109_ = new_n17968_ & new_n28963_;
  assign new_n29110_ = ~new_n29108_ & ~new_n29109_;
  assign new_n29111_ = pi0628 & ~new_n29110_;
  assign new_n29112_ = ~pi1156 & ~new_n29111_;
  assign new_n29113_ = ~new_n29107_ & new_n29112_;
  assign new_n29114_ = ~new_n17734_ & new_n29080_;
  assign new_n29115_ = new_n17734_ & new_n28963_;
  assign new_n29116_ = ~new_n29114_ & ~new_n29115_;
  assign new_n29117_ = pi0628 & ~new_n29116_;
  assign new_n29118_ = ~pi0628 & new_n28963_;
  assign new_n29119_ = pi1156 & ~new_n29118_;
  assign new_n29120_ = ~new_n29117_ & new_n29119_;
  assign new_n29121_ = ~pi0629 & ~new_n29120_;
  assign new_n29122_ = ~new_n29113_ & new_n29121_;
  assign new_n29123_ = pi0628 & new_n29106_;
  assign new_n29124_ = ~pi0628 & ~new_n29110_;
  assign new_n29125_ = pi1156 & ~new_n29124_;
  assign new_n29126_ = ~new_n29123_ & new_n29125_;
  assign new_n29127_ = ~pi0628 & ~new_n29116_;
  assign new_n29128_ = pi0628 & new_n28963_;
  assign new_n29129_ = ~pi1156 & ~new_n29128_;
  assign new_n29130_ = ~new_n29127_ & new_n29129_;
  assign new_n29131_ = pi0629 & ~new_n29130_;
  assign new_n29132_ = ~new_n29126_ & new_n29131_;
  assign new_n29133_ = ~new_n29122_ & ~new_n29132_;
  assign new_n29134_ = pi0792 & ~new_n29133_;
  assign new_n29135_ = ~pi0792 & new_n29106_;
  assign new_n29136_ = ~new_n29134_ & ~new_n29135_;
  assign new_n29137_ = ~pi0647 & ~new_n29136_;
  assign new_n29138_ = ~new_n17762_ & ~new_n29110_;
  assign new_n29139_ = new_n17762_ & new_n28963_;
  assign new_n29140_ = ~new_n29138_ & ~new_n29139_;
  assign new_n29141_ = pi0647 & ~new_n29140_;
  assign new_n29142_ = ~pi1157 & ~new_n29141_;
  assign new_n29143_ = ~new_n29137_ & new_n29142_;
  assign new_n29144_ = ~pi0792 & new_n29116_;
  assign new_n29145_ = ~new_n29120_ & ~new_n29130_;
  assign new_n29146_ = pi0792 & ~new_n29145_;
  assign new_n29147_ = ~new_n29144_ & ~new_n29146_;
  assign new_n29148_ = pi0647 & new_n29147_;
  assign new_n29149_ = ~pi0647 & new_n28963_;
  assign new_n29150_ = pi1157 & ~new_n29149_;
  assign new_n29151_ = ~new_n29148_ & new_n29150_;
  assign new_n29152_ = ~pi0630 & ~new_n29151_;
  assign new_n29153_ = ~new_n29143_ & new_n29152_;
  assign new_n29154_ = pi0647 & ~new_n29136_;
  assign new_n29155_ = ~pi0647 & ~new_n29140_;
  assign new_n29156_ = pi1157 & ~new_n29155_;
  assign new_n29157_ = ~new_n29154_ & new_n29156_;
  assign new_n29158_ = ~pi0647 & new_n29147_;
  assign new_n29159_ = pi0647 & new_n28963_;
  assign new_n29160_ = ~pi1157 & ~new_n29159_;
  assign new_n29161_ = ~new_n29158_ & new_n29160_;
  assign new_n29162_ = pi0630 & ~new_n29161_;
  assign new_n29163_ = ~new_n29157_ & new_n29162_;
  assign new_n29164_ = ~new_n29153_ & ~new_n29163_;
  assign new_n29165_ = pi0787 & ~new_n29164_;
  assign new_n29166_ = ~pi0787 & ~new_n29136_;
  assign new_n29167_ = ~new_n29165_ & ~new_n29166_;
  assign new_n29168_ = ~pi0644 & ~new_n29167_;
  assign new_n29169_ = ~pi0787 & ~new_n29147_;
  assign new_n29170_ = ~new_n29151_ & ~new_n29161_;
  assign new_n29171_ = pi0787 & ~new_n29170_;
  assign new_n29172_ = ~new_n29169_ & ~new_n29171_;
  assign new_n29173_ = pi0644 & new_n29172_;
  assign new_n29174_ = ~pi0715 & ~new_n29173_;
  assign new_n29175_ = ~new_n29168_ & new_n29174_;
  assign new_n29176_ = new_n17804_ & ~new_n28963_;
  assign new_n29177_ = ~new_n17804_ & new_n29140_;
  assign new_n29178_ = ~new_n29176_ & ~new_n29177_;
  assign new_n29179_ = ~pi0644 & new_n29178_;
  assign new_n29180_ = pi0644 & new_n28963_;
  assign new_n29181_ = pi0715 & ~new_n29180_;
  assign new_n29182_ = ~new_n29179_ & new_n29181_;
  assign new_n29183_ = ~pi1160 & ~new_n29182_;
  assign new_n29184_ = ~new_n29175_ & new_n29183_;
  assign new_n29185_ = pi0644 & ~new_n29167_;
  assign new_n29186_ = ~pi0644 & new_n29172_;
  assign new_n29187_ = pi0715 & ~new_n29186_;
  assign new_n29188_ = ~new_n29185_ & new_n29187_;
  assign new_n29189_ = pi0644 & new_n29178_;
  assign new_n29190_ = ~pi0644 & new_n28963_;
  assign new_n29191_ = ~pi0715 & ~new_n29190_;
  assign new_n29192_ = ~new_n29189_ & new_n29191_;
  assign new_n29193_ = pi1160 & ~new_n29192_;
  assign new_n29194_ = ~new_n29188_ & new_n29193_;
  assign new_n29195_ = pi0790 & ~new_n29194_;
  assign new_n29196_ = ~new_n29184_ & new_n29195_;
  assign new_n29197_ = ~pi0790 & new_n29167_;
  assign new_n29198_ = ~po1038 & ~new_n29197_;
  assign new_n29199_ = ~new_n29196_ & new_n29198_;
  assign new_n29200_ = ~pi0186 & po1038;
  assign new_n29201_ = ~pi0832 & ~new_n29200_;
  assign new_n29202_ = ~new_n29199_ & new_n29201_;
  assign new_n29203_ = ~pi0186 & ~new_n2754_;
  assign new_n29204_ = ~pi0752 & new_n16913_;
  assign new_n29205_ = ~new_n29203_ & ~new_n29204_;
  assign new_n29206_ = ~new_n17858_ & ~new_n29205_;
  assign new_n29207_ = ~pi0785 & ~new_n29206_;
  assign new_n29208_ = ~new_n17863_ & ~new_n29205_;
  assign new_n29209_ = pi1155 & ~new_n29208_;
  assign new_n29210_ = ~new_n17866_ & new_n29206_;
  assign new_n29211_ = ~pi1155 & ~new_n29210_;
  assign new_n29212_ = ~new_n29209_ & ~new_n29211_;
  assign new_n29213_ = pi0785 & ~new_n29212_;
  assign new_n29214_ = ~new_n29207_ & ~new_n29213_;
  assign new_n29215_ = ~pi0781 & ~new_n29214_;
  assign new_n29216_ = ~new_n17873_ & new_n29214_;
  assign new_n29217_ = pi1154 & ~new_n29216_;
  assign new_n29218_ = ~new_n17876_ & new_n29214_;
  assign new_n29219_ = ~pi1154 & ~new_n29218_;
  assign new_n29220_ = ~new_n29217_ & ~new_n29219_;
  assign new_n29221_ = pi0781 & ~new_n29220_;
  assign new_n29222_ = ~new_n29215_ & ~new_n29221_;
  assign new_n29223_ = ~pi0789 & ~new_n29222_;
  assign new_n29224_ = pi0619 & new_n29222_;
  assign new_n29225_ = ~pi0619 & new_n29203_;
  assign new_n29226_ = pi1159 & ~new_n29225_;
  assign new_n29227_ = ~new_n29224_ & new_n29226_;
  assign new_n29228_ = ~pi0619 & new_n29222_;
  assign new_n29229_ = pi0619 & new_n29203_;
  assign new_n29230_ = ~pi1159 & ~new_n29229_;
  assign new_n29231_ = ~new_n29228_ & new_n29230_;
  assign new_n29232_ = ~new_n29227_ & ~new_n29231_;
  assign new_n29233_ = pi0789 & ~new_n29232_;
  assign new_n29234_ = ~new_n29223_ & ~new_n29233_;
  assign new_n29235_ = ~new_n17968_ & new_n29234_;
  assign new_n29236_ = new_n17968_ & new_n29203_;
  assign new_n29237_ = ~new_n29235_ & ~new_n29236_;
  assign new_n29238_ = ~new_n17762_ & ~new_n29237_;
  assign new_n29239_ = new_n17762_ & new_n29203_;
  assign new_n29240_ = ~new_n29238_ & ~new_n29239_;
  assign new_n29241_ = ~new_n20556_ & new_n29240_;
  assign new_n29242_ = pi0703 & new_n16915_;
  assign new_n29243_ = ~new_n29203_ & ~new_n29242_;
  assign new_n29244_ = ~pi0778 & new_n29243_;
  assign new_n29245_ = ~pi0625 & new_n29242_;
  assign new_n29246_ = ~new_n29243_ & ~new_n29245_;
  assign new_n29247_ = pi1153 & ~new_n29246_;
  assign new_n29248_ = ~pi1153 & ~new_n29203_;
  assign new_n29249_ = ~new_n29245_ & new_n29248_;
  assign new_n29250_ = ~new_n29247_ & ~new_n29249_;
  assign new_n29251_ = pi0778 & ~new_n29250_;
  assign new_n29252_ = ~new_n29244_ & ~new_n29251_;
  assign new_n29253_ = ~new_n17844_ & new_n29252_;
  assign new_n29254_ = ~new_n17846_ & new_n29253_;
  assign new_n29255_ = ~new_n17848_ & new_n29254_;
  assign new_n29256_ = ~new_n17980_ & new_n29255_;
  assign new_n29257_ = ~new_n18011_ & new_n29256_;
  assign new_n29258_ = ~pi0647 & new_n29257_;
  assign new_n29259_ = pi0647 & new_n29203_;
  assign new_n29260_ = ~pi1157 & ~new_n29259_;
  assign new_n29261_ = ~new_n29258_ & new_n29260_;
  assign new_n29262_ = pi0630 & new_n29261_;
  assign new_n29263_ = pi0647 & ~new_n29257_;
  assign new_n29264_ = ~pi0647 & ~new_n29203_;
  assign new_n29265_ = ~new_n29263_ & ~new_n29264_;
  assign new_n29266_ = new_n17801_ & ~new_n29265_;
  assign new_n29267_ = ~new_n29262_ & ~new_n29266_;
  assign new_n29268_ = ~new_n29241_ & new_n29267_;
  assign new_n29269_ = pi0787 & ~new_n29268_;
  assign new_n29270_ = pi0626 & ~new_n29234_;
  assign new_n29271_ = ~pi0626 & ~new_n29203_;
  assign new_n29272_ = new_n17731_ & ~new_n29271_;
  assign new_n29273_ = ~new_n29270_ & new_n29272_;
  assign new_n29274_ = new_n17856_ & new_n29255_;
  assign new_n29275_ = ~pi0626 & ~new_n29234_;
  assign new_n29276_ = pi0626 & ~new_n29203_;
  assign new_n29277_ = new_n17732_ & ~new_n29276_;
  assign new_n29278_ = ~new_n29275_ & new_n29277_;
  assign new_n29279_ = ~new_n29274_ & ~new_n29278_;
  assign new_n29280_ = ~new_n29273_ & new_n29279_;
  assign new_n29281_ = pi0788 & ~new_n29280_;
  assign new_n29282_ = ~new_n16639_ & ~new_n29243_;
  assign new_n29283_ = pi0625 & new_n29282_;
  assign new_n29284_ = new_n29205_ & ~new_n29282_;
  assign new_n29285_ = ~new_n29283_ & ~new_n29284_;
  assign new_n29286_ = new_n29248_ & ~new_n29285_;
  assign new_n29287_ = ~pi0608 & ~new_n29247_;
  assign new_n29288_ = ~new_n29286_ & new_n29287_;
  assign new_n29289_ = pi1153 & new_n29205_;
  assign new_n29290_ = ~new_n29283_ & new_n29289_;
  assign new_n29291_ = pi0608 & ~new_n29249_;
  assign new_n29292_ = ~new_n29290_ & new_n29291_;
  assign new_n29293_ = ~new_n29288_ & ~new_n29292_;
  assign new_n29294_ = pi0778 & ~new_n29293_;
  assign new_n29295_ = ~pi0778 & ~new_n29284_;
  assign new_n29296_ = ~new_n29294_ & ~new_n29295_;
  assign new_n29297_ = ~pi0609 & ~new_n29296_;
  assign new_n29298_ = pi0609 & new_n29252_;
  assign new_n29299_ = ~pi1155 & ~new_n29298_;
  assign new_n29300_ = ~new_n29297_ & new_n29299_;
  assign new_n29301_ = ~pi0660 & ~new_n29209_;
  assign new_n29302_ = ~new_n29300_ & new_n29301_;
  assign new_n29303_ = pi0609 & ~new_n29296_;
  assign new_n29304_ = ~pi0609 & new_n29252_;
  assign new_n29305_ = pi1155 & ~new_n29304_;
  assign new_n29306_ = ~new_n29303_ & new_n29305_;
  assign new_n29307_ = pi0660 & ~new_n29211_;
  assign new_n29308_ = ~new_n29306_ & new_n29307_;
  assign new_n29309_ = ~new_n29302_ & ~new_n29308_;
  assign new_n29310_ = pi0785 & ~new_n29309_;
  assign new_n29311_ = ~pi0785 & ~new_n29296_;
  assign new_n29312_ = ~new_n29310_ & ~new_n29311_;
  assign new_n29313_ = ~pi0618 & ~new_n29312_;
  assign new_n29314_ = pi0618 & new_n29253_;
  assign new_n29315_ = ~pi1154 & ~new_n29314_;
  assign new_n29316_ = ~new_n29313_ & new_n29315_;
  assign new_n29317_ = ~pi0627 & ~new_n29217_;
  assign new_n29318_ = ~new_n29316_ & new_n29317_;
  assign new_n29319_ = pi0618 & ~new_n29312_;
  assign new_n29320_ = ~pi0618 & new_n29253_;
  assign new_n29321_ = pi1154 & ~new_n29320_;
  assign new_n29322_ = ~new_n29319_ & new_n29321_;
  assign new_n29323_ = pi0627 & ~new_n29219_;
  assign new_n29324_ = ~new_n29322_ & new_n29323_;
  assign new_n29325_ = ~new_n29318_ & ~new_n29324_;
  assign new_n29326_ = pi0781 & ~new_n29325_;
  assign new_n29327_ = ~pi0781 & ~new_n29312_;
  assign new_n29328_ = ~new_n29326_ & ~new_n29327_;
  assign new_n29329_ = pi0619 & ~new_n29328_;
  assign new_n29330_ = ~pi0619 & new_n29254_;
  assign new_n29331_ = pi1159 & ~new_n29330_;
  assign new_n29332_ = ~new_n29329_ & new_n29331_;
  assign new_n29333_ = pi0648 & ~new_n29231_;
  assign new_n29334_ = ~new_n29332_ & new_n29333_;
  assign new_n29335_ = ~pi0619 & ~new_n29328_;
  assign new_n29336_ = pi0619 & new_n29254_;
  assign new_n29337_ = ~pi1159 & ~new_n29336_;
  assign new_n29338_ = ~new_n29335_ & new_n29337_;
  assign new_n29339_ = ~pi0648 & ~new_n29227_;
  assign new_n29340_ = ~new_n29338_ & new_n29339_;
  assign new_n29341_ = pi0789 & ~new_n29340_;
  assign new_n29342_ = ~new_n29334_ & new_n29341_;
  assign new_n29343_ = ~pi0789 & new_n29328_;
  assign new_n29344_ = new_n17969_ & ~new_n29343_;
  assign new_n29345_ = ~new_n29342_ & new_n29344_;
  assign new_n29346_ = ~new_n29281_ & ~new_n29345_;
  assign new_n29347_ = ~new_n20364_ & ~new_n29346_;
  assign new_n29348_ = new_n18008_ & ~new_n29237_;
  assign new_n29349_ = new_n20851_ & new_n29256_;
  assign new_n29350_ = ~new_n29348_ & ~new_n29349_;
  assign new_n29351_ = ~pi0629 & ~new_n29350_;
  assign new_n29352_ = new_n20855_ & new_n29256_;
  assign new_n29353_ = new_n18007_ & ~new_n29237_;
  assign new_n29354_ = ~new_n29352_ & ~new_n29353_;
  assign new_n29355_ = pi0629 & ~new_n29354_;
  assign new_n29356_ = ~new_n29351_ & ~new_n29355_;
  assign new_n29357_ = pi0792 & ~new_n29356_;
  assign new_n29358_ = ~new_n20360_ & ~new_n29357_;
  assign new_n29359_ = ~new_n29347_ & new_n29358_;
  assign new_n29360_ = ~new_n29269_ & ~new_n29359_;
  assign new_n29361_ = pi0644 & new_n29360_;
  assign new_n29362_ = ~pi0787 & ~new_n29257_;
  assign new_n29363_ = pi1157 & ~new_n29265_;
  assign new_n29364_ = ~new_n29261_ & ~new_n29363_;
  assign new_n29365_ = pi0787 & ~new_n29364_;
  assign new_n29366_ = ~new_n29362_ & ~new_n29365_;
  assign new_n29367_ = ~pi0644 & new_n29366_;
  assign new_n29368_ = pi0715 & ~new_n29367_;
  assign new_n29369_ = ~new_n29361_ & new_n29368_;
  assign new_n29370_ = ~new_n17804_ & ~new_n29240_;
  assign new_n29371_ = new_n17804_ & new_n29203_;
  assign new_n29372_ = ~new_n29370_ & ~new_n29371_;
  assign new_n29373_ = pi0644 & ~new_n29372_;
  assign new_n29374_ = ~pi0644 & new_n29203_;
  assign new_n29375_ = ~pi0715 & ~new_n29374_;
  assign new_n29376_ = ~new_n29373_ & new_n29375_;
  assign new_n29377_ = pi1160 & ~new_n29376_;
  assign new_n29378_ = ~new_n29369_ & new_n29377_;
  assign new_n29379_ = ~pi0644 & new_n29360_;
  assign new_n29380_ = pi0644 & new_n29366_;
  assign new_n29381_ = ~pi0715 & ~new_n29380_;
  assign new_n29382_ = ~new_n29379_ & new_n29381_;
  assign new_n29383_ = ~pi0644 & ~new_n29372_;
  assign new_n29384_ = pi0644 & new_n29203_;
  assign new_n29385_ = pi0715 & ~new_n29384_;
  assign new_n29386_ = ~new_n29383_ & new_n29385_;
  assign new_n29387_ = ~pi1160 & ~new_n29386_;
  assign new_n29388_ = ~new_n29382_ & new_n29387_;
  assign new_n29389_ = ~new_n29378_ & ~new_n29388_;
  assign new_n29390_ = pi0790 & ~new_n29389_;
  assign new_n29391_ = ~pi0790 & new_n29360_;
  assign new_n29392_ = pi0832 & ~new_n29391_;
  assign new_n29393_ = ~new_n29390_ & new_n29392_;
  assign po0343 = ~new_n29202_ & ~new_n29393_;
  assign new_n29395_ = pi0187 & ~new_n3272_;
  assign new_n29396_ = ~pi0770 & ~new_n19376_;
  assign new_n29397_ = ~new_n21011_ & ~new_n29396_;
  assign new_n29398_ = ~pi0187 & ~new_n29397_;
  assign new_n29399_ = ~pi0187 & ~new_n19370_;
  assign new_n29400_ = ~pi0770 & ~new_n29399_;
  assign new_n29401_ = ~new_n24446_ & new_n29400_;
  assign new_n29402_ = ~new_n29398_ & ~new_n29401_;
  assign new_n29403_ = ~pi0726 & ~new_n29402_;
  assign new_n29404_ = ~pi0187 & new_n19389_;
  assign new_n29405_ = pi0187 & new_n19394_;
  assign new_n29406_ = pi0770 & ~new_n19396_;
  assign new_n29407_ = ~new_n29405_ & new_n29406_;
  assign new_n29408_ = ~new_n29404_ & new_n29407_;
  assign new_n29409_ = pi0187 & new_n19406_;
  assign new_n29410_ = ~pi0187 & ~new_n19414_;
  assign new_n29411_ = ~pi0770 & ~new_n29410_;
  assign new_n29412_ = ~new_n29409_ & new_n29411_;
  assign new_n29413_ = pi0726 & ~new_n29412_;
  assign new_n29414_ = ~new_n29408_ & new_n29413_;
  assign new_n29415_ = new_n3272_ & ~new_n29414_;
  assign new_n29416_ = ~new_n29403_ & new_n29415_;
  assign new_n29417_ = ~new_n29395_ & ~new_n29416_;
  assign new_n29418_ = ~pi0625 & new_n29417_;
  assign new_n29419_ = new_n3272_ & new_n29402_;
  assign new_n29420_ = ~new_n29395_ & ~new_n29419_;
  assign new_n29421_ = pi0625 & new_n29420_;
  assign new_n29422_ = ~pi1153 & ~new_n29421_;
  assign new_n29423_ = ~new_n29418_ & new_n29422_;
  assign new_n29424_ = ~pi0187 & new_n18124_;
  assign new_n29425_ = pi0187 & ~new_n18128_;
  assign new_n29426_ = ~pi0038 & ~new_n29425_;
  assign new_n29427_ = ~new_n29424_ & new_n29426_;
  assign new_n29428_ = ~pi0187 & ~new_n17431_;
  assign new_n29429_ = new_n17544_ & ~new_n29428_;
  assign new_n29430_ = pi0726 & ~new_n29429_;
  assign new_n29431_ = ~new_n29427_ & new_n29430_;
  assign new_n29432_ = ~pi0187 & ~pi0726;
  assign new_n29433_ = ~new_n17551_ & new_n29432_;
  assign new_n29434_ = new_n3272_ & ~new_n29433_;
  assign new_n29435_ = ~new_n29431_ & new_n29434_;
  assign new_n29436_ = ~new_n29395_ & ~new_n29435_;
  assign new_n29437_ = pi0625 & new_n29436_;
  assign new_n29438_ = ~pi0187 & ~new_n17558_;
  assign new_n29439_ = ~pi0625 & new_n29438_;
  assign new_n29440_ = pi1153 & ~new_n29439_;
  assign new_n29441_ = ~new_n29437_ & new_n29440_;
  assign new_n29442_ = ~pi0608 & ~new_n29441_;
  assign new_n29443_ = ~new_n29423_ & new_n29442_;
  assign new_n29444_ = pi0625 & new_n29417_;
  assign new_n29445_ = ~pi0625 & new_n29420_;
  assign new_n29446_ = pi1153 & ~new_n29445_;
  assign new_n29447_ = ~new_n29444_ & new_n29446_;
  assign new_n29448_ = ~pi0625 & new_n29436_;
  assign new_n29449_ = pi0625 & new_n29438_;
  assign new_n29450_ = ~pi1153 & ~new_n29449_;
  assign new_n29451_ = ~new_n29448_ & new_n29450_;
  assign new_n29452_ = pi0608 & ~new_n29451_;
  assign new_n29453_ = ~new_n29447_ & new_n29452_;
  assign new_n29454_ = ~new_n29443_ & ~new_n29453_;
  assign new_n29455_ = pi0778 & ~new_n29454_;
  assign new_n29456_ = ~pi0778 & new_n29417_;
  assign new_n29457_ = ~new_n29455_ & ~new_n29456_;
  assign new_n29458_ = ~pi0609 & ~new_n29457_;
  assign new_n29459_ = ~pi0778 & ~new_n29436_;
  assign new_n29460_ = ~new_n29441_ & ~new_n29451_;
  assign new_n29461_ = pi0778 & ~new_n29460_;
  assign new_n29462_ = ~new_n29459_ & ~new_n29461_;
  assign new_n29463_ = pi0609 & new_n29462_;
  assign new_n29464_ = ~pi1155 & ~new_n29463_;
  assign new_n29465_ = ~new_n29458_ & new_n29464_;
  assign new_n29466_ = ~new_n17591_ & ~new_n29438_;
  assign new_n29467_ = ~new_n17590_ & ~new_n29420_;
  assign new_n29468_ = pi0609 & new_n29467_;
  assign new_n29469_ = ~new_n29466_ & ~new_n29468_;
  assign new_n29470_ = pi1155 & ~new_n29469_;
  assign new_n29471_ = ~pi0660 & ~new_n29470_;
  assign new_n29472_ = ~new_n29465_ & new_n29471_;
  assign new_n29473_ = pi0609 & ~new_n29457_;
  assign new_n29474_ = ~pi0609 & new_n29462_;
  assign new_n29475_ = pi1155 & ~new_n29474_;
  assign new_n29476_ = ~new_n29473_ & new_n29475_;
  assign new_n29477_ = ~new_n17603_ & ~new_n29438_;
  assign new_n29478_ = ~pi0609 & new_n29467_;
  assign new_n29479_ = ~new_n29477_ & ~new_n29478_;
  assign new_n29480_ = ~pi1155 & ~new_n29479_;
  assign new_n29481_ = pi0660 & ~new_n29480_;
  assign new_n29482_ = ~new_n29476_ & new_n29481_;
  assign new_n29483_ = ~new_n29472_ & ~new_n29482_;
  assign new_n29484_ = pi0785 & ~new_n29483_;
  assign new_n29485_ = ~pi0785 & ~new_n29457_;
  assign new_n29486_ = ~new_n29484_ & ~new_n29485_;
  assign new_n29487_ = ~pi0618 & ~new_n29486_;
  assign new_n29488_ = ~new_n17618_ & ~new_n29462_;
  assign new_n29489_ = new_n17618_ & ~new_n29438_;
  assign new_n29490_ = ~new_n29488_ & ~new_n29489_;
  assign new_n29491_ = pi0618 & new_n29490_;
  assign new_n29492_ = ~pi1154 & ~new_n29491_;
  assign new_n29493_ = ~new_n29487_ & new_n29492_;
  assign new_n29494_ = new_n17590_ & ~new_n29438_;
  assign new_n29495_ = ~new_n29467_ & ~new_n29494_;
  assign new_n29496_ = ~pi0785 & ~new_n29495_;
  assign new_n29497_ = ~new_n29470_ & ~new_n29480_;
  assign new_n29498_ = pi0785 & ~new_n29497_;
  assign new_n29499_ = ~new_n29496_ & ~new_n29498_;
  assign new_n29500_ = pi0618 & new_n29499_;
  assign new_n29501_ = ~pi0618 & new_n29438_;
  assign new_n29502_ = pi1154 & ~new_n29501_;
  assign new_n29503_ = ~new_n29500_ & new_n29502_;
  assign new_n29504_ = ~pi0627 & ~new_n29503_;
  assign new_n29505_ = ~new_n29493_ & new_n29504_;
  assign new_n29506_ = pi0618 & ~new_n29486_;
  assign new_n29507_ = ~pi0618 & new_n29490_;
  assign new_n29508_ = pi1154 & ~new_n29507_;
  assign new_n29509_ = ~new_n29506_ & new_n29508_;
  assign new_n29510_ = ~pi0618 & new_n29499_;
  assign new_n29511_ = pi0618 & new_n29438_;
  assign new_n29512_ = ~pi1154 & ~new_n29511_;
  assign new_n29513_ = ~new_n29510_ & new_n29512_;
  assign new_n29514_ = pi0627 & ~new_n29513_;
  assign new_n29515_ = ~new_n29509_ & new_n29514_;
  assign new_n29516_ = ~new_n29505_ & ~new_n29515_;
  assign new_n29517_ = pi0781 & ~new_n29516_;
  assign new_n29518_ = ~pi0781 & ~new_n29486_;
  assign new_n29519_ = ~new_n29517_ & ~new_n29518_;
  assign new_n29520_ = ~pi0619 & ~new_n29519_;
  assign new_n29521_ = ~new_n17655_ & new_n29490_;
  assign new_n29522_ = new_n17655_ & new_n29438_;
  assign new_n29523_ = ~new_n29521_ & ~new_n29522_;
  assign new_n29524_ = pi0619 & ~new_n29523_;
  assign new_n29525_ = ~pi1159 & ~new_n29524_;
  assign new_n29526_ = ~new_n29520_ & new_n29525_;
  assign new_n29527_ = ~pi0781 & ~new_n29499_;
  assign new_n29528_ = ~new_n29503_ & ~new_n29513_;
  assign new_n29529_ = pi0781 & ~new_n29528_;
  assign new_n29530_ = ~new_n29527_ & ~new_n29529_;
  assign new_n29531_ = pi0619 & new_n29530_;
  assign new_n29532_ = ~pi0619 & new_n29438_;
  assign new_n29533_ = pi1159 & ~new_n29532_;
  assign new_n29534_ = ~new_n29531_ & new_n29533_;
  assign new_n29535_ = ~pi0648 & ~new_n29534_;
  assign new_n29536_ = ~new_n29526_ & new_n29535_;
  assign new_n29537_ = pi0619 & ~new_n29519_;
  assign new_n29538_ = ~pi0619 & ~new_n29523_;
  assign new_n29539_ = pi1159 & ~new_n29538_;
  assign new_n29540_ = ~new_n29537_ & new_n29539_;
  assign new_n29541_ = ~pi0619 & new_n29530_;
  assign new_n29542_ = pi0619 & new_n29438_;
  assign new_n29543_ = ~pi1159 & ~new_n29542_;
  assign new_n29544_ = ~new_n29541_ & new_n29543_;
  assign new_n29545_ = pi0648 & ~new_n29544_;
  assign new_n29546_ = ~new_n29540_ & new_n29545_;
  assign new_n29547_ = ~new_n29536_ & ~new_n29546_;
  assign new_n29548_ = pi0789 & ~new_n29547_;
  assign new_n29549_ = ~pi0789 & ~new_n29519_;
  assign new_n29550_ = ~new_n29548_ & ~new_n29549_;
  assign new_n29551_ = ~pi0788 & new_n29550_;
  assign new_n29552_ = ~pi0626 & new_n29550_;
  assign new_n29553_ = new_n17691_ & ~new_n29438_;
  assign new_n29554_ = ~new_n17691_ & new_n29523_;
  assign new_n29555_ = ~new_n29553_ & ~new_n29554_;
  assign new_n29556_ = pi0626 & ~new_n29555_;
  assign new_n29557_ = ~pi0641 & ~new_n29556_;
  assign new_n29558_ = ~new_n29552_ & new_n29557_;
  assign new_n29559_ = ~pi0789 & ~new_n29530_;
  assign new_n29560_ = ~new_n29534_ & ~new_n29544_;
  assign new_n29561_ = pi0789 & ~new_n29560_;
  assign new_n29562_ = ~new_n29559_ & ~new_n29561_;
  assign new_n29563_ = ~pi0626 & ~new_n29562_;
  assign new_n29564_ = pi0626 & ~new_n29438_;
  assign new_n29565_ = pi0641 & ~new_n29564_;
  assign new_n29566_ = ~new_n29563_ & new_n29565_;
  assign new_n29567_ = ~pi1158 & ~new_n29566_;
  assign new_n29568_ = ~new_n29558_ & new_n29567_;
  assign new_n29569_ = pi0626 & new_n29550_;
  assign new_n29570_ = ~pi0626 & ~new_n29555_;
  assign new_n29571_ = pi0641 & ~new_n29570_;
  assign new_n29572_ = ~new_n29569_ & new_n29571_;
  assign new_n29573_ = pi0626 & ~new_n29562_;
  assign new_n29574_ = ~pi0626 & ~new_n29438_;
  assign new_n29575_ = ~pi0641 & ~new_n29574_;
  assign new_n29576_ = ~new_n29573_ & new_n29575_;
  assign new_n29577_ = pi1158 & ~new_n29576_;
  assign new_n29578_ = ~new_n29572_ & new_n29577_;
  assign new_n29579_ = ~new_n29568_ & ~new_n29578_;
  assign new_n29580_ = pi0788 & ~new_n29579_;
  assign new_n29581_ = ~new_n29551_ & ~new_n29580_;
  assign new_n29582_ = ~pi0628 & new_n29581_;
  assign new_n29583_ = ~new_n17968_ & new_n29562_;
  assign new_n29584_ = new_n17968_ & new_n29438_;
  assign new_n29585_ = ~new_n29583_ & ~new_n29584_;
  assign new_n29586_ = pi0628 & ~new_n29585_;
  assign new_n29587_ = ~pi1156 & ~new_n29586_;
  assign new_n29588_ = ~new_n29582_ & new_n29587_;
  assign new_n29589_ = ~new_n17734_ & new_n29555_;
  assign new_n29590_ = new_n17734_ & new_n29438_;
  assign new_n29591_ = ~new_n29589_ & ~new_n29590_;
  assign new_n29592_ = pi0628 & ~new_n29591_;
  assign new_n29593_ = ~pi0628 & new_n29438_;
  assign new_n29594_ = pi1156 & ~new_n29593_;
  assign new_n29595_ = ~new_n29592_ & new_n29594_;
  assign new_n29596_ = ~pi0629 & ~new_n29595_;
  assign new_n29597_ = ~new_n29588_ & new_n29596_;
  assign new_n29598_ = pi0628 & new_n29581_;
  assign new_n29599_ = ~pi0628 & ~new_n29585_;
  assign new_n29600_ = pi1156 & ~new_n29599_;
  assign new_n29601_ = ~new_n29598_ & new_n29600_;
  assign new_n29602_ = ~pi0628 & ~new_n29591_;
  assign new_n29603_ = pi0628 & new_n29438_;
  assign new_n29604_ = ~pi1156 & ~new_n29603_;
  assign new_n29605_ = ~new_n29602_ & new_n29604_;
  assign new_n29606_ = pi0629 & ~new_n29605_;
  assign new_n29607_ = ~new_n29601_ & new_n29606_;
  assign new_n29608_ = ~new_n29597_ & ~new_n29607_;
  assign new_n29609_ = pi0792 & ~new_n29608_;
  assign new_n29610_ = ~pi0792 & new_n29581_;
  assign new_n29611_ = ~new_n29609_ & ~new_n29610_;
  assign new_n29612_ = ~pi0647 & ~new_n29611_;
  assign new_n29613_ = ~new_n17762_ & ~new_n29585_;
  assign new_n29614_ = new_n17762_ & new_n29438_;
  assign new_n29615_ = ~new_n29613_ & ~new_n29614_;
  assign new_n29616_ = pi0647 & ~new_n29615_;
  assign new_n29617_ = ~pi1157 & ~new_n29616_;
  assign new_n29618_ = ~new_n29612_ & new_n29617_;
  assign new_n29619_ = ~pi0792 & new_n29591_;
  assign new_n29620_ = ~new_n29595_ & ~new_n29605_;
  assign new_n29621_ = pi0792 & ~new_n29620_;
  assign new_n29622_ = ~new_n29619_ & ~new_n29621_;
  assign new_n29623_ = pi0647 & new_n29622_;
  assign new_n29624_ = ~pi0647 & new_n29438_;
  assign new_n29625_ = pi1157 & ~new_n29624_;
  assign new_n29626_ = ~new_n29623_ & new_n29625_;
  assign new_n29627_ = ~pi0630 & ~new_n29626_;
  assign new_n29628_ = ~new_n29618_ & new_n29627_;
  assign new_n29629_ = pi0647 & ~new_n29611_;
  assign new_n29630_ = ~pi0647 & ~new_n29615_;
  assign new_n29631_ = pi1157 & ~new_n29630_;
  assign new_n29632_ = ~new_n29629_ & new_n29631_;
  assign new_n29633_ = ~pi0647 & new_n29622_;
  assign new_n29634_ = pi0647 & new_n29438_;
  assign new_n29635_ = ~pi1157 & ~new_n29634_;
  assign new_n29636_ = ~new_n29633_ & new_n29635_;
  assign new_n29637_ = pi0630 & ~new_n29636_;
  assign new_n29638_ = ~new_n29632_ & new_n29637_;
  assign new_n29639_ = ~new_n29628_ & ~new_n29638_;
  assign new_n29640_ = pi0787 & ~new_n29639_;
  assign new_n29641_ = ~pi0787 & ~new_n29611_;
  assign new_n29642_ = ~new_n29640_ & ~new_n29641_;
  assign new_n29643_ = ~pi0644 & ~new_n29642_;
  assign new_n29644_ = ~pi0787 & ~new_n29622_;
  assign new_n29645_ = ~new_n29626_ & ~new_n29636_;
  assign new_n29646_ = pi0787 & ~new_n29645_;
  assign new_n29647_ = ~new_n29644_ & ~new_n29646_;
  assign new_n29648_ = pi0644 & new_n29647_;
  assign new_n29649_ = ~pi0715 & ~new_n29648_;
  assign new_n29650_ = ~new_n29643_ & new_n29649_;
  assign new_n29651_ = new_n17804_ & ~new_n29438_;
  assign new_n29652_ = ~new_n17804_ & new_n29615_;
  assign new_n29653_ = ~new_n29651_ & ~new_n29652_;
  assign new_n29654_ = ~pi0644 & new_n29653_;
  assign new_n29655_ = pi0644 & new_n29438_;
  assign new_n29656_ = pi0715 & ~new_n29655_;
  assign new_n29657_ = ~new_n29654_ & new_n29656_;
  assign new_n29658_ = ~pi1160 & ~new_n29657_;
  assign new_n29659_ = ~new_n29650_ & new_n29658_;
  assign new_n29660_ = pi0644 & ~new_n29642_;
  assign new_n29661_ = ~pi0644 & new_n29647_;
  assign new_n29662_ = pi0715 & ~new_n29661_;
  assign new_n29663_ = ~new_n29660_ & new_n29662_;
  assign new_n29664_ = pi0644 & new_n29653_;
  assign new_n29665_ = ~pi0644 & new_n29438_;
  assign new_n29666_ = ~pi0715 & ~new_n29665_;
  assign new_n29667_ = ~new_n29664_ & new_n29666_;
  assign new_n29668_ = pi1160 & ~new_n29667_;
  assign new_n29669_ = ~new_n29663_ & new_n29668_;
  assign new_n29670_ = pi0790 & ~new_n29669_;
  assign new_n29671_ = ~new_n29659_ & new_n29670_;
  assign new_n29672_ = ~pi0790 & new_n29642_;
  assign new_n29673_ = ~po1038 & ~new_n29672_;
  assign new_n29674_ = ~new_n29671_ & new_n29673_;
  assign new_n29675_ = ~pi0187 & po1038;
  assign new_n29676_ = ~pi0832 & ~new_n29675_;
  assign new_n29677_ = ~new_n29674_ & new_n29676_;
  assign new_n29678_ = ~pi0187 & ~new_n2754_;
  assign new_n29679_ = ~pi0770 & new_n16913_;
  assign new_n29680_ = ~new_n29678_ & ~new_n29679_;
  assign new_n29681_ = ~new_n17858_ & ~new_n29680_;
  assign new_n29682_ = ~pi0785 & ~new_n29681_;
  assign new_n29683_ = ~new_n17863_ & ~new_n29680_;
  assign new_n29684_ = pi1155 & ~new_n29683_;
  assign new_n29685_ = ~new_n17866_ & new_n29681_;
  assign new_n29686_ = ~pi1155 & ~new_n29685_;
  assign new_n29687_ = ~new_n29684_ & ~new_n29686_;
  assign new_n29688_ = pi0785 & ~new_n29687_;
  assign new_n29689_ = ~new_n29682_ & ~new_n29688_;
  assign new_n29690_ = ~pi0781 & ~new_n29689_;
  assign new_n29691_ = ~new_n17873_ & new_n29689_;
  assign new_n29692_ = pi1154 & ~new_n29691_;
  assign new_n29693_ = ~new_n17876_ & new_n29689_;
  assign new_n29694_ = ~pi1154 & ~new_n29693_;
  assign new_n29695_ = ~new_n29692_ & ~new_n29694_;
  assign new_n29696_ = pi0781 & ~new_n29695_;
  assign new_n29697_ = ~new_n29690_ & ~new_n29696_;
  assign new_n29698_ = ~pi0789 & ~new_n29697_;
  assign new_n29699_ = pi0619 & new_n29697_;
  assign new_n29700_ = ~pi0619 & new_n29678_;
  assign new_n29701_ = pi1159 & ~new_n29700_;
  assign new_n29702_ = ~new_n29699_ & new_n29701_;
  assign new_n29703_ = ~pi0619 & new_n29697_;
  assign new_n29704_ = pi0619 & new_n29678_;
  assign new_n29705_ = ~pi1159 & ~new_n29704_;
  assign new_n29706_ = ~new_n29703_ & new_n29705_;
  assign new_n29707_ = ~new_n29702_ & ~new_n29706_;
  assign new_n29708_ = pi0789 & ~new_n29707_;
  assign new_n29709_ = ~new_n29698_ & ~new_n29708_;
  assign new_n29710_ = ~new_n17968_ & new_n29709_;
  assign new_n29711_ = new_n17968_ & new_n29678_;
  assign new_n29712_ = ~new_n29710_ & ~new_n29711_;
  assign new_n29713_ = ~new_n17762_ & ~new_n29712_;
  assign new_n29714_ = new_n17762_ & new_n29678_;
  assign new_n29715_ = ~new_n29713_ & ~new_n29714_;
  assign new_n29716_ = ~new_n20556_ & new_n29715_;
  assign new_n29717_ = pi0726 & new_n16915_;
  assign new_n29718_ = ~new_n29678_ & ~new_n29717_;
  assign new_n29719_ = ~pi0778 & new_n29718_;
  assign new_n29720_ = ~pi0625 & new_n29717_;
  assign new_n29721_ = ~new_n29718_ & ~new_n29720_;
  assign new_n29722_ = pi1153 & ~new_n29721_;
  assign new_n29723_ = ~pi1153 & ~new_n29678_;
  assign new_n29724_ = ~new_n29720_ & new_n29723_;
  assign new_n29725_ = ~new_n29722_ & ~new_n29724_;
  assign new_n29726_ = pi0778 & ~new_n29725_;
  assign new_n29727_ = ~new_n29719_ & ~new_n29726_;
  assign new_n29728_ = ~new_n17844_ & new_n29727_;
  assign new_n29729_ = ~new_n17846_ & new_n29728_;
  assign new_n29730_ = ~new_n17848_ & new_n29729_;
  assign new_n29731_ = ~new_n17980_ & new_n29730_;
  assign new_n29732_ = ~new_n18011_ & new_n29731_;
  assign new_n29733_ = ~pi0647 & new_n29732_;
  assign new_n29734_ = pi0647 & new_n29678_;
  assign new_n29735_ = ~pi1157 & ~new_n29734_;
  assign new_n29736_ = ~new_n29733_ & new_n29735_;
  assign new_n29737_ = pi0630 & new_n29736_;
  assign new_n29738_ = pi0647 & ~new_n29732_;
  assign new_n29739_ = ~pi0647 & ~new_n29678_;
  assign new_n29740_ = ~new_n29738_ & ~new_n29739_;
  assign new_n29741_ = new_n17801_ & ~new_n29740_;
  assign new_n29742_ = ~new_n29737_ & ~new_n29741_;
  assign new_n29743_ = ~new_n29716_ & new_n29742_;
  assign new_n29744_ = pi0787 & ~new_n29743_;
  assign new_n29745_ = pi0626 & ~new_n29709_;
  assign new_n29746_ = ~pi0626 & ~new_n29678_;
  assign new_n29747_ = new_n17731_ & ~new_n29746_;
  assign new_n29748_ = ~new_n29745_ & new_n29747_;
  assign new_n29749_ = new_n17856_ & new_n29730_;
  assign new_n29750_ = ~pi0626 & ~new_n29709_;
  assign new_n29751_ = pi0626 & ~new_n29678_;
  assign new_n29752_ = new_n17732_ & ~new_n29751_;
  assign new_n29753_ = ~new_n29750_ & new_n29752_;
  assign new_n29754_ = ~new_n29749_ & ~new_n29753_;
  assign new_n29755_ = ~new_n29748_ & new_n29754_;
  assign new_n29756_ = pi0788 & ~new_n29755_;
  assign new_n29757_ = ~new_n16639_ & ~new_n29718_;
  assign new_n29758_ = pi0625 & new_n29757_;
  assign new_n29759_ = new_n29680_ & ~new_n29757_;
  assign new_n29760_ = ~new_n29758_ & ~new_n29759_;
  assign new_n29761_ = new_n29723_ & ~new_n29760_;
  assign new_n29762_ = ~pi0608 & ~new_n29722_;
  assign new_n29763_ = ~new_n29761_ & new_n29762_;
  assign new_n29764_ = pi1153 & new_n29680_;
  assign new_n29765_ = ~new_n29758_ & new_n29764_;
  assign new_n29766_ = pi0608 & ~new_n29724_;
  assign new_n29767_ = ~new_n29765_ & new_n29766_;
  assign new_n29768_ = ~new_n29763_ & ~new_n29767_;
  assign new_n29769_ = pi0778 & ~new_n29768_;
  assign new_n29770_ = ~pi0778 & ~new_n29759_;
  assign new_n29771_ = ~new_n29769_ & ~new_n29770_;
  assign new_n29772_ = ~pi0609 & ~new_n29771_;
  assign new_n29773_ = pi0609 & new_n29727_;
  assign new_n29774_ = ~pi1155 & ~new_n29773_;
  assign new_n29775_ = ~new_n29772_ & new_n29774_;
  assign new_n29776_ = ~pi0660 & ~new_n29684_;
  assign new_n29777_ = ~new_n29775_ & new_n29776_;
  assign new_n29778_ = pi0609 & ~new_n29771_;
  assign new_n29779_ = ~pi0609 & new_n29727_;
  assign new_n29780_ = pi1155 & ~new_n29779_;
  assign new_n29781_ = ~new_n29778_ & new_n29780_;
  assign new_n29782_ = pi0660 & ~new_n29686_;
  assign new_n29783_ = ~new_n29781_ & new_n29782_;
  assign new_n29784_ = ~new_n29777_ & ~new_n29783_;
  assign new_n29785_ = pi0785 & ~new_n29784_;
  assign new_n29786_ = ~pi0785 & ~new_n29771_;
  assign new_n29787_ = ~new_n29785_ & ~new_n29786_;
  assign new_n29788_ = ~pi0618 & ~new_n29787_;
  assign new_n29789_ = pi0618 & new_n29728_;
  assign new_n29790_ = ~pi1154 & ~new_n29789_;
  assign new_n29791_ = ~new_n29788_ & new_n29790_;
  assign new_n29792_ = ~pi0627 & ~new_n29692_;
  assign new_n29793_ = ~new_n29791_ & new_n29792_;
  assign new_n29794_ = pi0618 & ~new_n29787_;
  assign new_n29795_ = ~pi0618 & new_n29728_;
  assign new_n29796_ = pi1154 & ~new_n29795_;
  assign new_n29797_ = ~new_n29794_ & new_n29796_;
  assign new_n29798_ = pi0627 & ~new_n29694_;
  assign new_n29799_ = ~new_n29797_ & new_n29798_;
  assign new_n29800_ = ~new_n29793_ & ~new_n29799_;
  assign new_n29801_ = pi0781 & ~new_n29800_;
  assign new_n29802_ = ~pi0781 & ~new_n29787_;
  assign new_n29803_ = ~new_n29801_ & ~new_n29802_;
  assign new_n29804_ = pi0619 & ~new_n29803_;
  assign new_n29805_ = ~pi0619 & new_n29729_;
  assign new_n29806_ = pi1159 & ~new_n29805_;
  assign new_n29807_ = ~new_n29804_ & new_n29806_;
  assign new_n29808_ = pi0648 & ~new_n29706_;
  assign new_n29809_ = ~new_n29807_ & new_n29808_;
  assign new_n29810_ = ~pi0619 & ~new_n29803_;
  assign new_n29811_ = pi0619 & new_n29729_;
  assign new_n29812_ = ~pi1159 & ~new_n29811_;
  assign new_n29813_ = ~new_n29810_ & new_n29812_;
  assign new_n29814_ = ~pi0648 & ~new_n29702_;
  assign new_n29815_ = ~new_n29813_ & new_n29814_;
  assign new_n29816_ = pi0789 & ~new_n29815_;
  assign new_n29817_ = ~new_n29809_ & new_n29816_;
  assign new_n29818_ = ~pi0789 & new_n29803_;
  assign new_n29819_ = new_n17969_ & ~new_n29818_;
  assign new_n29820_ = ~new_n29817_ & new_n29819_;
  assign new_n29821_ = ~new_n29756_ & ~new_n29820_;
  assign new_n29822_ = ~new_n20364_ & ~new_n29821_;
  assign new_n29823_ = new_n18008_ & ~new_n29712_;
  assign new_n29824_ = new_n20851_ & new_n29731_;
  assign new_n29825_ = ~new_n29823_ & ~new_n29824_;
  assign new_n29826_ = ~pi0629 & ~new_n29825_;
  assign new_n29827_ = new_n20855_ & new_n29731_;
  assign new_n29828_ = new_n18007_ & ~new_n29712_;
  assign new_n29829_ = ~new_n29827_ & ~new_n29828_;
  assign new_n29830_ = pi0629 & ~new_n29829_;
  assign new_n29831_ = ~new_n29826_ & ~new_n29830_;
  assign new_n29832_ = pi0792 & ~new_n29831_;
  assign new_n29833_ = ~new_n20360_ & ~new_n29832_;
  assign new_n29834_ = ~new_n29822_ & new_n29833_;
  assign new_n29835_ = ~new_n29744_ & ~new_n29834_;
  assign new_n29836_ = pi0644 & new_n29835_;
  assign new_n29837_ = ~pi0787 & ~new_n29732_;
  assign new_n29838_ = pi1157 & ~new_n29740_;
  assign new_n29839_ = ~new_n29736_ & ~new_n29838_;
  assign new_n29840_ = pi0787 & ~new_n29839_;
  assign new_n29841_ = ~new_n29837_ & ~new_n29840_;
  assign new_n29842_ = ~pi0644 & new_n29841_;
  assign new_n29843_ = pi0715 & ~new_n29842_;
  assign new_n29844_ = ~new_n29836_ & new_n29843_;
  assign new_n29845_ = ~new_n17804_ & ~new_n29715_;
  assign new_n29846_ = new_n17804_ & new_n29678_;
  assign new_n29847_ = ~new_n29845_ & ~new_n29846_;
  assign new_n29848_ = pi0644 & ~new_n29847_;
  assign new_n29849_ = ~pi0644 & new_n29678_;
  assign new_n29850_ = ~pi0715 & ~new_n29849_;
  assign new_n29851_ = ~new_n29848_ & new_n29850_;
  assign new_n29852_ = pi1160 & ~new_n29851_;
  assign new_n29853_ = ~new_n29844_ & new_n29852_;
  assign new_n29854_ = ~pi0644 & new_n29835_;
  assign new_n29855_ = pi0644 & new_n29841_;
  assign new_n29856_ = ~pi0715 & ~new_n29855_;
  assign new_n29857_ = ~new_n29854_ & new_n29856_;
  assign new_n29858_ = ~pi0644 & ~new_n29847_;
  assign new_n29859_ = pi0644 & new_n29678_;
  assign new_n29860_ = pi0715 & ~new_n29859_;
  assign new_n29861_ = ~new_n29858_ & new_n29860_;
  assign new_n29862_ = ~pi1160 & ~new_n29861_;
  assign new_n29863_ = ~new_n29857_ & new_n29862_;
  assign new_n29864_ = ~new_n29853_ & ~new_n29863_;
  assign new_n29865_ = pi0790 & ~new_n29864_;
  assign new_n29866_ = ~pi0790 & new_n29835_;
  assign new_n29867_ = pi0832 & ~new_n29866_;
  assign new_n29868_ = ~new_n29865_ & new_n29867_;
  assign po0344 = ~new_n29677_ & ~new_n29868_;
  assign new_n29870_ = pi0188 & ~new_n3272_;
  assign new_n29871_ = ~pi0768 & ~new_n19376_;
  assign new_n29872_ = ~new_n22338_ & ~new_n29871_;
  assign new_n29873_ = ~pi0188 & ~new_n29872_;
  assign new_n29874_ = ~pi0188 & ~new_n19370_;
  assign new_n29875_ = ~pi0768 & ~new_n29874_;
  assign new_n29876_ = ~new_n24446_ & new_n29875_;
  assign new_n29877_ = ~new_n29873_ & ~new_n29876_;
  assign new_n29878_ = ~pi0705 & ~new_n29877_;
  assign new_n29879_ = ~pi0188 & new_n19389_;
  assign new_n29880_ = pi0188 & new_n19394_;
  assign new_n29881_ = pi0768 & ~new_n19396_;
  assign new_n29882_ = ~new_n29880_ & new_n29881_;
  assign new_n29883_ = ~new_n29879_ & new_n29882_;
  assign new_n29884_ = pi0188 & new_n19406_;
  assign new_n29885_ = ~pi0188 & ~new_n19414_;
  assign new_n29886_ = ~pi0768 & ~new_n29885_;
  assign new_n29887_ = ~new_n29884_ & new_n29886_;
  assign new_n29888_ = pi0705 & ~new_n29887_;
  assign new_n29889_ = ~new_n29883_ & new_n29888_;
  assign new_n29890_ = new_n3272_ & ~new_n29889_;
  assign new_n29891_ = ~new_n29878_ & new_n29890_;
  assign new_n29892_ = ~new_n29870_ & ~new_n29891_;
  assign new_n29893_ = ~pi0625 & new_n29892_;
  assign new_n29894_ = new_n3272_ & new_n29877_;
  assign new_n29895_ = ~new_n29870_ & ~new_n29894_;
  assign new_n29896_ = pi0625 & new_n29895_;
  assign new_n29897_ = ~pi1153 & ~new_n29896_;
  assign new_n29898_ = ~new_n29893_ & new_n29897_;
  assign new_n29899_ = ~pi0188 & new_n18124_;
  assign new_n29900_ = pi0188 & ~new_n18128_;
  assign new_n29901_ = ~pi0038 & ~new_n29900_;
  assign new_n29902_ = ~new_n29899_ & new_n29901_;
  assign new_n29903_ = ~pi0188 & ~new_n17431_;
  assign new_n29904_ = new_n17544_ & ~new_n29903_;
  assign new_n29905_ = pi0705 & ~new_n29904_;
  assign new_n29906_ = ~new_n29902_ & new_n29905_;
  assign new_n29907_ = ~pi0188 & ~pi0705;
  assign new_n29908_ = ~new_n17551_ & new_n29907_;
  assign new_n29909_ = new_n3272_ & ~new_n29908_;
  assign new_n29910_ = ~new_n29906_ & new_n29909_;
  assign new_n29911_ = ~new_n29870_ & ~new_n29910_;
  assign new_n29912_ = pi0625 & new_n29911_;
  assign new_n29913_ = ~pi0188 & ~new_n17558_;
  assign new_n29914_ = ~pi0625 & new_n29913_;
  assign new_n29915_ = pi1153 & ~new_n29914_;
  assign new_n29916_ = ~new_n29912_ & new_n29915_;
  assign new_n29917_ = ~pi0608 & ~new_n29916_;
  assign new_n29918_ = ~new_n29898_ & new_n29917_;
  assign new_n29919_ = pi0625 & new_n29892_;
  assign new_n29920_ = ~pi0625 & new_n29895_;
  assign new_n29921_ = pi1153 & ~new_n29920_;
  assign new_n29922_ = ~new_n29919_ & new_n29921_;
  assign new_n29923_ = ~pi0625 & new_n29911_;
  assign new_n29924_ = pi0625 & new_n29913_;
  assign new_n29925_ = ~pi1153 & ~new_n29924_;
  assign new_n29926_ = ~new_n29923_ & new_n29925_;
  assign new_n29927_ = pi0608 & ~new_n29926_;
  assign new_n29928_ = ~new_n29922_ & new_n29927_;
  assign new_n29929_ = ~new_n29918_ & ~new_n29928_;
  assign new_n29930_ = pi0778 & ~new_n29929_;
  assign new_n29931_ = ~pi0778 & new_n29892_;
  assign new_n29932_ = ~new_n29930_ & ~new_n29931_;
  assign new_n29933_ = ~pi0609 & ~new_n29932_;
  assign new_n29934_ = ~pi0778 & ~new_n29911_;
  assign new_n29935_ = ~new_n29916_ & ~new_n29926_;
  assign new_n29936_ = pi0778 & ~new_n29935_;
  assign new_n29937_ = ~new_n29934_ & ~new_n29936_;
  assign new_n29938_ = pi0609 & new_n29937_;
  assign new_n29939_ = ~pi1155 & ~new_n29938_;
  assign new_n29940_ = ~new_n29933_ & new_n29939_;
  assign new_n29941_ = ~new_n17591_ & ~new_n29913_;
  assign new_n29942_ = ~new_n17590_ & ~new_n29895_;
  assign new_n29943_ = pi0609 & new_n29942_;
  assign new_n29944_ = ~new_n29941_ & ~new_n29943_;
  assign new_n29945_ = pi1155 & ~new_n29944_;
  assign new_n29946_ = ~pi0660 & ~new_n29945_;
  assign new_n29947_ = ~new_n29940_ & new_n29946_;
  assign new_n29948_ = pi0609 & ~new_n29932_;
  assign new_n29949_ = ~pi0609 & new_n29937_;
  assign new_n29950_ = pi1155 & ~new_n29949_;
  assign new_n29951_ = ~new_n29948_ & new_n29950_;
  assign new_n29952_ = ~new_n17603_ & ~new_n29913_;
  assign new_n29953_ = ~pi0609 & new_n29942_;
  assign new_n29954_ = ~new_n29952_ & ~new_n29953_;
  assign new_n29955_ = ~pi1155 & ~new_n29954_;
  assign new_n29956_ = pi0660 & ~new_n29955_;
  assign new_n29957_ = ~new_n29951_ & new_n29956_;
  assign new_n29958_ = ~new_n29947_ & ~new_n29957_;
  assign new_n29959_ = pi0785 & ~new_n29958_;
  assign new_n29960_ = ~pi0785 & ~new_n29932_;
  assign new_n29961_ = ~new_n29959_ & ~new_n29960_;
  assign new_n29962_ = ~pi0618 & ~new_n29961_;
  assign new_n29963_ = ~new_n17618_ & ~new_n29937_;
  assign new_n29964_ = new_n17618_ & ~new_n29913_;
  assign new_n29965_ = ~new_n29963_ & ~new_n29964_;
  assign new_n29966_ = pi0618 & new_n29965_;
  assign new_n29967_ = ~pi1154 & ~new_n29966_;
  assign new_n29968_ = ~new_n29962_ & new_n29967_;
  assign new_n29969_ = new_n17590_ & ~new_n29913_;
  assign new_n29970_ = ~new_n29942_ & ~new_n29969_;
  assign new_n29971_ = ~pi0785 & ~new_n29970_;
  assign new_n29972_ = ~new_n29945_ & ~new_n29955_;
  assign new_n29973_ = pi0785 & ~new_n29972_;
  assign new_n29974_ = ~new_n29971_ & ~new_n29973_;
  assign new_n29975_ = pi0618 & new_n29974_;
  assign new_n29976_ = ~pi0618 & new_n29913_;
  assign new_n29977_ = pi1154 & ~new_n29976_;
  assign new_n29978_ = ~new_n29975_ & new_n29977_;
  assign new_n29979_ = ~pi0627 & ~new_n29978_;
  assign new_n29980_ = ~new_n29968_ & new_n29979_;
  assign new_n29981_ = pi0618 & ~new_n29961_;
  assign new_n29982_ = ~pi0618 & new_n29965_;
  assign new_n29983_ = pi1154 & ~new_n29982_;
  assign new_n29984_ = ~new_n29981_ & new_n29983_;
  assign new_n29985_ = ~pi0618 & new_n29974_;
  assign new_n29986_ = pi0618 & new_n29913_;
  assign new_n29987_ = ~pi1154 & ~new_n29986_;
  assign new_n29988_ = ~new_n29985_ & new_n29987_;
  assign new_n29989_ = pi0627 & ~new_n29988_;
  assign new_n29990_ = ~new_n29984_ & new_n29989_;
  assign new_n29991_ = ~new_n29980_ & ~new_n29990_;
  assign new_n29992_ = pi0781 & ~new_n29991_;
  assign new_n29993_ = ~pi0781 & ~new_n29961_;
  assign new_n29994_ = ~new_n29992_ & ~new_n29993_;
  assign new_n29995_ = ~pi0619 & ~new_n29994_;
  assign new_n29996_ = ~new_n17655_ & new_n29965_;
  assign new_n29997_ = new_n17655_ & new_n29913_;
  assign new_n29998_ = ~new_n29996_ & ~new_n29997_;
  assign new_n29999_ = pi0619 & ~new_n29998_;
  assign new_n30000_ = ~pi1159 & ~new_n29999_;
  assign new_n30001_ = ~new_n29995_ & new_n30000_;
  assign new_n30002_ = ~pi0781 & ~new_n29974_;
  assign new_n30003_ = ~new_n29978_ & ~new_n29988_;
  assign new_n30004_ = pi0781 & ~new_n30003_;
  assign new_n30005_ = ~new_n30002_ & ~new_n30004_;
  assign new_n30006_ = pi0619 & new_n30005_;
  assign new_n30007_ = ~pi0619 & new_n29913_;
  assign new_n30008_ = pi1159 & ~new_n30007_;
  assign new_n30009_ = ~new_n30006_ & new_n30008_;
  assign new_n30010_ = ~pi0648 & ~new_n30009_;
  assign new_n30011_ = ~new_n30001_ & new_n30010_;
  assign new_n30012_ = pi0619 & ~new_n29994_;
  assign new_n30013_ = ~pi0619 & ~new_n29998_;
  assign new_n30014_ = pi1159 & ~new_n30013_;
  assign new_n30015_ = ~new_n30012_ & new_n30014_;
  assign new_n30016_ = ~pi0619 & new_n30005_;
  assign new_n30017_ = pi0619 & new_n29913_;
  assign new_n30018_ = ~pi1159 & ~new_n30017_;
  assign new_n30019_ = ~new_n30016_ & new_n30018_;
  assign new_n30020_ = pi0648 & ~new_n30019_;
  assign new_n30021_ = ~new_n30015_ & new_n30020_;
  assign new_n30022_ = ~new_n30011_ & ~new_n30021_;
  assign new_n30023_ = pi0789 & ~new_n30022_;
  assign new_n30024_ = ~pi0789 & ~new_n29994_;
  assign new_n30025_ = ~new_n30023_ & ~new_n30024_;
  assign new_n30026_ = ~pi0788 & new_n30025_;
  assign new_n30027_ = ~pi0626 & new_n30025_;
  assign new_n30028_ = new_n17691_ & ~new_n29913_;
  assign new_n30029_ = ~new_n17691_ & new_n29998_;
  assign new_n30030_ = ~new_n30028_ & ~new_n30029_;
  assign new_n30031_ = pi0626 & ~new_n30030_;
  assign new_n30032_ = ~pi0641 & ~new_n30031_;
  assign new_n30033_ = ~new_n30027_ & new_n30032_;
  assign new_n30034_ = ~pi0789 & ~new_n30005_;
  assign new_n30035_ = ~new_n30009_ & ~new_n30019_;
  assign new_n30036_ = pi0789 & ~new_n30035_;
  assign new_n30037_ = ~new_n30034_ & ~new_n30036_;
  assign new_n30038_ = ~pi0626 & ~new_n30037_;
  assign new_n30039_ = pi0626 & ~new_n29913_;
  assign new_n30040_ = pi0641 & ~new_n30039_;
  assign new_n30041_ = ~new_n30038_ & new_n30040_;
  assign new_n30042_ = ~pi1158 & ~new_n30041_;
  assign new_n30043_ = ~new_n30033_ & new_n30042_;
  assign new_n30044_ = pi0626 & new_n30025_;
  assign new_n30045_ = ~pi0626 & ~new_n30030_;
  assign new_n30046_ = pi0641 & ~new_n30045_;
  assign new_n30047_ = ~new_n30044_ & new_n30046_;
  assign new_n30048_ = pi0626 & ~new_n30037_;
  assign new_n30049_ = ~pi0626 & ~new_n29913_;
  assign new_n30050_ = ~pi0641 & ~new_n30049_;
  assign new_n30051_ = ~new_n30048_ & new_n30050_;
  assign new_n30052_ = pi1158 & ~new_n30051_;
  assign new_n30053_ = ~new_n30047_ & new_n30052_;
  assign new_n30054_ = ~new_n30043_ & ~new_n30053_;
  assign new_n30055_ = pi0788 & ~new_n30054_;
  assign new_n30056_ = ~new_n30026_ & ~new_n30055_;
  assign new_n30057_ = ~pi0628 & new_n30056_;
  assign new_n30058_ = ~new_n17968_ & new_n30037_;
  assign new_n30059_ = new_n17968_ & new_n29913_;
  assign new_n30060_ = ~new_n30058_ & ~new_n30059_;
  assign new_n30061_ = pi0628 & ~new_n30060_;
  assign new_n30062_ = ~pi1156 & ~new_n30061_;
  assign new_n30063_ = ~new_n30057_ & new_n30062_;
  assign new_n30064_ = ~new_n17734_ & new_n30030_;
  assign new_n30065_ = new_n17734_ & new_n29913_;
  assign new_n30066_ = ~new_n30064_ & ~new_n30065_;
  assign new_n30067_ = pi0628 & ~new_n30066_;
  assign new_n30068_ = ~pi0628 & new_n29913_;
  assign new_n30069_ = pi1156 & ~new_n30068_;
  assign new_n30070_ = ~new_n30067_ & new_n30069_;
  assign new_n30071_ = ~pi0629 & ~new_n30070_;
  assign new_n30072_ = ~new_n30063_ & new_n30071_;
  assign new_n30073_ = pi0628 & new_n30056_;
  assign new_n30074_ = ~pi0628 & ~new_n30060_;
  assign new_n30075_ = pi1156 & ~new_n30074_;
  assign new_n30076_ = ~new_n30073_ & new_n30075_;
  assign new_n30077_ = ~pi0628 & ~new_n30066_;
  assign new_n30078_ = pi0628 & new_n29913_;
  assign new_n30079_ = ~pi1156 & ~new_n30078_;
  assign new_n30080_ = ~new_n30077_ & new_n30079_;
  assign new_n30081_ = pi0629 & ~new_n30080_;
  assign new_n30082_ = ~new_n30076_ & new_n30081_;
  assign new_n30083_ = ~new_n30072_ & ~new_n30082_;
  assign new_n30084_ = pi0792 & ~new_n30083_;
  assign new_n30085_ = ~pi0792 & new_n30056_;
  assign new_n30086_ = ~new_n30084_ & ~new_n30085_;
  assign new_n30087_ = ~pi0647 & ~new_n30086_;
  assign new_n30088_ = ~new_n17762_ & ~new_n30060_;
  assign new_n30089_ = new_n17762_ & new_n29913_;
  assign new_n30090_ = ~new_n30088_ & ~new_n30089_;
  assign new_n30091_ = pi0647 & ~new_n30090_;
  assign new_n30092_ = ~pi1157 & ~new_n30091_;
  assign new_n30093_ = ~new_n30087_ & new_n30092_;
  assign new_n30094_ = ~pi0792 & new_n30066_;
  assign new_n30095_ = ~new_n30070_ & ~new_n30080_;
  assign new_n30096_ = pi0792 & ~new_n30095_;
  assign new_n30097_ = ~new_n30094_ & ~new_n30096_;
  assign new_n30098_ = pi0647 & new_n30097_;
  assign new_n30099_ = ~pi0647 & new_n29913_;
  assign new_n30100_ = pi1157 & ~new_n30099_;
  assign new_n30101_ = ~new_n30098_ & new_n30100_;
  assign new_n30102_ = ~pi0630 & ~new_n30101_;
  assign new_n30103_ = ~new_n30093_ & new_n30102_;
  assign new_n30104_ = pi0647 & ~new_n30086_;
  assign new_n30105_ = ~pi0647 & ~new_n30090_;
  assign new_n30106_ = pi1157 & ~new_n30105_;
  assign new_n30107_ = ~new_n30104_ & new_n30106_;
  assign new_n30108_ = ~pi0647 & new_n30097_;
  assign new_n30109_ = pi0647 & new_n29913_;
  assign new_n30110_ = ~pi1157 & ~new_n30109_;
  assign new_n30111_ = ~new_n30108_ & new_n30110_;
  assign new_n30112_ = pi0630 & ~new_n30111_;
  assign new_n30113_ = ~new_n30107_ & new_n30112_;
  assign new_n30114_ = ~new_n30103_ & ~new_n30113_;
  assign new_n30115_ = pi0787 & ~new_n30114_;
  assign new_n30116_ = ~pi0787 & ~new_n30086_;
  assign new_n30117_ = ~new_n30115_ & ~new_n30116_;
  assign new_n30118_ = ~pi0644 & ~new_n30117_;
  assign new_n30119_ = ~pi0787 & ~new_n30097_;
  assign new_n30120_ = ~new_n30101_ & ~new_n30111_;
  assign new_n30121_ = pi0787 & ~new_n30120_;
  assign new_n30122_ = ~new_n30119_ & ~new_n30121_;
  assign new_n30123_ = pi0644 & new_n30122_;
  assign new_n30124_ = ~pi0715 & ~new_n30123_;
  assign new_n30125_ = ~new_n30118_ & new_n30124_;
  assign new_n30126_ = new_n17804_ & ~new_n29913_;
  assign new_n30127_ = ~new_n17804_ & new_n30090_;
  assign new_n30128_ = ~new_n30126_ & ~new_n30127_;
  assign new_n30129_ = ~pi0644 & new_n30128_;
  assign new_n30130_ = pi0644 & new_n29913_;
  assign new_n30131_ = pi0715 & ~new_n30130_;
  assign new_n30132_ = ~new_n30129_ & new_n30131_;
  assign new_n30133_ = ~pi1160 & ~new_n30132_;
  assign new_n30134_ = ~new_n30125_ & new_n30133_;
  assign new_n30135_ = pi0644 & ~new_n30117_;
  assign new_n30136_ = ~pi0644 & new_n30122_;
  assign new_n30137_ = pi0715 & ~new_n30136_;
  assign new_n30138_ = ~new_n30135_ & new_n30137_;
  assign new_n30139_ = pi0644 & new_n30128_;
  assign new_n30140_ = ~pi0644 & new_n29913_;
  assign new_n30141_ = ~pi0715 & ~new_n30140_;
  assign new_n30142_ = ~new_n30139_ & new_n30141_;
  assign new_n30143_ = pi1160 & ~new_n30142_;
  assign new_n30144_ = ~new_n30138_ & new_n30143_;
  assign new_n30145_ = pi0790 & ~new_n30144_;
  assign new_n30146_ = ~new_n30134_ & new_n30145_;
  assign new_n30147_ = ~pi0790 & new_n30117_;
  assign new_n30148_ = ~po1038 & ~new_n30147_;
  assign new_n30149_ = ~new_n30146_ & new_n30148_;
  assign new_n30150_ = ~pi0188 & po1038;
  assign new_n30151_ = ~pi0832 & ~new_n30150_;
  assign new_n30152_ = ~new_n30149_ & new_n30151_;
  assign new_n30153_ = ~pi0188 & ~new_n2754_;
  assign new_n30154_ = ~pi0768 & new_n16913_;
  assign new_n30155_ = ~new_n30153_ & ~new_n30154_;
  assign new_n30156_ = ~new_n17858_ & ~new_n30155_;
  assign new_n30157_ = ~pi0785 & ~new_n30156_;
  assign new_n30158_ = ~new_n17863_ & ~new_n30155_;
  assign new_n30159_ = pi1155 & ~new_n30158_;
  assign new_n30160_ = ~new_n17866_ & new_n30156_;
  assign new_n30161_ = ~pi1155 & ~new_n30160_;
  assign new_n30162_ = ~new_n30159_ & ~new_n30161_;
  assign new_n30163_ = pi0785 & ~new_n30162_;
  assign new_n30164_ = ~new_n30157_ & ~new_n30163_;
  assign new_n30165_ = ~pi0781 & ~new_n30164_;
  assign new_n30166_ = ~new_n17873_ & new_n30164_;
  assign new_n30167_ = pi1154 & ~new_n30166_;
  assign new_n30168_ = ~new_n17876_ & new_n30164_;
  assign new_n30169_ = ~pi1154 & ~new_n30168_;
  assign new_n30170_ = ~new_n30167_ & ~new_n30169_;
  assign new_n30171_ = pi0781 & ~new_n30170_;
  assign new_n30172_ = ~new_n30165_ & ~new_n30171_;
  assign new_n30173_ = ~pi0789 & ~new_n30172_;
  assign new_n30174_ = pi0619 & new_n30172_;
  assign new_n30175_ = ~pi0619 & new_n30153_;
  assign new_n30176_ = pi1159 & ~new_n30175_;
  assign new_n30177_ = ~new_n30174_ & new_n30176_;
  assign new_n30178_ = ~pi0619 & new_n30172_;
  assign new_n30179_ = pi0619 & new_n30153_;
  assign new_n30180_ = ~pi1159 & ~new_n30179_;
  assign new_n30181_ = ~new_n30178_ & new_n30180_;
  assign new_n30182_ = ~new_n30177_ & ~new_n30181_;
  assign new_n30183_ = pi0789 & ~new_n30182_;
  assign new_n30184_ = ~new_n30173_ & ~new_n30183_;
  assign new_n30185_ = ~new_n17968_ & new_n30184_;
  assign new_n30186_ = new_n17968_ & new_n30153_;
  assign new_n30187_ = ~new_n30185_ & ~new_n30186_;
  assign new_n30188_ = ~new_n17762_ & ~new_n30187_;
  assign new_n30189_ = new_n17762_ & new_n30153_;
  assign new_n30190_ = ~new_n30188_ & ~new_n30189_;
  assign new_n30191_ = ~new_n20556_ & new_n30190_;
  assign new_n30192_ = pi0705 & new_n16915_;
  assign new_n30193_ = ~new_n30153_ & ~new_n30192_;
  assign new_n30194_ = ~pi0778 & new_n30193_;
  assign new_n30195_ = ~pi0625 & new_n30192_;
  assign new_n30196_ = ~new_n30193_ & ~new_n30195_;
  assign new_n30197_ = pi1153 & ~new_n30196_;
  assign new_n30198_ = ~pi1153 & ~new_n30153_;
  assign new_n30199_ = ~new_n30195_ & new_n30198_;
  assign new_n30200_ = ~new_n30197_ & ~new_n30199_;
  assign new_n30201_ = pi0778 & ~new_n30200_;
  assign new_n30202_ = ~new_n30194_ & ~new_n30201_;
  assign new_n30203_ = ~new_n17844_ & new_n30202_;
  assign new_n30204_ = ~new_n17846_ & new_n30203_;
  assign new_n30205_ = ~new_n17848_ & new_n30204_;
  assign new_n30206_ = ~new_n17980_ & new_n30205_;
  assign new_n30207_ = ~new_n18011_ & new_n30206_;
  assign new_n30208_ = ~pi0647 & new_n30207_;
  assign new_n30209_ = pi0647 & new_n30153_;
  assign new_n30210_ = ~pi1157 & ~new_n30209_;
  assign new_n30211_ = ~new_n30208_ & new_n30210_;
  assign new_n30212_ = pi0630 & new_n30211_;
  assign new_n30213_ = pi0647 & ~new_n30207_;
  assign new_n30214_ = ~pi0647 & ~new_n30153_;
  assign new_n30215_ = ~new_n30213_ & ~new_n30214_;
  assign new_n30216_ = new_n17801_ & ~new_n30215_;
  assign new_n30217_ = ~new_n30212_ & ~new_n30216_;
  assign new_n30218_ = ~new_n30191_ & new_n30217_;
  assign new_n30219_ = pi0787 & ~new_n30218_;
  assign new_n30220_ = pi0626 & ~new_n30184_;
  assign new_n30221_ = ~pi0626 & ~new_n30153_;
  assign new_n30222_ = new_n17731_ & ~new_n30221_;
  assign new_n30223_ = ~new_n30220_ & new_n30222_;
  assign new_n30224_ = new_n17856_ & new_n30205_;
  assign new_n30225_ = ~pi0626 & ~new_n30184_;
  assign new_n30226_ = pi0626 & ~new_n30153_;
  assign new_n30227_ = new_n17732_ & ~new_n30226_;
  assign new_n30228_ = ~new_n30225_ & new_n30227_;
  assign new_n30229_ = ~new_n30224_ & ~new_n30228_;
  assign new_n30230_ = ~new_n30223_ & new_n30229_;
  assign new_n30231_ = pi0788 & ~new_n30230_;
  assign new_n30232_ = ~new_n16639_ & ~new_n30193_;
  assign new_n30233_ = pi0625 & new_n30232_;
  assign new_n30234_ = new_n30155_ & ~new_n30232_;
  assign new_n30235_ = ~new_n30233_ & ~new_n30234_;
  assign new_n30236_ = new_n30198_ & ~new_n30235_;
  assign new_n30237_ = ~pi0608 & ~new_n30197_;
  assign new_n30238_ = ~new_n30236_ & new_n30237_;
  assign new_n30239_ = pi1153 & new_n30155_;
  assign new_n30240_ = ~new_n30233_ & new_n30239_;
  assign new_n30241_ = pi0608 & ~new_n30199_;
  assign new_n30242_ = ~new_n30240_ & new_n30241_;
  assign new_n30243_ = ~new_n30238_ & ~new_n30242_;
  assign new_n30244_ = pi0778 & ~new_n30243_;
  assign new_n30245_ = ~pi0778 & ~new_n30234_;
  assign new_n30246_ = ~new_n30244_ & ~new_n30245_;
  assign new_n30247_ = ~pi0609 & ~new_n30246_;
  assign new_n30248_ = pi0609 & new_n30202_;
  assign new_n30249_ = ~pi1155 & ~new_n30248_;
  assign new_n30250_ = ~new_n30247_ & new_n30249_;
  assign new_n30251_ = ~pi0660 & ~new_n30159_;
  assign new_n30252_ = ~new_n30250_ & new_n30251_;
  assign new_n30253_ = pi0609 & ~new_n30246_;
  assign new_n30254_ = ~pi0609 & new_n30202_;
  assign new_n30255_ = pi1155 & ~new_n30254_;
  assign new_n30256_ = ~new_n30253_ & new_n30255_;
  assign new_n30257_ = pi0660 & ~new_n30161_;
  assign new_n30258_ = ~new_n30256_ & new_n30257_;
  assign new_n30259_ = ~new_n30252_ & ~new_n30258_;
  assign new_n30260_ = pi0785 & ~new_n30259_;
  assign new_n30261_ = ~pi0785 & ~new_n30246_;
  assign new_n30262_ = ~new_n30260_ & ~new_n30261_;
  assign new_n30263_ = ~pi0618 & ~new_n30262_;
  assign new_n30264_ = pi0618 & new_n30203_;
  assign new_n30265_ = ~pi1154 & ~new_n30264_;
  assign new_n30266_ = ~new_n30263_ & new_n30265_;
  assign new_n30267_ = ~pi0627 & ~new_n30167_;
  assign new_n30268_ = ~new_n30266_ & new_n30267_;
  assign new_n30269_ = pi0618 & ~new_n30262_;
  assign new_n30270_ = ~pi0618 & new_n30203_;
  assign new_n30271_ = pi1154 & ~new_n30270_;
  assign new_n30272_ = ~new_n30269_ & new_n30271_;
  assign new_n30273_ = pi0627 & ~new_n30169_;
  assign new_n30274_ = ~new_n30272_ & new_n30273_;
  assign new_n30275_ = ~new_n30268_ & ~new_n30274_;
  assign new_n30276_ = pi0781 & ~new_n30275_;
  assign new_n30277_ = ~pi0781 & ~new_n30262_;
  assign new_n30278_ = ~new_n30276_ & ~new_n30277_;
  assign new_n30279_ = pi0619 & ~new_n30278_;
  assign new_n30280_ = ~pi0619 & new_n30204_;
  assign new_n30281_ = pi1159 & ~new_n30280_;
  assign new_n30282_ = ~new_n30279_ & new_n30281_;
  assign new_n30283_ = pi0648 & ~new_n30181_;
  assign new_n30284_ = ~new_n30282_ & new_n30283_;
  assign new_n30285_ = ~pi0619 & ~new_n30278_;
  assign new_n30286_ = pi0619 & new_n30204_;
  assign new_n30287_ = ~pi1159 & ~new_n30286_;
  assign new_n30288_ = ~new_n30285_ & new_n30287_;
  assign new_n30289_ = ~pi0648 & ~new_n30177_;
  assign new_n30290_ = ~new_n30288_ & new_n30289_;
  assign new_n30291_ = pi0789 & ~new_n30290_;
  assign new_n30292_ = ~new_n30284_ & new_n30291_;
  assign new_n30293_ = ~pi0789 & new_n30278_;
  assign new_n30294_ = new_n17969_ & ~new_n30293_;
  assign new_n30295_ = ~new_n30292_ & new_n30294_;
  assign new_n30296_ = ~new_n30231_ & ~new_n30295_;
  assign new_n30297_ = ~new_n20364_ & ~new_n30296_;
  assign new_n30298_ = new_n18008_ & ~new_n30187_;
  assign new_n30299_ = new_n20851_ & new_n30206_;
  assign new_n30300_ = ~new_n30298_ & ~new_n30299_;
  assign new_n30301_ = ~pi0629 & ~new_n30300_;
  assign new_n30302_ = new_n20855_ & new_n30206_;
  assign new_n30303_ = new_n18007_ & ~new_n30187_;
  assign new_n30304_ = ~new_n30302_ & ~new_n30303_;
  assign new_n30305_ = pi0629 & ~new_n30304_;
  assign new_n30306_ = ~new_n30301_ & ~new_n30305_;
  assign new_n30307_ = pi0792 & ~new_n30306_;
  assign new_n30308_ = ~new_n20360_ & ~new_n30307_;
  assign new_n30309_ = ~new_n30297_ & new_n30308_;
  assign new_n30310_ = ~new_n30219_ & ~new_n30309_;
  assign new_n30311_ = pi0644 & new_n30310_;
  assign new_n30312_ = ~pi0787 & ~new_n30207_;
  assign new_n30313_ = pi1157 & ~new_n30215_;
  assign new_n30314_ = ~new_n30211_ & ~new_n30313_;
  assign new_n30315_ = pi0787 & ~new_n30314_;
  assign new_n30316_ = ~new_n30312_ & ~new_n30315_;
  assign new_n30317_ = ~pi0644 & new_n30316_;
  assign new_n30318_ = pi0715 & ~new_n30317_;
  assign new_n30319_ = ~new_n30311_ & new_n30318_;
  assign new_n30320_ = ~new_n17804_ & ~new_n30190_;
  assign new_n30321_ = new_n17804_ & new_n30153_;
  assign new_n30322_ = ~new_n30320_ & ~new_n30321_;
  assign new_n30323_ = pi0644 & ~new_n30322_;
  assign new_n30324_ = ~pi0644 & new_n30153_;
  assign new_n30325_ = ~pi0715 & ~new_n30324_;
  assign new_n30326_ = ~new_n30323_ & new_n30325_;
  assign new_n30327_ = pi1160 & ~new_n30326_;
  assign new_n30328_ = ~new_n30319_ & new_n30327_;
  assign new_n30329_ = ~pi0644 & new_n30310_;
  assign new_n30330_ = pi0644 & new_n30316_;
  assign new_n30331_ = ~pi0715 & ~new_n30330_;
  assign new_n30332_ = ~new_n30329_ & new_n30331_;
  assign new_n30333_ = ~pi0644 & ~new_n30322_;
  assign new_n30334_ = pi0644 & new_n30153_;
  assign new_n30335_ = pi0715 & ~new_n30334_;
  assign new_n30336_ = ~new_n30333_ & new_n30335_;
  assign new_n30337_ = ~pi1160 & ~new_n30336_;
  assign new_n30338_ = ~new_n30332_ & new_n30337_;
  assign new_n30339_ = ~new_n30328_ & ~new_n30338_;
  assign new_n30340_ = pi0790 & ~new_n30339_;
  assign new_n30341_ = ~pi0790 & new_n30310_;
  assign new_n30342_ = pi0832 & ~new_n30341_;
  assign new_n30343_ = ~new_n30340_ & new_n30342_;
  assign po0345 = ~new_n30152_ & ~new_n30343_;
  assign new_n30345_ = pi0189 & ~new_n3272_;
  assign new_n30346_ = pi0772 & new_n17391_;
  assign new_n30347_ = ~new_n22231_ & ~new_n30346_;
  assign new_n30348_ = pi0039 & ~new_n30347_;
  assign new_n30349_ = pi0772 & new_n17226_;
  assign new_n30350_ = ~pi0772 & new_n17260_;
  assign new_n30351_ = ~pi0039 & ~new_n30350_;
  assign new_n30352_ = ~new_n30349_ & new_n30351_;
  assign new_n30353_ = ~new_n30348_ & ~new_n30352_;
  assign new_n30354_ = pi0189 & ~new_n30353_;
  assign new_n30355_ = ~pi0189 & pi0772;
  assign new_n30356_ = new_n17426_ & new_n30355_;
  assign new_n30357_ = ~new_n30354_ & ~new_n30356_;
  assign new_n30358_ = ~pi0038 & ~new_n30357_;
  assign new_n30359_ = pi0772 & new_n16639_;
  assign new_n30360_ = new_n17431_ & ~new_n30359_;
  assign new_n30361_ = ~pi0189 & ~new_n17431_;
  assign new_n30362_ = pi0038 & ~new_n30361_;
  assign new_n30363_ = ~new_n30360_ & new_n30362_;
  assign new_n30364_ = ~new_n30358_ & ~new_n30363_;
  assign new_n30365_ = ~pi0727 & new_n30364_;
  assign new_n30366_ = pi0189 & ~new_n16810_;
  assign new_n30367_ = ~pi0189 & ~new_n16928_;
  assign new_n30368_ = ~pi0772 & ~new_n30367_;
  assign new_n30369_ = ~new_n30366_ & new_n30368_;
  assign new_n30370_ = ~pi0189 & ~new_n17007_;
  assign new_n30371_ = pi0189 & new_n17074_;
  assign new_n30372_ = pi0772 & ~new_n30371_;
  assign new_n30373_ = ~new_n30370_ & new_n30372_;
  assign new_n30374_ = pi0039 & ~new_n30373_;
  assign new_n30375_ = ~new_n30369_ & new_n30374_;
  assign new_n30376_ = pi0189 & ~new_n17217_;
  assign new_n30377_ = ~pi0189 & ~new_n17178_;
  assign new_n30378_ = ~pi0772 & ~new_n30377_;
  assign new_n30379_ = ~new_n30376_ & new_n30378_;
  assign new_n30380_ = pi0189 & new_n17227_;
  assign new_n30381_ = ~pi0189 & new_n17234_;
  assign new_n30382_ = pi0772 & ~new_n30381_;
  assign new_n30383_ = ~new_n30380_ & new_n30382_;
  assign new_n30384_ = ~pi0039 & ~new_n30383_;
  assign new_n30385_ = ~new_n30379_ & new_n30384_;
  assign new_n30386_ = ~pi0038 & ~new_n30385_;
  assign new_n30387_ = ~new_n30375_ & new_n30386_;
  assign new_n30388_ = pi0727 & ~new_n19396_;
  assign new_n30389_ = ~new_n30363_ & new_n30388_;
  assign new_n30390_ = ~new_n30387_ & new_n30389_;
  assign new_n30391_ = new_n3272_ & ~new_n30390_;
  assign new_n30392_ = ~new_n30365_ & new_n30391_;
  assign new_n30393_ = ~new_n30345_ & ~new_n30392_;
  assign new_n30394_ = ~pi0625 & new_n30393_;
  assign new_n30395_ = new_n3272_ & ~new_n30364_;
  assign new_n30396_ = ~new_n30345_ & ~new_n30395_;
  assign new_n30397_ = pi0625 & new_n30396_;
  assign new_n30398_ = ~pi1153 & ~new_n30397_;
  assign new_n30399_ = ~new_n30394_ & new_n30398_;
  assign new_n30400_ = pi0189 & ~new_n17558_;
  assign new_n30401_ = pi0727 & new_n3272_;
  assign new_n30402_ = ~new_n30400_ & ~new_n30401_;
  assign new_n30403_ = pi0189 & ~new_n18124_;
  assign new_n30404_ = ~pi0189 & new_n18128_;
  assign new_n30405_ = ~pi0038 & ~new_n30404_;
  assign new_n30406_ = ~new_n30403_ & new_n30405_;
  assign new_n30407_ = new_n19956_ & ~new_n30361_;
  assign new_n30408_ = new_n30401_ & ~new_n30407_;
  assign new_n30409_ = ~new_n30406_ & new_n30408_;
  assign new_n30410_ = ~new_n30402_ & ~new_n30409_;
  assign new_n30411_ = pi0625 & ~new_n30410_;
  assign new_n30412_ = ~pi0625 & ~new_n30400_;
  assign new_n30413_ = pi1153 & ~new_n30412_;
  assign new_n30414_ = ~new_n30411_ & new_n30413_;
  assign new_n30415_ = ~pi0608 & ~new_n30414_;
  assign new_n30416_ = ~new_n30399_ & new_n30415_;
  assign new_n30417_ = pi0625 & new_n30393_;
  assign new_n30418_ = ~pi0625 & new_n30396_;
  assign new_n30419_ = pi1153 & ~new_n30418_;
  assign new_n30420_ = ~new_n30417_ & new_n30419_;
  assign new_n30421_ = ~pi0625 & ~new_n30410_;
  assign new_n30422_ = pi0625 & ~new_n30400_;
  assign new_n30423_ = ~pi1153 & ~new_n30422_;
  assign new_n30424_ = ~new_n30421_ & new_n30423_;
  assign new_n30425_ = pi0608 & ~new_n30424_;
  assign new_n30426_ = ~new_n30420_ & new_n30425_;
  assign new_n30427_ = ~new_n30416_ & ~new_n30426_;
  assign new_n30428_ = pi0778 & ~new_n30427_;
  assign new_n30429_ = ~pi0778 & new_n30393_;
  assign new_n30430_ = ~new_n30428_ & ~new_n30429_;
  assign new_n30431_ = ~pi0609 & ~new_n30430_;
  assign new_n30432_ = ~pi0778 & new_n30410_;
  assign new_n30433_ = ~new_n30414_ & ~new_n30424_;
  assign new_n30434_ = pi0778 & ~new_n30433_;
  assign new_n30435_ = ~new_n30432_ & ~new_n30434_;
  assign new_n30436_ = pi0609 & new_n30435_;
  assign new_n30437_ = ~pi1155 & ~new_n30436_;
  assign new_n30438_ = ~new_n30431_ & new_n30437_;
  assign new_n30439_ = new_n17590_ & ~new_n30400_;
  assign new_n30440_ = ~new_n17590_ & new_n30396_;
  assign new_n30441_ = ~new_n30439_ & ~new_n30440_;
  assign new_n30442_ = pi0609 & ~new_n30441_;
  assign new_n30443_ = ~pi0609 & ~new_n30400_;
  assign new_n30444_ = pi1155 & ~new_n30443_;
  assign new_n30445_ = ~new_n30442_ & new_n30444_;
  assign new_n30446_ = ~pi0660 & ~new_n30445_;
  assign new_n30447_ = ~new_n30438_ & new_n30446_;
  assign new_n30448_ = pi0609 & ~new_n30430_;
  assign new_n30449_ = ~pi0609 & new_n30435_;
  assign new_n30450_ = pi1155 & ~new_n30449_;
  assign new_n30451_ = ~new_n30448_ & new_n30450_;
  assign new_n30452_ = ~pi0609 & ~new_n30441_;
  assign new_n30453_ = pi0609 & ~new_n30400_;
  assign new_n30454_ = ~pi1155 & ~new_n30453_;
  assign new_n30455_ = ~new_n30452_ & new_n30454_;
  assign new_n30456_ = pi0660 & ~new_n30455_;
  assign new_n30457_ = ~new_n30451_ & new_n30456_;
  assign new_n30458_ = ~new_n30447_ & ~new_n30457_;
  assign new_n30459_ = pi0785 & ~new_n30458_;
  assign new_n30460_ = ~pi0785 & ~new_n30430_;
  assign new_n30461_ = ~new_n30459_ & ~new_n30460_;
  assign new_n30462_ = ~pi0618 & ~new_n30461_;
  assign new_n30463_ = new_n17618_ & ~new_n30400_;
  assign new_n30464_ = ~new_n17618_ & new_n30435_;
  assign new_n30465_ = ~new_n30463_ & ~new_n30464_;
  assign new_n30466_ = pi0618 & ~new_n30465_;
  assign new_n30467_ = ~pi1154 & ~new_n30466_;
  assign new_n30468_ = ~new_n30462_ & new_n30467_;
  assign new_n30469_ = ~pi0785 & new_n30441_;
  assign new_n30470_ = ~new_n30445_ & ~new_n30455_;
  assign new_n30471_ = pi0785 & ~new_n30470_;
  assign new_n30472_ = ~new_n30469_ & ~new_n30471_;
  assign new_n30473_ = pi0618 & new_n30472_;
  assign new_n30474_ = ~pi0618 & ~new_n30400_;
  assign new_n30475_ = pi1154 & ~new_n30474_;
  assign new_n30476_ = ~new_n30473_ & new_n30475_;
  assign new_n30477_ = ~pi0627 & ~new_n30476_;
  assign new_n30478_ = ~new_n30468_ & new_n30477_;
  assign new_n30479_ = pi0618 & ~new_n30461_;
  assign new_n30480_ = ~pi0618 & ~new_n30465_;
  assign new_n30481_ = pi1154 & ~new_n30480_;
  assign new_n30482_ = ~new_n30479_ & new_n30481_;
  assign new_n30483_ = ~pi0618 & new_n30472_;
  assign new_n30484_ = pi0618 & ~new_n30400_;
  assign new_n30485_ = ~pi1154 & ~new_n30484_;
  assign new_n30486_ = ~new_n30483_ & new_n30485_;
  assign new_n30487_ = pi0627 & ~new_n30486_;
  assign new_n30488_ = ~new_n30482_ & new_n30487_;
  assign new_n30489_ = ~new_n30478_ & ~new_n30488_;
  assign new_n30490_ = pi0781 & ~new_n30489_;
  assign new_n30491_ = ~pi0781 & ~new_n30461_;
  assign new_n30492_ = ~new_n30490_ & ~new_n30491_;
  assign new_n30493_ = ~pi0619 & ~new_n30492_;
  assign new_n30494_ = ~new_n17655_ & new_n30465_;
  assign new_n30495_ = new_n17655_ & new_n30400_;
  assign new_n30496_ = ~new_n30494_ & ~new_n30495_;
  assign new_n30497_ = pi0619 & new_n30496_;
  assign new_n30498_ = ~pi1159 & ~new_n30497_;
  assign new_n30499_ = ~new_n30493_ & new_n30498_;
  assign new_n30500_ = ~pi0781 & ~new_n30472_;
  assign new_n30501_ = ~new_n30476_ & ~new_n30486_;
  assign new_n30502_ = pi0781 & ~new_n30501_;
  assign new_n30503_ = ~new_n30500_ & ~new_n30502_;
  assign new_n30504_ = pi0619 & new_n30503_;
  assign new_n30505_ = ~pi0619 & ~new_n30400_;
  assign new_n30506_ = pi1159 & ~new_n30505_;
  assign new_n30507_ = ~new_n30504_ & new_n30506_;
  assign new_n30508_ = ~pi0648 & ~new_n30507_;
  assign new_n30509_ = ~new_n30499_ & new_n30508_;
  assign new_n30510_ = pi0619 & ~new_n30492_;
  assign new_n30511_ = ~pi0619 & new_n30496_;
  assign new_n30512_ = pi1159 & ~new_n30511_;
  assign new_n30513_ = ~new_n30510_ & new_n30512_;
  assign new_n30514_ = ~pi0619 & new_n30503_;
  assign new_n30515_ = pi0619 & ~new_n30400_;
  assign new_n30516_ = ~pi1159 & ~new_n30515_;
  assign new_n30517_ = ~new_n30514_ & new_n30516_;
  assign new_n30518_ = pi0648 & ~new_n30517_;
  assign new_n30519_ = ~new_n30513_ & new_n30518_;
  assign new_n30520_ = ~new_n30509_ & ~new_n30519_;
  assign new_n30521_ = pi0789 & ~new_n30520_;
  assign new_n30522_ = ~pi0789 & ~new_n30492_;
  assign new_n30523_ = ~new_n30521_ & ~new_n30522_;
  assign new_n30524_ = ~pi0788 & new_n30523_;
  assign new_n30525_ = ~pi0626 & new_n30523_;
  assign new_n30526_ = new_n17691_ & ~new_n30400_;
  assign new_n30527_ = ~new_n17691_ & new_n30496_;
  assign new_n30528_ = ~new_n30526_ & ~new_n30527_;
  assign new_n30529_ = pi0626 & new_n30528_;
  assign new_n30530_ = ~pi0641 & ~new_n30529_;
  assign new_n30531_ = ~new_n30525_ & new_n30530_;
  assign new_n30532_ = ~pi0789 & ~new_n30503_;
  assign new_n30533_ = ~new_n30507_ & ~new_n30517_;
  assign new_n30534_ = pi0789 & ~new_n30533_;
  assign new_n30535_ = ~new_n30532_ & ~new_n30534_;
  assign new_n30536_ = ~pi0626 & ~new_n30535_;
  assign new_n30537_ = pi0626 & new_n30400_;
  assign new_n30538_ = pi0641 & ~new_n30537_;
  assign new_n30539_ = ~new_n30536_ & new_n30538_;
  assign new_n30540_ = ~pi1158 & ~new_n30539_;
  assign new_n30541_ = ~new_n30531_ & new_n30540_;
  assign new_n30542_ = pi0626 & new_n30523_;
  assign new_n30543_ = ~pi0626 & new_n30528_;
  assign new_n30544_ = pi0641 & ~new_n30543_;
  assign new_n30545_ = ~new_n30542_ & new_n30544_;
  assign new_n30546_ = pi0626 & ~new_n30535_;
  assign new_n30547_ = ~pi0626 & new_n30400_;
  assign new_n30548_ = ~pi0641 & ~new_n30547_;
  assign new_n30549_ = ~new_n30546_ & new_n30548_;
  assign new_n30550_ = pi1158 & ~new_n30549_;
  assign new_n30551_ = ~new_n30545_ & new_n30550_;
  assign new_n30552_ = ~new_n30541_ & ~new_n30551_;
  assign new_n30553_ = pi0788 & ~new_n30552_;
  assign new_n30554_ = ~new_n30524_ & ~new_n30553_;
  assign new_n30555_ = ~pi0628 & new_n30554_;
  assign new_n30556_ = ~new_n17968_ & ~new_n30535_;
  assign new_n30557_ = new_n17968_ & new_n30400_;
  assign new_n30558_ = ~new_n30556_ & ~new_n30557_;
  assign new_n30559_ = pi0628 & new_n30558_;
  assign new_n30560_ = ~pi1156 & ~new_n30559_;
  assign new_n30561_ = ~new_n30555_ & new_n30560_;
  assign new_n30562_ = ~new_n17734_ & new_n30528_;
  assign new_n30563_ = new_n17734_ & new_n30400_;
  assign new_n30564_ = ~new_n30562_ & ~new_n30563_;
  assign new_n30565_ = pi0628 & new_n30564_;
  assign new_n30566_ = ~pi0628 & ~new_n30400_;
  assign new_n30567_ = pi1156 & ~new_n30566_;
  assign new_n30568_ = ~new_n30565_ & new_n30567_;
  assign new_n30569_ = ~pi0629 & ~new_n30568_;
  assign new_n30570_ = ~new_n30561_ & new_n30569_;
  assign new_n30571_ = pi0628 & new_n30554_;
  assign new_n30572_ = ~pi0628 & new_n30558_;
  assign new_n30573_ = pi1156 & ~new_n30572_;
  assign new_n30574_ = ~new_n30571_ & new_n30573_;
  assign new_n30575_ = ~pi0628 & new_n30564_;
  assign new_n30576_ = pi0628 & ~new_n30400_;
  assign new_n30577_ = ~pi1156 & ~new_n30576_;
  assign new_n30578_ = ~new_n30575_ & new_n30577_;
  assign new_n30579_ = pi0629 & ~new_n30578_;
  assign new_n30580_ = ~new_n30574_ & new_n30579_;
  assign new_n30581_ = ~new_n30570_ & ~new_n30580_;
  assign new_n30582_ = pi0792 & ~new_n30581_;
  assign new_n30583_ = ~pi0792 & new_n30554_;
  assign new_n30584_ = ~new_n30582_ & ~new_n30583_;
  assign new_n30585_ = ~pi0647 & ~new_n30584_;
  assign new_n30586_ = ~new_n17762_ & ~new_n30558_;
  assign new_n30587_ = new_n17762_ & new_n30400_;
  assign new_n30588_ = ~new_n30586_ & ~new_n30587_;
  assign new_n30589_ = pi0647 & new_n30588_;
  assign new_n30590_ = ~pi1157 & ~new_n30589_;
  assign new_n30591_ = ~new_n30585_ & new_n30590_;
  assign new_n30592_ = ~pi0792 & ~new_n30564_;
  assign new_n30593_ = ~new_n30568_ & ~new_n30578_;
  assign new_n30594_ = pi0792 & ~new_n30593_;
  assign new_n30595_ = ~new_n30592_ & ~new_n30594_;
  assign new_n30596_ = pi0647 & new_n30595_;
  assign new_n30597_ = ~pi0647 & ~new_n30400_;
  assign new_n30598_ = pi1157 & ~new_n30597_;
  assign new_n30599_ = ~new_n30596_ & new_n30598_;
  assign new_n30600_ = ~pi0630 & ~new_n30599_;
  assign new_n30601_ = ~new_n30591_ & new_n30600_;
  assign new_n30602_ = pi0647 & ~new_n30584_;
  assign new_n30603_ = ~pi0647 & new_n30588_;
  assign new_n30604_ = pi1157 & ~new_n30603_;
  assign new_n30605_ = ~new_n30602_ & new_n30604_;
  assign new_n30606_ = ~pi0647 & new_n30595_;
  assign new_n30607_ = pi0647 & ~new_n30400_;
  assign new_n30608_ = ~pi1157 & ~new_n30607_;
  assign new_n30609_ = ~new_n30606_ & new_n30608_;
  assign new_n30610_ = pi0630 & ~new_n30609_;
  assign new_n30611_ = ~new_n30605_ & new_n30610_;
  assign new_n30612_ = ~new_n30601_ & ~new_n30611_;
  assign new_n30613_ = pi0787 & ~new_n30612_;
  assign new_n30614_ = ~pi0787 & ~new_n30584_;
  assign new_n30615_ = ~new_n30613_ & ~new_n30614_;
  assign new_n30616_ = ~pi0644 & ~new_n30615_;
  assign new_n30617_ = ~pi0787 & ~new_n30595_;
  assign new_n30618_ = ~new_n30599_ & ~new_n30609_;
  assign new_n30619_ = pi0787 & ~new_n30618_;
  assign new_n30620_ = ~new_n30617_ & ~new_n30619_;
  assign new_n30621_ = pi0644 & new_n30620_;
  assign new_n30622_ = ~pi0715 & ~new_n30621_;
  assign new_n30623_ = ~new_n30616_ & new_n30622_;
  assign new_n30624_ = new_n17804_ & ~new_n30400_;
  assign new_n30625_ = ~new_n17804_ & new_n30588_;
  assign new_n30626_ = ~new_n30624_ & ~new_n30625_;
  assign new_n30627_ = ~pi0644 & ~new_n30626_;
  assign new_n30628_ = pi0644 & ~new_n30400_;
  assign new_n30629_ = pi0715 & ~new_n30628_;
  assign new_n30630_ = ~new_n30627_ & new_n30629_;
  assign new_n30631_ = ~pi1160 & ~new_n30630_;
  assign new_n30632_ = ~new_n30623_ & new_n30631_;
  assign new_n30633_ = pi0644 & ~new_n30615_;
  assign new_n30634_ = ~pi0644 & new_n30620_;
  assign new_n30635_ = pi0715 & ~new_n30634_;
  assign new_n30636_ = ~new_n30633_ & new_n30635_;
  assign new_n30637_ = pi0644 & ~new_n30626_;
  assign new_n30638_ = ~pi0644 & ~new_n30400_;
  assign new_n30639_ = ~pi0715 & ~new_n30638_;
  assign new_n30640_ = ~new_n30637_ & new_n30639_;
  assign new_n30641_ = pi1160 & ~new_n30640_;
  assign new_n30642_ = ~new_n30636_ & new_n30641_;
  assign new_n30643_ = pi0790 & ~new_n30642_;
  assign new_n30644_ = ~new_n30632_ & new_n30643_;
  assign new_n30645_ = ~pi0790 & new_n30615_;
  assign new_n30646_ = new_n6305_ & ~new_n30645_;
  assign new_n30647_ = ~new_n30644_ & new_n30646_;
  assign new_n30648_ = ~pi0189 & ~new_n6305_;
  assign new_n30649_ = ~pi0057 & ~new_n30648_;
  assign new_n30650_ = ~new_n30647_ & new_n30649_;
  assign new_n30651_ = pi0057 & pi0189;
  assign new_n30652_ = ~pi0832 & ~new_n30651_;
  assign new_n30653_ = ~new_n30650_ & new_n30652_;
  assign new_n30654_ = pi0189 & ~new_n2754_;
  assign new_n30655_ = pi0772 & new_n16913_;
  assign new_n30656_ = ~new_n30654_ & ~new_n30655_;
  assign new_n30657_ = pi0727 & new_n16916_;
  assign new_n30658_ = new_n30656_ & ~new_n30657_;
  assign new_n30659_ = pi0625 & new_n30657_;
  assign new_n30660_ = ~new_n30658_ & ~new_n30659_;
  assign new_n30661_ = ~pi1153 & ~new_n30660_;
  assign new_n30662_ = pi0727 & new_n16915_;
  assign new_n30663_ = pi0625 & new_n30662_;
  assign new_n30664_ = pi1153 & ~new_n30654_;
  assign new_n30665_ = ~new_n30663_ & new_n30664_;
  assign new_n30666_ = ~pi0608 & ~new_n30665_;
  assign new_n30667_ = ~new_n30661_ & new_n30666_;
  assign new_n30668_ = pi1153 & new_n30656_;
  assign new_n30669_ = ~new_n30659_ & new_n30668_;
  assign new_n30670_ = ~new_n30654_ & ~new_n30662_;
  assign new_n30671_ = ~new_n30663_ & ~new_n30670_;
  assign new_n30672_ = ~pi1153 & ~new_n30671_;
  assign new_n30673_ = pi0608 & ~new_n30672_;
  assign new_n30674_ = ~new_n30669_ & new_n30673_;
  assign new_n30675_ = ~new_n30667_ & ~new_n30674_;
  assign new_n30676_ = pi0778 & ~new_n30675_;
  assign new_n30677_ = ~pi0778 & ~new_n30658_;
  assign new_n30678_ = ~new_n30676_ & ~new_n30677_;
  assign new_n30679_ = ~pi0609 & ~new_n30678_;
  assign new_n30680_ = ~pi0778 & new_n30670_;
  assign new_n30681_ = ~new_n30665_ & ~new_n30672_;
  assign new_n30682_ = pi0778 & ~new_n30681_;
  assign new_n30683_ = ~new_n30680_ & ~new_n30682_;
  assign new_n30684_ = pi0609 & new_n30683_;
  assign new_n30685_ = ~pi1155 & ~new_n30684_;
  assign new_n30686_ = ~new_n30679_ & new_n30685_;
  assign new_n30687_ = new_n17591_ & new_n30655_;
  assign new_n30688_ = pi1155 & ~new_n30654_;
  assign new_n30689_ = ~new_n30687_ & new_n30688_;
  assign new_n30690_ = ~pi0660 & ~new_n30689_;
  assign new_n30691_ = ~new_n30686_ & new_n30690_;
  assign new_n30692_ = pi0609 & ~new_n30678_;
  assign new_n30693_ = ~pi0609 & new_n30683_;
  assign new_n30694_ = pi1155 & ~new_n30693_;
  assign new_n30695_ = ~new_n30692_ & new_n30694_;
  assign new_n30696_ = new_n17603_ & new_n30655_;
  assign new_n30697_ = ~pi1155 & ~new_n30654_;
  assign new_n30698_ = ~new_n30696_ & new_n30697_;
  assign new_n30699_ = pi0660 & ~new_n30698_;
  assign new_n30700_ = ~new_n30695_ & new_n30699_;
  assign new_n30701_ = ~new_n30691_ & ~new_n30700_;
  assign new_n30702_ = pi0785 & ~new_n30701_;
  assign new_n30703_ = ~pi0785 & ~new_n30678_;
  assign new_n30704_ = ~new_n30702_ & ~new_n30703_;
  assign new_n30705_ = pi0618 & ~new_n30704_;
  assign new_n30706_ = ~new_n17618_ & new_n30683_;
  assign new_n30707_ = ~new_n30654_ & ~new_n30706_;
  assign new_n30708_ = ~pi0618 & ~new_n30707_;
  assign new_n30709_ = pi1154 & ~new_n30708_;
  assign new_n30710_ = ~new_n30705_ & new_n30709_;
  assign new_n30711_ = ~new_n20223_ & new_n30655_;
  assign new_n30712_ = new_n20321_ & new_n30711_;
  assign new_n30713_ = ~pi1154 & ~new_n30654_;
  assign new_n30714_ = ~new_n30712_ & new_n30713_;
  assign new_n30715_ = pi0627 & ~new_n30714_;
  assign new_n30716_ = ~new_n30710_ & new_n30715_;
  assign new_n30717_ = ~pi0618 & ~new_n30704_;
  assign new_n30718_ = pi0618 & ~new_n30707_;
  assign new_n30719_ = ~pi1154 & ~new_n30718_;
  assign new_n30720_ = ~new_n30717_ & new_n30719_;
  assign new_n30721_ = new_n20311_ & new_n30711_;
  assign new_n30722_ = pi1154 & ~new_n30654_;
  assign new_n30723_ = ~new_n30721_ & new_n30722_;
  assign new_n30724_ = ~pi0627 & ~new_n30723_;
  assign new_n30725_ = ~new_n30720_ & new_n30724_;
  assign new_n30726_ = ~new_n30716_ & ~new_n30725_;
  assign new_n30727_ = pi0781 & ~new_n30726_;
  assign new_n30728_ = ~pi0781 & ~new_n30704_;
  assign new_n30729_ = ~new_n23615_ & ~new_n30728_;
  assign new_n30730_ = ~new_n30727_ & new_n30729_;
  assign new_n30731_ = new_n19280_ & new_n30683_;
  assign new_n30732_ = ~new_n23613_ & ~new_n30731_;
  assign new_n30733_ = ~new_n20229_ & new_n30711_;
  assign new_n30734_ = new_n20336_ & new_n30733_;
  assign new_n30735_ = new_n17689_ & ~new_n30734_;
  assign new_n30736_ = new_n20346_ & new_n30733_;
  assign new_n30737_ = new_n17688_ & ~new_n30736_;
  assign new_n30738_ = ~new_n30735_ & ~new_n30737_;
  assign new_n30739_ = ~new_n30732_ & new_n30738_;
  assign new_n30740_ = pi0789 & ~new_n30654_;
  assign new_n30741_ = ~new_n30739_ & new_n30740_;
  assign new_n30742_ = new_n17969_ & ~new_n30741_;
  assign new_n30743_ = ~new_n30730_ & new_n30742_;
  assign new_n30744_ = ~new_n17691_ & new_n30731_;
  assign new_n30745_ = ~new_n30654_ & ~new_n30744_;
  assign new_n30746_ = new_n17851_ & ~new_n30745_;
  assign new_n30747_ = new_n20235_ & new_n30711_;
  assign new_n30748_ = pi0626 & new_n30747_;
  assign new_n30749_ = ~new_n30654_ & ~new_n30748_;
  assign new_n30750_ = pi1158 & ~new_n30749_;
  assign new_n30751_ = ~pi0641 & ~new_n30750_;
  assign new_n30752_ = ~new_n30746_ & new_n30751_;
  assign new_n30753_ = new_n17850_ & ~new_n30745_;
  assign new_n30754_ = ~pi0626 & new_n30747_;
  assign new_n30755_ = ~new_n30654_ & ~new_n30754_;
  assign new_n30756_ = ~pi1158 & ~new_n30755_;
  assign new_n30757_ = pi0641 & ~new_n30756_;
  assign new_n30758_ = ~new_n30753_ & new_n30757_;
  assign new_n30759_ = pi0788 & ~new_n30758_;
  assign new_n30760_ = ~new_n30752_ & new_n30759_;
  assign new_n30761_ = ~new_n20364_ & ~new_n30760_;
  assign new_n30762_ = ~new_n30743_ & new_n30761_;
  assign new_n30763_ = ~new_n17968_ & new_n30747_;
  assign new_n30764_ = ~pi0629 & new_n30763_;
  assign new_n30765_ = pi0628 & ~new_n30764_;
  assign new_n30766_ = new_n19281_ & new_n30683_;
  assign new_n30767_ = pi0629 & ~new_n30766_;
  assign new_n30768_ = ~new_n30765_ & ~new_n30767_;
  assign new_n30769_ = ~pi1156 & ~new_n30768_;
  assign new_n30770_ = pi0628 & new_n30766_;
  assign new_n30771_ = ~pi0628 & ~new_n30763_;
  assign new_n30772_ = pi0629 & ~new_n30771_;
  assign new_n30773_ = pi1156 & ~new_n30772_;
  assign new_n30774_ = ~new_n30770_ & new_n30773_;
  assign new_n30775_ = ~new_n30769_ & ~new_n30774_;
  assign new_n30776_ = pi0792 & ~new_n30654_;
  assign new_n30777_ = ~new_n30775_ & new_n30776_;
  assign new_n30778_ = ~new_n30762_ & ~new_n30777_;
  assign new_n30779_ = ~new_n20360_ & ~new_n30778_;
  assign new_n30780_ = ~new_n17762_ & new_n30763_;
  assign new_n30781_ = ~pi0630 & new_n30780_;
  assign new_n30782_ = pi0647 & ~new_n30781_;
  assign new_n30783_ = ~new_n19311_ & new_n30766_;
  assign new_n30784_ = pi0630 & ~new_n30783_;
  assign new_n30785_ = ~new_n30782_ & ~new_n30784_;
  assign new_n30786_ = ~pi1157 & ~new_n30785_;
  assign new_n30787_ = ~pi0630 & ~new_n30783_;
  assign new_n30788_ = pi0647 & ~new_n30787_;
  assign new_n30789_ = pi0630 & new_n30780_;
  assign new_n30790_ = pi1157 & ~new_n30789_;
  assign new_n30791_ = ~new_n30788_ & new_n30790_;
  assign new_n30792_ = ~new_n30786_ & ~new_n30791_;
  assign new_n30793_ = pi0787 & ~new_n30654_;
  assign new_n30794_ = ~new_n30792_ & new_n30793_;
  assign new_n30795_ = ~new_n30779_ & ~new_n30794_;
  assign new_n30796_ = pi0644 & new_n30795_;
  assign new_n30797_ = ~new_n19335_ & new_n30783_;
  assign new_n30798_ = ~new_n30654_ & ~new_n30797_;
  assign new_n30799_ = ~pi0644 & ~new_n30798_;
  assign new_n30800_ = pi0715 & ~new_n30799_;
  assign new_n30801_ = ~new_n30796_ & new_n30800_;
  assign new_n30802_ = ~new_n17968_ & new_n23689_;
  assign new_n30803_ = new_n30747_ & new_n30802_;
  assign new_n30804_ = pi0644 & new_n30803_;
  assign new_n30805_ = ~pi0715 & ~new_n30654_;
  assign new_n30806_ = ~new_n30804_ & new_n30805_;
  assign new_n30807_ = pi1160 & ~new_n30806_;
  assign new_n30808_ = ~new_n30801_ & new_n30807_;
  assign new_n30809_ = ~pi0644 & new_n30795_;
  assign new_n30810_ = pi0644 & ~new_n30798_;
  assign new_n30811_ = ~pi0715 & ~new_n30810_;
  assign new_n30812_ = ~new_n30809_ & new_n30811_;
  assign new_n30813_ = ~pi0644 & new_n30803_;
  assign new_n30814_ = pi0715 & ~new_n30654_;
  assign new_n30815_ = ~new_n30813_ & new_n30814_;
  assign new_n30816_ = ~pi1160 & ~new_n30815_;
  assign new_n30817_ = ~new_n30812_ & new_n30816_;
  assign new_n30818_ = ~new_n30808_ & ~new_n30817_;
  assign new_n30819_ = pi0790 & ~new_n30818_;
  assign new_n30820_ = ~pi0790 & new_n30795_;
  assign new_n30821_ = pi0832 & ~new_n30820_;
  assign new_n30822_ = ~new_n30819_ & new_n30821_;
  assign po0346 = ~new_n30653_ & ~new_n30822_;
  assign new_n30824_ = ~pi0190 & ~new_n2754_;
  assign new_n30825_ = pi0763 & new_n16913_;
  assign new_n30826_ = ~new_n30824_ & ~new_n30825_;
  assign new_n30827_ = ~new_n17858_ & ~new_n30826_;
  assign new_n30828_ = ~pi0785 & ~new_n30827_;
  assign new_n30829_ = new_n17603_ & new_n30825_;
  assign new_n30830_ = new_n30827_ & ~new_n30829_;
  assign new_n30831_ = pi1155 & ~new_n30830_;
  assign new_n30832_ = ~pi1155 & ~new_n30824_;
  assign new_n30833_ = ~new_n30829_ & new_n30832_;
  assign new_n30834_ = ~new_n30831_ & ~new_n30833_;
  assign new_n30835_ = pi0785 & ~new_n30834_;
  assign new_n30836_ = ~new_n30828_ & ~new_n30835_;
  assign new_n30837_ = ~pi0781 & ~new_n30836_;
  assign new_n30838_ = ~new_n17873_ & new_n30836_;
  assign new_n30839_ = pi1154 & ~new_n30838_;
  assign new_n30840_ = ~new_n17876_ & new_n30836_;
  assign new_n30841_ = ~pi1154 & ~new_n30840_;
  assign new_n30842_ = ~new_n30839_ & ~new_n30841_;
  assign new_n30843_ = pi0781 & ~new_n30842_;
  assign new_n30844_ = ~new_n30837_ & ~new_n30843_;
  assign new_n30845_ = ~pi0789 & ~new_n30844_;
  assign new_n30846_ = ~new_n23057_ & new_n30844_;
  assign new_n30847_ = pi1159 & ~new_n30846_;
  assign new_n30848_ = ~new_n23060_ & new_n30844_;
  assign new_n30849_ = ~pi1159 & ~new_n30848_;
  assign new_n30850_ = ~new_n30847_ & ~new_n30849_;
  assign new_n30851_ = pi0789 & ~new_n30850_;
  assign new_n30852_ = ~new_n30845_ & ~new_n30851_;
  assign new_n30853_ = ~new_n17968_ & new_n30852_;
  assign new_n30854_ = new_n17968_ & new_n30824_;
  assign new_n30855_ = ~new_n30853_ & ~new_n30854_;
  assign new_n30856_ = ~new_n17762_ & ~new_n30855_;
  assign new_n30857_ = new_n17762_ & new_n30824_;
  assign new_n30858_ = ~new_n30856_ & ~new_n30857_;
  assign new_n30859_ = ~new_n20556_ & new_n30858_;
  assign new_n30860_ = pi0699 & new_n16915_;
  assign new_n30861_ = ~new_n30824_ & ~new_n30860_;
  assign new_n30862_ = ~pi0778 & ~new_n30861_;
  assign new_n30863_ = ~pi0625 & new_n30860_;
  assign new_n30864_ = ~new_n30861_ & ~new_n30863_;
  assign new_n30865_ = pi1153 & ~new_n30864_;
  assign new_n30866_ = ~pi1153 & ~new_n30824_;
  assign new_n30867_ = ~new_n30863_ & new_n30866_;
  assign new_n30868_ = pi0778 & ~new_n30867_;
  assign new_n30869_ = ~new_n30865_ & new_n30868_;
  assign new_n30870_ = ~new_n30862_ & ~new_n30869_;
  assign new_n30871_ = ~new_n17844_ & ~new_n30870_;
  assign new_n30872_ = ~new_n17846_ & new_n30871_;
  assign new_n30873_ = ~new_n17848_ & new_n30872_;
  assign new_n30874_ = ~new_n17980_ & new_n30873_;
  assign new_n30875_ = ~new_n18011_ & new_n30874_;
  assign new_n30876_ = ~pi0647 & new_n30875_;
  assign new_n30877_ = pi0647 & new_n30824_;
  assign new_n30878_ = ~pi1157 & ~new_n30877_;
  assign new_n30879_ = ~new_n30876_ & new_n30878_;
  assign new_n30880_ = pi0630 & new_n30879_;
  assign new_n30881_ = pi0647 & ~new_n30875_;
  assign new_n30882_ = ~pi0647 & ~new_n30824_;
  assign new_n30883_ = ~new_n30881_ & ~new_n30882_;
  assign new_n30884_ = new_n17801_ & ~new_n30883_;
  assign new_n30885_ = ~new_n30880_ & ~new_n30884_;
  assign new_n30886_ = ~new_n30859_ & new_n30885_;
  assign new_n30887_ = pi0787 & ~new_n30886_;
  assign new_n30888_ = pi0626 & ~new_n30852_;
  assign new_n30889_ = ~pi0626 & ~new_n30824_;
  assign new_n30890_ = new_n17731_ & ~new_n30889_;
  assign new_n30891_ = ~new_n30888_ & new_n30890_;
  assign new_n30892_ = new_n17856_ & new_n30873_;
  assign new_n30893_ = ~pi0626 & ~new_n30852_;
  assign new_n30894_ = pi0626 & ~new_n30824_;
  assign new_n30895_ = new_n17732_ & ~new_n30894_;
  assign new_n30896_ = ~new_n30893_ & new_n30895_;
  assign new_n30897_ = ~new_n30892_ & ~new_n30896_;
  assign new_n30898_ = ~new_n30891_ & new_n30897_;
  assign new_n30899_ = pi0788 & ~new_n30898_;
  assign new_n30900_ = ~new_n16639_ & ~new_n30861_;
  assign new_n30901_ = pi0625 & new_n30900_;
  assign new_n30902_ = new_n30826_ & ~new_n30900_;
  assign new_n30903_ = ~new_n30901_ & ~new_n30902_;
  assign new_n30904_ = new_n30866_ & ~new_n30903_;
  assign new_n30905_ = ~pi0608 & ~new_n30865_;
  assign new_n30906_ = ~new_n30904_ & new_n30905_;
  assign new_n30907_ = pi1153 & new_n30826_;
  assign new_n30908_ = ~new_n30901_ & new_n30907_;
  assign new_n30909_ = pi0608 & ~new_n30867_;
  assign new_n30910_ = ~new_n30908_ & new_n30909_;
  assign new_n30911_ = ~new_n30906_ & ~new_n30910_;
  assign new_n30912_ = pi0778 & ~new_n30911_;
  assign new_n30913_ = ~pi0778 & ~new_n30902_;
  assign new_n30914_ = ~new_n30912_ & ~new_n30913_;
  assign new_n30915_ = ~pi0609 & ~new_n30914_;
  assign new_n30916_ = pi0609 & ~new_n30870_;
  assign new_n30917_ = ~pi1155 & ~new_n30916_;
  assign new_n30918_ = ~new_n30915_ & new_n30917_;
  assign new_n30919_ = ~pi0660 & ~new_n30831_;
  assign new_n30920_ = ~new_n30918_ & new_n30919_;
  assign new_n30921_ = pi0609 & ~new_n30914_;
  assign new_n30922_ = ~pi0609 & ~new_n30870_;
  assign new_n30923_ = pi1155 & ~new_n30922_;
  assign new_n30924_ = ~new_n30921_ & new_n30923_;
  assign new_n30925_ = pi0660 & ~new_n30833_;
  assign new_n30926_ = ~new_n30924_ & new_n30925_;
  assign new_n30927_ = ~new_n30920_ & ~new_n30926_;
  assign new_n30928_ = pi0785 & ~new_n30927_;
  assign new_n30929_ = ~pi0785 & ~new_n30914_;
  assign new_n30930_ = ~new_n30928_ & ~new_n30929_;
  assign new_n30931_ = ~pi0618 & ~new_n30930_;
  assign new_n30932_ = pi0618 & new_n30871_;
  assign new_n30933_ = ~pi1154 & ~new_n30932_;
  assign new_n30934_ = ~new_n30931_ & new_n30933_;
  assign new_n30935_ = ~pi0627 & ~new_n30839_;
  assign new_n30936_ = ~new_n30934_ & new_n30935_;
  assign new_n30937_ = pi0618 & ~new_n30930_;
  assign new_n30938_ = ~pi0618 & new_n30871_;
  assign new_n30939_ = pi1154 & ~new_n30938_;
  assign new_n30940_ = ~new_n30937_ & new_n30939_;
  assign new_n30941_ = pi0627 & ~new_n30841_;
  assign new_n30942_ = ~new_n30940_ & new_n30941_;
  assign new_n30943_ = ~new_n30936_ & ~new_n30942_;
  assign new_n30944_ = pi0781 & ~new_n30943_;
  assign new_n30945_ = ~pi0781 & ~new_n30930_;
  assign new_n30946_ = ~new_n30944_ & ~new_n30945_;
  assign new_n30947_ = pi0619 & ~new_n30946_;
  assign new_n30948_ = ~pi0619 & new_n30872_;
  assign new_n30949_ = pi1159 & ~new_n30948_;
  assign new_n30950_ = ~new_n30947_ & new_n30949_;
  assign new_n30951_ = pi0648 & ~new_n30849_;
  assign new_n30952_ = ~new_n30950_ & new_n30951_;
  assign new_n30953_ = ~pi0619 & ~new_n30946_;
  assign new_n30954_ = pi0619 & new_n30872_;
  assign new_n30955_ = ~pi1159 & ~new_n30954_;
  assign new_n30956_ = ~new_n30953_ & new_n30955_;
  assign new_n30957_ = ~pi0648 & ~new_n30847_;
  assign new_n30958_ = ~new_n30956_ & new_n30957_;
  assign new_n30959_ = pi0789 & ~new_n30958_;
  assign new_n30960_ = ~new_n30952_ & new_n30959_;
  assign new_n30961_ = ~pi0789 & new_n30946_;
  assign new_n30962_ = new_n17969_ & ~new_n30961_;
  assign new_n30963_ = ~new_n30960_ & new_n30962_;
  assign new_n30964_ = ~new_n30899_ & ~new_n30963_;
  assign new_n30965_ = ~new_n20364_ & ~new_n30964_;
  assign new_n30966_ = new_n18008_ & ~new_n30855_;
  assign new_n30967_ = new_n20851_ & new_n30874_;
  assign new_n30968_ = ~new_n30966_ & ~new_n30967_;
  assign new_n30969_ = ~pi0629 & ~new_n30968_;
  assign new_n30970_ = new_n20855_ & new_n30874_;
  assign new_n30971_ = new_n18007_ & ~new_n30855_;
  assign new_n30972_ = ~new_n30970_ & ~new_n30971_;
  assign new_n30973_ = pi0629 & ~new_n30972_;
  assign new_n30974_ = ~new_n30969_ & ~new_n30973_;
  assign new_n30975_ = pi0792 & ~new_n30974_;
  assign new_n30976_ = ~new_n20360_ & ~new_n30975_;
  assign new_n30977_ = ~new_n30965_ & new_n30976_;
  assign new_n30978_ = ~new_n30887_ & ~new_n30977_;
  assign new_n30979_ = pi0644 & new_n30978_;
  assign new_n30980_ = ~pi0787 & ~new_n30875_;
  assign new_n30981_ = pi1157 & ~new_n30883_;
  assign new_n30982_ = ~new_n30879_ & ~new_n30981_;
  assign new_n30983_ = pi0787 & ~new_n30982_;
  assign new_n30984_ = ~new_n30980_ & ~new_n30983_;
  assign new_n30985_ = ~pi0644 & new_n30984_;
  assign new_n30986_ = pi0715 & ~new_n30985_;
  assign new_n30987_ = ~new_n30979_ & new_n30986_;
  assign new_n30988_ = ~new_n17804_ & ~new_n30858_;
  assign new_n30989_ = new_n17804_ & new_n30824_;
  assign new_n30990_ = ~new_n30988_ & ~new_n30989_;
  assign new_n30991_ = pi0644 & ~new_n30990_;
  assign new_n30992_ = ~pi0644 & new_n30824_;
  assign new_n30993_ = ~pi0715 & ~new_n30992_;
  assign new_n30994_ = ~new_n30991_ & new_n30993_;
  assign new_n30995_ = pi1160 & ~new_n30994_;
  assign new_n30996_ = ~new_n30987_ & new_n30995_;
  assign new_n30997_ = ~pi0644 & new_n30978_;
  assign new_n30998_ = pi0644 & new_n30984_;
  assign new_n30999_ = ~pi0715 & ~new_n30998_;
  assign new_n31000_ = ~new_n30997_ & new_n30999_;
  assign new_n31001_ = ~pi0644 & ~new_n30990_;
  assign new_n31002_ = pi0644 & new_n30824_;
  assign new_n31003_ = pi0715 & ~new_n31002_;
  assign new_n31004_ = ~new_n31001_ & new_n31003_;
  assign new_n31005_ = ~pi1160 & ~new_n31004_;
  assign new_n31006_ = ~new_n31000_ & new_n31005_;
  assign new_n31007_ = ~new_n30996_ & ~new_n31006_;
  assign new_n31008_ = pi0790 & ~new_n31007_;
  assign new_n31009_ = ~pi0790 & new_n30978_;
  assign new_n31010_ = pi0832 & ~new_n31009_;
  assign new_n31011_ = ~new_n31008_ & new_n31010_;
  assign new_n31012_ = ~pi0190 & ~new_n17558_;
  assign new_n31013_ = new_n17691_ & ~new_n31012_;
  assign new_n31014_ = pi0190 & ~new_n3272_;
  assign new_n31015_ = ~pi0190 & new_n18124_;
  assign new_n31016_ = pi0190 & ~new_n18128_;
  assign new_n31017_ = ~pi0038 & ~new_n31016_;
  assign new_n31018_ = ~new_n31015_ & new_n31017_;
  assign new_n31019_ = ~pi0190 & ~new_n17431_;
  assign new_n31020_ = new_n17544_ & ~new_n31019_;
  assign new_n31021_ = pi0699 & ~new_n31020_;
  assign new_n31022_ = ~new_n31018_ & new_n31021_;
  assign new_n31023_ = ~pi0190 & ~pi0699;
  assign new_n31024_ = ~new_n17551_ & new_n31023_;
  assign new_n31025_ = new_n3272_ & ~new_n31024_;
  assign new_n31026_ = ~new_n31022_ & new_n31025_;
  assign new_n31027_ = ~new_n31014_ & ~new_n31026_;
  assign new_n31028_ = ~pi0778 & ~new_n31027_;
  assign new_n31029_ = pi0625 & new_n31027_;
  assign new_n31030_ = ~pi0625 & new_n31012_;
  assign new_n31031_ = pi1153 & ~new_n31030_;
  assign new_n31032_ = ~new_n31029_ & new_n31031_;
  assign new_n31033_ = ~pi0625 & new_n31027_;
  assign new_n31034_ = pi0625 & new_n31012_;
  assign new_n31035_ = ~pi1153 & ~new_n31034_;
  assign new_n31036_ = ~new_n31033_ & new_n31035_;
  assign new_n31037_ = ~new_n31032_ & ~new_n31036_;
  assign new_n31038_ = pi0778 & ~new_n31037_;
  assign new_n31039_ = ~new_n31028_ & ~new_n31038_;
  assign new_n31040_ = ~new_n17618_ & ~new_n31039_;
  assign new_n31041_ = new_n17618_ & ~new_n31012_;
  assign new_n31042_ = ~new_n31040_ & ~new_n31041_;
  assign new_n31043_ = ~new_n17655_ & new_n31042_;
  assign new_n31044_ = new_n17655_ & new_n31012_;
  assign new_n31045_ = ~new_n31043_ & ~new_n31044_;
  assign new_n31046_ = ~new_n17691_ & new_n31045_;
  assign new_n31047_ = ~new_n31013_ & ~new_n31046_;
  assign new_n31048_ = ~new_n17734_ & new_n31047_;
  assign new_n31049_ = new_n17734_ & new_n31012_;
  assign new_n31050_ = ~new_n31048_ & ~new_n31049_;
  assign new_n31051_ = ~pi0628 & ~new_n31050_;
  assign new_n31052_ = pi0628 & new_n31012_;
  assign new_n31053_ = ~new_n31051_ & ~new_n31052_;
  assign new_n31054_ = ~pi1156 & ~new_n31053_;
  assign new_n31055_ = pi0628 & ~new_n31050_;
  assign new_n31056_ = ~pi0628 & new_n31012_;
  assign new_n31057_ = ~new_n31055_ & ~new_n31056_;
  assign new_n31058_ = pi1156 & ~new_n31057_;
  assign new_n31059_ = ~new_n31054_ & ~new_n31058_;
  assign new_n31060_ = pi0792 & ~new_n31059_;
  assign new_n31061_ = ~pi0792 & ~new_n31050_;
  assign new_n31062_ = ~new_n31060_ & ~new_n31061_;
  assign new_n31063_ = ~pi0647 & ~new_n31062_;
  assign new_n31064_ = pi0647 & new_n31012_;
  assign new_n31065_ = ~new_n31063_ & ~new_n31064_;
  assign new_n31066_ = ~pi1157 & ~new_n31065_;
  assign new_n31067_ = pi0647 & ~new_n31062_;
  assign new_n31068_ = ~pi0647 & new_n31012_;
  assign new_n31069_ = ~new_n31067_ & ~new_n31068_;
  assign new_n31070_ = pi1157 & ~new_n31069_;
  assign new_n31071_ = ~new_n31066_ & ~new_n31070_;
  assign new_n31072_ = pi0787 & ~new_n31071_;
  assign new_n31073_ = ~pi0787 & ~new_n31062_;
  assign new_n31074_ = ~new_n31072_ & ~new_n31073_;
  assign new_n31075_ = ~pi0644 & ~new_n31074_;
  assign new_n31076_ = pi0715 & ~new_n31075_;
  assign new_n31077_ = ~pi0763 & new_n17347_;
  assign new_n31078_ = pi0190 & new_n17424_;
  assign new_n31079_ = ~new_n31077_ & ~new_n31078_;
  assign new_n31080_ = pi0039 & ~new_n31079_;
  assign new_n31081_ = ~pi0190 & pi0763;
  assign new_n31082_ = new_n17393_ & new_n31081_;
  assign new_n31083_ = pi0763 & ~new_n17397_;
  assign new_n31084_ = pi0190 & ~new_n31083_;
  assign new_n31085_ = ~new_n22356_ & ~new_n31084_;
  assign new_n31086_ = ~new_n31082_ & new_n31085_;
  assign new_n31087_ = ~new_n31080_ & new_n31086_;
  assign new_n31088_ = ~pi0038 & ~new_n31087_;
  assign new_n31089_ = pi0763 & new_n17433_;
  assign new_n31090_ = pi0038 & ~new_n31019_;
  assign new_n31091_ = ~new_n31089_ & new_n31090_;
  assign new_n31092_ = ~new_n31088_ & ~new_n31091_;
  assign new_n31093_ = new_n3272_ & ~new_n31092_;
  assign new_n31094_ = ~new_n31014_ & ~new_n31093_;
  assign new_n31095_ = ~new_n17590_ & ~new_n31094_;
  assign new_n31096_ = new_n17590_ & ~new_n31012_;
  assign new_n31097_ = ~new_n31095_ & ~new_n31096_;
  assign new_n31098_ = ~pi0785 & ~new_n31097_;
  assign new_n31099_ = ~new_n17591_ & ~new_n31012_;
  assign new_n31100_ = pi0609 & new_n31095_;
  assign new_n31101_ = ~new_n31099_ & ~new_n31100_;
  assign new_n31102_ = pi1155 & ~new_n31101_;
  assign new_n31103_ = ~new_n17603_ & ~new_n31012_;
  assign new_n31104_ = ~pi0609 & new_n31095_;
  assign new_n31105_ = ~new_n31103_ & ~new_n31104_;
  assign new_n31106_ = ~pi1155 & ~new_n31105_;
  assign new_n31107_ = ~new_n31102_ & ~new_n31106_;
  assign new_n31108_ = pi0785 & ~new_n31107_;
  assign new_n31109_ = ~new_n31098_ & ~new_n31108_;
  assign new_n31110_ = ~pi0781 & ~new_n31109_;
  assign new_n31111_ = pi0618 & new_n31109_;
  assign new_n31112_ = ~pi0618 & new_n31012_;
  assign new_n31113_ = pi1154 & ~new_n31112_;
  assign new_n31114_ = ~new_n31111_ & new_n31113_;
  assign new_n31115_ = ~pi0618 & new_n31109_;
  assign new_n31116_ = pi0618 & new_n31012_;
  assign new_n31117_ = ~pi1154 & ~new_n31116_;
  assign new_n31118_ = ~new_n31115_ & new_n31117_;
  assign new_n31119_ = ~new_n31114_ & ~new_n31118_;
  assign new_n31120_ = pi0781 & ~new_n31119_;
  assign new_n31121_ = ~new_n31110_ & ~new_n31120_;
  assign new_n31122_ = ~pi0789 & ~new_n31121_;
  assign new_n31123_ = pi0619 & new_n31121_;
  assign new_n31124_ = ~pi0619 & new_n31012_;
  assign new_n31125_ = pi1159 & ~new_n31124_;
  assign new_n31126_ = ~new_n31123_ & new_n31125_;
  assign new_n31127_ = ~pi0619 & new_n31121_;
  assign new_n31128_ = pi0619 & new_n31012_;
  assign new_n31129_ = ~pi1159 & ~new_n31128_;
  assign new_n31130_ = ~new_n31127_ & new_n31129_;
  assign new_n31131_ = ~new_n31126_ & ~new_n31130_;
  assign new_n31132_ = pi0789 & ~new_n31131_;
  assign new_n31133_ = ~new_n31122_ & ~new_n31132_;
  assign new_n31134_ = ~new_n17968_ & new_n31133_;
  assign new_n31135_ = new_n17968_ & new_n31012_;
  assign new_n31136_ = ~new_n31134_ & ~new_n31135_;
  assign new_n31137_ = ~new_n17762_ & ~new_n31136_;
  assign new_n31138_ = new_n17762_ & new_n31012_;
  assign new_n31139_ = ~new_n31137_ & ~new_n31138_;
  assign new_n31140_ = ~new_n17804_ & ~new_n31139_;
  assign new_n31141_ = new_n17804_ & new_n31012_;
  assign new_n31142_ = ~new_n31140_ & ~new_n31141_;
  assign new_n31143_ = pi0644 & ~new_n31142_;
  assign new_n31144_ = ~pi0644 & new_n31012_;
  assign new_n31145_ = ~pi0715 & ~new_n31144_;
  assign new_n31146_ = ~new_n31143_ & new_n31145_;
  assign new_n31147_ = pi1160 & ~new_n31146_;
  assign new_n31148_ = ~new_n31076_ & new_n31147_;
  assign new_n31149_ = pi0644 & ~new_n31074_;
  assign new_n31150_ = ~pi0715 & ~new_n31149_;
  assign new_n31151_ = ~pi0644 & ~new_n31142_;
  assign new_n31152_ = pi0644 & new_n31012_;
  assign new_n31153_ = pi0715 & ~new_n31152_;
  assign new_n31154_ = ~new_n31151_ & new_n31153_;
  assign new_n31155_ = ~pi1160 & ~new_n31154_;
  assign new_n31156_ = ~new_n31150_ & new_n31155_;
  assign new_n31157_ = ~new_n31148_ & ~new_n31156_;
  assign new_n31158_ = pi0790 & ~new_n31157_;
  assign new_n31159_ = pi0644 & new_n31147_;
  assign new_n31160_ = ~pi0644 & new_n31155_;
  assign new_n31161_ = pi0790 & ~new_n31160_;
  assign new_n31162_ = ~new_n31159_ & new_n31161_;
  assign new_n31163_ = ~new_n20567_ & new_n31136_;
  assign new_n31164_ = new_n17760_ & new_n31053_;
  assign new_n31165_ = new_n17759_ & new_n31057_;
  assign new_n31166_ = ~new_n31164_ & ~new_n31165_;
  assign new_n31167_ = ~new_n31163_ & new_n31166_;
  assign new_n31168_ = pi0792 & ~new_n31167_;
  assign new_n31169_ = ~pi0699 & new_n31092_;
  assign new_n31170_ = ~pi0190 & new_n16810_;
  assign new_n31171_ = pi0190 & new_n16928_;
  assign new_n31172_ = ~pi0763 & ~new_n31171_;
  assign new_n31173_ = ~new_n31170_ & new_n31172_;
  assign new_n31174_ = pi0190 & new_n17007_;
  assign new_n31175_ = ~pi0190 & ~new_n17074_;
  assign new_n31176_ = pi0763 & ~new_n31175_;
  assign new_n31177_ = ~new_n31174_ & new_n31176_;
  assign new_n31178_ = pi0039 & ~new_n31177_;
  assign new_n31179_ = ~new_n31173_ & new_n31178_;
  assign new_n31180_ = pi0190 & new_n17178_;
  assign new_n31181_ = ~pi0190 & new_n17217_;
  assign new_n31182_ = ~pi0763 & ~new_n31181_;
  assign new_n31183_ = ~new_n31180_ & new_n31182_;
  assign new_n31184_ = ~pi0190 & ~new_n17227_;
  assign new_n31185_ = pi0190 & ~new_n17234_;
  assign new_n31186_ = pi0763 & ~new_n31185_;
  assign new_n31187_ = ~new_n31184_ & new_n31186_;
  assign new_n31188_ = ~pi0039 & ~new_n31187_;
  assign new_n31189_ = ~new_n31183_ & new_n31188_;
  assign new_n31190_ = ~pi0038 & ~new_n31189_;
  assign new_n31191_ = ~new_n31179_ & new_n31190_;
  assign new_n31192_ = ~pi0763 & new_n24079_;
  assign new_n31193_ = ~new_n17035_ & ~new_n31192_;
  assign new_n31194_ = ~pi0039 & ~new_n31193_;
  assign new_n31195_ = ~pi0190 & ~new_n31194_;
  assign new_n31196_ = ~new_n16916_ & ~new_n30825_;
  assign new_n31197_ = pi0190 & ~new_n31196_;
  assign new_n31198_ = new_n6257_ & new_n31197_;
  assign new_n31199_ = pi0038 & ~new_n31198_;
  assign new_n31200_ = ~new_n31195_ & new_n31199_;
  assign new_n31201_ = pi0699 & ~new_n31200_;
  assign new_n31202_ = ~new_n31191_ & new_n31201_;
  assign new_n31203_ = new_n3272_ & ~new_n31202_;
  assign new_n31204_ = ~new_n31169_ & new_n31203_;
  assign new_n31205_ = ~new_n31014_ & ~new_n31204_;
  assign new_n31206_ = ~pi0625 & new_n31205_;
  assign new_n31207_ = pi0625 & new_n31094_;
  assign new_n31208_ = ~pi1153 & ~new_n31207_;
  assign new_n31209_ = ~new_n31206_ & new_n31208_;
  assign new_n31210_ = ~pi0608 & ~new_n31032_;
  assign new_n31211_ = ~new_n31209_ & new_n31210_;
  assign new_n31212_ = pi0625 & new_n31205_;
  assign new_n31213_ = ~pi0625 & new_n31094_;
  assign new_n31214_ = pi1153 & ~new_n31213_;
  assign new_n31215_ = ~new_n31212_ & new_n31214_;
  assign new_n31216_ = pi0608 & ~new_n31036_;
  assign new_n31217_ = ~new_n31215_ & new_n31216_;
  assign new_n31218_ = ~new_n31211_ & ~new_n31217_;
  assign new_n31219_ = pi0778 & ~new_n31218_;
  assign new_n31220_ = ~pi0778 & new_n31205_;
  assign new_n31221_ = ~new_n31219_ & ~new_n31220_;
  assign new_n31222_ = ~pi0609 & ~new_n31221_;
  assign new_n31223_ = pi0609 & new_n31039_;
  assign new_n31224_ = ~pi1155 & ~new_n31223_;
  assign new_n31225_ = ~new_n31222_ & new_n31224_;
  assign new_n31226_ = ~pi0660 & ~new_n31102_;
  assign new_n31227_ = ~new_n31225_ & new_n31226_;
  assign new_n31228_ = pi0609 & ~new_n31221_;
  assign new_n31229_ = ~pi0609 & new_n31039_;
  assign new_n31230_ = pi1155 & ~new_n31229_;
  assign new_n31231_ = ~new_n31228_ & new_n31230_;
  assign new_n31232_ = pi0660 & ~new_n31106_;
  assign new_n31233_ = ~new_n31231_ & new_n31232_;
  assign new_n31234_ = ~new_n31227_ & ~new_n31233_;
  assign new_n31235_ = pi0785 & ~new_n31234_;
  assign new_n31236_ = ~pi0785 & ~new_n31221_;
  assign new_n31237_ = ~new_n31235_ & ~new_n31236_;
  assign new_n31238_ = ~pi0618 & ~new_n31237_;
  assign new_n31239_ = pi0618 & new_n31042_;
  assign new_n31240_ = ~pi1154 & ~new_n31239_;
  assign new_n31241_ = ~new_n31238_ & new_n31240_;
  assign new_n31242_ = ~pi0627 & ~new_n31114_;
  assign new_n31243_ = ~new_n31241_ & new_n31242_;
  assign new_n31244_ = pi0618 & ~new_n31237_;
  assign new_n31245_ = ~pi0618 & new_n31042_;
  assign new_n31246_ = pi1154 & ~new_n31245_;
  assign new_n31247_ = ~new_n31244_ & new_n31246_;
  assign new_n31248_ = pi0627 & ~new_n31118_;
  assign new_n31249_ = ~new_n31247_ & new_n31248_;
  assign new_n31250_ = ~new_n31243_ & ~new_n31249_;
  assign new_n31251_ = pi0781 & ~new_n31250_;
  assign new_n31252_ = ~pi0781 & ~new_n31237_;
  assign new_n31253_ = ~new_n31251_ & ~new_n31252_;
  assign new_n31254_ = pi0619 & ~new_n31253_;
  assign new_n31255_ = ~pi0619 & ~new_n31045_;
  assign new_n31256_ = pi1159 & ~new_n31255_;
  assign new_n31257_ = ~new_n31254_ & new_n31256_;
  assign new_n31258_ = pi0648 & ~new_n31130_;
  assign new_n31259_ = ~new_n31257_ & new_n31258_;
  assign new_n31260_ = ~pi0619 & ~new_n31253_;
  assign new_n31261_ = pi0619 & ~new_n31045_;
  assign new_n31262_ = ~pi1159 & ~new_n31261_;
  assign new_n31263_ = ~new_n31260_ & new_n31262_;
  assign new_n31264_ = ~pi0648 & ~new_n31126_;
  assign new_n31265_ = ~new_n31263_ & new_n31264_;
  assign new_n31266_ = pi0789 & ~new_n31265_;
  assign new_n31267_ = ~new_n31259_ & new_n31266_;
  assign new_n31268_ = ~pi0789 & new_n31253_;
  assign new_n31269_ = new_n17969_ & ~new_n31268_;
  assign new_n31270_ = ~new_n31267_ & new_n31269_;
  assign new_n31271_ = pi0626 & ~new_n31133_;
  assign new_n31272_ = ~pi0626 & ~new_n31012_;
  assign new_n31273_ = new_n17731_ & ~new_n31272_;
  assign new_n31274_ = ~new_n31271_ & new_n31273_;
  assign new_n31275_ = new_n17856_ & new_n31047_;
  assign new_n31276_ = ~pi0626 & ~new_n31133_;
  assign new_n31277_ = pi0626 & ~new_n31012_;
  assign new_n31278_ = new_n17732_ & ~new_n31277_;
  assign new_n31279_ = ~new_n31276_ & new_n31278_;
  assign new_n31280_ = ~new_n31275_ & ~new_n31279_;
  assign new_n31281_ = ~new_n31274_ & new_n31280_;
  assign new_n31282_ = pi0788 & ~new_n31281_;
  assign new_n31283_ = ~new_n20364_ & ~new_n31282_;
  assign new_n31284_ = ~new_n31270_ & new_n31283_;
  assign new_n31285_ = ~new_n31168_ & ~new_n31284_;
  assign new_n31286_ = ~new_n20360_ & ~new_n31285_;
  assign new_n31287_ = new_n17801_ & new_n31069_;
  assign new_n31288_ = new_n17802_ & new_n31065_;
  assign new_n31289_ = ~new_n20556_ & new_n31139_;
  assign new_n31290_ = ~new_n31288_ & ~new_n31289_;
  assign new_n31291_ = ~new_n31287_ & new_n31290_;
  assign new_n31292_ = pi0787 & ~new_n31291_;
  assign new_n31293_ = ~new_n31286_ & ~new_n31292_;
  assign new_n31294_ = ~new_n31162_ & new_n31293_;
  assign new_n31295_ = ~new_n31158_ & ~new_n31294_;
  assign new_n31296_ = ~po1038 & ~new_n31295_;
  assign new_n31297_ = ~pi0190 & po1038;
  assign new_n31298_ = ~pi0832 & ~new_n31297_;
  assign new_n31299_ = ~new_n31296_ & new_n31298_;
  assign po0347 = ~new_n31011_ & ~new_n31299_;
  assign new_n31301_ = ~pi0191 & ~new_n2754_;
  assign new_n31302_ = pi0746 & new_n16913_;
  assign new_n31303_ = ~new_n31301_ & ~new_n31302_;
  assign new_n31304_ = ~new_n17858_ & ~new_n31303_;
  assign new_n31305_ = ~pi0785 & ~new_n31304_;
  assign new_n31306_ = new_n17603_ & new_n31302_;
  assign new_n31307_ = new_n31304_ & ~new_n31306_;
  assign new_n31308_ = pi1155 & ~new_n31307_;
  assign new_n31309_ = ~pi1155 & ~new_n31301_;
  assign new_n31310_ = ~new_n31306_ & new_n31309_;
  assign new_n31311_ = ~new_n31308_ & ~new_n31310_;
  assign new_n31312_ = pi0785 & ~new_n31311_;
  assign new_n31313_ = ~new_n31305_ & ~new_n31312_;
  assign new_n31314_ = ~pi0781 & ~new_n31313_;
  assign new_n31315_ = ~new_n17873_ & new_n31313_;
  assign new_n31316_ = pi1154 & ~new_n31315_;
  assign new_n31317_ = ~new_n17876_ & new_n31313_;
  assign new_n31318_ = ~pi1154 & ~new_n31317_;
  assign new_n31319_ = ~new_n31316_ & ~new_n31318_;
  assign new_n31320_ = pi0781 & ~new_n31319_;
  assign new_n31321_ = ~new_n31314_ & ~new_n31320_;
  assign new_n31322_ = ~pi0789 & ~new_n31321_;
  assign new_n31323_ = ~new_n23057_ & new_n31321_;
  assign new_n31324_ = pi1159 & ~new_n31323_;
  assign new_n31325_ = ~new_n23060_ & new_n31321_;
  assign new_n31326_ = ~pi1159 & ~new_n31325_;
  assign new_n31327_ = ~new_n31324_ & ~new_n31326_;
  assign new_n31328_ = pi0789 & ~new_n31327_;
  assign new_n31329_ = ~new_n31322_ & ~new_n31328_;
  assign new_n31330_ = ~new_n17968_ & new_n31329_;
  assign new_n31331_ = new_n17968_ & new_n31301_;
  assign new_n31332_ = ~new_n31330_ & ~new_n31331_;
  assign new_n31333_ = ~new_n17762_ & ~new_n31332_;
  assign new_n31334_ = new_n17762_ & new_n31301_;
  assign new_n31335_ = ~new_n31333_ & ~new_n31334_;
  assign new_n31336_ = ~new_n20556_ & new_n31335_;
  assign new_n31337_ = pi0729 & new_n16915_;
  assign new_n31338_ = ~new_n31301_ & ~new_n31337_;
  assign new_n31339_ = ~pi0778 & ~new_n31338_;
  assign new_n31340_ = ~pi0625 & new_n31337_;
  assign new_n31341_ = ~new_n31338_ & ~new_n31340_;
  assign new_n31342_ = pi1153 & ~new_n31341_;
  assign new_n31343_ = ~pi1153 & ~new_n31301_;
  assign new_n31344_ = ~new_n31340_ & new_n31343_;
  assign new_n31345_ = pi0778 & ~new_n31344_;
  assign new_n31346_ = ~new_n31342_ & new_n31345_;
  assign new_n31347_ = ~new_n31339_ & ~new_n31346_;
  assign new_n31348_ = ~new_n17844_ & ~new_n31347_;
  assign new_n31349_ = ~new_n17846_ & new_n31348_;
  assign new_n31350_ = ~new_n17848_ & new_n31349_;
  assign new_n31351_ = ~new_n17980_ & new_n31350_;
  assign new_n31352_ = ~new_n18011_ & new_n31351_;
  assign new_n31353_ = ~pi0647 & new_n31352_;
  assign new_n31354_ = pi0647 & new_n31301_;
  assign new_n31355_ = ~pi1157 & ~new_n31354_;
  assign new_n31356_ = ~new_n31353_ & new_n31355_;
  assign new_n31357_ = pi0630 & new_n31356_;
  assign new_n31358_ = pi0647 & ~new_n31352_;
  assign new_n31359_ = ~pi0647 & ~new_n31301_;
  assign new_n31360_ = ~new_n31358_ & ~new_n31359_;
  assign new_n31361_ = new_n17801_ & ~new_n31360_;
  assign new_n31362_ = ~new_n31357_ & ~new_n31361_;
  assign new_n31363_ = ~new_n31336_ & new_n31362_;
  assign new_n31364_ = pi0787 & ~new_n31363_;
  assign new_n31365_ = pi0626 & ~new_n31329_;
  assign new_n31366_ = ~pi0626 & ~new_n31301_;
  assign new_n31367_ = new_n17731_ & ~new_n31366_;
  assign new_n31368_ = ~new_n31365_ & new_n31367_;
  assign new_n31369_ = new_n17856_ & new_n31350_;
  assign new_n31370_ = ~pi0626 & ~new_n31329_;
  assign new_n31371_ = pi0626 & ~new_n31301_;
  assign new_n31372_ = new_n17732_ & ~new_n31371_;
  assign new_n31373_ = ~new_n31370_ & new_n31372_;
  assign new_n31374_ = ~new_n31369_ & ~new_n31373_;
  assign new_n31375_ = ~new_n31368_ & new_n31374_;
  assign new_n31376_ = pi0788 & ~new_n31375_;
  assign new_n31377_ = ~new_n16639_ & ~new_n31338_;
  assign new_n31378_ = pi0625 & new_n31377_;
  assign new_n31379_ = new_n31303_ & ~new_n31377_;
  assign new_n31380_ = ~new_n31378_ & ~new_n31379_;
  assign new_n31381_ = new_n31343_ & ~new_n31380_;
  assign new_n31382_ = ~pi0608 & ~new_n31342_;
  assign new_n31383_ = ~new_n31381_ & new_n31382_;
  assign new_n31384_ = pi1153 & new_n31303_;
  assign new_n31385_ = ~new_n31378_ & new_n31384_;
  assign new_n31386_ = pi0608 & ~new_n31344_;
  assign new_n31387_ = ~new_n31385_ & new_n31386_;
  assign new_n31388_ = ~new_n31383_ & ~new_n31387_;
  assign new_n31389_ = pi0778 & ~new_n31388_;
  assign new_n31390_ = ~pi0778 & ~new_n31379_;
  assign new_n31391_ = ~new_n31389_ & ~new_n31390_;
  assign new_n31392_ = ~pi0609 & ~new_n31391_;
  assign new_n31393_ = pi0609 & ~new_n31347_;
  assign new_n31394_ = ~pi1155 & ~new_n31393_;
  assign new_n31395_ = ~new_n31392_ & new_n31394_;
  assign new_n31396_ = ~pi0660 & ~new_n31308_;
  assign new_n31397_ = ~new_n31395_ & new_n31396_;
  assign new_n31398_ = pi0609 & ~new_n31391_;
  assign new_n31399_ = ~pi0609 & ~new_n31347_;
  assign new_n31400_ = pi1155 & ~new_n31399_;
  assign new_n31401_ = ~new_n31398_ & new_n31400_;
  assign new_n31402_ = pi0660 & ~new_n31310_;
  assign new_n31403_ = ~new_n31401_ & new_n31402_;
  assign new_n31404_ = ~new_n31397_ & ~new_n31403_;
  assign new_n31405_ = pi0785 & ~new_n31404_;
  assign new_n31406_ = ~pi0785 & ~new_n31391_;
  assign new_n31407_ = ~new_n31405_ & ~new_n31406_;
  assign new_n31408_ = ~pi0618 & ~new_n31407_;
  assign new_n31409_ = pi0618 & new_n31348_;
  assign new_n31410_ = ~pi1154 & ~new_n31409_;
  assign new_n31411_ = ~new_n31408_ & new_n31410_;
  assign new_n31412_ = ~pi0627 & ~new_n31316_;
  assign new_n31413_ = ~new_n31411_ & new_n31412_;
  assign new_n31414_ = pi0618 & ~new_n31407_;
  assign new_n31415_ = ~pi0618 & new_n31348_;
  assign new_n31416_ = pi1154 & ~new_n31415_;
  assign new_n31417_ = ~new_n31414_ & new_n31416_;
  assign new_n31418_ = pi0627 & ~new_n31318_;
  assign new_n31419_ = ~new_n31417_ & new_n31418_;
  assign new_n31420_ = ~new_n31413_ & ~new_n31419_;
  assign new_n31421_ = pi0781 & ~new_n31420_;
  assign new_n31422_ = ~pi0781 & ~new_n31407_;
  assign new_n31423_ = ~new_n31421_ & ~new_n31422_;
  assign new_n31424_ = pi0619 & ~new_n31423_;
  assign new_n31425_ = ~pi0619 & new_n31349_;
  assign new_n31426_ = pi1159 & ~new_n31425_;
  assign new_n31427_ = ~new_n31424_ & new_n31426_;
  assign new_n31428_ = pi0648 & ~new_n31326_;
  assign new_n31429_ = ~new_n31427_ & new_n31428_;
  assign new_n31430_ = ~pi0619 & ~new_n31423_;
  assign new_n31431_ = pi0619 & new_n31349_;
  assign new_n31432_ = ~pi1159 & ~new_n31431_;
  assign new_n31433_ = ~new_n31430_ & new_n31432_;
  assign new_n31434_ = ~pi0648 & ~new_n31324_;
  assign new_n31435_ = ~new_n31433_ & new_n31434_;
  assign new_n31436_ = pi0789 & ~new_n31435_;
  assign new_n31437_ = ~new_n31429_ & new_n31436_;
  assign new_n31438_ = ~pi0789 & new_n31423_;
  assign new_n31439_ = new_n17969_ & ~new_n31438_;
  assign new_n31440_ = ~new_n31437_ & new_n31439_;
  assign new_n31441_ = ~new_n31376_ & ~new_n31440_;
  assign new_n31442_ = ~new_n20364_ & ~new_n31441_;
  assign new_n31443_ = new_n18008_ & ~new_n31332_;
  assign new_n31444_ = new_n20851_ & new_n31351_;
  assign new_n31445_ = ~new_n31443_ & ~new_n31444_;
  assign new_n31446_ = ~pi0629 & ~new_n31445_;
  assign new_n31447_ = new_n20855_ & new_n31351_;
  assign new_n31448_ = new_n18007_ & ~new_n31332_;
  assign new_n31449_ = ~new_n31447_ & ~new_n31448_;
  assign new_n31450_ = pi0629 & ~new_n31449_;
  assign new_n31451_ = ~new_n31446_ & ~new_n31450_;
  assign new_n31452_ = pi0792 & ~new_n31451_;
  assign new_n31453_ = ~new_n20360_ & ~new_n31452_;
  assign new_n31454_ = ~new_n31442_ & new_n31453_;
  assign new_n31455_ = ~new_n31364_ & ~new_n31454_;
  assign new_n31456_ = pi0644 & new_n31455_;
  assign new_n31457_ = ~pi0787 & ~new_n31352_;
  assign new_n31458_ = pi1157 & ~new_n31360_;
  assign new_n31459_ = ~new_n31356_ & ~new_n31458_;
  assign new_n31460_ = pi0787 & ~new_n31459_;
  assign new_n31461_ = ~new_n31457_ & ~new_n31460_;
  assign new_n31462_ = ~pi0644 & new_n31461_;
  assign new_n31463_ = pi0715 & ~new_n31462_;
  assign new_n31464_ = ~new_n31456_ & new_n31463_;
  assign new_n31465_ = ~new_n17804_ & ~new_n31335_;
  assign new_n31466_ = new_n17804_ & new_n31301_;
  assign new_n31467_ = ~new_n31465_ & ~new_n31466_;
  assign new_n31468_ = pi0644 & ~new_n31467_;
  assign new_n31469_ = ~pi0644 & new_n31301_;
  assign new_n31470_ = ~pi0715 & ~new_n31469_;
  assign new_n31471_ = ~new_n31468_ & new_n31470_;
  assign new_n31472_ = pi1160 & ~new_n31471_;
  assign new_n31473_ = ~new_n31464_ & new_n31472_;
  assign new_n31474_ = ~pi0644 & new_n31455_;
  assign new_n31475_ = pi0644 & new_n31461_;
  assign new_n31476_ = ~pi0715 & ~new_n31475_;
  assign new_n31477_ = ~new_n31474_ & new_n31476_;
  assign new_n31478_ = ~pi0644 & ~new_n31467_;
  assign new_n31479_ = pi0644 & new_n31301_;
  assign new_n31480_ = pi0715 & ~new_n31479_;
  assign new_n31481_ = ~new_n31478_ & new_n31480_;
  assign new_n31482_ = ~pi1160 & ~new_n31481_;
  assign new_n31483_ = ~new_n31477_ & new_n31482_;
  assign new_n31484_ = ~new_n31473_ & ~new_n31483_;
  assign new_n31485_ = pi0790 & ~new_n31484_;
  assign new_n31486_ = ~pi0790 & new_n31455_;
  assign new_n31487_ = pi0832 & ~new_n31486_;
  assign new_n31488_ = ~new_n31485_ & new_n31487_;
  assign new_n31489_ = ~pi0191 & ~new_n17558_;
  assign new_n31490_ = new_n17691_ & ~new_n31489_;
  assign new_n31491_ = pi0191 & ~new_n3272_;
  assign new_n31492_ = ~pi0191 & new_n18124_;
  assign new_n31493_ = pi0191 & ~new_n18128_;
  assign new_n31494_ = ~pi0038 & ~new_n31493_;
  assign new_n31495_ = ~new_n31492_ & new_n31494_;
  assign new_n31496_ = ~pi0191 & ~new_n17431_;
  assign new_n31497_ = new_n17544_ & ~new_n31496_;
  assign new_n31498_ = pi0729 & ~new_n31497_;
  assign new_n31499_ = ~new_n31495_ & new_n31498_;
  assign new_n31500_ = ~pi0191 & ~pi0729;
  assign new_n31501_ = ~new_n17551_ & new_n31500_;
  assign new_n31502_ = new_n3272_ & ~new_n31501_;
  assign new_n31503_ = ~new_n31499_ & new_n31502_;
  assign new_n31504_ = ~new_n31491_ & ~new_n31503_;
  assign new_n31505_ = ~pi0778 & ~new_n31504_;
  assign new_n31506_ = pi0625 & new_n31504_;
  assign new_n31507_ = ~pi0625 & new_n31489_;
  assign new_n31508_ = pi1153 & ~new_n31507_;
  assign new_n31509_ = ~new_n31506_ & new_n31508_;
  assign new_n31510_ = ~pi0625 & new_n31504_;
  assign new_n31511_ = pi0625 & new_n31489_;
  assign new_n31512_ = ~pi1153 & ~new_n31511_;
  assign new_n31513_ = ~new_n31510_ & new_n31512_;
  assign new_n31514_ = ~new_n31509_ & ~new_n31513_;
  assign new_n31515_ = pi0778 & ~new_n31514_;
  assign new_n31516_ = ~new_n31505_ & ~new_n31515_;
  assign new_n31517_ = ~new_n17618_ & ~new_n31516_;
  assign new_n31518_ = new_n17618_ & ~new_n31489_;
  assign new_n31519_ = ~new_n31517_ & ~new_n31518_;
  assign new_n31520_ = ~new_n17655_ & new_n31519_;
  assign new_n31521_ = new_n17655_ & new_n31489_;
  assign new_n31522_ = ~new_n31520_ & ~new_n31521_;
  assign new_n31523_ = ~new_n17691_ & new_n31522_;
  assign new_n31524_ = ~new_n31490_ & ~new_n31523_;
  assign new_n31525_ = ~new_n17734_ & new_n31524_;
  assign new_n31526_ = new_n17734_ & new_n31489_;
  assign new_n31527_ = ~new_n31525_ & ~new_n31526_;
  assign new_n31528_ = ~pi0628 & ~new_n31527_;
  assign new_n31529_ = pi0628 & new_n31489_;
  assign new_n31530_ = ~new_n31528_ & ~new_n31529_;
  assign new_n31531_ = ~pi1156 & ~new_n31530_;
  assign new_n31532_ = pi0628 & ~new_n31527_;
  assign new_n31533_ = ~pi0628 & new_n31489_;
  assign new_n31534_ = ~new_n31532_ & ~new_n31533_;
  assign new_n31535_ = pi1156 & ~new_n31534_;
  assign new_n31536_ = ~new_n31531_ & ~new_n31535_;
  assign new_n31537_ = pi0792 & ~new_n31536_;
  assign new_n31538_ = ~pi0792 & ~new_n31527_;
  assign new_n31539_ = ~new_n31537_ & ~new_n31538_;
  assign new_n31540_ = ~pi0647 & ~new_n31539_;
  assign new_n31541_ = pi0647 & new_n31489_;
  assign new_n31542_ = ~new_n31540_ & ~new_n31541_;
  assign new_n31543_ = ~pi1157 & ~new_n31542_;
  assign new_n31544_ = pi0647 & ~new_n31539_;
  assign new_n31545_ = ~pi0647 & new_n31489_;
  assign new_n31546_ = ~new_n31544_ & ~new_n31545_;
  assign new_n31547_ = pi1157 & ~new_n31546_;
  assign new_n31548_ = ~new_n31543_ & ~new_n31547_;
  assign new_n31549_ = pi0787 & ~new_n31548_;
  assign new_n31550_ = ~pi0787 & ~new_n31539_;
  assign new_n31551_ = ~new_n31549_ & ~new_n31550_;
  assign new_n31552_ = ~pi0644 & ~new_n31551_;
  assign new_n31553_ = pi0715 & ~new_n31552_;
  assign new_n31554_ = ~pi0746 & new_n17347_;
  assign new_n31555_ = pi0191 & new_n17424_;
  assign new_n31556_ = ~new_n31554_ & ~new_n31555_;
  assign new_n31557_ = pi0039 & ~new_n31556_;
  assign new_n31558_ = ~pi0191 & pi0746;
  assign new_n31559_ = new_n17393_ & new_n31558_;
  assign new_n31560_ = pi0746 & ~new_n17397_;
  assign new_n31561_ = pi0191 & ~new_n31560_;
  assign new_n31562_ = ~new_n22437_ & ~new_n31561_;
  assign new_n31563_ = ~new_n31559_ & new_n31562_;
  assign new_n31564_ = ~new_n31557_ & new_n31563_;
  assign new_n31565_ = ~pi0038 & ~new_n31564_;
  assign new_n31566_ = pi0746 & new_n17433_;
  assign new_n31567_ = pi0038 & ~new_n31496_;
  assign new_n31568_ = ~new_n31566_ & new_n31567_;
  assign new_n31569_ = ~new_n31565_ & ~new_n31568_;
  assign new_n31570_ = new_n3272_ & ~new_n31569_;
  assign new_n31571_ = ~new_n31491_ & ~new_n31570_;
  assign new_n31572_ = ~new_n17590_ & ~new_n31571_;
  assign new_n31573_ = new_n17590_ & ~new_n31489_;
  assign new_n31574_ = ~new_n31572_ & ~new_n31573_;
  assign new_n31575_ = ~pi0785 & ~new_n31574_;
  assign new_n31576_ = ~new_n17591_ & ~new_n31489_;
  assign new_n31577_ = pi0609 & new_n31572_;
  assign new_n31578_ = ~new_n31576_ & ~new_n31577_;
  assign new_n31579_ = pi1155 & ~new_n31578_;
  assign new_n31580_ = ~new_n17603_ & ~new_n31489_;
  assign new_n31581_ = ~pi0609 & new_n31572_;
  assign new_n31582_ = ~new_n31580_ & ~new_n31581_;
  assign new_n31583_ = ~pi1155 & ~new_n31582_;
  assign new_n31584_ = ~new_n31579_ & ~new_n31583_;
  assign new_n31585_ = pi0785 & ~new_n31584_;
  assign new_n31586_ = ~new_n31575_ & ~new_n31585_;
  assign new_n31587_ = ~pi0781 & ~new_n31586_;
  assign new_n31588_ = pi0618 & new_n31586_;
  assign new_n31589_ = ~pi0618 & new_n31489_;
  assign new_n31590_ = pi1154 & ~new_n31589_;
  assign new_n31591_ = ~new_n31588_ & new_n31590_;
  assign new_n31592_ = ~pi0618 & new_n31586_;
  assign new_n31593_ = pi0618 & new_n31489_;
  assign new_n31594_ = ~pi1154 & ~new_n31593_;
  assign new_n31595_ = ~new_n31592_ & new_n31594_;
  assign new_n31596_ = ~new_n31591_ & ~new_n31595_;
  assign new_n31597_ = pi0781 & ~new_n31596_;
  assign new_n31598_ = ~new_n31587_ & ~new_n31597_;
  assign new_n31599_ = ~pi0789 & ~new_n31598_;
  assign new_n31600_ = pi0619 & new_n31598_;
  assign new_n31601_ = ~pi0619 & new_n31489_;
  assign new_n31602_ = pi1159 & ~new_n31601_;
  assign new_n31603_ = ~new_n31600_ & new_n31602_;
  assign new_n31604_ = ~pi0619 & new_n31598_;
  assign new_n31605_ = pi0619 & new_n31489_;
  assign new_n31606_ = ~pi1159 & ~new_n31605_;
  assign new_n31607_ = ~new_n31604_ & new_n31606_;
  assign new_n31608_ = ~new_n31603_ & ~new_n31607_;
  assign new_n31609_ = pi0789 & ~new_n31608_;
  assign new_n31610_ = ~new_n31599_ & ~new_n31609_;
  assign new_n31611_ = ~new_n17968_ & new_n31610_;
  assign new_n31612_ = new_n17968_ & new_n31489_;
  assign new_n31613_ = ~new_n31611_ & ~new_n31612_;
  assign new_n31614_ = ~new_n17762_ & ~new_n31613_;
  assign new_n31615_ = new_n17762_ & new_n31489_;
  assign new_n31616_ = ~new_n31614_ & ~new_n31615_;
  assign new_n31617_ = ~new_n17804_ & ~new_n31616_;
  assign new_n31618_ = new_n17804_ & new_n31489_;
  assign new_n31619_ = ~new_n31617_ & ~new_n31618_;
  assign new_n31620_ = pi0644 & ~new_n31619_;
  assign new_n31621_ = ~pi0644 & new_n31489_;
  assign new_n31622_ = ~pi0715 & ~new_n31621_;
  assign new_n31623_ = ~new_n31620_ & new_n31622_;
  assign new_n31624_ = pi1160 & ~new_n31623_;
  assign new_n31625_ = ~new_n31553_ & new_n31624_;
  assign new_n31626_ = pi0644 & ~new_n31551_;
  assign new_n31627_ = ~pi0715 & ~new_n31626_;
  assign new_n31628_ = ~pi0644 & ~new_n31619_;
  assign new_n31629_ = pi0644 & new_n31489_;
  assign new_n31630_ = pi0715 & ~new_n31629_;
  assign new_n31631_ = ~new_n31628_ & new_n31630_;
  assign new_n31632_ = ~pi1160 & ~new_n31631_;
  assign new_n31633_ = ~new_n31627_ & new_n31632_;
  assign new_n31634_ = ~new_n31625_ & ~new_n31633_;
  assign new_n31635_ = pi0790 & ~new_n31634_;
  assign new_n31636_ = pi0644 & new_n31624_;
  assign new_n31637_ = ~pi0644 & new_n31632_;
  assign new_n31638_ = pi0790 & ~new_n31637_;
  assign new_n31639_ = ~new_n31636_ & new_n31638_;
  assign new_n31640_ = ~new_n20567_ & new_n31613_;
  assign new_n31641_ = new_n17760_ & new_n31530_;
  assign new_n31642_ = new_n17759_ & new_n31534_;
  assign new_n31643_ = ~new_n31641_ & ~new_n31642_;
  assign new_n31644_ = ~new_n31640_ & new_n31643_;
  assign new_n31645_ = pi0792 & ~new_n31644_;
  assign new_n31646_ = ~pi0729 & new_n31569_;
  assign new_n31647_ = ~pi0191 & new_n16810_;
  assign new_n31648_ = pi0191 & new_n16928_;
  assign new_n31649_ = ~pi0746 & ~new_n31648_;
  assign new_n31650_ = ~new_n31647_ & new_n31649_;
  assign new_n31651_ = pi0191 & new_n17007_;
  assign new_n31652_ = ~pi0191 & ~new_n17074_;
  assign new_n31653_ = pi0746 & ~new_n31652_;
  assign new_n31654_ = ~new_n31651_ & new_n31653_;
  assign new_n31655_ = pi0039 & ~new_n31654_;
  assign new_n31656_ = ~new_n31650_ & new_n31655_;
  assign new_n31657_ = pi0191 & new_n17178_;
  assign new_n31658_ = ~pi0191 & new_n17217_;
  assign new_n31659_ = ~pi0746 & ~new_n31658_;
  assign new_n31660_ = ~new_n31657_ & new_n31659_;
  assign new_n31661_ = ~pi0191 & ~new_n17227_;
  assign new_n31662_ = pi0191 & ~new_n17234_;
  assign new_n31663_ = pi0746 & ~new_n31662_;
  assign new_n31664_ = ~new_n31661_ & new_n31663_;
  assign new_n31665_ = ~pi0039 & ~new_n31664_;
  assign new_n31666_ = ~new_n31660_ & new_n31665_;
  assign new_n31667_ = ~pi0038 & ~new_n31666_;
  assign new_n31668_ = ~new_n31656_ & new_n31667_;
  assign new_n31669_ = ~pi0746 & new_n24079_;
  assign new_n31670_ = ~new_n17035_ & ~new_n31669_;
  assign new_n31671_ = ~pi0039 & ~new_n31670_;
  assign new_n31672_ = ~pi0191 & ~new_n31671_;
  assign new_n31673_ = ~new_n16916_ & ~new_n31302_;
  assign new_n31674_ = pi0191 & ~new_n31673_;
  assign new_n31675_ = new_n6257_ & new_n31674_;
  assign new_n31676_ = pi0038 & ~new_n31675_;
  assign new_n31677_ = ~new_n31672_ & new_n31676_;
  assign new_n31678_ = pi0729 & ~new_n31677_;
  assign new_n31679_ = ~new_n31668_ & new_n31678_;
  assign new_n31680_ = new_n3272_ & ~new_n31679_;
  assign new_n31681_ = ~new_n31646_ & new_n31680_;
  assign new_n31682_ = ~new_n31491_ & ~new_n31681_;
  assign new_n31683_ = ~pi0625 & new_n31682_;
  assign new_n31684_ = pi0625 & new_n31571_;
  assign new_n31685_ = ~pi1153 & ~new_n31684_;
  assign new_n31686_ = ~new_n31683_ & new_n31685_;
  assign new_n31687_ = ~pi0608 & ~new_n31509_;
  assign new_n31688_ = ~new_n31686_ & new_n31687_;
  assign new_n31689_ = pi0625 & new_n31682_;
  assign new_n31690_ = ~pi0625 & new_n31571_;
  assign new_n31691_ = pi1153 & ~new_n31690_;
  assign new_n31692_ = ~new_n31689_ & new_n31691_;
  assign new_n31693_ = pi0608 & ~new_n31513_;
  assign new_n31694_ = ~new_n31692_ & new_n31693_;
  assign new_n31695_ = ~new_n31688_ & ~new_n31694_;
  assign new_n31696_ = pi0778 & ~new_n31695_;
  assign new_n31697_ = ~pi0778 & new_n31682_;
  assign new_n31698_ = ~new_n31696_ & ~new_n31697_;
  assign new_n31699_ = ~pi0609 & ~new_n31698_;
  assign new_n31700_ = pi0609 & new_n31516_;
  assign new_n31701_ = ~pi1155 & ~new_n31700_;
  assign new_n31702_ = ~new_n31699_ & new_n31701_;
  assign new_n31703_ = ~pi0660 & ~new_n31579_;
  assign new_n31704_ = ~new_n31702_ & new_n31703_;
  assign new_n31705_ = pi0609 & ~new_n31698_;
  assign new_n31706_ = ~pi0609 & new_n31516_;
  assign new_n31707_ = pi1155 & ~new_n31706_;
  assign new_n31708_ = ~new_n31705_ & new_n31707_;
  assign new_n31709_ = pi0660 & ~new_n31583_;
  assign new_n31710_ = ~new_n31708_ & new_n31709_;
  assign new_n31711_ = ~new_n31704_ & ~new_n31710_;
  assign new_n31712_ = pi0785 & ~new_n31711_;
  assign new_n31713_ = ~pi0785 & ~new_n31698_;
  assign new_n31714_ = ~new_n31712_ & ~new_n31713_;
  assign new_n31715_ = ~pi0618 & ~new_n31714_;
  assign new_n31716_ = pi0618 & new_n31519_;
  assign new_n31717_ = ~pi1154 & ~new_n31716_;
  assign new_n31718_ = ~new_n31715_ & new_n31717_;
  assign new_n31719_ = ~pi0627 & ~new_n31591_;
  assign new_n31720_ = ~new_n31718_ & new_n31719_;
  assign new_n31721_ = pi0618 & ~new_n31714_;
  assign new_n31722_ = ~pi0618 & new_n31519_;
  assign new_n31723_ = pi1154 & ~new_n31722_;
  assign new_n31724_ = ~new_n31721_ & new_n31723_;
  assign new_n31725_ = pi0627 & ~new_n31595_;
  assign new_n31726_ = ~new_n31724_ & new_n31725_;
  assign new_n31727_ = ~new_n31720_ & ~new_n31726_;
  assign new_n31728_ = pi0781 & ~new_n31727_;
  assign new_n31729_ = ~pi0781 & ~new_n31714_;
  assign new_n31730_ = ~new_n31728_ & ~new_n31729_;
  assign new_n31731_ = pi0619 & ~new_n31730_;
  assign new_n31732_ = ~pi0619 & ~new_n31522_;
  assign new_n31733_ = pi1159 & ~new_n31732_;
  assign new_n31734_ = ~new_n31731_ & new_n31733_;
  assign new_n31735_ = pi0648 & ~new_n31607_;
  assign new_n31736_ = ~new_n31734_ & new_n31735_;
  assign new_n31737_ = ~pi0619 & ~new_n31730_;
  assign new_n31738_ = pi0619 & ~new_n31522_;
  assign new_n31739_ = ~pi1159 & ~new_n31738_;
  assign new_n31740_ = ~new_n31737_ & new_n31739_;
  assign new_n31741_ = ~pi0648 & ~new_n31603_;
  assign new_n31742_ = ~new_n31740_ & new_n31741_;
  assign new_n31743_ = pi0789 & ~new_n31742_;
  assign new_n31744_ = ~new_n31736_ & new_n31743_;
  assign new_n31745_ = ~pi0789 & new_n31730_;
  assign new_n31746_ = new_n17969_ & ~new_n31745_;
  assign new_n31747_ = ~new_n31744_ & new_n31746_;
  assign new_n31748_ = pi0626 & ~new_n31610_;
  assign new_n31749_ = ~pi0626 & ~new_n31489_;
  assign new_n31750_ = new_n17731_ & ~new_n31749_;
  assign new_n31751_ = ~new_n31748_ & new_n31750_;
  assign new_n31752_ = new_n17856_ & new_n31524_;
  assign new_n31753_ = ~pi0626 & ~new_n31610_;
  assign new_n31754_ = pi0626 & ~new_n31489_;
  assign new_n31755_ = new_n17732_ & ~new_n31754_;
  assign new_n31756_ = ~new_n31753_ & new_n31755_;
  assign new_n31757_ = ~new_n31752_ & ~new_n31756_;
  assign new_n31758_ = ~new_n31751_ & new_n31757_;
  assign new_n31759_ = pi0788 & ~new_n31758_;
  assign new_n31760_ = ~new_n20364_ & ~new_n31759_;
  assign new_n31761_ = ~new_n31747_ & new_n31760_;
  assign new_n31762_ = ~new_n31645_ & ~new_n31761_;
  assign new_n31763_ = ~new_n20360_ & ~new_n31762_;
  assign new_n31764_ = new_n17801_ & new_n31546_;
  assign new_n31765_ = new_n17802_ & new_n31542_;
  assign new_n31766_ = ~new_n20556_ & new_n31616_;
  assign new_n31767_ = ~new_n31765_ & ~new_n31766_;
  assign new_n31768_ = ~new_n31764_ & new_n31767_;
  assign new_n31769_ = pi0787 & ~new_n31768_;
  assign new_n31770_ = ~new_n31763_ & ~new_n31769_;
  assign new_n31771_ = ~new_n31639_ & new_n31770_;
  assign new_n31772_ = ~new_n31635_ & ~new_n31771_;
  assign new_n31773_ = ~po1038 & ~new_n31772_;
  assign new_n31774_ = ~pi0191 & po1038;
  assign new_n31775_ = ~pi0832 & ~new_n31774_;
  assign new_n31776_ = ~new_n31773_ & new_n31775_;
  assign po0348 = ~new_n31488_ & ~new_n31776_;
  assign new_n31778_ = ~pi0192 & ~new_n2754_;
  assign new_n31779_ = pi0764 & new_n16913_;
  assign new_n31780_ = ~new_n31778_ & ~new_n31779_;
  assign new_n31781_ = ~new_n17858_ & ~new_n31780_;
  assign new_n31782_ = ~pi0785 & ~new_n31781_;
  assign new_n31783_ = new_n17603_ & new_n31779_;
  assign new_n31784_ = new_n31781_ & ~new_n31783_;
  assign new_n31785_ = pi1155 & ~new_n31784_;
  assign new_n31786_ = ~pi1155 & ~new_n31778_;
  assign new_n31787_ = ~new_n31783_ & new_n31786_;
  assign new_n31788_ = ~new_n31785_ & ~new_n31787_;
  assign new_n31789_ = pi0785 & ~new_n31788_;
  assign new_n31790_ = ~new_n31782_ & ~new_n31789_;
  assign new_n31791_ = ~pi0781 & ~new_n31790_;
  assign new_n31792_ = ~new_n17873_ & new_n31790_;
  assign new_n31793_ = pi1154 & ~new_n31792_;
  assign new_n31794_ = ~new_n17876_ & new_n31790_;
  assign new_n31795_ = ~pi1154 & ~new_n31794_;
  assign new_n31796_ = ~new_n31793_ & ~new_n31795_;
  assign new_n31797_ = pi0781 & ~new_n31796_;
  assign new_n31798_ = ~new_n31791_ & ~new_n31797_;
  assign new_n31799_ = ~pi0789 & ~new_n31798_;
  assign new_n31800_ = ~new_n23057_ & new_n31798_;
  assign new_n31801_ = pi1159 & ~new_n31800_;
  assign new_n31802_ = ~new_n23060_ & new_n31798_;
  assign new_n31803_ = ~pi1159 & ~new_n31802_;
  assign new_n31804_ = ~new_n31801_ & ~new_n31803_;
  assign new_n31805_ = pi0789 & ~new_n31804_;
  assign new_n31806_ = ~new_n31799_ & ~new_n31805_;
  assign new_n31807_ = ~new_n17968_ & new_n31806_;
  assign new_n31808_ = new_n17968_ & new_n31778_;
  assign new_n31809_ = ~new_n31807_ & ~new_n31808_;
  assign new_n31810_ = ~new_n17762_ & ~new_n31809_;
  assign new_n31811_ = new_n17762_ & new_n31778_;
  assign new_n31812_ = ~new_n31810_ & ~new_n31811_;
  assign new_n31813_ = ~new_n20556_ & new_n31812_;
  assign new_n31814_ = pi0691 & new_n16915_;
  assign new_n31815_ = ~new_n31778_ & ~new_n31814_;
  assign new_n31816_ = ~pi0778 & ~new_n31815_;
  assign new_n31817_ = ~pi0625 & new_n31814_;
  assign new_n31818_ = ~new_n31815_ & ~new_n31817_;
  assign new_n31819_ = pi1153 & ~new_n31818_;
  assign new_n31820_ = ~pi1153 & ~new_n31778_;
  assign new_n31821_ = ~new_n31817_ & new_n31820_;
  assign new_n31822_ = pi0778 & ~new_n31821_;
  assign new_n31823_ = ~new_n31819_ & new_n31822_;
  assign new_n31824_ = ~new_n31816_ & ~new_n31823_;
  assign new_n31825_ = ~new_n17844_ & ~new_n31824_;
  assign new_n31826_ = ~new_n17846_ & new_n31825_;
  assign new_n31827_ = ~new_n17848_ & new_n31826_;
  assign new_n31828_ = ~new_n17980_ & new_n31827_;
  assign new_n31829_ = ~new_n18011_ & new_n31828_;
  assign new_n31830_ = ~pi0647 & new_n31829_;
  assign new_n31831_ = pi0647 & new_n31778_;
  assign new_n31832_ = ~pi1157 & ~new_n31831_;
  assign new_n31833_ = ~new_n31830_ & new_n31832_;
  assign new_n31834_ = pi0630 & new_n31833_;
  assign new_n31835_ = pi0647 & ~new_n31829_;
  assign new_n31836_ = ~pi0647 & ~new_n31778_;
  assign new_n31837_ = ~new_n31835_ & ~new_n31836_;
  assign new_n31838_ = new_n17801_ & ~new_n31837_;
  assign new_n31839_ = ~new_n31834_ & ~new_n31838_;
  assign new_n31840_ = ~new_n31813_ & new_n31839_;
  assign new_n31841_ = pi0787 & ~new_n31840_;
  assign new_n31842_ = pi0626 & ~new_n31806_;
  assign new_n31843_ = ~pi0626 & ~new_n31778_;
  assign new_n31844_ = new_n17731_ & ~new_n31843_;
  assign new_n31845_ = ~new_n31842_ & new_n31844_;
  assign new_n31846_ = new_n17856_ & new_n31827_;
  assign new_n31847_ = ~pi0626 & ~new_n31806_;
  assign new_n31848_ = pi0626 & ~new_n31778_;
  assign new_n31849_ = new_n17732_ & ~new_n31848_;
  assign new_n31850_ = ~new_n31847_ & new_n31849_;
  assign new_n31851_ = ~new_n31846_ & ~new_n31850_;
  assign new_n31852_ = ~new_n31845_ & new_n31851_;
  assign new_n31853_ = pi0788 & ~new_n31852_;
  assign new_n31854_ = ~new_n16639_ & ~new_n31815_;
  assign new_n31855_ = pi0625 & new_n31854_;
  assign new_n31856_ = new_n31780_ & ~new_n31854_;
  assign new_n31857_ = ~new_n31855_ & ~new_n31856_;
  assign new_n31858_ = new_n31820_ & ~new_n31857_;
  assign new_n31859_ = ~pi0608 & ~new_n31819_;
  assign new_n31860_ = ~new_n31858_ & new_n31859_;
  assign new_n31861_ = pi1153 & new_n31780_;
  assign new_n31862_ = ~new_n31855_ & new_n31861_;
  assign new_n31863_ = pi0608 & ~new_n31821_;
  assign new_n31864_ = ~new_n31862_ & new_n31863_;
  assign new_n31865_ = ~new_n31860_ & ~new_n31864_;
  assign new_n31866_ = pi0778 & ~new_n31865_;
  assign new_n31867_ = ~pi0778 & ~new_n31856_;
  assign new_n31868_ = ~new_n31866_ & ~new_n31867_;
  assign new_n31869_ = ~pi0609 & ~new_n31868_;
  assign new_n31870_ = pi0609 & ~new_n31824_;
  assign new_n31871_ = ~pi1155 & ~new_n31870_;
  assign new_n31872_ = ~new_n31869_ & new_n31871_;
  assign new_n31873_ = ~pi0660 & ~new_n31785_;
  assign new_n31874_ = ~new_n31872_ & new_n31873_;
  assign new_n31875_ = pi0609 & ~new_n31868_;
  assign new_n31876_ = ~pi0609 & ~new_n31824_;
  assign new_n31877_ = pi1155 & ~new_n31876_;
  assign new_n31878_ = ~new_n31875_ & new_n31877_;
  assign new_n31879_ = pi0660 & ~new_n31787_;
  assign new_n31880_ = ~new_n31878_ & new_n31879_;
  assign new_n31881_ = ~new_n31874_ & ~new_n31880_;
  assign new_n31882_ = pi0785 & ~new_n31881_;
  assign new_n31883_ = ~pi0785 & ~new_n31868_;
  assign new_n31884_ = ~new_n31882_ & ~new_n31883_;
  assign new_n31885_ = ~pi0618 & ~new_n31884_;
  assign new_n31886_ = pi0618 & new_n31825_;
  assign new_n31887_ = ~pi1154 & ~new_n31886_;
  assign new_n31888_ = ~new_n31885_ & new_n31887_;
  assign new_n31889_ = ~pi0627 & ~new_n31793_;
  assign new_n31890_ = ~new_n31888_ & new_n31889_;
  assign new_n31891_ = pi0618 & ~new_n31884_;
  assign new_n31892_ = ~pi0618 & new_n31825_;
  assign new_n31893_ = pi1154 & ~new_n31892_;
  assign new_n31894_ = ~new_n31891_ & new_n31893_;
  assign new_n31895_ = pi0627 & ~new_n31795_;
  assign new_n31896_ = ~new_n31894_ & new_n31895_;
  assign new_n31897_ = ~new_n31890_ & ~new_n31896_;
  assign new_n31898_ = pi0781 & ~new_n31897_;
  assign new_n31899_ = ~pi0781 & ~new_n31884_;
  assign new_n31900_ = ~new_n31898_ & ~new_n31899_;
  assign new_n31901_ = pi0619 & ~new_n31900_;
  assign new_n31902_ = ~pi0619 & new_n31826_;
  assign new_n31903_ = pi1159 & ~new_n31902_;
  assign new_n31904_ = ~new_n31901_ & new_n31903_;
  assign new_n31905_ = pi0648 & ~new_n31803_;
  assign new_n31906_ = ~new_n31904_ & new_n31905_;
  assign new_n31907_ = ~pi0619 & ~new_n31900_;
  assign new_n31908_ = pi0619 & new_n31826_;
  assign new_n31909_ = ~pi1159 & ~new_n31908_;
  assign new_n31910_ = ~new_n31907_ & new_n31909_;
  assign new_n31911_ = ~pi0648 & ~new_n31801_;
  assign new_n31912_ = ~new_n31910_ & new_n31911_;
  assign new_n31913_ = pi0789 & ~new_n31912_;
  assign new_n31914_ = ~new_n31906_ & new_n31913_;
  assign new_n31915_ = ~pi0789 & new_n31900_;
  assign new_n31916_ = new_n17969_ & ~new_n31915_;
  assign new_n31917_ = ~new_n31914_ & new_n31916_;
  assign new_n31918_ = ~new_n31853_ & ~new_n31917_;
  assign new_n31919_ = ~new_n20364_ & ~new_n31918_;
  assign new_n31920_ = new_n18008_ & ~new_n31809_;
  assign new_n31921_ = new_n20851_ & new_n31828_;
  assign new_n31922_ = ~new_n31920_ & ~new_n31921_;
  assign new_n31923_ = ~pi0629 & ~new_n31922_;
  assign new_n31924_ = new_n20855_ & new_n31828_;
  assign new_n31925_ = new_n18007_ & ~new_n31809_;
  assign new_n31926_ = ~new_n31924_ & ~new_n31925_;
  assign new_n31927_ = pi0629 & ~new_n31926_;
  assign new_n31928_ = ~new_n31923_ & ~new_n31927_;
  assign new_n31929_ = pi0792 & ~new_n31928_;
  assign new_n31930_ = ~new_n20360_ & ~new_n31929_;
  assign new_n31931_ = ~new_n31919_ & new_n31930_;
  assign new_n31932_ = ~new_n31841_ & ~new_n31931_;
  assign new_n31933_ = pi0644 & new_n31932_;
  assign new_n31934_ = ~pi0787 & ~new_n31829_;
  assign new_n31935_ = pi1157 & ~new_n31837_;
  assign new_n31936_ = ~new_n31833_ & ~new_n31935_;
  assign new_n31937_ = pi0787 & ~new_n31936_;
  assign new_n31938_ = ~new_n31934_ & ~new_n31937_;
  assign new_n31939_ = ~pi0644 & new_n31938_;
  assign new_n31940_ = pi0715 & ~new_n31939_;
  assign new_n31941_ = ~new_n31933_ & new_n31940_;
  assign new_n31942_ = ~new_n17804_ & ~new_n31812_;
  assign new_n31943_ = new_n17804_ & new_n31778_;
  assign new_n31944_ = ~new_n31942_ & ~new_n31943_;
  assign new_n31945_ = pi0644 & ~new_n31944_;
  assign new_n31946_ = ~pi0644 & new_n31778_;
  assign new_n31947_ = ~pi0715 & ~new_n31946_;
  assign new_n31948_ = ~new_n31945_ & new_n31947_;
  assign new_n31949_ = pi1160 & ~new_n31948_;
  assign new_n31950_ = ~new_n31941_ & new_n31949_;
  assign new_n31951_ = ~pi0644 & new_n31932_;
  assign new_n31952_ = pi0644 & new_n31938_;
  assign new_n31953_ = ~pi0715 & ~new_n31952_;
  assign new_n31954_ = ~new_n31951_ & new_n31953_;
  assign new_n31955_ = ~pi0644 & ~new_n31944_;
  assign new_n31956_ = pi0644 & new_n31778_;
  assign new_n31957_ = pi0715 & ~new_n31956_;
  assign new_n31958_ = ~new_n31955_ & new_n31957_;
  assign new_n31959_ = ~pi1160 & ~new_n31958_;
  assign new_n31960_ = ~new_n31954_ & new_n31959_;
  assign new_n31961_ = ~new_n31950_ & ~new_n31960_;
  assign new_n31962_ = pi0790 & ~new_n31961_;
  assign new_n31963_ = ~pi0790 & new_n31932_;
  assign new_n31964_ = pi0832 & ~new_n31963_;
  assign new_n31965_ = ~new_n31962_ & new_n31964_;
  assign new_n31966_ = ~pi0192 & ~new_n17558_;
  assign new_n31967_ = new_n17691_ & ~new_n31966_;
  assign new_n31968_ = pi0192 & ~new_n3272_;
  assign new_n31969_ = ~pi0192 & new_n18124_;
  assign new_n31970_ = pi0192 & ~new_n18128_;
  assign new_n31971_ = ~pi0038 & ~new_n31970_;
  assign new_n31972_ = ~new_n31969_ & new_n31971_;
  assign new_n31973_ = ~pi0192 & ~new_n17431_;
  assign new_n31974_ = new_n17544_ & ~new_n31973_;
  assign new_n31975_ = pi0691 & ~new_n31974_;
  assign new_n31976_ = ~new_n31972_ & new_n31975_;
  assign new_n31977_ = ~pi0192 & ~pi0691;
  assign new_n31978_ = ~new_n17551_ & new_n31977_;
  assign new_n31979_ = new_n3272_ & ~new_n31978_;
  assign new_n31980_ = ~new_n31976_ & new_n31979_;
  assign new_n31981_ = ~new_n31968_ & ~new_n31980_;
  assign new_n31982_ = ~pi0778 & ~new_n31981_;
  assign new_n31983_ = pi0625 & new_n31981_;
  assign new_n31984_ = ~pi0625 & new_n31966_;
  assign new_n31985_ = pi1153 & ~new_n31984_;
  assign new_n31986_ = ~new_n31983_ & new_n31985_;
  assign new_n31987_ = ~pi0625 & new_n31981_;
  assign new_n31988_ = pi0625 & new_n31966_;
  assign new_n31989_ = ~pi1153 & ~new_n31988_;
  assign new_n31990_ = ~new_n31987_ & new_n31989_;
  assign new_n31991_ = ~new_n31986_ & ~new_n31990_;
  assign new_n31992_ = pi0778 & ~new_n31991_;
  assign new_n31993_ = ~new_n31982_ & ~new_n31992_;
  assign new_n31994_ = ~new_n17618_ & ~new_n31993_;
  assign new_n31995_ = new_n17618_ & ~new_n31966_;
  assign new_n31996_ = ~new_n31994_ & ~new_n31995_;
  assign new_n31997_ = ~new_n17655_ & new_n31996_;
  assign new_n31998_ = new_n17655_ & new_n31966_;
  assign new_n31999_ = ~new_n31997_ & ~new_n31998_;
  assign new_n32000_ = ~new_n17691_ & new_n31999_;
  assign new_n32001_ = ~new_n31967_ & ~new_n32000_;
  assign new_n32002_ = ~new_n17734_ & new_n32001_;
  assign new_n32003_ = new_n17734_ & new_n31966_;
  assign new_n32004_ = ~new_n32002_ & ~new_n32003_;
  assign new_n32005_ = ~pi0628 & ~new_n32004_;
  assign new_n32006_ = pi0628 & new_n31966_;
  assign new_n32007_ = ~new_n32005_ & ~new_n32006_;
  assign new_n32008_ = ~pi1156 & ~new_n32007_;
  assign new_n32009_ = pi0628 & ~new_n32004_;
  assign new_n32010_ = ~pi0628 & new_n31966_;
  assign new_n32011_ = ~new_n32009_ & ~new_n32010_;
  assign new_n32012_ = pi1156 & ~new_n32011_;
  assign new_n32013_ = ~new_n32008_ & ~new_n32012_;
  assign new_n32014_ = pi0792 & ~new_n32013_;
  assign new_n32015_ = ~pi0792 & ~new_n32004_;
  assign new_n32016_ = ~new_n32014_ & ~new_n32015_;
  assign new_n32017_ = ~pi0647 & ~new_n32016_;
  assign new_n32018_ = pi0647 & new_n31966_;
  assign new_n32019_ = ~new_n32017_ & ~new_n32018_;
  assign new_n32020_ = ~pi1157 & ~new_n32019_;
  assign new_n32021_ = pi0647 & ~new_n32016_;
  assign new_n32022_ = ~pi0647 & new_n31966_;
  assign new_n32023_ = ~new_n32021_ & ~new_n32022_;
  assign new_n32024_ = pi1157 & ~new_n32023_;
  assign new_n32025_ = ~new_n32020_ & ~new_n32024_;
  assign new_n32026_ = pi0787 & ~new_n32025_;
  assign new_n32027_ = ~pi0787 & ~new_n32016_;
  assign new_n32028_ = ~new_n32026_ & ~new_n32027_;
  assign new_n32029_ = ~pi0644 & ~new_n32028_;
  assign new_n32030_ = pi0715 & ~new_n32029_;
  assign new_n32031_ = ~pi0764 & new_n17347_;
  assign new_n32032_ = pi0192 & new_n17424_;
  assign new_n32033_ = ~new_n32031_ & ~new_n32032_;
  assign new_n32034_ = pi0039 & ~new_n32033_;
  assign new_n32035_ = ~pi0192 & pi0764;
  assign new_n32036_ = new_n17393_ & new_n32035_;
  assign new_n32037_ = pi0764 & ~new_n17397_;
  assign new_n32038_ = pi0192 & ~new_n32037_;
  assign new_n32039_ = ~new_n22598_ & ~new_n32038_;
  assign new_n32040_ = ~new_n32036_ & new_n32039_;
  assign new_n32041_ = ~new_n32034_ & new_n32040_;
  assign new_n32042_ = ~pi0038 & ~new_n32041_;
  assign new_n32043_ = pi0764 & new_n17433_;
  assign new_n32044_ = pi0038 & ~new_n31973_;
  assign new_n32045_ = ~new_n32043_ & new_n32044_;
  assign new_n32046_ = ~new_n32042_ & ~new_n32045_;
  assign new_n32047_ = new_n3272_ & ~new_n32046_;
  assign new_n32048_ = ~new_n31968_ & ~new_n32047_;
  assign new_n32049_ = ~new_n17590_ & ~new_n32048_;
  assign new_n32050_ = new_n17590_ & ~new_n31966_;
  assign new_n32051_ = ~new_n32049_ & ~new_n32050_;
  assign new_n32052_ = ~pi0785 & ~new_n32051_;
  assign new_n32053_ = ~new_n17591_ & ~new_n31966_;
  assign new_n32054_ = pi0609 & new_n32049_;
  assign new_n32055_ = ~new_n32053_ & ~new_n32054_;
  assign new_n32056_ = pi1155 & ~new_n32055_;
  assign new_n32057_ = ~new_n17603_ & ~new_n31966_;
  assign new_n32058_ = ~pi0609 & new_n32049_;
  assign new_n32059_ = ~new_n32057_ & ~new_n32058_;
  assign new_n32060_ = ~pi1155 & ~new_n32059_;
  assign new_n32061_ = ~new_n32056_ & ~new_n32060_;
  assign new_n32062_ = pi0785 & ~new_n32061_;
  assign new_n32063_ = ~new_n32052_ & ~new_n32062_;
  assign new_n32064_ = ~pi0781 & ~new_n32063_;
  assign new_n32065_ = pi0618 & new_n32063_;
  assign new_n32066_ = ~pi0618 & new_n31966_;
  assign new_n32067_ = pi1154 & ~new_n32066_;
  assign new_n32068_ = ~new_n32065_ & new_n32067_;
  assign new_n32069_ = ~pi0618 & new_n32063_;
  assign new_n32070_ = pi0618 & new_n31966_;
  assign new_n32071_ = ~pi1154 & ~new_n32070_;
  assign new_n32072_ = ~new_n32069_ & new_n32071_;
  assign new_n32073_ = ~new_n32068_ & ~new_n32072_;
  assign new_n32074_ = pi0781 & ~new_n32073_;
  assign new_n32075_ = ~new_n32064_ & ~new_n32074_;
  assign new_n32076_ = ~pi0789 & ~new_n32075_;
  assign new_n32077_ = pi0619 & new_n32075_;
  assign new_n32078_ = ~pi0619 & new_n31966_;
  assign new_n32079_ = pi1159 & ~new_n32078_;
  assign new_n32080_ = ~new_n32077_ & new_n32079_;
  assign new_n32081_ = ~pi0619 & new_n32075_;
  assign new_n32082_ = pi0619 & new_n31966_;
  assign new_n32083_ = ~pi1159 & ~new_n32082_;
  assign new_n32084_ = ~new_n32081_ & new_n32083_;
  assign new_n32085_ = ~new_n32080_ & ~new_n32084_;
  assign new_n32086_ = pi0789 & ~new_n32085_;
  assign new_n32087_ = ~new_n32076_ & ~new_n32086_;
  assign new_n32088_ = ~new_n17968_ & new_n32087_;
  assign new_n32089_ = new_n17968_ & new_n31966_;
  assign new_n32090_ = ~new_n32088_ & ~new_n32089_;
  assign new_n32091_ = ~new_n17762_ & ~new_n32090_;
  assign new_n32092_ = new_n17762_ & new_n31966_;
  assign new_n32093_ = ~new_n32091_ & ~new_n32092_;
  assign new_n32094_ = ~new_n17804_ & ~new_n32093_;
  assign new_n32095_ = new_n17804_ & new_n31966_;
  assign new_n32096_ = ~new_n32094_ & ~new_n32095_;
  assign new_n32097_ = pi0644 & ~new_n32096_;
  assign new_n32098_ = ~pi0644 & new_n31966_;
  assign new_n32099_ = ~pi0715 & ~new_n32098_;
  assign new_n32100_ = ~new_n32097_ & new_n32099_;
  assign new_n32101_ = pi1160 & ~new_n32100_;
  assign new_n32102_ = ~new_n32030_ & new_n32101_;
  assign new_n32103_ = pi0644 & ~new_n32028_;
  assign new_n32104_ = ~pi0715 & ~new_n32103_;
  assign new_n32105_ = ~pi0644 & ~new_n32096_;
  assign new_n32106_ = pi0644 & new_n31966_;
  assign new_n32107_ = pi0715 & ~new_n32106_;
  assign new_n32108_ = ~new_n32105_ & new_n32107_;
  assign new_n32109_ = ~pi1160 & ~new_n32108_;
  assign new_n32110_ = ~new_n32104_ & new_n32109_;
  assign new_n32111_ = ~new_n32102_ & ~new_n32110_;
  assign new_n32112_ = pi0790 & ~new_n32111_;
  assign new_n32113_ = pi0644 & new_n32101_;
  assign new_n32114_ = ~pi0644 & new_n32109_;
  assign new_n32115_ = pi0790 & ~new_n32114_;
  assign new_n32116_ = ~new_n32113_ & new_n32115_;
  assign new_n32117_ = ~new_n20567_ & new_n32090_;
  assign new_n32118_ = new_n17760_ & new_n32007_;
  assign new_n32119_ = new_n17759_ & new_n32011_;
  assign new_n32120_ = ~new_n32118_ & ~new_n32119_;
  assign new_n32121_ = ~new_n32117_ & new_n32120_;
  assign new_n32122_ = pi0792 & ~new_n32121_;
  assign new_n32123_ = ~pi0691 & new_n32046_;
  assign new_n32124_ = ~pi0192 & new_n16810_;
  assign new_n32125_ = pi0192 & new_n16928_;
  assign new_n32126_ = ~pi0764 & ~new_n32125_;
  assign new_n32127_ = ~new_n32124_ & new_n32126_;
  assign new_n32128_ = pi0192 & new_n17007_;
  assign new_n32129_ = ~pi0192 & ~new_n17074_;
  assign new_n32130_ = pi0764 & ~new_n32129_;
  assign new_n32131_ = ~new_n32128_ & new_n32130_;
  assign new_n32132_ = pi0039 & ~new_n32131_;
  assign new_n32133_ = ~new_n32127_ & new_n32132_;
  assign new_n32134_ = pi0192 & new_n17178_;
  assign new_n32135_ = ~pi0192 & new_n17217_;
  assign new_n32136_ = ~pi0764 & ~new_n32135_;
  assign new_n32137_ = ~new_n32134_ & new_n32136_;
  assign new_n32138_ = ~pi0192 & ~new_n17227_;
  assign new_n32139_ = pi0192 & ~new_n17234_;
  assign new_n32140_ = pi0764 & ~new_n32139_;
  assign new_n32141_ = ~new_n32138_ & new_n32140_;
  assign new_n32142_ = ~pi0039 & ~new_n32141_;
  assign new_n32143_ = ~new_n32137_ & new_n32142_;
  assign new_n32144_ = ~pi0038 & ~new_n32143_;
  assign new_n32145_ = ~new_n32133_ & new_n32144_;
  assign new_n32146_ = ~pi0764 & new_n24079_;
  assign new_n32147_ = ~new_n17035_ & ~new_n32146_;
  assign new_n32148_ = ~pi0039 & ~new_n32147_;
  assign new_n32149_ = ~pi0192 & ~new_n32148_;
  assign new_n32150_ = ~new_n16916_ & ~new_n31779_;
  assign new_n32151_ = pi0192 & ~new_n32150_;
  assign new_n32152_ = new_n6257_ & new_n32151_;
  assign new_n32153_ = pi0038 & ~new_n32152_;
  assign new_n32154_ = ~new_n32149_ & new_n32153_;
  assign new_n32155_ = pi0691 & ~new_n32154_;
  assign new_n32156_ = ~new_n32145_ & new_n32155_;
  assign new_n32157_ = new_n3272_ & ~new_n32156_;
  assign new_n32158_ = ~new_n32123_ & new_n32157_;
  assign new_n32159_ = ~new_n31968_ & ~new_n32158_;
  assign new_n32160_ = ~pi0625 & new_n32159_;
  assign new_n32161_ = pi0625 & new_n32048_;
  assign new_n32162_ = ~pi1153 & ~new_n32161_;
  assign new_n32163_ = ~new_n32160_ & new_n32162_;
  assign new_n32164_ = ~pi0608 & ~new_n31986_;
  assign new_n32165_ = ~new_n32163_ & new_n32164_;
  assign new_n32166_ = pi0625 & new_n32159_;
  assign new_n32167_ = ~pi0625 & new_n32048_;
  assign new_n32168_ = pi1153 & ~new_n32167_;
  assign new_n32169_ = ~new_n32166_ & new_n32168_;
  assign new_n32170_ = pi0608 & ~new_n31990_;
  assign new_n32171_ = ~new_n32169_ & new_n32170_;
  assign new_n32172_ = ~new_n32165_ & ~new_n32171_;
  assign new_n32173_ = pi0778 & ~new_n32172_;
  assign new_n32174_ = ~pi0778 & new_n32159_;
  assign new_n32175_ = ~new_n32173_ & ~new_n32174_;
  assign new_n32176_ = ~pi0609 & ~new_n32175_;
  assign new_n32177_ = pi0609 & new_n31993_;
  assign new_n32178_ = ~pi1155 & ~new_n32177_;
  assign new_n32179_ = ~new_n32176_ & new_n32178_;
  assign new_n32180_ = ~pi0660 & ~new_n32056_;
  assign new_n32181_ = ~new_n32179_ & new_n32180_;
  assign new_n32182_ = pi0609 & ~new_n32175_;
  assign new_n32183_ = ~pi0609 & new_n31993_;
  assign new_n32184_ = pi1155 & ~new_n32183_;
  assign new_n32185_ = ~new_n32182_ & new_n32184_;
  assign new_n32186_ = pi0660 & ~new_n32060_;
  assign new_n32187_ = ~new_n32185_ & new_n32186_;
  assign new_n32188_ = ~new_n32181_ & ~new_n32187_;
  assign new_n32189_ = pi0785 & ~new_n32188_;
  assign new_n32190_ = ~pi0785 & ~new_n32175_;
  assign new_n32191_ = ~new_n32189_ & ~new_n32190_;
  assign new_n32192_ = ~pi0618 & ~new_n32191_;
  assign new_n32193_ = pi0618 & new_n31996_;
  assign new_n32194_ = ~pi1154 & ~new_n32193_;
  assign new_n32195_ = ~new_n32192_ & new_n32194_;
  assign new_n32196_ = ~pi0627 & ~new_n32068_;
  assign new_n32197_ = ~new_n32195_ & new_n32196_;
  assign new_n32198_ = pi0618 & ~new_n32191_;
  assign new_n32199_ = ~pi0618 & new_n31996_;
  assign new_n32200_ = pi1154 & ~new_n32199_;
  assign new_n32201_ = ~new_n32198_ & new_n32200_;
  assign new_n32202_ = pi0627 & ~new_n32072_;
  assign new_n32203_ = ~new_n32201_ & new_n32202_;
  assign new_n32204_ = ~new_n32197_ & ~new_n32203_;
  assign new_n32205_ = pi0781 & ~new_n32204_;
  assign new_n32206_ = ~pi0781 & ~new_n32191_;
  assign new_n32207_ = ~new_n32205_ & ~new_n32206_;
  assign new_n32208_ = pi0619 & ~new_n32207_;
  assign new_n32209_ = ~pi0619 & ~new_n31999_;
  assign new_n32210_ = pi1159 & ~new_n32209_;
  assign new_n32211_ = ~new_n32208_ & new_n32210_;
  assign new_n32212_ = pi0648 & ~new_n32084_;
  assign new_n32213_ = ~new_n32211_ & new_n32212_;
  assign new_n32214_ = ~pi0619 & ~new_n32207_;
  assign new_n32215_ = pi0619 & ~new_n31999_;
  assign new_n32216_ = ~pi1159 & ~new_n32215_;
  assign new_n32217_ = ~new_n32214_ & new_n32216_;
  assign new_n32218_ = ~pi0648 & ~new_n32080_;
  assign new_n32219_ = ~new_n32217_ & new_n32218_;
  assign new_n32220_ = pi0789 & ~new_n32219_;
  assign new_n32221_ = ~new_n32213_ & new_n32220_;
  assign new_n32222_ = ~pi0789 & new_n32207_;
  assign new_n32223_ = new_n17969_ & ~new_n32222_;
  assign new_n32224_ = ~new_n32221_ & new_n32223_;
  assign new_n32225_ = pi0626 & ~new_n32087_;
  assign new_n32226_ = ~pi0626 & ~new_n31966_;
  assign new_n32227_ = new_n17731_ & ~new_n32226_;
  assign new_n32228_ = ~new_n32225_ & new_n32227_;
  assign new_n32229_ = new_n17856_ & new_n32001_;
  assign new_n32230_ = ~pi0626 & ~new_n32087_;
  assign new_n32231_ = pi0626 & ~new_n31966_;
  assign new_n32232_ = new_n17732_ & ~new_n32231_;
  assign new_n32233_ = ~new_n32230_ & new_n32232_;
  assign new_n32234_ = ~new_n32229_ & ~new_n32233_;
  assign new_n32235_ = ~new_n32228_ & new_n32234_;
  assign new_n32236_ = pi0788 & ~new_n32235_;
  assign new_n32237_ = ~new_n20364_ & ~new_n32236_;
  assign new_n32238_ = ~new_n32224_ & new_n32237_;
  assign new_n32239_ = ~new_n32122_ & ~new_n32238_;
  assign new_n32240_ = ~new_n20360_ & ~new_n32239_;
  assign new_n32241_ = new_n17801_ & new_n32023_;
  assign new_n32242_ = new_n17802_ & new_n32019_;
  assign new_n32243_ = ~new_n20556_ & new_n32093_;
  assign new_n32244_ = ~new_n32242_ & ~new_n32243_;
  assign new_n32245_ = ~new_n32241_ & new_n32244_;
  assign new_n32246_ = pi0787 & ~new_n32245_;
  assign new_n32247_ = ~new_n32240_ & ~new_n32246_;
  assign new_n32248_ = ~new_n32116_ & new_n32247_;
  assign new_n32249_ = ~new_n32112_ & ~new_n32248_;
  assign new_n32250_ = ~po1038 & ~new_n32249_;
  assign new_n32251_ = ~pi0192 & po1038;
  assign new_n32252_ = ~pi0832 & ~new_n32251_;
  assign new_n32253_ = ~new_n32250_ & new_n32252_;
  assign po0349 = ~new_n31965_ & ~new_n32253_;
  assign new_n32255_ = ~pi0193 & ~new_n2754_;
  assign new_n32256_ = pi0739 & new_n16913_;
  assign new_n32257_ = ~new_n32255_ & ~new_n32256_;
  assign new_n32258_ = ~new_n17858_ & ~new_n32257_;
  assign new_n32259_ = ~pi0785 & ~new_n32258_;
  assign new_n32260_ = new_n17603_ & new_n32256_;
  assign new_n32261_ = new_n32258_ & ~new_n32260_;
  assign new_n32262_ = pi1155 & ~new_n32261_;
  assign new_n32263_ = ~pi1155 & ~new_n32255_;
  assign new_n32264_ = ~new_n32260_ & new_n32263_;
  assign new_n32265_ = ~new_n32262_ & ~new_n32264_;
  assign new_n32266_ = pi0785 & ~new_n32265_;
  assign new_n32267_ = ~new_n32259_ & ~new_n32266_;
  assign new_n32268_ = ~pi0781 & ~new_n32267_;
  assign new_n32269_ = ~new_n17873_ & new_n32267_;
  assign new_n32270_ = pi1154 & ~new_n32269_;
  assign new_n32271_ = ~new_n17876_ & new_n32267_;
  assign new_n32272_ = ~pi1154 & ~new_n32271_;
  assign new_n32273_ = ~new_n32270_ & ~new_n32272_;
  assign new_n32274_ = pi0781 & ~new_n32273_;
  assign new_n32275_ = ~new_n32268_ & ~new_n32274_;
  assign new_n32276_ = ~pi0789 & ~new_n32275_;
  assign new_n32277_ = ~new_n23057_ & new_n32275_;
  assign new_n32278_ = pi1159 & ~new_n32277_;
  assign new_n32279_ = ~new_n23060_ & new_n32275_;
  assign new_n32280_ = ~pi1159 & ~new_n32279_;
  assign new_n32281_ = ~new_n32278_ & ~new_n32280_;
  assign new_n32282_ = pi0789 & ~new_n32281_;
  assign new_n32283_ = ~new_n32276_ & ~new_n32282_;
  assign new_n32284_ = ~new_n17968_ & new_n32283_;
  assign new_n32285_ = new_n17968_ & new_n32255_;
  assign new_n32286_ = ~new_n32284_ & ~new_n32285_;
  assign new_n32287_ = ~new_n17762_ & ~new_n32286_;
  assign new_n32288_ = new_n17762_ & new_n32255_;
  assign new_n32289_ = ~new_n32287_ & ~new_n32288_;
  assign new_n32290_ = ~new_n20556_ & new_n32289_;
  assign new_n32291_ = pi0690 & new_n16915_;
  assign new_n32292_ = ~new_n32255_ & ~new_n32291_;
  assign new_n32293_ = ~pi0778 & ~new_n32292_;
  assign new_n32294_ = ~pi0625 & new_n32291_;
  assign new_n32295_ = ~new_n32292_ & ~new_n32294_;
  assign new_n32296_ = pi1153 & ~new_n32295_;
  assign new_n32297_ = ~pi1153 & ~new_n32255_;
  assign new_n32298_ = ~new_n32294_ & new_n32297_;
  assign new_n32299_ = pi0778 & ~new_n32298_;
  assign new_n32300_ = ~new_n32296_ & new_n32299_;
  assign new_n32301_ = ~new_n32293_ & ~new_n32300_;
  assign new_n32302_ = ~new_n17844_ & ~new_n32301_;
  assign new_n32303_ = ~new_n17846_ & new_n32302_;
  assign new_n32304_ = ~new_n17848_ & new_n32303_;
  assign new_n32305_ = ~new_n17980_ & new_n32304_;
  assign new_n32306_ = ~new_n18011_ & new_n32305_;
  assign new_n32307_ = ~pi0647 & new_n32306_;
  assign new_n32308_ = pi0647 & new_n32255_;
  assign new_n32309_ = ~pi1157 & ~new_n32308_;
  assign new_n32310_ = ~new_n32307_ & new_n32309_;
  assign new_n32311_ = pi0630 & new_n32310_;
  assign new_n32312_ = pi0647 & ~new_n32306_;
  assign new_n32313_ = ~pi0647 & ~new_n32255_;
  assign new_n32314_ = ~new_n32312_ & ~new_n32313_;
  assign new_n32315_ = new_n17801_ & ~new_n32314_;
  assign new_n32316_ = ~new_n32311_ & ~new_n32315_;
  assign new_n32317_ = ~new_n32290_ & new_n32316_;
  assign new_n32318_ = pi0787 & ~new_n32317_;
  assign new_n32319_ = pi0626 & ~new_n32283_;
  assign new_n32320_ = ~pi0626 & ~new_n32255_;
  assign new_n32321_ = new_n17731_ & ~new_n32320_;
  assign new_n32322_ = ~new_n32319_ & new_n32321_;
  assign new_n32323_ = new_n17856_ & new_n32304_;
  assign new_n32324_ = ~pi0626 & ~new_n32283_;
  assign new_n32325_ = pi0626 & ~new_n32255_;
  assign new_n32326_ = new_n17732_ & ~new_n32325_;
  assign new_n32327_ = ~new_n32324_ & new_n32326_;
  assign new_n32328_ = ~new_n32323_ & ~new_n32327_;
  assign new_n32329_ = ~new_n32322_ & new_n32328_;
  assign new_n32330_ = pi0788 & ~new_n32329_;
  assign new_n32331_ = ~new_n16639_ & ~new_n32292_;
  assign new_n32332_ = pi0625 & new_n32331_;
  assign new_n32333_ = new_n32257_ & ~new_n32331_;
  assign new_n32334_ = ~new_n32332_ & ~new_n32333_;
  assign new_n32335_ = new_n32297_ & ~new_n32334_;
  assign new_n32336_ = ~pi0608 & ~new_n32296_;
  assign new_n32337_ = ~new_n32335_ & new_n32336_;
  assign new_n32338_ = pi1153 & new_n32257_;
  assign new_n32339_ = ~new_n32332_ & new_n32338_;
  assign new_n32340_ = pi0608 & ~new_n32298_;
  assign new_n32341_ = ~new_n32339_ & new_n32340_;
  assign new_n32342_ = ~new_n32337_ & ~new_n32341_;
  assign new_n32343_ = pi0778 & ~new_n32342_;
  assign new_n32344_ = ~pi0778 & ~new_n32333_;
  assign new_n32345_ = ~new_n32343_ & ~new_n32344_;
  assign new_n32346_ = ~pi0609 & ~new_n32345_;
  assign new_n32347_ = pi0609 & ~new_n32301_;
  assign new_n32348_ = ~pi1155 & ~new_n32347_;
  assign new_n32349_ = ~new_n32346_ & new_n32348_;
  assign new_n32350_ = ~pi0660 & ~new_n32262_;
  assign new_n32351_ = ~new_n32349_ & new_n32350_;
  assign new_n32352_ = pi0609 & ~new_n32345_;
  assign new_n32353_ = ~pi0609 & ~new_n32301_;
  assign new_n32354_ = pi1155 & ~new_n32353_;
  assign new_n32355_ = ~new_n32352_ & new_n32354_;
  assign new_n32356_ = pi0660 & ~new_n32264_;
  assign new_n32357_ = ~new_n32355_ & new_n32356_;
  assign new_n32358_ = ~new_n32351_ & ~new_n32357_;
  assign new_n32359_ = pi0785 & ~new_n32358_;
  assign new_n32360_ = ~pi0785 & ~new_n32345_;
  assign new_n32361_ = ~new_n32359_ & ~new_n32360_;
  assign new_n32362_ = ~pi0618 & ~new_n32361_;
  assign new_n32363_ = pi0618 & new_n32302_;
  assign new_n32364_ = ~pi1154 & ~new_n32363_;
  assign new_n32365_ = ~new_n32362_ & new_n32364_;
  assign new_n32366_ = ~pi0627 & ~new_n32270_;
  assign new_n32367_ = ~new_n32365_ & new_n32366_;
  assign new_n32368_ = pi0618 & ~new_n32361_;
  assign new_n32369_ = ~pi0618 & new_n32302_;
  assign new_n32370_ = pi1154 & ~new_n32369_;
  assign new_n32371_ = ~new_n32368_ & new_n32370_;
  assign new_n32372_ = pi0627 & ~new_n32272_;
  assign new_n32373_ = ~new_n32371_ & new_n32372_;
  assign new_n32374_ = ~new_n32367_ & ~new_n32373_;
  assign new_n32375_ = pi0781 & ~new_n32374_;
  assign new_n32376_ = ~pi0781 & ~new_n32361_;
  assign new_n32377_ = ~new_n32375_ & ~new_n32376_;
  assign new_n32378_ = pi0619 & ~new_n32377_;
  assign new_n32379_ = ~pi0619 & new_n32303_;
  assign new_n32380_ = pi1159 & ~new_n32379_;
  assign new_n32381_ = ~new_n32378_ & new_n32380_;
  assign new_n32382_ = pi0648 & ~new_n32280_;
  assign new_n32383_ = ~new_n32381_ & new_n32382_;
  assign new_n32384_ = ~pi0619 & ~new_n32377_;
  assign new_n32385_ = pi0619 & new_n32303_;
  assign new_n32386_ = ~pi1159 & ~new_n32385_;
  assign new_n32387_ = ~new_n32384_ & new_n32386_;
  assign new_n32388_ = ~pi0648 & ~new_n32278_;
  assign new_n32389_ = ~new_n32387_ & new_n32388_;
  assign new_n32390_ = pi0789 & ~new_n32389_;
  assign new_n32391_ = ~new_n32383_ & new_n32390_;
  assign new_n32392_ = ~pi0789 & new_n32377_;
  assign new_n32393_ = new_n17969_ & ~new_n32392_;
  assign new_n32394_ = ~new_n32391_ & new_n32393_;
  assign new_n32395_ = ~new_n32330_ & ~new_n32394_;
  assign new_n32396_ = ~new_n20364_ & ~new_n32395_;
  assign new_n32397_ = new_n18008_ & ~new_n32286_;
  assign new_n32398_ = new_n20851_ & new_n32305_;
  assign new_n32399_ = ~new_n32397_ & ~new_n32398_;
  assign new_n32400_ = ~pi0629 & ~new_n32399_;
  assign new_n32401_ = new_n20855_ & new_n32305_;
  assign new_n32402_ = new_n18007_ & ~new_n32286_;
  assign new_n32403_ = ~new_n32401_ & ~new_n32402_;
  assign new_n32404_ = pi0629 & ~new_n32403_;
  assign new_n32405_ = ~new_n32400_ & ~new_n32404_;
  assign new_n32406_ = pi0792 & ~new_n32405_;
  assign new_n32407_ = ~new_n20360_ & ~new_n32406_;
  assign new_n32408_ = ~new_n32396_ & new_n32407_;
  assign new_n32409_ = ~new_n32318_ & ~new_n32408_;
  assign new_n32410_ = pi0644 & new_n32409_;
  assign new_n32411_ = ~pi0787 & ~new_n32306_;
  assign new_n32412_ = pi1157 & ~new_n32314_;
  assign new_n32413_ = ~new_n32310_ & ~new_n32412_;
  assign new_n32414_ = pi0787 & ~new_n32413_;
  assign new_n32415_ = ~new_n32411_ & ~new_n32414_;
  assign new_n32416_ = ~pi0644 & new_n32415_;
  assign new_n32417_ = pi0715 & ~new_n32416_;
  assign new_n32418_ = ~new_n32410_ & new_n32417_;
  assign new_n32419_ = ~new_n17804_ & ~new_n32289_;
  assign new_n32420_ = new_n17804_ & new_n32255_;
  assign new_n32421_ = ~new_n32419_ & ~new_n32420_;
  assign new_n32422_ = pi0644 & ~new_n32421_;
  assign new_n32423_ = ~pi0644 & new_n32255_;
  assign new_n32424_ = ~pi0715 & ~new_n32423_;
  assign new_n32425_ = ~new_n32422_ & new_n32424_;
  assign new_n32426_ = pi1160 & ~new_n32425_;
  assign new_n32427_ = ~new_n32418_ & new_n32426_;
  assign new_n32428_ = ~pi0644 & new_n32409_;
  assign new_n32429_ = pi0644 & new_n32415_;
  assign new_n32430_ = ~pi0715 & ~new_n32429_;
  assign new_n32431_ = ~new_n32428_ & new_n32430_;
  assign new_n32432_ = ~pi0644 & ~new_n32421_;
  assign new_n32433_ = pi0644 & new_n32255_;
  assign new_n32434_ = pi0715 & ~new_n32433_;
  assign new_n32435_ = ~new_n32432_ & new_n32434_;
  assign new_n32436_ = ~pi1160 & ~new_n32435_;
  assign new_n32437_ = ~new_n32431_ & new_n32436_;
  assign new_n32438_ = ~new_n32427_ & ~new_n32437_;
  assign new_n32439_ = pi0790 & ~new_n32438_;
  assign new_n32440_ = ~pi0790 & new_n32409_;
  assign new_n32441_ = pi0832 & ~new_n32440_;
  assign new_n32442_ = ~new_n32439_ & new_n32441_;
  assign new_n32443_ = ~pi0193 & ~new_n17558_;
  assign new_n32444_ = new_n17691_ & ~new_n32443_;
  assign new_n32445_ = pi0690 & new_n3272_;
  assign new_n32446_ = new_n32443_ & ~new_n32445_;
  assign new_n32447_ = pi0193 & ~new_n18128_;
  assign new_n32448_ = ~pi0038 & ~new_n32447_;
  assign new_n32449_ = new_n3272_ & ~new_n32448_;
  assign new_n32450_ = ~pi0193 & new_n18124_;
  assign new_n32451_ = ~new_n32449_ & ~new_n32450_;
  assign new_n32452_ = ~pi0193 & ~new_n17431_;
  assign new_n32453_ = new_n17544_ & ~new_n32452_;
  assign new_n32454_ = pi0690 & ~new_n32453_;
  assign new_n32455_ = ~new_n32451_ & new_n32454_;
  assign new_n32456_ = ~new_n32446_ & ~new_n32455_;
  assign new_n32457_ = ~pi0778 & new_n32456_;
  assign new_n32458_ = pi0625 & ~new_n32456_;
  assign new_n32459_ = ~pi0625 & new_n32443_;
  assign new_n32460_ = pi1153 & ~new_n32459_;
  assign new_n32461_ = ~new_n32458_ & new_n32460_;
  assign new_n32462_ = ~pi0625 & ~new_n32456_;
  assign new_n32463_ = pi0625 & new_n32443_;
  assign new_n32464_ = ~pi1153 & ~new_n32463_;
  assign new_n32465_ = ~new_n32462_ & new_n32464_;
  assign new_n32466_ = ~new_n32461_ & ~new_n32465_;
  assign new_n32467_ = pi0778 & ~new_n32466_;
  assign new_n32468_ = ~new_n32457_ & ~new_n32467_;
  assign new_n32469_ = ~new_n17618_ & ~new_n32468_;
  assign new_n32470_ = new_n17618_ & ~new_n32443_;
  assign new_n32471_ = ~new_n32469_ & ~new_n32470_;
  assign new_n32472_ = ~new_n17655_ & new_n32471_;
  assign new_n32473_ = new_n17655_ & new_n32443_;
  assign new_n32474_ = ~new_n32472_ & ~new_n32473_;
  assign new_n32475_ = ~new_n17691_ & new_n32474_;
  assign new_n32476_ = ~new_n32444_ & ~new_n32475_;
  assign new_n32477_ = ~new_n17734_ & new_n32476_;
  assign new_n32478_ = new_n17734_ & new_n32443_;
  assign new_n32479_ = ~new_n32477_ & ~new_n32478_;
  assign new_n32480_ = ~pi0792 & new_n32479_;
  assign new_n32481_ = pi0628 & ~new_n32479_;
  assign new_n32482_ = ~pi0628 & new_n32443_;
  assign new_n32483_ = pi1156 & ~new_n32482_;
  assign new_n32484_ = ~new_n32481_ & new_n32483_;
  assign new_n32485_ = ~pi0628 & ~new_n32479_;
  assign new_n32486_ = pi0628 & new_n32443_;
  assign new_n32487_ = ~pi1156 & ~new_n32486_;
  assign new_n32488_ = ~new_n32485_ & new_n32487_;
  assign new_n32489_ = ~new_n32484_ & ~new_n32488_;
  assign new_n32490_ = pi0792 & ~new_n32489_;
  assign new_n32491_ = ~new_n32480_ & ~new_n32490_;
  assign new_n32492_ = ~pi0647 & ~new_n32491_;
  assign new_n32493_ = pi0647 & ~new_n32443_;
  assign new_n32494_ = ~new_n32492_ & ~new_n32493_;
  assign new_n32495_ = ~pi1157 & new_n32494_;
  assign new_n32496_ = pi0647 & ~new_n32491_;
  assign new_n32497_ = ~pi0647 & ~new_n32443_;
  assign new_n32498_ = ~new_n32496_ & ~new_n32497_;
  assign new_n32499_ = pi1157 & new_n32498_;
  assign new_n32500_ = ~new_n32495_ & ~new_n32499_;
  assign new_n32501_ = pi0787 & ~new_n32500_;
  assign new_n32502_ = ~pi0787 & new_n32491_;
  assign new_n32503_ = ~new_n32501_ & ~new_n32502_;
  assign new_n32504_ = ~pi0644 & ~new_n32503_;
  assign new_n32505_ = pi0715 & ~new_n32504_;
  assign new_n32506_ = pi0193 & ~new_n3272_;
  assign new_n32507_ = pi0739 & new_n17433_;
  assign new_n32508_ = ~new_n32452_ & ~new_n32507_;
  assign new_n32509_ = pi0038 & ~new_n32508_;
  assign new_n32510_ = ~pi0193 & new_n17393_;
  assign new_n32511_ = pi0193 & ~new_n17426_;
  assign new_n32512_ = pi0739 & ~new_n32511_;
  assign new_n32513_ = ~new_n32510_ & new_n32512_;
  assign new_n32514_ = ~pi0193 & ~pi0739;
  assign new_n32515_ = ~new_n17349_ & new_n32514_;
  assign new_n32516_ = ~new_n32513_ & ~new_n32515_;
  assign new_n32517_ = ~pi0038 & ~new_n32516_;
  assign new_n32518_ = ~new_n32509_ & ~new_n32517_;
  assign new_n32519_ = new_n3272_ & new_n32518_;
  assign new_n32520_ = ~new_n32506_ & ~new_n32519_;
  assign new_n32521_ = ~new_n17590_ & ~new_n32520_;
  assign new_n32522_ = new_n17590_ & ~new_n32443_;
  assign new_n32523_ = ~new_n32521_ & ~new_n32522_;
  assign new_n32524_ = ~pi0785 & ~new_n32523_;
  assign new_n32525_ = ~new_n17591_ & ~new_n32443_;
  assign new_n32526_ = pi0609 & new_n32521_;
  assign new_n32527_ = ~new_n32525_ & ~new_n32526_;
  assign new_n32528_ = pi1155 & ~new_n32527_;
  assign new_n32529_ = ~new_n17603_ & ~new_n32443_;
  assign new_n32530_ = ~pi0609 & new_n32521_;
  assign new_n32531_ = ~new_n32529_ & ~new_n32530_;
  assign new_n32532_ = ~pi1155 & ~new_n32531_;
  assign new_n32533_ = ~new_n32528_ & ~new_n32532_;
  assign new_n32534_ = pi0785 & ~new_n32533_;
  assign new_n32535_ = ~new_n32524_ & ~new_n32534_;
  assign new_n32536_ = ~pi0781 & ~new_n32535_;
  assign new_n32537_ = pi0618 & new_n32535_;
  assign new_n32538_ = ~pi0618 & new_n32443_;
  assign new_n32539_ = pi1154 & ~new_n32538_;
  assign new_n32540_ = ~new_n32537_ & new_n32539_;
  assign new_n32541_ = ~pi0618 & new_n32535_;
  assign new_n32542_ = pi0618 & new_n32443_;
  assign new_n32543_ = ~pi1154 & ~new_n32542_;
  assign new_n32544_ = ~new_n32541_ & new_n32543_;
  assign new_n32545_ = ~new_n32540_ & ~new_n32544_;
  assign new_n32546_ = pi0781 & ~new_n32545_;
  assign new_n32547_ = ~new_n32536_ & ~new_n32546_;
  assign new_n32548_ = ~pi0789 & ~new_n32547_;
  assign new_n32549_ = pi0619 & new_n32547_;
  assign new_n32550_ = ~pi0619 & new_n32443_;
  assign new_n32551_ = pi1159 & ~new_n32550_;
  assign new_n32552_ = ~new_n32549_ & new_n32551_;
  assign new_n32553_ = ~pi0619 & new_n32547_;
  assign new_n32554_ = pi0619 & new_n32443_;
  assign new_n32555_ = ~pi1159 & ~new_n32554_;
  assign new_n32556_ = ~new_n32553_ & new_n32555_;
  assign new_n32557_ = ~new_n32552_ & ~new_n32556_;
  assign new_n32558_ = pi0789 & ~new_n32557_;
  assign new_n32559_ = ~new_n32548_ & ~new_n32558_;
  assign new_n32560_ = ~new_n17968_ & new_n32559_;
  assign new_n32561_ = new_n17968_ & new_n32443_;
  assign new_n32562_ = ~new_n32560_ & ~new_n32561_;
  assign new_n32563_ = ~new_n17762_ & ~new_n32562_;
  assign new_n32564_ = new_n17762_ & new_n32443_;
  assign new_n32565_ = ~new_n32563_ & ~new_n32564_;
  assign new_n32566_ = ~new_n17804_ & ~new_n32565_;
  assign new_n32567_ = new_n17804_ & new_n32443_;
  assign new_n32568_ = ~new_n32566_ & ~new_n32567_;
  assign new_n32569_ = pi0644 & ~new_n32568_;
  assign new_n32570_ = ~pi0644 & new_n32443_;
  assign new_n32571_ = ~pi0715 & ~new_n32570_;
  assign new_n32572_ = ~new_n32569_ & new_n32571_;
  assign new_n32573_ = pi1160 & ~new_n32572_;
  assign new_n32574_ = ~new_n32505_ & new_n32573_;
  assign new_n32575_ = pi0644 & ~new_n32503_;
  assign new_n32576_ = ~pi0715 & ~new_n32575_;
  assign new_n32577_ = ~pi0644 & ~new_n32568_;
  assign new_n32578_ = pi0644 & new_n32443_;
  assign new_n32579_ = pi0715 & ~new_n32578_;
  assign new_n32580_ = ~new_n32577_ & new_n32579_;
  assign new_n32581_ = ~pi1160 & ~new_n32580_;
  assign new_n32582_ = ~new_n32576_ & new_n32581_;
  assign new_n32583_ = ~new_n32574_ & ~new_n32582_;
  assign new_n32584_ = pi0790 & ~new_n32583_;
  assign new_n32585_ = pi0644 & new_n32573_;
  assign new_n32586_ = ~pi0644 & new_n32581_;
  assign new_n32587_ = pi0790 & ~new_n32586_;
  assign new_n32588_ = ~new_n32585_ & new_n32587_;
  assign new_n32589_ = ~new_n20567_ & new_n32562_;
  assign new_n32590_ = ~pi0629 & new_n32484_;
  assign new_n32591_ = pi0629 & new_n32488_;
  assign new_n32592_ = ~new_n32590_ & ~new_n32591_;
  assign new_n32593_ = ~new_n32589_ & new_n32592_;
  assign new_n32594_ = pi0792 & ~new_n32593_;
  assign new_n32595_ = ~pi0690 & ~new_n32518_;
  assign new_n32596_ = ~pi0193 & new_n16810_;
  assign new_n32597_ = pi0193 & new_n16928_;
  assign new_n32598_ = ~pi0739 & ~new_n32597_;
  assign new_n32599_ = ~new_n32596_ & new_n32598_;
  assign new_n32600_ = pi0193 & new_n17007_;
  assign new_n32601_ = ~pi0193 & ~new_n17074_;
  assign new_n32602_ = pi0739 & ~new_n32601_;
  assign new_n32603_ = ~new_n32600_ & new_n32602_;
  assign new_n32604_ = pi0039 & ~new_n32603_;
  assign new_n32605_ = ~new_n32599_ & new_n32604_;
  assign new_n32606_ = ~pi0193 & new_n17227_;
  assign new_n32607_ = pi0193 & new_n17234_;
  assign new_n32608_ = pi0739 & ~new_n32607_;
  assign new_n32609_ = ~new_n32606_ & new_n32608_;
  assign new_n32610_ = ~pi0193 & ~new_n17217_;
  assign new_n32611_ = pi0193 & ~new_n17178_;
  assign new_n32612_ = ~pi0739 & ~new_n32611_;
  assign new_n32613_ = ~new_n32610_ & new_n32612_;
  assign new_n32614_ = ~new_n32609_ & ~new_n32613_;
  assign new_n32615_ = ~pi0039 & ~new_n32614_;
  assign new_n32616_ = ~pi0038 & ~new_n32615_;
  assign new_n32617_ = ~new_n32605_ & new_n32616_;
  assign new_n32618_ = ~pi0739 & new_n24079_;
  assign new_n32619_ = ~new_n17035_ & ~new_n32618_;
  assign new_n32620_ = ~pi0039 & ~new_n32619_;
  assign new_n32621_ = ~pi0193 & ~new_n32620_;
  assign new_n32622_ = ~new_n16916_ & ~new_n32256_;
  assign new_n32623_ = pi0193 & ~new_n32622_;
  assign new_n32624_ = new_n6257_ & new_n32623_;
  assign new_n32625_ = pi0038 & ~new_n32624_;
  assign new_n32626_ = ~new_n32621_ & new_n32625_;
  assign new_n32627_ = pi0690 & ~new_n32626_;
  assign new_n32628_ = ~new_n32617_ & new_n32627_;
  assign new_n32629_ = new_n3272_ & ~new_n32628_;
  assign new_n32630_ = ~new_n32595_ & new_n32629_;
  assign new_n32631_ = ~new_n32506_ & ~new_n32630_;
  assign new_n32632_ = ~pi0625 & new_n32631_;
  assign new_n32633_ = pi0625 & new_n32520_;
  assign new_n32634_ = ~pi1153 & ~new_n32633_;
  assign new_n32635_ = ~new_n32632_ & new_n32634_;
  assign new_n32636_ = ~pi0608 & ~new_n32461_;
  assign new_n32637_ = ~new_n32635_ & new_n32636_;
  assign new_n32638_ = pi0625 & new_n32631_;
  assign new_n32639_ = ~pi0625 & new_n32520_;
  assign new_n32640_ = pi1153 & ~new_n32639_;
  assign new_n32641_ = ~new_n32638_ & new_n32640_;
  assign new_n32642_ = pi0608 & ~new_n32465_;
  assign new_n32643_ = ~new_n32641_ & new_n32642_;
  assign new_n32644_ = ~new_n32637_ & ~new_n32643_;
  assign new_n32645_ = pi0778 & ~new_n32644_;
  assign new_n32646_ = ~pi0778 & new_n32631_;
  assign new_n32647_ = ~new_n32645_ & ~new_n32646_;
  assign new_n32648_ = ~pi0609 & ~new_n32647_;
  assign new_n32649_ = pi0609 & new_n32468_;
  assign new_n32650_ = ~pi1155 & ~new_n32649_;
  assign new_n32651_ = ~new_n32648_ & new_n32650_;
  assign new_n32652_ = ~pi0660 & ~new_n32528_;
  assign new_n32653_ = ~new_n32651_ & new_n32652_;
  assign new_n32654_ = pi0609 & ~new_n32647_;
  assign new_n32655_ = ~pi0609 & new_n32468_;
  assign new_n32656_ = pi1155 & ~new_n32655_;
  assign new_n32657_ = ~new_n32654_ & new_n32656_;
  assign new_n32658_ = pi0660 & ~new_n32532_;
  assign new_n32659_ = ~new_n32657_ & new_n32658_;
  assign new_n32660_ = ~new_n32653_ & ~new_n32659_;
  assign new_n32661_ = pi0785 & ~new_n32660_;
  assign new_n32662_ = ~pi0785 & ~new_n32647_;
  assign new_n32663_ = ~new_n32661_ & ~new_n32662_;
  assign new_n32664_ = ~pi0618 & ~new_n32663_;
  assign new_n32665_ = pi0618 & new_n32471_;
  assign new_n32666_ = ~pi1154 & ~new_n32665_;
  assign new_n32667_ = ~new_n32664_ & new_n32666_;
  assign new_n32668_ = ~pi0627 & ~new_n32540_;
  assign new_n32669_ = ~new_n32667_ & new_n32668_;
  assign new_n32670_ = pi0618 & ~new_n32663_;
  assign new_n32671_ = ~pi0618 & new_n32471_;
  assign new_n32672_ = pi1154 & ~new_n32671_;
  assign new_n32673_ = ~new_n32670_ & new_n32672_;
  assign new_n32674_ = pi0627 & ~new_n32544_;
  assign new_n32675_ = ~new_n32673_ & new_n32674_;
  assign new_n32676_ = ~new_n32669_ & ~new_n32675_;
  assign new_n32677_ = pi0781 & ~new_n32676_;
  assign new_n32678_ = ~pi0781 & ~new_n32663_;
  assign new_n32679_ = ~new_n32677_ & ~new_n32678_;
  assign new_n32680_ = pi0619 & ~new_n32679_;
  assign new_n32681_ = ~pi0619 & ~new_n32474_;
  assign new_n32682_ = pi1159 & ~new_n32681_;
  assign new_n32683_ = ~new_n32680_ & new_n32682_;
  assign new_n32684_ = pi0648 & ~new_n32556_;
  assign new_n32685_ = ~new_n32683_ & new_n32684_;
  assign new_n32686_ = ~pi0619 & ~new_n32679_;
  assign new_n32687_ = pi0619 & ~new_n32474_;
  assign new_n32688_ = ~pi1159 & ~new_n32687_;
  assign new_n32689_ = ~new_n32686_ & new_n32688_;
  assign new_n32690_ = ~pi0648 & ~new_n32552_;
  assign new_n32691_ = ~new_n32689_ & new_n32690_;
  assign new_n32692_ = pi0789 & ~new_n32691_;
  assign new_n32693_ = ~new_n32685_ & new_n32692_;
  assign new_n32694_ = ~pi0789 & new_n32679_;
  assign new_n32695_ = new_n17969_ & ~new_n32694_;
  assign new_n32696_ = ~new_n32693_ & new_n32695_;
  assign new_n32697_ = pi0626 & ~new_n32559_;
  assign new_n32698_ = ~pi0626 & ~new_n32443_;
  assign new_n32699_ = new_n17731_ & ~new_n32698_;
  assign new_n32700_ = ~new_n32697_ & new_n32699_;
  assign new_n32701_ = new_n17856_ & new_n32476_;
  assign new_n32702_ = ~pi0626 & ~new_n32559_;
  assign new_n32703_ = pi0626 & ~new_n32443_;
  assign new_n32704_ = new_n17732_ & ~new_n32703_;
  assign new_n32705_ = ~new_n32702_ & new_n32704_;
  assign new_n32706_ = ~new_n32701_ & ~new_n32705_;
  assign new_n32707_ = ~new_n32700_ & new_n32706_;
  assign new_n32708_ = pi0788 & ~new_n32707_;
  assign new_n32709_ = ~new_n20364_ & ~new_n32708_;
  assign new_n32710_ = ~new_n32696_ & new_n32709_;
  assign new_n32711_ = ~new_n32594_ & ~new_n32710_;
  assign new_n32712_ = ~new_n20360_ & ~new_n32711_;
  assign new_n32713_ = ~new_n20556_ & new_n32565_;
  assign new_n32714_ = new_n17802_ & ~new_n32494_;
  assign new_n32715_ = new_n17801_ & ~new_n32498_;
  assign new_n32716_ = ~new_n32714_ & ~new_n32715_;
  assign new_n32717_ = ~new_n32713_ & new_n32716_;
  assign new_n32718_ = pi0787 & ~new_n32717_;
  assign new_n32719_ = ~new_n32712_ & ~new_n32718_;
  assign new_n32720_ = ~new_n32588_ & new_n32719_;
  assign new_n32721_ = ~new_n32584_ & ~new_n32720_;
  assign new_n32722_ = ~po1038 & ~new_n32721_;
  assign new_n32723_ = ~pi0193 & po1038;
  assign new_n32724_ = ~pi0832 & ~new_n32723_;
  assign new_n32725_ = ~new_n32722_ & new_n32724_;
  assign po0350 = ~new_n32442_ & ~new_n32725_;
  assign new_n32727_ = pi0194 & ~new_n3272_;
  assign new_n32728_ = ~pi0194 & new_n19389_;
  assign new_n32729_ = pi0194 & ~new_n24548_;
  assign new_n32730_ = ~pi0748 & ~new_n32729_;
  assign new_n32731_ = ~new_n32728_ & new_n32730_;
  assign new_n32732_ = pi0194 & new_n19406_;
  assign new_n32733_ = ~pi0194 & ~new_n19414_;
  assign new_n32734_ = pi0748 & ~new_n32733_;
  assign new_n32735_ = ~new_n32732_ & new_n32734_;
  assign new_n32736_ = pi0730 & ~new_n32735_;
  assign new_n32737_ = ~new_n32731_ & new_n32736_;
  assign new_n32738_ = ~pi0194 & new_n19376_;
  assign new_n32739_ = pi0194 & new_n24446_;
  assign new_n32740_ = ~new_n32738_ & ~new_n32739_;
  assign new_n32741_ = pi0748 & ~new_n32740_;
  assign new_n32742_ = ~pi0194 & ~new_n17551_;
  assign new_n32743_ = ~pi0748 & ~new_n32742_;
  assign new_n32744_ = ~new_n32741_ & ~new_n32743_;
  assign new_n32745_ = ~pi0730 & new_n32744_;
  assign new_n32746_ = new_n3272_ & ~new_n32745_;
  assign new_n32747_ = ~new_n32737_ & new_n32746_;
  assign new_n32748_ = ~new_n32727_ & ~new_n32747_;
  assign new_n32749_ = ~pi0625 & new_n32748_;
  assign new_n32750_ = new_n3272_ & ~new_n32744_;
  assign new_n32751_ = ~new_n32727_ & ~new_n32750_;
  assign new_n32752_ = pi0625 & new_n32751_;
  assign new_n32753_ = ~pi1153 & ~new_n32752_;
  assign new_n32754_ = ~new_n32749_ & new_n32753_;
  assign new_n32755_ = pi0194 & ~new_n24384_;
  assign new_n32756_ = ~pi0194 & new_n24387_;
  assign new_n32757_ = pi0730 & ~new_n32756_;
  assign new_n32758_ = ~pi0730 & new_n32742_;
  assign new_n32759_ = new_n3272_ & ~new_n32758_;
  assign new_n32760_ = ~new_n32757_ & new_n32759_;
  assign new_n32761_ = ~new_n32755_ & ~new_n32760_;
  assign new_n32762_ = pi0625 & new_n32761_;
  assign new_n32763_ = ~pi0194 & ~new_n17558_;
  assign new_n32764_ = ~pi0625 & new_n32763_;
  assign new_n32765_ = pi1153 & ~new_n32764_;
  assign new_n32766_ = ~new_n32762_ & new_n32765_;
  assign new_n32767_ = ~pi0608 & ~new_n32766_;
  assign new_n32768_ = ~new_n32754_ & new_n32767_;
  assign new_n32769_ = pi0625 & new_n32748_;
  assign new_n32770_ = ~pi0625 & new_n32751_;
  assign new_n32771_ = pi1153 & ~new_n32770_;
  assign new_n32772_ = ~new_n32769_ & new_n32771_;
  assign new_n32773_ = ~pi0625 & new_n32761_;
  assign new_n32774_ = pi0625 & new_n32763_;
  assign new_n32775_ = ~pi1153 & ~new_n32774_;
  assign new_n32776_ = ~new_n32773_ & new_n32775_;
  assign new_n32777_ = pi0608 & ~new_n32776_;
  assign new_n32778_ = ~new_n32772_ & new_n32777_;
  assign new_n32779_ = ~new_n32768_ & ~new_n32778_;
  assign new_n32780_ = pi0778 & ~new_n32779_;
  assign new_n32781_ = ~pi0778 & new_n32748_;
  assign new_n32782_ = ~new_n32780_ & ~new_n32781_;
  assign new_n32783_ = ~pi0609 & ~new_n32782_;
  assign new_n32784_ = ~pi0778 & ~new_n32761_;
  assign new_n32785_ = ~new_n32766_ & ~new_n32776_;
  assign new_n32786_ = pi0778 & ~new_n32785_;
  assign new_n32787_ = ~new_n32784_ & ~new_n32786_;
  assign new_n32788_ = pi0609 & new_n32787_;
  assign new_n32789_ = ~pi1155 & ~new_n32788_;
  assign new_n32790_ = ~new_n32783_ & new_n32789_;
  assign new_n32791_ = ~new_n17591_ & ~new_n32763_;
  assign new_n32792_ = ~new_n17590_ & ~new_n32751_;
  assign new_n32793_ = pi0609 & new_n32792_;
  assign new_n32794_ = ~new_n32791_ & ~new_n32793_;
  assign new_n32795_ = pi1155 & ~new_n32794_;
  assign new_n32796_ = ~pi0660 & ~new_n32795_;
  assign new_n32797_ = ~new_n32790_ & new_n32796_;
  assign new_n32798_ = pi0609 & ~new_n32782_;
  assign new_n32799_ = ~pi0609 & new_n32787_;
  assign new_n32800_ = pi1155 & ~new_n32799_;
  assign new_n32801_ = ~new_n32798_ & new_n32800_;
  assign new_n32802_ = ~new_n17603_ & ~new_n32763_;
  assign new_n32803_ = ~pi0609 & new_n32792_;
  assign new_n32804_ = ~new_n32802_ & ~new_n32803_;
  assign new_n32805_ = ~pi1155 & ~new_n32804_;
  assign new_n32806_ = pi0660 & ~new_n32805_;
  assign new_n32807_ = ~new_n32801_ & new_n32806_;
  assign new_n32808_ = ~new_n32797_ & ~new_n32807_;
  assign new_n32809_ = pi0785 & ~new_n32808_;
  assign new_n32810_ = ~pi0785 & ~new_n32782_;
  assign new_n32811_ = ~new_n32809_ & ~new_n32810_;
  assign new_n32812_ = ~pi0618 & ~new_n32811_;
  assign new_n32813_ = ~new_n17618_ & ~new_n32787_;
  assign new_n32814_ = new_n17618_ & ~new_n32763_;
  assign new_n32815_ = ~new_n32813_ & ~new_n32814_;
  assign new_n32816_ = pi0618 & new_n32815_;
  assign new_n32817_ = ~pi1154 & ~new_n32816_;
  assign new_n32818_ = ~new_n32812_ & new_n32817_;
  assign new_n32819_ = new_n17590_ & ~new_n32763_;
  assign new_n32820_ = ~new_n32792_ & ~new_n32819_;
  assign new_n32821_ = ~pi0785 & ~new_n32820_;
  assign new_n32822_ = ~new_n32795_ & ~new_n32805_;
  assign new_n32823_ = pi0785 & ~new_n32822_;
  assign new_n32824_ = ~new_n32821_ & ~new_n32823_;
  assign new_n32825_ = pi0618 & new_n32824_;
  assign new_n32826_ = ~pi0618 & new_n32763_;
  assign new_n32827_ = pi1154 & ~new_n32826_;
  assign new_n32828_ = ~new_n32825_ & new_n32827_;
  assign new_n32829_ = ~pi0627 & ~new_n32828_;
  assign new_n32830_ = ~new_n32818_ & new_n32829_;
  assign new_n32831_ = pi0618 & ~new_n32811_;
  assign new_n32832_ = ~pi0618 & new_n32815_;
  assign new_n32833_ = pi1154 & ~new_n32832_;
  assign new_n32834_ = ~new_n32831_ & new_n32833_;
  assign new_n32835_ = ~pi0618 & new_n32824_;
  assign new_n32836_ = pi0618 & new_n32763_;
  assign new_n32837_ = ~pi1154 & ~new_n32836_;
  assign new_n32838_ = ~new_n32835_ & new_n32837_;
  assign new_n32839_ = pi0627 & ~new_n32838_;
  assign new_n32840_ = ~new_n32834_ & new_n32839_;
  assign new_n32841_ = ~new_n32830_ & ~new_n32840_;
  assign new_n32842_ = pi0781 & ~new_n32841_;
  assign new_n32843_ = ~pi0781 & ~new_n32811_;
  assign new_n32844_ = ~new_n32842_ & ~new_n32843_;
  assign new_n32845_ = ~pi0619 & ~new_n32844_;
  assign new_n32846_ = ~new_n17655_ & new_n32815_;
  assign new_n32847_ = new_n17655_ & new_n32763_;
  assign new_n32848_ = ~new_n32846_ & ~new_n32847_;
  assign new_n32849_ = pi0619 & ~new_n32848_;
  assign new_n32850_ = ~pi1159 & ~new_n32849_;
  assign new_n32851_ = ~new_n32845_ & new_n32850_;
  assign new_n32852_ = ~pi0781 & ~new_n32824_;
  assign new_n32853_ = ~new_n32828_ & ~new_n32838_;
  assign new_n32854_ = pi0781 & ~new_n32853_;
  assign new_n32855_ = ~new_n32852_ & ~new_n32854_;
  assign new_n32856_ = pi0619 & new_n32855_;
  assign new_n32857_ = ~pi0619 & new_n32763_;
  assign new_n32858_ = pi1159 & ~new_n32857_;
  assign new_n32859_ = ~new_n32856_ & new_n32858_;
  assign new_n32860_ = ~pi0648 & ~new_n32859_;
  assign new_n32861_ = ~new_n32851_ & new_n32860_;
  assign new_n32862_ = pi0619 & ~new_n32844_;
  assign new_n32863_ = ~pi0619 & ~new_n32848_;
  assign new_n32864_ = pi1159 & ~new_n32863_;
  assign new_n32865_ = ~new_n32862_ & new_n32864_;
  assign new_n32866_ = ~pi0619 & new_n32855_;
  assign new_n32867_ = pi0619 & new_n32763_;
  assign new_n32868_ = ~pi1159 & ~new_n32867_;
  assign new_n32869_ = ~new_n32866_ & new_n32868_;
  assign new_n32870_ = pi0648 & ~new_n32869_;
  assign new_n32871_ = ~new_n32865_ & new_n32870_;
  assign new_n32872_ = ~new_n32861_ & ~new_n32871_;
  assign new_n32873_ = pi0789 & ~new_n32872_;
  assign new_n32874_ = ~pi0789 & ~new_n32844_;
  assign new_n32875_ = ~new_n32873_ & ~new_n32874_;
  assign new_n32876_ = ~pi0788 & new_n32875_;
  assign new_n32877_ = ~pi0626 & new_n32875_;
  assign new_n32878_ = new_n17691_ & ~new_n32763_;
  assign new_n32879_ = ~new_n17691_ & new_n32848_;
  assign new_n32880_ = ~new_n32878_ & ~new_n32879_;
  assign new_n32881_ = pi0626 & ~new_n32880_;
  assign new_n32882_ = ~pi0641 & ~new_n32881_;
  assign new_n32883_ = ~new_n32877_ & new_n32882_;
  assign new_n32884_ = ~pi0789 & ~new_n32855_;
  assign new_n32885_ = ~new_n32859_ & ~new_n32869_;
  assign new_n32886_ = pi0789 & ~new_n32885_;
  assign new_n32887_ = ~new_n32884_ & ~new_n32886_;
  assign new_n32888_ = ~pi0626 & ~new_n32887_;
  assign new_n32889_ = pi0626 & ~new_n32763_;
  assign new_n32890_ = pi0641 & ~new_n32889_;
  assign new_n32891_ = ~new_n32888_ & new_n32890_;
  assign new_n32892_ = ~pi1158 & ~new_n32891_;
  assign new_n32893_ = ~new_n32883_ & new_n32892_;
  assign new_n32894_ = pi0626 & new_n32875_;
  assign new_n32895_ = ~pi0626 & ~new_n32880_;
  assign new_n32896_ = pi0641 & ~new_n32895_;
  assign new_n32897_ = ~new_n32894_ & new_n32896_;
  assign new_n32898_ = pi0626 & ~new_n32887_;
  assign new_n32899_ = ~pi0626 & ~new_n32763_;
  assign new_n32900_ = ~pi0641 & ~new_n32899_;
  assign new_n32901_ = ~new_n32898_ & new_n32900_;
  assign new_n32902_ = pi1158 & ~new_n32901_;
  assign new_n32903_ = ~new_n32897_ & new_n32902_;
  assign new_n32904_ = ~new_n32893_ & ~new_n32903_;
  assign new_n32905_ = pi0788 & ~new_n32904_;
  assign new_n32906_ = ~new_n32876_ & ~new_n32905_;
  assign new_n32907_ = ~pi0628 & new_n32906_;
  assign new_n32908_ = ~new_n17968_ & new_n32887_;
  assign new_n32909_ = new_n17968_ & new_n32763_;
  assign new_n32910_ = ~new_n32908_ & ~new_n32909_;
  assign new_n32911_ = pi0628 & ~new_n32910_;
  assign new_n32912_ = ~pi1156 & ~new_n32911_;
  assign new_n32913_ = ~new_n32907_ & new_n32912_;
  assign new_n32914_ = ~new_n17734_ & new_n32880_;
  assign new_n32915_ = new_n17734_ & new_n32763_;
  assign new_n32916_ = ~new_n32914_ & ~new_n32915_;
  assign new_n32917_ = pi0628 & ~new_n32916_;
  assign new_n32918_ = ~pi0628 & new_n32763_;
  assign new_n32919_ = pi1156 & ~new_n32918_;
  assign new_n32920_ = ~new_n32917_ & new_n32919_;
  assign new_n32921_ = ~pi0629 & ~new_n32920_;
  assign new_n32922_ = ~new_n32913_ & new_n32921_;
  assign new_n32923_ = pi0628 & new_n32906_;
  assign new_n32924_ = ~pi0628 & ~new_n32910_;
  assign new_n32925_ = pi1156 & ~new_n32924_;
  assign new_n32926_ = ~new_n32923_ & new_n32925_;
  assign new_n32927_ = ~pi0628 & ~new_n32916_;
  assign new_n32928_ = pi0628 & new_n32763_;
  assign new_n32929_ = ~pi1156 & ~new_n32928_;
  assign new_n32930_ = ~new_n32927_ & new_n32929_;
  assign new_n32931_ = pi0629 & ~new_n32930_;
  assign new_n32932_ = ~new_n32926_ & new_n32931_;
  assign new_n32933_ = ~new_n32922_ & ~new_n32932_;
  assign new_n32934_ = pi0792 & ~new_n32933_;
  assign new_n32935_ = ~pi0792 & new_n32906_;
  assign new_n32936_ = ~new_n32934_ & ~new_n32935_;
  assign new_n32937_ = ~pi0647 & ~new_n32936_;
  assign new_n32938_ = ~new_n17762_ & ~new_n32910_;
  assign new_n32939_ = new_n17762_ & new_n32763_;
  assign new_n32940_ = ~new_n32938_ & ~new_n32939_;
  assign new_n32941_ = pi0647 & ~new_n32940_;
  assign new_n32942_ = ~pi1157 & ~new_n32941_;
  assign new_n32943_ = ~new_n32937_ & new_n32942_;
  assign new_n32944_ = ~pi0792 & new_n32916_;
  assign new_n32945_ = ~new_n32920_ & ~new_n32930_;
  assign new_n32946_ = pi0792 & ~new_n32945_;
  assign new_n32947_ = ~new_n32944_ & ~new_n32946_;
  assign new_n32948_ = pi0647 & new_n32947_;
  assign new_n32949_ = ~pi0647 & new_n32763_;
  assign new_n32950_ = pi1157 & ~new_n32949_;
  assign new_n32951_ = ~new_n32948_ & new_n32950_;
  assign new_n32952_ = ~pi0630 & ~new_n32951_;
  assign new_n32953_ = ~new_n32943_ & new_n32952_;
  assign new_n32954_ = pi0647 & ~new_n32936_;
  assign new_n32955_ = ~pi0647 & ~new_n32940_;
  assign new_n32956_ = pi1157 & ~new_n32955_;
  assign new_n32957_ = ~new_n32954_ & new_n32956_;
  assign new_n32958_ = ~pi0647 & new_n32947_;
  assign new_n32959_ = pi0647 & new_n32763_;
  assign new_n32960_ = ~pi1157 & ~new_n32959_;
  assign new_n32961_ = ~new_n32958_ & new_n32960_;
  assign new_n32962_ = pi0630 & ~new_n32961_;
  assign new_n32963_ = ~new_n32957_ & new_n32962_;
  assign new_n32964_ = ~new_n32953_ & ~new_n32963_;
  assign new_n32965_ = pi0787 & ~new_n32964_;
  assign new_n32966_ = ~pi0787 & ~new_n32936_;
  assign new_n32967_ = ~new_n32965_ & ~new_n32966_;
  assign new_n32968_ = ~pi0644 & ~new_n32967_;
  assign new_n32969_ = ~pi0787 & ~new_n32947_;
  assign new_n32970_ = ~new_n32951_ & ~new_n32961_;
  assign new_n32971_ = pi0787 & ~new_n32970_;
  assign new_n32972_ = ~new_n32969_ & ~new_n32971_;
  assign new_n32973_ = pi0644 & new_n32972_;
  assign new_n32974_ = ~pi0715 & ~new_n32973_;
  assign new_n32975_ = ~new_n32968_ & new_n32974_;
  assign new_n32976_ = new_n17804_ & ~new_n32763_;
  assign new_n32977_ = ~new_n17804_ & new_n32940_;
  assign new_n32978_ = ~new_n32976_ & ~new_n32977_;
  assign new_n32979_ = ~pi0644 & new_n32978_;
  assign new_n32980_ = pi0644 & new_n32763_;
  assign new_n32981_ = pi0715 & ~new_n32980_;
  assign new_n32982_ = ~new_n32979_ & new_n32981_;
  assign new_n32983_ = ~pi1160 & ~new_n32982_;
  assign new_n32984_ = ~new_n32975_ & new_n32983_;
  assign new_n32985_ = pi0644 & ~new_n32967_;
  assign new_n32986_ = ~pi0644 & new_n32972_;
  assign new_n32987_ = pi0715 & ~new_n32986_;
  assign new_n32988_ = ~new_n32985_ & new_n32987_;
  assign new_n32989_ = pi0644 & new_n32978_;
  assign new_n32990_ = ~pi0644 & new_n32763_;
  assign new_n32991_ = ~pi0715 & ~new_n32990_;
  assign new_n32992_ = ~new_n32989_ & new_n32991_;
  assign new_n32993_ = pi1160 & ~new_n32992_;
  assign new_n32994_ = ~new_n32988_ & new_n32993_;
  assign new_n32995_ = pi0790 & ~new_n32994_;
  assign new_n32996_ = ~new_n32984_ & new_n32995_;
  assign new_n32997_ = ~pi0790 & new_n32967_;
  assign new_n32998_ = ~po1038 & ~new_n32997_;
  assign new_n32999_ = ~new_n32996_ & new_n32998_;
  assign new_n33000_ = ~pi0194 & po1038;
  assign new_n33001_ = ~pi0832 & ~new_n33000_;
  assign new_n33002_ = ~new_n32999_ & new_n33001_;
  assign new_n33003_ = ~pi0194 & ~new_n2754_;
  assign new_n33004_ = pi0748 & new_n16913_;
  assign new_n33005_ = ~new_n33003_ & ~new_n33004_;
  assign new_n33006_ = ~new_n17858_ & ~new_n33005_;
  assign new_n33007_ = ~pi0785 & ~new_n33006_;
  assign new_n33008_ = ~new_n17863_ & ~new_n33005_;
  assign new_n33009_ = pi1155 & ~new_n33008_;
  assign new_n33010_ = ~new_n17866_ & new_n33006_;
  assign new_n33011_ = ~pi1155 & ~new_n33010_;
  assign new_n33012_ = ~new_n33009_ & ~new_n33011_;
  assign new_n33013_ = pi0785 & ~new_n33012_;
  assign new_n33014_ = ~new_n33007_ & ~new_n33013_;
  assign new_n33015_ = ~pi0781 & ~new_n33014_;
  assign new_n33016_ = ~new_n17873_ & new_n33014_;
  assign new_n33017_ = pi1154 & ~new_n33016_;
  assign new_n33018_ = ~new_n17876_ & new_n33014_;
  assign new_n33019_ = ~pi1154 & ~new_n33018_;
  assign new_n33020_ = ~new_n33017_ & ~new_n33019_;
  assign new_n33021_ = pi0781 & ~new_n33020_;
  assign new_n33022_ = ~new_n33015_ & ~new_n33021_;
  assign new_n33023_ = ~pi0789 & ~new_n33022_;
  assign new_n33024_ = pi0619 & new_n33022_;
  assign new_n33025_ = ~pi0619 & new_n33003_;
  assign new_n33026_ = pi1159 & ~new_n33025_;
  assign new_n33027_ = ~new_n33024_ & new_n33026_;
  assign new_n33028_ = ~pi0619 & new_n33022_;
  assign new_n33029_ = pi0619 & new_n33003_;
  assign new_n33030_ = ~pi1159 & ~new_n33029_;
  assign new_n33031_ = ~new_n33028_ & new_n33030_;
  assign new_n33032_ = ~new_n33027_ & ~new_n33031_;
  assign new_n33033_ = pi0789 & ~new_n33032_;
  assign new_n33034_ = ~new_n33023_ & ~new_n33033_;
  assign new_n33035_ = ~new_n17968_ & new_n33034_;
  assign new_n33036_ = new_n17968_ & new_n33003_;
  assign new_n33037_ = ~new_n33035_ & ~new_n33036_;
  assign new_n33038_ = ~new_n17762_ & ~new_n33037_;
  assign new_n33039_ = new_n17762_ & new_n33003_;
  assign new_n33040_ = ~new_n33038_ & ~new_n33039_;
  assign new_n33041_ = ~new_n20556_ & new_n33040_;
  assign new_n33042_ = pi0730 & new_n16915_;
  assign new_n33043_ = ~new_n33003_ & ~new_n33042_;
  assign new_n33044_ = ~pi0778 & new_n33043_;
  assign new_n33045_ = ~pi0625 & new_n33042_;
  assign new_n33046_ = ~new_n33043_ & ~new_n33045_;
  assign new_n33047_ = pi1153 & ~new_n33046_;
  assign new_n33048_ = ~pi1153 & ~new_n33003_;
  assign new_n33049_ = ~new_n33045_ & new_n33048_;
  assign new_n33050_ = ~new_n33047_ & ~new_n33049_;
  assign new_n33051_ = pi0778 & ~new_n33050_;
  assign new_n33052_ = ~new_n33044_ & ~new_n33051_;
  assign new_n33053_ = ~new_n17844_ & new_n33052_;
  assign new_n33054_ = ~new_n17846_ & new_n33053_;
  assign new_n33055_ = ~new_n17848_ & new_n33054_;
  assign new_n33056_ = ~new_n17980_ & new_n33055_;
  assign new_n33057_ = ~new_n18011_ & new_n33056_;
  assign new_n33058_ = ~pi0647 & new_n33057_;
  assign new_n33059_ = pi0647 & new_n33003_;
  assign new_n33060_ = ~pi1157 & ~new_n33059_;
  assign new_n33061_ = ~new_n33058_ & new_n33060_;
  assign new_n33062_ = pi0630 & new_n33061_;
  assign new_n33063_ = pi0647 & ~new_n33057_;
  assign new_n33064_ = ~pi0647 & ~new_n33003_;
  assign new_n33065_ = ~new_n33063_ & ~new_n33064_;
  assign new_n33066_ = new_n17801_ & ~new_n33065_;
  assign new_n33067_ = ~new_n33062_ & ~new_n33066_;
  assign new_n33068_ = ~new_n33041_ & new_n33067_;
  assign new_n33069_ = pi0787 & ~new_n33068_;
  assign new_n33070_ = pi0626 & ~new_n33034_;
  assign new_n33071_ = ~pi0626 & ~new_n33003_;
  assign new_n33072_ = new_n17731_ & ~new_n33071_;
  assign new_n33073_ = ~new_n33070_ & new_n33072_;
  assign new_n33074_ = new_n17856_ & new_n33055_;
  assign new_n33075_ = ~pi0626 & ~new_n33034_;
  assign new_n33076_ = pi0626 & ~new_n33003_;
  assign new_n33077_ = new_n17732_ & ~new_n33076_;
  assign new_n33078_ = ~new_n33075_ & new_n33077_;
  assign new_n33079_ = ~new_n33074_ & ~new_n33078_;
  assign new_n33080_ = ~new_n33073_ & new_n33079_;
  assign new_n33081_ = pi0788 & ~new_n33080_;
  assign new_n33082_ = ~new_n16639_ & ~new_n33043_;
  assign new_n33083_ = pi0625 & new_n33082_;
  assign new_n33084_ = new_n33005_ & ~new_n33082_;
  assign new_n33085_ = ~new_n33083_ & ~new_n33084_;
  assign new_n33086_ = new_n33048_ & ~new_n33085_;
  assign new_n33087_ = ~pi0608 & ~new_n33047_;
  assign new_n33088_ = ~new_n33086_ & new_n33087_;
  assign new_n33089_ = pi1153 & new_n33005_;
  assign new_n33090_ = ~new_n33083_ & new_n33089_;
  assign new_n33091_ = pi0608 & ~new_n33049_;
  assign new_n33092_ = ~new_n33090_ & new_n33091_;
  assign new_n33093_ = ~new_n33088_ & ~new_n33092_;
  assign new_n33094_ = pi0778 & ~new_n33093_;
  assign new_n33095_ = ~pi0778 & ~new_n33084_;
  assign new_n33096_ = ~new_n33094_ & ~new_n33095_;
  assign new_n33097_ = ~pi0609 & ~new_n33096_;
  assign new_n33098_ = pi0609 & new_n33052_;
  assign new_n33099_ = ~pi1155 & ~new_n33098_;
  assign new_n33100_ = ~new_n33097_ & new_n33099_;
  assign new_n33101_ = ~pi0660 & ~new_n33009_;
  assign new_n33102_ = ~new_n33100_ & new_n33101_;
  assign new_n33103_ = pi0609 & ~new_n33096_;
  assign new_n33104_ = ~pi0609 & new_n33052_;
  assign new_n33105_ = pi1155 & ~new_n33104_;
  assign new_n33106_ = ~new_n33103_ & new_n33105_;
  assign new_n33107_ = pi0660 & ~new_n33011_;
  assign new_n33108_ = ~new_n33106_ & new_n33107_;
  assign new_n33109_ = ~new_n33102_ & ~new_n33108_;
  assign new_n33110_ = pi0785 & ~new_n33109_;
  assign new_n33111_ = ~pi0785 & ~new_n33096_;
  assign new_n33112_ = ~new_n33110_ & ~new_n33111_;
  assign new_n33113_ = ~pi0618 & ~new_n33112_;
  assign new_n33114_ = pi0618 & new_n33053_;
  assign new_n33115_ = ~pi1154 & ~new_n33114_;
  assign new_n33116_ = ~new_n33113_ & new_n33115_;
  assign new_n33117_ = ~pi0627 & ~new_n33017_;
  assign new_n33118_ = ~new_n33116_ & new_n33117_;
  assign new_n33119_ = pi0618 & ~new_n33112_;
  assign new_n33120_ = ~pi0618 & new_n33053_;
  assign new_n33121_ = pi1154 & ~new_n33120_;
  assign new_n33122_ = ~new_n33119_ & new_n33121_;
  assign new_n33123_ = pi0627 & ~new_n33019_;
  assign new_n33124_ = ~new_n33122_ & new_n33123_;
  assign new_n33125_ = ~new_n33118_ & ~new_n33124_;
  assign new_n33126_ = pi0781 & ~new_n33125_;
  assign new_n33127_ = ~pi0781 & ~new_n33112_;
  assign new_n33128_ = ~new_n33126_ & ~new_n33127_;
  assign new_n33129_ = pi0619 & ~new_n33128_;
  assign new_n33130_ = ~pi0619 & new_n33054_;
  assign new_n33131_ = pi1159 & ~new_n33130_;
  assign new_n33132_ = ~new_n33129_ & new_n33131_;
  assign new_n33133_ = pi0648 & ~new_n33031_;
  assign new_n33134_ = ~new_n33132_ & new_n33133_;
  assign new_n33135_ = ~pi0619 & ~new_n33128_;
  assign new_n33136_ = pi0619 & new_n33054_;
  assign new_n33137_ = ~pi1159 & ~new_n33136_;
  assign new_n33138_ = ~new_n33135_ & new_n33137_;
  assign new_n33139_ = ~pi0648 & ~new_n33027_;
  assign new_n33140_ = ~new_n33138_ & new_n33139_;
  assign new_n33141_ = pi0789 & ~new_n33140_;
  assign new_n33142_ = ~new_n33134_ & new_n33141_;
  assign new_n33143_ = ~pi0789 & new_n33128_;
  assign new_n33144_ = new_n17969_ & ~new_n33143_;
  assign new_n33145_ = ~new_n33142_ & new_n33144_;
  assign new_n33146_ = ~new_n33081_ & ~new_n33145_;
  assign new_n33147_ = ~new_n20364_ & ~new_n33146_;
  assign new_n33148_ = new_n18008_ & ~new_n33037_;
  assign new_n33149_ = new_n20851_ & new_n33056_;
  assign new_n33150_ = ~new_n33148_ & ~new_n33149_;
  assign new_n33151_ = ~pi0629 & ~new_n33150_;
  assign new_n33152_ = new_n20855_ & new_n33056_;
  assign new_n33153_ = new_n18007_ & ~new_n33037_;
  assign new_n33154_ = ~new_n33152_ & ~new_n33153_;
  assign new_n33155_ = pi0629 & ~new_n33154_;
  assign new_n33156_ = ~new_n33151_ & ~new_n33155_;
  assign new_n33157_ = pi0792 & ~new_n33156_;
  assign new_n33158_ = ~new_n20360_ & ~new_n33157_;
  assign new_n33159_ = ~new_n33147_ & new_n33158_;
  assign new_n33160_ = ~new_n33069_ & ~new_n33159_;
  assign new_n33161_ = pi0644 & new_n33160_;
  assign new_n33162_ = ~pi0787 & ~new_n33057_;
  assign new_n33163_ = pi1157 & ~new_n33065_;
  assign new_n33164_ = ~new_n33061_ & ~new_n33163_;
  assign new_n33165_ = pi0787 & ~new_n33164_;
  assign new_n33166_ = ~new_n33162_ & ~new_n33165_;
  assign new_n33167_ = ~pi0644 & new_n33166_;
  assign new_n33168_ = pi0715 & ~new_n33167_;
  assign new_n33169_ = ~new_n33161_ & new_n33168_;
  assign new_n33170_ = ~new_n17804_ & ~new_n33040_;
  assign new_n33171_ = new_n17804_ & new_n33003_;
  assign new_n33172_ = ~new_n33170_ & ~new_n33171_;
  assign new_n33173_ = pi0644 & ~new_n33172_;
  assign new_n33174_ = ~pi0644 & new_n33003_;
  assign new_n33175_ = ~pi0715 & ~new_n33174_;
  assign new_n33176_ = ~new_n33173_ & new_n33175_;
  assign new_n33177_ = pi1160 & ~new_n33176_;
  assign new_n33178_ = ~new_n33169_ & new_n33177_;
  assign new_n33179_ = ~pi0644 & new_n33160_;
  assign new_n33180_ = pi0644 & new_n33166_;
  assign new_n33181_ = ~pi0715 & ~new_n33180_;
  assign new_n33182_ = ~new_n33179_ & new_n33181_;
  assign new_n33183_ = ~pi0644 & ~new_n33172_;
  assign new_n33184_ = pi0644 & new_n33003_;
  assign new_n33185_ = pi0715 & ~new_n33184_;
  assign new_n33186_ = ~new_n33183_ & new_n33185_;
  assign new_n33187_ = ~pi1160 & ~new_n33186_;
  assign new_n33188_ = ~new_n33182_ & new_n33187_;
  assign new_n33189_ = ~new_n33178_ & ~new_n33188_;
  assign new_n33190_ = pi0790 & ~new_n33189_;
  assign new_n33191_ = ~pi0790 & new_n33160_;
  assign new_n33192_ = pi0832 & ~new_n33191_;
  assign new_n33193_ = ~new_n33190_ & new_n33192_;
  assign po0351 = ~new_n33002_ & ~new_n33193_;
  assign new_n33195_ = ~new_n6221_ & new_n16194_;
  assign new_n33196_ = ~new_n11476_ & ~new_n33195_;
  assign new_n33197_ = ~new_n11473_ & new_n16171_;
  assign new_n33198_ = new_n16168_ & ~new_n16551_;
  assign new_n33199_ = ~new_n33197_ & ~new_n33198_;
  assign new_n33200_ = new_n33196_ & new_n33199_;
  assign new_n33201_ = pi0232 & ~new_n33200_;
  assign new_n33202_ = ~new_n16548_ & ~new_n33201_;
  assign new_n33203_ = pi0039 & ~new_n33202_;
  assign new_n33204_ = new_n13901_ & ~new_n16196_;
  assign new_n33205_ = ~pi0039 & ~new_n33204_;
  assign new_n33206_ = ~pi0138 & new_n16565_;
  assign new_n33207_ = ~pi0196 & new_n33206_;
  assign new_n33208_ = pi0195 & ~new_n33207_;
  assign new_n33209_ = new_n10200_ & ~new_n33208_;
  assign new_n33210_ = ~new_n33205_ & new_n33209_;
  assign new_n33211_ = ~new_n33203_ & new_n33210_;
  assign new_n33212_ = ~new_n9402_ & ~new_n16162_;
  assign new_n33213_ = pi0171 & new_n13721_;
  assign new_n33214_ = ~new_n33212_ & ~new_n33213_;
  assign new_n33215_ = pi0299 & ~new_n33214_;
  assign new_n33216_ = pi0192 & new_n16505_;
  assign new_n33217_ = ~pi0192 & new_n16493_;
  assign new_n33218_ = pi0232 & ~new_n33217_;
  assign new_n33219_ = ~new_n33216_ & new_n33218_;
  assign new_n33220_ = ~new_n33215_ & new_n33219_;
  assign new_n33221_ = new_n16497_ & ~new_n33220_;
  assign new_n33222_ = pi0192 & new_n16528_;
  assign new_n33223_ = ~pi0171 & new_n9074_;
  assign new_n33224_ = ~new_n16521_ & ~new_n33223_;
  assign new_n33225_ = new_n9069_ & ~new_n33224_;
  assign new_n33226_ = new_n9071_ & ~new_n33225_;
  assign new_n33227_ = ~pi0192 & new_n16514_;
  assign new_n33228_ = ~new_n33226_ & ~new_n33227_;
  assign new_n33229_ = ~new_n33222_ & new_n33228_;
  assign new_n33230_ = pi0232 & ~new_n33229_;
  assign new_n33231_ = ~new_n16520_ & ~new_n33230_;
  assign new_n33232_ = pi0039 & ~new_n33231_;
  assign new_n33233_ = new_n3211_ & ~new_n33232_;
  assign new_n33234_ = ~new_n33221_ & new_n33233_;
  assign new_n33235_ = ~pi0087 & ~new_n33234_;
  assign new_n33236_ = new_n16492_ & ~new_n33235_;
  assign new_n33237_ = ~pi0092 & ~new_n33236_;
  assign new_n33238_ = new_n16491_ & ~new_n33237_;
  assign new_n33239_ = ~pi0055 & ~new_n33238_;
  assign new_n33240_ = ~new_n16543_ & ~new_n33239_;
  assign new_n33241_ = new_n3298_ & ~new_n33240_;
  assign new_n33242_ = new_n9722_ & new_n33208_;
  assign new_n33243_ = ~new_n33241_ & new_n33242_;
  assign po0352 = new_n33211_ | new_n33243_;
  assign new_n33245_ = ~pi0170 & new_n9074_;
  assign new_n33246_ = ~new_n16521_ & ~new_n33245_;
  assign new_n33247_ = new_n9069_ & ~new_n33246_;
  assign new_n33248_ = new_n9071_ & ~new_n33247_;
  assign new_n33249_ = ~new_n16514_ & ~new_n33248_;
  assign new_n33250_ = pi0232 & ~new_n33249_;
  assign new_n33251_ = ~new_n16520_ & ~new_n33250_;
  assign new_n33252_ = pi0232 & new_n16528_;
  assign new_n33253_ = new_n33251_ & ~new_n33252_;
  assign new_n33254_ = pi0039 & ~new_n33253_;
  assign new_n33255_ = ~pi0038 & pi0194;
  assign new_n33256_ = ~new_n33254_ & new_n33255_;
  assign new_n33257_ = pi0039 & ~new_n33251_;
  assign new_n33258_ = ~pi0038 & ~pi0194;
  assign new_n33259_ = ~new_n33257_ & new_n33258_;
  assign new_n33260_ = ~new_n33256_ & ~new_n33259_;
  assign new_n33261_ = ~new_n16497_ & ~new_n33260_;
  assign new_n33262_ = ~new_n16505_ & new_n33256_;
  assign new_n33263_ = ~new_n16493_ & new_n33259_;
  assign new_n33264_ = ~new_n33262_ & ~new_n33263_;
  assign new_n33265_ = ~new_n9402_ & ~new_n16271_;
  assign new_n33266_ = pi0170 & new_n13721_;
  assign new_n33267_ = ~new_n33265_ & ~new_n33266_;
  assign new_n33268_ = pi0299 & ~new_n33267_;
  assign new_n33269_ = pi0232 & ~new_n33268_;
  assign new_n33270_ = ~new_n33264_ & new_n33269_;
  assign new_n33271_ = ~new_n33261_ & ~new_n33270_;
  assign new_n33272_ = ~pi0100 & ~new_n33271_;
  assign new_n33273_ = ~pi0087 & ~new_n33272_;
  assign new_n33274_ = new_n16492_ & ~new_n33273_;
  assign new_n33275_ = ~pi0092 & ~new_n33274_;
  assign new_n33276_ = new_n16491_ & ~new_n33275_;
  assign new_n33277_ = ~pi0055 & ~new_n33276_;
  assign new_n33278_ = ~new_n16543_ & ~new_n33277_;
  assign new_n33279_ = new_n3298_ & ~new_n33278_;
  assign new_n33280_ = new_n9722_ & ~new_n33279_;
  assign new_n33281_ = pi0196 & ~new_n33280_;
  assign new_n33282_ = ~pi0170 & new_n9546_;
  assign new_n33283_ = ~new_n16550_ & ~new_n33282_;
  assign new_n33284_ = new_n13130_ & ~new_n33283_;
  assign new_n33285_ = new_n13132_ & new_n16550_;
  assign new_n33286_ = pi0232 & ~new_n33285_;
  assign new_n33287_ = ~new_n33284_ & new_n33286_;
  assign new_n33288_ = ~new_n16548_ & ~new_n33287_;
  assign new_n33289_ = pi0299 & ~new_n33288_;
  assign new_n33290_ = ~new_n11474_ & ~new_n33289_;
  assign new_n33291_ = pi0039 & ~new_n33290_;
  assign new_n33292_ = new_n13901_ & ~new_n16272_;
  assign new_n33293_ = ~pi0039 & ~new_n33292_;
  assign new_n33294_ = ~pi0038 & ~new_n33293_;
  assign new_n33295_ = ~new_n33291_ & new_n33294_;
  assign new_n33296_ = ~pi0194 & ~new_n33295_;
  assign new_n33297_ = pi0039 & ~new_n33288_;
  assign new_n33298_ = new_n13901_ & new_n16331_;
  assign new_n33299_ = ~pi0039 & ~new_n33298_;
  assign new_n33300_ = ~pi0038 & ~new_n33299_;
  assign new_n33301_ = ~new_n33297_ & new_n33300_;
  assign new_n33302_ = pi0194 & ~new_n33301_;
  assign new_n33303_ = new_n10197_ & ~new_n33302_;
  assign new_n33304_ = ~new_n33296_ & new_n33303_;
  assign new_n33305_ = ~pi0196 & ~new_n33304_;
  assign new_n33306_ = ~new_n33206_ & ~new_n33305_;
  assign new_n33307_ = ~new_n33281_ & new_n33306_;
  assign new_n33308_ = pi0195 & ~pi0196;
  assign new_n33309_ = ~new_n33280_ & new_n33308_;
  assign new_n33310_ = ~new_n33304_ & ~new_n33308_;
  assign new_n33311_ = new_n33206_ & ~new_n33310_;
  assign new_n33312_ = ~new_n33309_ & new_n33311_;
  assign po0353 = new_n33307_ | new_n33312_;
  assign new_n33314_ = ~pi0767 & pi0947;
  assign new_n33315_ = ~pi0698 & new_n20915_;
  assign new_n33316_ = ~new_n33314_ & ~new_n33315_;
  assign new_n33317_ = new_n2754_ & ~new_n33316_;
  assign new_n33318_ = ~pi0197 & ~new_n2754_;
  assign new_n33319_ = pi0832 & ~new_n33318_;
  assign new_n33320_ = ~new_n33317_ & new_n33319_;
  assign new_n33321_ = pi0197 & ~new_n17549_;
  assign new_n33322_ = new_n17431_ & ~new_n33314_;
  assign new_n33323_ = pi0038 & ~new_n33322_;
  assign new_n33324_ = ~new_n33321_ & new_n33323_;
  assign new_n33325_ = ~pi0197 & ~new_n21000_;
  assign new_n33326_ = pi0197 & ~new_n21155_;
  assign new_n33327_ = pi0299 & ~new_n33326_;
  assign new_n33328_ = ~new_n33325_ & new_n33327_;
  assign new_n33329_ = ~pi0197 & ~new_n17326_;
  assign new_n33330_ = new_n21018_ & ~new_n33329_;
  assign new_n33331_ = ~pi0767 & ~new_n33330_;
  assign new_n33332_ = ~new_n33328_ & new_n33331_;
  assign new_n33333_ = ~pi0197 & pi0767;
  assign new_n33334_ = ~new_n17347_ & new_n33333_;
  assign new_n33335_ = pi0039 & ~new_n33334_;
  assign new_n33336_ = ~new_n33332_ & new_n33335_;
  assign new_n33337_ = new_n17260_ & new_n33314_;
  assign new_n33338_ = ~pi0197 & ~new_n17260_;
  assign new_n33339_ = ~pi0039 & ~new_n33338_;
  assign new_n33340_ = ~new_n33337_ & new_n33339_;
  assign new_n33341_ = ~pi0038 & ~new_n33340_;
  assign new_n33342_ = ~new_n33336_ & new_n33341_;
  assign new_n33343_ = ~new_n33324_ & ~new_n33342_;
  assign new_n33344_ = pi0698 & ~new_n33343_;
  assign new_n33345_ = ~new_n21066_ & new_n33340_;
  assign new_n33346_ = ~pi0197 & new_n21092_;
  assign new_n33347_ = pi0197 & new_n21108_;
  assign new_n33348_ = ~pi0767 & ~new_n33347_;
  assign new_n33349_ = ~new_n33346_ & new_n33348_;
  assign new_n33350_ = ~pi0197 & new_n21044_;
  assign new_n33351_ = pi0197 & new_n21060_;
  assign new_n33352_ = pi0299 & ~new_n33351_;
  assign new_n33353_ = ~new_n33350_ & new_n33352_;
  assign new_n33354_ = new_n21063_ & ~new_n33329_;
  assign new_n33355_ = pi0767 & ~new_n33354_;
  assign new_n33356_ = ~new_n33353_ & new_n33355_;
  assign new_n33357_ = pi0039 & ~new_n33356_;
  assign new_n33358_ = ~new_n33349_ & new_n33357_;
  assign new_n33359_ = ~new_n33345_ & ~new_n33358_;
  assign new_n33360_ = ~pi0038 & ~new_n33359_;
  assign new_n33361_ = pi0767 & pi0947;
  assign new_n33362_ = ~pi0039 & ~new_n33361_;
  assign new_n33363_ = new_n21237_ & new_n33362_;
  assign new_n33364_ = ~pi0197 & ~new_n17431_;
  assign new_n33365_ = pi0038 & ~new_n33364_;
  assign new_n33366_ = ~new_n33363_ & new_n33365_;
  assign new_n33367_ = ~pi0698 & ~new_n33366_;
  assign new_n33368_ = ~new_n33360_ & new_n33367_;
  assign new_n33369_ = ~new_n33344_ & ~new_n33368_;
  assign new_n33370_ = new_n10197_ & ~new_n33369_;
  assign new_n33371_ = ~pi0197 & ~new_n10197_;
  assign new_n33372_ = ~pi0832 & ~new_n33371_;
  assign new_n33373_ = ~new_n33370_ & new_n33372_;
  assign po0354 = ~new_n33320_ & ~new_n33373_;
  assign new_n33375_ = new_n3186_ & ~new_n17260_;
  assign new_n33376_ = new_n18873_ & ~new_n33375_;
  assign new_n33377_ = pi0198 & ~new_n33376_;
  assign new_n33378_ = pi0198 & ~new_n16941_;
  assign new_n33379_ = ~new_n6238_ & new_n33378_;
  assign new_n33380_ = pi0198 & ~new_n16636_;
  assign new_n33381_ = ~po1101 & ~new_n33380_;
  assign new_n33382_ = pi0198 & ~new_n16740_;
  assign new_n33383_ = po1101 & ~new_n33382_;
  assign new_n33384_ = ~new_n33381_ & ~new_n33383_;
  assign new_n33385_ = new_n6238_ & new_n33384_;
  assign new_n33386_ = ~new_n3057_ & ~new_n33385_;
  assign new_n33387_ = ~new_n33379_ & new_n33386_;
  assign new_n33388_ = new_n3057_ & ~new_n33380_;
  assign new_n33389_ = ~pi0223 & ~new_n33388_;
  assign new_n33390_ = ~new_n33387_ & new_n33389_;
  assign new_n33391_ = pi0198 & ~new_n16687_;
  assign new_n33392_ = ~new_n33381_ & new_n33391_;
  assign new_n33393_ = ~new_n6180_ & ~new_n16701_;
  assign new_n33394_ = new_n6180_ & ~new_n16660_;
  assign new_n33395_ = pi0198 & ~new_n33394_;
  assign new_n33396_ = ~new_n33393_ & new_n33395_;
  assign new_n33397_ = ~new_n6238_ & new_n33396_;
  assign new_n33398_ = ~new_n33392_ & ~new_n33397_;
  assign new_n33399_ = pi0223 & ~new_n33398_;
  assign new_n33400_ = ~pi0299 & ~new_n33399_;
  assign new_n33401_ = ~new_n33390_ & new_n33400_;
  assign new_n33402_ = ~new_n6212_ & new_n33378_;
  assign new_n33403_ = new_n6212_ & new_n33384_;
  assign new_n33404_ = ~new_n3467_ & ~new_n33403_;
  assign new_n33405_ = ~new_n33402_ & new_n33404_;
  assign new_n33406_ = new_n3467_ & ~new_n33380_;
  assign new_n33407_ = ~pi0215 & ~new_n33406_;
  assign new_n33408_ = ~new_n33405_ & new_n33407_;
  assign new_n33409_ = ~new_n6212_ & new_n33396_;
  assign new_n33410_ = ~new_n33392_ & ~new_n33409_;
  assign new_n33411_ = pi0215 & ~new_n33410_;
  assign new_n33412_ = pi0299 & ~new_n33411_;
  assign new_n33413_ = ~new_n33408_ & new_n33412_;
  assign new_n33414_ = new_n3272_ & new_n10982_;
  assign new_n33415_ = ~new_n33413_ & new_n33414_;
  assign new_n33416_ = ~new_n33401_ & new_n33415_;
  assign new_n33417_ = ~new_n33377_ & ~new_n33416_;
  assign new_n33418_ = new_n17762_ & ~new_n33417_;
  assign new_n33419_ = pi0198 & ~new_n3272_;
  assign new_n33420_ = pi0198 & ~new_n17193_;
  assign new_n33421_ = pi0603 & pi0633;
  assign new_n33422_ = ~new_n33420_ & ~new_n33421_;
  assign new_n33423_ = pi0198 & ~new_n17172_;
  assign new_n33424_ = ~pi0198 & new_n17212_;
  assign new_n33425_ = ~new_n33423_ & ~new_n33424_;
  assign new_n33426_ = new_n33421_ & new_n33425_;
  assign new_n33427_ = ~new_n33422_ & ~new_n33426_;
  assign new_n33428_ = pi0299 & new_n33427_;
  assign new_n33429_ = ~new_n17159_ & ~new_n17203_;
  assign new_n33430_ = pi0633 & ~new_n33429_;
  assign new_n33431_ = ~new_n17181_ & ~new_n33430_;
  assign new_n33432_ = ~new_n17223_ & ~new_n33431_;
  assign new_n33433_ = ~pi0299 & new_n33432_;
  assign new_n33434_ = ~pi0039 & ~new_n33433_;
  assign new_n33435_ = ~new_n33428_ & new_n33434_;
  assign new_n33436_ = pi0633 & new_n16636_;
  assign new_n33437_ = ~new_n16638_ & new_n33436_;
  assign new_n33438_ = ~new_n33380_ & ~new_n33437_;
  assign new_n33439_ = pi0603 & ~new_n33438_;
  assign new_n33440_ = ~pi0603 & new_n33380_;
  assign new_n33441_ = ~new_n33439_ & ~new_n33440_;
  assign new_n33442_ = ~new_n16707_ & new_n33441_;
  assign new_n33443_ = new_n6185_ & ~new_n33438_;
  assign new_n33444_ = ~new_n16660_ & new_n33437_;
  assign new_n33445_ = ~new_n33391_ & ~new_n33444_;
  assign new_n33446_ = ~new_n33443_ & new_n33445_;
  assign new_n33447_ = pi0603 & ~new_n33446_;
  assign new_n33448_ = new_n16707_ & ~new_n33440_;
  assign new_n33449_ = ~new_n33447_ & new_n33448_;
  assign new_n33450_ = ~new_n33442_ & ~new_n33449_;
  assign new_n33451_ = ~new_n6183_ & new_n33450_;
  assign new_n33452_ = ~new_n33391_ & ~new_n33447_;
  assign new_n33453_ = new_n6183_ & ~new_n33452_;
  assign new_n33454_ = ~new_n33451_ & ~new_n33453_;
  assign new_n33455_ = new_n6212_ & new_n33454_;
  assign new_n33456_ = pi0633 & new_n16976_;
  assign new_n33457_ = ~new_n33396_ & ~new_n33456_;
  assign new_n33458_ = ~new_n6183_ & ~new_n33457_;
  assign new_n33459_ = pi0198 & new_n16660_;
  assign new_n33460_ = ~new_n33444_ & ~new_n33459_;
  assign new_n33461_ = new_n17371_ & ~new_n33460_;
  assign new_n33462_ = ~new_n33458_ & ~new_n33461_;
  assign new_n33463_ = ~new_n6212_ & new_n33462_;
  assign new_n33464_ = pi0215 & ~new_n33463_;
  assign new_n33465_ = ~new_n33455_ & new_n33464_;
  assign new_n33466_ = pi0198 & new_n16738_;
  assign new_n33467_ = pi0633 & new_n16779_;
  assign new_n33468_ = ~new_n33466_ & ~new_n33467_;
  assign new_n33469_ = ~new_n6185_ & ~new_n33468_;
  assign new_n33470_ = ~new_n33443_ & ~new_n33469_;
  assign new_n33471_ = pi0603 & ~new_n33470_;
  assign new_n33472_ = ~pi0642 & ~new_n33471_;
  assign new_n33473_ = pi0642 & ~new_n33439_;
  assign new_n33474_ = new_n6179_ & ~new_n33473_;
  assign new_n33475_ = ~new_n33472_ & new_n33474_;
  assign new_n33476_ = ~new_n6179_ & new_n33439_;
  assign new_n33477_ = ~new_n33440_ & ~new_n33476_;
  assign new_n33478_ = ~new_n33475_ & new_n33477_;
  assign new_n33479_ = ~new_n6183_ & new_n33478_;
  assign new_n33480_ = ~pi0603 & new_n33382_;
  assign new_n33481_ = new_n6183_ & ~new_n33480_;
  assign new_n33482_ = ~new_n33471_ & new_n33481_;
  assign new_n33483_ = ~new_n33479_ & ~new_n33482_;
  assign new_n33484_ = new_n6212_ & new_n33483_;
  assign new_n33485_ = new_n6185_ & new_n33468_;
  assign new_n33486_ = ~new_n6185_ & new_n33438_;
  assign new_n33487_ = pi0603 & ~new_n16707_;
  assign new_n33488_ = ~new_n33486_ & new_n33487_;
  assign new_n33489_ = ~new_n33485_ & new_n33488_;
  assign new_n33490_ = pi0603 & ~new_n33468_;
  assign new_n33491_ = new_n16707_ & new_n33490_;
  assign new_n33492_ = pi0198 & new_n16816_;
  assign new_n33493_ = ~new_n33491_ & ~new_n33492_;
  assign new_n33494_ = ~new_n33489_ & new_n33493_;
  assign new_n33495_ = ~new_n6183_ & new_n33494_;
  assign new_n33496_ = new_n6183_ & ~new_n33466_;
  assign new_n33497_ = ~new_n33490_ & new_n33496_;
  assign new_n33498_ = ~new_n33495_ & ~new_n33497_;
  assign new_n33499_ = ~new_n6212_ & new_n33498_;
  assign new_n33500_ = ~new_n3467_ & ~new_n33499_;
  assign new_n33501_ = ~new_n33484_ & new_n33500_;
  assign new_n33502_ = new_n3467_ & new_n33441_;
  assign new_n33503_ = ~pi0215 & ~new_n33502_;
  assign new_n33504_ = ~new_n33501_ & new_n33503_;
  assign new_n33505_ = ~new_n33465_ & ~new_n33504_;
  assign new_n33506_ = pi0299 & ~new_n33505_;
  assign new_n33507_ = new_n6238_ & new_n33454_;
  assign new_n33508_ = ~new_n6238_ & new_n33462_;
  assign new_n33509_ = pi0223 & ~new_n33508_;
  assign new_n33510_ = ~new_n33507_ & new_n33509_;
  assign new_n33511_ = new_n6238_ & new_n33483_;
  assign new_n33512_ = ~new_n6238_ & new_n33498_;
  assign new_n33513_ = ~new_n3057_ & ~new_n33512_;
  assign new_n33514_ = ~new_n33511_ & new_n33513_;
  assign new_n33515_ = new_n3057_ & new_n33441_;
  assign new_n33516_ = ~pi0223 & ~new_n33515_;
  assign new_n33517_ = ~new_n33514_ & new_n33516_;
  assign new_n33518_ = ~new_n33510_ & ~new_n33517_;
  assign new_n33519_ = ~pi0299 & ~new_n33518_;
  assign new_n33520_ = pi0039 & ~new_n33519_;
  assign new_n33521_ = ~new_n33506_ & new_n33520_;
  assign new_n33522_ = ~new_n33435_ & ~new_n33521_;
  assign new_n33523_ = ~pi0038 & ~new_n33522_;
  assign new_n33524_ = pi0039 & pi0198;
  assign new_n33525_ = pi0038 & ~new_n33524_;
  assign new_n33526_ = pi0198 & ~new_n16647_;
  assign new_n33527_ = pi0633 & new_n16639_;
  assign new_n33528_ = new_n16647_ & new_n33527_;
  assign new_n33529_ = ~new_n33526_ & ~new_n33528_;
  assign new_n33530_ = ~pi0039 & ~new_n33529_;
  assign new_n33531_ = new_n33525_ & ~new_n33530_;
  assign new_n33532_ = new_n3272_ & ~new_n33531_;
  assign new_n33533_ = ~new_n33523_ & new_n33532_;
  assign new_n33534_ = ~new_n33419_ & ~new_n33533_;
  assign new_n33535_ = ~new_n17590_ & ~new_n33534_;
  assign new_n33536_ = new_n17590_ & ~new_n33417_;
  assign new_n33537_ = ~new_n33535_ & ~new_n33536_;
  assign new_n33538_ = ~pi0785 & ~new_n33537_;
  assign new_n33539_ = ~new_n17591_ & ~new_n33417_;
  assign new_n33540_ = pi0609 & new_n33535_;
  assign new_n33541_ = ~new_n33539_ & ~new_n33540_;
  assign new_n33542_ = pi1155 & ~new_n33541_;
  assign new_n33543_ = ~new_n17603_ & ~new_n33417_;
  assign new_n33544_ = ~pi0609 & new_n33535_;
  assign new_n33545_ = ~new_n33543_ & ~new_n33544_;
  assign new_n33546_ = ~pi1155 & ~new_n33545_;
  assign new_n33547_ = ~new_n33542_ & ~new_n33546_;
  assign new_n33548_ = pi0785 & ~new_n33547_;
  assign new_n33549_ = ~new_n33538_ & ~new_n33548_;
  assign new_n33550_ = ~pi0781 & ~new_n33549_;
  assign new_n33551_ = pi0618 & new_n33549_;
  assign new_n33552_ = ~pi0618 & new_n33417_;
  assign new_n33553_ = pi1154 & ~new_n33552_;
  assign new_n33554_ = ~new_n33551_ & new_n33553_;
  assign new_n33555_ = ~pi0618 & new_n33549_;
  assign new_n33556_ = pi0618 & new_n33417_;
  assign new_n33557_ = ~pi1154 & ~new_n33556_;
  assign new_n33558_ = ~new_n33555_ & new_n33557_;
  assign new_n33559_ = ~new_n33554_ & ~new_n33558_;
  assign new_n33560_ = pi0781 & ~new_n33559_;
  assign new_n33561_ = ~new_n33550_ & ~new_n33560_;
  assign new_n33562_ = ~pi0789 & ~new_n33561_;
  assign new_n33563_ = pi0619 & new_n33561_;
  assign new_n33564_ = ~pi0619 & new_n33417_;
  assign new_n33565_ = pi1159 & ~new_n33564_;
  assign new_n33566_ = ~new_n33563_ & new_n33565_;
  assign new_n33567_ = ~pi0619 & new_n33561_;
  assign new_n33568_ = pi0619 & new_n33417_;
  assign new_n33569_ = ~pi1159 & ~new_n33568_;
  assign new_n33570_ = ~new_n33567_ & new_n33569_;
  assign new_n33571_ = ~new_n33566_ & ~new_n33570_;
  assign new_n33572_ = pi0789 & ~new_n33571_;
  assign new_n33573_ = ~new_n33562_ & ~new_n33572_;
  assign new_n33574_ = ~new_n17968_ & new_n33573_;
  assign new_n33575_ = new_n17968_ & new_n33417_;
  assign new_n33576_ = ~new_n33574_ & ~new_n33575_;
  assign new_n33577_ = ~new_n17762_ & new_n33576_;
  assign new_n33578_ = ~new_n33418_ & ~new_n33577_;
  assign new_n33579_ = ~new_n20556_ & ~new_n33578_;
  assign new_n33580_ = ~new_n19279_ & new_n33417_;
  assign new_n33581_ = new_n17655_ & ~new_n33417_;
  assign new_n33582_ = ~new_n16812_ & ~new_n33380_;
  assign new_n33583_ = pi0634 & ~new_n33582_;
  assign new_n33584_ = ~new_n33380_ & ~new_n33583_;
  assign new_n33585_ = ~new_n6185_ & new_n33584_;
  assign new_n33586_ = pi0634 & new_n16814_;
  assign new_n33587_ = ~new_n33466_ & ~new_n33586_;
  assign new_n33588_ = new_n6185_ & new_n33587_;
  assign new_n33589_ = ~new_n33585_ & ~new_n33588_;
  assign new_n33590_ = ~new_n6180_ & ~new_n33589_;
  assign new_n33591_ = new_n6180_ & new_n33587_;
  assign new_n33592_ = new_n16631_ & ~new_n33591_;
  assign new_n33593_ = ~new_n33590_ & new_n33592_;
  assign new_n33594_ = pi0198 & new_n16777_;
  assign new_n33595_ = new_n6183_ & ~new_n33587_;
  assign new_n33596_ = ~new_n33594_ & ~new_n33595_;
  assign new_n33597_ = ~new_n33593_ & new_n33596_;
  assign new_n33598_ = ~new_n6238_ & ~new_n33597_;
  assign new_n33599_ = ~new_n6180_ & new_n33584_;
  assign new_n33600_ = new_n16631_ & ~new_n33599_;
  assign new_n33601_ = new_n6185_ & ~new_n33584_;
  assign new_n33602_ = ~new_n6185_ & ~new_n33587_;
  assign new_n33603_ = ~new_n33601_ & ~new_n33602_;
  assign new_n33604_ = new_n6180_ & new_n33603_;
  assign new_n33605_ = new_n33600_ & ~new_n33604_;
  assign new_n33606_ = new_n6183_ & ~new_n33603_;
  assign new_n33607_ = new_n6180_ & ~new_n33382_;
  assign new_n33608_ = ~new_n6180_ & ~new_n33380_;
  assign new_n33609_ = ~pi0680 & ~new_n33608_;
  assign new_n33610_ = ~new_n33607_ & new_n33609_;
  assign new_n33611_ = ~new_n33606_ & ~new_n33610_;
  assign new_n33612_ = ~new_n33605_ & new_n33611_;
  assign new_n33613_ = new_n6238_ & ~new_n33612_;
  assign new_n33614_ = ~new_n3057_ & ~new_n33613_;
  assign new_n33615_ = ~new_n33598_ & new_n33614_;
  assign new_n33616_ = pi0680 & new_n33583_;
  assign new_n33617_ = ~new_n33380_ & ~new_n33616_;
  assign new_n33618_ = new_n3057_ & new_n33617_;
  assign new_n33619_ = ~pi0223 & ~new_n33618_;
  assign new_n33620_ = ~new_n33615_ & new_n33619_;
  assign new_n33621_ = pi0634 & ~new_n16660_;
  assign new_n33622_ = new_n16812_ & new_n33621_;
  assign new_n33623_ = ~new_n33459_ & ~new_n33622_;
  assign new_n33624_ = ~new_n6185_ & ~new_n33623_;
  assign new_n33625_ = ~new_n33601_ & ~new_n33624_;
  assign new_n33626_ = new_n6180_ & new_n33625_;
  assign new_n33627_ = new_n33600_ & ~new_n33626_;
  assign new_n33628_ = ~pi0680 & new_n33396_;
  assign new_n33629_ = new_n33391_ & new_n33628_;
  assign new_n33630_ = new_n6183_ & ~new_n33625_;
  assign new_n33631_ = ~new_n33629_ & ~new_n33630_;
  assign new_n33632_ = ~new_n33627_ & new_n33631_;
  assign new_n33633_ = new_n6238_ & new_n33632_;
  assign new_n33634_ = new_n6185_ & new_n33623_;
  assign new_n33635_ = ~new_n33585_ & ~new_n33634_;
  assign new_n33636_ = ~new_n6180_ & ~new_n33635_;
  assign new_n33637_ = new_n6180_ & new_n33623_;
  assign new_n33638_ = new_n16631_ & ~new_n33637_;
  assign new_n33639_ = ~new_n33636_ & new_n33638_;
  assign new_n33640_ = new_n6183_ & ~new_n33623_;
  assign new_n33641_ = ~new_n33628_ & ~new_n33640_;
  assign new_n33642_ = ~new_n33639_ & new_n33641_;
  assign new_n33643_ = ~new_n6238_ & new_n33642_;
  assign new_n33644_ = pi0223 & ~new_n33643_;
  assign new_n33645_ = ~new_n33633_ & new_n33644_;
  assign new_n33646_ = ~pi0299 & ~new_n33645_;
  assign new_n33647_ = ~new_n33620_ & new_n33646_;
  assign new_n33648_ = new_n6212_ & ~new_n33612_;
  assign new_n33649_ = ~new_n6212_ & ~new_n33597_;
  assign new_n33650_ = ~new_n3467_ & ~new_n33649_;
  assign new_n33651_ = ~new_n33648_ & new_n33650_;
  assign new_n33652_ = new_n3467_ & new_n33617_;
  assign new_n33653_ = ~pi0215 & ~new_n33652_;
  assign new_n33654_ = ~new_n33651_ & new_n33653_;
  assign new_n33655_ = new_n6212_ & new_n33632_;
  assign new_n33656_ = ~new_n6212_ & new_n33642_;
  assign new_n33657_ = pi0215 & ~new_n33656_;
  assign new_n33658_ = ~new_n33655_ & new_n33657_;
  assign new_n33659_ = pi0299 & ~new_n33658_;
  assign new_n33660_ = ~new_n33654_ & new_n33659_;
  assign new_n33661_ = ~new_n33647_ & ~new_n33660_;
  assign new_n33662_ = pi0039 & ~new_n33661_;
  assign new_n33663_ = pi0634 & pi0680;
  assign new_n33664_ = ~pi0198 & new_n17168_;
  assign new_n33665_ = pi0198 & ~new_n17196_;
  assign new_n33666_ = ~new_n33664_ & ~new_n33665_;
  assign new_n33667_ = new_n33663_ & ~new_n33666_;
  assign new_n33668_ = new_n33420_ & ~new_n33663_;
  assign new_n33669_ = ~new_n33667_ & ~new_n33668_;
  assign new_n33670_ = pi0299 & ~new_n33669_;
  assign new_n33671_ = pi0198 & new_n17183_;
  assign new_n33672_ = ~new_n17132_ & new_n33663_;
  assign new_n33673_ = ~new_n33671_ & new_n33672_;
  assign new_n33674_ = ~new_n17181_ & ~new_n33673_;
  assign new_n33675_ = ~pi0299 & ~new_n33674_;
  assign new_n33676_ = ~pi0039 & ~new_n33675_;
  assign new_n33677_ = ~new_n33670_ & new_n33676_;
  assign new_n33678_ = ~new_n33662_ & ~new_n33677_;
  assign new_n33679_ = ~pi0038 & ~new_n33678_;
  assign new_n33680_ = pi0634 & new_n16914_;
  assign new_n33681_ = new_n16647_ & new_n33680_;
  assign new_n33682_ = ~new_n33526_ & ~new_n33681_;
  assign new_n33683_ = ~pi0039 & ~new_n33682_;
  assign new_n33684_ = new_n33525_ & ~new_n33683_;
  assign new_n33685_ = new_n3272_ & ~new_n33684_;
  assign new_n33686_ = ~new_n33679_ & new_n33685_;
  assign new_n33687_ = ~new_n33419_ & ~new_n33686_;
  assign new_n33688_ = ~pi0778 & ~new_n33687_;
  assign new_n33689_ = pi0625 & new_n33687_;
  assign new_n33690_ = ~pi0625 & new_n33417_;
  assign new_n33691_ = pi1153 & ~new_n33690_;
  assign new_n33692_ = ~new_n33689_ & new_n33691_;
  assign new_n33693_ = ~pi0625 & new_n33687_;
  assign new_n33694_ = pi0625 & new_n33417_;
  assign new_n33695_ = ~pi1153 & ~new_n33694_;
  assign new_n33696_ = ~new_n33693_ & new_n33695_;
  assign new_n33697_ = ~new_n33692_ & ~new_n33696_;
  assign new_n33698_ = pi0778 & ~new_n33697_;
  assign new_n33699_ = ~new_n33688_ & ~new_n33698_;
  assign new_n33700_ = ~new_n17618_ & new_n33699_;
  assign new_n33701_ = new_n17618_ & new_n33417_;
  assign new_n33702_ = ~new_n33700_ & ~new_n33701_;
  assign new_n33703_ = ~new_n17655_ & new_n33702_;
  assign new_n33704_ = ~new_n33581_ & ~new_n33703_;
  assign new_n33705_ = ~new_n17691_ & new_n33704_;
  assign new_n33706_ = ~new_n17734_ & new_n33705_;
  assign new_n33707_ = ~new_n33580_ & ~new_n33706_;
  assign new_n33708_ = ~pi0792 & new_n33707_;
  assign new_n33709_ = pi0628 & ~new_n33707_;
  assign new_n33710_ = ~pi0628 & new_n33417_;
  assign new_n33711_ = ~new_n33709_ & ~new_n33710_;
  assign new_n33712_ = pi1156 & new_n33711_;
  assign new_n33713_ = ~pi0628 & ~new_n33707_;
  assign new_n33714_ = pi0628 & new_n33417_;
  assign new_n33715_ = ~pi1156 & ~new_n33714_;
  assign new_n33716_ = ~new_n33713_ & new_n33715_;
  assign new_n33717_ = ~new_n33712_ & ~new_n33716_;
  assign new_n33718_ = pi0792 & ~new_n33717_;
  assign new_n33719_ = ~new_n33708_ & ~new_n33718_;
  assign new_n33720_ = ~pi0647 & new_n33719_;
  assign new_n33721_ = pi0647 & new_n33417_;
  assign new_n33722_ = ~pi1157 & ~new_n33721_;
  assign new_n33723_ = ~new_n33720_ & new_n33722_;
  assign new_n33724_ = pi0630 & new_n33723_;
  assign new_n33725_ = pi0647 & ~new_n33719_;
  assign new_n33726_ = ~pi0647 & ~new_n33417_;
  assign new_n33727_ = ~new_n33725_ & ~new_n33726_;
  assign new_n33728_ = new_n17801_ & ~new_n33727_;
  assign new_n33729_ = ~new_n33724_ & ~new_n33728_;
  assign new_n33730_ = ~new_n33579_ & new_n33729_;
  assign new_n33731_ = pi0787 & ~new_n33730_;
  assign new_n33732_ = ~new_n20567_ & new_n33576_;
  assign new_n33733_ = pi0629 & new_n33716_;
  assign new_n33734_ = new_n17759_ & new_n33711_;
  assign new_n33735_ = ~new_n33733_ & ~new_n33734_;
  assign new_n33736_ = ~new_n33732_ & new_n33735_;
  assign new_n33737_ = pi0792 & ~new_n33736_;
  assign new_n33738_ = pi0626 & ~new_n33573_;
  assign new_n33739_ = ~pi0626 & ~new_n33417_;
  assign new_n33740_ = new_n17731_ & ~new_n33739_;
  assign new_n33741_ = ~new_n33738_ & new_n33740_;
  assign new_n33742_ = new_n17691_ & new_n33417_;
  assign new_n33743_ = ~new_n33705_ & ~new_n33742_;
  assign new_n33744_ = new_n17856_ & ~new_n33743_;
  assign new_n33745_ = ~pi0626 & ~new_n33573_;
  assign new_n33746_ = pi0626 & ~new_n33417_;
  assign new_n33747_ = new_n17732_ & ~new_n33746_;
  assign new_n33748_ = ~new_n33745_ & new_n33747_;
  assign new_n33749_ = ~new_n33744_ & ~new_n33748_;
  assign new_n33750_ = ~new_n33741_ & new_n33749_;
  assign new_n33751_ = pi0788 & ~new_n33750_;
  assign new_n33752_ = ~pi0603 & ~new_n33666_;
  assign new_n33753_ = pi0198 & ~pi0665;
  assign new_n33754_ = pi0633 & ~new_n33753_;
  assign new_n33755_ = ~new_n33664_ & new_n33754_;
  assign new_n33756_ = new_n33425_ & new_n33755_;
  assign new_n33757_ = ~new_n17212_ & new_n33665_;
  assign new_n33758_ = ~pi0198 & ~pi0665;
  assign new_n33759_ = new_n17172_ & new_n33758_;
  assign new_n33760_ = ~pi0633 & ~new_n33759_;
  assign new_n33761_ = ~new_n33757_ & new_n33760_;
  assign new_n33762_ = pi0603 & ~new_n33761_;
  assign new_n33763_ = ~new_n33756_ & new_n33762_;
  assign new_n33764_ = ~new_n33752_ & ~new_n33763_;
  assign new_n33765_ = new_n33663_ & ~new_n33764_;
  assign new_n33766_ = new_n33427_ & ~new_n33663_;
  assign new_n33767_ = pi0299 & ~new_n33766_;
  assign new_n33768_ = ~new_n33765_ & new_n33767_;
  assign new_n33769_ = ~pi0634 & new_n17181_;
  assign new_n33770_ = pi0634 & new_n17184_;
  assign new_n33771_ = ~new_n17205_ & new_n33770_;
  assign new_n33772_ = ~new_n33769_ & ~new_n33771_;
  assign new_n33773_ = ~pi0633 & ~new_n33772_;
  assign new_n33774_ = pi0198 & ~pi0633;
  assign new_n33775_ = pi0634 & ~pi0665;
  assign new_n33776_ = ~new_n33774_ & new_n33775_;
  assign new_n33777_ = ~new_n17157_ & new_n33776_;
  assign new_n33778_ = pi0603 & ~new_n33777_;
  assign new_n33779_ = ~new_n33430_ & new_n33778_;
  assign new_n33780_ = ~new_n33773_ & new_n33779_;
  assign new_n33781_ = ~pi0603 & new_n33674_;
  assign new_n33782_ = pi0680 & ~new_n33781_;
  assign new_n33783_ = ~new_n33780_ & new_n33782_;
  assign new_n33784_ = ~pi0680 & new_n33432_;
  assign new_n33785_ = ~pi0299 & ~new_n33784_;
  assign new_n33786_ = ~new_n33783_ & new_n33785_;
  assign new_n33787_ = ~new_n33768_ & ~new_n33786_;
  assign new_n33788_ = ~pi0039 & ~new_n33787_;
  assign new_n33789_ = ~pi0680 & new_n33478_;
  assign new_n33790_ = new_n16846_ & new_n33775_;
  assign new_n33791_ = new_n33438_ & ~new_n33790_;
  assign new_n33792_ = new_n6185_ & ~new_n33791_;
  assign new_n33793_ = pi0634 & new_n16825_;
  assign new_n33794_ = new_n33468_ & ~new_n33793_;
  assign new_n33795_ = ~new_n6185_ & ~new_n33794_;
  assign new_n33796_ = ~new_n33792_ & ~new_n33795_;
  assign new_n33797_ = pi0603 & ~new_n33796_;
  assign new_n33798_ = ~pi0642 & new_n33797_;
  assign new_n33799_ = ~pi0603 & ~new_n33584_;
  assign new_n33800_ = pi0603 & ~new_n33791_;
  assign new_n33801_ = pi0642 & new_n33800_;
  assign new_n33802_ = ~new_n33799_ & ~new_n33801_;
  assign new_n33803_ = ~new_n33798_ & new_n33802_;
  assign new_n33804_ = new_n6179_ & ~new_n33803_;
  assign new_n33805_ = ~new_n33799_ & ~new_n33800_;
  assign new_n33806_ = ~new_n6179_ & ~new_n33805_;
  assign new_n33807_ = ~new_n16630_ & ~new_n33806_;
  assign new_n33808_ = ~new_n33804_ & new_n33807_;
  assign new_n33809_ = ~pi0603 & ~new_n33603_;
  assign new_n33810_ = new_n16630_ & ~new_n33809_;
  assign new_n33811_ = ~new_n33797_ & new_n33810_;
  assign new_n33812_ = ~new_n33808_ & ~new_n33811_;
  assign new_n33813_ = pi0680 & ~new_n33812_;
  assign new_n33814_ = ~new_n33789_ & ~new_n33813_;
  assign new_n33815_ = new_n6212_ & new_n33814_;
  assign new_n33816_ = ~pi0603 & new_n33589_;
  assign new_n33817_ = ~new_n16707_ & new_n33800_;
  assign new_n33818_ = ~new_n33488_ & ~new_n33817_;
  assign new_n33819_ = ~new_n6180_ & new_n33818_;
  assign new_n33820_ = ~new_n6185_ & ~new_n33818_;
  assign new_n33821_ = new_n33794_ & ~new_n33820_;
  assign new_n33822_ = ~new_n33819_ & ~new_n33821_;
  assign new_n33823_ = ~new_n33816_ & ~new_n33822_;
  assign new_n33824_ = new_n16631_ & ~new_n33823_;
  assign new_n33825_ = ~pi0680 & ~new_n33494_;
  assign new_n33826_ = ~new_n16639_ & ~new_n33587_;
  assign new_n33827_ = ~new_n33490_ & ~new_n33826_;
  assign new_n33828_ = new_n6183_ & ~new_n33827_;
  assign new_n33829_ = ~new_n33825_ & ~new_n33828_;
  assign new_n33830_ = ~new_n33824_ & new_n33829_;
  assign new_n33831_ = ~new_n6212_ & ~new_n33830_;
  assign new_n33832_ = ~new_n3467_ & ~new_n33831_;
  assign new_n33833_ = ~new_n33815_ & new_n33832_;
  assign new_n33834_ = new_n16790_ & new_n33583_;
  assign new_n33835_ = new_n33441_ & ~new_n33834_;
  assign new_n33836_ = new_n3467_ & new_n33835_;
  assign new_n33837_ = ~pi0215 & ~new_n33836_;
  assign new_n33838_ = ~new_n33833_ & new_n33837_;
  assign new_n33839_ = new_n16875_ & new_n33758_;
  assign new_n33840_ = new_n16638_ & new_n33753_;
  assign new_n33841_ = ~new_n33459_ & ~new_n33840_;
  assign new_n33842_ = ~new_n33839_ & new_n33841_;
  assign new_n33843_ = pi0634 & ~new_n33842_;
  assign new_n33844_ = ~pi0634 & new_n33459_;
  assign new_n33845_ = ~new_n33444_ & ~new_n33844_;
  assign new_n33846_ = ~new_n33843_ & new_n33845_;
  assign new_n33847_ = ~new_n6185_ & ~new_n33846_;
  assign new_n33848_ = ~new_n33792_ & ~new_n33847_;
  assign new_n33849_ = pi0603 & ~new_n33848_;
  assign new_n33850_ = new_n16707_ & ~new_n33799_;
  assign new_n33851_ = ~new_n33849_ & new_n33850_;
  assign new_n33852_ = ~new_n16707_ & new_n33805_;
  assign new_n33853_ = new_n16631_ & ~new_n33852_;
  assign new_n33854_ = ~new_n33851_ & new_n33853_;
  assign new_n33855_ = ~pi0680 & new_n33450_;
  assign new_n33856_ = ~pi0603 & ~new_n33625_;
  assign new_n33857_ = ~new_n33849_ & ~new_n33856_;
  assign new_n33858_ = new_n6183_ & ~new_n33857_;
  assign new_n33859_ = ~new_n33855_ & ~new_n33858_;
  assign new_n33860_ = ~new_n33854_ & new_n33859_;
  assign new_n33861_ = new_n6212_ & new_n33860_;
  assign new_n33862_ = ~pi0603 & new_n33635_;
  assign new_n33863_ = ~new_n33820_ & ~new_n33862_;
  assign new_n33864_ = pi0603 & ~new_n33846_;
  assign new_n33865_ = new_n16707_ & new_n33864_;
  assign new_n33866_ = ~new_n33818_ & ~new_n33846_;
  assign new_n33867_ = ~new_n33865_ & ~new_n33866_;
  assign new_n33868_ = new_n33863_ & new_n33867_;
  assign new_n33869_ = new_n16631_ & ~new_n33868_;
  assign new_n33870_ = ~pi0680 & ~new_n33457_;
  assign new_n33871_ = ~pi0603 & ~new_n33623_;
  assign new_n33872_ = ~new_n33864_ & ~new_n33871_;
  assign new_n33873_ = new_n6183_ & ~new_n33872_;
  assign new_n33874_ = ~new_n33870_ & ~new_n33873_;
  assign new_n33875_ = ~new_n33869_ & new_n33874_;
  assign new_n33876_ = ~new_n6212_ & new_n33875_;
  assign new_n33877_ = pi0215 & ~new_n33876_;
  assign new_n33878_ = ~new_n33861_ & new_n33877_;
  assign new_n33879_ = ~new_n33838_ & ~new_n33878_;
  assign new_n33880_ = pi0299 & ~new_n33879_;
  assign new_n33881_ = new_n6238_ & new_n33814_;
  assign new_n33882_ = ~new_n6238_ & ~new_n33830_;
  assign new_n33883_ = ~new_n3057_ & ~new_n33882_;
  assign new_n33884_ = ~new_n33881_ & new_n33883_;
  assign new_n33885_ = new_n3057_ & new_n33835_;
  assign new_n33886_ = ~pi0223 & ~new_n33885_;
  assign new_n33887_ = ~new_n33884_ & new_n33886_;
  assign new_n33888_ = new_n6238_ & new_n33860_;
  assign new_n33889_ = ~new_n6238_ & new_n33875_;
  assign new_n33890_ = pi0223 & ~new_n33889_;
  assign new_n33891_ = ~new_n33888_ & new_n33890_;
  assign new_n33892_ = ~new_n33887_ & ~new_n33891_;
  assign new_n33893_ = ~pi0299 & ~new_n33892_;
  assign new_n33894_ = pi0039 & ~new_n33893_;
  assign new_n33895_ = ~new_n33880_ & new_n33894_;
  assign new_n33896_ = ~new_n33788_ & ~new_n33895_;
  assign new_n33897_ = ~pi0038 & ~new_n33896_;
  assign new_n33898_ = pi0634 & new_n17247_;
  assign new_n33899_ = new_n33529_ & ~new_n33898_;
  assign new_n33900_ = ~pi0039 & ~new_n33899_;
  assign new_n33901_ = new_n33525_ & ~new_n33900_;
  assign new_n33902_ = new_n3272_ & ~new_n33901_;
  assign new_n33903_ = ~new_n33897_ & new_n33902_;
  assign new_n33904_ = ~new_n33419_ & ~new_n33903_;
  assign new_n33905_ = ~pi0625 & new_n33904_;
  assign new_n33906_ = pi0625 & new_n33534_;
  assign new_n33907_ = ~pi1153 & ~new_n33906_;
  assign new_n33908_ = ~new_n33905_ & new_n33907_;
  assign new_n33909_ = ~pi0608 & ~new_n33692_;
  assign new_n33910_ = ~new_n33908_ & new_n33909_;
  assign new_n33911_ = pi0625 & new_n33904_;
  assign new_n33912_ = ~pi0625 & new_n33534_;
  assign new_n33913_ = pi1153 & ~new_n33912_;
  assign new_n33914_ = ~new_n33911_ & new_n33913_;
  assign new_n33915_ = pi0608 & ~new_n33696_;
  assign new_n33916_ = ~new_n33914_ & new_n33915_;
  assign new_n33917_ = ~new_n33910_ & ~new_n33916_;
  assign new_n33918_ = pi0778 & ~new_n33917_;
  assign new_n33919_ = ~pi0778 & new_n33904_;
  assign new_n33920_ = ~new_n33918_ & ~new_n33919_;
  assign new_n33921_ = ~pi0609 & ~new_n33920_;
  assign new_n33922_ = pi0609 & new_n33699_;
  assign new_n33923_ = ~pi1155 & ~new_n33922_;
  assign new_n33924_ = ~new_n33921_ & new_n33923_;
  assign new_n33925_ = ~pi0660 & ~new_n33542_;
  assign new_n33926_ = ~new_n33924_ & new_n33925_;
  assign new_n33927_ = pi0609 & ~new_n33920_;
  assign new_n33928_ = ~pi0609 & new_n33699_;
  assign new_n33929_ = pi1155 & ~new_n33928_;
  assign new_n33930_ = ~new_n33927_ & new_n33929_;
  assign new_n33931_ = pi0660 & ~new_n33546_;
  assign new_n33932_ = ~new_n33930_ & new_n33931_;
  assign new_n33933_ = ~new_n33926_ & ~new_n33932_;
  assign new_n33934_ = pi0785 & ~new_n33933_;
  assign new_n33935_ = ~pi0785 & ~new_n33920_;
  assign new_n33936_ = ~new_n33934_ & ~new_n33935_;
  assign new_n33937_ = ~pi0618 & ~new_n33936_;
  assign new_n33938_ = pi0618 & ~new_n33702_;
  assign new_n33939_ = ~pi1154 & ~new_n33938_;
  assign new_n33940_ = ~new_n33937_ & new_n33939_;
  assign new_n33941_ = ~pi0627 & ~new_n33554_;
  assign new_n33942_ = ~new_n33940_ & new_n33941_;
  assign new_n33943_ = pi0618 & ~new_n33936_;
  assign new_n33944_ = ~pi0618 & ~new_n33702_;
  assign new_n33945_ = pi1154 & ~new_n33944_;
  assign new_n33946_ = ~new_n33943_ & new_n33945_;
  assign new_n33947_ = pi0627 & ~new_n33558_;
  assign new_n33948_ = ~new_n33946_ & new_n33947_;
  assign new_n33949_ = ~new_n33942_ & ~new_n33948_;
  assign new_n33950_ = pi0781 & ~new_n33949_;
  assign new_n33951_ = ~pi0781 & ~new_n33936_;
  assign new_n33952_ = ~new_n33950_ & ~new_n33951_;
  assign new_n33953_ = pi0619 & ~new_n33952_;
  assign new_n33954_ = ~pi0619 & new_n33704_;
  assign new_n33955_ = pi1159 & ~new_n33954_;
  assign new_n33956_ = ~new_n33953_ & new_n33955_;
  assign new_n33957_ = pi0648 & ~new_n33570_;
  assign new_n33958_ = ~new_n33956_ & new_n33957_;
  assign new_n33959_ = ~pi0619 & ~new_n33952_;
  assign new_n33960_ = pi0619 & new_n33704_;
  assign new_n33961_ = ~pi1159 & ~new_n33960_;
  assign new_n33962_ = ~new_n33959_ & new_n33961_;
  assign new_n33963_ = ~pi0648 & ~new_n33566_;
  assign new_n33964_ = ~new_n33962_ & new_n33963_;
  assign new_n33965_ = pi0789 & ~new_n33964_;
  assign new_n33966_ = ~new_n33958_ & new_n33965_;
  assign new_n33967_ = ~pi0789 & new_n33952_;
  assign new_n33968_ = new_n17969_ & ~new_n33967_;
  assign new_n33969_ = ~new_n33966_ & new_n33968_;
  assign new_n33970_ = ~new_n33751_ & ~new_n33969_;
  assign new_n33971_ = ~new_n33737_ & ~new_n33970_;
  assign new_n33972_ = new_n20364_ & new_n33736_;
  assign new_n33973_ = ~new_n20360_ & ~new_n33972_;
  assign new_n33974_ = ~new_n33971_ & new_n33973_;
  assign new_n33975_ = ~new_n33731_ & ~new_n33974_;
  assign new_n33976_ = ~pi0790 & ~new_n33975_;
  assign new_n33977_ = ~pi0644 & new_n33975_;
  assign new_n33978_ = ~pi0787 & ~new_n33719_;
  assign new_n33979_ = pi1157 & ~new_n33727_;
  assign new_n33980_ = ~new_n33723_ & ~new_n33979_;
  assign new_n33981_ = pi0787 & ~new_n33980_;
  assign new_n33982_ = ~new_n33978_ & ~new_n33981_;
  assign new_n33983_ = pi0644 & new_n33982_;
  assign new_n33984_ = ~pi0715 & ~new_n33983_;
  assign new_n33985_ = ~new_n33977_ & new_n33984_;
  assign new_n33986_ = ~new_n17804_ & new_n33578_;
  assign new_n33987_ = new_n17804_ & new_n33417_;
  assign new_n33988_ = ~new_n33986_ & ~new_n33987_;
  assign new_n33989_ = ~pi0644 & ~new_n33988_;
  assign new_n33990_ = pi0644 & new_n33417_;
  assign new_n33991_ = pi0715 & ~new_n33990_;
  assign new_n33992_ = ~new_n33989_ & new_n33991_;
  assign new_n33993_ = ~pi1160 & ~new_n33992_;
  assign new_n33994_ = ~new_n33985_ & new_n33993_;
  assign new_n33995_ = pi0644 & new_n33975_;
  assign new_n33996_ = ~pi0644 & new_n33982_;
  assign new_n33997_ = pi0715 & ~new_n33996_;
  assign new_n33998_ = ~new_n33995_ & new_n33997_;
  assign new_n33999_ = pi0644 & ~new_n33988_;
  assign new_n34000_ = ~pi0644 & new_n33417_;
  assign new_n34001_ = ~pi0715 & ~new_n34000_;
  assign new_n34002_ = ~new_n33999_ & new_n34001_;
  assign new_n34003_ = pi1160 & ~new_n34002_;
  assign new_n34004_ = ~new_n33998_ & new_n34003_;
  assign new_n34005_ = pi0790 & ~new_n34004_;
  assign new_n34006_ = ~new_n33994_ & new_n34005_;
  assign new_n34007_ = ~new_n33976_ & ~new_n34006_;
  assign new_n34008_ = ~po1038 & ~new_n34007_;
  assign new_n34009_ = pi0198 & po1038;
  assign po0355 = new_n34008_ | new_n34009_;
  assign new_n34011_ = pi0199 & ~new_n17558_;
  assign new_n34012_ = ~pi0617 & ~new_n34011_;
  assign new_n34013_ = ~pi0199 & ~new_n19369_;
  assign new_n34014_ = new_n19375_ & ~new_n34013_;
  assign new_n34015_ = pi0199 & new_n17393_;
  assign new_n34016_ = ~pi0199 & ~new_n17426_;
  assign new_n34017_ = ~pi0038 & ~new_n34016_;
  assign new_n34018_ = ~new_n34015_ & new_n34017_;
  assign new_n34019_ = ~new_n34014_ & ~new_n34018_;
  assign new_n34020_ = new_n3272_ & ~new_n34019_;
  assign new_n34021_ = pi0199 & ~new_n3272_;
  assign new_n34022_ = pi0617 & ~new_n34021_;
  assign new_n34023_ = ~new_n34020_ & new_n34022_;
  assign new_n34024_ = ~new_n34012_ & ~new_n34023_;
  assign new_n34025_ = ~pi0637 & new_n34024_;
  assign new_n34026_ = pi0199 & new_n19388_;
  assign new_n34027_ = new_n3272_ & ~new_n24548_;
  assign new_n34028_ = ~pi0199 & ~new_n34027_;
  assign new_n34029_ = ~pi0617 & ~new_n19384_;
  assign new_n34030_ = ~new_n34028_ & new_n34029_;
  assign new_n34031_ = ~new_n34026_ & new_n34030_;
  assign new_n34032_ = new_n3272_ & new_n19406_;
  assign new_n34033_ = ~pi0199 & ~new_n34032_;
  assign new_n34034_ = pi0199 & new_n19414_;
  assign new_n34035_ = pi0617 & ~new_n34034_;
  assign new_n34036_ = ~new_n34033_ & new_n34035_;
  assign new_n34037_ = ~new_n34021_ & ~new_n34036_;
  assign new_n34038_ = ~new_n34031_ & new_n34037_;
  assign new_n34039_ = pi0637 & ~new_n34038_;
  assign new_n34040_ = ~new_n34025_ & ~new_n34039_;
  assign new_n34041_ = ~pi0625 & new_n34040_;
  assign new_n34042_ = pi0625 & ~new_n34024_;
  assign new_n34043_ = ~pi1153 & ~new_n34042_;
  assign new_n34044_ = ~new_n34041_ & new_n34043_;
  assign new_n34045_ = ~pi0637 & ~new_n34011_;
  assign new_n34046_ = ~pi0199 & ~new_n17431_;
  assign new_n34047_ = new_n19956_ & ~new_n34046_;
  assign new_n34048_ = pi0199 & ~new_n17533_;
  assign new_n34049_ = ~pi0199 & ~new_n17483_;
  assign new_n34050_ = pi0039 & ~new_n34049_;
  assign new_n34051_ = ~new_n34048_ & new_n34050_;
  assign new_n34052_ = ~pi0199 & new_n17233_;
  assign new_n34053_ = pi0199 & ~new_n17200_;
  assign new_n34054_ = ~pi0039 & ~new_n34053_;
  assign new_n34055_ = ~new_n34052_ & new_n34054_;
  assign new_n34056_ = ~pi0038 & ~new_n34055_;
  assign new_n34057_ = ~new_n34051_ & new_n34056_;
  assign new_n34058_ = ~new_n34047_ & ~new_n34057_;
  assign new_n34059_ = new_n3272_ & ~new_n34058_;
  assign new_n34060_ = pi0637 & ~new_n34021_;
  assign new_n34061_ = ~new_n34059_ & new_n34060_;
  assign new_n34062_ = ~new_n34045_ & ~new_n34061_;
  assign new_n34063_ = pi0625 & ~new_n34062_;
  assign new_n34064_ = ~pi0625 & ~new_n34011_;
  assign new_n34065_ = pi1153 & ~new_n34064_;
  assign new_n34066_ = ~new_n34063_ & new_n34065_;
  assign new_n34067_ = ~pi0608 & ~new_n34066_;
  assign new_n34068_ = ~new_n34044_ & new_n34067_;
  assign new_n34069_ = pi0625 & new_n34040_;
  assign new_n34070_ = ~pi0625 & ~new_n34024_;
  assign new_n34071_ = pi1153 & ~new_n34070_;
  assign new_n34072_ = ~new_n34069_ & new_n34071_;
  assign new_n34073_ = ~pi0625 & ~new_n34062_;
  assign new_n34074_ = pi0625 & ~new_n34011_;
  assign new_n34075_ = ~pi1153 & ~new_n34074_;
  assign new_n34076_ = ~new_n34073_ & new_n34075_;
  assign new_n34077_ = pi0608 & ~new_n34076_;
  assign new_n34078_ = ~new_n34072_ & new_n34077_;
  assign new_n34079_ = ~new_n34068_ & ~new_n34078_;
  assign new_n34080_ = pi0778 & ~new_n34079_;
  assign new_n34081_ = ~pi0778 & new_n34040_;
  assign new_n34082_ = ~new_n34080_ & ~new_n34081_;
  assign new_n34083_ = ~pi0609 & ~new_n34082_;
  assign new_n34084_ = ~pi0778 & new_n34062_;
  assign new_n34085_ = ~new_n34066_ & ~new_n34076_;
  assign new_n34086_ = pi0778 & ~new_n34085_;
  assign new_n34087_ = ~new_n34084_ & ~new_n34086_;
  assign new_n34088_ = pi0609 & new_n34087_;
  assign new_n34089_ = ~pi1155 & ~new_n34088_;
  assign new_n34090_ = ~new_n34083_ & new_n34089_;
  assign new_n34091_ = ~new_n17590_ & ~new_n34024_;
  assign new_n34092_ = new_n17590_ & ~new_n34011_;
  assign new_n34093_ = ~new_n34091_ & ~new_n34092_;
  assign new_n34094_ = pi0609 & ~new_n34093_;
  assign new_n34095_ = ~pi0609 & ~new_n34011_;
  assign new_n34096_ = pi1155 & ~new_n34095_;
  assign new_n34097_ = ~new_n34094_ & new_n34096_;
  assign new_n34098_ = ~pi0660 & ~new_n34097_;
  assign new_n34099_ = ~new_n34090_ & new_n34098_;
  assign new_n34100_ = pi0609 & ~new_n34082_;
  assign new_n34101_ = ~pi0609 & new_n34087_;
  assign new_n34102_ = pi1155 & ~new_n34101_;
  assign new_n34103_ = ~new_n34100_ & new_n34102_;
  assign new_n34104_ = ~pi0609 & ~new_n34093_;
  assign new_n34105_ = pi0609 & ~new_n34011_;
  assign new_n34106_ = ~pi1155 & ~new_n34105_;
  assign new_n34107_ = ~new_n34104_ & new_n34106_;
  assign new_n34108_ = pi0660 & ~new_n34107_;
  assign new_n34109_ = ~new_n34103_ & new_n34108_;
  assign new_n34110_ = ~new_n34099_ & ~new_n34109_;
  assign new_n34111_ = pi0785 & ~new_n34110_;
  assign new_n34112_ = ~pi0785 & ~new_n34082_;
  assign new_n34113_ = ~new_n34111_ & ~new_n34112_;
  assign new_n34114_ = ~pi0618 & ~new_n34113_;
  assign new_n34115_ = new_n17618_ & ~new_n34011_;
  assign new_n34116_ = ~new_n17618_ & new_n34087_;
  assign new_n34117_ = ~new_n34115_ & ~new_n34116_;
  assign new_n34118_ = pi0618 & ~new_n34117_;
  assign new_n34119_ = ~pi1154 & ~new_n34118_;
  assign new_n34120_ = ~new_n34114_ & new_n34119_;
  assign new_n34121_ = ~pi0785 & new_n34093_;
  assign new_n34122_ = ~new_n34097_ & ~new_n34107_;
  assign new_n34123_ = pi0785 & ~new_n34122_;
  assign new_n34124_ = ~new_n34121_ & ~new_n34123_;
  assign new_n34125_ = pi0618 & new_n34124_;
  assign new_n34126_ = ~pi0618 & ~new_n34011_;
  assign new_n34127_ = pi1154 & ~new_n34126_;
  assign new_n34128_ = ~new_n34125_ & new_n34127_;
  assign new_n34129_ = ~pi0627 & ~new_n34128_;
  assign new_n34130_ = ~new_n34120_ & new_n34129_;
  assign new_n34131_ = pi0618 & ~new_n34113_;
  assign new_n34132_ = ~pi0618 & ~new_n34117_;
  assign new_n34133_ = pi1154 & ~new_n34132_;
  assign new_n34134_ = ~new_n34131_ & new_n34133_;
  assign new_n34135_ = ~pi0618 & new_n34124_;
  assign new_n34136_ = pi0618 & ~new_n34011_;
  assign new_n34137_ = ~pi1154 & ~new_n34136_;
  assign new_n34138_ = ~new_n34135_ & new_n34137_;
  assign new_n34139_ = pi0627 & ~new_n34138_;
  assign new_n34140_ = ~new_n34134_ & new_n34139_;
  assign new_n34141_ = ~new_n34130_ & ~new_n34140_;
  assign new_n34142_ = pi0781 & ~new_n34141_;
  assign new_n34143_ = ~pi0781 & ~new_n34113_;
  assign new_n34144_ = ~new_n34142_ & ~new_n34143_;
  assign new_n34145_ = ~pi0619 & ~new_n34144_;
  assign new_n34146_ = ~new_n17655_ & new_n34117_;
  assign new_n34147_ = new_n17655_ & new_n34011_;
  assign new_n34148_ = ~new_n34146_ & ~new_n34147_;
  assign new_n34149_ = pi0619 & new_n34148_;
  assign new_n34150_ = ~pi1159 & ~new_n34149_;
  assign new_n34151_ = ~new_n34145_ & new_n34150_;
  assign new_n34152_ = ~pi0781 & ~new_n34124_;
  assign new_n34153_ = ~new_n34128_ & ~new_n34138_;
  assign new_n34154_ = pi0781 & ~new_n34153_;
  assign new_n34155_ = ~new_n34152_ & ~new_n34154_;
  assign new_n34156_ = pi0619 & new_n34155_;
  assign new_n34157_ = ~pi0619 & ~new_n34011_;
  assign new_n34158_ = pi1159 & ~new_n34157_;
  assign new_n34159_ = ~new_n34156_ & new_n34158_;
  assign new_n34160_ = ~pi0648 & ~new_n34159_;
  assign new_n34161_ = ~new_n34151_ & new_n34160_;
  assign new_n34162_ = pi0619 & ~new_n34144_;
  assign new_n34163_ = ~pi0619 & new_n34148_;
  assign new_n34164_ = pi1159 & ~new_n34163_;
  assign new_n34165_ = ~new_n34162_ & new_n34164_;
  assign new_n34166_ = ~pi0619 & new_n34155_;
  assign new_n34167_ = pi0619 & ~new_n34011_;
  assign new_n34168_ = ~pi1159 & ~new_n34167_;
  assign new_n34169_ = ~new_n34166_ & new_n34168_;
  assign new_n34170_ = pi0648 & ~new_n34169_;
  assign new_n34171_ = ~new_n34165_ & new_n34170_;
  assign new_n34172_ = ~new_n34161_ & ~new_n34171_;
  assign new_n34173_ = pi0789 & ~new_n34172_;
  assign new_n34174_ = ~pi0789 & ~new_n34144_;
  assign new_n34175_ = ~new_n34173_ & ~new_n34174_;
  assign new_n34176_ = ~pi0788 & new_n34175_;
  assign new_n34177_ = ~pi0626 & new_n34175_;
  assign new_n34178_ = new_n17691_ & ~new_n34011_;
  assign new_n34179_ = ~new_n17691_ & new_n34148_;
  assign new_n34180_ = ~new_n34178_ & ~new_n34179_;
  assign new_n34181_ = pi0626 & new_n34180_;
  assign new_n34182_ = ~pi0641 & ~new_n34181_;
  assign new_n34183_ = ~new_n34177_ & new_n34182_;
  assign new_n34184_ = ~pi0789 & ~new_n34155_;
  assign new_n34185_ = ~new_n34159_ & ~new_n34169_;
  assign new_n34186_ = pi0789 & ~new_n34185_;
  assign new_n34187_ = ~new_n34184_ & ~new_n34186_;
  assign new_n34188_ = ~pi0626 & ~new_n34187_;
  assign new_n34189_ = pi0626 & new_n34011_;
  assign new_n34190_ = pi0641 & ~new_n34189_;
  assign new_n34191_ = ~new_n34188_ & new_n34190_;
  assign new_n34192_ = ~pi1158 & ~new_n34191_;
  assign new_n34193_ = ~new_n34183_ & new_n34192_;
  assign new_n34194_ = pi0626 & new_n34175_;
  assign new_n34195_ = ~pi0626 & new_n34180_;
  assign new_n34196_ = pi0641 & ~new_n34195_;
  assign new_n34197_ = ~new_n34194_ & new_n34196_;
  assign new_n34198_ = pi0626 & ~new_n34187_;
  assign new_n34199_ = ~pi0626 & new_n34011_;
  assign new_n34200_ = ~pi0641 & ~new_n34199_;
  assign new_n34201_ = ~new_n34198_ & new_n34200_;
  assign new_n34202_ = pi1158 & ~new_n34201_;
  assign new_n34203_ = ~new_n34197_ & new_n34202_;
  assign new_n34204_ = ~new_n34193_ & ~new_n34203_;
  assign new_n34205_ = pi0788 & ~new_n34204_;
  assign new_n34206_ = ~new_n34176_ & ~new_n34205_;
  assign new_n34207_ = ~pi0628 & new_n34206_;
  assign new_n34208_ = ~new_n17968_ & ~new_n34187_;
  assign new_n34209_ = new_n17968_ & new_n34011_;
  assign new_n34210_ = ~new_n34208_ & ~new_n34209_;
  assign new_n34211_ = pi0628 & new_n34210_;
  assign new_n34212_ = ~pi1156 & ~new_n34211_;
  assign new_n34213_ = ~new_n34207_ & new_n34212_;
  assign new_n34214_ = ~new_n17734_ & new_n34180_;
  assign new_n34215_ = new_n17734_ & new_n34011_;
  assign new_n34216_ = ~new_n34214_ & ~new_n34215_;
  assign new_n34217_ = pi0628 & new_n34216_;
  assign new_n34218_ = ~pi0628 & ~new_n34011_;
  assign new_n34219_ = pi1156 & ~new_n34218_;
  assign new_n34220_ = ~new_n34217_ & new_n34219_;
  assign new_n34221_ = ~pi0629 & ~new_n34220_;
  assign new_n34222_ = ~new_n34213_ & new_n34221_;
  assign new_n34223_ = pi0628 & new_n34206_;
  assign new_n34224_ = ~pi0628 & new_n34210_;
  assign new_n34225_ = pi1156 & ~new_n34224_;
  assign new_n34226_ = ~new_n34223_ & new_n34225_;
  assign new_n34227_ = ~pi0628 & new_n34216_;
  assign new_n34228_ = pi0628 & ~new_n34011_;
  assign new_n34229_ = ~pi1156 & ~new_n34228_;
  assign new_n34230_ = ~new_n34227_ & new_n34229_;
  assign new_n34231_ = pi0629 & ~new_n34230_;
  assign new_n34232_ = ~new_n34226_ & new_n34231_;
  assign new_n34233_ = ~new_n34222_ & ~new_n34232_;
  assign new_n34234_ = pi0792 & ~new_n34233_;
  assign new_n34235_ = ~pi0792 & new_n34206_;
  assign new_n34236_ = ~new_n34234_ & ~new_n34235_;
  assign new_n34237_ = ~pi0647 & ~new_n34236_;
  assign new_n34238_ = ~new_n17762_ & ~new_n34210_;
  assign new_n34239_ = new_n17762_ & new_n34011_;
  assign new_n34240_ = ~new_n34238_ & ~new_n34239_;
  assign new_n34241_ = pi0647 & new_n34240_;
  assign new_n34242_ = ~pi1157 & ~new_n34241_;
  assign new_n34243_ = ~new_n34237_ & new_n34242_;
  assign new_n34244_ = ~pi0792 & ~new_n34216_;
  assign new_n34245_ = ~new_n34220_ & ~new_n34230_;
  assign new_n34246_ = pi0792 & ~new_n34245_;
  assign new_n34247_ = ~new_n34244_ & ~new_n34246_;
  assign new_n34248_ = pi0647 & new_n34247_;
  assign new_n34249_ = ~pi0647 & ~new_n34011_;
  assign new_n34250_ = pi1157 & ~new_n34249_;
  assign new_n34251_ = ~new_n34248_ & new_n34250_;
  assign new_n34252_ = ~pi0630 & ~new_n34251_;
  assign new_n34253_ = ~new_n34243_ & new_n34252_;
  assign new_n34254_ = pi0647 & ~new_n34236_;
  assign new_n34255_ = ~pi0647 & new_n34240_;
  assign new_n34256_ = pi1157 & ~new_n34255_;
  assign new_n34257_ = ~new_n34254_ & new_n34256_;
  assign new_n34258_ = ~pi0647 & new_n34247_;
  assign new_n34259_ = pi0647 & ~new_n34011_;
  assign new_n34260_ = ~pi1157 & ~new_n34259_;
  assign new_n34261_ = ~new_n34258_ & new_n34260_;
  assign new_n34262_ = pi0630 & ~new_n34261_;
  assign new_n34263_ = ~new_n34257_ & new_n34262_;
  assign new_n34264_ = ~new_n34253_ & ~new_n34263_;
  assign new_n34265_ = pi0787 & ~new_n34264_;
  assign new_n34266_ = ~pi0787 & ~new_n34236_;
  assign new_n34267_ = ~new_n34265_ & ~new_n34266_;
  assign new_n34268_ = ~pi0790 & new_n34267_;
  assign new_n34269_ = ~pi0644 & ~new_n34267_;
  assign new_n34270_ = ~pi0787 & ~new_n34247_;
  assign new_n34271_ = ~new_n34251_ & ~new_n34261_;
  assign new_n34272_ = pi0787 & ~new_n34271_;
  assign new_n34273_ = ~new_n34270_ & ~new_n34272_;
  assign new_n34274_ = pi0644 & new_n34273_;
  assign new_n34275_ = ~pi0715 & ~new_n34274_;
  assign new_n34276_ = ~new_n34269_ & new_n34275_;
  assign new_n34277_ = new_n17804_ & ~new_n34011_;
  assign new_n34278_ = ~new_n17804_ & new_n34240_;
  assign new_n34279_ = ~new_n34277_ & ~new_n34278_;
  assign new_n34280_ = ~pi0644 & ~new_n34279_;
  assign new_n34281_ = pi0644 & ~new_n34011_;
  assign new_n34282_ = pi0715 & ~new_n34281_;
  assign new_n34283_ = ~new_n34280_ & new_n34282_;
  assign new_n34284_ = ~pi1160 & ~new_n34283_;
  assign new_n34285_ = ~new_n34276_ & new_n34284_;
  assign new_n34286_ = pi0644 & ~new_n34267_;
  assign new_n34287_ = ~pi0644 & new_n34273_;
  assign new_n34288_ = pi0715 & ~new_n34287_;
  assign new_n34289_ = ~new_n34286_ & new_n34288_;
  assign new_n34290_ = pi0644 & ~new_n34279_;
  assign new_n34291_ = ~pi0644 & ~new_n34011_;
  assign new_n34292_ = ~pi0715 & ~new_n34291_;
  assign new_n34293_ = ~new_n34290_ & new_n34292_;
  assign new_n34294_ = pi1160 & ~new_n34293_;
  assign new_n34295_ = ~new_n34289_ & new_n34294_;
  assign new_n34296_ = pi0790 & ~new_n34295_;
  assign new_n34297_ = ~new_n34285_ & new_n34296_;
  assign new_n34298_ = ~new_n34268_ & ~new_n34297_;
  assign new_n34299_ = ~po1038 & ~new_n34298_;
  assign new_n34300_ = pi0199 & po1038;
  assign po0356 = new_n34299_ | new_n34300_;
  assign new_n34302_ = pi0200 & ~new_n17558_;
  assign new_n34303_ = ~pi0606 & ~new_n34302_;
  assign new_n34304_ = ~pi0200 & ~new_n19369_;
  assign new_n34305_ = new_n19375_ & ~new_n34304_;
  assign new_n34306_ = pi0200 & new_n17393_;
  assign new_n34307_ = ~pi0200 & ~new_n17426_;
  assign new_n34308_ = ~pi0038 & ~new_n34307_;
  assign new_n34309_ = ~new_n34306_ & new_n34308_;
  assign new_n34310_ = ~new_n34305_ & ~new_n34309_;
  assign new_n34311_ = new_n3272_ & ~new_n34310_;
  assign new_n34312_ = pi0200 & ~new_n3272_;
  assign new_n34313_ = pi0606 & ~new_n34312_;
  assign new_n34314_ = ~new_n34311_ & new_n34313_;
  assign new_n34315_ = ~new_n34303_ & ~new_n34314_;
  assign new_n34316_ = ~new_n17590_ & ~new_n34315_;
  assign new_n34317_ = new_n17590_ & ~new_n34302_;
  assign new_n34318_ = ~new_n34316_ & ~new_n34317_;
  assign new_n34319_ = ~pi0785 & new_n34318_;
  assign new_n34320_ = pi0609 & ~new_n34318_;
  assign new_n34321_ = ~pi0609 & ~new_n34302_;
  assign new_n34322_ = pi1155 & ~new_n34321_;
  assign new_n34323_ = ~new_n34320_ & new_n34322_;
  assign new_n34324_ = ~pi0609 & ~new_n34318_;
  assign new_n34325_ = pi0609 & ~new_n34302_;
  assign new_n34326_ = ~pi1155 & ~new_n34325_;
  assign new_n34327_ = ~new_n34324_ & new_n34326_;
  assign new_n34328_ = ~new_n34323_ & ~new_n34327_;
  assign new_n34329_ = pi0785 & ~new_n34328_;
  assign new_n34330_ = ~new_n34319_ & ~new_n34329_;
  assign new_n34331_ = ~pi0781 & ~new_n34330_;
  assign new_n34332_ = pi0618 & new_n34330_;
  assign new_n34333_ = ~pi0618 & ~new_n34302_;
  assign new_n34334_ = pi1154 & ~new_n34333_;
  assign new_n34335_ = ~new_n34332_ & new_n34334_;
  assign new_n34336_ = ~pi0618 & new_n34330_;
  assign new_n34337_ = pi0618 & ~new_n34302_;
  assign new_n34338_ = ~pi1154 & ~new_n34337_;
  assign new_n34339_ = ~new_n34336_ & new_n34338_;
  assign new_n34340_ = ~new_n34335_ & ~new_n34339_;
  assign new_n34341_ = pi0781 & ~new_n34340_;
  assign new_n34342_ = ~new_n34331_ & ~new_n34341_;
  assign new_n34343_ = ~pi0789 & ~new_n34342_;
  assign new_n34344_ = pi0619 & new_n34342_;
  assign new_n34345_ = ~pi0619 & ~new_n34302_;
  assign new_n34346_ = pi1159 & ~new_n34345_;
  assign new_n34347_ = ~new_n34344_ & new_n34346_;
  assign new_n34348_ = ~pi0619 & new_n34342_;
  assign new_n34349_ = pi0619 & ~new_n34302_;
  assign new_n34350_ = ~pi1159 & ~new_n34349_;
  assign new_n34351_ = ~new_n34348_ & new_n34350_;
  assign new_n34352_ = ~new_n34347_ & ~new_n34351_;
  assign new_n34353_ = pi0789 & ~new_n34352_;
  assign new_n34354_ = ~new_n34343_ & ~new_n34353_;
  assign new_n34355_ = ~new_n17968_ & ~new_n34354_;
  assign new_n34356_ = new_n17968_ & new_n34302_;
  assign new_n34357_ = ~new_n34355_ & ~new_n34356_;
  assign new_n34358_ = ~new_n20567_ & ~new_n34357_;
  assign new_n34359_ = new_n17691_ & ~new_n34302_;
  assign new_n34360_ = new_n17618_ & ~new_n34302_;
  assign new_n34361_ = ~pi0643 & ~new_n34302_;
  assign new_n34362_ = ~pi0200 & ~new_n17431_;
  assign new_n34363_ = new_n19956_ & ~new_n34362_;
  assign new_n34364_ = pi0200 & new_n17517_;
  assign new_n34365_ = ~pi0200 & new_n17468_;
  assign new_n34366_ = ~pi0299 & ~new_n34365_;
  assign new_n34367_ = ~new_n34364_ & new_n34366_;
  assign new_n34368_ = pi0200 & new_n17531_;
  assign new_n34369_ = ~pi0200 & new_n17481_;
  assign new_n34370_ = pi0299 & ~new_n34369_;
  assign new_n34371_ = ~new_n34368_ & new_n34370_;
  assign new_n34372_ = ~new_n34367_ & ~new_n34371_;
  assign new_n34373_ = pi0039 & ~new_n34372_;
  assign new_n34374_ = pi0200 & new_n17200_;
  assign new_n34375_ = ~pi0200 & ~new_n17233_;
  assign new_n34376_ = ~pi0039 & ~new_n34375_;
  assign new_n34377_ = ~new_n34374_ & new_n34376_;
  assign new_n34378_ = ~new_n34373_ & ~new_n34377_;
  assign new_n34379_ = ~pi0038 & ~new_n34378_;
  assign new_n34380_ = ~new_n34363_ & ~new_n34379_;
  assign new_n34381_ = new_n3272_ & ~new_n34380_;
  assign new_n34382_ = pi0643 & ~new_n34312_;
  assign new_n34383_ = ~new_n34381_ & new_n34382_;
  assign new_n34384_ = ~new_n34361_ & ~new_n34383_;
  assign new_n34385_ = ~pi0778 & new_n34384_;
  assign new_n34386_ = pi0625 & ~new_n34384_;
  assign new_n34387_ = ~pi0625 & ~new_n34302_;
  assign new_n34388_ = pi1153 & ~new_n34387_;
  assign new_n34389_ = ~new_n34386_ & new_n34388_;
  assign new_n34390_ = ~pi0625 & ~new_n34384_;
  assign new_n34391_ = pi0625 & ~new_n34302_;
  assign new_n34392_ = ~pi1153 & ~new_n34391_;
  assign new_n34393_ = ~new_n34390_ & new_n34392_;
  assign new_n34394_ = ~new_n34389_ & ~new_n34393_;
  assign new_n34395_ = pi0778 & ~new_n34394_;
  assign new_n34396_ = ~new_n34385_ & ~new_n34395_;
  assign new_n34397_ = ~new_n17618_ & new_n34396_;
  assign new_n34398_ = ~new_n34360_ & ~new_n34397_;
  assign new_n34399_ = ~new_n17655_ & new_n34398_;
  assign new_n34400_ = new_n17655_ & new_n34302_;
  assign new_n34401_ = ~new_n34399_ & ~new_n34400_;
  assign new_n34402_ = ~new_n17691_ & new_n34401_;
  assign new_n34403_ = ~new_n34359_ & ~new_n34402_;
  assign new_n34404_ = ~new_n17734_ & new_n34403_;
  assign new_n34405_ = new_n17734_ & new_n34302_;
  assign new_n34406_ = ~new_n34404_ & ~new_n34405_;
  assign new_n34407_ = pi0628 & new_n34406_;
  assign new_n34408_ = ~pi0628 & ~new_n34302_;
  assign new_n34409_ = pi1156 & ~new_n34408_;
  assign new_n34410_ = ~new_n34407_ & new_n34409_;
  assign new_n34411_ = ~pi0629 & new_n34410_;
  assign new_n34412_ = ~pi0628 & new_n34406_;
  assign new_n34413_ = pi0628 & ~new_n34302_;
  assign new_n34414_ = ~pi1156 & ~new_n34413_;
  assign new_n34415_ = ~new_n34412_ & new_n34414_;
  assign new_n34416_ = pi0629 & new_n34415_;
  assign new_n34417_ = ~new_n34411_ & ~new_n34416_;
  assign new_n34418_ = ~new_n34358_ & new_n34417_;
  assign new_n34419_ = pi0792 & ~new_n34418_;
  assign new_n34420_ = ~pi0643 & new_n34315_;
  assign new_n34421_ = ~new_n16790_ & ~new_n17544_;
  assign new_n34422_ = new_n34363_ & ~new_n34421_;
  assign new_n34423_ = pi0200 & ~new_n19387_;
  assign new_n34424_ = ~pi0200 & ~new_n19393_;
  assign new_n34425_ = ~pi0038 & ~new_n34424_;
  assign new_n34426_ = ~new_n34423_ & new_n34425_;
  assign new_n34427_ = ~new_n34422_ & ~new_n34426_;
  assign new_n34428_ = ~pi0606 & new_n3272_;
  assign new_n34429_ = ~new_n34427_ & new_n34428_;
  assign new_n34430_ = pi0200 & ~new_n24657_;
  assign new_n34431_ = ~pi0200 & ~new_n19403_;
  assign new_n34432_ = ~pi0038 & ~new_n34431_;
  assign new_n34433_ = ~new_n34430_ & new_n34432_;
  assign new_n34434_ = ~new_n19401_ & ~new_n19402_;
  assign new_n34435_ = ~pi0200 & ~new_n34434_;
  assign new_n34436_ = pi0038 & pi0200;
  assign new_n34437_ = new_n19411_ & new_n34436_;
  assign new_n34438_ = pi0606 & new_n3272_;
  assign new_n34439_ = ~new_n34437_ & new_n34438_;
  assign new_n34440_ = ~new_n34435_ & new_n34439_;
  assign new_n34441_ = ~new_n34433_ & new_n34440_;
  assign new_n34442_ = ~new_n34312_ & ~new_n34441_;
  assign new_n34443_ = ~new_n34429_ & new_n34442_;
  assign new_n34444_ = pi0643 & ~new_n34443_;
  assign new_n34445_ = ~new_n34420_ & ~new_n34444_;
  assign new_n34446_ = ~pi0625 & new_n34445_;
  assign new_n34447_ = pi0625 & ~new_n34315_;
  assign new_n34448_ = ~pi1153 & ~new_n34447_;
  assign new_n34449_ = ~new_n34446_ & new_n34448_;
  assign new_n34450_ = ~pi0608 & ~new_n34389_;
  assign new_n34451_ = ~new_n34449_ & new_n34450_;
  assign new_n34452_ = pi0625 & new_n34445_;
  assign new_n34453_ = ~pi0625 & ~new_n34315_;
  assign new_n34454_ = pi1153 & ~new_n34453_;
  assign new_n34455_ = ~new_n34452_ & new_n34454_;
  assign new_n34456_ = pi0608 & ~new_n34393_;
  assign new_n34457_ = ~new_n34455_ & new_n34456_;
  assign new_n34458_ = ~new_n34451_ & ~new_n34457_;
  assign new_n34459_ = pi0778 & ~new_n34458_;
  assign new_n34460_ = ~pi0778 & new_n34445_;
  assign new_n34461_ = ~new_n34459_ & ~new_n34460_;
  assign new_n34462_ = ~pi0609 & ~new_n34461_;
  assign new_n34463_ = pi0609 & new_n34396_;
  assign new_n34464_ = ~pi1155 & ~new_n34463_;
  assign new_n34465_ = ~new_n34462_ & new_n34464_;
  assign new_n34466_ = ~pi0660 & ~new_n34323_;
  assign new_n34467_ = ~new_n34465_ & new_n34466_;
  assign new_n34468_ = pi0609 & ~new_n34461_;
  assign new_n34469_ = ~pi0609 & new_n34396_;
  assign new_n34470_ = pi1155 & ~new_n34469_;
  assign new_n34471_ = ~new_n34468_ & new_n34470_;
  assign new_n34472_ = pi0660 & ~new_n34327_;
  assign new_n34473_ = ~new_n34471_ & new_n34472_;
  assign new_n34474_ = ~new_n34467_ & ~new_n34473_;
  assign new_n34475_ = pi0785 & ~new_n34474_;
  assign new_n34476_ = ~pi0785 & ~new_n34461_;
  assign new_n34477_ = ~new_n34475_ & ~new_n34476_;
  assign new_n34478_ = ~pi0618 & ~new_n34477_;
  assign new_n34479_ = pi0618 & ~new_n34398_;
  assign new_n34480_ = ~pi1154 & ~new_n34479_;
  assign new_n34481_ = ~new_n34478_ & new_n34480_;
  assign new_n34482_ = ~pi0627 & ~new_n34335_;
  assign new_n34483_ = ~new_n34481_ & new_n34482_;
  assign new_n34484_ = pi0618 & ~new_n34477_;
  assign new_n34485_ = ~pi0618 & ~new_n34398_;
  assign new_n34486_ = pi1154 & ~new_n34485_;
  assign new_n34487_ = ~new_n34484_ & new_n34486_;
  assign new_n34488_ = pi0627 & ~new_n34339_;
  assign new_n34489_ = ~new_n34487_ & new_n34488_;
  assign new_n34490_ = ~new_n34483_ & ~new_n34489_;
  assign new_n34491_ = pi0781 & ~new_n34490_;
  assign new_n34492_ = ~pi0781 & ~new_n34477_;
  assign new_n34493_ = ~new_n34491_ & ~new_n34492_;
  assign new_n34494_ = pi0619 & ~new_n34493_;
  assign new_n34495_ = ~pi0619 & new_n34401_;
  assign new_n34496_ = pi1159 & ~new_n34495_;
  assign new_n34497_ = ~new_n34494_ & new_n34496_;
  assign new_n34498_ = pi0648 & ~new_n34351_;
  assign new_n34499_ = ~new_n34497_ & new_n34498_;
  assign new_n34500_ = ~pi0619 & ~new_n34493_;
  assign new_n34501_ = pi0619 & new_n34401_;
  assign new_n34502_ = ~pi1159 & ~new_n34501_;
  assign new_n34503_ = ~new_n34500_ & new_n34502_;
  assign new_n34504_ = ~pi0648 & ~new_n34347_;
  assign new_n34505_ = ~new_n34503_ & new_n34504_;
  assign new_n34506_ = pi0789 & ~new_n34505_;
  assign new_n34507_ = ~new_n34499_ & new_n34506_;
  assign new_n34508_ = ~pi0789 & new_n34493_;
  assign new_n34509_ = new_n17969_ & ~new_n34508_;
  assign new_n34510_ = ~new_n34507_ & new_n34509_;
  assign new_n34511_ = pi0626 & ~new_n34354_;
  assign new_n34512_ = ~pi0626 & new_n34302_;
  assign new_n34513_ = new_n17731_ & ~new_n34512_;
  assign new_n34514_ = ~new_n34511_ & new_n34513_;
  assign new_n34515_ = new_n17856_ & ~new_n34403_;
  assign new_n34516_ = ~pi0626 & ~new_n34354_;
  assign new_n34517_ = pi0626 & new_n34302_;
  assign new_n34518_ = new_n17732_ & ~new_n34517_;
  assign new_n34519_ = ~new_n34516_ & new_n34518_;
  assign new_n34520_ = ~new_n34515_ & ~new_n34519_;
  assign new_n34521_ = ~new_n34514_ & new_n34520_;
  assign new_n34522_ = pi0788 & ~new_n34521_;
  assign new_n34523_ = ~new_n20364_ & ~new_n34522_;
  assign new_n34524_ = ~new_n34510_ & new_n34523_;
  assign new_n34525_ = ~new_n34419_ & ~new_n34524_;
  assign new_n34526_ = ~new_n20360_ & ~new_n34525_;
  assign new_n34527_ = ~pi0792 & ~new_n34406_;
  assign new_n34528_ = ~new_n34410_ & ~new_n34415_;
  assign new_n34529_ = pi0792 & ~new_n34528_;
  assign new_n34530_ = ~new_n34527_ & ~new_n34529_;
  assign new_n34531_ = pi0647 & ~new_n34530_;
  assign new_n34532_ = ~pi0647 & new_n34302_;
  assign new_n34533_ = ~new_n34531_ & ~new_n34532_;
  assign new_n34534_ = new_n17801_ & ~new_n34533_;
  assign new_n34535_ = ~pi0647 & new_n34530_;
  assign new_n34536_ = pi0647 & ~new_n34302_;
  assign new_n34537_ = ~pi1157 & ~new_n34536_;
  assign new_n34538_ = ~new_n34535_ & new_n34537_;
  assign new_n34539_ = pi0630 & new_n34538_;
  assign new_n34540_ = ~new_n17762_ & ~new_n34357_;
  assign new_n34541_ = new_n17762_ & new_n34302_;
  assign new_n34542_ = ~new_n34540_ & ~new_n34541_;
  assign new_n34543_ = ~new_n20556_ & ~new_n34542_;
  assign new_n34544_ = ~new_n34539_ & ~new_n34543_;
  assign new_n34545_ = ~new_n34534_ & new_n34544_;
  assign new_n34546_ = pi0787 & ~new_n34545_;
  assign new_n34547_ = ~new_n34526_ & ~new_n34546_;
  assign new_n34548_ = ~pi0644 & new_n34547_;
  assign new_n34549_ = ~pi0787 & ~new_n34530_;
  assign new_n34550_ = pi1157 & ~new_n34533_;
  assign new_n34551_ = ~new_n34538_ & ~new_n34550_;
  assign new_n34552_ = pi0787 & ~new_n34551_;
  assign new_n34553_ = ~new_n34549_ & ~new_n34552_;
  assign new_n34554_ = pi0644 & new_n34553_;
  assign new_n34555_ = ~pi0715 & ~new_n34554_;
  assign new_n34556_ = ~new_n34548_ & new_n34555_;
  assign new_n34557_ = ~new_n17804_ & ~new_n34542_;
  assign new_n34558_ = new_n17804_ & new_n34302_;
  assign new_n34559_ = ~new_n34557_ & ~new_n34558_;
  assign new_n34560_ = ~pi0644 & new_n34559_;
  assign new_n34561_ = pi0644 & ~new_n34302_;
  assign new_n34562_ = pi0715 & ~new_n34561_;
  assign new_n34563_ = ~new_n34560_ & new_n34562_;
  assign new_n34564_ = ~pi1160 & ~new_n34563_;
  assign new_n34565_ = ~new_n34556_ & new_n34564_;
  assign new_n34566_ = pi0644 & new_n34547_;
  assign new_n34567_ = ~pi0644 & new_n34553_;
  assign new_n34568_ = pi0715 & ~new_n34567_;
  assign new_n34569_ = ~new_n34566_ & new_n34568_;
  assign new_n34570_ = pi0644 & new_n34559_;
  assign new_n34571_ = ~pi0644 & ~new_n34302_;
  assign new_n34572_ = ~pi0715 & ~new_n34571_;
  assign new_n34573_ = ~new_n34570_ & new_n34572_;
  assign new_n34574_ = pi1160 & ~new_n34573_;
  assign new_n34575_ = ~new_n34569_ & new_n34574_;
  assign new_n34576_ = ~new_n34565_ & ~new_n34575_;
  assign new_n34577_ = pi0790 & ~new_n34576_;
  assign new_n34578_ = ~pi0790 & new_n34547_;
  assign new_n34579_ = ~new_n34577_ & ~new_n34578_;
  assign new_n34580_ = ~po1038 & ~new_n34579_;
  assign new_n34581_ = ~pi0200 & po1038;
  assign po0357 = ~new_n34580_ & ~new_n34581_;
  assign new_n34583_ = pi0233 & pi0237;
  assign new_n34584_ = pi0057 & pi0332;
  assign new_n34585_ = pi0332 & ~new_n3298_;
  assign new_n34586_ = ~pi0059 & ~new_n34585_;
  assign new_n34587_ = pi0074 & pi0332;
  assign new_n34588_ = ~pi0055 & ~new_n34587_;
  assign new_n34589_ = new_n2516_ & new_n11086_;
  assign new_n34590_ = pi0468 & new_n6180_;
  assign new_n34591_ = ~pi0299 & pi0587;
  assign new_n34592_ = ~new_n21089_ & ~new_n34591_;
  assign new_n34593_ = ~pi0468 & ~new_n34592_;
  assign new_n34594_ = ~new_n34590_ & ~new_n34593_;
  assign new_n34595_ = new_n34589_ & ~new_n34594_;
  assign new_n34596_ = ~pi0332 & ~new_n34595_;
  assign new_n34597_ = new_n7390_ & ~new_n34596_;
  assign new_n34598_ = new_n3100_ & new_n6617_;
  assign new_n34599_ = ~pi0332 & ~new_n34598_;
  assign new_n34600_ = new_n15692_ & ~new_n34599_;
  assign new_n34601_ = pi0332 & ~new_n3243_;
  assign new_n34602_ = ~new_n34600_ & ~new_n34601_;
  assign new_n34603_ = ~new_n34597_ & new_n34602_;
  assign new_n34604_ = ~pi0074 & ~new_n34603_;
  assign new_n34605_ = new_n34588_ & ~new_n34604_;
  assign new_n34606_ = new_n3273_ & new_n6573_;
  assign new_n34607_ = new_n3100_ & new_n34606_;
  assign new_n34608_ = ~pi0332 & ~new_n34607_;
  assign new_n34609_ = pi0055 & new_n34608_;
  assign new_n34610_ = new_n3298_ & ~new_n34609_;
  assign new_n34611_ = ~new_n34605_ & new_n34610_;
  assign new_n34612_ = new_n34586_ & ~new_n34611_;
  assign new_n34613_ = new_n6304_ & ~new_n34608_;
  assign new_n34614_ = pi0332 & ~new_n6304_;
  assign new_n34615_ = pi0059 & ~new_n34614_;
  assign new_n34616_ = ~new_n34613_ & new_n34615_;
  assign new_n34617_ = ~pi0057 & ~new_n34616_;
  assign new_n34618_ = ~new_n34612_ & new_n34617_;
  assign new_n34619_ = ~new_n34584_ & ~new_n34618_;
  assign new_n34620_ = ~new_n34583_ & ~new_n34619_;
  assign new_n34621_ = ~pi0332 & ~new_n6180_;
  assign new_n34622_ = ~pi0947 & ~new_n34621_;
  assign new_n34623_ = pi0096 & pi0210;
  assign new_n34624_ = pi0332 & new_n34623_;
  assign new_n34625_ = ~pi0032 & pi0070;
  assign new_n34626_ = ~pi0070 & ~pi0841;
  assign new_n34627_ = pi0032 & new_n34626_;
  assign new_n34628_ = ~new_n34625_ & ~new_n34627_;
  assign new_n34629_ = ~pi0210 & ~new_n34628_;
  assign new_n34630_ = ~pi0032 & ~pi0096;
  assign new_n34631_ = pi0070 & new_n34630_;
  assign new_n34632_ = ~pi0332 & ~new_n34631_;
  assign new_n34633_ = ~new_n34629_ & new_n34632_;
  assign new_n34634_ = ~new_n34624_ & ~new_n34633_;
  assign new_n34635_ = ~new_n6185_ & new_n34634_;
  assign new_n34636_ = new_n6180_ & ~new_n34635_;
  assign new_n34637_ = new_n34622_ & ~new_n34636_;
  assign new_n34638_ = pi0332 & pi0468;
  assign new_n34639_ = ~pi0468 & ~new_n34633_;
  assign new_n34640_ = ~new_n34638_ & ~new_n34639_;
  assign new_n34641_ = ~new_n6180_ & new_n34640_;
  assign new_n34642_ = new_n6180_ & ~new_n34634_;
  assign new_n34643_ = pi0947 & ~new_n34642_;
  assign new_n34644_ = ~new_n34641_ & new_n34643_;
  assign new_n34645_ = ~new_n34637_ & ~new_n34644_;
  assign new_n34646_ = pi0057 & ~new_n34645_;
  assign new_n34647_ = ~new_n3273_ & new_n34645_;
  assign new_n34648_ = ~pi0095 & new_n2719_;
  assign new_n34649_ = ~pi0070 & ~new_n34648_;
  assign new_n34650_ = new_n34630_ & ~new_n34649_;
  assign new_n34651_ = pi0210 & new_n34650_;
  assign new_n34652_ = pi0032 & ~new_n34626_;
  assign new_n34653_ = ~pi0095 & new_n2782_;
  assign new_n34654_ = ~new_n34652_ & new_n34653_;
  assign new_n34655_ = new_n2495_ & new_n34654_;
  assign new_n34656_ = new_n2523_ & new_n34655_;
  assign new_n34657_ = new_n34628_ & ~new_n34656_;
  assign new_n34658_ = ~pi0210 & ~new_n34657_;
  assign new_n34659_ = ~pi0332 & ~new_n34658_;
  assign new_n34660_ = ~new_n34651_ & new_n34659_;
  assign new_n34661_ = ~new_n34624_ & ~new_n34660_;
  assign new_n34662_ = ~new_n6185_ & new_n34661_;
  assign new_n34663_ = new_n6180_ & ~new_n34662_;
  assign new_n34664_ = new_n34622_ & ~new_n34663_;
  assign new_n34665_ = ~pi0468 & ~new_n34660_;
  assign new_n34666_ = ~new_n34638_ & ~new_n34665_;
  assign new_n34667_ = ~new_n6180_ & new_n34666_;
  assign new_n34668_ = new_n6180_ & ~new_n34661_;
  assign new_n34669_ = pi0947 & ~new_n34668_;
  assign new_n34670_ = ~new_n34667_ & new_n34669_;
  assign new_n34671_ = ~new_n34664_ & ~new_n34670_;
  assign new_n34672_ = new_n3273_ & new_n34671_;
  assign new_n34673_ = ~new_n34647_ & ~new_n34672_;
  assign new_n34674_ = new_n6304_ & ~new_n34673_;
  assign new_n34675_ = ~new_n6304_ & new_n34645_;
  assign new_n34676_ = pi0059 & ~new_n34675_;
  assign new_n34677_ = ~new_n34674_ & new_n34676_;
  assign new_n34678_ = new_n2516_ & new_n2535_;
  assign new_n34679_ = ~pi0095 & new_n2450_;
  assign new_n34680_ = new_n34678_ & new_n34679_;
  assign new_n34681_ = ~pi0070 & ~new_n34680_;
  assign new_n34682_ = new_n34630_ & ~new_n34681_;
  assign new_n34683_ = pi0210 & new_n34682_;
  assign new_n34684_ = new_n34654_ & new_n34678_;
  assign new_n34685_ = new_n34628_ & ~new_n34684_;
  assign new_n34686_ = ~pi0210 & ~new_n34685_;
  assign new_n34687_ = ~pi0332 & ~new_n34686_;
  assign new_n34688_ = ~new_n34683_ & new_n34687_;
  assign new_n34689_ = ~pi0468 & ~new_n34688_;
  assign new_n34690_ = ~new_n34638_ & ~new_n34689_;
  assign new_n34691_ = ~new_n6180_ & new_n34690_;
  assign new_n34692_ = ~new_n34624_ & ~new_n34688_;
  assign new_n34693_ = new_n6180_ & ~new_n34692_;
  assign new_n34694_ = pi0947 & ~new_n34693_;
  assign new_n34695_ = ~new_n34691_ & new_n34694_;
  assign new_n34696_ = ~new_n6185_ & new_n34692_;
  assign new_n34697_ = new_n6180_ & ~new_n34696_;
  assign new_n34698_ = new_n34622_ & ~new_n34697_;
  assign new_n34699_ = pi0299 & ~new_n34698_;
  assign new_n34700_ = ~new_n34695_ & new_n34699_;
  assign new_n34701_ = pi0198 & new_n34682_;
  assign new_n34702_ = ~pi0198 & ~new_n34685_;
  assign new_n34703_ = ~pi0332 & ~new_n34702_;
  assign new_n34704_ = ~new_n34701_ & new_n34703_;
  assign new_n34705_ = ~pi0468 & ~new_n34704_;
  assign new_n34706_ = ~new_n6180_ & ~new_n34638_;
  assign new_n34707_ = ~new_n34705_ & new_n34706_;
  assign new_n34708_ = pi0096 & pi0198;
  assign new_n34709_ = pi0332 & new_n34708_;
  assign new_n34710_ = ~new_n34704_ & ~new_n34709_;
  assign new_n34711_ = new_n6180_ & ~new_n34710_;
  assign new_n34712_ = pi0587 & ~new_n34711_;
  assign new_n34713_ = ~new_n34707_ & new_n34712_;
  assign new_n34714_ = ~pi0587 & ~new_n34621_;
  assign new_n34715_ = ~new_n6185_ & new_n34710_;
  assign new_n34716_ = new_n6180_ & ~new_n34715_;
  assign new_n34717_ = new_n34714_ & ~new_n34716_;
  assign new_n34718_ = ~pi0299 & ~new_n34717_;
  assign new_n34719_ = ~new_n34713_ & new_n34718_;
  assign new_n34720_ = ~new_n34700_ & ~new_n34719_;
  assign new_n34721_ = new_n7390_ & ~new_n34720_;
  assign new_n34722_ = pi0198 & new_n34650_;
  assign new_n34723_ = ~pi0198 & ~new_n34657_;
  assign new_n34724_ = ~pi0332 & ~new_n34723_;
  assign new_n34725_ = ~new_n34722_ & new_n34724_;
  assign new_n34726_ = ~new_n34709_ & ~new_n34725_;
  assign new_n34727_ = ~new_n6185_ & new_n34726_;
  assign new_n34728_ = new_n6180_ & ~new_n34727_;
  assign new_n34729_ = new_n34714_ & ~new_n34728_;
  assign new_n34730_ = ~pi0468 & ~new_n34725_;
  assign new_n34731_ = new_n34706_ & ~new_n34730_;
  assign new_n34732_ = new_n6180_ & ~new_n34726_;
  assign new_n34733_ = pi0587 & ~new_n34732_;
  assign new_n34734_ = ~new_n34731_ & new_n34733_;
  assign new_n34735_ = ~new_n34729_ & ~new_n34734_;
  assign new_n34736_ = ~pi0299 & ~new_n34735_;
  assign new_n34737_ = pi0299 & ~new_n34671_;
  assign new_n34738_ = new_n15692_ & ~new_n34737_;
  assign new_n34739_ = ~new_n34736_ & new_n34738_;
  assign new_n34740_ = ~new_n34721_ & ~new_n34739_;
  assign new_n34741_ = ~pi0074 & ~new_n34740_;
  assign new_n34742_ = pi0299 & ~new_n34645_;
  assign new_n34743_ = ~pi0074 & new_n3243_;
  assign new_n34744_ = ~pi0198 & ~new_n34628_;
  assign new_n34745_ = new_n34632_ & ~new_n34744_;
  assign new_n34746_ = new_n6577_ & ~new_n34745_;
  assign new_n34747_ = new_n34621_ & ~new_n34746_;
  assign new_n34748_ = ~new_n34709_ & ~new_n34745_;
  assign new_n34749_ = new_n6180_ & ~new_n34748_;
  assign new_n34750_ = ~pi0299 & ~new_n6576_;
  assign new_n34751_ = ~new_n34749_ & new_n34750_;
  assign new_n34752_ = ~new_n34747_ & new_n34751_;
  assign new_n34753_ = ~new_n34743_ & ~new_n34752_;
  assign new_n34754_ = ~new_n34742_ & new_n34753_;
  assign new_n34755_ = ~pi0055 & ~new_n34754_;
  assign new_n34756_ = ~new_n34741_ & new_n34755_;
  assign new_n34757_ = pi0055 & new_n34673_;
  assign new_n34758_ = new_n3298_ & ~new_n34757_;
  assign new_n34759_ = ~new_n34756_ & new_n34758_;
  assign new_n34760_ = ~new_n3298_ & new_n34645_;
  assign new_n34761_ = ~pi0059 & ~new_n34760_;
  assign new_n34762_ = ~new_n34759_ & new_n34761_;
  assign new_n34763_ = ~new_n34677_ & ~new_n34762_;
  assign new_n34764_ = ~pi0057 & ~new_n34763_;
  assign new_n34765_ = ~new_n34646_ & ~new_n34764_;
  assign new_n34766_ = new_n34583_ & ~new_n34765_;
  assign new_n34767_ = ~new_n34620_ & ~new_n34766_;
  assign new_n34768_ = ~pi0201 & ~new_n34767_;
  assign new_n34769_ = ~new_n16479_ & ~new_n34623_;
  assign new_n34770_ = ~new_n6573_ & ~new_n16479_;
  assign new_n34771_ = new_n6577_ & new_n34708_;
  assign new_n34772_ = new_n16479_ & ~new_n34771_;
  assign new_n34773_ = ~new_n34770_ & ~new_n34772_;
  assign new_n34774_ = ~new_n34769_ & new_n34773_;
  assign new_n34775_ = new_n34583_ & new_n34774_;
  assign new_n34776_ = pi0201 & ~new_n34775_;
  assign po0358 = ~new_n34768_ & ~new_n34776_;
  assign new_n34778_ = ~pi0233 & pi0237;
  assign new_n34779_ = ~new_n34619_ & ~new_n34778_;
  assign new_n34780_ = ~new_n34765_ & new_n34778_;
  assign new_n34781_ = ~new_n34779_ & ~new_n34780_;
  assign new_n34782_ = ~pi0202 & ~new_n34781_;
  assign new_n34783_ = new_n34774_ & new_n34778_;
  assign new_n34784_ = pi0202 & ~new_n34783_;
  assign po0359 = ~new_n34782_ & ~new_n34784_;
  assign new_n34786_ = ~pi0233 & ~pi0237;
  assign new_n34787_ = ~new_n34619_ & ~new_n34786_;
  assign new_n34788_ = ~new_n34765_ & new_n34786_;
  assign new_n34789_ = ~new_n34787_ & ~new_n34788_;
  assign new_n34790_ = ~pi0203 & ~new_n34789_;
  assign new_n34791_ = new_n34774_ & new_n34786_;
  assign new_n34792_ = pi0203 & ~new_n34791_;
  assign po0360 = ~new_n34790_ & ~new_n34792_;
  assign new_n34794_ = ~pi0468 & pi0602;
  assign new_n34795_ = pi0468 & new_n6183_;
  assign new_n34796_ = ~new_n34794_ & ~new_n34795_;
  assign new_n34797_ = ~pi0299 & ~new_n34796_;
  assign new_n34798_ = ~new_n6492_ & ~new_n34797_;
  assign new_n34799_ = new_n3100_ & ~new_n34798_;
  assign new_n34800_ = ~pi0332 & ~new_n34799_;
  assign new_n34801_ = new_n15692_ & ~new_n34800_;
  assign new_n34802_ = pi0299 & ~pi0907;
  assign new_n34803_ = ~pi0299 & ~pi0602;
  assign new_n34804_ = ~pi0468 & ~new_n34803_;
  assign new_n34805_ = ~new_n34802_ & new_n34804_;
  assign new_n34806_ = ~new_n34795_ & ~new_n34805_;
  assign new_n34807_ = new_n34589_ & ~new_n34806_;
  assign new_n34808_ = ~pi0332 & ~new_n34807_;
  assign new_n34809_ = new_n7390_ & ~new_n34808_;
  assign new_n34810_ = ~new_n34801_ & ~new_n34809_;
  assign new_n34811_ = ~pi0074 & ~new_n34810_;
  assign new_n34812_ = new_n34588_ & ~new_n34601_;
  assign new_n34813_ = ~new_n34811_ & new_n34812_;
  assign new_n34814_ = new_n3273_ & new_n6310_;
  assign new_n34815_ = new_n3100_ & new_n34814_;
  assign new_n34816_ = ~pi0332 & ~new_n34815_;
  assign new_n34817_ = pi0055 & new_n34816_;
  assign new_n34818_ = new_n3298_ & ~new_n34817_;
  assign new_n34819_ = ~new_n34813_ & new_n34818_;
  assign new_n34820_ = new_n34586_ & ~new_n34819_;
  assign new_n34821_ = new_n6304_ & ~new_n34816_;
  assign new_n34822_ = new_n34615_ & ~new_n34821_;
  assign new_n34823_ = ~pi0057 & ~new_n34822_;
  assign new_n34824_ = ~new_n34820_ & new_n34823_;
  assign new_n34825_ = ~new_n34584_ & ~new_n34824_;
  assign new_n34826_ = ~new_n34583_ & ~new_n34825_;
  assign new_n34827_ = ~pi0332 & ~new_n6183_;
  assign new_n34828_ = ~pi0907 & ~new_n34827_;
  assign new_n34829_ = new_n6183_ & ~new_n34635_;
  assign new_n34830_ = new_n34828_ & ~new_n34829_;
  assign new_n34831_ = ~new_n6183_ & new_n34640_;
  assign new_n34832_ = new_n6183_ & ~new_n34634_;
  assign new_n34833_ = pi0907 & ~new_n34832_;
  assign new_n34834_ = ~new_n34831_ & new_n34833_;
  assign new_n34835_ = ~new_n34830_ & ~new_n34834_;
  assign new_n34836_ = pi0057 & ~new_n34835_;
  assign new_n34837_ = ~new_n3273_ & new_n34835_;
  assign new_n34838_ = ~new_n6183_ & new_n34666_;
  assign new_n34839_ = new_n6183_ & ~new_n34661_;
  assign new_n34840_ = pi0907 & ~new_n34839_;
  assign new_n34841_ = ~new_n34838_ & new_n34840_;
  assign new_n34842_ = pi0332 & ~new_n16630_;
  assign new_n34843_ = pi0680 & ~new_n34842_;
  assign new_n34844_ = ~new_n34662_ & new_n34843_;
  assign new_n34845_ = new_n34828_ & ~new_n34844_;
  assign new_n34846_ = ~new_n34841_ & ~new_n34845_;
  assign new_n34847_ = new_n3273_ & new_n34846_;
  assign new_n34848_ = ~new_n34837_ & ~new_n34847_;
  assign new_n34849_ = new_n6304_ & ~new_n34848_;
  assign new_n34850_ = ~new_n6304_ & new_n34835_;
  assign new_n34851_ = pi0059 & ~new_n34850_;
  assign new_n34852_ = ~new_n34849_ & new_n34851_;
  assign new_n34853_ = pi0299 & new_n34846_;
  assign new_n34854_ = new_n6183_ & new_n34708_;
  assign new_n34855_ = pi0332 & ~new_n34854_;
  assign new_n34856_ = ~pi0299 & ~new_n34855_;
  assign new_n34857_ = new_n6318_ & new_n34726_;
  assign new_n34858_ = new_n34856_ & ~new_n34857_;
  assign new_n34859_ = ~new_n34853_ & ~new_n34858_;
  assign new_n34860_ = new_n15692_ & ~new_n34859_;
  assign new_n34861_ = new_n6318_ & new_n34710_;
  assign new_n34862_ = new_n34856_ & ~new_n34861_;
  assign new_n34863_ = ~new_n6183_ & new_n34690_;
  assign new_n34864_ = new_n6183_ & ~new_n34692_;
  assign new_n34865_ = pi0907 & ~new_n34864_;
  assign new_n34866_ = ~new_n34863_ & new_n34865_;
  assign new_n34867_ = new_n6183_ & ~new_n34696_;
  assign new_n34868_ = new_n34828_ & ~new_n34867_;
  assign new_n34869_ = pi0299 & ~new_n34868_;
  assign new_n34870_ = ~new_n34866_ & new_n34869_;
  assign new_n34871_ = ~new_n34862_ & ~new_n34870_;
  assign new_n34872_ = new_n7390_ & ~new_n34871_;
  assign new_n34873_ = ~new_n34860_ & ~new_n34872_;
  assign new_n34874_ = ~pi0074 & ~new_n34873_;
  assign new_n34875_ = pi0299 & ~new_n34835_;
  assign new_n34876_ = new_n34748_ & ~new_n34796_;
  assign new_n34877_ = ~new_n34855_ & ~new_n34876_;
  assign new_n34878_ = ~pi0299 & ~new_n34877_;
  assign new_n34879_ = ~new_n34743_ & ~new_n34878_;
  assign new_n34880_ = ~new_n34875_ & new_n34879_;
  assign new_n34881_ = ~pi0055 & ~new_n34880_;
  assign new_n34882_ = ~new_n34874_ & new_n34881_;
  assign new_n34883_ = pi0055 & new_n34848_;
  assign new_n34884_ = new_n3298_ & ~new_n34883_;
  assign new_n34885_ = ~new_n34882_ & new_n34884_;
  assign new_n34886_ = ~new_n3298_ & new_n34835_;
  assign new_n34887_ = ~pi0059 & ~new_n34886_;
  assign new_n34888_ = ~new_n34885_ & new_n34887_;
  assign new_n34889_ = ~new_n34852_ & ~new_n34888_;
  assign new_n34890_ = ~pi0057 & ~new_n34889_;
  assign new_n34891_ = ~new_n34836_ & ~new_n34890_;
  assign new_n34892_ = new_n34583_ & ~new_n34891_;
  assign new_n34893_ = ~new_n34826_ & ~new_n34892_;
  assign new_n34894_ = ~pi0204 & ~new_n34893_;
  assign new_n34895_ = new_n6318_ & new_n34708_;
  assign new_n34896_ = new_n16479_ & ~new_n34895_;
  assign new_n34897_ = ~new_n6310_ & ~new_n16479_;
  assign new_n34898_ = ~new_n34769_ & ~new_n34897_;
  assign new_n34899_ = ~new_n34896_ & new_n34898_;
  assign new_n34900_ = new_n34583_ & new_n34899_;
  assign new_n34901_ = pi0204 & ~new_n34900_;
  assign po0361 = ~new_n34894_ & ~new_n34901_;
  assign new_n34903_ = ~new_n34778_ & ~new_n34825_;
  assign new_n34904_ = new_n34778_ & ~new_n34891_;
  assign new_n34905_ = ~new_n34903_ & ~new_n34904_;
  assign new_n34906_ = ~pi0205 & ~new_n34905_;
  assign new_n34907_ = new_n34778_ & new_n34899_;
  assign new_n34908_ = pi0205 & ~new_n34907_;
  assign po0362 = ~new_n34906_ & ~new_n34908_;
  assign new_n34910_ = pi0233 & ~pi0237;
  assign new_n34911_ = ~new_n34825_ & ~new_n34910_;
  assign new_n34912_ = ~new_n34891_ & new_n34910_;
  assign new_n34913_ = ~new_n34911_ & ~new_n34912_;
  assign new_n34914_ = ~pi0206 & ~new_n34913_;
  assign new_n34915_ = new_n34899_ & new_n34910_;
  assign new_n34916_ = pi0206 & ~new_n34915_;
  assign po0363 = ~new_n34914_ & ~new_n34916_;
  assign new_n34918_ = ~new_n19188_ & new_n24384_;
  assign new_n34919_ = new_n19281_ & new_n34918_;
  assign new_n34920_ = ~new_n19311_ & new_n34919_;
  assign new_n34921_ = pi0207 & ~new_n34920_;
  assign new_n34922_ = ~new_n17558_ & new_n17691_;
  assign new_n34923_ = new_n3272_ & new_n24387_;
  assign new_n34924_ = ~pi0778 & ~new_n34923_;
  assign new_n34925_ = ~pi0625 & ~new_n17558_;
  assign new_n34926_ = pi0625 & ~new_n34923_;
  assign new_n34927_ = ~new_n34925_ & ~new_n34926_;
  assign new_n34928_ = pi1153 & ~new_n34927_;
  assign new_n34929_ = pi0625 & ~new_n17558_;
  assign new_n34930_ = ~pi0625 & ~new_n34923_;
  assign new_n34931_ = ~new_n34929_ & ~new_n34930_;
  assign new_n34932_ = ~pi1153 & ~new_n34931_;
  assign new_n34933_ = ~new_n34928_ & ~new_n34932_;
  assign new_n34934_ = pi0778 & ~new_n34933_;
  assign new_n34935_ = ~new_n34924_ & ~new_n34934_;
  assign new_n34936_ = ~new_n17618_ & ~new_n34935_;
  assign new_n34937_ = ~new_n17558_ & new_n17618_;
  assign new_n34938_ = ~new_n34936_ & ~new_n34937_;
  assign new_n34939_ = ~new_n17655_ & new_n34938_;
  assign new_n34940_ = new_n17558_ & new_n17655_;
  assign new_n34941_ = ~new_n34939_ & ~new_n34940_;
  assign new_n34942_ = ~new_n17691_ & new_n34941_;
  assign new_n34943_ = ~new_n34922_ & ~new_n34942_;
  assign new_n34944_ = ~new_n17734_ & new_n34943_;
  assign new_n34945_ = new_n17558_ & new_n17734_;
  assign new_n34946_ = ~new_n34944_ & ~new_n34945_;
  assign new_n34947_ = ~new_n19311_ & ~new_n34946_;
  assign new_n34948_ = new_n17558_ & new_n18010_;
  assign new_n34949_ = ~new_n34947_ & ~new_n34948_;
  assign new_n34950_ = ~pi0207 & ~new_n34949_;
  assign new_n34951_ = ~new_n34921_ & ~new_n34950_;
  assign new_n34952_ = pi0710 & ~new_n34951_;
  assign new_n34953_ = ~pi0207 & ~new_n17558_;
  assign new_n34954_ = ~pi0710 & ~new_n34953_;
  assign new_n34955_ = ~new_n34952_ & ~new_n34954_;
  assign new_n34956_ = ~pi0647 & new_n34955_;
  assign new_n34957_ = pi0647 & new_n34953_;
  assign new_n34958_ = ~pi1157 & ~new_n34957_;
  assign new_n34959_ = ~new_n34956_ & new_n34958_;
  assign new_n34960_ = pi0630 & new_n34959_;
  assign new_n34961_ = pi0647 & new_n34955_;
  assign new_n34962_ = ~pi0647 & new_n34953_;
  assign new_n34963_ = pi1157 & ~new_n34962_;
  assign new_n34964_ = ~new_n34961_ & new_n34963_;
  assign new_n34965_ = ~pi0630 & new_n34964_;
  assign new_n34966_ = ~new_n17558_ & new_n17590_;
  assign new_n34967_ = new_n3272_ & new_n19376_;
  assign new_n34968_ = ~new_n17590_ & ~new_n34967_;
  assign new_n34969_ = ~new_n34966_ & ~new_n34968_;
  assign new_n34970_ = ~pi0785 & ~new_n34969_;
  assign new_n34971_ = ~new_n17558_ & ~new_n17603_;
  assign new_n34972_ = ~pi0609 & new_n34968_;
  assign new_n34973_ = ~new_n34971_ & ~new_n34972_;
  assign new_n34974_ = ~pi1155 & ~new_n34973_;
  assign new_n34975_ = ~new_n17558_ & ~new_n17591_;
  assign new_n34976_ = pi0609 & new_n34968_;
  assign new_n34977_ = ~new_n34975_ & ~new_n34976_;
  assign new_n34978_ = pi1155 & ~new_n34977_;
  assign new_n34979_ = ~new_n34974_ & ~new_n34978_;
  assign new_n34980_ = pi0785 & ~new_n34979_;
  assign new_n34981_ = ~new_n34970_ & ~new_n34980_;
  assign new_n34982_ = ~pi0781 & ~new_n34981_;
  assign new_n34983_ = ~pi0618 & new_n34981_;
  assign new_n34984_ = pi0618 & new_n17558_;
  assign new_n34985_ = ~pi1154 & ~new_n34984_;
  assign new_n34986_ = ~new_n34983_ & new_n34985_;
  assign new_n34987_ = pi0618 & new_n34981_;
  assign new_n34988_ = ~pi0618 & new_n17558_;
  assign new_n34989_ = pi1154 & ~new_n34988_;
  assign new_n34990_ = ~new_n34987_ & new_n34989_;
  assign new_n34991_ = ~new_n34986_ & ~new_n34990_;
  assign new_n34992_ = pi0781 & ~new_n34991_;
  assign new_n34993_ = ~new_n34982_ & ~new_n34992_;
  assign new_n34994_ = ~pi0789 & ~new_n34993_;
  assign new_n34995_ = ~pi0619 & new_n34993_;
  assign new_n34996_ = pi0619 & new_n17558_;
  assign new_n34997_ = ~pi1159 & ~new_n34996_;
  assign new_n34998_ = ~new_n34995_ & new_n34997_;
  assign new_n34999_ = pi0619 & new_n34993_;
  assign new_n35000_ = ~pi0619 & new_n17558_;
  assign new_n35001_ = pi1159 & ~new_n35000_;
  assign new_n35002_ = ~new_n34999_ & new_n35001_;
  assign new_n35003_ = ~new_n34998_ & ~new_n35002_;
  assign new_n35004_ = pi0789 & ~new_n35003_;
  assign new_n35005_ = ~new_n34994_ & ~new_n35004_;
  assign new_n35006_ = ~new_n17968_ & new_n35005_;
  assign new_n35007_ = new_n17558_ & new_n17968_;
  assign new_n35008_ = ~new_n35006_ & ~new_n35007_;
  assign new_n35009_ = ~new_n17762_ & ~new_n35008_;
  assign new_n35010_ = new_n17558_ & new_n17762_;
  assign new_n35011_ = ~new_n35009_ & ~new_n35010_;
  assign new_n35012_ = ~pi0207 & ~new_n35011_;
  assign new_n35013_ = new_n3272_ & ~new_n24446_;
  assign new_n35014_ = ~new_n17590_ & new_n35013_;
  assign new_n35015_ = ~new_n20223_ & new_n35014_;
  assign new_n35016_ = ~new_n20229_ & new_n35015_;
  assign new_n35017_ = ~new_n20233_ & new_n35016_;
  assign new_n35018_ = ~new_n17968_ & new_n35017_;
  assign new_n35019_ = ~new_n17762_ & new_n35018_;
  assign new_n35020_ = pi0207 & ~new_n35019_;
  assign new_n35021_ = pi0623 & ~new_n35020_;
  assign new_n35022_ = ~new_n35012_ & new_n35021_;
  assign new_n35023_ = ~pi0623 & new_n34953_;
  assign new_n35024_ = ~new_n35022_ & ~new_n35023_;
  assign new_n35025_ = ~new_n20556_ & new_n35024_;
  assign new_n35026_ = ~new_n34965_ & ~new_n35025_;
  assign new_n35027_ = ~new_n34960_ & new_n35026_;
  assign new_n35028_ = pi0787 & ~new_n35027_;
  assign new_n35029_ = ~pi0628 & ~new_n17558_;
  assign new_n35030_ = pi0628 & new_n34946_;
  assign new_n35031_ = ~new_n35029_ & ~new_n35030_;
  assign new_n35032_ = ~pi0629 & ~new_n35031_;
  assign new_n35033_ = ~new_n35029_ & ~new_n35032_;
  assign new_n35034_ = pi1156 & ~new_n35033_;
  assign new_n35035_ = pi0628 & ~new_n17558_;
  assign new_n35036_ = ~pi1156 & new_n35035_;
  assign new_n35037_ = ~pi0628 & new_n34946_;
  assign new_n35038_ = ~new_n35035_ & ~new_n35037_;
  assign new_n35039_ = new_n17760_ & ~new_n35038_;
  assign new_n35040_ = ~new_n35036_ & ~new_n35039_;
  assign new_n35041_ = ~new_n35034_ & new_n35040_;
  assign new_n35042_ = pi0792 & ~new_n35041_;
  assign new_n35043_ = pi0619 & new_n34941_;
  assign new_n35044_ = pi0618 & ~new_n34938_;
  assign new_n35045_ = pi0609 & ~new_n34935_;
  assign new_n35046_ = new_n3272_ & ~new_n19389_;
  assign new_n35047_ = ~pi0778 & ~new_n35046_;
  assign new_n35048_ = pi0625 & ~new_n35046_;
  assign new_n35049_ = ~new_n34925_ & ~new_n35048_;
  assign new_n35050_ = pi1153 & ~new_n35049_;
  assign new_n35051_ = pi0608 & ~new_n34932_;
  assign new_n35052_ = ~new_n35050_ & new_n35051_;
  assign new_n35053_ = ~pi0625 & ~new_n35046_;
  assign new_n35054_ = ~new_n34929_ & ~new_n35053_;
  assign new_n35055_ = ~pi1153 & ~new_n35054_;
  assign new_n35056_ = ~pi0608 & ~new_n34928_;
  assign new_n35057_ = ~new_n35055_ & new_n35056_;
  assign new_n35058_ = pi0778 & ~new_n35057_;
  assign new_n35059_ = ~new_n35052_ & new_n35058_;
  assign new_n35060_ = ~new_n35047_ & ~new_n35059_;
  assign new_n35061_ = ~pi0609 & ~new_n35060_;
  assign new_n35062_ = ~new_n35045_ & ~new_n35061_;
  assign new_n35063_ = ~pi1155 & ~new_n35062_;
  assign new_n35064_ = pi1155 & ~new_n17558_;
  assign new_n35065_ = ~pi0660 & ~new_n35064_;
  assign new_n35066_ = ~new_n35063_ & new_n35065_;
  assign new_n35067_ = ~pi0609 & ~new_n34935_;
  assign new_n35068_ = pi0609 & ~new_n35060_;
  assign new_n35069_ = ~new_n35067_ & ~new_n35068_;
  assign new_n35070_ = pi1155 & ~new_n35069_;
  assign new_n35071_ = ~pi1155 & ~new_n17558_;
  assign new_n35072_ = pi0660 & ~new_n35071_;
  assign new_n35073_ = ~new_n35070_ & new_n35072_;
  assign new_n35074_ = ~new_n35066_ & ~new_n35073_;
  assign new_n35075_ = pi0785 & ~new_n35074_;
  assign new_n35076_ = ~pi0785 & new_n35060_;
  assign new_n35077_ = ~new_n35075_ & ~new_n35076_;
  assign new_n35078_ = ~pi0618 & new_n35077_;
  assign new_n35079_ = ~new_n35044_ & ~new_n35078_;
  assign new_n35080_ = ~pi1154 & ~new_n35079_;
  assign new_n35081_ = pi1154 & ~new_n17558_;
  assign new_n35082_ = ~pi0627 & ~new_n35081_;
  assign new_n35083_ = ~new_n35080_ & new_n35082_;
  assign new_n35084_ = ~pi0618 & ~new_n34938_;
  assign new_n35085_ = pi0618 & new_n35077_;
  assign new_n35086_ = ~new_n35084_ & ~new_n35085_;
  assign new_n35087_ = pi1154 & ~new_n35086_;
  assign new_n35088_ = ~pi1154 & ~new_n17558_;
  assign new_n35089_ = pi0627 & ~new_n35088_;
  assign new_n35090_ = ~new_n35087_ & new_n35089_;
  assign new_n35091_ = ~new_n35083_ & ~new_n35090_;
  assign new_n35092_ = pi0781 & ~new_n35091_;
  assign new_n35093_ = ~pi0781 & ~new_n35077_;
  assign new_n35094_ = ~new_n35092_ & ~new_n35093_;
  assign new_n35095_ = ~pi0619 & new_n35094_;
  assign new_n35096_ = ~new_n35043_ & ~new_n35095_;
  assign new_n35097_ = ~pi1159 & ~new_n35096_;
  assign new_n35098_ = pi1159 & ~new_n17558_;
  assign new_n35099_ = ~pi0648 & ~new_n35098_;
  assign new_n35100_ = ~new_n35097_ & new_n35099_;
  assign new_n35101_ = ~pi0619 & new_n34941_;
  assign new_n35102_ = pi0619 & new_n35094_;
  assign new_n35103_ = ~new_n35101_ & ~new_n35102_;
  assign new_n35104_ = pi1159 & ~new_n35103_;
  assign new_n35105_ = ~pi1159 & ~new_n17558_;
  assign new_n35106_ = pi0648 & ~new_n35105_;
  assign new_n35107_ = ~new_n35104_ & new_n35106_;
  assign new_n35108_ = ~new_n35100_ & ~new_n35107_;
  assign new_n35109_ = pi0789 & ~new_n35108_;
  assign new_n35110_ = ~pi0789 & ~new_n35094_;
  assign new_n35111_ = ~new_n35109_ & ~new_n35110_;
  assign new_n35112_ = ~pi0626 & ~new_n35111_;
  assign new_n35113_ = pi0626 & new_n34943_;
  assign new_n35114_ = ~pi0641 & ~new_n35113_;
  assign new_n35115_ = ~new_n35112_ & new_n35114_;
  assign new_n35116_ = pi0641 & ~new_n17558_;
  assign new_n35117_ = ~pi1158 & ~new_n35116_;
  assign new_n35118_ = ~new_n35115_ & new_n35117_;
  assign new_n35119_ = pi0626 & ~new_n35111_;
  assign new_n35120_ = ~pi0626 & new_n34943_;
  assign new_n35121_ = pi0641 & ~new_n35120_;
  assign new_n35122_ = ~new_n35119_ & new_n35121_;
  assign new_n35123_ = ~pi0641 & ~new_n17558_;
  assign new_n35124_ = pi1158 & ~new_n35123_;
  assign new_n35125_ = ~new_n35122_ & new_n35124_;
  assign new_n35126_ = ~new_n35118_ & ~new_n35125_;
  assign new_n35127_ = pi0788 & ~new_n35126_;
  assign new_n35128_ = ~pi0788 & ~new_n35111_;
  assign new_n35129_ = ~new_n20364_ & ~new_n35128_;
  assign new_n35130_ = ~new_n35127_ & new_n35129_;
  assign new_n35131_ = ~new_n35042_ & ~new_n35130_;
  assign new_n35132_ = ~pi0207 & ~new_n35131_;
  assign new_n35133_ = ~pi0778 & ~new_n34027_;
  assign new_n35134_ = pi0625 & new_n34027_;
  assign new_n35135_ = pi1153 & ~new_n35134_;
  assign new_n35136_ = ~pi0625 & new_n24384_;
  assign new_n35137_ = ~pi1153 & ~new_n35136_;
  assign new_n35138_ = pi0608 & ~new_n35137_;
  assign new_n35139_ = ~new_n35135_ & new_n35138_;
  assign new_n35140_ = ~pi0625 & new_n34027_;
  assign new_n35141_ = ~pi1153 & ~new_n35140_;
  assign new_n35142_ = pi0625 & new_n24384_;
  assign new_n35143_ = pi1153 & ~new_n35142_;
  assign new_n35144_ = ~pi0608 & ~new_n35143_;
  assign new_n35145_ = ~new_n35141_ & new_n35144_;
  assign new_n35146_ = pi0778 & ~new_n35145_;
  assign new_n35147_ = ~new_n35139_ & new_n35146_;
  assign new_n35148_ = ~new_n35133_ & ~new_n35147_;
  assign new_n35149_ = ~pi0609 & ~new_n35148_;
  assign new_n35150_ = pi0609 & ~new_n34918_;
  assign new_n35151_ = new_n17615_ & ~new_n35150_;
  assign new_n35152_ = ~new_n35149_ & new_n35151_;
  assign new_n35153_ = pi0609 & ~new_n35148_;
  assign new_n35154_ = ~pi0609 & ~new_n34918_;
  assign new_n35155_ = new_n17616_ & ~new_n35154_;
  assign new_n35156_ = ~new_n35153_ & new_n35155_;
  assign new_n35157_ = ~new_n35152_ & ~new_n35156_;
  assign new_n35158_ = pi0785 & ~new_n35157_;
  assign new_n35159_ = ~pi0785 & new_n35148_;
  assign new_n35160_ = ~new_n35158_ & ~new_n35159_;
  assign new_n35161_ = pi0618 & new_n35160_;
  assign new_n35162_ = ~new_n17618_ & new_n34918_;
  assign new_n35163_ = ~pi0618 & ~new_n35162_;
  assign new_n35164_ = new_n17653_ & ~new_n35163_;
  assign new_n35165_ = ~new_n35161_ & new_n35164_;
  assign new_n35166_ = ~pi0618 & new_n35160_;
  assign new_n35167_ = pi0618 & ~new_n35162_;
  assign new_n35168_ = new_n17652_ & ~new_n35167_;
  assign new_n35169_ = ~new_n35166_ & new_n35168_;
  assign new_n35170_ = pi0781 & ~new_n35169_;
  assign new_n35171_ = ~new_n35165_ & new_n35170_;
  assign new_n35172_ = ~pi0781 & new_n35160_;
  assign new_n35173_ = ~new_n23615_ & ~new_n35172_;
  assign new_n35174_ = ~new_n35171_ & new_n35173_;
  assign new_n35175_ = new_n19280_ & new_n34918_;
  assign new_n35176_ = new_n17690_ & new_n20233_;
  assign new_n35177_ = new_n35175_ & new_n35176_;
  assign new_n35178_ = ~new_n35174_ & ~new_n35177_;
  assign new_n35179_ = pi0626 & new_n35178_;
  assign new_n35180_ = ~new_n17691_ & new_n35175_;
  assign new_n35181_ = ~pi0626 & ~new_n35180_;
  assign new_n35182_ = pi0641 & ~new_n35181_;
  assign new_n35183_ = pi1158 & new_n35182_;
  assign new_n35184_ = ~new_n35179_ & new_n35183_;
  assign new_n35185_ = ~pi0626 & new_n35178_;
  assign new_n35186_ = pi0626 & ~new_n35180_;
  assign new_n35187_ = ~pi0641 & ~new_n35186_;
  assign new_n35188_ = ~pi1158 & new_n35187_;
  assign new_n35189_ = ~new_n35185_ & new_n35188_;
  assign new_n35190_ = pi0788 & ~new_n35189_;
  assign new_n35191_ = ~new_n35184_ & new_n35190_;
  assign new_n35192_ = ~pi0788 & new_n35178_;
  assign new_n35193_ = ~new_n20364_ & ~new_n35192_;
  assign new_n35194_ = ~new_n35191_ & new_n35193_;
  assign new_n35195_ = new_n17762_ & new_n18009_;
  assign new_n35196_ = new_n34919_ & new_n35195_;
  assign new_n35197_ = ~new_n35194_ & ~new_n35196_;
  assign new_n35198_ = pi0207 & ~new_n35197_;
  assign new_n35199_ = ~pi0623 & ~new_n35198_;
  assign new_n35200_ = ~new_n35132_ & new_n35199_;
  assign new_n35201_ = new_n3272_ & new_n19414_;
  assign new_n35202_ = ~pi0778 & ~new_n35201_;
  assign new_n35203_ = pi0625 & new_n34967_;
  assign new_n35204_ = ~pi0625 & new_n35201_;
  assign new_n35205_ = ~pi1153 & ~new_n35204_;
  assign new_n35206_ = ~new_n35203_ & new_n35205_;
  assign new_n35207_ = new_n35056_ & ~new_n35206_;
  assign new_n35208_ = ~pi0625 & new_n34967_;
  assign new_n35209_ = pi0625 & new_n35201_;
  assign new_n35210_ = pi1153 & ~new_n35209_;
  assign new_n35211_ = ~new_n35208_ & new_n35210_;
  assign new_n35212_ = new_n35051_ & ~new_n35211_;
  assign new_n35213_ = pi0778 & ~new_n35212_;
  assign new_n35214_ = ~new_n35207_ & new_n35213_;
  assign new_n35215_ = ~new_n35202_ & ~new_n35214_;
  assign new_n35216_ = ~pi0609 & ~new_n35215_;
  assign new_n35217_ = ~new_n35045_ & ~new_n35216_;
  assign new_n35218_ = ~pi1155 & ~new_n35217_;
  assign new_n35219_ = ~pi0660 & ~new_n34978_;
  assign new_n35220_ = ~new_n35218_ & new_n35219_;
  assign new_n35221_ = pi0609 & ~new_n35215_;
  assign new_n35222_ = ~new_n35067_ & ~new_n35221_;
  assign new_n35223_ = pi1155 & ~new_n35222_;
  assign new_n35224_ = pi0660 & ~new_n34974_;
  assign new_n35225_ = ~new_n35223_ & new_n35224_;
  assign new_n35226_ = ~new_n35220_ & ~new_n35225_;
  assign new_n35227_ = pi0785 & ~new_n35226_;
  assign new_n35228_ = ~pi0785 & new_n35215_;
  assign new_n35229_ = ~new_n35227_ & ~new_n35228_;
  assign new_n35230_ = ~pi0618 & new_n35229_;
  assign new_n35231_ = ~new_n35044_ & ~new_n35230_;
  assign new_n35232_ = ~pi1154 & ~new_n35231_;
  assign new_n35233_ = ~pi0627 & ~new_n34990_;
  assign new_n35234_ = ~new_n35232_ & new_n35233_;
  assign new_n35235_ = pi0618 & new_n35229_;
  assign new_n35236_ = ~new_n35084_ & ~new_n35235_;
  assign new_n35237_ = pi1154 & ~new_n35236_;
  assign new_n35238_ = pi0627 & ~new_n34986_;
  assign new_n35239_ = ~new_n35237_ & new_n35238_;
  assign new_n35240_ = ~new_n35234_ & ~new_n35239_;
  assign new_n35241_ = pi0781 & ~new_n35240_;
  assign new_n35242_ = ~pi0781 & ~new_n35229_;
  assign new_n35243_ = ~new_n35241_ & ~new_n35242_;
  assign new_n35244_ = pi0619 & new_n35243_;
  assign new_n35245_ = ~new_n35101_ & ~new_n35244_;
  assign new_n35246_ = pi1159 & ~new_n35245_;
  assign new_n35247_ = pi0648 & ~new_n34998_;
  assign new_n35248_ = ~new_n35246_ & new_n35247_;
  assign new_n35249_ = ~pi0619 & new_n35243_;
  assign new_n35250_ = ~new_n35043_ & ~new_n35249_;
  assign new_n35251_ = ~pi1159 & ~new_n35250_;
  assign new_n35252_ = ~pi0648 & ~new_n35002_;
  assign new_n35253_ = ~new_n35251_ & new_n35252_;
  assign new_n35254_ = pi0789 & ~new_n35253_;
  assign new_n35255_ = ~new_n35248_ & new_n35254_;
  assign new_n35256_ = ~pi0789 & new_n35243_;
  assign new_n35257_ = new_n17969_ & ~new_n35256_;
  assign new_n35258_ = ~new_n35255_ & new_n35257_;
  assign new_n35259_ = ~new_n17733_ & ~new_n17855_;
  assign new_n35260_ = new_n35005_ & new_n35259_;
  assign new_n35261_ = pi0641 & ~new_n34943_;
  assign new_n35262_ = new_n17850_ & ~new_n35123_;
  assign new_n35263_ = ~new_n35261_ & new_n35262_;
  assign new_n35264_ = ~pi0641 & ~new_n34943_;
  assign new_n35265_ = new_n17851_ & ~new_n35116_;
  assign new_n35266_ = ~new_n35264_ & new_n35265_;
  assign new_n35267_ = ~new_n35263_ & ~new_n35266_;
  assign new_n35268_ = ~new_n35260_ & new_n35267_;
  assign new_n35269_ = pi0788 & ~new_n35268_;
  assign new_n35270_ = ~new_n20364_ & ~new_n35269_;
  assign new_n35271_ = ~new_n35258_ & new_n35270_;
  assign new_n35272_ = pi1156 & new_n35032_;
  assign new_n35273_ = ~new_n20567_ & new_n35008_;
  assign new_n35274_ = ~new_n35039_ & ~new_n35273_;
  assign new_n35275_ = ~new_n35272_ & new_n35274_;
  assign new_n35276_ = pi0792 & ~new_n35275_;
  assign new_n35277_ = ~new_n35271_ & ~new_n35276_;
  assign new_n35278_ = ~pi0207 & ~new_n35277_;
  assign new_n35279_ = pi1156 & ~new_n35018_;
  assign new_n35280_ = ~pi1156 & ~new_n34919_;
  assign new_n35281_ = new_n20563_ & ~new_n35280_;
  assign new_n35282_ = ~new_n35279_ & new_n35281_;
  assign new_n35283_ = ~pi1156 & ~new_n35018_;
  assign new_n35284_ = pi1156 & ~new_n34919_;
  assign new_n35285_ = new_n20565_ & ~new_n35284_;
  assign new_n35286_ = ~new_n35283_ & new_n35285_;
  assign new_n35287_ = ~new_n35282_ & ~new_n35286_;
  assign new_n35288_ = pi0792 & ~new_n35287_;
  assign new_n35289_ = ~pi1159 & ~new_n35175_;
  assign new_n35290_ = pi1159 & ~new_n35016_;
  assign new_n35291_ = pi0619 & ~pi0648;
  assign new_n35292_ = ~new_n35290_ & new_n35291_;
  assign new_n35293_ = ~new_n35289_ & new_n35292_;
  assign new_n35294_ = pi1159 & ~new_n35175_;
  assign new_n35295_ = ~pi1159 & ~new_n35016_;
  assign new_n35296_ = ~pi0619 & pi0648;
  assign new_n35297_ = ~new_n35295_ & new_n35296_;
  assign new_n35298_ = ~new_n35294_ & new_n35297_;
  assign new_n35299_ = pi0789 & ~new_n35298_;
  assign new_n35300_ = ~new_n35293_ & new_n35299_;
  assign new_n35301_ = pi0789 & ~new_n35300_;
  assign new_n35302_ = ~pi1154 & ~new_n35167_;
  assign new_n35303_ = new_n20226_ & new_n35015_;
  assign new_n35304_ = ~pi0627 & ~new_n35303_;
  assign new_n35305_ = ~new_n35302_ & new_n35304_;
  assign new_n35306_ = ~pi0778 & ~new_n34032_;
  assign new_n35307_ = pi0625 & new_n34032_;
  assign new_n35308_ = ~pi0625 & new_n35013_;
  assign new_n35309_ = pi1153 & ~new_n35308_;
  assign new_n35310_ = ~new_n35307_ & new_n35309_;
  assign new_n35311_ = new_n35138_ & ~new_n35310_;
  assign new_n35312_ = ~pi0625 & new_n34032_;
  assign new_n35313_ = pi0625 & new_n35013_;
  assign new_n35314_ = ~pi1153 & ~new_n35313_;
  assign new_n35315_ = ~new_n35312_ & new_n35314_;
  assign new_n35316_ = new_n35144_ & ~new_n35315_;
  assign new_n35317_ = pi0778 & ~new_n35316_;
  assign new_n35318_ = ~new_n35311_ & new_n35317_;
  assign new_n35319_ = ~new_n35306_ & ~new_n35318_;
  assign new_n35320_ = ~pi0785 & ~new_n35319_;
  assign new_n35321_ = ~pi0609 & ~new_n35319_;
  assign new_n35322_ = ~pi1155 & ~new_n35150_;
  assign new_n35323_ = ~new_n35321_ & new_n35322_;
  assign new_n35324_ = new_n20220_ & new_n35014_;
  assign new_n35325_ = ~pi0660 & ~new_n35324_;
  assign new_n35326_ = ~new_n35323_ & new_n35325_;
  assign new_n35327_ = pi0609 & ~new_n35319_;
  assign new_n35328_ = pi1155 & ~new_n35154_;
  assign new_n35329_ = ~new_n35327_ & new_n35328_;
  assign new_n35330_ = new_n20221_ & new_n35014_;
  assign new_n35331_ = pi0660 & ~new_n35330_;
  assign new_n35332_ = ~new_n35329_ & new_n35331_;
  assign new_n35333_ = ~new_n35326_ & ~new_n35332_;
  assign new_n35334_ = pi0785 & ~new_n35333_;
  assign new_n35335_ = ~new_n35320_ & ~new_n35334_;
  assign new_n35336_ = pi0618 & ~new_n35335_;
  assign new_n35337_ = pi1154 & ~new_n35163_;
  assign new_n35338_ = ~new_n35336_ & new_n35337_;
  assign new_n35339_ = new_n20227_ & new_n35015_;
  assign new_n35340_ = pi0627 & ~new_n35339_;
  assign new_n35341_ = ~new_n35338_ & new_n35340_;
  assign new_n35342_ = ~new_n35305_ & ~new_n35341_;
  assign new_n35343_ = pi0781 & ~new_n35342_;
  assign new_n35344_ = ~pi0618 & ~pi0627;
  assign new_n35345_ = pi0781 & ~new_n35344_;
  assign new_n35346_ = ~new_n35335_ & ~new_n35345_;
  assign new_n35347_ = ~new_n23614_ & new_n35300_;
  assign new_n35348_ = ~new_n35346_ & ~new_n35347_;
  assign new_n35349_ = ~new_n35343_ & new_n35348_;
  assign new_n35350_ = ~new_n35301_ & ~new_n35349_;
  assign new_n35351_ = ~pi0626 & new_n35350_;
  assign new_n35352_ = new_n35187_ & ~new_n35351_;
  assign new_n35353_ = new_n17853_ & new_n35017_;
  assign new_n35354_ = ~pi1158 & ~new_n35353_;
  assign new_n35355_ = ~new_n35352_ & new_n35354_;
  assign new_n35356_ = pi0626 & new_n35350_;
  assign new_n35357_ = new_n35182_ & ~new_n35356_;
  assign new_n35358_ = new_n17854_ & new_n35017_;
  assign new_n35359_ = pi1158 & ~new_n35358_;
  assign new_n35360_ = ~new_n35357_ & new_n35359_;
  assign new_n35361_ = ~new_n35355_ & ~new_n35360_;
  assign new_n35362_ = pi0788 & ~new_n35361_;
  assign new_n35363_ = ~pi0788 & new_n35350_;
  assign new_n35364_ = ~new_n20364_ & ~new_n35363_;
  assign new_n35365_ = ~new_n35362_ & new_n35364_;
  assign new_n35366_ = ~new_n35288_ & ~new_n35365_;
  assign new_n35367_ = pi0207 & ~new_n35366_;
  assign new_n35368_ = pi0623 & ~new_n35367_;
  assign new_n35369_ = ~new_n35278_ & new_n35368_;
  assign new_n35370_ = pi0710 & ~new_n35369_;
  assign new_n35371_ = ~new_n35200_ & new_n35370_;
  assign new_n35372_ = ~pi0710 & ~new_n35024_;
  assign new_n35373_ = ~new_n20360_ & ~new_n35372_;
  assign new_n35374_ = ~new_n35371_ & new_n35373_;
  assign new_n35375_ = ~new_n35028_ & ~new_n35374_;
  assign new_n35376_ = pi0644 & new_n35375_;
  assign new_n35377_ = ~pi0787 & ~new_n34955_;
  assign new_n35378_ = ~new_n34959_ & ~new_n34964_;
  assign new_n35379_ = pi0787 & ~new_n35378_;
  assign new_n35380_ = ~new_n35377_ & ~new_n35379_;
  assign new_n35381_ = ~pi0644 & new_n35380_;
  assign new_n35382_ = pi0715 & ~new_n35381_;
  assign new_n35383_ = ~new_n35376_ & new_n35382_;
  assign new_n35384_ = new_n17804_ & ~new_n34953_;
  assign new_n35385_ = ~new_n17804_ & new_n35024_;
  assign new_n35386_ = ~new_n35384_ & ~new_n35385_;
  assign new_n35387_ = pi0644 & new_n35386_;
  assign new_n35388_ = ~pi0644 & new_n34953_;
  assign new_n35389_ = ~pi0715 & ~new_n35388_;
  assign new_n35390_ = ~new_n35387_ & new_n35389_;
  assign new_n35391_ = pi1160 & ~new_n35390_;
  assign new_n35392_ = ~new_n35383_ & new_n35391_;
  assign new_n35393_ = ~pi0644 & new_n35375_;
  assign new_n35394_ = pi0644 & new_n35380_;
  assign new_n35395_ = ~pi0715 & ~new_n35394_;
  assign new_n35396_ = ~new_n35393_ & new_n35395_;
  assign new_n35397_ = ~pi0644 & new_n35386_;
  assign new_n35398_ = pi0644 & new_n34953_;
  assign new_n35399_ = pi0715 & ~new_n35398_;
  assign new_n35400_ = ~new_n35397_ & new_n35399_;
  assign new_n35401_ = ~pi1160 & ~new_n35400_;
  assign new_n35402_ = ~new_n35396_ & new_n35401_;
  assign new_n35403_ = ~new_n35392_ & ~new_n35402_;
  assign new_n35404_ = pi0790 & ~new_n35403_;
  assign new_n35405_ = ~pi0790 & new_n35375_;
  assign new_n35406_ = ~new_n35404_ & ~new_n35405_;
  assign new_n35407_ = ~po1038 & ~new_n35406_;
  assign new_n35408_ = ~pi0207 & po1038;
  assign po0364 = new_n35407_ | new_n35408_;
  assign new_n35410_ = pi0208 & ~new_n34920_;
  assign new_n35411_ = ~pi0208 & ~new_n34949_;
  assign new_n35412_ = ~new_n35410_ & ~new_n35411_;
  assign new_n35413_ = pi0638 & ~new_n35412_;
  assign new_n35414_ = ~pi0208 & ~new_n17558_;
  assign new_n35415_ = ~pi0638 & ~new_n35414_;
  assign new_n35416_ = ~new_n35413_ & ~new_n35415_;
  assign new_n35417_ = ~pi0647 & new_n35416_;
  assign new_n35418_ = pi0647 & new_n35414_;
  assign new_n35419_ = ~pi1157 & ~new_n35418_;
  assign new_n35420_ = ~new_n35417_ & new_n35419_;
  assign new_n35421_ = pi0630 & new_n35420_;
  assign new_n35422_ = pi0647 & new_n35416_;
  assign new_n35423_ = ~pi0647 & new_n35414_;
  assign new_n35424_ = pi1157 & ~new_n35423_;
  assign new_n35425_ = ~new_n35422_ & new_n35424_;
  assign new_n35426_ = ~pi0630 & new_n35425_;
  assign new_n35427_ = ~pi0208 & ~new_n35011_;
  assign new_n35428_ = pi0208 & ~new_n35019_;
  assign new_n35429_ = pi0607 & ~new_n35428_;
  assign new_n35430_ = ~new_n35427_ & new_n35429_;
  assign new_n35431_ = ~pi0607 & new_n35414_;
  assign new_n35432_ = ~new_n35430_ & ~new_n35431_;
  assign new_n35433_ = ~new_n20556_ & new_n35432_;
  assign new_n35434_ = ~new_n35426_ & ~new_n35433_;
  assign new_n35435_ = ~new_n35421_ & new_n35434_;
  assign new_n35436_ = pi0787 & ~new_n35435_;
  assign new_n35437_ = ~pi0208 & ~new_n35131_;
  assign new_n35438_ = pi0208 & ~new_n35197_;
  assign new_n35439_ = ~pi0607 & ~new_n35438_;
  assign new_n35440_ = ~new_n35437_ & new_n35439_;
  assign new_n35441_ = ~pi0208 & ~new_n35277_;
  assign new_n35442_ = pi0208 & ~new_n35366_;
  assign new_n35443_ = pi0607 & ~new_n35442_;
  assign new_n35444_ = ~new_n35441_ & new_n35443_;
  assign new_n35445_ = pi0638 & ~new_n35444_;
  assign new_n35446_ = ~new_n35440_ & new_n35445_;
  assign new_n35447_ = ~pi0638 & ~new_n35432_;
  assign new_n35448_ = ~new_n20360_ & ~new_n35447_;
  assign new_n35449_ = ~new_n35446_ & new_n35448_;
  assign new_n35450_ = ~new_n35436_ & ~new_n35449_;
  assign new_n35451_ = pi0644 & new_n35450_;
  assign new_n35452_ = ~pi0787 & ~new_n35416_;
  assign new_n35453_ = ~new_n35420_ & ~new_n35425_;
  assign new_n35454_ = pi0787 & ~new_n35453_;
  assign new_n35455_ = ~new_n35452_ & ~new_n35454_;
  assign new_n35456_ = ~pi0644 & new_n35455_;
  assign new_n35457_ = pi0715 & ~new_n35456_;
  assign new_n35458_ = ~new_n35451_ & new_n35457_;
  assign new_n35459_ = new_n17804_ & ~new_n35414_;
  assign new_n35460_ = ~new_n17804_ & new_n35432_;
  assign new_n35461_ = ~new_n35459_ & ~new_n35460_;
  assign new_n35462_ = pi0644 & new_n35461_;
  assign new_n35463_ = ~pi0644 & new_n35414_;
  assign new_n35464_ = ~pi0715 & ~new_n35463_;
  assign new_n35465_ = ~new_n35462_ & new_n35464_;
  assign new_n35466_ = pi1160 & ~new_n35465_;
  assign new_n35467_ = ~new_n35458_ & new_n35466_;
  assign new_n35468_ = ~pi0644 & new_n35450_;
  assign new_n35469_ = pi0644 & new_n35455_;
  assign new_n35470_ = ~pi0715 & ~new_n35469_;
  assign new_n35471_ = ~new_n35468_ & new_n35470_;
  assign new_n35472_ = ~pi0644 & new_n35461_;
  assign new_n35473_ = pi0644 & new_n35414_;
  assign new_n35474_ = pi0715 & ~new_n35473_;
  assign new_n35475_ = ~new_n35472_ & new_n35474_;
  assign new_n35476_ = ~pi1160 & ~new_n35475_;
  assign new_n35477_ = ~new_n35471_ & new_n35476_;
  assign new_n35478_ = ~new_n35467_ & ~new_n35477_;
  assign new_n35479_ = pi0790 & ~new_n35478_;
  assign new_n35480_ = ~pi0790 & new_n35450_;
  assign new_n35481_ = ~new_n35479_ & ~new_n35480_;
  assign new_n35482_ = ~po1038 & ~new_n35481_;
  assign new_n35483_ = ~pi0208 & po1038;
  assign po0365 = new_n35482_ | new_n35483_;
  assign new_n35485_ = ~new_n20360_ & ~new_n35131_;
  assign new_n35486_ = ~pi0647 & ~new_n17558_;
  assign new_n35487_ = pi0647 & new_n34949_;
  assign new_n35488_ = ~new_n35486_ & ~new_n35487_;
  assign new_n35489_ = ~pi0630 & ~new_n35488_;
  assign new_n35490_ = ~new_n35486_ & ~new_n35489_;
  assign new_n35491_ = pi1157 & ~new_n35490_;
  assign new_n35492_ = pi0647 & ~new_n17558_;
  assign new_n35493_ = ~pi1157 & new_n35492_;
  assign new_n35494_ = ~pi0647 & new_n34949_;
  assign new_n35495_ = ~new_n35492_ & ~new_n35494_;
  assign new_n35496_ = new_n17802_ & ~new_n35495_;
  assign new_n35497_ = ~new_n35493_ & ~new_n35496_;
  assign new_n35498_ = ~new_n35491_ & new_n35497_;
  assign new_n35499_ = pi0787 & ~new_n35498_;
  assign new_n35500_ = ~new_n35485_ & ~new_n35499_;
  assign new_n35501_ = ~pi0644 & ~new_n35500_;
  assign new_n35502_ = ~new_n19335_ & new_n34949_;
  assign new_n35503_ = ~new_n17558_ & new_n19335_;
  assign new_n35504_ = ~new_n35502_ & ~new_n35503_;
  assign new_n35505_ = pi0644 & ~new_n35504_;
  assign new_n35506_ = ~pi0715 & ~new_n35505_;
  assign new_n35507_ = ~new_n35501_ & new_n35506_;
  assign new_n35508_ = pi0715 & new_n17558_;
  assign new_n35509_ = ~pi1160 & ~new_n35508_;
  assign new_n35510_ = ~new_n35507_ & new_n35509_;
  assign new_n35511_ = pi0644 & ~new_n35500_;
  assign new_n35512_ = ~pi0644 & ~new_n35504_;
  assign new_n35513_ = pi0715 & ~new_n35512_;
  assign new_n35514_ = ~new_n35511_ & new_n35513_;
  assign new_n35515_ = ~pi0715 & new_n17558_;
  assign new_n35516_ = pi1160 & ~new_n35515_;
  assign new_n35517_ = ~new_n35514_ & new_n35516_;
  assign new_n35518_ = ~new_n35510_ & ~new_n35517_;
  assign new_n35519_ = pi0790 & ~new_n35518_;
  assign new_n35520_ = ~pi0790 & ~new_n35500_;
  assign new_n35521_ = ~po1038 & ~new_n35520_;
  assign new_n35522_ = ~new_n35519_ & new_n35521_;
  assign new_n35523_ = pi0639 & new_n35522_;
  assign new_n35524_ = new_n10197_ & new_n17551_;
  assign new_n35525_ = ~pi0639 & new_n35524_;
  assign new_n35526_ = ~pi0622 & ~new_n35525_;
  assign new_n35527_ = ~new_n35523_ & new_n35526_;
  assign new_n35528_ = ~new_n20360_ & ~new_n35277_;
  assign new_n35529_ = pi1157 & new_n35489_;
  assign new_n35530_ = ~new_n20556_ & new_n35011_;
  assign new_n35531_ = ~new_n35496_ & ~new_n35530_;
  assign new_n35532_ = ~new_n35529_ & new_n35531_;
  assign new_n35533_ = pi0787 & ~new_n35532_;
  assign new_n35534_ = ~new_n35528_ & ~new_n35533_;
  assign new_n35535_ = ~pi0644 & ~new_n35534_;
  assign new_n35536_ = new_n35506_ & ~new_n35535_;
  assign new_n35537_ = ~new_n17558_ & new_n17804_;
  assign new_n35538_ = ~new_n17804_ & new_n35011_;
  assign new_n35539_ = ~new_n35537_ & ~new_n35538_;
  assign new_n35540_ = ~pi0644 & ~new_n35539_;
  assign new_n35541_ = pi0644 & ~new_n17558_;
  assign new_n35542_ = ~new_n35540_ & ~new_n35541_;
  assign new_n35543_ = pi0715 & new_n35542_;
  assign new_n35544_ = ~pi1160 & ~new_n35543_;
  assign new_n35545_ = ~new_n35536_ & new_n35544_;
  assign new_n35546_ = pi0644 & ~new_n35534_;
  assign new_n35547_ = new_n35513_ & ~new_n35546_;
  assign new_n35548_ = pi0644 & ~new_n35539_;
  assign new_n35549_ = ~pi0644 & ~new_n17558_;
  assign new_n35550_ = ~new_n35548_ & ~new_n35549_;
  assign new_n35551_ = ~pi0715 & new_n35550_;
  assign new_n35552_ = pi1160 & ~new_n35551_;
  assign new_n35553_ = ~new_n35547_ & new_n35552_;
  assign new_n35554_ = ~new_n35545_ & ~new_n35553_;
  assign new_n35555_ = pi0790 & ~new_n35554_;
  assign new_n35556_ = ~pi0790 & ~new_n35534_;
  assign new_n35557_ = ~po1038 & ~new_n35556_;
  assign new_n35558_ = ~new_n35555_ & new_n35557_;
  assign new_n35559_ = pi0639 & new_n35558_;
  assign new_n35560_ = ~pi1160 & new_n35542_;
  assign new_n35561_ = pi1160 & new_n35550_;
  assign new_n35562_ = pi0790 & ~new_n35561_;
  assign new_n35563_ = ~new_n35560_ & new_n35562_;
  assign new_n35564_ = ~pi0790 & ~new_n35539_;
  assign new_n35565_ = ~po1038 & ~new_n35564_;
  assign new_n35566_ = ~new_n35563_ & new_n35565_;
  assign new_n35567_ = ~pi0639 & new_n35566_;
  assign new_n35568_ = pi0622 & ~new_n35567_;
  assign new_n35569_ = ~new_n35559_ & new_n35568_;
  assign new_n35570_ = ~new_n35527_ & ~new_n35569_;
  assign new_n35571_ = ~pi0209 & ~new_n35570_;
  assign new_n35572_ = ~new_n19335_ & new_n34920_;
  assign new_n35573_ = pi0644 & ~new_n35572_;
  assign new_n35574_ = ~pi0715 & ~new_n35573_;
  assign new_n35575_ = ~pi0647 & ~new_n35366_;
  assign new_n35576_ = pi0647 & new_n35019_;
  assign new_n35577_ = ~pi1157 & ~new_n35576_;
  assign new_n35578_ = ~new_n35575_ & new_n35577_;
  assign new_n35579_ = pi0647 & new_n34920_;
  assign new_n35580_ = pi1157 & ~new_n35579_;
  assign new_n35581_ = ~pi0630 & ~new_n35580_;
  assign new_n35582_ = ~new_n35578_ & new_n35581_;
  assign new_n35583_ = pi0647 & ~new_n35366_;
  assign new_n35584_ = ~pi0647 & new_n35019_;
  assign new_n35585_ = pi1157 & ~new_n35584_;
  assign new_n35586_ = ~new_n35583_ & new_n35585_;
  assign new_n35587_ = ~pi0647 & new_n34920_;
  assign new_n35588_ = ~pi1157 & ~new_n35587_;
  assign new_n35589_ = pi0630 & ~new_n35588_;
  assign new_n35590_ = ~new_n35586_ & new_n35589_;
  assign new_n35591_ = ~new_n35582_ & ~new_n35590_;
  assign new_n35592_ = pi0787 & ~new_n35591_;
  assign new_n35593_ = ~pi0787 & ~new_n35366_;
  assign new_n35594_ = ~new_n35592_ & ~new_n35593_;
  assign new_n35595_ = ~pi0644 & new_n35594_;
  assign new_n35596_ = new_n35574_ & ~new_n35595_;
  assign new_n35597_ = new_n23689_ & new_n35018_;
  assign new_n35598_ = ~pi0644 & pi0715;
  assign new_n35599_ = new_n35597_ & new_n35598_;
  assign new_n35600_ = ~pi1160 & ~new_n35599_;
  assign new_n35601_ = ~new_n35596_ & new_n35600_;
  assign new_n35602_ = ~pi0644 & ~new_n35572_;
  assign new_n35603_ = pi0715 & ~new_n35602_;
  assign new_n35604_ = pi0644 & new_n35594_;
  assign new_n35605_ = new_n35603_ & ~new_n35604_;
  assign new_n35606_ = pi0644 & ~pi0715;
  assign new_n35607_ = new_n35597_ & new_n35606_;
  assign new_n35608_ = pi1160 & ~new_n35607_;
  assign new_n35609_ = ~new_n35605_ & new_n35608_;
  assign new_n35610_ = ~new_n35601_ & ~new_n35609_;
  assign new_n35611_ = pi0790 & ~new_n35610_;
  assign new_n35612_ = ~pi0790 & new_n35594_;
  assign new_n35613_ = ~po1038 & ~new_n35612_;
  assign new_n35614_ = ~new_n35611_ & new_n35613_;
  assign new_n35615_ = pi0622 & pi0639;
  assign new_n35616_ = ~new_n35614_ & new_n35615_;
  assign new_n35617_ = ~new_n20360_ & ~new_n35197_;
  assign new_n35618_ = new_n17804_ & new_n19334_;
  assign new_n35619_ = new_n34920_ & new_n35618_;
  assign new_n35620_ = ~new_n35617_ & ~new_n35619_;
  assign new_n35621_ = ~pi0644 & new_n35620_;
  assign new_n35622_ = ~pi1160 & new_n35574_;
  assign new_n35623_ = ~new_n35621_ & new_n35622_;
  assign new_n35624_ = pi0644 & new_n35620_;
  assign new_n35625_ = pi1160 & new_n35603_;
  assign new_n35626_ = ~new_n35624_ & new_n35625_;
  assign new_n35627_ = pi0790 & ~new_n35626_;
  assign new_n35628_ = ~new_n35623_ & new_n35627_;
  assign new_n35629_ = ~pi0790 & new_n35620_;
  assign new_n35630_ = ~po1038 & ~new_n35629_;
  assign new_n35631_ = ~new_n35628_ & new_n35630_;
  assign new_n35632_ = ~pi0622 & ~new_n35631_;
  assign new_n35633_ = ~pi0644 & pi1160;
  assign new_n35634_ = pi0644 & ~pi1160;
  assign new_n35635_ = ~new_n35633_ & ~new_n35634_;
  assign new_n35636_ = pi0790 & ~new_n35635_;
  assign new_n35637_ = ~po1038 & ~new_n35636_;
  assign new_n35638_ = new_n35597_ & new_n35637_;
  assign new_n35639_ = pi0622 & new_n35638_;
  assign new_n35640_ = ~pi0639 & ~new_n35639_;
  assign new_n35641_ = pi0209 & ~new_n35640_;
  assign new_n35642_ = ~new_n35632_ & new_n35641_;
  assign new_n35643_ = ~new_n35616_ & new_n35642_;
  assign po0366 = new_n35571_ | new_n35643_;
  assign new_n35645_ = pi0634 & new_n20915_;
  assign new_n35646_ = pi0633 & pi0947;
  assign new_n35647_ = ~new_n35645_ & ~new_n35646_;
  assign new_n35648_ = new_n17431_ & ~new_n35647_;
  assign new_n35649_ = pi0210 & ~new_n17431_;
  assign new_n35650_ = pi0038 & ~new_n35649_;
  assign new_n35651_ = ~new_n35648_ & new_n35650_;
  assign new_n35652_ = pi0210 & ~new_n16636_;
  assign new_n35653_ = ~po1101 & new_n35652_;
  assign new_n35654_ = pi0210 & po1101;
  assign new_n35655_ = ~new_n16740_ & new_n35654_;
  assign new_n35656_ = ~new_n35653_ & ~new_n35655_;
  assign new_n35657_ = ~pi0907 & new_n35656_;
  assign new_n35658_ = pi0634 & new_n16636_;
  assign new_n35659_ = ~new_n35652_ & ~new_n35658_;
  assign new_n35660_ = ~new_n6221_ & ~new_n35659_;
  assign new_n35661_ = pi0907 & ~new_n35660_;
  assign new_n35662_ = pi0210 & new_n16738_;
  assign new_n35663_ = pi0634 & ~new_n16738_;
  assign new_n35664_ = ~new_n35662_ & ~new_n35663_;
  assign new_n35665_ = new_n6221_ & ~new_n35664_;
  assign new_n35666_ = new_n35661_ & ~new_n35665_;
  assign new_n35667_ = ~pi0947 & ~new_n35666_;
  assign new_n35668_ = ~new_n35657_ & new_n35667_;
  assign new_n35669_ = ~new_n33436_ & ~new_n35652_;
  assign new_n35670_ = ~po1101 & new_n35669_;
  assign new_n35671_ = pi0947 & ~new_n35670_;
  assign new_n35672_ = po1101 & new_n35669_;
  assign new_n35673_ = ~new_n6221_ & ~new_n35672_;
  assign new_n35674_ = pi0633 & ~new_n16738_;
  assign new_n35675_ = ~new_n35662_ & ~new_n35674_;
  assign new_n35676_ = ~new_n6185_ & ~new_n35675_;
  assign new_n35677_ = ~new_n35673_ & ~new_n35676_;
  assign new_n35678_ = new_n35671_ & ~new_n35677_;
  assign new_n35679_ = new_n6238_ & ~new_n35678_;
  assign new_n35680_ = ~new_n35668_ & new_n35679_;
  assign new_n35681_ = new_n6215_ & new_n35659_;
  assign new_n35682_ = pi0907 & ~new_n35681_;
  assign new_n35683_ = ~new_n6215_ & new_n35664_;
  assign new_n35684_ = new_n35682_ & ~new_n35683_;
  assign new_n35685_ = pi0210 & ~new_n16941_;
  assign new_n35686_ = ~pi0907 & new_n35685_;
  assign new_n35687_ = ~new_n35684_ & ~new_n35686_;
  assign new_n35688_ = ~pi0947 & ~new_n35687_;
  assign new_n35689_ = new_n6215_ & new_n35669_;
  assign new_n35690_ = pi0947 & ~new_n35689_;
  assign new_n35691_ = ~new_n6215_ & new_n35675_;
  assign new_n35692_ = new_n35690_ & ~new_n35691_;
  assign new_n35693_ = ~new_n6238_ & ~new_n35692_;
  assign new_n35694_ = ~new_n35688_ & new_n35693_;
  assign new_n35695_ = ~new_n35680_ & ~new_n35694_;
  assign new_n35696_ = ~new_n3057_ & ~new_n35695_;
  assign new_n35697_ = new_n16636_ & ~new_n35647_;
  assign new_n35698_ = ~new_n35652_ & ~new_n35697_;
  assign new_n35699_ = new_n3057_ & new_n35698_;
  assign new_n35700_ = ~pi0223 & ~new_n35699_;
  assign new_n35701_ = ~new_n35696_ & new_n35700_;
  assign new_n35702_ = ~new_n16687_ & new_n35654_;
  assign new_n35703_ = ~new_n35653_ & ~new_n35702_;
  assign new_n35704_ = ~pi0907 & new_n35703_;
  assign new_n35705_ = pi0210 & new_n16660_;
  assign new_n35706_ = ~new_n33621_ & ~new_n35705_;
  assign new_n35707_ = new_n6221_ & ~new_n35706_;
  assign new_n35708_ = new_n35661_ & ~new_n35707_;
  assign new_n35709_ = ~pi0947 & ~new_n35708_;
  assign new_n35710_ = ~new_n35704_ & new_n35709_;
  assign new_n35711_ = pi0633 & ~new_n16660_;
  assign new_n35712_ = ~new_n35705_ & ~new_n35711_;
  assign new_n35713_ = ~new_n6185_ & ~new_n35712_;
  assign new_n35714_ = ~new_n35673_ & ~new_n35713_;
  assign new_n35715_ = new_n35671_ & ~new_n35714_;
  assign new_n35716_ = new_n6238_ & ~new_n35715_;
  assign new_n35717_ = ~new_n35710_ & new_n35716_;
  assign new_n35718_ = ~new_n6215_ & new_n35706_;
  assign new_n35719_ = new_n35682_ & ~new_n35718_;
  assign new_n35720_ = new_n6215_ & new_n16635_;
  assign new_n35721_ = new_n2754_ & new_n35720_;
  assign new_n35722_ = new_n35705_ & ~new_n35721_;
  assign new_n35723_ = ~new_n35719_ & ~new_n35722_;
  assign new_n35724_ = ~pi0947 & ~new_n35723_;
  assign new_n35725_ = ~new_n6215_ & new_n35712_;
  assign new_n35726_ = new_n35690_ & ~new_n35725_;
  assign new_n35727_ = ~new_n6238_ & ~new_n35726_;
  assign new_n35728_ = ~new_n35724_ & new_n35727_;
  assign new_n35729_ = pi0223 & ~new_n35728_;
  assign new_n35730_ = ~new_n35717_ & new_n35729_;
  assign new_n35731_ = ~pi0299 & ~new_n35730_;
  assign new_n35732_ = ~new_n35701_ & new_n35731_;
  assign new_n35733_ = ~new_n6211_ & ~new_n35685_;
  assign new_n35734_ = new_n6211_ & new_n35656_;
  assign new_n35735_ = ~pi0907 & ~new_n35734_;
  assign new_n35736_ = ~new_n35733_ & new_n35735_;
  assign new_n35737_ = ~new_n35684_ & ~new_n35736_;
  assign new_n35738_ = ~pi0947 & ~new_n35737_;
  assign new_n35739_ = ~new_n3467_ & ~new_n35692_;
  assign new_n35740_ = ~new_n35738_ & new_n35739_;
  assign new_n35741_ = new_n3467_ & new_n35698_;
  assign new_n35742_ = ~pi0215 & ~new_n35741_;
  assign new_n35743_ = ~new_n35740_ & new_n35742_;
  assign new_n35744_ = new_n6211_ & new_n35703_;
  assign new_n35745_ = ~new_n6211_ & ~new_n35722_;
  assign new_n35746_ = ~pi0907 & ~new_n35745_;
  assign new_n35747_ = ~new_n35744_ & new_n35746_;
  assign new_n35748_ = ~new_n35719_ & ~new_n35747_;
  assign new_n35749_ = ~pi0947 & ~new_n35748_;
  assign new_n35750_ = ~new_n35726_ & ~new_n35749_;
  assign new_n35751_ = pi0215 & ~new_n35750_;
  assign new_n35752_ = pi0299 & ~new_n35751_;
  assign new_n35753_ = ~new_n35743_ & new_n35752_;
  assign new_n35754_ = pi0039 & ~new_n35753_;
  assign new_n35755_ = ~new_n35732_ & new_n35754_;
  assign new_n35756_ = new_n17182_ & ~new_n35647_;
  assign new_n35757_ = pi0210 & ~new_n17182_;
  assign new_n35758_ = ~pi0299 & ~new_n35757_;
  assign new_n35759_ = ~new_n35756_ & new_n35758_;
  assign new_n35760_ = ~new_n17191_ & ~new_n35647_;
  assign new_n35761_ = pi0299 & ~new_n35760_;
  assign new_n35762_ = ~new_n17192_ & new_n35761_;
  assign new_n35763_ = ~pi0039 & ~new_n35762_;
  assign new_n35764_ = ~new_n35759_ & new_n35763_;
  assign new_n35765_ = ~pi0038 & ~new_n35764_;
  assign new_n35766_ = ~new_n35755_ & new_n35765_;
  assign new_n35767_ = ~new_n35651_ & ~new_n35766_;
  assign new_n35768_ = new_n10197_ & ~new_n35767_;
  assign new_n35769_ = ~pi0210 & ~new_n10197_;
  assign po0367 = ~new_n35768_ & ~new_n35769_;
  assign new_n35771_ = new_n3272_ & ~new_n21641_;
  assign new_n35772_ = pi0606 & new_n35771_;
  assign new_n35773_ = new_n3272_ & ~new_n21637_;
  assign new_n35774_ = ~pi0606 & new_n35773_;
  assign new_n35775_ = pi0643 & ~new_n35774_;
  assign new_n35776_ = ~new_n35772_ & new_n35775_;
  assign new_n35777_ = new_n3272_ & ~new_n21009_;
  assign new_n35778_ = pi0606 & new_n35777_;
  assign new_n35779_ = ~pi0606 & new_n17558_;
  assign new_n35780_ = ~pi0643 & ~new_n35779_;
  assign new_n35781_ = ~new_n35778_ & new_n35780_;
  assign new_n35782_ = ~po1038 & ~new_n35781_;
  assign new_n35783_ = ~new_n35776_ & new_n35782_;
  assign new_n35784_ = pi0211 & ~new_n35783_;
  assign new_n35785_ = new_n3272_ & new_n21626_;
  assign new_n35786_ = pi0606 & ~new_n35785_;
  assign new_n35787_ = new_n3272_ & new_n21623_;
  assign new_n35788_ = ~pi0606 & ~new_n35787_;
  assign new_n35789_ = pi0643 & ~new_n35788_;
  assign new_n35790_ = ~new_n35786_ & new_n35789_;
  assign new_n35791_ = new_n3272_ & new_n21033_;
  assign new_n35792_ = pi0606 & ~pi0643;
  assign new_n35793_ = new_n35791_ & new_n35792_;
  assign new_n35794_ = ~new_n35790_ & ~new_n35793_;
  assign new_n35795_ = ~pi0211 & ~po1038;
  assign new_n35796_ = ~new_n35794_ & new_n35795_;
  assign po0368 = new_n35784_ | new_n35796_;
  assign new_n35798_ = pi0607 & new_n35771_;
  assign new_n35799_ = ~pi0607 & new_n35773_;
  assign new_n35800_ = pi0638 & ~new_n35799_;
  assign new_n35801_ = ~new_n35798_ & new_n35800_;
  assign new_n35802_ = pi0607 & new_n35777_;
  assign new_n35803_ = ~pi0607 & new_n17558_;
  assign new_n35804_ = ~pi0638 & ~new_n35803_;
  assign new_n35805_ = ~new_n35802_ & new_n35804_;
  assign new_n35806_ = ~po1038 & ~new_n35805_;
  assign new_n35807_ = ~new_n35801_ & new_n35806_;
  assign new_n35808_ = ~pi0212 & ~new_n35807_;
  assign new_n35809_ = ~pi0607 & ~new_n35787_;
  assign new_n35810_ = pi0607 & ~new_n35785_;
  assign new_n35811_ = pi0638 & ~new_n35810_;
  assign new_n35812_ = ~new_n35809_ & new_n35811_;
  assign new_n35813_ = pi0607 & ~pi0638;
  assign new_n35814_ = new_n35791_ & new_n35813_;
  assign new_n35815_ = ~new_n35812_ & ~new_n35814_;
  assign new_n35816_ = pi0212 & ~po1038;
  assign new_n35817_ = ~new_n35815_ & new_n35816_;
  assign po0369 = new_n35808_ | new_n35817_;
  assign new_n35819_ = pi0213 & ~po1038;
  assign new_n35820_ = ~pi0622 & ~new_n35787_;
  assign new_n35821_ = pi0622 & ~new_n35785_;
  assign new_n35822_ = pi0639 & ~new_n35821_;
  assign new_n35823_ = ~new_n35820_ & new_n35822_;
  assign new_n35824_ = pi0622 & ~pi0639;
  assign new_n35825_ = new_n35791_ & new_n35824_;
  assign new_n35826_ = ~new_n35823_ & ~new_n35825_;
  assign new_n35827_ = new_n35819_ & ~new_n35826_;
  assign new_n35828_ = pi0639 & new_n35771_;
  assign new_n35829_ = ~pi0639 & new_n35777_;
  assign new_n35830_ = pi0622 & ~new_n35829_;
  assign new_n35831_ = ~new_n35828_ & new_n35830_;
  assign new_n35832_ = pi0639 & new_n35773_;
  assign new_n35833_ = ~pi0639 & new_n17558_;
  assign new_n35834_ = ~pi0622 & ~new_n35833_;
  assign new_n35835_ = ~new_n35832_ & new_n35834_;
  assign new_n35836_ = ~po1038 & ~new_n35835_;
  assign new_n35837_ = ~new_n35831_ & new_n35836_;
  assign new_n35838_ = ~pi0213 & ~new_n35837_;
  assign po0370 = new_n35827_ | new_n35838_;
  assign new_n35840_ = pi0623 & new_n35771_;
  assign new_n35841_ = ~pi0623 & new_n35773_;
  assign new_n35842_ = pi0710 & ~new_n35841_;
  assign new_n35843_ = ~new_n35840_ & new_n35842_;
  assign new_n35844_ = pi0623 & new_n35777_;
  assign new_n35845_ = ~pi0623 & new_n17558_;
  assign new_n35846_ = ~pi0710 & ~new_n35845_;
  assign new_n35847_ = ~new_n35844_ & new_n35846_;
  assign new_n35848_ = ~po1038 & ~new_n35847_;
  assign new_n35849_ = ~new_n35843_ & new_n35848_;
  assign new_n35850_ = ~pi0214 & ~new_n35849_;
  assign new_n35851_ = ~pi0623 & ~new_n35787_;
  assign new_n35852_ = pi0623 & ~new_n35785_;
  assign new_n35853_ = pi0710 & ~new_n35852_;
  assign new_n35854_ = ~new_n35851_ & new_n35853_;
  assign new_n35855_ = pi0623 & ~pi0710;
  assign new_n35856_ = new_n35791_ & new_n35855_;
  assign new_n35857_ = ~new_n35854_ & ~new_n35856_;
  assign new_n35858_ = pi0214 & ~po1038;
  assign new_n35859_ = ~new_n35857_ & new_n35858_;
  assign po0371 = new_n35850_ | new_n35859_;
  assign new_n35861_ = pi0215 & ~new_n10197_;
  assign new_n35862_ = ~pi0947 & new_n21319_;
  assign new_n35863_ = pi0681 & pi0907;
  assign new_n35864_ = ~pi0947 & new_n35863_;
  assign new_n35865_ = ~new_n6183_ & ~new_n16703_;
  assign new_n35866_ = new_n16629_ & new_n17264_;
  assign new_n35867_ = ~pi0642 & ~new_n35866_;
  assign new_n35868_ = ~new_n35865_ & new_n35867_;
  assign new_n35869_ = pi0947 & ~new_n35868_;
  assign new_n35870_ = ~new_n35864_ & ~new_n35869_;
  assign new_n35871_ = ~new_n35862_ & new_n35870_;
  assign new_n35872_ = pi0299 & ~new_n35871_;
  assign new_n35873_ = new_n21387_ & ~new_n35863_;
  assign new_n35874_ = ~pi0642 & new_n16740_;
  assign new_n35875_ = new_n6183_ & ~new_n35874_;
  assign new_n35876_ = new_n16707_ & new_n16742_;
  assign new_n35877_ = ~new_n6179_ & new_n16636_;
  assign new_n35878_ = ~pi0642 & new_n35877_;
  assign new_n35879_ = ~new_n6183_ & ~new_n35878_;
  assign new_n35880_ = ~new_n35876_ & new_n35879_;
  assign new_n35881_ = ~new_n35875_ & ~new_n35880_;
  assign new_n35882_ = new_n6238_ & ~new_n35881_;
  assign new_n35883_ = ~pi0642 & new_n16941_;
  assign new_n35884_ = ~new_n6238_ & ~new_n35883_;
  assign new_n35885_ = pi0947 & ~new_n35884_;
  assign new_n35886_ = ~new_n35882_ & new_n35885_;
  assign new_n35887_ = ~new_n3057_ & ~new_n35886_;
  assign new_n35888_ = ~new_n35873_ & new_n35887_;
  assign new_n35889_ = new_n3057_ & ~new_n16636_;
  assign new_n35890_ = pi0642 & pi0947;
  assign new_n35891_ = ~new_n35864_ & ~new_n35890_;
  assign new_n35892_ = new_n3057_ & ~new_n35891_;
  assign new_n35893_ = ~pi0223 & ~new_n35892_;
  assign new_n35894_ = ~new_n35889_ & new_n35893_;
  assign new_n35895_ = ~new_n35888_ & new_n35894_;
  assign new_n35896_ = ~new_n6183_ & ~new_n16693_;
  assign new_n35897_ = new_n6183_ & ~new_n16687_;
  assign new_n35898_ = ~pi0642 & ~new_n35897_;
  assign new_n35899_ = ~new_n35896_ & new_n35898_;
  assign new_n35900_ = new_n6238_ & ~new_n35899_;
  assign new_n35901_ = ~new_n6238_ & ~new_n35868_;
  assign new_n35902_ = pi0947 & ~new_n35901_;
  assign new_n35903_ = ~new_n35900_ & new_n35902_;
  assign new_n35904_ = ~new_n21082_ & ~new_n35903_;
  assign new_n35905_ = pi0223 & ~new_n35864_;
  assign new_n35906_ = ~new_n35904_ & new_n35905_;
  assign new_n35907_ = ~pi0299 & ~new_n35906_;
  assign new_n35908_ = ~new_n35895_ & new_n35907_;
  assign new_n35909_ = ~new_n35872_ & ~new_n35908_;
  assign new_n35910_ = pi0215 & ~new_n35909_;
  assign new_n35911_ = new_n16756_ & new_n35864_;
  assign new_n35912_ = pi0642 & ~new_n16630_;
  assign new_n35913_ = new_n16636_ & new_n35912_;
  assign new_n35914_ = pi0642 & new_n16630_;
  assign new_n35915_ = ~new_n17283_ & new_n35914_;
  assign new_n35916_ = ~new_n17304_ & new_n35915_;
  assign new_n35917_ = ~new_n35913_ & ~new_n35916_;
  assign new_n35918_ = pi0947 & ~new_n35917_;
  assign new_n35919_ = new_n6238_ & ~new_n35918_;
  assign new_n35920_ = ~new_n35911_ & new_n35919_;
  assign new_n35921_ = new_n16774_ & new_n35863_;
  assign new_n35922_ = ~pi0947 & ~new_n35921_;
  assign new_n35923_ = ~new_n6183_ & new_n16771_;
  assign new_n35924_ = ~new_n16940_ & ~new_n35923_;
  assign new_n35925_ = new_n35914_ & new_n35924_;
  assign new_n35926_ = ~new_n16771_ & new_n35912_;
  assign new_n35927_ = pi0947 & ~new_n35926_;
  assign new_n35928_ = ~new_n35925_ & new_n35927_;
  assign new_n35929_ = ~new_n35922_ & ~new_n35928_;
  assign new_n35930_ = ~new_n6238_ & ~new_n35929_;
  assign new_n35931_ = ~new_n3057_ & ~new_n35930_;
  assign new_n35932_ = ~new_n35920_ & new_n35931_;
  assign new_n35933_ = new_n16636_ & new_n35892_;
  assign new_n35934_ = ~pi0223 & ~new_n35933_;
  assign new_n35935_ = ~new_n35932_ & new_n35934_;
  assign new_n35936_ = new_n6238_ & ~new_n16693_;
  assign new_n35937_ = new_n35863_ & ~new_n35936_;
  assign new_n35938_ = ~pi0947 & ~new_n35937_;
  assign new_n35939_ = pi0947 & ~new_n16701_;
  assign new_n35940_ = ~new_n16703_ & ~new_n35939_;
  assign new_n35941_ = ~new_n6238_ & new_n35940_;
  assign new_n35942_ = ~new_n17278_ & new_n35915_;
  assign new_n35943_ = pi0947 & ~new_n35913_;
  assign new_n35944_ = ~new_n35942_ & new_n35943_;
  assign new_n35945_ = ~new_n35941_ & ~new_n35944_;
  assign new_n35946_ = ~new_n35938_ & new_n35945_;
  assign new_n35947_ = pi0223 & ~new_n35946_;
  assign new_n35948_ = ~new_n35935_ & ~new_n35947_;
  assign new_n35949_ = ~pi0299 & ~new_n35948_;
  assign new_n35950_ = ~new_n3467_ & new_n35929_;
  assign new_n35951_ = new_n16865_ & ~new_n35891_;
  assign new_n35952_ = pi0299 & ~new_n35951_;
  assign new_n35953_ = ~new_n35950_ & new_n35952_;
  assign new_n35954_ = ~pi0215 & ~new_n35953_;
  assign new_n35955_ = ~new_n35949_ & new_n35954_;
  assign new_n35956_ = ~new_n35910_ & ~new_n35955_;
  assign new_n35957_ = pi0039 & ~new_n35956_;
  assign new_n35958_ = pi0215 & ~new_n17182_;
  assign new_n35959_ = new_n17182_ & ~new_n35891_;
  assign new_n35960_ = ~pi0299 & ~new_n35959_;
  assign new_n35961_ = ~new_n35958_ & new_n35960_;
  assign new_n35962_ = new_n17193_ & ~new_n35891_;
  assign new_n35963_ = pi0215 & ~new_n17193_;
  assign new_n35964_ = pi0299 & ~new_n35963_;
  assign new_n35965_ = ~new_n35962_ & new_n35964_;
  assign new_n35966_ = ~pi0039 & ~new_n35965_;
  assign new_n35967_ = ~new_n35961_ & new_n35966_;
  assign new_n35968_ = ~pi0038 & ~new_n35967_;
  assign new_n35969_ = ~new_n35957_ & new_n35968_;
  assign new_n35970_ = pi0215 & ~new_n17431_;
  assign new_n35971_ = new_n17431_ & ~new_n35891_;
  assign new_n35972_ = pi0038 & ~new_n35971_;
  assign new_n35973_ = ~new_n35970_ & new_n35972_;
  assign new_n35974_ = new_n10197_ & ~new_n35973_;
  assign new_n35975_ = ~new_n35969_ & new_n35974_;
  assign po0372 = new_n35861_ | new_n35975_;
  assign new_n35977_ = pi0216 & ~new_n17431_;
  assign new_n35978_ = pi0662 & pi0907;
  assign new_n35979_ = ~pi0947 & new_n35978_;
  assign new_n35980_ = pi0614 & pi0947;
  assign new_n35981_ = ~new_n35979_ & ~new_n35980_;
  assign new_n35982_ = new_n17431_ & ~new_n35981_;
  assign new_n35983_ = pi0038 & ~new_n35982_;
  assign new_n35984_ = ~new_n35977_ & new_n35983_;
  assign new_n35985_ = ~pi0947 & new_n20993_;
  assign new_n35986_ = ~pi0614 & new_n16941_;
  assign new_n35987_ = pi0947 & ~new_n35986_;
  assign new_n35988_ = ~new_n35979_ & ~new_n35987_;
  assign new_n35989_ = ~new_n35985_ & new_n35988_;
  assign new_n35990_ = pi0216 & ~new_n35989_;
  assign new_n35991_ = new_n35924_ & new_n35980_;
  assign new_n35992_ = new_n16774_ & new_n35979_;
  assign new_n35993_ = ~new_n35991_ & ~new_n35992_;
  assign new_n35994_ = new_n5766_ & ~new_n35993_;
  assign new_n35995_ = new_n16865_ & ~new_n35981_;
  assign new_n35996_ = ~new_n35994_ & ~new_n35995_;
  assign new_n35997_ = ~new_n35990_ & new_n35996_;
  assign new_n35998_ = ~pi0215 & ~new_n35997_;
  assign new_n35999_ = ~new_n16873_ & ~new_n33394_;
  assign new_n36000_ = ~new_n33393_ & new_n35999_;
  assign new_n36001_ = new_n17298_ & ~new_n36000_;
  assign new_n36002_ = ~pi0614 & ~new_n16660_;
  assign new_n36003_ = new_n6183_ & new_n36002_;
  assign new_n36004_ = ~new_n36001_ & ~new_n36003_;
  assign new_n36005_ = pi0947 & new_n36004_;
  assign new_n36006_ = pi0216 & ~new_n35979_;
  assign new_n36007_ = ~new_n36005_ & new_n36006_;
  assign new_n36008_ = ~new_n35862_ & new_n36007_;
  assign new_n36009_ = new_n16703_ & new_n35978_;
  assign new_n36010_ = ~pi0947 & ~new_n36009_;
  assign new_n36011_ = ~new_n17278_ & new_n17306_;
  assign new_n36012_ = pi0947 & ~new_n17309_;
  assign new_n36013_ = ~new_n36011_ & new_n36012_;
  assign new_n36014_ = pi0947 & new_n16701_;
  assign new_n36015_ = ~new_n36013_ & ~new_n36014_;
  assign new_n36016_ = ~new_n36010_ & new_n36015_;
  assign new_n36017_ = ~pi0216 & ~new_n36016_;
  assign new_n36018_ = pi0215 & ~new_n36017_;
  assign new_n36019_ = ~new_n36008_ & new_n36018_;
  assign new_n36020_ = pi0299 & ~new_n36019_;
  assign new_n36021_ = ~new_n35998_ & new_n36020_;
  assign new_n36022_ = pi0947 & ~new_n17303_;
  assign new_n36023_ = ~pi0947 & new_n17313_;
  assign new_n36024_ = ~new_n35978_ & new_n36023_;
  assign new_n36025_ = ~new_n36022_ & ~new_n36024_;
  assign new_n36026_ = new_n6238_ & ~new_n36025_;
  assign new_n36027_ = ~pi0947 & ~new_n17320_;
  assign new_n36028_ = ~new_n6238_ & ~new_n35979_;
  assign new_n36029_ = ~new_n35987_ & new_n36028_;
  assign new_n36030_ = ~new_n36027_ & new_n36029_;
  assign new_n36031_ = ~new_n3057_ & ~new_n36030_;
  assign new_n36032_ = ~new_n36026_ & new_n36031_;
  assign new_n36033_ = new_n3057_ & ~new_n35981_;
  assign new_n36034_ = ~pi0223 & ~new_n36033_;
  assign new_n36035_ = ~new_n35889_ & new_n36034_;
  assign new_n36036_ = ~new_n36032_ & new_n36035_;
  assign new_n36037_ = ~pi0616 & new_n16689_;
  assign new_n36038_ = ~new_n6183_ & ~new_n17287_;
  assign new_n36039_ = ~new_n36037_ & new_n36038_;
  assign new_n36040_ = ~pi0614 & ~new_n35897_;
  assign new_n36041_ = ~new_n36039_ & new_n36040_;
  assign new_n36042_ = new_n6238_ & ~new_n36041_;
  assign new_n36043_ = ~new_n6238_ & new_n36004_;
  assign new_n36044_ = pi0947 & ~new_n36043_;
  assign new_n36045_ = ~new_n36042_ & new_n36044_;
  assign new_n36046_ = ~new_n21082_ & ~new_n36045_;
  assign new_n36047_ = pi0223 & ~new_n35979_;
  assign new_n36048_ = ~new_n36046_ & new_n36047_;
  assign new_n36049_ = pi0216 & ~new_n36048_;
  assign new_n36050_ = ~new_n36036_ & new_n36049_;
  assign new_n36051_ = new_n16756_ & new_n35979_;
  assign new_n36052_ = pi0947 & ~new_n17310_;
  assign new_n36053_ = new_n6238_ & ~new_n36052_;
  assign new_n36054_ = ~new_n36051_ & new_n36053_;
  assign new_n36055_ = ~new_n6238_ & new_n35993_;
  assign new_n36056_ = ~new_n3057_ & ~new_n36055_;
  assign new_n36057_ = ~new_n36054_ & new_n36056_;
  assign new_n36058_ = new_n16636_ & new_n36033_;
  assign new_n36059_ = ~pi0223 & ~new_n36058_;
  assign new_n36060_ = ~new_n36057_ & new_n36059_;
  assign new_n36061_ = ~new_n35936_ & new_n35978_;
  assign new_n36062_ = ~pi0947 & ~new_n36061_;
  assign new_n36063_ = ~new_n35941_ & ~new_n36013_;
  assign new_n36064_ = ~new_n36062_ & new_n36063_;
  assign new_n36065_ = pi0223 & ~new_n36064_;
  assign new_n36066_ = ~pi0216 & ~new_n36065_;
  assign new_n36067_ = ~new_n36060_ & new_n36066_;
  assign new_n36068_ = ~pi0299 & ~new_n36067_;
  assign new_n36069_ = ~new_n36050_ & new_n36068_;
  assign new_n36070_ = pi0039 & ~new_n36069_;
  assign new_n36071_ = ~new_n36021_ & new_n36070_;
  assign new_n36072_ = pi0216 & ~new_n17182_;
  assign new_n36073_ = new_n17182_ & ~new_n35981_;
  assign new_n36074_ = ~pi0299 & ~new_n36073_;
  assign new_n36075_ = ~new_n36072_ & new_n36074_;
  assign new_n36076_ = new_n17193_ & ~new_n35981_;
  assign new_n36077_ = pi0216 & ~new_n17193_;
  assign new_n36078_ = pi0299 & ~new_n36077_;
  assign new_n36079_ = ~new_n36076_ & new_n36078_;
  assign new_n36080_ = ~pi0039 & ~new_n36079_;
  assign new_n36081_ = ~new_n36075_ & new_n36080_;
  assign new_n36082_ = ~pi0038 & ~new_n36081_;
  assign new_n36083_ = ~new_n36071_ & new_n36082_;
  assign new_n36084_ = ~new_n35984_ & ~new_n36083_;
  assign new_n36085_ = new_n10197_ & ~new_n36084_;
  assign new_n36086_ = ~pi0216 & ~new_n10197_;
  assign po0373 = ~new_n36085_ & ~new_n36086_;
  assign new_n36088_ = ~pi0695 & ~new_n35522_;
  assign new_n36089_ = pi0695 & ~new_n35524_;
  assign new_n36090_ = ~pi0217 & ~new_n36089_;
  assign new_n36091_ = ~new_n36088_ & new_n36090_;
  assign new_n36092_ = ~pi0695 & new_n35631_;
  assign new_n36093_ = pi0217 & ~new_n36092_;
  assign new_n36094_ = ~pi0612 & ~new_n36093_;
  assign new_n36095_ = ~new_n36091_ & new_n36094_;
  assign new_n36096_ = ~pi0695 & ~new_n35558_;
  assign new_n36097_ = pi0695 & ~new_n35566_;
  assign new_n36098_ = ~pi0217 & ~new_n36097_;
  assign new_n36099_ = ~new_n36096_ & new_n36098_;
  assign new_n36100_ = ~pi0695 & new_n35614_;
  assign new_n36101_ = pi0695 & new_n35638_;
  assign new_n36102_ = pi0217 & ~new_n36101_;
  assign new_n36103_ = ~new_n36100_ & new_n36102_;
  assign new_n36104_ = pi0612 & ~new_n36103_;
  assign new_n36105_ = ~new_n36099_ & new_n36104_;
  assign po0374 = new_n36095_ | new_n36105_;
  assign new_n36107_ = ~new_n34786_ & ~new_n34825_;
  assign new_n36108_ = new_n34786_ & ~new_n34891_;
  assign new_n36109_ = ~new_n36107_ & ~new_n36108_;
  assign new_n36110_ = ~pi0218 & ~new_n36109_;
  assign new_n36111_ = new_n34786_ & new_n34899_;
  assign new_n36112_ = pi0218 & ~new_n36111_;
  assign po0375 = ~new_n36110_ & ~new_n36112_;
  assign new_n36114_ = ~pi0219 & ~po1038;
  assign new_n36115_ = ~pi0617 & ~new_n35787_;
  assign new_n36116_ = pi0617 & ~new_n35785_;
  assign new_n36117_ = pi0637 & ~new_n36116_;
  assign new_n36118_ = ~new_n36115_ & new_n36117_;
  assign new_n36119_ = pi0617 & ~pi0637;
  assign new_n36120_ = new_n35791_ & new_n36119_;
  assign new_n36121_ = ~new_n36118_ & ~new_n36120_;
  assign new_n36122_ = new_n36114_ & ~new_n36121_;
  assign new_n36123_ = pi0617 & new_n35771_;
  assign new_n36124_ = ~pi0617 & new_n35773_;
  assign new_n36125_ = pi0637 & ~new_n36124_;
  assign new_n36126_ = ~new_n36123_ & new_n36125_;
  assign new_n36127_ = pi0617 & new_n35777_;
  assign new_n36128_ = ~pi0617 & new_n17558_;
  assign new_n36129_ = ~pi0637 & ~new_n36128_;
  assign new_n36130_ = ~new_n36127_ & new_n36129_;
  assign new_n36131_ = ~po1038 & ~new_n36130_;
  assign new_n36132_ = ~new_n36126_ & new_n36131_;
  assign new_n36133_ = pi0219 & ~new_n36132_;
  assign po0376 = new_n36122_ | new_n36133_;
  assign new_n36135_ = ~new_n34619_ & ~new_n34910_;
  assign new_n36136_ = ~new_n34765_ & new_n34910_;
  assign new_n36137_ = ~new_n36135_ & ~new_n36136_;
  assign new_n36138_ = ~pi0220 & ~new_n36137_;
  assign new_n36139_ = new_n34774_ & new_n34910_;
  assign new_n36140_ = pi0220 & ~new_n36139_;
  assign po0377 = ~new_n36138_ & ~new_n36140_;
  assign new_n36142_ = pi0221 & ~new_n17431_;
  assign new_n36143_ = pi0661 & pi0907;
  assign new_n36144_ = ~pi0947 & new_n36143_;
  assign new_n36145_ = pi0616 & pi0947;
  assign new_n36146_ = ~new_n36144_ & ~new_n36145_;
  assign new_n36147_ = new_n17431_ & ~new_n36146_;
  assign new_n36148_ = pi0038 & ~new_n36147_;
  assign new_n36149_ = ~new_n36142_ & new_n36148_;
  assign new_n36150_ = ~new_n20993_ & ~new_n36143_;
  assign new_n36151_ = ~pi0947 & ~new_n36150_;
  assign new_n36152_ = ~new_n6185_ & new_n16754_;
  assign new_n36153_ = ~new_n16770_ & ~new_n36152_;
  assign new_n36154_ = new_n17275_ & ~new_n36153_;
  assign new_n36155_ = ~new_n35883_ & ~new_n35925_;
  assign new_n36156_ = new_n17279_ & ~new_n36155_;
  assign new_n36157_ = pi0947 & ~new_n36156_;
  assign new_n36158_ = ~new_n36154_ & new_n36157_;
  assign new_n36159_ = pi0221 & ~new_n36158_;
  assign new_n36160_ = ~new_n36151_ & new_n36159_;
  assign new_n36161_ = new_n35924_ & new_n36145_;
  assign new_n36162_ = new_n16774_ & new_n36144_;
  assign new_n36163_ = ~new_n36161_ & ~new_n36162_;
  assign new_n36164_ = pi0216 & ~new_n36163_;
  assign new_n36165_ = new_n16636_ & ~new_n36146_;
  assign new_n36166_ = ~pi0216 & new_n36165_;
  assign new_n36167_ = ~pi0221 & ~new_n36166_;
  assign new_n36168_ = ~new_n36164_ & new_n36167_;
  assign new_n36169_ = ~pi0215 & ~new_n36168_;
  assign new_n36170_ = ~new_n36160_ & new_n36169_;
  assign new_n36171_ = ~new_n16690_ & ~new_n16701_;
  assign new_n36172_ = ~new_n6183_ & ~new_n36171_;
  assign new_n36173_ = ~pi0616 & ~new_n35866_;
  assign new_n36174_ = ~new_n36172_ & new_n36173_;
  assign new_n36175_ = pi0947 & ~new_n36174_;
  assign new_n36176_ = pi0221 & ~new_n36144_;
  assign new_n36177_ = ~new_n36175_ & new_n36176_;
  assign new_n36178_ = ~new_n35862_ & new_n36177_;
  assign new_n36179_ = pi0947 & ~new_n17289_;
  assign new_n36180_ = ~new_n36144_ & ~new_n36179_;
  assign new_n36181_ = ~new_n35940_ & ~new_n36180_;
  assign new_n36182_ = ~pi0221 & ~new_n36181_;
  assign new_n36183_ = pi0215 & ~new_n36182_;
  assign new_n36184_ = ~new_n36178_ & new_n36183_;
  assign new_n36185_ = pi0299 & ~new_n36184_;
  assign new_n36186_ = ~new_n36170_ & new_n36185_;
  assign new_n36187_ = new_n16754_ & new_n17275_;
  assign new_n36188_ = new_n17303_ & ~new_n17307_;
  assign new_n36189_ = new_n17279_ & ~new_n36188_;
  assign new_n36190_ = ~new_n36187_ & ~new_n36189_;
  assign new_n36191_ = pi0947 & ~new_n36190_;
  assign new_n36192_ = new_n6238_ & ~new_n36023_;
  assign new_n36193_ = ~new_n36191_ & new_n36192_;
  assign new_n36194_ = ~new_n36027_ & ~new_n36158_;
  assign new_n36195_ = ~new_n6238_ & ~new_n36194_;
  assign new_n36196_ = ~new_n36144_ & ~new_n36195_;
  assign new_n36197_ = ~new_n36193_ & new_n36196_;
  assign new_n36198_ = ~new_n3057_ & ~new_n36197_;
  assign new_n36199_ = new_n3057_ & new_n36165_;
  assign new_n36200_ = ~pi0223 & ~new_n36199_;
  assign new_n36201_ = ~new_n35889_ & new_n36200_;
  assign new_n36202_ = ~new_n36198_ & new_n36201_;
  assign new_n36203_ = ~pi0947 & ~new_n17272_;
  assign new_n36204_ = ~new_n36175_ & ~new_n36203_;
  assign new_n36205_ = ~new_n6238_ & ~new_n36204_;
  assign new_n36206_ = ~pi0947 & new_n17292_;
  assign new_n36207_ = pi0947 & ~new_n17282_;
  assign new_n36208_ = new_n6238_ & ~new_n36207_;
  assign new_n36209_ = ~new_n36206_ & new_n36208_;
  assign new_n36210_ = pi0223 & ~new_n36144_;
  assign new_n36211_ = ~new_n36209_ & new_n36210_;
  assign new_n36212_ = ~new_n36205_ & new_n36211_;
  assign new_n36213_ = pi0221 & ~new_n36212_;
  assign new_n36214_ = ~new_n36202_ & new_n36213_;
  assign new_n36215_ = new_n16756_ & new_n36144_;
  assign new_n36216_ = new_n17285_ & ~new_n17304_;
  assign new_n36217_ = ~new_n17288_ & ~new_n36216_;
  assign new_n36218_ = pi0947 & ~new_n36217_;
  assign new_n36219_ = new_n6238_ & ~new_n36218_;
  assign new_n36220_ = ~new_n36215_ & new_n36219_;
  assign new_n36221_ = ~new_n6238_ & new_n36163_;
  assign new_n36222_ = ~new_n3057_ & ~new_n36221_;
  assign new_n36223_ = ~new_n36220_ & new_n36222_;
  assign new_n36224_ = new_n36200_ & ~new_n36223_;
  assign new_n36225_ = new_n35936_ & ~new_n36179_;
  assign new_n36226_ = ~new_n35941_ & ~new_n36180_;
  assign new_n36227_ = ~new_n36225_ & new_n36226_;
  assign new_n36228_ = pi0223 & ~new_n36227_;
  assign new_n36229_ = ~pi0221 & ~new_n36228_;
  assign new_n36230_ = ~new_n36224_ & new_n36229_;
  assign new_n36231_ = ~pi0299 & ~new_n36230_;
  assign new_n36232_ = ~new_n36214_ & new_n36231_;
  assign new_n36233_ = pi0039 & ~new_n36232_;
  assign new_n36234_ = ~new_n36186_ & new_n36233_;
  assign new_n36235_ = pi0221 & ~new_n17182_;
  assign new_n36236_ = new_n17182_ & ~new_n36146_;
  assign new_n36237_ = ~pi0299 & ~new_n36236_;
  assign new_n36238_ = ~new_n36235_ & new_n36237_;
  assign new_n36239_ = new_n17193_ & ~new_n36146_;
  assign new_n36240_ = pi0221 & ~new_n17193_;
  assign new_n36241_ = pi0299 & ~new_n36240_;
  assign new_n36242_ = ~new_n36239_ & new_n36241_;
  assign new_n36243_ = ~pi0039 & ~new_n36242_;
  assign new_n36244_ = ~new_n36238_ & new_n36243_;
  assign new_n36245_ = ~pi0038 & ~new_n36244_;
  assign new_n36246_ = ~new_n36234_ & new_n36245_;
  assign new_n36247_ = ~new_n36149_ & ~new_n36246_;
  assign new_n36248_ = new_n10197_ & ~new_n36247_;
  assign new_n36249_ = ~pi0221 & ~new_n10197_;
  assign po0378 = ~new_n36248_ & ~new_n36249_;
  assign new_n36251_ = ~pi0223 & ~new_n17322_;
  assign new_n36252_ = ~new_n17295_ & ~new_n36251_;
  assign new_n36253_ = ~pi0299 & ~new_n36252_;
  assign new_n36254_ = pi0039 & ~new_n36253_;
  assign new_n36255_ = ~new_n17346_ & new_n36254_;
  assign new_n36256_ = ~pi0038 & ~new_n18106_;
  assign new_n36257_ = ~new_n36255_ & new_n36256_;
  assign new_n36258_ = new_n18873_ & ~new_n36257_;
  assign new_n36259_ = pi0222 & ~new_n36258_;
  assign new_n36260_ = new_n17968_ & ~new_n36259_;
  assign new_n36261_ = pi0222 & ~new_n3272_;
  assign new_n36262_ = pi0616 & ~new_n16822_;
  assign new_n36263_ = ~pi0616 & new_n36153_;
  assign new_n36264_ = ~new_n36262_ & ~new_n36263_;
  assign new_n36265_ = ~new_n16629_ & ~new_n36264_;
  assign new_n36266_ = ~new_n6181_ & new_n36264_;
  assign new_n36267_ = pi0616 & new_n16639_;
  assign new_n36268_ = new_n16779_ & ~new_n36267_;
  assign new_n36269_ = ~new_n16817_ & ~new_n36268_;
  assign new_n36270_ = new_n6181_ & ~new_n36269_;
  assign new_n36271_ = new_n16629_ & ~new_n36270_;
  assign new_n36272_ = ~new_n36266_ & new_n36271_;
  assign new_n36273_ = ~new_n36265_ & ~new_n36272_;
  assign new_n36274_ = ~new_n6238_ & new_n36273_;
  assign new_n36275_ = pi0616 & ~new_n16842_;
  assign new_n36276_ = ~new_n16755_ & ~new_n36275_;
  assign new_n36277_ = ~new_n16629_ & ~new_n36276_;
  assign new_n36278_ = ~new_n6181_ & new_n36276_;
  assign new_n36279_ = new_n6181_ & ~new_n36267_;
  assign new_n36280_ = new_n16740_ & new_n36279_;
  assign new_n36281_ = new_n16629_ & ~new_n36280_;
  assign new_n36282_ = ~new_n36278_ & new_n36281_;
  assign new_n36283_ = ~new_n36277_ & ~new_n36282_;
  assign new_n36284_ = new_n6238_ & new_n36283_;
  assign new_n36285_ = pi0222 & ~new_n36284_;
  assign new_n36286_ = ~new_n36274_ & new_n36285_;
  assign new_n36287_ = ~new_n16771_ & new_n36267_;
  assign new_n36288_ = ~new_n16629_ & ~new_n36287_;
  assign new_n36289_ = ~new_n6181_ & new_n36287_;
  assign new_n36290_ = pi0616 & new_n6181_;
  assign new_n36291_ = new_n16780_ & new_n36290_;
  assign new_n36292_ = new_n16629_ & ~new_n36291_;
  assign new_n36293_ = ~new_n36289_ & new_n36292_;
  assign new_n36294_ = ~new_n36288_ & ~new_n36293_;
  assign new_n36295_ = ~new_n6238_ & new_n36294_;
  assign new_n36296_ = ~new_n6183_ & new_n16661_;
  assign new_n36297_ = ~new_n17399_ & ~new_n36296_;
  assign new_n36298_ = pi0616 & ~new_n36297_;
  assign new_n36299_ = new_n6238_ & new_n36298_;
  assign new_n36300_ = pi0224 & ~new_n36299_;
  assign new_n36301_ = ~new_n36295_ & new_n36300_;
  assign new_n36302_ = new_n16639_ & new_n17287_;
  assign new_n36303_ = ~pi0224 & ~new_n36302_;
  assign new_n36304_ = ~pi0222 & ~new_n36303_;
  assign new_n36305_ = ~new_n36301_ & new_n36304_;
  assign new_n36306_ = ~pi0223 & ~new_n36305_;
  assign new_n36307_ = ~new_n36286_ & new_n36306_;
  assign new_n36308_ = ~new_n16692_ & ~new_n36275_;
  assign new_n36309_ = ~new_n16629_ & ~new_n36308_;
  assign new_n36310_ = ~new_n6181_ & new_n36308_;
  assign new_n36311_ = new_n16687_ & new_n36279_;
  assign new_n36312_ = new_n16629_ & ~new_n36311_;
  assign new_n36313_ = ~new_n36310_ & new_n36312_;
  assign new_n36314_ = ~new_n36309_ & ~new_n36313_;
  assign new_n36315_ = new_n6238_ & new_n36314_;
  assign new_n36316_ = pi0616 & ~new_n16869_;
  assign new_n36317_ = new_n16703_ & ~new_n36316_;
  assign new_n36318_ = ~new_n16629_ & ~new_n36317_;
  assign new_n36319_ = ~new_n6181_ & ~new_n16703_;
  assign new_n36320_ = ~new_n17264_ & ~new_n36316_;
  assign new_n36321_ = ~new_n36319_ & new_n36320_;
  assign new_n36322_ = new_n16629_ & ~new_n36321_;
  assign new_n36323_ = ~new_n36318_ & ~new_n36322_;
  assign new_n36324_ = ~new_n6238_ & new_n36323_;
  assign new_n36325_ = pi0222 & ~new_n36324_;
  assign new_n36326_ = ~new_n36315_ & new_n36325_;
  assign new_n36327_ = ~new_n16669_ & ~new_n36296_;
  assign new_n36328_ = pi0616 & ~new_n36327_;
  assign new_n36329_ = ~pi0222 & new_n36328_;
  assign new_n36330_ = ~new_n17419_ & new_n36329_;
  assign new_n36331_ = pi0223 & ~new_n36330_;
  assign new_n36332_ = ~new_n36326_ & new_n36331_;
  assign new_n36333_ = ~new_n36307_ & ~new_n36332_;
  assign new_n36334_ = ~pi0299 & ~new_n36333_;
  assign new_n36335_ = ~new_n6212_ & new_n36273_;
  assign new_n36336_ = new_n6212_ & new_n36283_;
  assign new_n36337_ = pi0222 & ~new_n36336_;
  assign new_n36338_ = ~new_n36335_ & new_n36337_;
  assign new_n36339_ = ~new_n6212_ & ~new_n36294_;
  assign new_n36340_ = new_n6212_ & ~new_n36298_;
  assign new_n36341_ = ~pi0222 & ~new_n36340_;
  assign new_n36342_ = ~new_n36339_ & new_n36341_;
  assign new_n36343_ = ~new_n3467_ & ~new_n36342_;
  assign new_n36344_ = ~new_n36338_ & new_n36343_;
  assign new_n36345_ = pi0222 & ~new_n16636_;
  assign new_n36346_ = new_n3467_ & ~new_n36345_;
  assign new_n36347_ = ~new_n36302_ & new_n36346_;
  assign new_n36348_ = ~pi0215 & ~new_n36347_;
  assign new_n36349_ = ~new_n36344_ & new_n36348_;
  assign new_n36350_ = ~new_n17409_ & new_n36329_;
  assign new_n36351_ = new_n6212_ & new_n36314_;
  assign new_n36352_ = ~new_n6212_ & new_n36323_;
  assign new_n36353_ = pi0222 & ~new_n36352_;
  assign new_n36354_ = ~new_n36351_ & new_n36353_;
  assign new_n36355_ = ~new_n36350_ & ~new_n36354_;
  assign new_n36356_ = pi0215 & ~new_n36355_;
  assign new_n36357_ = pi0299 & ~new_n36356_;
  assign new_n36358_ = ~new_n36349_ & new_n36357_;
  assign new_n36359_ = pi0039 & ~new_n36358_;
  assign new_n36360_ = ~new_n36334_ & new_n36359_;
  assign new_n36361_ = pi0222 & new_n17226_;
  assign new_n36362_ = ~pi0222 & ~new_n17215_;
  assign new_n36363_ = ~pi0616 & new_n17215_;
  assign new_n36364_ = ~pi0039 & ~new_n36363_;
  assign new_n36365_ = ~new_n36362_ & new_n36364_;
  assign new_n36366_ = ~new_n36361_ & new_n36365_;
  assign new_n36367_ = ~pi0038 & ~new_n36366_;
  assign new_n36368_ = ~new_n36360_ & new_n36367_;
  assign new_n36369_ = pi0222 & ~new_n17431_;
  assign new_n36370_ = pi0038 & ~new_n36369_;
  assign new_n36371_ = pi0616 & new_n17433_;
  assign new_n36372_ = new_n36370_ & ~new_n36371_;
  assign new_n36373_ = new_n3272_ & ~new_n36372_;
  assign new_n36374_ = ~new_n36368_ & new_n36373_;
  assign new_n36375_ = ~new_n36261_ & ~new_n36374_;
  assign new_n36376_ = ~new_n17590_ & ~new_n36375_;
  assign new_n36377_ = new_n17590_ & new_n36259_;
  assign new_n36378_ = ~new_n36376_ & ~new_n36377_;
  assign new_n36379_ = ~pi0785 & ~new_n36378_;
  assign new_n36380_ = pi0609 & new_n36378_;
  assign new_n36381_ = ~pi0609 & ~new_n36259_;
  assign new_n36382_ = pi1155 & ~new_n36381_;
  assign new_n36383_ = ~new_n36380_ & new_n36382_;
  assign new_n36384_ = ~pi0609 & new_n36378_;
  assign new_n36385_ = pi0609 & ~new_n36259_;
  assign new_n36386_ = ~pi1155 & ~new_n36385_;
  assign new_n36387_ = ~new_n36384_ & new_n36386_;
  assign new_n36388_ = ~new_n36383_ & ~new_n36387_;
  assign new_n36389_ = pi0785 & ~new_n36388_;
  assign new_n36390_ = ~new_n36379_ & ~new_n36389_;
  assign new_n36391_ = ~pi0781 & ~new_n36390_;
  assign new_n36392_ = pi0618 & new_n36390_;
  assign new_n36393_ = ~pi0618 & ~new_n36259_;
  assign new_n36394_ = pi1154 & ~new_n36393_;
  assign new_n36395_ = ~new_n36392_ & new_n36394_;
  assign new_n36396_ = ~pi0618 & new_n36390_;
  assign new_n36397_ = pi0618 & ~new_n36259_;
  assign new_n36398_ = ~pi1154 & ~new_n36397_;
  assign new_n36399_ = ~new_n36396_ & new_n36398_;
  assign new_n36400_ = ~new_n36395_ & ~new_n36399_;
  assign new_n36401_ = pi0781 & ~new_n36400_;
  assign new_n36402_ = ~new_n36391_ & ~new_n36401_;
  assign new_n36403_ = ~pi0789 & ~new_n36402_;
  assign new_n36404_ = pi0619 & new_n36402_;
  assign new_n36405_ = ~pi0619 & ~new_n36259_;
  assign new_n36406_ = pi1159 & ~new_n36405_;
  assign new_n36407_ = ~new_n36404_ & new_n36406_;
  assign new_n36408_ = ~pi0619 & new_n36402_;
  assign new_n36409_ = pi0619 & ~new_n36259_;
  assign new_n36410_ = ~pi1159 & ~new_n36409_;
  assign new_n36411_ = ~new_n36408_ & new_n36410_;
  assign new_n36412_ = ~new_n36407_ & ~new_n36411_;
  assign new_n36413_ = pi0789 & ~new_n36412_;
  assign new_n36414_ = ~new_n36403_ & ~new_n36413_;
  assign new_n36415_ = ~new_n17968_ & new_n36414_;
  assign new_n36416_ = ~new_n36260_ & ~new_n36415_;
  assign new_n36417_ = ~new_n20567_ & new_n36416_;
  assign new_n36418_ = ~new_n19279_ & ~new_n36259_;
  assign new_n36419_ = ~pi0222 & ~new_n17168_;
  assign new_n36420_ = pi0661 & pi0680;
  assign new_n36421_ = new_n17168_ & ~new_n36420_;
  assign new_n36422_ = pi0222 & new_n17196_;
  assign new_n36423_ = pi0299 & ~new_n36422_;
  assign new_n36424_ = ~new_n36421_ & new_n36423_;
  assign new_n36425_ = ~new_n36419_ & new_n36424_;
  assign new_n36426_ = ~pi0222 & ~new_n17154_;
  assign new_n36427_ = new_n17154_ & ~new_n36420_;
  assign new_n36428_ = pi0222 & new_n17187_;
  assign new_n36429_ = ~pi0299 & ~new_n36428_;
  assign new_n36430_ = ~new_n36427_ & new_n36429_;
  assign new_n36431_ = ~new_n36426_ & new_n36430_;
  assign new_n36432_ = ~pi0039 & ~new_n36431_;
  assign new_n36433_ = ~new_n36425_ & new_n36432_;
  assign new_n36434_ = pi0661 & ~new_n17489_;
  assign new_n36435_ = ~pi0661 & new_n17296_;
  assign new_n36436_ = ~new_n6181_ & ~new_n16756_;
  assign new_n36437_ = ~pi0662 & new_n17304_;
  assign new_n36438_ = ~new_n36436_ & ~new_n36437_;
  assign new_n36439_ = new_n16629_ & ~new_n36438_;
  assign new_n36440_ = ~new_n36435_ & ~new_n36439_;
  assign new_n36441_ = ~new_n36434_ & new_n36440_;
  assign new_n36442_ = new_n6238_ & new_n36441_;
  assign new_n36443_ = ~pi0661 & ~new_n17320_;
  assign new_n36444_ = pi0680 & new_n17013_;
  assign new_n36445_ = ~new_n16777_ & ~new_n36444_;
  assign new_n36446_ = pi0661 & ~new_n36445_;
  assign new_n36447_ = ~new_n36443_ & ~new_n36446_;
  assign new_n36448_ = ~new_n6238_ & new_n36447_;
  assign new_n36449_ = pi0222 & ~new_n36448_;
  assign new_n36450_ = ~new_n36442_ & new_n36449_;
  assign new_n36451_ = pi0661 & new_n17449_;
  assign new_n36452_ = ~new_n6238_ & new_n36451_;
  assign new_n36453_ = ~new_n17454_ & new_n36420_;
  assign new_n36454_ = new_n6238_ & new_n36453_;
  assign new_n36455_ = pi0224 & ~new_n36454_;
  assign new_n36456_ = ~new_n36452_ & new_n36455_;
  assign new_n36457_ = pi0661 & new_n17474_;
  assign new_n36458_ = ~pi0224 & ~new_n36457_;
  assign new_n36459_ = ~pi0222 & ~new_n36458_;
  assign new_n36460_ = ~new_n36456_ & new_n36459_;
  assign new_n36461_ = ~pi0223 & ~new_n36460_;
  assign new_n36462_ = ~new_n36450_ & new_n36461_;
  assign new_n36463_ = ~pi0661 & ~new_n17292_;
  assign new_n36464_ = ~new_n16694_ & ~new_n17507_;
  assign new_n36465_ = pi0661 & ~new_n36464_;
  assign new_n36466_ = ~new_n36463_ & ~new_n36465_;
  assign new_n36467_ = new_n6238_ & new_n36466_;
  assign new_n36468_ = new_n16629_ & new_n17267_;
  assign new_n36469_ = ~pi0661 & new_n17262_;
  assign new_n36470_ = pi0661 & ~new_n17510_;
  assign new_n36471_ = ~new_n36469_ & ~new_n36470_;
  assign new_n36472_ = ~new_n36468_ & new_n36471_;
  assign new_n36473_ = ~new_n6238_ & new_n36472_;
  assign new_n36474_ = pi0222 & ~new_n36473_;
  assign new_n36475_ = ~new_n36467_ & new_n36474_;
  assign new_n36476_ = ~pi0222 & pi0661;
  assign new_n36477_ = new_n17465_ & new_n36476_;
  assign new_n36478_ = pi0223 & ~new_n36477_;
  assign new_n36479_ = ~new_n36475_ & new_n36478_;
  assign new_n36480_ = ~new_n36462_ & ~new_n36479_;
  assign new_n36481_ = ~pi0299 & ~new_n36480_;
  assign new_n36482_ = new_n6212_ & new_n36441_;
  assign new_n36483_ = ~new_n6212_ & new_n36447_;
  assign new_n36484_ = pi0222 & ~new_n36483_;
  assign new_n36485_ = ~new_n36482_ & new_n36484_;
  assign new_n36486_ = new_n6212_ & ~new_n36453_;
  assign new_n36487_ = ~new_n6212_ & ~new_n36451_;
  assign new_n36488_ = ~pi0222 & ~new_n36487_;
  assign new_n36489_ = ~new_n36486_ & new_n36488_;
  assign new_n36490_ = ~new_n3467_ & ~new_n36489_;
  assign new_n36491_ = ~new_n36485_ & new_n36490_;
  assign new_n36492_ = new_n36346_ & ~new_n36457_;
  assign new_n36493_ = ~pi0215 & ~new_n36492_;
  assign new_n36494_ = ~new_n36491_ & new_n36493_;
  assign new_n36495_ = new_n17478_ & new_n36476_;
  assign new_n36496_ = new_n6212_ & new_n36466_;
  assign new_n36497_ = ~new_n6212_ & new_n36472_;
  assign new_n36498_ = pi0222 & ~new_n36497_;
  assign new_n36499_ = ~new_n36496_ & new_n36498_;
  assign new_n36500_ = ~new_n36495_ & ~new_n36499_;
  assign new_n36501_ = pi0215 & ~new_n36500_;
  assign new_n36502_ = pi0299 & ~new_n36501_;
  assign new_n36503_ = ~new_n36494_ & new_n36502_;
  assign new_n36504_ = ~new_n36481_ & ~new_n36503_;
  assign new_n36505_ = pi0039 & ~new_n36504_;
  assign new_n36506_ = ~new_n36433_ & ~new_n36505_;
  assign new_n36507_ = ~pi0038 & ~new_n36506_;
  assign new_n36508_ = pi0661 & new_n17543_;
  assign new_n36509_ = new_n36370_ & ~new_n36508_;
  assign new_n36510_ = new_n3272_ & ~new_n36509_;
  assign new_n36511_ = ~new_n36507_ & new_n36510_;
  assign new_n36512_ = ~new_n36261_ & ~new_n36511_;
  assign new_n36513_ = ~pi0778 & ~new_n36512_;
  assign new_n36514_ = pi0625 & new_n36512_;
  assign new_n36515_ = ~pi0625 & ~new_n36259_;
  assign new_n36516_ = pi1153 & ~new_n36515_;
  assign new_n36517_ = ~new_n36514_ & new_n36516_;
  assign new_n36518_ = ~pi0625 & new_n36512_;
  assign new_n36519_ = pi0625 & ~new_n36259_;
  assign new_n36520_ = ~pi1153 & ~new_n36519_;
  assign new_n36521_ = ~new_n36518_ & new_n36520_;
  assign new_n36522_ = ~new_n36517_ & ~new_n36521_;
  assign new_n36523_ = pi0778 & ~new_n36522_;
  assign new_n36524_ = ~new_n36513_ & ~new_n36523_;
  assign new_n36525_ = ~new_n17618_ & ~new_n36524_;
  assign new_n36526_ = new_n17618_ & new_n36259_;
  assign new_n36527_ = ~new_n36525_ & ~new_n36526_;
  assign new_n36528_ = ~new_n17655_ & ~new_n36527_;
  assign new_n36529_ = new_n17655_ & new_n36259_;
  assign new_n36530_ = ~new_n36528_ & ~new_n36529_;
  assign new_n36531_ = ~new_n17691_ & new_n36530_;
  assign new_n36532_ = ~new_n17734_ & new_n36531_;
  assign new_n36533_ = ~new_n36418_ & ~new_n36532_;
  assign new_n36534_ = ~pi0628 & ~new_n36533_;
  assign new_n36535_ = pi0628 & ~new_n36259_;
  assign new_n36536_ = new_n17760_ & ~new_n36535_;
  assign new_n36537_ = ~new_n36534_ & new_n36536_;
  assign new_n36538_ = pi0628 & ~new_n36533_;
  assign new_n36539_ = ~pi0628 & ~new_n36259_;
  assign new_n36540_ = new_n17759_ & ~new_n36539_;
  assign new_n36541_ = ~new_n36538_ & new_n36540_;
  assign new_n36542_ = ~new_n36537_ & ~new_n36541_;
  assign new_n36543_ = ~new_n36417_ & new_n36542_;
  assign new_n36544_ = pi0792 & ~new_n36543_;
  assign new_n36545_ = ~pi0680 & new_n36264_;
  assign new_n36546_ = new_n6185_ & new_n16758_;
  assign new_n36547_ = ~new_n16665_ & ~new_n36546_;
  assign new_n36548_ = ~new_n16934_ & new_n36547_;
  assign new_n36549_ = pi0642 & ~new_n36548_;
  assign new_n36550_ = ~pi0603 & new_n36547_;
  assign new_n36551_ = pi0603 & new_n16738_;
  assign new_n36552_ = ~new_n16763_ & ~new_n36551_;
  assign new_n36553_ = ~new_n36550_ & new_n36552_;
  assign new_n36554_ = ~pi0642 & new_n36553_;
  assign new_n36555_ = new_n6179_ & ~new_n36554_;
  assign new_n36556_ = ~new_n36549_ & new_n36555_;
  assign new_n36557_ = new_n16873_ & new_n36548_;
  assign new_n36558_ = new_n16947_ & ~new_n36547_;
  assign new_n36559_ = pi0616 & ~new_n36558_;
  assign new_n36560_ = pi0680 & ~new_n36559_;
  assign new_n36561_ = ~new_n36557_ & new_n36560_;
  assign new_n36562_ = ~new_n36556_ & new_n36561_;
  assign new_n36563_ = pi0661 & ~new_n36562_;
  assign new_n36564_ = ~new_n36545_ & new_n36563_;
  assign new_n36565_ = ~pi0661 & pi0681;
  assign new_n36566_ = ~new_n36264_ & new_n36565_;
  assign new_n36567_ = ~new_n36272_ & ~new_n36566_;
  assign new_n36568_ = ~new_n36564_ & new_n36567_;
  assign new_n36569_ = ~new_n6212_ & ~new_n36568_;
  assign new_n36570_ = pi0616 & ~new_n17021_;
  assign new_n36571_ = pi0680 & ~new_n36570_;
  assign new_n36572_ = ~new_n16748_ & new_n36571_;
  assign new_n36573_ = ~pi0680 & new_n36276_;
  assign new_n36574_ = pi0661 & ~new_n36573_;
  assign new_n36575_ = ~new_n36572_ & new_n36574_;
  assign new_n36576_ = ~new_n36276_ & new_n36565_;
  assign new_n36577_ = ~new_n36282_ & ~new_n36576_;
  assign new_n36578_ = ~new_n36575_ & new_n36577_;
  assign new_n36579_ = new_n6212_ & ~new_n36578_;
  assign new_n36580_ = pi0222 & ~new_n36579_;
  assign new_n36581_ = ~new_n36569_ & new_n36580_;
  assign new_n36582_ = pi0616 & new_n16935_;
  assign new_n36583_ = pi0680 & ~new_n36582_;
  assign new_n36584_ = ~new_n16834_ & new_n36583_;
  assign new_n36585_ = ~pi0680 & new_n36287_;
  assign new_n36586_ = pi0661 & ~new_n36585_;
  assign new_n36587_ = ~new_n36584_ & new_n36586_;
  assign new_n36588_ = ~new_n36287_ & new_n36565_;
  assign new_n36589_ = ~new_n36293_ & ~new_n36588_;
  assign new_n36590_ = ~new_n36587_ & new_n36589_;
  assign new_n36591_ = ~new_n6212_ & new_n36590_;
  assign new_n36592_ = pi0616 & ~new_n16948_;
  assign new_n36593_ = pi0680 & ~new_n16858_;
  assign new_n36594_ = ~new_n36592_ & new_n36593_;
  assign new_n36595_ = ~pi0680 & new_n36302_;
  assign new_n36596_ = pi0661 & ~new_n36595_;
  assign new_n36597_ = ~new_n36594_ & new_n36596_;
  assign new_n36598_ = new_n16951_ & new_n36290_;
  assign new_n36599_ = ~new_n6181_ & new_n36302_;
  assign new_n36600_ = new_n16629_ & ~new_n36599_;
  assign new_n36601_ = ~new_n36598_ & new_n36600_;
  assign new_n36602_ = ~new_n36302_ & new_n36565_;
  assign new_n36603_ = ~new_n36601_ & ~new_n36602_;
  assign new_n36604_ = ~new_n36597_ & new_n36603_;
  assign new_n36605_ = new_n6212_ & new_n36604_;
  assign new_n36606_ = ~pi0222 & ~new_n36605_;
  assign new_n36607_ = ~new_n36591_ & new_n36606_;
  assign new_n36608_ = ~new_n36581_ & ~new_n36607_;
  assign new_n36609_ = ~new_n3467_ & ~new_n36608_;
  assign new_n36610_ = ~new_n36267_ & ~new_n36420_;
  assign new_n36611_ = ~pi0616 & ~new_n16843_;
  assign new_n36612_ = ~new_n36592_ & ~new_n36611_;
  assign new_n36613_ = ~new_n36610_ & new_n36612_;
  assign new_n36614_ = new_n36346_ & ~new_n36613_;
  assign new_n36615_ = ~pi0215 & ~new_n36614_;
  assign new_n36616_ = ~new_n36609_ & new_n36615_;
  assign new_n36617_ = ~pi0680 & new_n36317_;
  assign new_n36618_ = ~new_n16709_ & new_n16947_;
  assign new_n36619_ = pi0616 & ~new_n36618_;
  assign new_n36620_ = pi0680 & ~new_n36619_;
  assign new_n36621_ = new_n16713_ & new_n36620_;
  assign new_n36622_ = pi0661 & ~new_n36621_;
  assign new_n36623_ = ~new_n36617_ & new_n36622_;
  assign new_n36624_ = ~new_n36317_ & new_n36565_;
  assign new_n36625_ = ~new_n36322_ & ~new_n36624_;
  assign new_n36626_ = ~new_n36623_ & new_n36625_;
  assign new_n36627_ = ~new_n6212_ & ~new_n36626_;
  assign new_n36628_ = ~new_n16680_ & new_n36571_;
  assign new_n36629_ = ~pi0680 & new_n36308_;
  assign new_n36630_ = pi0661 & ~new_n36629_;
  assign new_n36631_ = ~new_n36628_ & new_n36630_;
  assign new_n36632_ = ~new_n36308_ & new_n36565_;
  assign new_n36633_ = ~new_n36313_ & ~new_n36632_;
  assign new_n36634_ = ~new_n36631_ & new_n36633_;
  assign new_n36635_ = new_n6212_ & ~new_n36634_;
  assign new_n36636_ = pi0222 & ~new_n36635_;
  assign new_n36637_ = ~new_n36627_ & new_n36636_;
  assign new_n36638_ = ~new_n16708_ & ~new_n16985_;
  assign new_n36639_ = pi0616 & new_n36638_;
  assign new_n36640_ = pi0680 & ~new_n36639_;
  assign new_n36641_ = new_n16883_ & new_n36640_;
  assign new_n36642_ = pi0616 & new_n16708_;
  assign new_n36643_ = ~pi0680 & new_n36642_;
  assign new_n36644_ = pi0661 & ~new_n36643_;
  assign new_n36645_ = ~new_n36641_ & new_n36644_;
  assign new_n36646_ = ~pi0661 & ~new_n36642_;
  assign new_n36647_ = ~new_n16660_ & new_n36302_;
  assign new_n36648_ = new_n6183_ & ~new_n36647_;
  assign new_n36649_ = ~new_n36646_ & ~new_n36648_;
  assign new_n36650_ = ~new_n36645_ & new_n36649_;
  assign new_n36651_ = ~new_n6212_ & new_n36650_;
  assign new_n36652_ = new_n16894_ & new_n36420_;
  assign new_n36653_ = ~new_n36328_ & ~new_n36652_;
  assign new_n36654_ = new_n6212_ & ~new_n36653_;
  assign new_n36655_ = ~pi0222 & ~new_n36654_;
  assign new_n36656_ = ~new_n36651_ & new_n36655_;
  assign new_n36657_ = pi0215 & ~new_n36656_;
  assign new_n36658_ = ~new_n36637_ & new_n36657_;
  assign new_n36659_ = pi0299 & ~new_n36658_;
  assign new_n36660_ = ~new_n36616_ & new_n36659_;
  assign new_n36661_ = new_n36420_ & ~new_n36612_;
  assign new_n36662_ = ~new_n36302_ & ~new_n36420_;
  assign new_n36663_ = ~pi0222 & ~new_n36662_;
  assign new_n36664_ = ~new_n36661_ & new_n36663_;
  assign new_n36665_ = ~new_n3313_ & ~new_n36664_;
  assign new_n36666_ = ~new_n6238_ & new_n36590_;
  assign new_n36667_ = new_n6238_ & new_n36604_;
  assign new_n36668_ = pi0224 & ~new_n36667_;
  assign new_n36669_ = ~new_n36666_ & new_n36668_;
  assign new_n36670_ = ~new_n36665_ & ~new_n36669_;
  assign new_n36671_ = ~new_n6238_ & new_n36568_;
  assign new_n36672_ = new_n6238_ & new_n36578_;
  assign new_n36673_ = pi0222 & ~new_n36672_;
  assign new_n36674_ = ~new_n36671_ & new_n36673_;
  assign new_n36675_ = ~new_n36670_ & ~new_n36674_;
  assign new_n36676_ = ~pi0223 & ~new_n36675_;
  assign new_n36677_ = ~new_n6238_ & ~new_n36626_;
  assign new_n36678_ = new_n6238_ & ~new_n36634_;
  assign new_n36679_ = pi0222 & ~new_n36678_;
  assign new_n36680_ = ~new_n36677_ & new_n36679_;
  assign new_n36681_ = ~new_n6238_ & new_n36650_;
  assign new_n36682_ = new_n6238_ & ~new_n36653_;
  assign new_n36683_ = ~pi0222 & ~new_n36682_;
  assign new_n36684_ = ~new_n36681_ & new_n36683_;
  assign new_n36685_ = pi0223 & ~new_n36684_;
  assign new_n36686_ = ~new_n36680_ & new_n36685_;
  assign new_n36687_ = ~pi0299 & ~new_n36686_;
  assign new_n36688_ = ~new_n36676_ & new_n36687_;
  assign new_n36689_ = pi0039 & ~new_n36688_;
  assign new_n36690_ = ~new_n36660_ & new_n36689_;
  assign new_n36691_ = new_n17175_ & ~new_n36420_;
  assign new_n36692_ = ~pi0616 & new_n17213_;
  assign new_n36693_ = ~pi0603 & ~new_n17196_;
  assign new_n36694_ = ~new_n16762_ & ~new_n17173_;
  assign new_n36695_ = ~new_n36693_ & new_n36694_;
  assign new_n36696_ = ~new_n36692_ & ~new_n36695_;
  assign new_n36697_ = ~new_n36691_ & new_n36696_;
  assign new_n36698_ = pi0222 & ~new_n36697_;
  assign new_n36699_ = pi0661 & new_n17176_;
  assign new_n36700_ = pi0616 & new_n17213_;
  assign new_n36701_ = ~pi0222 & ~new_n36700_;
  assign new_n36702_ = ~new_n36699_ & new_n36701_;
  assign new_n36703_ = ~new_n36698_ & ~new_n36702_;
  assign new_n36704_ = pi0299 & ~new_n36703_;
  assign new_n36705_ = pi0661 & new_n17164_;
  assign new_n36706_ = pi0616 & new_n17208_;
  assign new_n36707_ = ~pi0222 & ~new_n36706_;
  assign new_n36708_ = ~new_n36705_ & new_n36707_;
  assign new_n36709_ = new_n17163_ & ~new_n36420_;
  assign new_n36710_ = ~pi0616 & new_n17208_;
  assign new_n36711_ = ~pi0603 & ~new_n17187_;
  assign new_n36712_ = ~new_n16762_ & ~new_n17161_;
  assign new_n36713_ = ~new_n36711_ & new_n36712_;
  assign new_n36714_ = ~new_n36710_ & ~new_n36713_;
  assign new_n36715_ = ~new_n36709_ & new_n36714_;
  assign new_n36716_ = pi0222 & ~new_n36715_;
  assign new_n36717_ = ~new_n36708_ & ~new_n36716_;
  assign new_n36718_ = ~pi0299 & ~new_n36717_;
  assign new_n36719_ = ~pi0039 & ~new_n36718_;
  assign new_n36720_ = ~new_n36704_ & new_n36719_;
  assign new_n36721_ = ~pi0038 & ~new_n36720_;
  assign new_n36722_ = ~new_n36690_ & new_n36721_;
  assign new_n36723_ = new_n16647_ & new_n16947_;
  assign new_n36724_ = ~pi0222 & ~pi0616;
  assign new_n36725_ = ~pi0039 & pi0616;
  assign new_n36726_ = new_n36420_ & new_n36725_;
  assign new_n36727_ = ~new_n36724_ & ~new_n36726_;
  assign new_n36728_ = new_n36723_ & ~new_n36727_;
  assign new_n36729_ = ~pi0616 & ~new_n16790_;
  assign new_n36730_ = ~new_n36610_ & ~new_n36729_;
  assign new_n36731_ = new_n17431_ & new_n36730_;
  assign new_n36732_ = ~new_n36369_ & ~new_n36731_;
  assign new_n36733_ = ~new_n36728_ & ~new_n36732_;
  assign new_n36734_ = pi0038 & ~new_n36733_;
  assign new_n36735_ = new_n3272_ & ~new_n36734_;
  assign new_n36736_ = ~new_n36722_ & new_n36735_;
  assign new_n36737_ = ~new_n36261_ & ~new_n36736_;
  assign new_n36738_ = ~pi0625 & new_n36737_;
  assign new_n36739_ = pi0625 & new_n36375_;
  assign new_n36740_ = ~pi1153 & ~new_n36739_;
  assign new_n36741_ = ~new_n36738_ & new_n36740_;
  assign new_n36742_ = ~pi0608 & ~new_n36517_;
  assign new_n36743_ = ~new_n36741_ & new_n36742_;
  assign new_n36744_ = pi0625 & new_n36737_;
  assign new_n36745_ = ~pi0625 & new_n36375_;
  assign new_n36746_ = pi1153 & ~new_n36745_;
  assign new_n36747_ = ~new_n36744_ & new_n36746_;
  assign new_n36748_ = pi0608 & ~new_n36521_;
  assign new_n36749_ = ~new_n36747_ & new_n36748_;
  assign new_n36750_ = ~new_n36743_ & ~new_n36749_;
  assign new_n36751_ = pi0778 & ~new_n36750_;
  assign new_n36752_ = ~pi0778 & new_n36737_;
  assign new_n36753_ = ~new_n36751_ & ~new_n36752_;
  assign new_n36754_ = ~pi0609 & ~new_n36753_;
  assign new_n36755_ = pi0609 & new_n36524_;
  assign new_n36756_ = ~pi1155 & ~new_n36755_;
  assign new_n36757_ = ~new_n36754_ & new_n36756_;
  assign new_n36758_ = ~pi0660 & ~new_n36383_;
  assign new_n36759_ = ~new_n36757_ & new_n36758_;
  assign new_n36760_ = pi0609 & ~new_n36753_;
  assign new_n36761_ = ~pi0609 & new_n36524_;
  assign new_n36762_ = pi1155 & ~new_n36761_;
  assign new_n36763_ = ~new_n36760_ & new_n36762_;
  assign new_n36764_ = pi0660 & ~new_n36387_;
  assign new_n36765_ = ~new_n36763_ & new_n36764_;
  assign new_n36766_ = ~new_n36759_ & ~new_n36765_;
  assign new_n36767_ = pi0785 & ~new_n36766_;
  assign new_n36768_ = ~pi0785 & ~new_n36753_;
  assign new_n36769_ = ~new_n36767_ & ~new_n36768_;
  assign new_n36770_ = ~pi0618 & ~new_n36769_;
  assign new_n36771_ = pi0618 & new_n36527_;
  assign new_n36772_ = ~pi1154 & ~new_n36771_;
  assign new_n36773_ = ~new_n36770_ & new_n36772_;
  assign new_n36774_ = ~pi0627 & ~new_n36395_;
  assign new_n36775_ = ~new_n36773_ & new_n36774_;
  assign new_n36776_ = pi0618 & ~new_n36769_;
  assign new_n36777_ = ~pi0618 & new_n36527_;
  assign new_n36778_ = pi1154 & ~new_n36777_;
  assign new_n36779_ = ~new_n36776_ & new_n36778_;
  assign new_n36780_ = pi0627 & ~new_n36399_;
  assign new_n36781_ = ~new_n36779_ & new_n36780_;
  assign new_n36782_ = ~new_n36775_ & ~new_n36781_;
  assign new_n36783_ = pi0781 & ~new_n36782_;
  assign new_n36784_ = ~pi0781 & ~new_n36769_;
  assign new_n36785_ = ~new_n36783_ & ~new_n36784_;
  assign new_n36786_ = pi0619 & ~new_n36785_;
  assign new_n36787_ = ~pi0619 & new_n36530_;
  assign new_n36788_ = pi1159 & ~new_n36787_;
  assign new_n36789_ = ~new_n36786_ & new_n36788_;
  assign new_n36790_ = pi0648 & ~new_n36411_;
  assign new_n36791_ = ~new_n36789_ & new_n36790_;
  assign new_n36792_ = ~pi0619 & ~new_n36785_;
  assign new_n36793_ = pi0619 & new_n36530_;
  assign new_n36794_ = ~pi1159 & ~new_n36793_;
  assign new_n36795_ = ~new_n36792_ & new_n36794_;
  assign new_n36796_ = ~pi0648 & ~new_n36407_;
  assign new_n36797_ = ~new_n36795_ & new_n36796_;
  assign new_n36798_ = pi0789 & ~new_n36797_;
  assign new_n36799_ = ~new_n36791_ & new_n36798_;
  assign new_n36800_ = ~pi0789 & new_n36785_;
  assign new_n36801_ = pi0626 & new_n36414_;
  assign new_n36802_ = ~pi0626 & ~new_n36259_;
  assign new_n36803_ = new_n17731_ & ~new_n36802_;
  assign new_n36804_ = ~new_n36801_ & new_n36803_;
  assign new_n36805_ = ~pi0626 & new_n36414_;
  assign new_n36806_ = pi0626 & ~new_n36259_;
  assign new_n36807_ = new_n17732_ & ~new_n36806_;
  assign new_n36808_ = ~new_n36805_ & new_n36807_;
  assign new_n36809_ = new_n17691_ & ~new_n36259_;
  assign new_n36810_ = new_n17856_ & ~new_n36809_;
  assign new_n36811_ = ~new_n36531_ & new_n36810_;
  assign new_n36812_ = ~new_n36808_ & ~new_n36811_;
  assign new_n36813_ = ~new_n36804_ & new_n36812_;
  assign new_n36814_ = pi0788 & ~new_n36813_;
  assign new_n36815_ = ~new_n36800_ & ~new_n36814_;
  assign new_n36816_ = ~new_n36799_ & new_n36815_;
  assign new_n36817_ = ~new_n17969_ & new_n36813_;
  assign new_n36818_ = ~new_n20364_ & ~new_n36817_;
  assign new_n36819_ = ~new_n36816_ & new_n36818_;
  assign new_n36820_ = ~new_n36544_ & ~new_n36819_;
  assign new_n36821_ = ~new_n20360_ & ~new_n36820_;
  assign new_n36822_ = ~new_n17762_ & new_n36416_;
  assign new_n36823_ = new_n17762_ & new_n36259_;
  assign new_n36824_ = ~new_n36822_ & ~new_n36823_;
  assign new_n36825_ = ~new_n20556_ & ~new_n36824_;
  assign new_n36826_ = ~new_n19311_ & ~new_n36533_;
  assign new_n36827_ = new_n18010_ & ~new_n36259_;
  assign new_n36828_ = ~new_n36826_ & ~new_n36827_;
  assign new_n36829_ = pi0647 & ~new_n36828_;
  assign new_n36830_ = ~pi0647 & ~new_n36259_;
  assign new_n36831_ = pi1157 & ~new_n36830_;
  assign new_n36832_ = ~new_n36829_ & new_n36831_;
  assign new_n36833_ = ~pi0630 & new_n36832_;
  assign new_n36834_ = ~pi0647 & ~new_n36828_;
  assign new_n36835_ = pi0647 & ~new_n36259_;
  assign new_n36836_ = ~pi1157 & ~new_n36835_;
  assign new_n36837_ = ~new_n36834_ & new_n36836_;
  assign new_n36838_ = pi0630 & new_n36837_;
  assign new_n36839_ = ~new_n36833_ & ~new_n36838_;
  assign new_n36840_ = ~new_n36825_ & new_n36839_;
  assign new_n36841_ = pi0787 & ~new_n36840_;
  assign new_n36842_ = ~new_n36821_ & ~new_n36841_;
  assign new_n36843_ = pi0644 & new_n36842_;
  assign new_n36844_ = ~pi0787 & new_n36828_;
  assign new_n36845_ = ~new_n36832_ & ~new_n36837_;
  assign new_n36846_ = pi0787 & ~new_n36845_;
  assign new_n36847_ = ~new_n36844_ & ~new_n36846_;
  assign new_n36848_ = ~pi0644 & new_n36847_;
  assign new_n36849_ = pi0715 & ~new_n36848_;
  assign new_n36850_ = ~new_n36843_ & new_n36849_;
  assign new_n36851_ = new_n17804_ & ~new_n36259_;
  assign new_n36852_ = ~new_n17804_ & new_n36824_;
  assign new_n36853_ = ~new_n36851_ & ~new_n36852_;
  assign new_n36854_ = pi0644 & ~new_n36853_;
  assign new_n36855_ = ~pi0644 & ~new_n36259_;
  assign new_n36856_ = ~pi0715 & ~new_n36855_;
  assign new_n36857_ = ~new_n36854_ & new_n36856_;
  assign new_n36858_ = pi1160 & ~new_n36857_;
  assign new_n36859_ = ~new_n36850_ & new_n36858_;
  assign new_n36860_ = ~pi0644 & new_n36842_;
  assign new_n36861_ = pi0644 & new_n36847_;
  assign new_n36862_ = ~pi0715 & ~new_n36861_;
  assign new_n36863_ = ~new_n36860_ & new_n36862_;
  assign new_n36864_ = ~pi0644 & ~new_n36853_;
  assign new_n36865_ = pi0644 & ~new_n36259_;
  assign new_n36866_ = pi0715 & ~new_n36865_;
  assign new_n36867_ = ~new_n36864_ & new_n36866_;
  assign new_n36868_ = ~pi1160 & ~new_n36867_;
  assign new_n36869_ = ~new_n36863_ & new_n36868_;
  assign new_n36870_ = ~new_n36859_ & ~new_n36869_;
  assign new_n36871_ = pi0790 & ~new_n36870_;
  assign new_n36872_ = ~pi0790 & new_n36842_;
  assign new_n36873_ = ~new_n36871_ & ~new_n36872_;
  assign new_n36874_ = ~po1038 & ~new_n36873_;
  assign new_n36875_ = ~pi0222 & po1038;
  assign po0379 = ~new_n36874_ & ~new_n36875_;
  assign new_n36877_ = ~pi0299 & ~new_n17294_;
  assign new_n36878_ = pi0039 & ~new_n36877_;
  assign new_n36879_ = ~new_n17346_ & new_n36878_;
  assign new_n36880_ = new_n14865_ & ~new_n18106_;
  assign new_n36881_ = ~new_n36879_ & new_n36880_;
  assign new_n36882_ = new_n18873_ & ~new_n36881_;
  assign new_n36883_ = pi0223 & ~new_n36882_;
  assign new_n36884_ = new_n17968_ & ~new_n36883_;
  assign new_n36885_ = new_n17590_ & ~new_n36883_;
  assign new_n36886_ = pi0223 & ~new_n3272_;
  assign new_n36887_ = pi0642 & new_n16639_;
  assign new_n36888_ = new_n35877_ & ~new_n36887_;
  assign new_n36889_ = pi0642 & ~new_n16842_;
  assign new_n36890_ = new_n6179_ & ~new_n36889_;
  assign new_n36891_ = ~new_n16751_ & new_n36890_;
  assign new_n36892_ = ~new_n36888_ & ~new_n36891_;
  assign new_n36893_ = pi0681 & new_n36892_;
  assign new_n36894_ = ~new_n6182_ & ~new_n36892_;
  assign new_n36895_ = ~new_n17352_ & ~new_n35874_;
  assign new_n36896_ = new_n6182_ & ~new_n36895_;
  assign new_n36897_ = ~pi0681 & ~new_n36896_;
  assign new_n36898_ = ~new_n36894_ & new_n36897_;
  assign new_n36899_ = new_n6212_ & ~new_n36898_;
  assign new_n36900_ = ~new_n36893_ & new_n36899_;
  assign new_n36901_ = pi0642 & ~new_n16822_;
  assign new_n36902_ = ~pi0642 & ~new_n16774_;
  assign new_n36903_ = ~new_n36901_ & ~new_n36902_;
  assign new_n36904_ = pi0681 & ~new_n36903_;
  assign new_n36905_ = ~new_n6182_ & new_n36903_;
  assign new_n36906_ = new_n17317_ & ~new_n36887_;
  assign new_n36907_ = ~pi0681 & ~new_n36906_;
  assign new_n36908_ = ~new_n36905_ & new_n36907_;
  assign new_n36909_ = ~new_n6212_ & ~new_n36908_;
  assign new_n36910_ = ~new_n36904_ & new_n36909_;
  assign new_n36911_ = pi0223 & ~new_n36910_;
  assign new_n36912_ = ~new_n36900_ & new_n36911_;
  assign new_n36913_ = ~new_n16771_ & new_n36887_;
  assign new_n36914_ = pi0681 & ~new_n36913_;
  assign new_n36915_ = ~new_n6182_ & new_n36913_;
  assign new_n36916_ = pi0642 & new_n6182_;
  assign new_n36917_ = new_n16780_ & new_n36916_;
  assign new_n36918_ = ~pi0681 & ~new_n36917_;
  assign new_n36919_ = ~new_n36915_ & new_n36918_;
  assign new_n36920_ = ~new_n36914_ & ~new_n36919_;
  assign new_n36921_ = ~new_n20899_ & new_n36920_;
  assign new_n36922_ = pi0642 & new_n16661_;
  assign new_n36923_ = ~new_n6182_ & new_n36922_;
  assign new_n36924_ = ~pi0681 & ~new_n36923_;
  assign new_n36925_ = new_n16951_ & new_n36916_;
  assign new_n36926_ = new_n36924_ & ~new_n36925_;
  assign new_n36927_ = pi0681 & ~new_n36922_;
  assign new_n36928_ = ~new_n36926_ & ~new_n36927_;
  assign new_n36929_ = new_n20899_ & new_n36928_;
  assign new_n36930_ = ~pi0947 & ~new_n36929_;
  assign new_n36931_ = ~new_n36921_ & new_n36930_;
  assign new_n36932_ = pi0947 & ~new_n36920_;
  assign new_n36933_ = ~pi0223 & ~new_n36932_;
  assign new_n36934_ = ~new_n36931_ & new_n36933_;
  assign new_n36935_ = ~new_n3467_ & ~new_n36934_;
  assign new_n36936_ = ~new_n36912_ & new_n36935_;
  assign new_n36937_ = pi0223 & ~new_n16636_;
  assign new_n36938_ = new_n3467_ & ~new_n36937_;
  assign new_n36939_ = ~new_n36922_ & new_n36938_;
  assign new_n36940_ = ~pi0215 & ~new_n36939_;
  assign new_n36941_ = ~new_n36936_ & new_n36940_;
  assign new_n36942_ = new_n16669_ & new_n36916_;
  assign new_n36943_ = new_n36924_ & ~new_n36942_;
  assign new_n36944_ = pi0642 & ~new_n16869_;
  assign new_n36945_ = new_n6182_ & ~new_n36944_;
  assign new_n36946_ = ~new_n16660_ & new_n36945_;
  assign new_n36947_ = ~pi0681 & ~new_n36946_;
  assign new_n36948_ = new_n16701_ & new_n36947_;
  assign new_n36949_ = ~new_n36943_ & ~new_n36948_;
  assign new_n36950_ = pi0642 & new_n16708_;
  assign new_n36951_ = pi0681 & ~new_n36950_;
  assign new_n36952_ = new_n36949_ & ~new_n36951_;
  assign new_n36953_ = ~new_n20899_ & new_n36952_;
  assign new_n36954_ = new_n6212_ & ~new_n36943_;
  assign new_n36955_ = new_n36922_ & new_n36954_;
  assign new_n36956_ = ~pi0947 & ~new_n36955_;
  assign new_n36957_ = ~new_n36953_ & new_n36956_;
  assign new_n36958_ = pi0947 & ~new_n36952_;
  assign new_n36959_ = ~pi0223 & ~new_n36958_;
  assign new_n36960_ = ~new_n36957_ & new_n36959_;
  assign new_n36961_ = new_n36308_ & ~new_n36889_;
  assign new_n36962_ = ~new_n36888_ & ~new_n36961_;
  assign new_n36963_ = pi0681 & new_n36962_;
  assign new_n36964_ = ~new_n6182_ & ~new_n36962_;
  assign new_n36965_ = new_n16647_ & ~new_n36887_;
  assign new_n36966_ = new_n6182_ & new_n36965_;
  assign new_n36967_ = new_n16687_ & new_n36966_;
  assign new_n36968_ = ~pi0681 & ~new_n36967_;
  assign new_n36969_ = ~new_n36964_ & new_n36968_;
  assign new_n36970_ = ~new_n36963_ & ~new_n36969_;
  assign new_n36971_ = new_n6212_ & new_n36970_;
  assign new_n36972_ = ~pi0642 & ~new_n16703_;
  assign new_n36973_ = pi0642 & ~new_n16870_;
  assign new_n36974_ = ~new_n36972_ & ~new_n36973_;
  assign new_n36975_ = ~new_n6182_ & new_n36974_;
  assign new_n36976_ = new_n36947_ & ~new_n36975_;
  assign new_n36977_ = pi0681 & ~new_n36974_;
  assign new_n36978_ = ~new_n36976_ & ~new_n36977_;
  assign new_n36979_ = ~new_n6212_ & new_n36978_;
  assign new_n36980_ = pi0223 & ~new_n36979_;
  assign new_n36981_ = ~new_n36971_ & new_n36980_;
  assign new_n36982_ = ~new_n36960_ & ~new_n36981_;
  assign new_n36983_ = pi0215 & ~new_n36982_;
  assign new_n36984_ = pi0299 & ~new_n36983_;
  assign new_n36985_ = ~new_n36941_ & new_n36984_;
  assign new_n36986_ = ~new_n6238_ & new_n36920_;
  assign new_n36987_ = new_n6238_ & new_n36928_;
  assign new_n36988_ = ~new_n3057_ & ~new_n36987_;
  assign new_n36989_ = ~new_n36986_ & new_n36988_;
  assign new_n36990_ = new_n3057_ & ~new_n36922_;
  assign new_n36991_ = ~pi0223 & ~new_n36990_;
  assign new_n36992_ = ~new_n36989_ & new_n36991_;
  assign new_n36993_ = new_n6238_ & new_n36970_;
  assign new_n36994_ = ~new_n6238_ & new_n36978_;
  assign new_n36995_ = pi0223 & ~new_n36994_;
  assign new_n36996_ = ~new_n36993_ & new_n36995_;
  assign new_n36997_ = ~pi0299 & ~new_n36996_;
  assign new_n36998_ = ~new_n36992_ & new_n36997_;
  assign new_n36999_ = pi0039 & ~new_n36998_;
  assign new_n37000_ = ~new_n36985_ & new_n36999_;
  assign new_n37001_ = ~pi0223 & pi0642;
  assign new_n37002_ = new_n17208_ & new_n37001_;
  assign new_n37003_ = ~pi0299 & ~new_n37002_;
  assign new_n37004_ = ~pi0642 & new_n17208_;
  assign new_n37005_ = pi0223 & ~new_n37004_;
  assign new_n37006_ = new_n17224_ & new_n37005_;
  assign new_n37007_ = new_n37003_ & ~new_n37006_;
  assign new_n37008_ = new_n17213_ & new_n37001_;
  assign new_n37009_ = pi0299 & ~new_n37008_;
  assign new_n37010_ = new_n6178_ & new_n17212_;
  assign new_n37011_ = pi0223 & ~new_n17221_;
  assign new_n37012_ = ~new_n37010_ & new_n37011_;
  assign new_n37013_ = new_n37009_ & ~new_n37012_;
  assign new_n37014_ = ~pi0039 & ~new_n37013_;
  assign new_n37015_ = ~new_n37007_ & new_n37014_;
  assign new_n37016_ = ~pi0038 & ~new_n37015_;
  assign new_n37017_ = ~new_n37000_ & new_n37016_;
  assign new_n37018_ = pi0039 & pi0223;
  assign new_n37019_ = pi0038 & ~new_n37018_;
  assign new_n37020_ = ~pi0223 & ~new_n16647_;
  assign new_n37021_ = ~pi0039 & ~new_n37020_;
  assign new_n37022_ = ~new_n36965_ & new_n37021_;
  assign new_n37023_ = new_n37019_ & ~new_n37022_;
  assign new_n37024_ = new_n3272_ & ~new_n37023_;
  assign new_n37025_ = ~new_n37017_ & new_n37024_;
  assign new_n37026_ = ~new_n36886_ & ~new_n37025_;
  assign new_n37027_ = ~new_n17590_ & new_n37026_;
  assign new_n37028_ = ~new_n36885_ & ~new_n37027_;
  assign new_n37029_ = ~pi0785 & new_n37028_;
  assign new_n37030_ = pi0609 & ~new_n37028_;
  assign new_n37031_ = ~pi0609 & ~new_n36883_;
  assign new_n37032_ = pi1155 & ~new_n37031_;
  assign new_n37033_ = ~new_n37030_ & new_n37032_;
  assign new_n37034_ = ~pi0609 & ~new_n37028_;
  assign new_n37035_ = pi0609 & ~new_n36883_;
  assign new_n37036_ = ~pi1155 & ~new_n37035_;
  assign new_n37037_ = ~new_n37034_ & new_n37036_;
  assign new_n37038_ = ~new_n37033_ & ~new_n37037_;
  assign new_n37039_ = pi0785 & ~new_n37038_;
  assign new_n37040_ = ~new_n37029_ & ~new_n37039_;
  assign new_n37041_ = ~pi0781 & ~new_n37040_;
  assign new_n37042_ = pi0618 & new_n37040_;
  assign new_n37043_ = ~pi0618 & ~new_n36883_;
  assign new_n37044_ = pi1154 & ~new_n37043_;
  assign new_n37045_ = ~new_n37042_ & new_n37044_;
  assign new_n37046_ = ~pi0618 & new_n37040_;
  assign new_n37047_ = pi0618 & ~new_n36883_;
  assign new_n37048_ = ~pi1154 & ~new_n37047_;
  assign new_n37049_ = ~new_n37046_ & new_n37048_;
  assign new_n37050_ = ~new_n37045_ & ~new_n37049_;
  assign new_n37051_ = pi0781 & ~new_n37050_;
  assign new_n37052_ = ~new_n37041_ & ~new_n37051_;
  assign new_n37053_ = ~pi0789 & ~new_n37052_;
  assign new_n37054_ = pi0619 & new_n37052_;
  assign new_n37055_ = ~pi0619 & ~new_n36883_;
  assign new_n37056_ = pi1159 & ~new_n37055_;
  assign new_n37057_ = ~new_n37054_ & new_n37056_;
  assign new_n37058_ = ~pi0619 & new_n37052_;
  assign new_n37059_ = pi0619 & ~new_n36883_;
  assign new_n37060_ = ~pi1159 & ~new_n37059_;
  assign new_n37061_ = ~new_n37058_ & new_n37060_;
  assign new_n37062_ = ~new_n37057_ & ~new_n37061_;
  assign new_n37063_ = pi0789 & ~new_n37062_;
  assign new_n37064_ = ~new_n37053_ & ~new_n37063_;
  assign new_n37065_ = ~new_n17968_ & new_n37064_;
  assign new_n37066_ = ~new_n36884_ & ~new_n37065_;
  assign new_n37067_ = ~new_n17762_ & new_n37066_;
  assign new_n37068_ = new_n17762_ & new_n36883_;
  assign new_n37069_ = ~new_n37067_ & ~new_n37068_;
  assign new_n37070_ = ~new_n20556_ & ~new_n37069_;
  assign new_n37071_ = ~new_n19279_ & ~new_n36883_;
  assign new_n37072_ = new_n17618_ & ~new_n36883_;
  assign new_n37073_ = ~pi0223 & ~new_n17168_;
  assign new_n37074_ = pi0680 & pi0681;
  assign new_n37075_ = new_n17168_ & ~new_n37074_;
  assign new_n37076_ = pi0223 & new_n17196_;
  assign new_n37077_ = pi0299 & ~new_n37076_;
  assign new_n37078_ = ~new_n37075_ & new_n37077_;
  assign new_n37079_ = ~new_n37073_ & new_n37078_;
  assign new_n37080_ = ~pi0223 & ~new_n17154_;
  assign new_n37081_ = new_n17154_ & ~new_n37074_;
  assign new_n37082_ = pi0223 & new_n17187_;
  assign new_n37083_ = ~pi0299 & ~new_n37082_;
  assign new_n37084_ = ~new_n37081_ & new_n37083_;
  assign new_n37085_ = ~new_n37080_ & new_n37084_;
  assign new_n37086_ = ~pi0039 & ~new_n37085_;
  assign new_n37087_ = ~new_n37079_ & new_n37086_;
  assign new_n37088_ = pi0681 & new_n17474_;
  assign new_n37089_ = new_n36938_ & ~new_n37088_;
  assign new_n37090_ = pi0681 & ~new_n17489_;
  assign new_n37091_ = new_n6212_ & ~new_n17312_;
  assign new_n37092_ = ~new_n37090_ & new_n37091_;
  assign new_n37093_ = pi0681 & ~new_n36445_;
  assign new_n37094_ = ~new_n6212_ & ~new_n17319_;
  assign new_n37095_ = ~new_n37093_ & new_n37094_;
  assign new_n37096_ = pi0223 & ~new_n37095_;
  assign new_n37097_ = ~new_n37092_ & new_n37096_;
  assign new_n37098_ = ~new_n17454_ & new_n37074_;
  assign new_n37099_ = new_n6212_ & ~new_n37098_;
  assign new_n37100_ = pi0681 & new_n17449_;
  assign new_n37101_ = ~new_n6212_ & ~new_n37100_;
  assign new_n37102_ = ~pi0223 & ~new_n37101_;
  assign new_n37103_ = ~new_n37099_ & new_n37102_;
  assign new_n37104_ = ~new_n3467_ & ~new_n37103_;
  assign new_n37105_ = ~new_n37097_ & new_n37104_;
  assign new_n37106_ = ~new_n37089_ & ~new_n37105_;
  assign new_n37107_ = ~pi0215 & ~new_n37106_;
  assign new_n37108_ = pi0681 & ~new_n17510_;
  assign new_n37109_ = ~new_n17271_ & ~new_n37108_;
  assign new_n37110_ = ~new_n6212_ & new_n37109_;
  assign new_n37111_ = pi0681 & ~new_n36464_;
  assign new_n37112_ = ~new_n17291_ & ~new_n37111_;
  assign new_n37113_ = new_n6212_ & new_n37112_;
  assign new_n37114_ = pi0223 & ~new_n37113_;
  assign new_n37115_ = ~new_n37110_ & new_n37114_;
  assign new_n37116_ = ~pi0223 & pi0681;
  assign new_n37117_ = new_n17478_ & new_n37116_;
  assign new_n37118_ = pi0215 & ~new_n37117_;
  assign new_n37119_ = ~new_n37115_ & new_n37118_;
  assign new_n37120_ = pi0299 & ~new_n37119_;
  assign new_n37121_ = ~new_n37107_ & new_n37120_;
  assign new_n37122_ = new_n3057_ & ~new_n37088_;
  assign new_n37123_ = ~new_n6238_ & new_n37100_;
  assign new_n37124_ = new_n6238_ & new_n37098_;
  assign new_n37125_ = ~new_n3057_ & ~new_n37124_;
  assign new_n37126_ = ~new_n37123_ & new_n37125_;
  assign new_n37127_ = ~new_n37122_ & ~new_n37126_;
  assign new_n37128_ = ~pi0223 & ~new_n37127_;
  assign new_n37129_ = ~new_n6238_ & ~new_n37109_;
  assign new_n37130_ = new_n6238_ & ~new_n37112_;
  assign new_n37131_ = pi0223 & ~new_n37130_;
  assign new_n37132_ = ~new_n37129_ & new_n37131_;
  assign new_n37133_ = ~pi0299 & ~new_n37132_;
  assign new_n37134_ = ~new_n37128_ & new_n37133_;
  assign new_n37135_ = pi0039 & ~new_n37134_;
  assign new_n37136_ = ~new_n37121_ & new_n37135_;
  assign new_n37137_ = ~new_n37087_ & ~new_n37136_;
  assign new_n37138_ = ~pi0038 & ~new_n37137_;
  assign new_n37139_ = pi0223 & ~new_n17431_;
  assign new_n37140_ = pi0681 & new_n17543_;
  assign new_n37141_ = pi0038 & ~new_n37140_;
  assign new_n37142_ = ~new_n37139_ & new_n37141_;
  assign new_n37143_ = new_n3272_ & ~new_n37142_;
  assign new_n37144_ = ~new_n37138_ & new_n37143_;
  assign new_n37145_ = ~new_n36886_ & ~new_n37144_;
  assign new_n37146_ = ~pi0778 & ~new_n37145_;
  assign new_n37147_ = pi0625 & new_n37145_;
  assign new_n37148_ = ~pi0625 & ~new_n36883_;
  assign new_n37149_ = pi1153 & ~new_n37148_;
  assign new_n37150_ = ~new_n37147_ & new_n37149_;
  assign new_n37151_ = ~pi0625 & new_n37145_;
  assign new_n37152_ = pi0625 & ~new_n36883_;
  assign new_n37153_ = ~pi1153 & ~new_n37152_;
  assign new_n37154_ = ~new_n37151_ & new_n37153_;
  assign new_n37155_ = ~new_n37150_ & ~new_n37154_;
  assign new_n37156_ = pi0778 & ~new_n37155_;
  assign new_n37157_ = ~new_n37146_ & ~new_n37156_;
  assign new_n37158_ = ~new_n17618_ & new_n37157_;
  assign new_n37159_ = ~new_n37072_ & ~new_n37158_;
  assign new_n37160_ = ~new_n17655_ & new_n37159_;
  assign new_n37161_ = new_n17655_ & new_n36883_;
  assign new_n37162_ = ~new_n37160_ & ~new_n37161_;
  assign new_n37163_ = ~new_n17691_ & new_n37162_;
  assign new_n37164_ = ~new_n17734_ & new_n37163_;
  assign new_n37165_ = ~new_n37071_ & ~new_n37164_;
  assign new_n37166_ = ~new_n19311_ & ~new_n37165_;
  assign new_n37167_ = new_n18010_ & ~new_n36883_;
  assign new_n37168_ = ~new_n37166_ & ~new_n37167_;
  assign new_n37169_ = pi0647 & ~new_n37168_;
  assign new_n37170_ = ~pi0647 & ~new_n36883_;
  assign new_n37171_ = pi1157 & ~new_n37170_;
  assign new_n37172_ = ~new_n37169_ & new_n37171_;
  assign new_n37173_ = ~pi0630 & new_n37172_;
  assign new_n37174_ = ~pi0647 & ~new_n37168_;
  assign new_n37175_ = pi0647 & ~new_n36883_;
  assign new_n37176_ = ~pi1157 & ~new_n37175_;
  assign new_n37177_ = ~new_n37174_ & new_n37176_;
  assign new_n37178_ = pi0630 & new_n37177_;
  assign new_n37179_ = ~new_n37173_ & ~new_n37178_;
  assign new_n37180_ = ~new_n37070_ & new_n37179_;
  assign new_n37181_ = pi0787 & ~new_n37180_;
  assign new_n37182_ = ~new_n20567_ & new_n37066_;
  assign new_n37183_ = ~pi0628 & ~new_n37165_;
  assign new_n37184_ = pi0628 & ~new_n36883_;
  assign new_n37185_ = new_n17760_ & ~new_n37184_;
  assign new_n37186_ = ~new_n37183_ & new_n37185_;
  assign new_n37187_ = pi0628 & ~new_n37165_;
  assign new_n37188_ = ~pi0628 & ~new_n36883_;
  assign new_n37189_ = new_n17759_ & ~new_n37188_;
  assign new_n37190_ = ~new_n37187_ & new_n37189_;
  assign new_n37191_ = ~new_n37186_ & ~new_n37190_;
  assign new_n37192_ = ~new_n37182_ & new_n37191_;
  assign new_n37193_ = pi0792 & ~new_n37192_;
  assign new_n37194_ = ~pi0626 & ~new_n37064_;
  assign new_n37195_ = pi0626 & new_n36883_;
  assign new_n37196_ = new_n17732_ & ~new_n37195_;
  assign new_n37197_ = ~new_n37194_ & new_n37196_;
  assign new_n37198_ = new_n17691_ & ~new_n36883_;
  assign new_n37199_ = ~new_n37163_ & ~new_n37198_;
  assign new_n37200_ = new_n17856_ & ~new_n37199_;
  assign new_n37201_ = pi0626 & ~new_n37064_;
  assign new_n37202_ = ~pi0626 & new_n36883_;
  assign new_n37203_ = new_n17731_ & ~new_n37202_;
  assign new_n37204_ = ~new_n37201_ & new_n37203_;
  assign new_n37205_ = ~new_n37200_ & ~new_n37204_;
  assign new_n37206_ = ~new_n37197_ & new_n37205_;
  assign new_n37207_ = pi0788 & ~new_n37206_;
  assign new_n37208_ = ~new_n36914_ & ~new_n37074_;
  assign new_n37209_ = ~pi0642 & ~new_n6179_;
  assign new_n37210_ = ~new_n16823_ & new_n37209_;
  assign new_n37211_ = pi0642 & new_n16935_;
  assign new_n37212_ = pi0680 & ~new_n37211_;
  assign new_n37213_ = ~new_n16830_ & new_n37212_;
  assign new_n37214_ = ~new_n37210_ & new_n37213_;
  assign new_n37215_ = ~new_n37208_ & ~new_n37214_;
  assign new_n37216_ = ~new_n36919_ & ~new_n37215_;
  assign new_n37217_ = ~new_n6212_ & ~new_n37216_;
  assign new_n37218_ = ~pi0680 & ~new_n36922_;
  assign new_n37219_ = pi0642 & ~new_n17021_;
  assign new_n37220_ = ~new_n16640_ & ~new_n37219_;
  assign new_n37221_ = new_n35877_ & ~new_n37220_;
  assign new_n37222_ = pi0680 & ~new_n37221_;
  assign new_n37223_ = pi0642 & ~new_n16948_;
  assign new_n37224_ = new_n6179_ & ~new_n37223_;
  assign new_n37225_ = ~pi0642 & ~new_n16854_;
  assign new_n37226_ = new_n37224_ & ~new_n37225_;
  assign new_n37227_ = new_n37222_ & ~new_n37226_;
  assign new_n37228_ = ~new_n37218_ & ~new_n37227_;
  assign new_n37229_ = pi0681 & ~new_n37228_;
  assign new_n37230_ = ~new_n36926_ & ~new_n37229_;
  assign new_n37231_ = new_n6212_ & ~new_n37230_;
  assign new_n37232_ = ~pi0223 & ~new_n37231_;
  assign new_n37233_ = ~new_n37217_ & new_n37232_;
  assign new_n37234_ = ~new_n36893_ & ~new_n37074_;
  assign new_n37235_ = ~pi0642 & ~new_n16640_;
  assign new_n37236_ = pi0642 & new_n16947_;
  assign new_n37237_ = ~new_n37235_ & ~new_n37236_;
  assign new_n37238_ = new_n16647_ & ~new_n37237_;
  assign new_n37239_ = ~new_n16633_ & new_n37238_;
  assign new_n37240_ = ~new_n6179_ & ~new_n37239_;
  assign new_n37241_ = pi0680 & ~new_n37240_;
  assign new_n37242_ = ~new_n16744_ & ~new_n37219_;
  assign new_n37243_ = new_n6179_ & ~new_n37242_;
  assign new_n37244_ = new_n37241_ & ~new_n37243_;
  assign new_n37245_ = ~new_n37234_ & ~new_n37244_;
  assign new_n37246_ = new_n36899_ & ~new_n37245_;
  assign new_n37247_ = ~new_n36904_ & ~new_n37074_;
  assign new_n37248_ = new_n36548_ & new_n37209_;
  assign new_n37249_ = new_n16707_ & ~new_n36553_;
  assign new_n37250_ = pi0642 & ~new_n36558_;
  assign new_n37251_ = pi0680 & ~new_n37250_;
  assign new_n37252_ = ~new_n37249_ & new_n37251_;
  assign new_n37253_ = ~new_n37248_ & new_n37252_;
  assign new_n37254_ = ~new_n37247_ & ~new_n37253_;
  assign new_n37255_ = new_n36909_ & ~new_n37254_;
  assign new_n37256_ = pi0223 & ~new_n37255_;
  assign new_n37257_ = ~new_n37246_ & new_n37256_;
  assign new_n37258_ = ~new_n3467_ & ~new_n37257_;
  assign new_n37259_ = ~new_n37233_ & new_n37258_;
  assign new_n37260_ = new_n36887_ & ~new_n37074_;
  assign new_n37261_ = new_n37074_ & ~new_n37235_;
  assign new_n37262_ = ~new_n36723_ & new_n37261_;
  assign new_n37263_ = ~new_n37260_ & ~new_n37262_;
  assign new_n37264_ = new_n16636_ & ~new_n37263_;
  assign new_n37265_ = ~pi0223 & new_n37264_;
  assign new_n37266_ = new_n37074_ & new_n37238_;
  assign new_n37267_ = new_n36965_ & ~new_n37074_;
  assign new_n37268_ = pi0223 & ~new_n37267_;
  assign new_n37269_ = ~new_n37266_ & new_n37268_;
  assign new_n37270_ = new_n36938_ & ~new_n37269_;
  assign new_n37271_ = ~new_n37265_ & new_n37270_;
  assign new_n37272_ = ~pi0215 & ~new_n37271_;
  assign new_n37273_ = ~new_n37259_ & new_n37272_;
  assign new_n37274_ = ~new_n36963_ & ~new_n37074_;
  assign new_n37275_ = ~pi0614 & new_n16676_;
  assign new_n37276_ = ~new_n37219_ & ~new_n37275_;
  assign new_n37277_ = ~pi0616 & ~new_n37276_;
  assign new_n37278_ = new_n37241_ & ~new_n37277_;
  assign new_n37279_ = ~new_n37274_ & ~new_n37278_;
  assign new_n37280_ = ~new_n36969_ & ~new_n37279_;
  assign new_n37281_ = new_n6212_ & ~new_n37280_;
  assign new_n37282_ = ~pi0680 & new_n36974_;
  assign new_n37283_ = ~new_n6179_ & new_n16710_;
  assign new_n37284_ = pi0642 & ~new_n36618_;
  assign new_n37285_ = pi0680 & ~new_n16712_;
  assign new_n37286_ = ~new_n37284_ & new_n37285_;
  assign new_n37287_ = ~new_n37283_ & new_n37286_;
  assign new_n37288_ = pi0681 & ~new_n37287_;
  assign new_n37289_ = ~new_n37282_ & new_n37288_;
  assign new_n37290_ = ~new_n36976_ & ~new_n37289_;
  assign new_n37291_ = ~new_n6212_ & ~new_n37290_;
  assign new_n37292_ = pi0223 & ~new_n37291_;
  assign new_n37293_ = ~new_n37281_ & new_n37292_;
  assign new_n37294_ = ~new_n36951_ & ~new_n37074_;
  assign new_n37295_ = new_n16879_ & new_n16985_;
  assign new_n37296_ = new_n16707_ & ~new_n37295_;
  assign new_n37297_ = pi0642 & new_n36638_;
  assign new_n37298_ = ~new_n16871_ & new_n37209_;
  assign new_n37299_ = pi0680 & ~new_n37298_;
  assign new_n37300_ = ~new_n37297_ & new_n37299_;
  assign new_n37301_ = ~new_n37296_ & new_n37300_;
  assign new_n37302_ = ~new_n37294_ & ~new_n37301_;
  assign new_n37303_ = ~new_n6212_ & new_n36949_;
  assign new_n37304_ = ~new_n37302_ & new_n37303_;
  assign new_n37305_ = ~new_n16880_ & new_n37224_;
  assign new_n37306_ = new_n37222_ & ~new_n37305_;
  assign new_n37307_ = ~new_n37218_ & ~new_n37306_;
  assign new_n37308_ = pi0681 & ~new_n37307_;
  assign new_n37309_ = new_n36954_ & ~new_n37308_;
  assign new_n37310_ = ~pi0223 & ~new_n37309_;
  assign new_n37311_ = ~new_n37304_ & new_n37310_;
  assign new_n37312_ = pi0215 & ~new_n37311_;
  assign new_n37313_ = ~new_n37293_ & new_n37312_;
  assign new_n37314_ = pi0299 & ~new_n37313_;
  assign new_n37315_ = ~new_n37273_ & new_n37314_;
  assign new_n37316_ = new_n6238_ & new_n37230_;
  assign new_n37317_ = ~new_n6238_ & new_n37216_;
  assign new_n37318_ = ~new_n3057_ & ~new_n37317_;
  assign new_n37319_ = ~new_n37316_ & new_n37318_;
  assign new_n37320_ = new_n3057_ & ~new_n37264_;
  assign new_n37321_ = ~pi0223 & ~new_n37320_;
  assign new_n37322_ = ~new_n37319_ & new_n37321_;
  assign new_n37323_ = new_n6238_ & new_n37280_;
  assign new_n37324_ = ~new_n6238_ & new_n37290_;
  assign new_n37325_ = pi0223 & ~new_n37324_;
  assign new_n37326_ = ~new_n37323_ & new_n37325_;
  assign new_n37327_ = ~pi0299 & ~new_n37326_;
  assign new_n37328_ = ~new_n37322_ & new_n37327_;
  assign new_n37329_ = pi0039 & ~new_n37328_;
  assign new_n37330_ = ~new_n37315_ & new_n37329_;
  assign new_n37331_ = new_n17175_ & ~new_n37074_;
  assign new_n37332_ = pi0223 & ~new_n37010_;
  assign new_n37333_ = ~new_n36695_ & new_n37332_;
  assign new_n37334_ = ~new_n37331_ & new_n37333_;
  assign new_n37335_ = new_n17176_ & new_n37116_;
  assign new_n37336_ = new_n37009_ & ~new_n37335_;
  assign new_n37337_ = ~new_n37334_ & new_n37336_;
  assign new_n37338_ = new_n17163_ & ~new_n37074_;
  assign new_n37339_ = ~new_n36713_ & new_n37005_;
  assign new_n37340_ = ~new_n37338_ & new_n37339_;
  assign new_n37341_ = new_n17164_ & new_n37116_;
  assign new_n37342_ = new_n37003_ & ~new_n37341_;
  assign new_n37343_ = ~new_n37340_ & new_n37342_;
  assign new_n37344_ = ~pi0039 & ~new_n37343_;
  assign new_n37345_ = ~new_n37337_ & new_n37344_;
  assign new_n37346_ = ~pi0038 & ~new_n37345_;
  assign new_n37347_ = ~new_n37330_ & new_n37346_;
  assign new_n37348_ = new_n37263_ & ~new_n37269_;
  assign new_n37349_ = new_n37021_ & ~new_n37348_;
  assign new_n37350_ = new_n37019_ & ~new_n37349_;
  assign new_n37351_ = new_n3272_ & ~new_n37350_;
  assign new_n37352_ = ~new_n37347_ & new_n37351_;
  assign new_n37353_ = ~new_n36886_ & ~new_n37352_;
  assign new_n37354_ = ~pi0625 & new_n37353_;
  assign new_n37355_ = pi0625 & new_n37026_;
  assign new_n37356_ = ~pi1153 & ~new_n37355_;
  assign new_n37357_ = ~new_n37354_ & new_n37356_;
  assign new_n37358_ = ~pi0608 & ~new_n37357_;
  assign new_n37359_ = ~new_n37150_ & new_n37358_;
  assign new_n37360_ = pi0625 & new_n37353_;
  assign new_n37361_ = ~pi0625 & new_n37026_;
  assign new_n37362_ = pi1153 & ~new_n37361_;
  assign new_n37363_ = ~new_n37360_ & new_n37362_;
  assign new_n37364_ = pi0608 & ~new_n37363_;
  assign new_n37365_ = ~new_n37154_ & new_n37364_;
  assign new_n37366_ = ~new_n37359_ & ~new_n37365_;
  assign new_n37367_ = pi0778 & ~new_n37366_;
  assign new_n37368_ = ~pi0778 & new_n37353_;
  assign new_n37369_ = ~new_n37367_ & ~new_n37368_;
  assign new_n37370_ = ~pi0609 & ~new_n37369_;
  assign new_n37371_ = pi0609 & new_n37157_;
  assign new_n37372_ = ~pi1155 & ~new_n37371_;
  assign new_n37373_ = ~new_n37370_ & new_n37372_;
  assign new_n37374_ = ~pi0660 & ~new_n37033_;
  assign new_n37375_ = ~new_n37373_ & new_n37374_;
  assign new_n37376_ = pi0609 & ~new_n37369_;
  assign new_n37377_ = ~pi0609 & new_n37157_;
  assign new_n37378_ = pi1155 & ~new_n37377_;
  assign new_n37379_ = ~new_n37376_ & new_n37378_;
  assign new_n37380_ = pi0660 & ~new_n37037_;
  assign new_n37381_ = ~new_n37379_ & new_n37380_;
  assign new_n37382_ = ~new_n37375_ & ~new_n37381_;
  assign new_n37383_ = pi0785 & ~new_n37382_;
  assign new_n37384_ = ~pi0785 & ~new_n37369_;
  assign new_n37385_ = ~new_n37383_ & ~new_n37384_;
  assign new_n37386_ = ~pi0618 & ~new_n37385_;
  assign new_n37387_ = pi0618 & ~new_n37159_;
  assign new_n37388_ = ~pi1154 & ~new_n37387_;
  assign new_n37389_ = ~new_n37386_ & new_n37388_;
  assign new_n37390_ = ~pi0627 & ~new_n37045_;
  assign new_n37391_ = ~new_n37389_ & new_n37390_;
  assign new_n37392_ = pi0618 & ~new_n37385_;
  assign new_n37393_ = ~pi0618 & ~new_n37159_;
  assign new_n37394_ = pi1154 & ~new_n37393_;
  assign new_n37395_ = ~new_n37392_ & new_n37394_;
  assign new_n37396_ = pi0627 & ~new_n37049_;
  assign new_n37397_ = ~new_n37395_ & new_n37396_;
  assign new_n37398_ = ~new_n37391_ & ~new_n37397_;
  assign new_n37399_ = pi0781 & ~new_n37398_;
  assign new_n37400_ = ~pi0781 & ~new_n37385_;
  assign new_n37401_ = ~new_n37399_ & ~new_n37400_;
  assign new_n37402_ = pi0619 & ~new_n37401_;
  assign new_n37403_ = ~pi0619 & new_n37162_;
  assign new_n37404_ = pi1159 & ~new_n37403_;
  assign new_n37405_ = ~new_n37402_ & new_n37404_;
  assign new_n37406_ = pi0648 & ~new_n37061_;
  assign new_n37407_ = ~new_n37405_ & new_n37406_;
  assign new_n37408_ = ~pi0619 & ~new_n37401_;
  assign new_n37409_ = pi0619 & new_n37162_;
  assign new_n37410_ = ~pi1159 & ~new_n37409_;
  assign new_n37411_ = ~new_n37408_ & new_n37410_;
  assign new_n37412_ = ~pi0648 & ~new_n37057_;
  assign new_n37413_ = ~new_n37411_ & new_n37412_;
  assign new_n37414_ = pi0789 & ~new_n37413_;
  assign new_n37415_ = ~new_n37407_ & new_n37414_;
  assign new_n37416_ = ~pi0789 & new_n37401_;
  assign new_n37417_ = new_n17969_ & ~new_n37416_;
  assign new_n37418_ = ~new_n37415_ & new_n37417_;
  assign new_n37419_ = ~new_n37207_ & ~new_n37418_;
  assign new_n37420_ = ~new_n37193_ & ~new_n37419_;
  assign new_n37421_ = new_n20364_ & new_n37192_;
  assign new_n37422_ = ~new_n20360_ & ~new_n37421_;
  assign new_n37423_ = ~new_n37420_ & new_n37422_;
  assign new_n37424_ = ~new_n37181_ & ~new_n37423_;
  assign new_n37425_ = pi0644 & new_n37424_;
  assign new_n37426_ = ~pi0787 & new_n37168_;
  assign new_n37427_ = ~new_n37172_ & ~new_n37177_;
  assign new_n37428_ = pi0787 & ~new_n37427_;
  assign new_n37429_ = ~new_n37426_ & ~new_n37428_;
  assign new_n37430_ = ~pi0644 & new_n37429_;
  assign new_n37431_ = pi0715 & ~new_n37430_;
  assign new_n37432_ = ~new_n37425_ & new_n37431_;
  assign new_n37433_ = new_n17804_ & ~new_n36883_;
  assign new_n37434_ = ~new_n17804_ & new_n37069_;
  assign new_n37435_ = ~new_n37433_ & ~new_n37434_;
  assign new_n37436_ = pi0644 & ~new_n37435_;
  assign new_n37437_ = ~pi0644 & ~new_n36883_;
  assign new_n37438_ = ~pi0715 & ~new_n37437_;
  assign new_n37439_ = ~new_n37436_ & new_n37438_;
  assign new_n37440_ = pi1160 & ~new_n37439_;
  assign new_n37441_ = ~new_n37432_ & new_n37440_;
  assign new_n37442_ = ~pi0644 & new_n37424_;
  assign new_n37443_ = pi0644 & new_n37429_;
  assign new_n37444_ = ~pi0715 & ~new_n37443_;
  assign new_n37445_ = ~new_n37442_ & new_n37444_;
  assign new_n37446_ = ~pi0644 & ~new_n37435_;
  assign new_n37447_ = pi0644 & ~new_n36883_;
  assign new_n37448_ = pi0715 & ~new_n37447_;
  assign new_n37449_ = ~new_n37446_ & new_n37448_;
  assign new_n37450_ = ~pi1160 & ~new_n37449_;
  assign new_n37451_ = ~new_n37445_ & new_n37450_;
  assign new_n37452_ = ~new_n37441_ & ~new_n37451_;
  assign new_n37453_ = pi0790 & ~new_n37452_;
  assign new_n37454_ = ~pi0790 & new_n37424_;
  assign new_n37455_ = ~new_n37453_ & ~new_n37454_;
  assign new_n37456_ = ~po1038 & ~new_n37455_;
  assign new_n37457_ = ~pi0223 & po1038;
  assign po0380 = ~new_n37456_ & ~new_n37457_;
  assign new_n37459_ = pi0224 & ~new_n36258_;
  assign new_n37460_ = new_n17968_ & ~new_n37459_;
  assign new_n37461_ = pi0224 & ~new_n3272_;
  assign new_n37462_ = pi0614 & new_n16639_;
  assign new_n37463_ = new_n16636_ & ~new_n37462_;
  assign new_n37464_ = ~new_n6180_ & ~new_n37463_;
  assign new_n37465_ = ~new_n16692_ & ~new_n37464_;
  assign new_n37466_ = ~new_n16630_ & ~new_n37465_;
  assign new_n37467_ = ~pi0680 & ~new_n37465_;
  assign new_n37468_ = pi0680 & new_n37462_;
  assign new_n37469_ = ~new_n17278_ & ~new_n37468_;
  assign new_n37470_ = ~new_n37467_ & new_n37469_;
  assign new_n37471_ = new_n16630_ & ~new_n37470_;
  assign new_n37472_ = ~new_n37466_ & ~new_n37471_;
  assign new_n37473_ = new_n6238_ & new_n37472_;
  assign new_n37474_ = pi0614 & ~new_n16870_;
  assign new_n37475_ = ~new_n36000_ & ~new_n37474_;
  assign new_n37476_ = ~pi0680 & ~new_n37475_;
  assign new_n37477_ = pi0680 & ~new_n17370_;
  assign new_n37478_ = ~new_n36002_ & new_n37477_;
  assign new_n37479_ = ~new_n37476_ & ~new_n37478_;
  assign new_n37480_ = new_n16630_ & ~new_n37479_;
  assign new_n37481_ = ~new_n16630_ & ~new_n37475_;
  assign new_n37482_ = ~new_n37480_ & ~new_n37481_;
  assign new_n37483_ = ~new_n6238_ & new_n37482_;
  assign new_n37484_ = pi0224 & ~new_n37483_;
  assign new_n37485_ = ~new_n37473_ & new_n37484_;
  assign new_n37486_ = pi0614 & ~new_n36327_;
  assign new_n37487_ = ~pi0224 & new_n37486_;
  assign new_n37488_ = ~new_n17419_ & new_n37487_;
  assign new_n37489_ = pi0223 & ~new_n37488_;
  assign new_n37490_ = ~new_n37485_ & new_n37489_;
  assign new_n37491_ = ~new_n16755_ & ~new_n37464_;
  assign new_n37492_ = ~new_n16630_ & ~new_n37491_;
  assign new_n37493_ = ~pi0680 & ~new_n37491_;
  assign new_n37494_ = ~new_n17304_ & ~new_n37468_;
  assign new_n37495_ = ~new_n37493_ & new_n37494_;
  assign new_n37496_ = new_n16630_ & ~new_n37495_;
  assign new_n37497_ = ~new_n37492_ & ~new_n37496_;
  assign new_n37498_ = new_n6238_ & new_n37497_;
  assign new_n37499_ = ~new_n6185_ & new_n16752_;
  assign new_n37500_ = new_n6179_ & ~new_n16770_;
  assign new_n37501_ = ~new_n37499_ & new_n37500_;
  assign new_n37502_ = pi0614 & ~new_n16822_;
  assign new_n37503_ = ~pi0614 & pi0616;
  assign new_n37504_ = new_n16771_ & new_n37503_;
  assign new_n37505_ = ~new_n37502_ & ~new_n37504_;
  assign new_n37506_ = ~new_n37501_ & new_n37505_;
  assign new_n37507_ = ~new_n16630_ & ~new_n37506_;
  assign new_n37508_ = ~pi0680 & ~new_n37506_;
  assign new_n37509_ = pi0614 & new_n16780_;
  assign new_n37510_ = pi0680 & ~new_n37509_;
  assign new_n37511_ = new_n16738_ & new_n37510_;
  assign new_n37512_ = ~new_n37468_ & ~new_n37511_;
  assign new_n37513_ = ~new_n37508_ & new_n37512_;
  assign new_n37514_ = new_n16630_ & ~new_n37513_;
  assign new_n37515_ = ~new_n37507_ & ~new_n37514_;
  assign new_n37516_ = ~new_n6238_ & new_n37515_;
  assign new_n37517_ = pi0224 & ~new_n37516_;
  assign new_n37518_ = ~new_n37498_ & new_n37517_;
  assign new_n37519_ = ~new_n16771_ & new_n37462_;
  assign new_n37520_ = ~pi0680 & ~new_n37519_;
  assign new_n37521_ = ~new_n37510_ & ~new_n37520_;
  assign new_n37522_ = new_n16630_ & ~new_n37521_;
  assign new_n37523_ = ~new_n16630_ & ~new_n37519_;
  assign new_n37524_ = ~new_n37522_ & ~new_n37523_;
  assign new_n37525_ = ~new_n6238_ & ~new_n37524_;
  assign new_n37526_ = pi0614 & ~new_n36297_;
  assign new_n37527_ = new_n6238_ & ~new_n37526_;
  assign new_n37528_ = new_n5791_ & ~new_n37527_;
  assign new_n37529_ = ~new_n37525_ & new_n37528_;
  assign new_n37530_ = pi0614 & new_n16911_;
  assign new_n37531_ = ~pi0223 & ~new_n37530_;
  assign new_n37532_ = ~new_n37529_ & new_n37531_;
  assign new_n37533_ = ~new_n37518_ & new_n37532_;
  assign new_n37534_ = ~new_n37490_ & ~new_n37533_;
  assign new_n37535_ = ~pi0299 & ~new_n37534_;
  assign new_n37536_ = new_n6212_ & new_n37497_;
  assign new_n37537_ = ~new_n6212_ & new_n37515_;
  assign new_n37538_ = pi0224 & ~new_n37537_;
  assign new_n37539_ = ~new_n37536_ & new_n37538_;
  assign new_n37540_ = ~new_n6212_ & ~new_n37524_;
  assign new_n37541_ = new_n6212_ & ~new_n37526_;
  assign new_n37542_ = ~pi0224 & ~new_n37541_;
  assign new_n37543_ = ~new_n37540_ & new_n37542_;
  assign new_n37544_ = ~new_n3467_ & ~new_n37543_;
  assign new_n37545_ = ~new_n37539_ & new_n37544_;
  assign new_n37546_ = pi0224 & ~new_n16636_;
  assign new_n37547_ = new_n3467_ & ~new_n37546_;
  assign new_n37548_ = new_n16639_ & new_n17308_;
  assign new_n37549_ = new_n37547_ & ~new_n37548_;
  assign new_n37550_ = ~pi0215 & ~new_n37549_;
  assign new_n37551_ = ~new_n37545_ & new_n37550_;
  assign new_n37552_ = ~new_n17409_ & new_n37487_;
  assign new_n37553_ = new_n6212_ & new_n37472_;
  assign new_n37554_ = ~new_n6212_ & new_n37482_;
  assign new_n37555_ = pi0224 & ~new_n37554_;
  assign new_n37556_ = ~new_n37553_ & new_n37555_;
  assign new_n37557_ = ~new_n37552_ & ~new_n37556_;
  assign new_n37558_ = pi0215 & ~new_n37557_;
  assign new_n37559_ = pi0299 & ~new_n37558_;
  assign new_n37560_ = ~new_n37551_ & new_n37559_;
  assign new_n37561_ = pi0039 & ~new_n37560_;
  assign new_n37562_ = ~new_n37535_ & new_n37561_;
  assign new_n37563_ = pi0614 & new_n17213_;
  assign new_n37564_ = pi0224 & new_n17172_;
  assign new_n37565_ = new_n37563_ & ~new_n37564_;
  assign new_n37566_ = pi0224 & ~new_n17193_;
  assign new_n37567_ = ~new_n37565_ & ~new_n37566_;
  assign new_n37568_ = pi0299 & new_n37567_;
  assign new_n37569_ = ~pi0614 & new_n17208_;
  assign new_n37570_ = pi0224 & ~new_n37569_;
  assign new_n37571_ = new_n17224_ & new_n37570_;
  assign new_n37572_ = pi0614 & new_n17208_;
  assign new_n37573_ = ~pi0224 & new_n37572_;
  assign new_n37574_ = ~pi0299 & ~new_n37573_;
  assign new_n37575_ = ~new_n37571_ & new_n37574_;
  assign new_n37576_ = ~pi0039 & ~new_n37575_;
  assign new_n37577_ = ~new_n37568_ & new_n37576_;
  assign new_n37578_ = ~pi0038 & ~new_n37577_;
  assign new_n37579_ = ~new_n37562_ & new_n37578_;
  assign new_n37580_ = pi0224 & ~new_n17431_;
  assign new_n37581_ = pi0038 & ~new_n37580_;
  assign new_n37582_ = pi0614 & new_n17433_;
  assign new_n37583_ = new_n37581_ & ~new_n37582_;
  assign new_n37584_ = new_n3272_ & ~new_n37583_;
  assign new_n37585_ = ~new_n37579_ & new_n37584_;
  assign new_n37586_ = ~new_n37461_ & ~new_n37585_;
  assign new_n37587_ = ~new_n17590_ & ~new_n37586_;
  assign new_n37588_ = new_n17590_ & new_n37459_;
  assign new_n37589_ = ~new_n37587_ & ~new_n37588_;
  assign new_n37590_ = ~pi0785 & ~new_n37589_;
  assign new_n37591_ = pi0609 & new_n37589_;
  assign new_n37592_ = ~pi0609 & ~new_n37459_;
  assign new_n37593_ = pi1155 & ~new_n37592_;
  assign new_n37594_ = ~new_n37591_ & new_n37593_;
  assign new_n37595_ = ~pi0609 & new_n37589_;
  assign new_n37596_ = pi0609 & ~new_n37459_;
  assign new_n37597_ = ~pi1155 & ~new_n37596_;
  assign new_n37598_ = ~new_n37595_ & new_n37597_;
  assign new_n37599_ = ~new_n37594_ & ~new_n37598_;
  assign new_n37600_ = pi0785 & ~new_n37599_;
  assign new_n37601_ = ~new_n37590_ & ~new_n37600_;
  assign new_n37602_ = ~pi0781 & ~new_n37601_;
  assign new_n37603_ = pi0618 & new_n37601_;
  assign new_n37604_ = ~pi0618 & ~new_n37459_;
  assign new_n37605_ = pi1154 & ~new_n37604_;
  assign new_n37606_ = ~new_n37603_ & new_n37605_;
  assign new_n37607_ = ~pi0618 & new_n37601_;
  assign new_n37608_ = pi0618 & ~new_n37459_;
  assign new_n37609_ = ~pi1154 & ~new_n37608_;
  assign new_n37610_ = ~new_n37607_ & new_n37609_;
  assign new_n37611_ = ~new_n37606_ & ~new_n37610_;
  assign new_n37612_ = pi0781 & ~new_n37611_;
  assign new_n37613_ = ~new_n37602_ & ~new_n37612_;
  assign new_n37614_ = ~pi0789 & ~new_n37613_;
  assign new_n37615_ = pi0619 & new_n37613_;
  assign new_n37616_ = ~pi0619 & ~new_n37459_;
  assign new_n37617_ = pi1159 & ~new_n37616_;
  assign new_n37618_ = ~new_n37615_ & new_n37617_;
  assign new_n37619_ = ~pi0619 & new_n37613_;
  assign new_n37620_ = pi0619 & ~new_n37459_;
  assign new_n37621_ = ~pi1159 & ~new_n37620_;
  assign new_n37622_ = ~new_n37619_ & new_n37621_;
  assign new_n37623_ = ~new_n37618_ & ~new_n37622_;
  assign new_n37624_ = pi0789 & ~new_n37623_;
  assign new_n37625_ = ~new_n37614_ & ~new_n37624_;
  assign new_n37626_ = ~new_n17968_ & new_n37625_;
  assign new_n37627_ = ~new_n37460_ & ~new_n37626_;
  assign new_n37628_ = ~new_n20567_ & new_n37627_;
  assign new_n37629_ = ~new_n19279_ & ~new_n37459_;
  assign new_n37630_ = ~pi0224 & ~new_n17168_;
  assign new_n37631_ = pi0662 & pi0680;
  assign new_n37632_ = new_n17168_ & ~new_n37631_;
  assign new_n37633_ = pi0224 & new_n17196_;
  assign new_n37634_ = pi0299 & ~new_n37633_;
  assign new_n37635_ = ~new_n37632_ & new_n37634_;
  assign new_n37636_ = ~new_n37630_ & new_n37635_;
  assign new_n37637_ = ~pi0224 & ~new_n17154_;
  assign new_n37638_ = new_n17154_ & ~new_n37631_;
  assign new_n37639_ = pi0224 & new_n17187_;
  assign new_n37640_ = ~pi0299 & ~new_n37639_;
  assign new_n37641_ = ~new_n37638_ & new_n37640_;
  assign new_n37642_ = ~new_n37637_ & new_n37641_;
  assign new_n37643_ = ~pi0039 & ~new_n37642_;
  assign new_n37644_ = ~new_n37636_ & new_n37643_;
  assign new_n37645_ = new_n16812_ & new_n37631_;
  assign new_n37646_ = new_n37547_ & ~new_n37645_;
  assign new_n37647_ = pi0662 & ~new_n17489_;
  assign new_n37648_ = ~pi0662 & ~new_n17313_;
  assign new_n37649_ = ~new_n37647_ & ~new_n37648_;
  assign new_n37650_ = new_n6212_ & new_n37649_;
  assign new_n37651_ = ~new_n6181_ & ~new_n36445_;
  assign new_n37652_ = new_n17320_ & ~new_n37651_;
  assign new_n37653_ = ~new_n6212_ & new_n37652_;
  assign new_n37654_ = pi0224 & ~new_n37653_;
  assign new_n37655_ = ~new_n37650_ & new_n37654_;
  assign new_n37656_ = ~new_n17454_ & new_n37631_;
  assign new_n37657_ = new_n6212_ & ~new_n37656_;
  assign new_n37658_ = pi0662 & new_n17449_;
  assign new_n37659_ = ~new_n6212_ & ~new_n37658_;
  assign new_n37660_ = ~pi0224 & ~new_n37659_;
  assign new_n37661_ = ~new_n37657_ & new_n37660_;
  assign new_n37662_ = ~new_n3467_ & ~new_n37661_;
  assign new_n37663_ = ~new_n37655_ & new_n37662_;
  assign new_n37664_ = ~new_n37646_ & ~new_n37663_;
  assign new_n37665_ = ~pi0215 & ~new_n37664_;
  assign new_n37666_ = ~pi0662 & ~new_n17272_;
  assign new_n37667_ = pi0662 & ~new_n17510_;
  assign new_n37668_ = ~new_n37666_ & ~new_n37667_;
  assign new_n37669_ = ~new_n6212_ & new_n37668_;
  assign new_n37670_ = ~pi0662 & ~new_n17292_;
  assign new_n37671_ = pi0662 & ~new_n36464_;
  assign new_n37672_ = ~new_n37670_ & ~new_n37671_;
  assign new_n37673_ = new_n6212_ & new_n37672_;
  assign new_n37674_ = pi0224 & ~new_n37673_;
  assign new_n37675_ = ~new_n37669_ & new_n37674_;
  assign new_n37676_ = ~pi0224 & pi0662;
  assign new_n37677_ = new_n17478_ & new_n37676_;
  assign new_n37678_ = pi0215 & ~new_n37677_;
  assign new_n37679_ = ~new_n37675_ & new_n37678_;
  assign new_n37680_ = pi0299 & ~new_n37679_;
  assign new_n37681_ = ~new_n37665_ & new_n37680_;
  assign new_n37682_ = new_n6238_ & new_n37649_;
  assign new_n37683_ = ~new_n6238_ & new_n37652_;
  assign new_n37684_ = pi0224 & ~new_n37683_;
  assign new_n37685_ = ~new_n37682_ & new_n37684_;
  assign new_n37686_ = new_n6238_ & ~new_n37656_;
  assign new_n37687_ = ~new_n6238_ & ~new_n37658_;
  assign new_n37688_ = new_n5791_ & ~new_n37687_;
  assign new_n37689_ = ~new_n37686_ & new_n37688_;
  assign new_n37690_ = pi0662 & new_n17448_;
  assign new_n37691_ = ~pi0223 & ~new_n37690_;
  assign new_n37692_ = ~new_n37689_ & new_n37691_;
  assign new_n37693_ = ~new_n37685_ & new_n37692_;
  assign new_n37694_ = ~new_n6238_ & new_n37668_;
  assign new_n37695_ = new_n6238_ & new_n37672_;
  assign new_n37696_ = pi0224 & ~new_n37695_;
  assign new_n37697_ = ~new_n37694_ & new_n37696_;
  assign new_n37698_ = new_n17465_ & new_n37676_;
  assign new_n37699_ = pi0223 & ~new_n37698_;
  assign new_n37700_ = ~new_n37697_ & new_n37699_;
  assign new_n37701_ = ~pi0299 & ~new_n37700_;
  assign new_n37702_ = ~new_n37693_ & new_n37701_;
  assign new_n37703_ = pi0039 & ~new_n37702_;
  assign new_n37704_ = ~new_n37681_ & new_n37703_;
  assign new_n37705_ = ~new_n37644_ & ~new_n37704_;
  assign new_n37706_ = ~pi0038 & ~new_n37705_;
  assign new_n37707_ = pi0662 & new_n17543_;
  assign new_n37708_ = new_n37581_ & ~new_n37707_;
  assign new_n37709_ = new_n3272_ & ~new_n37708_;
  assign new_n37710_ = ~new_n37706_ & new_n37709_;
  assign new_n37711_ = ~new_n37461_ & ~new_n37710_;
  assign new_n37712_ = ~pi0778 & ~new_n37711_;
  assign new_n37713_ = pi0625 & new_n37711_;
  assign new_n37714_ = ~pi0625 & ~new_n37459_;
  assign new_n37715_ = pi1153 & ~new_n37714_;
  assign new_n37716_ = ~new_n37713_ & new_n37715_;
  assign new_n37717_ = ~pi0625 & new_n37711_;
  assign new_n37718_ = pi0625 & ~new_n37459_;
  assign new_n37719_ = ~pi1153 & ~new_n37718_;
  assign new_n37720_ = ~new_n37717_ & new_n37719_;
  assign new_n37721_ = ~new_n37716_ & ~new_n37720_;
  assign new_n37722_ = pi0778 & ~new_n37721_;
  assign new_n37723_ = ~new_n37712_ & ~new_n37722_;
  assign new_n37724_ = ~new_n17618_ & ~new_n37723_;
  assign new_n37725_ = new_n17618_ & new_n37459_;
  assign new_n37726_ = ~new_n37724_ & ~new_n37725_;
  assign new_n37727_ = ~new_n17655_ & ~new_n37726_;
  assign new_n37728_ = new_n17655_ & new_n37459_;
  assign new_n37729_ = ~new_n37727_ & ~new_n37728_;
  assign new_n37730_ = ~new_n17691_ & new_n37729_;
  assign new_n37731_ = ~new_n17734_ & new_n37730_;
  assign new_n37732_ = ~new_n37629_ & ~new_n37731_;
  assign new_n37733_ = ~pi0628 & ~new_n37732_;
  assign new_n37734_ = pi0628 & ~new_n37459_;
  assign new_n37735_ = new_n17760_ & ~new_n37734_;
  assign new_n37736_ = ~new_n37733_ & new_n37735_;
  assign new_n37737_ = pi0628 & ~new_n37732_;
  assign new_n37738_ = ~pi0628 & ~new_n37459_;
  assign new_n37739_ = new_n17759_ & ~new_n37738_;
  assign new_n37740_ = ~new_n37737_ & new_n37739_;
  assign new_n37741_ = ~new_n37736_ & ~new_n37740_;
  assign new_n37742_ = ~new_n37628_ & new_n37741_;
  assign new_n37743_ = pi0792 & ~new_n37742_;
  assign new_n37744_ = pi0614 & ~new_n36558_;
  assign new_n37745_ = new_n36548_ & new_n37503_;
  assign new_n37746_ = ~new_n37744_ & ~new_n37745_;
  assign new_n37747_ = ~new_n36556_ & new_n37746_;
  assign new_n37748_ = pi0680 & ~new_n37747_;
  assign new_n37749_ = ~new_n37508_ & ~new_n37748_;
  assign new_n37750_ = pi0662 & ~new_n37749_;
  assign new_n37751_ = ~pi0662 & ~new_n16629_;
  assign new_n37752_ = ~new_n37506_ & new_n37751_;
  assign new_n37753_ = ~new_n37514_ & ~new_n37752_;
  assign new_n37754_ = ~new_n37750_ & new_n37753_;
  assign new_n37755_ = pi0224 & new_n37754_;
  assign new_n37756_ = ~pi0614 & new_n16835_;
  assign new_n37757_ = pi0614 & ~new_n16935_;
  assign new_n37758_ = pi0680 & ~new_n37757_;
  assign new_n37759_ = ~new_n37756_ & new_n37758_;
  assign new_n37760_ = ~new_n37520_ & ~new_n37759_;
  assign new_n37761_ = pi0662 & ~new_n37760_;
  assign new_n37762_ = ~new_n37519_ & new_n37751_;
  assign new_n37763_ = ~new_n37522_ & ~new_n37762_;
  assign new_n37764_ = ~new_n37761_ & new_n37763_;
  assign new_n37765_ = ~pi0224 & ~new_n37764_;
  assign new_n37766_ = ~new_n6212_ & ~new_n37765_;
  assign new_n37767_ = ~new_n37755_ & new_n37766_;
  assign new_n37768_ = ~pi0614 & ~new_n24079_;
  assign new_n37769_ = pi0614 & ~new_n36723_;
  assign new_n37770_ = ~new_n37768_ & ~new_n37769_;
  assign new_n37771_ = ~new_n16633_ & new_n37770_;
  assign new_n37772_ = pi0616 & ~new_n37771_;
  assign new_n37773_ = pi0614 & ~new_n17021_;
  assign new_n37774_ = ~new_n16746_ & ~new_n37773_;
  assign new_n37775_ = ~pi0616 & ~new_n37774_;
  assign new_n37776_ = ~new_n37772_ & ~new_n37775_;
  assign new_n37777_ = pi0680 & ~new_n37776_;
  assign new_n37778_ = ~new_n37493_ & ~new_n37777_;
  assign new_n37779_ = pi0662 & ~new_n37778_;
  assign new_n37780_ = ~new_n37491_ & new_n37751_;
  assign new_n37781_ = ~new_n37496_ & ~new_n37780_;
  assign new_n37782_ = ~new_n37779_ & new_n37781_;
  assign new_n37783_ = pi0224 & new_n37782_;
  assign new_n37784_ = ~new_n16843_ & new_n37503_;
  assign new_n37785_ = ~new_n36592_ & ~new_n37784_;
  assign new_n37786_ = pi0680 & ~new_n37785_;
  assign new_n37787_ = ~new_n36593_ & ~new_n37548_;
  assign new_n37788_ = ~new_n37786_ & ~new_n37787_;
  assign new_n37789_ = pi0662 & ~new_n37788_;
  assign new_n37790_ = ~pi0662 & ~new_n37526_;
  assign new_n37791_ = ~new_n37789_ & ~new_n37790_;
  assign new_n37792_ = ~pi0224 & ~new_n37791_;
  assign new_n37793_ = new_n6212_ & ~new_n37792_;
  assign new_n37794_ = ~new_n37783_ & new_n37793_;
  assign new_n37795_ = ~new_n3467_ & ~new_n37794_;
  assign new_n37796_ = ~new_n37767_ & new_n37795_;
  assign new_n37797_ = new_n16843_ & new_n37631_;
  assign new_n37798_ = ~new_n37548_ & ~new_n37797_;
  assign new_n37799_ = ~pi0224 & ~new_n37798_;
  assign new_n37800_ = new_n37631_ & new_n37770_;
  assign new_n37801_ = ~new_n37462_ & ~new_n37631_;
  assign new_n37802_ = new_n16647_ & new_n37801_;
  assign new_n37803_ = pi0224 & ~new_n37802_;
  assign new_n37804_ = ~new_n37800_ & new_n37803_;
  assign new_n37805_ = new_n37547_ & ~new_n37804_;
  assign new_n37806_ = ~new_n37799_ & new_n37805_;
  assign new_n37807_ = ~pi0215 & ~new_n37806_;
  assign new_n37808_ = ~new_n37796_ & new_n37807_;
  assign new_n37809_ = ~new_n16678_ & ~new_n37773_;
  assign new_n37810_ = ~pi0616 & ~new_n37809_;
  assign new_n37811_ = ~new_n37772_ & ~new_n37810_;
  assign new_n37812_ = pi0680 & ~new_n37811_;
  assign new_n37813_ = ~new_n37467_ & ~new_n37812_;
  assign new_n37814_ = pi0662 & ~new_n37813_;
  assign new_n37815_ = ~new_n37465_ & new_n37751_;
  assign new_n37816_ = ~new_n37471_ & ~new_n37815_;
  assign new_n37817_ = ~new_n37814_ & new_n37816_;
  assign new_n37818_ = new_n6212_ & ~new_n37817_;
  assign new_n37819_ = pi0614 & ~new_n36618_;
  assign new_n37820_ = new_n16713_ & ~new_n37819_;
  assign new_n37821_ = pi0680 & ~new_n37820_;
  assign new_n37822_ = ~new_n37476_ & ~new_n37821_;
  assign new_n37823_ = pi0662 & ~new_n37822_;
  assign new_n37824_ = ~new_n37475_ & new_n37751_;
  assign new_n37825_ = ~new_n37480_ & ~new_n37824_;
  assign new_n37826_ = ~new_n37823_ & new_n37825_;
  assign new_n37827_ = ~new_n6212_ & ~new_n37826_;
  assign new_n37828_ = pi0224 & ~new_n37827_;
  assign new_n37829_ = ~new_n37818_ & new_n37828_;
  assign new_n37830_ = pi0680 & ~new_n16895_;
  assign new_n37831_ = ~new_n37548_ & ~new_n37830_;
  assign new_n37832_ = ~new_n37786_ & ~new_n37831_;
  assign new_n37833_ = pi0662 & ~new_n37832_;
  assign new_n37834_ = ~pi0662 & ~new_n37486_;
  assign new_n37835_ = ~new_n37833_ & ~new_n37834_;
  assign new_n37836_ = new_n6212_ & new_n37835_;
  assign new_n37837_ = ~new_n16701_ & new_n37486_;
  assign new_n37838_ = ~pi0662 & ~new_n37837_;
  assign new_n37839_ = ~pi0614 & new_n16872_;
  assign new_n37840_ = pi0614 & new_n36638_;
  assign new_n37841_ = pi0680 & ~new_n37840_;
  assign new_n37842_ = ~new_n37839_ & new_n37841_;
  assign new_n37843_ = ~new_n16882_ & new_n37842_;
  assign new_n37844_ = pi0614 & ~pi0680;
  assign new_n37845_ = new_n16708_ & new_n37844_;
  assign new_n37846_ = pi0662 & ~new_n37845_;
  assign new_n37847_ = ~new_n37843_ & new_n37846_;
  assign new_n37848_ = ~new_n37838_ & ~new_n37847_;
  assign new_n37849_ = ~new_n6212_ & new_n37848_;
  assign new_n37850_ = ~pi0224 & ~new_n37849_;
  assign new_n37851_ = ~new_n37836_ & new_n37850_;
  assign new_n37852_ = pi0215 & ~new_n37851_;
  assign new_n37853_ = ~new_n37829_ & new_n37852_;
  assign new_n37854_ = pi0299 & ~new_n37853_;
  assign new_n37855_ = ~new_n37808_ & new_n37854_;
  assign new_n37856_ = new_n6238_ & new_n37782_;
  assign new_n37857_ = ~new_n6238_ & new_n37754_;
  assign new_n37858_ = pi0224 & ~new_n37857_;
  assign new_n37859_ = ~new_n37856_ & new_n37858_;
  assign new_n37860_ = ~new_n6238_ & ~new_n37764_;
  assign new_n37861_ = new_n6238_ & ~new_n37791_;
  assign new_n37862_ = new_n5791_ & ~new_n37861_;
  assign new_n37863_ = ~new_n37860_ & new_n37862_;
  assign new_n37864_ = ~pi0222 & new_n37799_;
  assign new_n37865_ = ~pi0223 & ~new_n37864_;
  assign new_n37866_ = ~new_n37863_ & new_n37865_;
  assign new_n37867_ = ~new_n37859_ & new_n37866_;
  assign new_n37868_ = pi0224 & new_n37817_;
  assign new_n37869_ = ~pi0224 & ~new_n37835_;
  assign new_n37870_ = new_n6238_ & ~new_n37869_;
  assign new_n37871_ = ~new_n37868_ & new_n37870_;
  assign new_n37872_ = pi0224 & new_n37826_;
  assign new_n37873_ = ~pi0224 & ~new_n37848_;
  assign new_n37874_ = ~new_n6238_ & ~new_n37873_;
  assign new_n37875_ = ~new_n37872_ & new_n37874_;
  assign new_n37876_ = pi0223 & ~new_n37875_;
  assign new_n37877_ = ~new_n37871_ & new_n37876_;
  assign new_n37878_ = ~new_n37867_ & ~new_n37877_;
  assign new_n37879_ = ~pi0299 & ~new_n37878_;
  assign new_n37880_ = pi0039 & ~new_n37879_;
  assign new_n37881_ = ~new_n37855_ & new_n37880_;
  assign new_n37882_ = new_n17163_ & new_n37631_;
  assign new_n37883_ = ~new_n37572_ & ~new_n37882_;
  assign new_n37884_ = ~pi0224 & ~new_n37883_;
  assign new_n37885_ = new_n17163_ & ~new_n37631_;
  assign new_n37886_ = ~new_n36713_ & new_n37570_;
  assign new_n37887_ = ~new_n37885_ & new_n37886_;
  assign new_n37888_ = ~new_n37884_ & ~new_n37887_;
  assign new_n37889_ = ~pi0299 & ~new_n37888_;
  assign new_n37890_ = ~pi0614 & new_n17213_;
  assign new_n37891_ = ~new_n36695_ & ~new_n37890_;
  assign new_n37892_ = pi0224 & ~new_n37891_;
  assign new_n37893_ = ~pi0224 & ~new_n17175_;
  assign new_n37894_ = ~new_n37563_ & new_n37893_;
  assign new_n37895_ = ~new_n37892_ & ~new_n37894_;
  assign new_n37896_ = new_n37631_ & ~new_n37895_;
  assign new_n37897_ = new_n37567_ & ~new_n37631_;
  assign new_n37898_ = pi0299 & ~new_n37897_;
  assign new_n37899_ = ~new_n37896_ & new_n37898_;
  assign new_n37900_ = ~new_n37889_ & ~new_n37899_;
  assign new_n37901_ = ~pi0039 & ~new_n37900_;
  assign new_n37902_ = ~pi0038 & ~new_n37901_;
  assign new_n37903_ = ~new_n37881_ & new_n37902_;
  assign new_n37904_ = pi0662 & new_n16790_;
  assign new_n37905_ = new_n17431_ & new_n37904_;
  assign new_n37906_ = new_n37583_ & ~new_n37905_;
  assign new_n37907_ = new_n3272_ & ~new_n37906_;
  assign new_n37908_ = ~new_n37903_ & new_n37907_;
  assign new_n37909_ = ~new_n37461_ & ~new_n37908_;
  assign new_n37910_ = ~pi0625 & new_n37909_;
  assign new_n37911_ = pi0625 & new_n37586_;
  assign new_n37912_ = ~pi1153 & ~new_n37911_;
  assign new_n37913_ = ~new_n37910_ & new_n37912_;
  assign new_n37914_ = ~pi0608 & ~new_n37716_;
  assign new_n37915_ = ~new_n37913_ & new_n37914_;
  assign new_n37916_ = pi0625 & new_n37909_;
  assign new_n37917_ = ~pi0625 & new_n37586_;
  assign new_n37918_ = pi1153 & ~new_n37917_;
  assign new_n37919_ = ~new_n37916_ & new_n37918_;
  assign new_n37920_ = pi0608 & ~new_n37720_;
  assign new_n37921_ = ~new_n37919_ & new_n37920_;
  assign new_n37922_ = ~new_n37915_ & ~new_n37921_;
  assign new_n37923_ = pi0778 & ~new_n37922_;
  assign new_n37924_ = ~pi0778 & new_n37909_;
  assign new_n37925_ = ~new_n37923_ & ~new_n37924_;
  assign new_n37926_ = ~pi0609 & ~new_n37925_;
  assign new_n37927_ = pi0609 & new_n37723_;
  assign new_n37928_ = ~pi1155 & ~new_n37927_;
  assign new_n37929_ = ~new_n37926_ & new_n37928_;
  assign new_n37930_ = ~pi0660 & ~new_n37594_;
  assign new_n37931_ = ~new_n37929_ & new_n37930_;
  assign new_n37932_ = pi0609 & ~new_n37925_;
  assign new_n37933_ = ~pi0609 & new_n37723_;
  assign new_n37934_ = pi1155 & ~new_n37933_;
  assign new_n37935_ = ~new_n37932_ & new_n37934_;
  assign new_n37936_ = pi0660 & ~new_n37598_;
  assign new_n37937_ = ~new_n37935_ & new_n37936_;
  assign new_n37938_ = ~new_n37931_ & ~new_n37937_;
  assign new_n37939_ = pi0785 & ~new_n37938_;
  assign new_n37940_ = ~pi0785 & ~new_n37925_;
  assign new_n37941_ = ~new_n37939_ & ~new_n37940_;
  assign new_n37942_ = ~pi0618 & ~new_n37941_;
  assign new_n37943_ = pi0618 & new_n37726_;
  assign new_n37944_ = ~pi1154 & ~new_n37943_;
  assign new_n37945_ = ~new_n37942_ & new_n37944_;
  assign new_n37946_ = ~pi0627 & ~new_n37606_;
  assign new_n37947_ = ~new_n37945_ & new_n37946_;
  assign new_n37948_ = pi0618 & ~new_n37941_;
  assign new_n37949_ = ~pi0618 & new_n37726_;
  assign new_n37950_ = pi1154 & ~new_n37949_;
  assign new_n37951_ = ~new_n37948_ & new_n37950_;
  assign new_n37952_ = pi0627 & ~new_n37610_;
  assign new_n37953_ = ~new_n37951_ & new_n37952_;
  assign new_n37954_ = ~new_n37947_ & ~new_n37953_;
  assign new_n37955_ = pi0781 & ~new_n37954_;
  assign new_n37956_ = ~pi0781 & ~new_n37941_;
  assign new_n37957_ = ~new_n37955_ & ~new_n37956_;
  assign new_n37958_ = pi0619 & ~new_n37957_;
  assign new_n37959_ = ~pi0619 & new_n37729_;
  assign new_n37960_ = pi1159 & ~new_n37959_;
  assign new_n37961_ = ~new_n37958_ & new_n37960_;
  assign new_n37962_ = pi0648 & ~new_n37622_;
  assign new_n37963_ = ~new_n37961_ & new_n37962_;
  assign new_n37964_ = ~pi0619 & ~new_n37957_;
  assign new_n37965_ = pi0619 & new_n37729_;
  assign new_n37966_ = ~pi1159 & ~new_n37965_;
  assign new_n37967_ = ~new_n37964_ & new_n37966_;
  assign new_n37968_ = ~pi0648 & ~new_n37618_;
  assign new_n37969_ = ~new_n37967_ & new_n37968_;
  assign new_n37970_ = pi0789 & ~new_n37969_;
  assign new_n37971_ = ~new_n37963_ & new_n37970_;
  assign new_n37972_ = ~pi0789 & new_n37957_;
  assign new_n37973_ = new_n17969_ & ~new_n37972_;
  assign new_n37974_ = ~new_n37971_ & new_n37973_;
  assign new_n37975_ = ~pi0626 & ~new_n37625_;
  assign new_n37976_ = pi0626 & new_n37459_;
  assign new_n37977_ = new_n17732_ & ~new_n37976_;
  assign new_n37978_ = ~new_n37975_ & new_n37977_;
  assign new_n37979_ = new_n17691_ & ~new_n37459_;
  assign new_n37980_ = ~new_n37730_ & ~new_n37979_;
  assign new_n37981_ = new_n17856_ & ~new_n37980_;
  assign new_n37982_ = pi0626 & ~new_n37625_;
  assign new_n37983_ = ~pi0626 & new_n37459_;
  assign new_n37984_ = new_n17731_ & ~new_n37983_;
  assign new_n37985_ = ~new_n37982_ & new_n37984_;
  assign new_n37986_ = ~new_n37981_ & ~new_n37985_;
  assign new_n37987_ = ~new_n37978_ & new_n37986_;
  assign new_n37988_ = pi0788 & ~new_n37987_;
  assign new_n37989_ = ~new_n20364_ & ~new_n37988_;
  assign new_n37990_ = ~new_n37974_ & new_n37989_;
  assign new_n37991_ = ~new_n37743_ & ~new_n37990_;
  assign new_n37992_ = ~new_n20360_ & ~new_n37991_;
  assign new_n37993_ = ~new_n17762_ & new_n37627_;
  assign new_n37994_ = new_n17762_ & new_n37459_;
  assign new_n37995_ = ~new_n37993_ & ~new_n37994_;
  assign new_n37996_ = ~new_n20556_ & ~new_n37995_;
  assign new_n37997_ = ~new_n19311_ & ~new_n37732_;
  assign new_n37998_ = new_n18010_ & ~new_n37459_;
  assign new_n37999_ = ~new_n37997_ & ~new_n37998_;
  assign new_n38000_ = pi0647 & ~new_n37999_;
  assign new_n38001_ = ~pi0647 & ~new_n37459_;
  assign new_n38002_ = pi1157 & ~new_n38001_;
  assign new_n38003_ = ~new_n38000_ & new_n38002_;
  assign new_n38004_ = ~pi0630 & new_n38003_;
  assign new_n38005_ = ~pi0647 & ~new_n37999_;
  assign new_n38006_ = pi0647 & ~new_n37459_;
  assign new_n38007_ = ~pi1157 & ~new_n38006_;
  assign new_n38008_ = ~new_n38005_ & new_n38007_;
  assign new_n38009_ = pi0630 & new_n38008_;
  assign new_n38010_ = ~new_n38004_ & ~new_n38009_;
  assign new_n38011_ = ~new_n37996_ & new_n38010_;
  assign new_n38012_ = pi0787 & ~new_n38011_;
  assign new_n38013_ = ~new_n37992_ & ~new_n38012_;
  assign new_n38014_ = pi0644 & new_n38013_;
  assign new_n38015_ = ~pi0787 & new_n37999_;
  assign new_n38016_ = ~new_n38003_ & ~new_n38008_;
  assign new_n38017_ = pi0787 & ~new_n38016_;
  assign new_n38018_ = ~new_n38015_ & ~new_n38017_;
  assign new_n38019_ = ~pi0644 & new_n38018_;
  assign new_n38020_ = pi0715 & ~new_n38019_;
  assign new_n38021_ = ~new_n38014_ & new_n38020_;
  assign new_n38022_ = new_n17804_ & ~new_n37459_;
  assign new_n38023_ = ~new_n17804_ & new_n37995_;
  assign new_n38024_ = ~new_n38022_ & ~new_n38023_;
  assign new_n38025_ = pi0644 & ~new_n38024_;
  assign new_n38026_ = ~pi0644 & ~new_n37459_;
  assign new_n38027_ = ~pi0715 & ~new_n38026_;
  assign new_n38028_ = ~new_n38025_ & new_n38027_;
  assign new_n38029_ = pi1160 & ~new_n38028_;
  assign new_n38030_ = ~new_n38021_ & new_n38029_;
  assign new_n38031_ = ~pi0644 & new_n38013_;
  assign new_n38032_ = pi0644 & new_n38018_;
  assign new_n38033_ = ~pi0715 & ~new_n38032_;
  assign new_n38034_ = ~new_n38031_ & new_n38033_;
  assign new_n38035_ = ~pi0644 & ~new_n38024_;
  assign new_n38036_ = pi0644 & ~new_n37459_;
  assign new_n38037_ = pi0715 & ~new_n38036_;
  assign new_n38038_ = ~new_n38035_ & new_n38037_;
  assign new_n38039_ = ~pi1160 & ~new_n38038_;
  assign new_n38040_ = ~new_n38034_ & new_n38039_;
  assign new_n38041_ = ~new_n38030_ & ~new_n38040_;
  assign new_n38042_ = pi0790 & ~new_n38041_;
  assign new_n38043_ = ~pi0790 & new_n38013_;
  assign new_n38044_ = ~new_n38042_ & ~new_n38043_;
  assign new_n38045_ = ~po1038 & ~new_n38044_;
  assign new_n38046_ = ~pi0224 & po1038;
  assign po0381 = ~new_n38045_ & ~new_n38046_;
  assign new_n38048_ = ~new_n6166_ & new_n6263_;
  assign new_n38049_ = ~pi0137 & ~new_n38048_;
  assign new_n38050_ = new_n6259_ & ~new_n38049_;
  assign new_n38051_ = new_n2926_ & ~new_n11417_;
  assign new_n38052_ = ~new_n2712_ & new_n38051_;
  assign new_n38053_ = new_n2556_ & ~new_n38052_;
  assign new_n38054_ = new_n2554_ & ~new_n38053_;
  assign new_n38055_ = ~new_n2741_ & ~new_n38054_;
  assign new_n38056_ = ~pi0095 & ~new_n38055_;
  assign new_n38057_ = ~new_n2726_ & ~new_n38056_;
  assign new_n38058_ = pi0137 & ~new_n38057_;
  assign new_n38059_ = new_n2450_ & new_n11417_;
  assign new_n38060_ = new_n2784_ & ~new_n38059_;
  assign new_n38061_ = new_n2794_ & ~new_n38060_;
  assign new_n38062_ = ~pi0137 & ~new_n38061_;
  assign new_n38063_ = ~new_n38058_ & ~new_n38062_;
  assign new_n38064_ = pi0332 & ~new_n38063_;
  assign new_n38065_ = ~new_n2726_ & ~new_n2743_;
  assign new_n38066_ = pi0137 & ~new_n38065_;
  assign new_n38067_ = ~new_n2828_ & ~new_n38066_;
  assign new_n38068_ = ~pi0332 & ~new_n38067_;
  assign new_n38069_ = ~new_n38064_ & ~new_n38068_;
  assign new_n38070_ = new_n2993_ & new_n38069_;
  assign new_n38071_ = pi1093 & ~new_n38061_;
  assign new_n38072_ = new_n2794_ & new_n2800_;
  assign new_n38073_ = new_n2450_ & ~new_n7481_;
  assign new_n38074_ = ~new_n2531_ & new_n38073_;
  assign new_n38075_ = ~pi0032 & ~new_n38074_;
  assign new_n38076_ = new_n38072_ & ~new_n38075_;
  assign new_n38077_ = ~pi1093 & ~new_n38076_;
  assign new_n38078_ = ~new_n2800_ & new_n38061_;
  assign new_n38079_ = new_n11416_ & new_n38073_;
  assign new_n38080_ = new_n38072_ & new_n38079_;
  assign new_n38081_ = ~new_n38078_ & ~new_n38080_;
  assign new_n38082_ = new_n38077_ & new_n38081_;
  assign new_n38083_ = ~new_n38071_ & ~new_n38082_;
  assign new_n38084_ = new_n11547_ & ~new_n38083_;
  assign new_n38085_ = ~new_n2800_ & new_n2827_;
  assign new_n38086_ = new_n38077_ & ~new_n38085_;
  assign new_n38087_ = ~new_n2767_ & new_n38073_;
  assign new_n38088_ = ~pi0032 & ~new_n38087_;
  assign new_n38089_ = new_n38072_ & ~new_n38088_;
  assign new_n38090_ = pi1093 & ~new_n38085_;
  assign new_n38091_ = ~new_n38089_ & new_n38090_;
  assign new_n38092_ = ~new_n38086_ & ~new_n38091_;
  assign new_n38093_ = new_n11514_ & ~new_n38092_;
  assign new_n38094_ = new_n38081_ & new_n38093_;
  assign new_n38095_ = ~new_n38084_ & ~new_n38094_;
  assign new_n38096_ = ~new_n38058_ & new_n38095_;
  assign new_n38097_ = pi0332 & ~new_n38096_;
  assign new_n38098_ = pi1093 & ~new_n2827_;
  assign new_n38099_ = ~new_n38086_ & ~new_n38098_;
  assign new_n38100_ = new_n11547_ & ~new_n38099_;
  assign new_n38101_ = ~new_n38093_ & ~new_n38100_;
  assign new_n38102_ = ~new_n38066_ & new_n38101_;
  assign new_n38103_ = ~pi0332 & ~new_n38102_;
  assign new_n38104_ = ~new_n38097_ & ~new_n38103_;
  assign new_n38105_ = ~new_n2993_ & new_n38104_;
  assign new_n38106_ = ~pi0210 & ~new_n38105_;
  assign new_n38107_ = ~new_n38070_ & new_n38106_;
  assign new_n38108_ = ~new_n2723_ & ~new_n2726_;
  assign new_n38109_ = pi0137 & ~new_n38108_;
  assign new_n38110_ = ~new_n2786_ & ~new_n38109_;
  assign new_n38111_ = ~pi0332 & ~new_n38110_;
  assign new_n38112_ = ~new_n2501_ & ~new_n38054_;
  assign new_n38113_ = ~pi0095 & ~new_n38112_;
  assign new_n38114_ = new_n3025_ & ~new_n38113_;
  assign new_n38115_ = ~pi0137 & new_n2502_;
  assign new_n38116_ = ~new_n38060_ & new_n38115_;
  assign new_n38117_ = pi0332 & ~new_n38116_;
  assign new_n38118_ = ~new_n38114_ & new_n38117_;
  assign new_n38119_ = ~new_n38111_ & ~new_n38118_;
  assign new_n38120_ = pi0210 & ~new_n38119_;
  assign new_n38121_ = pi0299 & ~new_n38120_;
  assign new_n38122_ = ~new_n38107_ & new_n38121_;
  assign new_n38123_ = ~new_n6260_ & new_n38104_;
  assign new_n38124_ = new_n6260_ & new_n38069_;
  assign new_n38125_ = ~pi0198 & ~new_n38124_;
  assign new_n38126_ = ~new_n38123_ & new_n38125_;
  assign new_n38127_ = pi0198 & ~new_n38119_;
  assign new_n38128_ = ~pi0299 & ~new_n38127_;
  assign new_n38129_ = ~new_n38126_ & new_n38128_;
  assign new_n38130_ = ~new_n38122_ & ~new_n38129_;
  assign new_n38131_ = ~pi0039 & ~new_n38130_;
  assign new_n38132_ = pi0039 & new_n3115_;
  assign new_n38133_ = ~pi0038 & ~new_n38132_;
  assign new_n38134_ = ~new_n38131_ & new_n38133_;
  assign new_n38135_ = pi0038 & ~pi0137;
  assign new_n38136_ = new_n6134_ & ~new_n38135_;
  assign new_n38137_ = ~new_n38134_ & new_n38136_;
  assign new_n38138_ = ~new_n38050_ & ~new_n38137_;
  assign new_n38139_ = ~pi0087 & ~new_n38138_;
  assign new_n38140_ = new_n3115_ & new_n3212_;
  assign new_n38141_ = pi0087 & new_n38140_;
  assign new_n38142_ = ~pi0075 & ~new_n38141_;
  assign new_n38143_ = ~new_n38139_ & new_n38142_;
  assign new_n38144_ = new_n7301_ & ~new_n38049_;
  assign new_n38145_ = pi0075 & ~new_n38144_;
  assign new_n38146_ = ~pi0092 & ~new_n38145_;
  assign new_n38147_ = ~new_n38143_ & new_n38146_;
  assign new_n38148_ = pi0092 & new_n3235_;
  assign new_n38149_ = new_n38140_ & new_n38148_;
  assign new_n38150_ = ~pi0054 & ~new_n38149_;
  assign new_n38151_ = ~new_n38147_ & new_n38150_;
  assign new_n38152_ = new_n3282_ & new_n38140_;
  assign new_n38153_ = pi0054 & ~new_n38152_;
  assign new_n38154_ = ~pi0074 & ~new_n38153_;
  assign new_n38155_ = ~new_n38151_ & new_n38154_;
  assign new_n38156_ = pi0074 & new_n6128_;
  assign new_n38157_ = new_n38140_ & new_n38156_;
  assign new_n38158_ = ~pi0055 & ~new_n38157_;
  assign new_n38159_ = ~new_n38155_ & new_n38158_;
  assign new_n38160_ = new_n7348_ & ~new_n38159_;
  assign new_n38161_ = pi0056 & new_n3284_;
  assign new_n38162_ = new_n38140_ & new_n38161_;
  assign new_n38163_ = ~new_n38160_ & ~new_n38162_;
  assign new_n38164_ = ~pi0062 & ~new_n38163_;
  assign new_n38165_ = new_n3437_ & new_n38140_;
  assign new_n38166_ = pi0062 & new_n38165_;
  assign new_n38167_ = new_n3436_ & ~new_n38166_;
  assign new_n38168_ = ~new_n38164_ & new_n38167_;
  assign new_n38169_ = ~pi0062 & new_n38165_;
  assign new_n38170_ = ~new_n3436_ & ~new_n38169_;
  assign new_n38171_ = ~new_n6120_ & ~new_n38170_;
  assign po0382 = ~new_n38168_ & new_n38171_;
  assign new_n38173_ = pi0228 & pi0231;
  assign new_n38174_ = ~new_n2525_ & ~new_n2872_;
  assign new_n38175_ = ~pi0070 & ~new_n38174_;
  assign new_n38176_ = ~pi0051 & ~new_n38175_;
  assign new_n38177_ = new_n2559_ & ~new_n38176_;
  assign new_n38178_ = new_n2926_ & ~new_n38177_;
  assign new_n38179_ = new_n2556_ & ~new_n38178_;
  assign new_n38180_ = new_n2554_ & ~new_n38179_;
  assign new_n38181_ = ~new_n6173_ & ~new_n38180_;
  assign new_n38182_ = ~pi0095 & ~new_n38181_;
  assign new_n38183_ = new_n2787_ & ~new_n38182_;
  assign new_n38184_ = ~pi0039 & ~new_n38183_;
  assign new_n38185_ = ~pi0038 & ~new_n3357_;
  assign new_n38186_ = ~new_n38184_ & new_n38185_;
  assign new_n38187_ = ~pi0228 & new_n38186_;
  assign new_n38188_ = ~new_n38173_ & ~new_n38187_;
  assign new_n38189_ = ~pi0100 & ~new_n38188_;
  assign new_n38190_ = ~new_n14006_ & ~new_n38173_;
  assign new_n38191_ = pi0100 & ~new_n38190_;
  assign new_n38192_ = ~pi0087 & ~new_n38191_;
  assign new_n38193_ = ~new_n38189_ & new_n38192_;
  assign new_n38194_ = pi0087 & ~new_n38173_;
  assign new_n38195_ = ~new_n7356_ & new_n38194_;
  assign new_n38196_ = ~pi0075 & ~new_n38195_;
  assign new_n38197_ = ~new_n38193_ & new_n38196_;
  assign new_n38198_ = ~new_n14014_ & ~new_n38173_;
  assign new_n38199_ = pi0075 & ~new_n38198_;
  assign new_n38200_ = ~pi0092 & ~new_n38199_;
  assign new_n38201_ = ~new_n38197_ & new_n38200_;
  assign new_n38202_ = pi0092 & ~new_n38173_;
  assign new_n38203_ = ~new_n7382_ & new_n38202_;
  assign new_n38204_ = ~new_n38201_ & ~new_n38203_;
  assign new_n38205_ = ~pi0054 & ~new_n38204_;
  assign new_n38206_ = pi0054 & ~new_n38173_;
  assign new_n38207_ = ~pi0074 & ~new_n38206_;
  assign new_n38208_ = ~new_n38205_ & new_n38207_;
  assign new_n38209_ = ~new_n7391_ & ~new_n38173_;
  assign new_n38210_ = pi0074 & ~new_n38209_;
  assign new_n38211_ = ~pi0055 & ~new_n38210_;
  assign new_n38212_ = ~new_n38208_ & new_n38211_;
  assign new_n38213_ = pi0055 & ~new_n38173_;
  assign new_n38214_ = ~pi0056 & ~new_n38213_;
  assign new_n38215_ = ~new_n38212_ & new_n38214_;
  assign new_n38216_ = ~new_n7397_ & ~new_n38173_;
  assign new_n38217_ = pi0056 & ~new_n38216_;
  assign new_n38218_ = ~pi0062 & ~new_n38217_;
  assign new_n38219_ = ~new_n38215_ & new_n38218_;
  assign new_n38220_ = pi0062 & ~new_n38173_;
  assign new_n38221_ = ~new_n7357_ & new_n38220_;
  assign new_n38222_ = ~new_n38219_ & ~new_n38221_;
  assign new_n38223_ = new_n3436_ & ~new_n38222_;
  assign new_n38224_ = ~new_n3436_ & ~new_n38173_;
  assign po0383 = ~new_n38223_ & ~new_n38224_;
  assign new_n38226_ = new_n2497_ & new_n6356_;
  assign new_n38227_ = new_n2532_ & new_n11032_;
  assign new_n38228_ = new_n11030_ & new_n38227_;
  assign new_n38229_ = ~pi0091 & ~new_n2570_;
  assign new_n38230_ = ~new_n2799_ & new_n11022_;
  assign new_n38231_ = new_n38229_ & ~new_n38230_;
  assign new_n38232_ = ~new_n38228_ & new_n38231_;
  assign new_n38233_ = new_n38226_ & ~new_n38232_;
  assign new_n38234_ = ~pi0072 & ~new_n38233_;
  assign new_n38235_ = new_n6380_ & ~new_n38234_;
  assign new_n38236_ = pi0829 & ~new_n6196_;
  assign new_n38237_ = ~new_n38235_ & new_n38236_;
  assign new_n38238_ = new_n13091_ & ~new_n13116_;
  assign new_n38239_ = new_n6380_ & new_n38238_;
  assign new_n38240_ = ~new_n6469_ & ~new_n38239_;
  assign new_n38241_ = pi1093 & ~new_n38240_;
  assign new_n38242_ = new_n11022_ & new_n38226_;
  assign new_n38243_ = ~new_n7511_ & new_n38242_;
  assign new_n38244_ = new_n38226_ & ~new_n38229_;
  assign new_n38245_ = ~pi0072 & ~new_n38244_;
  assign new_n38246_ = ~new_n8903_ & new_n38245_;
  assign new_n38247_ = ~new_n38243_ & new_n38246_;
  assign new_n38248_ = new_n6380_ & ~new_n38247_;
  assign new_n38249_ = ~new_n38241_ & ~new_n38248_;
  assign new_n38250_ = ~new_n38242_ & new_n38245_;
  assign new_n38251_ = new_n6380_ & ~new_n38250_;
  assign new_n38252_ = new_n10068_ & ~new_n38251_;
  assign new_n38253_ = ~new_n38249_ & ~new_n38252_;
  assign new_n38254_ = ~new_n38237_ & new_n38253_;
  assign new_n38255_ = ~pi0039 & ~new_n38254_;
  assign po0384 = ~new_n11471_ | new_n38255_;
  assign new_n38257_ = ~pi0039 & pi0228;
  assign new_n38258_ = ~new_n11420_ & ~new_n11425_;
  assign new_n38259_ = pi0039 & ~new_n38258_;
  assign new_n38260_ = new_n6465_ & new_n38259_;
  assign new_n38261_ = ~new_n2797_ & ~new_n8904_;
  assign new_n38262_ = ~pi0032 & new_n10235_;
  assign new_n38263_ = ~new_n38261_ & new_n38262_;
  assign new_n38264_ = new_n2541_ & new_n38263_;
  assign new_n38265_ = ~new_n11487_ & new_n38264_;
  assign new_n38266_ = ~new_n38260_ & ~new_n38265_;
  assign new_n38267_ = new_n10200_ & ~new_n38266_;
  assign po0385 = new_n38257_ | new_n38267_;
  assign new_n38269_ = ~new_n6133_ & new_n10197_;
  assign new_n38270_ = pi0824 & ~new_n17138_;
  assign new_n38271_ = pi0829 & pi1091;
  assign new_n38272_ = new_n17143_ & new_n38271_;
  assign new_n38273_ = ~pi0824 & ~new_n38272_;
  assign new_n38274_ = new_n38271_ & new_n38273_;
  assign new_n38275_ = ~new_n38270_ & ~new_n38274_;
  assign new_n38276_ = new_n2799_ & ~new_n6461_;
  assign new_n38277_ = ~new_n38275_ & new_n38276_;
  assign new_n38278_ = ~new_n6166_ & ~new_n6461_;
  assign new_n38279_ = ~new_n6461_ & ~new_n38273_;
  assign new_n38280_ = ~new_n38270_ & new_n38279_;
  assign new_n38281_ = ~new_n17102_ & ~new_n38280_;
  assign new_n38282_ = ~new_n38278_ & ~new_n38281_;
  assign new_n38283_ = ~new_n38277_ & new_n38282_;
  assign new_n38284_ = ~new_n7511_ & new_n17102_;
  assign new_n38285_ = ~new_n17119_ & ~new_n38284_;
  assign new_n38286_ = new_n38278_ & ~new_n38285_;
  assign new_n38287_ = pi1093 & ~new_n38286_;
  assign new_n38288_ = ~new_n38283_ & new_n38287_;
  assign new_n38289_ = ~new_n6277_ & new_n17102_;
  assign new_n38290_ = new_n6167_ & new_n17090_;
  assign new_n38291_ = ~new_n17092_ & new_n38290_;
  assign new_n38292_ = ~pi0040 & ~new_n38291_;
  assign new_n38293_ = new_n10281_ & ~new_n38292_;
  assign new_n38294_ = pi0252 & ~new_n38293_;
  assign new_n38295_ = new_n6277_ & ~new_n17089_;
  assign new_n38296_ = ~new_n38294_ & new_n38295_;
  assign new_n38297_ = ~pi1093 & ~new_n38296_;
  assign new_n38298_ = ~new_n38289_ & new_n38297_;
  assign new_n38299_ = ~pi0039 & ~new_n38298_;
  assign new_n38300_ = ~new_n38288_ & new_n38299_;
  assign new_n38301_ = ~new_n6221_ & new_n16635_;
  assign new_n38302_ = ~new_n6194_ & new_n7510_;
  assign new_n38303_ = new_n16632_ & ~new_n38302_;
  assign new_n38304_ = new_n16722_ & new_n38302_;
  assign new_n38305_ = pi1091 & ~new_n38304_;
  assign new_n38306_ = ~new_n38303_ & new_n38305_;
  assign new_n38307_ = ~new_n6457_ & new_n16632_;
  assign new_n38308_ = new_n6457_ & new_n16722_;
  assign new_n38309_ = ~pi1091 & ~new_n38308_;
  assign new_n38310_ = ~new_n38307_ & new_n38309_;
  assign new_n38311_ = ~new_n38306_ & ~new_n38310_;
  assign new_n38312_ = ~pi0120 & ~new_n38311_;
  assign new_n38313_ = ~new_n16634_ & ~new_n38312_;
  assign new_n38314_ = new_n6221_ & new_n38313_;
  assign new_n38315_ = ~new_n38301_ & ~new_n38314_;
  assign new_n38316_ = new_n6238_ & new_n38315_;
  assign new_n38317_ = ~new_n6215_ & new_n38313_;
  assign new_n38318_ = ~new_n35720_ & ~new_n38317_;
  assign new_n38319_ = ~new_n6238_ & new_n38318_;
  assign new_n38320_ = ~new_n3057_ & ~new_n38319_;
  assign new_n38321_ = ~new_n38316_ & new_n38320_;
  assign new_n38322_ = new_n3057_ & new_n16635_;
  assign new_n38323_ = ~pi0223 & ~new_n38322_;
  assign new_n38324_ = ~new_n38321_ & new_n38323_;
  assign new_n38325_ = pi0120 & new_n6199_;
  assign new_n38326_ = new_n16635_ & ~new_n38325_;
  assign new_n38327_ = ~new_n38301_ & ~new_n38326_;
  assign new_n38328_ = new_n6238_ & ~new_n38327_;
  assign new_n38329_ = ~new_n35720_ & ~new_n38326_;
  assign new_n38330_ = ~new_n6238_ & ~new_n38329_;
  assign new_n38331_ = pi0223 & ~new_n38330_;
  assign new_n38332_ = ~new_n38328_ & new_n38331_;
  assign new_n38333_ = ~pi0299 & ~new_n38332_;
  assign new_n38334_ = ~new_n38324_ & new_n38333_;
  assign new_n38335_ = new_n6212_ & new_n38315_;
  assign new_n38336_ = ~new_n6212_ & new_n38318_;
  assign new_n38337_ = ~new_n3467_ & ~new_n38336_;
  assign new_n38338_ = ~new_n38335_ & new_n38337_;
  assign new_n38339_ = ~pi0215 & ~new_n17405_;
  assign new_n38340_ = ~new_n38338_ & new_n38339_;
  assign new_n38341_ = new_n6212_ & ~new_n38327_;
  assign new_n38342_ = ~new_n6212_ & ~new_n38329_;
  assign new_n38343_ = pi0215 & ~new_n38342_;
  assign new_n38344_ = ~new_n38341_ & new_n38343_;
  assign new_n38345_ = pi0299 & ~new_n38344_;
  assign new_n38346_ = ~new_n38340_ & new_n38345_;
  assign new_n38347_ = ~new_n38334_ & ~new_n38346_;
  assign new_n38348_ = pi0039 & ~new_n38347_;
  assign new_n38349_ = ~pi0038 & ~new_n38348_;
  assign new_n38350_ = ~new_n38300_ & new_n38349_;
  assign po0387 = new_n38269_ & ~new_n38350_;
  assign new_n38352_ = ~pi0081 & ~new_n2674_;
  assign new_n38353_ = new_n6341_ & ~new_n38352_;
  assign new_n38354_ = new_n2451_ & ~new_n38353_;
  assign new_n38355_ = new_n2682_ & ~new_n38354_;
  assign new_n38356_ = new_n2594_ & ~new_n38355_;
  assign new_n38357_ = new_n2686_ & ~new_n38356_;
  assign new_n38358_ = new_n2504_ & ~new_n38357_;
  assign new_n38359_ = ~new_n2507_ & ~new_n38358_;
  assign new_n38360_ = ~pi0086 & ~new_n38359_;
  assign new_n38361_ = new_n2592_ & ~new_n38360_;
  assign new_n38362_ = new_n2590_ & ~new_n38361_;
  assign new_n38363_ = ~new_n2585_ & ~new_n38362_;
  assign new_n38364_ = ~pi0108 & ~new_n38363_;
  assign new_n38365_ = new_n2584_ & ~new_n38364_;
  assign new_n38366_ = new_n2698_ & ~new_n38365_;
  assign new_n38367_ = ~new_n2575_ & ~new_n38366_;
  assign new_n38368_ = new_n2574_ & ~new_n38367_;
  assign new_n38369_ = new_n2573_ & ~new_n38368_;
  assign new_n38370_ = new_n2566_ & ~new_n38369_;
  assign new_n38371_ = new_n2857_ & ~new_n38370_;
  assign new_n38372_ = new_n2547_ & ~new_n38371_;
  assign new_n38373_ = new_n15622_ & ~new_n38372_;
  assign new_n38374_ = ~pi0070 & ~new_n38373_;
  assign new_n38375_ = ~new_n2848_ & ~new_n38374_;
  assign new_n38376_ = ~pi0051 & ~new_n38375_;
  assign new_n38377_ = new_n2559_ & ~new_n38376_;
  assign new_n38378_ = new_n2926_ & ~new_n38377_;
  assign new_n38379_ = new_n2556_ & ~new_n38378_;
  assign new_n38380_ = ~pi1082 & new_n2553_;
  assign new_n38381_ = ~pi0032 & ~new_n38380_;
  assign new_n38382_ = ~new_n38379_ & new_n38381_;
  assign new_n38383_ = ~new_n3367_ & ~new_n38382_;
  assign new_n38384_ = ~pi0095 & ~new_n38383_;
  assign new_n38385_ = ~new_n2726_ & ~new_n38384_;
  assign new_n38386_ = ~pi0039 & ~new_n38385_;
  assign new_n38387_ = ~new_n7307_ & ~new_n7309_;
  assign po0950 = ~new_n2799_ | ~new_n6198_;
  assign new_n38389_ = new_n6455_ & ~po0950;
  assign new_n38390_ = ~new_n38387_ & new_n38389_;
  assign new_n38391_ = new_n6190_ & new_n11369_;
  assign new_n38392_ = ~new_n38390_ & new_n38391_;
  assign new_n38393_ = ~new_n3357_ & ~new_n38392_;
  assign new_n38394_ = ~new_n38386_ & new_n38393_;
  assign new_n38395_ = ~pi0038 & ~new_n38394_;
  assign new_n38396_ = new_n6134_ & ~new_n38395_;
  assign new_n38397_ = ~pi0087 & ~new_n6259_;
  assign new_n38398_ = ~new_n38396_ & new_n38397_;
  assign new_n38399_ = ~new_n6288_ & ~new_n38398_;
  assign new_n38400_ = new_n3242_ & ~new_n38399_;
  assign new_n38401_ = new_n7306_ & ~new_n38400_;
  assign new_n38402_ = ~pi0054 & ~new_n38401_;
  assign new_n38403_ = ~new_n7341_ & ~new_n38402_;
  assign new_n38404_ = new_n8879_ & ~new_n38403_;
  assign new_n38405_ = new_n15712_ & ~new_n38404_;
  assign new_n38406_ = ~pi0056 & ~new_n38405_;
  assign new_n38407_ = ~new_n6127_ & ~new_n38406_;
  assign new_n38408_ = ~pi0062 & ~new_n38407_;
  assign new_n38409_ = ~new_n6299_ & ~new_n38408_;
  assign new_n38410_ = new_n3436_ & ~new_n38409_;
  assign po0389 = new_n6123_ & ~new_n38410_;
  assign new_n38412_ = ~pi0230 & ~pi0233;
  assign new_n38413_ = ~pi0212 & ~pi0214;
  assign new_n38414_ = ~pi0211 & ~new_n38413_;
  assign new_n38415_ = pi0219 & ~new_n38414_;
  assign new_n38416_ = po1038 & ~new_n38415_;
  assign new_n38417_ = pi1142 & ~new_n10486_;
  assign new_n38418_ = pi0211 & pi1143;
  assign new_n38419_ = ~pi0211 & pi1144;
  assign new_n38420_ = ~new_n38418_ & ~new_n38419_;
  assign new_n38421_ = ~pi0212 & pi0214;
  assign new_n38422_ = pi0212 & ~pi0214;
  assign new_n38423_ = ~new_n38421_ & ~new_n38422_;
  assign new_n38424_ = ~new_n38420_ & ~new_n38423_;
  assign new_n38425_ = ~pi0211 & pi1143;
  assign new_n38426_ = new_n10729_ & new_n38425_;
  assign new_n38427_ = ~new_n38424_ & ~new_n38426_;
  assign new_n38428_ = ~pi0219 & ~new_n38427_;
  assign new_n38429_ = ~new_n38417_ & ~new_n38428_;
  assign new_n38430_ = new_n38416_ & ~new_n38429_;
  assign new_n38431_ = pi0299 & ~new_n38420_;
  assign new_n38432_ = pi0199 & pi1142;
  assign new_n38433_ = ~pi0200 & ~new_n38432_;
  assign new_n38434_ = ~pi0199 & pi1144;
  assign new_n38435_ = new_n38433_ & ~new_n38434_;
  assign new_n38436_ = ~pi0199 & pi1143;
  assign new_n38437_ = pi0200 & ~new_n38436_;
  assign new_n38438_ = ~new_n38435_ & ~new_n38437_;
  assign new_n38439_ = ~pi0299 & ~new_n38438_;
  assign new_n38440_ = ~pi0207 & ~new_n38439_;
  assign new_n38441_ = new_n38433_ & ~new_n38436_;
  assign new_n38442_ = pi0207 & ~pi0299;
  assign new_n38443_ = ~pi0199 & pi1142;
  assign new_n38444_ = pi0200 & ~new_n38443_;
  assign new_n38445_ = new_n38442_ & ~new_n38444_;
  assign new_n38446_ = ~new_n38441_ & new_n38445_;
  assign new_n38447_ = ~new_n38440_ & ~new_n38446_;
  assign new_n38448_ = pi0208 & ~new_n38447_;
  assign new_n38449_ = pi0207 & ~pi0208;
  assign new_n38450_ = new_n38438_ & new_n38449_;
  assign new_n38451_ = ~new_n38448_ & ~new_n38450_;
  assign new_n38452_ = ~pi0299 & ~new_n38451_;
  assign new_n38453_ = ~new_n38431_ & ~new_n38452_;
  assign new_n38454_ = ~pi0214 & ~new_n38452_;
  assign new_n38455_ = ~pi0212 & ~new_n38454_;
  assign new_n38456_ = ~new_n38453_ & new_n38455_;
  assign new_n38457_ = ~new_n38431_ & new_n38454_;
  assign new_n38458_ = pi0211 & pi1142;
  assign new_n38459_ = ~new_n38425_ & ~new_n38458_;
  assign new_n38460_ = pi0299 & ~new_n38459_;
  assign new_n38461_ = pi0214 & ~new_n38460_;
  assign new_n38462_ = ~new_n38452_ & new_n38461_;
  assign new_n38463_ = pi0212 & ~new_n38462_;
  assign new_n38464_ = ~new_n38457_ & new_n38463_;
  assign new_n38465_ = ~pi0219 & ~new_n38464_;
  assign new_n38466_ = ~new_n38456_ & new_n38465_;
  assign new_n38467_ = ~pi0299 & new_n38451_;
  assign new_n38468_ = pi0299 & ~pi1142;
  assign new_n38469_ = new_n38414_ & ~new_n38468_;
  assign new_n38470_ = ~new_n38467_ & new_n38469_;
  assign new_n38471_ = ~new_n38414_ & new_n38452_;
  assign new_n38472_ = pi0219 & ~new_n38471_;
  assign new_n38473_ = ~new_n38470_ & new_n38472_;
  assign new_n38474_ = ~po1038 & ~new_n38473_;
  assign new_n38475_ = ~new_n38466_ & new_n38474_;
  assign new_n38476_ = ~new_n38430_ & ~new_n38475_;
  assign new_n38477_ = pi0213 & new_n38476_;
  assign new_n38478_ = ~pi0211 & pi1157;
  assign new_n38479_ = pi0211 & pi1156;
  assign new_n38480_ = ~new_n38478_ & ~new_n38479_;
  assign new_n38481_ = pi0214 & ~new_n38480_;
  assign new_n38482_ = ~pi0212 & ~new_n38481_;
  assign new_n38483_ = ~pi0211 & pi1156;
  assign new_n38484_ = pi0211 & pi1155;
  assign new_n38485_ = ~new_n38483_ & ~new_n38484_;
  assign new_n38486_ = ~pi0214 & ~new_n38485_;
  assign new_n38487_ = ~pi0211 & pi1155;
  assign new_n38488_ = pi0211 & pi1154;
  assign new_n38489_ = ~new_n38487_ & ~new_n38488_;
  assign new_n38490_ = pi0214 & ~new_n38489_;
  assign new_n38491_ = ~new_n38486_ & ~new_n38490_;
  assign new_n38492_ = pi0212 & new_n38491_;
  assign new_n38493_ = ~new_n38482_ & ~new_n38492_;
  assign new_n38494_ = ~pi0219 & ~new_n38493_;
  assign new_n38495_ = ~pi0211 & pi0214;
  assign new_n38496_ = pi1155 & new_n38495_;
  assign new_n38497_ = ~pi0212 & ~new_n38496_;
  assign new_n38498_ = ~pi0211 & pi1154;
  assign new_n38499_ = ~pi0214 & ~new_n38498_;
  assign new_n38500_ = ~pi0211 & pi1153;
  assign new_n38501_ = new_n10729_ & ~new_n38500_;
  assign new_n38502_ = ~new_n38499_ & ~new_n38501_;
  assign new_n38503_ = ~new_n38497_ & new_n38502_;
  assign new_n38504_ = pi0219 & ~new_n38503_;
  assign new_n38505_ = po1038 & ~new_n38504_;
  assign new_n38506_ = ~new_n38494_ & new_n38505_;
  assign new_n38507_ = ~pi0213 & ~new_n38506_;
  assign new_n38508_ = ~pi0219 & pi0299;
  assign new_n38509_ = new_n38493_ & new_n38508_;
  assign new_n38510_ = pi0299 & pi1155;
  assign new_n38511_ = new_n38421_ & new_n38510_;
  assign new_n38512_ = pi0299 & pi1154;
  assign new_n38513_ = ~pi0214 & ~new_n38512_;
  assign new_n38514_ = pi0299 & pi1153;
  assign new_n38515_ = pi0214 & ~new_n38514_;
  assign new_n38516_ = pi0212 & ~new_n38515_;
  assign new_n38517_ = ~new_n38513_ & new_n38516_;
  assign new_n38518_ = ~new_n38511_ & ~new_n38517_;
  assign new_n38519_ = ~pi0211 & pi0219;
  assign new_n38520_ = ~new_n38518_ & new_n38519_;
  assign new_n38521_ = ~new_n38509_ & ~new_n38520_;
  assign new_n38522_ = ~new_n38452_ & new_n38521_;
  assign new_n38523_ = ~po1038 & ~new_n38522_;
  assign new_n38524_ = new_n38507_ & ~new_n38523_;
  assign new_n38525_ = pi0209 & ~new_n38524_;
  assign new_n38526_ = ~new_n38477_ & new_n38525_;
  assign new_n38527_ = ~pi0200 & pi1155;
  assign new_n38528_ = pi0199 & new_n38527_;
  assign new_n38529_ = ~pi0299 & new_n38528_;
  assign new_n38530_ = ~pi1156 & ~new_n38529_;
  assign new_n38531_ = ~pi0200 & ~pi1155;
  assign new_n38532_ = pi0199 & pi0200;
  assign new_n38533_ = ~new_n10817_ & ~new_n38532_;
  assign new_n38534_ = ~pi0299 & new_n38533_;
  assign new_n38535_ = ~new_n38531_ & new_n38534_;
  assign new_n38536_ = ~new_n38530_ & new_n38535_;
  assign new_n38537_ = pi0207 & new_n38536_;
  assign new_n38538_ = ~pi0208 & ~new_n38537_;
  assign new_n38539_ = ~pi0299 & ~new_n38532_;
  assign new_n38540_ = pi1153 & ~new_n38539_;
  assign new_n38541_ = pi1154 & ~new_n38540_;
  assign new_n38542_ = new_n11373_ & new_n38527_;
  assign new_n38543_ = ~pi1153 & ~new_n11373_;
  assign new_n38544_ = pi1154 & new_n38533_;
  assign new_n38545_ = ~new_n38543_ & new_n38544_;
  assign new_n38546_ = ~new_n38542_ & ~new_n38545_;
  assign new_n38547_ = new_n38541_ & ~new_n38546_;
  assign new_n38548_ = ~pi0200 & ~pi0299;
  assign new_n38549_ = pi0199 & ~pi1153;
  assign new_n38550_ = new_n38548_ & ~new_n38549_;
  assign new_n38551_ = ~pi0199 & ~pi1155;
  assign new_n38552_ = ~pi1154 & ~new_n38551_;
  assign new_n38553_ = new_n38550_ & new_n38552_;
  assign new_n38554_ = ~new_n38547_ & ~new_n38553_;
  assign new_n38555_ = pi0207 & new_n38554_;
  assign new_n38556_ = pi0200 & ~pi0299;
  assign new_n38557_ = ~pi0199 & pi1155;
  assign new_n38558_ = new_n38556_ & new_n38557_;
  assign new_n38559_ = ~pi1154 & ~new_n38558_;
  assign new_n38560_ = pi0200 & ~new_n38557_;
  assign new_n38561_ = new_n10820_ & ~new_n38560_;
  assign new_n38562_ = ~new_n38559_ & new_n38561_;
  assign new_n38563_ = pi0200 & ~pi1155;
  assign new_n38564_ = new_n11373_ & ~new_n38563_;
  assign new_n38565_ = pi1156 & new_n38564_;
  assign new_n38566_ = ~new_n38562_ & ~new_n38565_;
  assign new_n38567_ = ~pi0207 & new_n38566_;
  assign new_n38568_ = ~new_n38555_ & ~new_n38567_;
  assign new_n38569_ = pi0208 & ~new_n38568_;
  assign new_n38570_ = ~new_n38538_ & ~new_n38569_;
  assign new_n38571_ = ~pi1157 & ~new_n38570_;
  assign new_n38572_ = pi0199 & ~pi1155;
  assign new_n38573_ = pi1156 & ~new_n38572_;
  assign new_n38574_ = new_n38539_ & new_n38573_;
  assign new_n38575_ = ~pi1156 & ~new_n38572_;
  assign new_n38576_ = new_n38548_ & new_n38575_;
  assign new_n38577_ = ~new_n38574_ & ~new_n38576_;
  assign new_n38578_ = pi0207 & ~new_n38577_;
  assign new_n38579_ = ~pi0208 & ~new_n38578_;
  assign new_n38580_ = ~new_n38569_ & ~new_n38579_;
  assign new_n38581_ = pi1157 & ~new_n38580_;
  assign new_n38582_ = ~new_n38571_ & ~new_n38581_;
  assign new_n38583_ = pi0211 & ~new_n38582_;
  assign new_n38584_ = ~pi0214 & ~new_n38582_;
  assign new_n38585_ = ~pi0212 & ~new_n38584_;
  assign new_n38586_ = new_n11383_ & new_n38531_;
  assign new_n38587_ = pi1153 & new_n38586_;
  assign new_n38588_ = pi1153 & ~new_n38556_;
  assign new_n38589_ = ~pi1153 & ~new_n10820_;
  assign new_n38590_ = ~new_n38588_ & ~new_n38589_;
  assign new_n38591_ = pi1155 & ~new_n38590_;
  assign new_n38592_ = ~new_n38587_ & ~new_n38591_;
  assign new_n38593_ = ~pi1154 & ~new_n38592_;
  assign new_n38594_ = pi1155 & ~new_n11383_;
  assign new_n38595_ = new_n38534_ & ~new_n38549_;
  assign new_n38596_ = ~new_n38594_ & ~new_n38595_;
  assign new_n38597_ = pi1154 & ~new_n38596_;
  assign new_n38598_ = ~new_n38593_ & ~new_n38597_;
  assign new_n38599_ = pi0207 & new_n38598_;
  assign new_n38600_ = ~pi0207 & ~new_n38510_;
  assign new_n38601_ = new_n38566_ & new_n38600_;
  assign new_n38602_ = pi0208 & ~new_n38601_;
  assign new_n38603_ = ~new_n38599_ & new_n38602_;
  assign new_n38604_ = pi1155 & ~new_n38556_;
  assign new_n38605_ = ~new_n11373_ & ~new_n38604_;
  assign new_n38606_ = pi1156 & ~new_n38605_;
  assign new_n38607_ = pi0199 & ~pi0200;
  assign new_n38608_ = ~pi0299 & ~new_n38607_;
  assign new_n38609_ = ~pi1155 & ~new_n38608_;
  assign new_n38610_ = ~pi1156 & ~new_n38556_;
  assign new_n38611_ = ~new_n38609_ & new_n38610_;
  assign new_n38612_ = ~new_n38606_ & ~new_n38611_;
  assign new_n38613_ = pi0207 & new_n38612_;
  assign new_n38614_ = ~pi0208 & ~new_n38600_;
  assign new_n38615_ = pi1157 & new_n38614_;
  assign new_n38616_ = ~new_n38613_ & new_n38615_;
  assign new_n38617_ = ~pi0299 & new_n38530_;
  assign new_n38618_ = ~pi0299 & ~new_n38533_;
  assign new_n38619_ = ~pi1155 & ~new_n11373_;
  assign new_n38620_ = ~new_n38618_ & ~new_n38619_;
  assign new_n38621_ = ~new_n38617_ & new_n38620_;
  assign new_n38622_ = new_n38614_ & new_n38621_;
  assign new_n38623_ = ~new_n38616_ & ~new_n38622_;
  assign new_n38624_ = ~new_n38603_ & new_n38623_;
  assign new_n38625_ = new_n38495_ & new_n38624_;
  assign new_n38626_ = new_n38585_ & ~new_n38625_;
  assign new_n38627_ = ~pi1155 & ~new_n10820_;
  assign new_n38628_ = ~new_n38604_ & ~new_n38627_;
  assign new_n38629_ = ~pi1156 & ~new_n38628_;
  assign new_n38630_ = new_n11383_ & ~new_n38527_;
  assign new_n38631_ = pi1156 & ~new_n38630_;
  assign new_n38632_ = ~new_n38629_ & ~new_n38631_;
  assign new_n38633_ = pi0207 & new_n38632_;
  assign new_n38634_ = ~pi0207 & ~pi0299;
  assign new_n38635_ = ~pi0208 & ~new_n38634_;
  assign new_n38636_ = ~new_n38633_ & new_n38635_;
  assign new_n38637_ = pi1157 & ~new_n38636_;
  assign new_n38638_ = ~pi0299 & ~new_n11444_;
  assign new_n38639_ = pi1156 & ~new_n38528_;
  assign new_n38640_ = new_n38638_ & new_n38639_;
  assign new_n38641_ = ~new_n38530_ & ~new_n38640_;
  assign new_n38642_ = pi0207 & new_n38641_;
  assign new_n38643_ = ~pi0299 & ~new_n38642_;
  assign new_n38644_ = ~pi0208 & ~new_n38643_;
  assign new_n38645_ = ~pi1157 & ~new_n38644_;
  assign new_n38646_ = pi0299 & ~pi1153;
  assign new_n38647_ = ~new_n38645_ & ~new_n38646_;
  assign new_n38648_ = ~new_n38637_ & new_n38647_;
  assign new_n38649_ = pi1153 & ~new_n38608_;
  assign new_n38650_ = new_n38546_ & ~new_n38649_;
  assign new_n38651_ = pi0207 & ~new_n38650_;
  assign new_n38652_ = ~new_n38594_ & ~new_n38627_;
  assign new_n38653_ = pi1156 & ~new_n38652_;
  assign new_n38654_ = pi1155 & ~new_n38618_;
  assign new_n38655_ = ~new_n38609_ & ~new_n38654_;
  assign new_n38656_ = pi1154 & ~new_n38655_;
  assign new_n38657_ = ~new_n38653_ & ~new_n38656_;
  assign new_n38658_ = pi0299 & ~pi1155;
  assign new_n38659_ = pi1155 & ~new_n38638_;
  assign new_n38660_ = ~new_n38658_ & ~new_n38659_;
  assign new_n38661_ = new_n38657_ & new_n38660_;
  assign new_n38662_ = ~pi0207 & ~new_n38646_;
  assign new_n38663_ = ~new_n38661_ & new_n38662_;
  assign new_n38664_ = ~new_n38651_ & ~new_n38663_;
  assign new_n38665_ = pi0208 & ~new_n38664_;
  assign new_n38666_ = new_n38495_ & ~new_n38665_;
  assign new_n38667_ = ~new_n38648_ & new_n38666_;
  assign new_n38668_ = ~pi0211 & ~pi0214;
  assign new_n38669_ = new_n38566_ & ~new_n38656_;
  assign new_n38670_ = ~pi0207 & ~new_n38669_;
  assign new_n38671_ = ~pi0299 & new_n38596_;
  assign new_n38672_ = pi1154 & ~new_n38671_;
  assign new_n38673_ = ~new_n38553_ & ~new_n38672_;
  assign new_n38674_ = pi0207 & ~new_n38673_;
  assign new_n38675_ = ~new_n38670_ & ~new_n38674_;
  assign new_n38676_ = pi0208 & ~new_n38675_;
  assign new_n38677_ = pi0299 & ~pi1154;
  assign new_n38678_ = pi1157 & ~new_n38677_;
  assign new_n38679_ = new_n38636_ & new_n38678_;
  assign new_n38680_ = ~new_n38512_ & ~new_n38537_;
  assign new_n38681_ = ~pi0208 & ~new_n38680_;
  assign new_n38682_ = ~pi1157 & new_n38681_;
  assign new_n38683_ = ~new_n38679_ & ~new_n38682_;
  assign new_n38684_ = ~new_n38676_ & new_n38683_;
  assign new_n38685_ = new_n38668_ & new_n38684_;
  assign new_n38686_ = pi0212 & ~new_n38685_;
  assign new_n38687_ = ~new_n38667_ & new_n38686_;
  assign new_n38688_ = ~new_n38626_ & ~new_n38687_;
  assign new_n38689_ = ~new_n38583_ & ~new_n38688_;
  assign new_n38690_ = pi0219 & ~new_n38689_;
  assign new_n38691_ = ~pi0207 & new_n38661_;
  assign new_n38692_ = new_n38442_ & new_n38650_;
  assign new_n38693_ = pi0208 & ~new_n38692_;
  assign new_n38694_ = ~new_n38691_ & new_n38693_;
  assign new_n38695_ = new_n38637_ & ~new_n38694_;
  assign new_n38696_ = ~pi0211 & ~new_n38695_;
  assign new_n38697_ = ~new_n38571_ & new_n38696_;
  assign new_n38698_ = pi0207 & ~new_n38554_;
  assign new_n38699_ = ~new_n38562_ & ~new_n38653_;
  assign new_n38700_ = ~pi0207 & ~new_n38699_;
  assign new_n38701_ = pi0299 & pi1156;
  assign new_n38702_ = pi0207 & new_n38701_;
  assign new_n38703_ = ~new_n38700_ & ~new_n38702_;
  assign new_n38704_ = ~new_n38698_ & new_n38703_;
  assign new_n38705_ = pi0208 & ~new_n38704_;
  assign new_n38706_ = ~new_n38530_ & new_n38644_;
  assign new_n38707_ = ~pi0208 & pi1157;
  assign new_n38708_ = ~new_n38578_ & ~new_n38701_;
  assign new_n38709_ = new_n38707_ & ~new_n38708_;
  assign new_n38710_ = ~new_n38706_ & ~new_n38709_;
  assign new_n38711_ = ~new_n38705_ & new_n38710_;
  assign new_n38712_ = pi0211 & ~new_n38711_;
  assign new_n38713_ = pi0214 & ~new_n38712_;
  assign new_n38714_ = ~new_n38697_ & new_n38713_;
  assign new_n38715_ = new_n38585_ & ~new_n38714_;
  assign new_n38716_ = new_n10484_ & ~new_n38684_;
  assign new_n38717_ = ~new_n10484_ & ~new_n38668_;
  assign new_n38718_ = ~new_n38624_ & new_n38717_;
  assign new_n38719_ = new_n38668_ & ~new_n38711_;
  assign new_n38720_ = ~new_n38718_ & ~new_n38719_;
  assign new_n38721_ = ~new_n38716_ & new_n38720_;
  assign new_n38722_ = pi0212 & ~new_n38721_;
  assign new_n38723_ = ~pi0219 & ~new_n38722_;
  assign new_n38724_ = ~new_n38715_ & new_n38723_;
  assign new_n38725_ = ~po1038 & ~new_n38724_;
  assign new_n38726_ = ~new_n38690_ & new_n38725_;
  assign new_n38727_ = new_n38507_ & ~new_n38726_;
  assign new_n38728_ = ~pi0211 & new_n10729_;
  assign new_n38729_ = pi0299 & ~pi1143;
  assign new_n38730_ = new_n38654_ & ~new_n38729_;
  assign new_n38731_ = pi0299 & pi1143;
  assign new_n38732_ = ~pi1155 & new_n38731_;
  assign new_n38733_ = pi1154 & ~new_n38586_;
  assign new_n38734_ = ~new_n38732_ & new_n38733_;
  assign new_n38735_ = ~new_n38730_ & new_n38734_;
  assign new_n38736_ = new_n38559_ & ~new_n38731_;
  assign new_n38737_ = ~pi1156 & ~new_n38736_;
  assign new_n38738_ = ~new_n38735_ & new_n38737_;
  assign new_n38739_ = ~new_n38652_ & ~new_n38729_;
  assign new_n38740_ = ~pi1154 & ~new_n38739_;
  assign new_n38741_ = ~pi0299 & ~new_n38560_;
  assign new_n38742_ = pi1154 & ~new_n38741_;
  assign new_n38743_ = ~new_n38731_ & new_n38742_;
  assign new_n38744_ = pi1156 & ~new_n38743_;
  assign new_n38745_ = ~new_n38740_ & new_n38744_;
  assign new_n38746_ = ~new_n38738_ & ~new_n38745_;
  assign new_n38747_ = ~pi0207 & new_n38746_;
  assign new_n38748_ = new_n38555_ & ~new_n38731_;
  assign new_n38749_ = pi0208 & ~new_n38748_;
  assign new_n38750_ = ~new_n38747_ & new_n38749_;
  assign new_n38751_ = ~pi1157 & new_n38644_;
  assign new_n38752_ = ~new_n38729_ & new_n38751_;
  assign new_n38753_ = ~new_n38574_ & new_n38628_;
  assign new_n38754_ = pi0207 & ~new_n38729_;
  assign new_n38755_ = ~new_n38753_ & new_n38754_;
  assign new_n38756_ = ~new_n38731_ & ~new_n38755_;
  assign new_n38757_ = new_n38707_ & ~new_n38756_;
  assign new_n38758_ = ~new_n38752_ & ~new_n38757_;
  assign new_n38759_ = ~new_n38750_ & new_n38758_;
  assign new_n38760_ = new_n38728_ & new_n38759_;
  assign new_n38761_ = pi0299 & ~pi1144;
  assign new_n38762_ = new_n38654_ & ~new_n38761_;
  assign new_n38763_ = pi0299 & pi1144;
  assign new_n38764_ = ~pi1155 & new_n38763_;
  assign new_n38765_ = new_n38733_ & ~new_n38764_;
  assign new_n38766_ = ~new_n38762_ & new_n38765_;
  assign new_n38767_ = new_n38559_ & ~new_n38763_;
  assign new_n38768_ = ~pi1156 & ~new_n38767_;
  assign new_n38769_ = ~new_n38766_ & new_n38768_;
  assign new_n38770_ = ~new_n38652_ & ~new_n38761_;
  assign new_n38771_ = ~pi1154 & ~new_n38770_;
  assign new_n38772_ = new_n38742_ & ~new_n38763_;
  assign new_n38773_ = pi1156 & ~new_n38772_;
  assign new_n38774_ = ~new_n38771_ & new_n38773_;
  assign new_n38775_ = ~new_n38769_ & ~new_n38774_;
  assign new_n38776_ = ~pi0207 & new_n38775_;
  assign new_n38777_ = new_n38555_ & ~new_n38763_;
  assign new_n38778_ = pi0208 & ~new_n38777_;
  assign new_n38779_ = ~new_n38776_ & new_n38778_;
  assign new_n38780_ = new_n38751_ & ~new_n38761_;
  assign new_n38781_ = pi0207 & ~new_n38761_;
  assign new_n38782_ = ~new_n38753_ & new_n38781_;
  assign new_n38783_ = ~new_n38763_ & ~new_n38782_;
  assign new_n38784_ = new_n38707_ & ~new_n38783_;
  assign new_n38785_ = ~new_n38780_ & ~new_n38784_;
  assign new_n38786_ = ~new_n38779_ & new_n38785_;
  assign new_n38787_ = ~pi0211 & ~new_n38786_;
  assign new_n38788_ = ~new_n10729_ & ~new_n38413_;
  assign new_n38789_ = pi0211 & ~new_n38759_;
  assign new_n38790_ = new_n38788_ & ~new_n38789_;
  assign new_n38791_ = ~new_n38787_ & new_n38790_;
  assign new_n38792_ = ~new_n38760_ & ~new_n38791_;
  assign new_n38793_ = ~pi0219 & ~new_n38792_;
  assign new_n38794_ = ~pi0219 & ~new_n38413_;
  assign new_n38795_ = ~new_n38414_ & ~new_n38794_;
  assign new_n38796_ = ~new_n38582_ & new_n38795_;
  assign new_n38797_ = ~pi0299 & ~new_n38598_;
  assign new_n38798_ = pi0299 & pi1142;
  assign new_n38799_ = pi0207 & ~new_n38798_;
  assign new_n38800_ = ~new_n38797_ & new_n38799_;
  assign new_n38801_ = ~new_n38468_ & ~new_n38657_;
  assign new_n38802_ = ~new_n38558_ & ~new_n38798_;
  assign new_n38803_ = ~pi1154 & ~pi1156;
  assign new_n38804_ = ~new_n38802_ & new_n38803_;
  assign new_n38805_ = ~pi0207 & ~new_n38804_;
  assign new_n38806_ = ~new_n38801_ & new_n38805_;
  assign new_n38807_ = pi0208 & ~new_n38806_;
  assign new_n38808_ = ~new_n38800_ & new_n38807_;
  assign new_n38809_ = ~new_n38468_ & ~new_n38645_;
  assign new_n38810_ = ~new_n38637_ & new_n38809_;
  assign new_n38811_ = ~new_n10486_ & ~new_n38795_;
  assign new_n38812_ = ~new_n38810_ & new_n38811_;
  assign new_n38813_ = ~new_n38808_ & new_n38812_;
  assign new_n38814_ = ~po1038 & ~new_n38813_;
  assign new_n38815_ = ~new_n38796_ & new_n38814_;
  assign new_n38816_ = ~new_n38793_ & new_n38815_;
  assign new_n38817_ = pi0213 & ~new_n38430_;
  assign new_n38818_ = ~new_n38816_ & new_n38817_;
  assign new_n38819_ = ~pi0209 & ~new_n38818_;
  assign new_n38820_ = ~new_n38727_ & new_n38819_;
  assign new_n38821_ = ~new_n38526_ & ~new_n38820_;
  assign new_n38822_ = pi0230 & ~new_n38821_;
  assign po0390 = new_n38412_ | new_n38822_;
  assign new_n38824_ = pi1153 & ~new_n38668_;
  assign new_n38825_ = ~new_n38495_ & ~new_n38499_;
  assign new_n38826_ = ~new_n38824_ & ~new_n38825_;
  assign new_n38827_ = pi0212 & ~new_n38826_;
  assign new_n38828_ = pi0211 & pi1153;
  assign new_n38829_ = ~new_n38498_ & ~new_n38828_;
  assign new_n38830_ = new_n38421_ & ~new_n38829_;
  assign new_n38831_ = ~pi0219 & ~new_n38830_;
  assign new_n38832_ = ~new_n38827_ & new_n38831_;
  assign new_n38833_ = new_n38416_ & ~new_n38832_;
  assign new_n38834_ = pi1152 & ~new_n38833_;
  assign new_n38835_ = ~new_n10624_ & new_n38566_;
  assign new_n38836_ = ~pi0207 & ~pi0208;
  assign new_n38837_ = ~new_n10624_ & ~new_n38836_;
  assign new_n38838_ = ~pi1154 & ~new_n38542_;
  assign new_n38839_ = ~pi0199 & new_n38531_;
  assign new_n38840_ = new_n38539_ & ~new_n38839_;
  assign new_n38841_ = ~new_n38838_ & new_n38840_;
  assign new_n38842_ = pi0207 & new_n38841_;
  assign new_n38843_ = ~new_n38837_ & ~new_n38842_;
  assign new_n38844_ = ~new_n38835_ & ~new_n38843_;
  assign new_n38845_ = ~pi0214 & ~new_n38844_;
  assign new_n38846_ = ~pi0212 & ~new_n38845_;
  assign new_n38847_ = ~pi0207 & new_n38512_;
  assign new_n38848_ = pi0207 & ~new_n38669_;
  assign new_n38849_ = ~new_n38847_ & ~new_n38848_;
  assign new_n38850_ = ~pi0208 & ~new_n38849_;
  assign new_n38851_ = ~pi1155 & new_n10817_;
  assign new_n38852_ = ~new_n38532_ & ~new_n38851_;
  assign new_n38853_ = ~pi0299 & ~new_n38852_;
  assign new_n38854_ = ~new_n38838_ & ~new_n38853_;
  assign new_n38855_ = pi0207 & new_n38854_;
  assign new_n38856_ = ~new_n38670_ & ~new_n38855_;
  assign new_n38857_ = pi0208 & ~new_n38856_;
  assign new_n38858_ = ~new_n38850_ & ~new_n38857_;
  assign new_n38859_ = ~pi0211 & ~new_n38858_;
  assign new_n38860_ = pi0207 & new_n38660_;
  assign new_n38861_ = new_n38657_ & new_n38860_;
  assign new_n38862_ = new_n38635_ & ~new_n38861_;
  assign new_n38863_ = new_n38442_ & ~new_n38854_;
  assign new_n38864_ = pi0208 & ~new_n38863_;
  assign new_n38865_ = ~new_n38691_ & new_n38864_;
  assign new_n38866_ = ~new_n38862_ & ~new_n38865_;
  assign new_n38867_ = ~new_n38646_ & ~new_n38866_;
  assign new_n38868_ = pi0211 & new_n38867_;
  assign new_n38869_ = ~new_n38859_ & ~new_n38868_;
  assign new_n38870_ = pi0214 & new_n38869_;
  assign new_n38871_ = new_n38846_ & ~new_n38870_;
  assign new_n38872_ = ~pi0219 & ~new_n38871_;
  assign new_n38873_ = ~pi0214 & ~new_n38869_;
  assign new_n38874_ = ~pi0211 & ~new_n38867_;
  assign new_n38875_ = pi0214 & ~new_n38874_;
  assign new_n38876_ = ~new_n38866_ & new_n38875_;
  assign new_n38877_ = ~new_n38873_ & ~new_n38876_;
  assign new_n38878_ = pi0212 & ~new_n38877_;
  assign new_n38879_ = new_n38872_ & ~new_n38878_;
  assign new_n38880_ = ~new_n38414_ & new_n38844_;
  assign new_n38881_ = pi0219 & ~new_n38880_;
  assign new_n38882_ = new_n38414_ & ~new_n38866_;
  assign new_n38883_ = new_n38881_ & ~new_n38882_;
  assign new_n38884_ = ~po1038 & ~new_n38883_;
  assign new_n38885_ = ~new_n38879_ & new_n38884_;
  assign new_n38886_ = new_n38834_ & ~new_n38885_;
  assign new_n38887_ = ~new_n10729_ & new_n38829_;
  assign new_n38888_ = new_n38794_ & ~new_n38887_;
  assign new_n38889_ = ~new_n38501_ & new_n38888_;
  assign new_n38890_ = po1038 & new_n38889_;
  assign new_n38891_ = ~pi1152 & ~new_n38890_;
  assign new_n38892_ = pi0211 & ~new_n38844_;
  assign new_n38893_ = new_n38875_ & ~new_n38892_;
  assign new_n38894_ = ~new_n38873_ & ~new_n38893_;
  assign new_n38895_ = pi0212 & ~new_n38894_;
  assign new_n38896_ = new_n38872_ & ~new_n38895_;
  assign new_n38897_ = pi0219 & ~new_n38844_;
  assign new_n38898_ = ~po1038 & ~new_n38897_;
  assign new_n38899_ = ~new_n38896_ & new_n38898_;
  assign new_n38900_ = new_n38891_ & ~new_n38899_;
  assign new_n38901_ = ~pi0213 & ~new_n38900_;
  assign new_n38902_ = ~new_n38886_ & new_n38901_;
  assign new_n38903_ = pi0207 & ~new_n38699_;
  assign new_n38904_ = ~new_n38701_ & ~new_n38903_;
  assign new_n38905_ = ~pi0208 & ~new_n38904_;
  assign new_n38906_ = new_n38703_ & ~new_n38842_;
  assign new_n38907_ = pi0208 & ~new_n38906_;
  assign new_n38908_ = ~new_n38905_ & ~new_n38907_;
  assign new_n38909_ = ~pi0211 & ~new_n38908_;
  assign new_n38910_ = ~new_n38510_ & new_n38566_;
  assign new_n38911_ = new_n38614_ & ~new_n38910_;
  assign new_n38912_ = pi0207 & ~new_n38510_;
  assign new_n38913_ = ~new_n38841_ & new_n38912_;
  assign new_n38914_ = pi0208 & ~new_n38913_;
  assign new_n38915_ = ~new_n38601_ & new_n38914_;
  assign new_n38916_ = ~new_n38911_ & ~new_n38915_;
  assign new_n38917_ = pi0211 & ~new_n38916_;
  assign new_n38918_ = ~new_n38909_ & ~new_n38917_;
  assign new_n38919_ = ~pi0214 & new_n38918_;
  assign new_n38920_ = pi0211 & ~new_n38858_;
  assign new_n38921_ = ~pi0211 & ~new_n38916_;
  assign new_n38922_ = pi0214 & ~new_n38921_;
  assign new_n38923_ = ~new_n38920_ & new_n38922_;
  assign new_n38924_ = pi0212 & ~new_n38923_;
  assign new_n38925_ = ~new_n38919_ & new_n38924_;
  assign new_n38926_ = pi0214 & new_n38918_;
  assign new_n38927_ = new_n38846_ & ~new_n38926_;
  assign new_n38928_ = ~pi0219 & ~new_n38927_;
  assign new_n38929_ = ~new_n38925_ & new_n38928_;
  assign new_n38930_ = ~new_n38413_ & new_n38859_;
  assign new_n38931_ = new_n38881_ & ~new_n38930_;
  assign new_n38932_ = new_n35819_ & ~new_n38931_;
  assign new_n38933_ = ~new_n38929_ & new_n38932_;
  assign new_n38934_ = pi0209 & ~new_n38933_;
  assign new_n38935_ = ~new_n38902_ & new_n38934_;
  assign new_n38936_ = ~pi0199 & pi1153;
  assign new_n38937_ = pi0200 & new_n38936_;
  assign new_n38938_ = ~pi0299 & new_n38937_;
  assign new_n38939_ = ~pi1154 & ~new_n38938_;
  assign new_n38940_ = pi1154 & new_n38556_;
  assign new_n38941_ = ~new_n38936_ & new_n38940_;
  assign new_n38942_ = ~new_n38939_ & ~new_n38941_;
  assign new_n38943_ = new_n38608_ & ~new_n38942_;
  assign new_n38944_ = new_n38635_ & ~new_n38943_;
  assign new_n38945_ = ~pi0207 & new_n38943_;
  assign new_n38946_ = ~pi0200 & ~pi1153;
  assign new_n38947_ = ~pi0199 & ~new_n38946_;
  assign new_n38948_ = ~pi0299 & ~new_n38947_;
  assign new_n38949_ = ~new_n38607_ & new_n38948_;
  assign new_n38950_ = pi0207 & new_n38949_;
  assign new_n38951_ = pi0208 & ~new_n38950_;
  assign new_n38952_ = ~new_n38945_ & new_n38951_;
  assign new_n38953_ = ~new_n38944_ & ~new_n38952_;
  assign new_n38954_ = ~pi0211 & new_n38953_;
  assign new_n38955_ = ~pi0299 & new_n10817_;
  assign new_n38956_ = ~pi1153 & ~new_n38955_;
  assign new_n38957_ = new_n38541_ & ~new_n38956_;
  assign new_n38958_ = ~pi0199 & ~pi1153;
  assign new_n38959_ = new_n38534_ & ~new_n38958_;
  assign new_n38960_ = ~new_n38957_ & ~new_n38959_;
  assign new_n38961_ = ~new_n10624_ & new_n38960_;
  assign new_n38962_ = ~pi1153 & new_n10817_;
  assign new_n38963_ = new_n38539_ & ~new_n38962_;
  assign new_n38964_ = new_n10624_ & ~new_n38963_;
  assign new_n38965_ = ~new_n38836_ & ~new_n38964_;
  assign new_n38966_ = ~new_n38961_ & new_n38965_;
  assign new_n38967_ = pi0211 & ~new_n38966_;
  assign new_n38968_ = ~new_n38954_ & ~new_n38967_;
  assign new_n38969_ = ~new_n38413_ & new_n38968_;
  assign new_n38970_ = pi0219 & ~new_n38413_;
  assign new_n38971_ = pi0219 & ~new_n38966_;
  assign new_n38972_ = ~new_n38970_ & ~new_n38971_;
  assign new_n38973_ = ~new_n38969_ & ~new_n38972_;
  assign new_n38974_ = ~po1038 & ~new_n38973_;
  assign new_n38975_ = ~pi0214 & ~new_n38966_;
  assign new_n38976_ = ~pi0212 & ~new_n38975_;
  assign new_n38977_ = pi0207 & ~new_n38960_;
  assign new_n38978_ = ~new_n38512_ & ~new_n38977_;
  assign new_n38979_ = ~pi0208 & ~new_n38978_;
  assign new_n38980_ = pi0207 & ~new_n38949_;
  assign new_n38981_ = ~new_n38677_ & new_n38980_;
  assign new_n38982_ = pi1154 & ~new_n10820_;
  assign new_n38983_ = ~new_n38957_ & ~new_n38982_;
  assign new_n38984_ = ~new_n38959_ & new_n38983_;
  assign new_n38985_ = ~pi0207 & ~new_n38984_;
  assign new_n38986_ = ~new_n38981_ & ~new_n38985_;
  assign new_n38987_ = pi0208 & ~new_n38986_;
  assign new_n38988_ = ~new_n38979_ & ~new_n38987_;
  assign new_n38989_ = ~pi0211 & ~new_n38988_;
  assign new_n38990_ = ~pi0207 & new_n38514_;
  assign new_n38991_ = ~pi1153 & ~new_n38548_;
  assign new_n38992_ = ~new_n38618_ & ~new_n38991_;
  assign new_n38993_ = pi1154 & ~new_n11383_;
  assign new_n38994_ = ~new_n38991_ & new_n38993_;
  assign new_n38995_ = ~new_n38992_ & ~new_n38994_;
  assign new_n38996_ = pi0207 & ~new_n38995_;
  assign new_n38997_ = ~new_n38990_ & ~new_n38996_;
  assign new_n38998_ = ~pi0208 & ~new_n38997_;
  assign new_n38999_ = ~pi0207 & ~new_n38995_;
  assign new_n39000_ = ~pi0299 & new_n38532_;
  assign new_n39001_ = pi0207 & ~new_n39000_;
  assign new_n39002_ = ~new_n38589_ & new_n39001_;
  assign new_n39003_ = ~new_n38999_ & ~new_n39002_;
  assign new_n39004_ = pi0208 & ~new_n39003_;
  assign new_n39005_ = ~new_n38998_ & ~new_n39004_;
  assign new_n39006_ = pi0211 & ~new_n39005_;
  assign new_n39007_ = ~new_n38989_ & ~new_n39006_;
  assign new_n39008_ = pi0214 & new_n39007_;
  assign new_n39009_ = new_n38976_ & ~new_n39008_;
  assign new_n39010_ = ~pi0214 & new_n39007_;
  assign new_n39011_ = pi0211 & ~new_n38953_;
  assign new_n39012_ = ~pi0211 & ~new_n39005_;
  assign new_n39013_ = pi0214 & ~new_n39012_;
  assign new_n39014_ = ~new_n39011_ & new_n39013_;
  assign new_n39015_ = pi0212 & ~new_n39014_;
  assign new_n39016_ = ~new_n39010_ & new_n39015_;
  assign new_n39017_ = ~pi0219 & ~new_n39016_;
  assign new_n39018_ = ~new_n39009_ & new_n39017_;
  assign new_n39019_ = new_n38974_ & ~new_n39018_;
  assign new_n39020_ = new_n38834_ & ~new_n39019_;
  assign new_n39021_ = pi1153 & ~pi1154;
  assign new_n39022_ = ~new_n38638_ & new_n39021_;
  assign new_n39023_ = ~new_n38994_ & ~new_n39022_;
  assign new_n39024_ = pi0207 & ~new_n39023_;
  assign new_n39025_ = ~new_n38990_ & ~new_n39024_;
  assign new_n39026_ = ~pi0208 & ~new_n39025_;
  assign new_n39027_ = ~pi0207 & ~new_n39023_;
  assign new_n39028_ = pi0207 & ~new_n10820_;
  assign new_n39029_ = pi1153 & new_n39028_;
  assign new_n39030_ = ~new_n39027_ & ~new_n39029_;
  assign new_n39031_ = pi0208 & ~new_n39030_;
  assign new_n39032_ = ~new_n39026_ & ~new_n39031_;
  assign new_n39033_ = new_n38728_ & new_n39032_;
  assign new_n39034_ = pi1153 & ~new_n11383_;
  assign new_n39035_ = ~new_n38589_ & ~new_n39034_;
  assign new_n39036_ = pi1154 & ~new_n39035_;
  assign new_n39037_ = ~new_n38938_ & ~new_n39036_;
  assign new_n39038_ = pi0207 & ~new_n39037_;
  assign new_n39039_ = ~new_n38847_ & ~new_n39038_;
  assign new_n39040_ = ~pi0208 & ~new_n39039_;
  assign new_n39041_ = ~pi0207 & new_n39037_;
  assign new_n39042_ = ~pi0299 & ~pi1153;
  assign new_n39043_ = ~new_n10820_ & ~new_n39042_;
  assign new_n39044_ = ~new_n38677_ & new_n39043_;
  assign new_n39045_ = pi0207 & ~new_n39044_;
  assign new_n39046_ = pi0208 & ~new_n39045_;
  assign new_n39047_ = ~new_n39041_ & new_n39046_;
  assign new_n39048_ = ~new_n39040_ & ~new_n39047_;
  assign new_n39049_ = ~pi0211 & new_n39048_;
  assign new_n39050_ = pi0211 & new_n39032_;
  assign new_n39051_ = ~new_n39049_ & ~new_n39050_;
  assign new_n39052_ = new_n38788_ & ~new_n39051_;
  assign new_n39053_ = ~new_n39033_ & ~new_n39052_;
  assign new_n39054_ = ~pi0219 & ~new_n39053_;
  assign new_n39055_ = pi0200 & ~pi1153;
  assign new_n39056_ = new_n11373_ & ~new_n39055_;
  assign new_n39057_ = pi1154 & ~new_n39056_;
  assign new_n39058_ = ~new_n38939_ & ~new_n39057_;
  assign new_n39059_ = new_n38837_ & new_n39058_;
  assign new_n39060_ = pi0208 & new_n38442_;
  assign new_n39061_ = pi1153 & ~new_n10820_;
  assign new_n39062_ = new_n39060_ & new_n39061_;
  assign new_n39063_ = ~new_n39059_ & ~new_n39062_;
  assign new_n39064_ = pi0219 & new_n39063_;
  assign new_n39065_ = ~po1038 & ~new_n39064_;
  assign new_n39066_ = ~new_n38495_ & ~new_n38788_;
  assign new_n39067_ = new_n39063_ & new_n39066_;
  assign new_n39068_ = new_n39065_ & ~new_n39067_;
  assign new_n39069_ = ~new_n39054_ & new_n39068_;
  assign new_n39070_ = new_n38891_ & ~new_n39069_;
  assign new_n39071_ = ~new_n39020_ & ~new_n39070_;
  assign new_n39072_ = ~pi0213 & new_n39071_;
  assign new_n39073_ = ~pi1152 & ~po1038;
  assign new_n39074_ = pi0211 & new_n39048_;
  assign new_n39075_ = ~pi0299 & ~new_n38937_;
  assign new_n39076_ = ~pi1154 & ~new_n39075_;
  assign new_n39077_ = ~new_n38658_ & new_n39076_;
  assign new_n39078_ = ~new_n38619_ & new_n39036_;
  assign new_n39079_ = ~new_n39077_ & ~new_n39078_;
  assign new_n39080_ = pi0207 & new_n39079_;
  assign new_n39081_ = new_n38614_ & ~new_n39080_;
  assign new_n39082_ = ~pi0207 & new_n39079_;
  assign new_n39083_ = ~new_n38658_ & new_n39043_;
  assign new_n39084_ = pi0207 & ~new_n39083_;
  assign new_n39085_ = pi0208 & ~new_n39084_;
  assign new_n39086_ = ~new_n39082_ & new_n39085_;
  assign new_n39087_ = ~new_n39081_ & ~new_n39086_;
  assign new_n39088_ = ~pi0211 & new_n39087_;
  assign new_n39089_ = new_n10729_ & ~new_n39088_;
  assign new_n39090_ = ~new_n39074_ & new_n39089_;
  assign new_n39091_ = pi0211 & new_n39087_;
  assign new_n39092_ = ~pi0211 & ~new_n38701_;
  assign new_n39093_ = new_n39063_ & new_n39092_;
  assign new_n39094_ = ~new_n38423_ & ~new_n39093_;
  assign new_n39095_ = ~new_n39091_ & new_n39094_;
  assign new_n39096_ = ~new_n39090_ & ~new_n39095_;
  assign new_n39097_ = ~pi0219 & ~new_n39096_;
  assign new_n39098_ = new_n38413_ & ~new_n39063_;
  assign new_n39099_ = pi0211 & new_n39063_;
  assign new_n39100_ = new_n38970_ & ~new_n39099_;
  assign new_n39101_ = ~new_n39049_ & new_n39100_;
  assign new_n39102_ = ~new_n39098_ & ~new_n39101_;
  assign new_n39103_ = ~new_n39097_ & new_n39102_;
  assign new_n39104_ = new_n39073_ & ~new_n39103_;
  assign new_n39105_ = ~new_n38414_ & new_n38966_;
  assign new_n39106_ = ~new_n38413_ & new_n38989_;
  assign new_n39107_ = ~new_n39105_ & ~new_n39106_;
  assign new_n39108_ = pi0219 & ~new_n39107_;
  assign new_n39109_ = pi0211 & ~new_n38988_;
  assign new_n39110_ = new_n38614_ & ~new_n38943_;
  assign new_n39111_ = ~new_n38952_ & ~new_n39110_;
  assign new_n39112_ = ~pi0199 & ~pi1154;
  assign new_n39113_ = ~pi0200 & new_n39112_;
  assign new_n39114_ = new_n38634_ & new_n39113_;
  assign new_n39115_ = ~new_n38658_ & ~new_n39114_;
  assign new_n39116_ = ~new_n39111_ & new_n39115_;
  assign new_n39117_ = ~pi0211 & new_n39116_;
  assign new_n39118_ = new_n10729_ & ~new_n39117_;
  assign new_n39119_ = ~new_n39109_ & new_n39118_;
  assign new_n39120_ = pi0211 & new_n39116_;
  assign new_n39121_ = ~new_n38701_ & new_n38960_;
  assign new_n39122_ = ~pi0207 & ~new_n39121_;
  assign new_n39123_ = pi0299 & ~pi1156;
  assign new_n39124_ = new_n38980_ & ~new_n39123_;
  assign new_n39125_ = pi0208 & ~new_n39124_;
  assign new_n39126_ = ~new_n39122_ & new_n39125_;
  assign new_n39127_ = ~pi0208 & ~new_n38701_;
  assign new_n39128_ = ~new_n38977_ & new_n39127_;
  assign new_n39129_ = ~pi0211 & ~new_n39128_;
  assign new_n39130_ = ~new_n39126_ & new_n39129_;
  assign new_n39131_ = ~new_n38423_ & ~new_n39130_;
  assign new_n39132_ = ~new_n39120_ & new_n39131_;
  assign new_n39133_ = ~pi0212 & new_n38975_;
  assign new_n39134_ = ~pi0219 & ~new_n39133_;
  assign new_n39135_ = ~new_n39132_ & new_n39134_;
  assign new_n39136_ = ~new_n39119_ & new_n39135_;
  assign new_n39137_ = ~new_n39108_ & ~new_n39136_;
  assign new_n39138_ = pi1152 & ~po1038;
  assign new_n39139_ = ~new_n39137_ & new_n39138_;
  assign new_n39140_ = ~new_n39104_ & ~new_n39139_;
  assign new_n39141_ = pi0213 & ~new_n39140_;
  assign new_n39142_ = ~pi0209 & ~new_n39141_;
  assign new_n39143_ = ~new_n39072_ & new_n39142_;
  assign new_n39144_ = ~new_n38935_ & ~new_n39143_;
  assign new_n39145_ = pi0212 & ~new_n38491_;
  assign new_n39146_ = pi0214 & ~new_n38485_;
  assign new_n39147_ = ~pi0212 & new_n39146_;
  assign new_n39148_ = ~pi0219 & ~new_n39147_;
  assign new_n39149_ = ~new_n39145_ & new_n39148_;
  assign new_n39150_ = pi0219 & ~new_n38498_;
  assign new_n39151_ = pi0213 & ~new_n39150_;
  assign new_n39152_ = new_n38416_ & new_n39151_;
  assign new_n39153_ = ~new_n39149_ & new_n39152_;
  assign new_n39154_ = ~new_n39144_ & ~new_n39153_;
  assign new_n39155_ = pi0230 & ~new_n39154_;
  assign new_n39156_ = ~pi0230 & pi0234;
  assign po0391 = new_n39155_ | new_n39156_;
  assign new_n39158_ = ~pi1156 & new_n38558_;
  assign new_n39159_ = ~new_n38653_ & ~new_n39158_;
  assign new_n39160_ = pi0207 & ~new_n39159_;
  assign new_n39161_ = ~pi0207 & new_n38641_;
  assign new_n39162_ = ~new_n39160_ & ~new_n39161_;
  assign new_n39163_ = pi0208 & ~new_n39162_;
  assign new_n39164_ = ~new_n38706_ & ~new_n39163_;
  assign new_n39165_ = ~pi1157 & ~new_n39164_;
  assign new_n39166_ = pi0208 & pi1157;
  assign new_n39167_ = ~new_n38576_ & ~new_n38631_;
  assign new_n39168_ = ~pi0207 & ~new_n39167_;
  assign new_n39169_ = ~new_n39160_ & ~new_n39168_;
  assign new_n39170_ = new_n39166_ & ~new_n39169_;
  assign new_n39171_ = ~new_n38709_ & ~new_n39170_;
  assign new_n39172_ = ~new_n39165_ & new_n39171_;
  assign new_n39173_ = ~pi0211 & ~new_n39172_;
  assign new_n39174_ = ~new_n38565_ & ~new_n38659_;
  assign new_n39175_ = pi0207 & ~new_n39174_;
  assign new_n39176_ = ~pi0207 & new_n38621_;
  assign new_n39177_ = ~new_n39175_ & ~new_n39176_;
  assign new_n39178_ = pi0208 & ~new_n39177_;
  assign new_n39179_ = ~new_n38622_ & ~new_n39178_;
  assign new_n39180_ = ~pi1157 & ~new_n39179_;
  assign new_n39181_ = ~pi0207 & ~new_n38612_;
  assign new_n39182_ = ~new_n39175_ & ~new_n39181_;
  assign new_n39183_ = new_n39166_ & ~new_n39182_;
  assign new_n39184_ = ~new_n38616_ & ~new_n39183_;
  assign new_n39185_ = ~new_n39180_ & new_n39184_;
  assign new_n39186_ = pi0211 & ~new_n39185_;
  assign new_n39187_ = new_n10729_ & ~new_n39186_;
  assign new_n39188_ = ~new_n39173_ & new_n39187_;
  assign new_n39189_ = new_n10624_ & ~new_n38565_;
  assign new_n39190_ = ~new_n39158_ & new_n39189_;
  assign new_n39191_ = ~pi0207 & ~new_n38536_;
  assign new_n39192_ = ~new_n39190_ & ~new_n39191_;
  assign new_n39193_ = ~new_n38538_ & new_n39192_;
  assign new_n39194_ = ~pi1157 & ~new_n39193_;
  assign new_n39195_ = ~pi0207 & new_n38577_;
  assign new_n39196_ = ~new_n39190_ & ~new_n39195_;
  assign new_n39197_ = ~new_n38579_ & new_n39196_;
  assign new_n39198_ = pi1157 & ~new_n39197_;
  assign new_n39199_ = ~new_n39194_ & ~new_n39198_;
  assign new_n39200_ = new_n38413_ & ~new_n39199_;
  assign new_n39201_ = pi0211 & ~new_n39172_;
  assign new_n39202_ = ~pi0207 & new_n38632_;
  assign new_n39203_ = pi0208 & ~new_n39202_;
  assign new_n39204_ = ~new_n38653_ & new_n38860_;
  assign new_n39205_ = new_n39203_ & ~new_n39204_;
  assign new_n39206_ = ~new_n38636_ & ~new_n39205_;
  assign new_n39207_ = pi1157 & new_n39206_;
  assign new_n39208_ = ~pi0211 & ~new_n39194_;
  assign new_n39209_ = ~new_n39207_ & new_n39208_;
  assign new_n39210_ = new_n38788_ & ~new_n39209_;
  assign new_n39211_ = ~new_n39201_ & new_n39210_;
  assign new_n39212_ = ~new_n39200_ & ~new_n39211_;
  assign new_n39213_ = ~new_n39188_ & new_n39212_;
  assign new_n39214_ = ~pi0219 & ~new_n39213_;
  assign new_n39215_ = ~pi0211 & new_n39185_;
  assign new_n39216_ = pi0211 & ~new_n39199_;
  assign new_n39217_ = ~new_n38423_ & ~new_n39216_;
  assign new_n39218_ = ~new_n39215_ & new_n39217_;
  assign new_n39219_ = new_n38423_ & new_n39199_;
  assign new_n39220_ = pi0219 & ~new_n39219_;
  assign new_n39221_ = ~new_n39218_ & new_n39220_;
  assign new_n39222_ = pi0209 & ~new_n39221_;
  assign new_n39223_ = ~new_n39214_ & new_n39222_;
  assign new_n39224_ = new_n10624_ & ~new_n39058_;
  assign new_n39225_ = ~new_n38554_ & ~new_n38836_;
  assign new_n39226_ = ~new_n10624_ & ~new_n39225_;
  assign new_n39227_ = ~new_n39224_ & ~new_n39226_;
  assign new_n39228_ = ~pi1157 & new_n39227_;
  assign new_n39229_ = new_n38635_ & ~new_n38692_;
  assign new_n39230_ = ~new_n39036_ & ~new_n39076_;
  assign new_n39231_ = pi0207 & new_n39230_;
  assign new_n39232_ = new_n38634_ & new_n38650_;
  assign new_n39233_ = pi0208 & ~new_n39232_;
  assign new_n39234_ = ~new_n39231_ & new_n39233_;
  assign new_n39235_ = ~new_n39229_ & ~new_n39234_;
  assign new_n39236_ = pi1157 & ~new_n39235_;
  assign new_n39237_ = ~pi0211 & ~new_n39236_;
  assign new_n39238_ = ~new_n39228_ & new_n39237_;
  assign new_n39239_ = ~new_n38701_ & ~new_n39227_;
  assign new_n39240_ = pi0211 & new_n39239_;
  assign new_n39241_ = ~new_n39238_ & ~new_n39240_;
  assign new_n39242_ = new_n38788_ & ~new_n39241_;
  assign new_n39243_ = ~pi0211 & ~new_n39239_;
  assign new_n39244_ = ~new_n38598_ & new_n38614_;
  assign new_n39245_ = ~pi0207 & new_n38598_;
  assign new_n39246_ = pi0208 & ~new_n39080_;
  assign new_n39247_ = ~new_n39245_ & new_n39246_;
  assign new_n39248_ = ~new_n39244_ & ~new_n39247_;
  assign new_n39249_ = pi0211 & ~new_n39248_;
  assign new_n39250_ = new_n10729_ & ~new_n39249_;
  assign new_n39251_ = ~new_n39243_ & new_n39250_;
  assign new_n39252_ = new_n38413_ & ~new_n39227_;
  assign new_n39253_ = ~new_n39251_ & ~new_n39252_;
  assign new_n39254_ = ~new_n39242_ & new_n39253_;
  assign new_n39255_ = ~pi0219 & ~new_n39254_;
  assign new_n39256_ = ~pi0211 & new_n39248_;
  assign new_n39257_ = pi0211 & ~new_n39227_;
  assign new_n39258_ = ~new_n38423_ & ~new_n39257_;
  assign new_n39259_ = ~new_n39256_ & new_n39258_;
  assign new_n39260_ = new_n38423_ & new_n39227_;
  assign new_n39261_ = pi0219 & ~new_n39260_;
  assign new_n39262_ = ~new_n39259_ & new_n39261_;
  assign new_n39263_ = ~pi0209 & ~new_n39262_;
  assign new_n39264_ = ~new_n39255_ & new_n39263_;
  assign new_n39265_ = ~new_n39223_ & ~new_n39264_;
  assign new_n39266_ = ~po1038 & ~new_n39265_;
  assign new_n39267_ = ~pi0212 & new_n38481_;
  assign new_n39268_ = ~pi0214 & ~new_n38480_;
  assign new_n39269_ = ~new_n39146_ & ~new_n39268_;
  assign new_n39270_ = pi0212 & ~new_n39269_;
  assign new_n39271_ = ~pi0219 & ~new_n39270_;
  assign new_n39272_ = ~new_n39267_ & new_n39271_;
  assign new_n39273_ = pi0219 & ~new_n38487_;
  assign new_n39274_ = pi0219 & ~new_n38788_;
  assign new_n39275_ = ~new_n39273_ & ~new_n39274_;
  assign new_n39276_ = po1038 & new_n39275_;
  assign new_n39277_ = ~new_n39272_ & new_n39276_;
  assign new_n39278_ = pi0213 & ~new_n39277_;
  assign new_n39279_ = ~new_n39266_ & new_n39278_;
  assign new_n39280_ = pi1157 & ~new_n39206_;
  assign new_n39281_ = pi0299 & ~pi1157;
  assign new_n39282_ = ~new_n39165_ & ~new_n39281_;
  assign new_n39283_ = ~new_n39280_ & new_n39282_;
  assign new_n39284_ = ~new_n38646_ & ~new_n39283_;
  assign new_n39285_ = ~pi0211 & ~new_n39284_;
  assign new_n39286_ = new_n39217_ & ~new_n39285_;
  assign new_n39287_ = new_n39220_ & ~new_n39286_;
  assign new_n39288_ = pi0211 & new_n39284_;
  assign new_n39289_ = ~new_n38559_ & ~new_n38660_;
  assign new_n39290_ = ~new_n38565_ & ~new_n39289_;
  assign new_n39291_ = pi0207 & ~new_n39290_;
  assign new_n39292_ = pi1154 & ~new_n38640_;
  assign new_n39293_ = ~new_n38535_ & ~new_n39292_;
  assign new_n39294_ = ~pi0207 & ~new_n38617_;
  assign new_n39295_ = ~new_n39293_ & new_n39294_;
  assign new_n39296_ = ~new_n39291_ & ~new_n39295_;
  assign new_n39297_ = pi0208 & ~new_n39296_;
  assign new_n39298_ = ~new_n38681_ & ~new_n39297_;
  assign new_n39299_ = ~pi1157 & ~new_n39298_;
  assign new_n39300_ = new_n38678_ & ~new_n39206_;
  assign new_n39301_ = ~new_n39299_ & ~new_n39300_;
  assign new_n39302_ = ~pi0211 & ~new_n39301_;
  assign new_n39303_ = new_n10729_ & ~new_n39302_;
  assign new_n39304_ = ~new_n39288_ & new_n39303_;
  assign new_n39305_ = pi0211 & new_n39301_;
  assign new_n39306_ = ~new_n39215_ & ~new_n39305_;
  assign new_n39307_ = new_n38788_ & ~new_n39306_;
  assign new_n39308_ = ~new_n39200_ & ~new_n39307_;
  assign new_n39309_ = ~new_n39304_ & new_n39308_;
  assign new_n39310_ = ~pi0219 & ~new_n39309_;
  assign new_n39311_ = ~new_n39287_ & ~new_n39310_;
  assign new_n39312_ = pi0209 & ~new_n39311_;
  assign new_n39313_ = ~new_n38651_ & ~new_n38990_;
  assign new_n39314_ = ~pi0208 & ~new_n39313_;
  assign new_n39315_ = ~pi0207 & ~new_n38650_;
  assign new_n39316_ = ~new_n39024_ & ~new_n39315_;
  assign new_n39317_ = pi0208 & ~new_n39316_;
  assign new_n39318_ = ~new_n39314_ & ~new_n39317_;
  assign new_n39319_ = ~pi0211 & new_n39318_;
  assign new_n39320_ = new_n39258_ & ~new_n39319_;
  assign new_n39321_ = new_n39261_ & ~new_n39320_;
  assign new_n39322_ = ~new_n38674_ & ~new_n38847_;
  assign new_n39323_ = ~pi0208 & ~new_n39322_;
  assign new_n39324_ = ~pi0207 & ~new_n38673_;
  assign new_n39325_ = ~new_n39038_ & ~new_n39324_;
  assign new_n39326_ = pi0208 & ~new_n39325_;
  assign new_n39327_ = ~new_n39323_ & ~new_n39326_;
  assign new_n39328_ = pi0211 & new_n39327_;
  assign new_n39329_ = ~new_n39256_ & ~new_n39328_;
  assign new_n39330_ = ~new_n38423_ & ~new_n39329_;
  assign new_n39331_ = ~pi0211 & ~new_n39327_;
  assign new_n39332_ = pi0211 & ~new_n39318_;
  assign new_n39333_ = new_n10729_ & ~new_n39332_;
  assign new_n39334_ = ~new_n39331_ & new_n39333_;
  assign new_n39335_ = ~new_n39252_ & ~new_n39334_;
  assign new_n39336_ = ~new_n39330_ & new_n39335_;
  assign new_n39337_ = ~pi0219 & ~new_n39336_;
  assign new_n39338_ = ~new_n39321_ & ~new_n39337_;
  assign new_n39339_ = ~pi0209 & ~new_n39338_;
  assign new_n39340_ = ~po1038 & ~new_n39339_;
  assign new_n39341_ = ~new_n39312_ & new_n39340_;
  assign new_n39342_ = new_n10729_ & ~new_n38829_;
  assign new_n39343_ = ~new_n38489_ & new_n38788_;
  assign new_n39344_ = ~pi0219 & ~new_n39343_;
  assign new_n39345_ = ~new_n39342_ & new_n39344_;
  assign new_n39346_ = pi0219 & ~new_n38500_;
  assign new_n39347_ = po1038 & ~new_n39346_;
  assign new_n39348_ = ~new_n39274_ & new_n39347_;
  assign new_n39349_ = ~new_n39345_ & new_n39348_;
  assign new_n39350_ = ~pi0213 & ~new_n39349_;
  assign new_n39351_ = ~new_n39341_ & new_n39350_;
  assign new_n39352_ = ~new_n39279_ & ~new_n39351_;
  assign new_n39353_ = pi0230 & ~new_n39352_;
  assign new_n39354_ = ~pi0230 & ~pi0235;
  assign po0392 = ~new_n39353_ & ~new_n39354_;
  assign new_n39356_ = ~pi0100 & new_n38186_;
  assign new_n39357_ = new_n38397_ & ~new_n39356_;
  assign new_n39358_ = ~new_n6288_ & ~new_n39357_;
  assign new_n39359_ = ~pi0075 & ~new_n39358_;
  assign new_n39360_ = ~new_n7302_ & ~new_n39359_;
  assign new_n39361_ = ~pi0092 & ~new_n39360_;
  assign new_n39362_ = new_n13654_ & ~new_n39361_;
  assign new_n39363_ = ~pi0074 & ~new_n39362_;
  assign new_n39364_ = new_n6131_ & ~new_n39363_;
  assign new_n39365_ = ~pi0056 & ~new_n39364_;
  assign new_n39366_ = ~new_n6127_ & ~new_n39365_;
  assign new_n39367_ = ~pi0062 & ~new_n39366_;
  assign po0393 = new_n13662_ & ~new_n39367_;
  assign new_n39369_ = ~pi0211 & pi1145;
  assign new_n39370_ = pi0211 & pi1144;
  assign new_n39371_ = ~new_n39369_ & ~new_n39370_;
  assign new_n39372_ = ~new_n10729_ & new_n39371_;
  assign new_n39373_ = new_n10729_ & new_n38420_;
  assign new_n39374_ = ~new_n38413_ & ~new_n39373_;
  assign new_n39375_ = ~new_n39372_ & new_n39374_;
  assign new_n39376_ = ~pi0219 & ~new_n39375_;
  assign new_n39377_ = pi0219 & ~new_n38425_;
  assign new_n39378_ = new_n38416_ & ~new_n39377_;
  assign new_n39379_ = ~new_n39376_ & new_n39378_;
  assign new_n39380_ = new_n38508_ & new_n39375_;
  assign new_n39381_ = pi0199 & pi1143;
  assign new_n39382_ = ~pi0200 & ~new_n39381_;
  assign new_n39383_ = ~new_n38434_ & new_n39382_;
  assign new_n39384_ = ~new_n38437_ & new_n39060_;
  assign new_n39385_ = ~new_n39383_ & new_n39384_;
  assign new_n39386_ = ~pi0199 & pi1145;
  assign new_n39387_ = new_n39382_ & ~new_n39386_;
  assign new_n39388_ = pi0200 & ~new_n38434_;
  assign new_n39389_ = new_n38837_ & ~new_n39388_;
  assign new_n39390_ = ~new_n39387_ & new_n39389_;
  assign new_n39391_ = ~new_n39385_ & ~new_n39390_;
  assign new_n39392_ = ~pi0299 & ~new_n39391_;
  assign new_n39393_ = pi0299 & new_n38970_;
  assign new_n39394_ = new_n38425_ & new_n39393_;
  assign new_n39395_ = ~new_n39392_ & ~new_n39394_;
  assign new_n39396_ = ~new_n39380_ & new_n39395_;
  assign new_n39397_ = ~po1038 & ~new_n39396_;
  assign new_n39398_ = ~new_n39379_ & ~new_n39397_;
  assign new_n39399_ = pi0213 & new_n39398_;
  assign new_n39400_ = pi0211 & pi1157;
  assign new_n39401_ = ~pi0211 & pi1158;
  assign new_n39402_ = ~new_n39400_ & ~new_n39401_;
  assign new_n39403_ = new_n38421_ & ~new_n39402_;
  assign new_n39404_ = new_n39271_ & ~new_n39403_;
  assign new_n39405_ = ~pi0219 & po1038;
  assign new_n39406_ = new_n38421_ & new_n38483_;
  assign new_n39407_ = po1038 & new_n39406_;
  assign new_n39408_ = ~new_n39405_ & ~new_n39407_;
  assign new_n39409_ = pi0214 & new_n38498_;
  assign new_n39410_ = pi1155 & new_n38668_;
  assign new_n39411_ = ~new_n39409_ & ~new_n39410_;
  assign new_n39412_ = pi0212 & ~new_n39411_;
  assign new_n39413_ = po1038 & new_n39412_;
  assign new_n39414_ = new_n39408_ & ~new_n39413_;
  assign new_n39415_ = ~new_n39404_ & ~new_n39414_;
  assign new_n39416_ = ~pi0213 & ~new_n39415_;
  assign new_n39417_ = new_n38508_ & ~new_n39404_;
  assign new_n39418_ = new_n38421_ & new_n38701_;
  assign new_n39419_ = ~pi0214 & ~new_n38510_;
  assign new_n39420_ = pi0214 & ~new_n38512_;
  assign new_n39421_ = pi0212 & ~new_n39420_;
  assign new_n39422_ = ~new_n39419_ & new_n39421_;
  assign new_n39423_ = ~new_n39418_ & ~new_n39422_;
  assign new_n39424_ = new_n38519_ & ~new_n39423_;
  assign new_n39425_ = ~new_n39392_ & ~new_n39424_;
  assign new_n39426_ = ~new_n39417_ & new_n39425_;
  assign new_n39427_ = ~po1038 & ~new_n39426_;
  assign new_n39428_ = new_n39416_ & ~new_n39427_;
  assign new_n39429_ = pi0209 & ~new_n39428_;
  assign new_n39430_ = ~new_n39399_ & new_n39429_;
  assign new_n39431_ = new_n38449_ & new_n38548_;
  assign new_n39432_ = pi1158 & new_n38955_;
  assign new_n39433_ = ~pi0199 & ~pi1158;
  assign new_n39434_ = pi1156 & ~new_n39433_;
  assign new_n39435_ = ~new_n39432_ & ~new_n39434_;
  assign new_n39436_ = new_n39431_ & ~new_n39435_;
  assign new_n39437_ = pi0207 & new_n38566_;
  assign new_n39438_ = pi0208 & ~new_n39191_;
  assign new_n39439_ = ~new_n39437_ & new_n39438_;
  assign new_n39440_ = ~new_n39436_ & ~new_n39439_;
  assign new_n39441_ = ~pi1157 & ~new_n39440_;
  assign new_n39442_ = pi1156 & new_n38607_;
  assign new_n39443_ = ~pi0200 & ~pi1158;
  assign new_n39444_ = ~pi0199 & ~new_n39443_;
  assign new_n39445_ = ~new_n39442_ & ~new_n39444_;
  assign new_n39446_ = new_n38442_ & ~new_n39445_;
  assign new_n39447_ = ~pi0208 & new_n39446_;
  assign new_n39448_ = pi0208 & ~new_n39195_;
  assign new_n39449_ = ~new_n39437_ & new_n39448_;
  assign new_n39450_ = ~new_n39447_ & ~new_n39449_;
  assign new_n39451_ = pi1157 & ~new_n39450_;
  assign new_n39452_ = ~new_n39441_ & ~new_n39451_;
  assign new_n39453_ = ~pi0214 & new_n39452_;
  assign new_n39454_ = ~pi0212 & ~new_n39453_;
  assign new_n39455_ = ~pi0299 & new_n39445_;
  assign new_n39456_ = new_n38635_ & ~new_n39455_;
  assign new_n39457_ = ~new_n38861_ & new_n39203_;
  assign new_n39458_ = ~new_n39456_ & ~new_n39457_;
  assign new_n39459_ = pi1157 & ~new_n39458_;
  assign new_n39460_ = ~new_n39441_ & ~new_n39459_;
  assign new_n39461_ = pi0211 & new_n39460_;
  assign new_n39462_ = pi1158 & new_n38661_;
  assign new_n39463_ = ~pi1158 & new_n38566_;
  assign new_n39464_ = pi0207 & ~new_n39463_;
  assign new_n39465_ = ~new_n39462_ & new_n39464_;
  assign new_n39466_ = ~pi0207 & ~new_n38632_;
  assign new_n39467_ = pi0299 & ~pi1158;
  assign new_n39468_ = new_n39466_ & ~new_n39467_;
  assign new_n39469_ = ~new_n39465_ & ~new_n39468_;
  assign new_n39470_ = new_n39166_ & ~new_n39469_;
  assign new_n39471_ = ~pi0299 & ~new_n38641_;
  assign new_n39472_ = ~pi0207 & ~new_n39467_;
  assign new_n39473_ = ~new_n39471_ & new_n39472_;
  assign new_n39474_ = pi0208 & ~new_n39473_;
  assign new_n39475_ = ~new_n39465_ & new_n39474_;
  assign new_n39476_ = ~pi0299 & ~new_n39028_;
  assign new_n39477_ = pi1158 & ~new_n39476_;
  assign new_n39478_ = new_n38442_ & new_n39442_;
  assign new_n39479_ = ~pi0208 & ~new_n39478_;
  assign new_n39480_ = ~new_n39477_ & new_n39479_;
  assign new_n39481_ = ~pi1157 & ~new_n39480_;
  assign new_n39482_ = ~new_n39475_ & new_n39481_;
  assign new_n39483_ = new_n38534_ & ~new_n38610_;
  assign new_n39484_ = pi1157 & ~new_n39432_;
  assign new_n39485_ = ~new_n39483_ & new_n39484_;
  assign new_n39486_ = pi0207 & ~new_n39485_;
  assign new_n39487_ = ~new_n39477_ & ~new_n39486_;
  assign new_n39488_ = new_n38707_ & ~new_n39487_;
  assign new_n39489_ = ~pi0211 & ~new_n39488_;
  assign new_n39490_ = ~new_n39482_ & new_n39489_;
  assign new_n39491_ = ~new_n39470_ & new_n39490_;
  assign new_n39492_ = ~new_n39461_ & ~new_n39491_;
  assign new_n39493_ = pi0214 & ~new_n39492_;
  assign new_n39494_ = new_n39454_ & ~new_n39493_;
  assign new_n39495_ = new_n38668_ & ~new_n39460_;
  assign new_n39496_ = pi0208 & ~new_n39161_;
  assign new_n39497_ = ~new_n38903_ & new_n39496_;
  assign new_n39498_ = ~pi0200 & pi0207;
  assign new_n39499_ = ~new_n39435_ & new_n39498_;
  assign new_n39500_ = new_n39127_ & ~new_n39499_;
  assign new_n39501_ = ~pi1157 & ~new_n39500_;
  assign new_n39502_ = ~new_n39497_ & new_n39501_;
  assign new_n39503_ = ~new_n38903_ & ~new_n39168_;
  assign new_n39504_ = new_n39166_ & ~new_n39503_;
  assign new_n39505_ = ~new_n38701_ & ~new_n39446_;
  assign new_n39506_ = new_n38707_ & ~new_n39505_;
  assign new_n39507_ = ~new_n39504_ & ~new_n39506_;
  assign new_n39508_ = ~new_n39502_ & new_n39507_;
  assign new_n39509_ = new_n38717_ & ~new_n39508_;
  assign new_n39510_ = pi0207 & ~new_n38910_;
  assign new_n39511_ = ~new_n39176_ & ~new_n39510_;
  assign new_n39512_ = pi0208 & ~new_n39511_;
  assign new_n39513_ = ~pi0208 & new_n38510_;
  assign new_n39514_ = ~new_n39436_ & ~new_n39513_;
  assign new_n39515_ = ~new_n39512_ & new_n39514_;
  assign new_n39516_ = ~pi1157 & ~new_n39515_;
  assign new_n39517_ = ~new_n39181_ & ~new_n39510_;
  assign new_n39518_ = new_n39166_ & ~new_n39517_;
  assign new_n39519_ = pi1156 & ~new_n39000_;
  assign new_n39520_ = ~pi1158 & ~new_n38534_;
  assign new_n39521_ = new_n39519_ & ~new_n39520_;
  assign new_n39522_ = ~new_n39444_ & ~new_n39521_;
  assign new_n39523_ = new_n38442_ & ~new_n39522_;
  assign new_n39524_ = ~new_n38510_ & ~new_n39523_;
  assign new_n39525_ = new_n38707_ & ~new_n39524_;
  assign new_n39526_ = ~new_n39518_ & ~new_n39525_;
  assign new_n39527_ = ~new_n39516_ & new_n39526_;
  assign new_n39528_ = new_n10484_ & ~new_n39527_;
  assign new_n39529_ = ~new_n39509_ & ~new_n39528_;
  assign new_n39530_ = ~new_n39495_ & new_n39529_;
  assign new_n39531_ = pi0212 & ~new_n39530_;
  assign new_n39532_ = ~pi0219 & ~new_n39531_;
  assign new_n39533_ = ~new_n39494_ & new_n39532_;
  assign new_n39534_ = ~new_n38414_ & new_n39452_;
  assign new_n39535_ = new_n38421_ & new_n39508_;
  assign new_n39536_ = ~pi0214 & ~new_n39527_;
  assign new_n39537_ = ~new_n38677_ & new_n39466_;
  assign new_n39538_ = pi1157 & ~new_n39537_;
  assign new_n39539_ = ~pi1157 & ~new_n39436_;
  assign new_n39540_ = ~new_n39295_ & new_n39539_;
  assign new_n39541_ = ~new_n39538_ & ~new_n39540_;
  assign new_n39542_ = pi0208 & ~new_n38848_;
  assign new_n39543_ = ~new_n39541_ & new_n39542_;
  assign new_n39544_ = new_n39523_ & ~new_n39539_;
  assign new_n39545_ = ~pi0208 & ~new_n38512_;
  assign new_n39546_ = ~new_n39544_ & new_n39545_;
  assign new_n39547_ = pi0214 & ~new_n39546_;
  assign new_n39548_ = ~new_n39543_ & new_n39547_;
  assign new_n39549_ = pi0212 & ~new_n39548_;
  assign new_n39550_ = ~new_n39536_ & new_n39549_;
  assign new_n39551_ = ~new_n39535_ & ~new_n39550_;
  assign new_n39552_ = ~pi0211 & ~new_n39551_;
  assign new_n39553_ = ~new_n39534_ & ~new_n39552_;
  assign new_n39554_ = pi0219 & ~new_n39553_;
  assign new_n39555_ = ~po1038 & ~new_n39554_;
  assign new_n39556_ = ~new_n39533_ & new_n39555_;
  assign new_n39557_ = new_n39416_ & ~new_n39556_;
  assign new_n39558_ = pi0299 & ~pi1145;
  assign new_n39559_ = ~new_n38655_ & ~new_n39558_;
  assign new_n39560_ = pi1154 & ~new_n39559_;
  assign new_n39561_ = pi0299 & pi1145;
  assign new_n39562_ = new_n38559_ & ~new_n39561_;
  assign new_n39563_ = ~pi1156 & ~new_n39562_;
  assign new_n39564_ = ~new_n39560_ & new_n39563_;
  assign new_n39565_ = ~new_n38652_ & ~new_n39558_;
  assign new_n39566_ = ~pi1154 & ~new_n39565_;
  assign new_n39567_ = new_n38742_ & ~new_n39561_;
  assign new_n39568_ = pi1156 & ~new_n39567_;
  assign new_n39569_ = ~new_n39566_ & new_n39568_;
  assign new_n39570_ = ~new_n39564_ & ~new_n39569_;
  assign new_n39571_ = pi0207 & ~new_n39570_;
  assign new_n39572_ = ~pi0200 & pi1157;
  assign new_n39573_ = ~pi0199 & new_n39572_;
  assign new_n39574_ = new_n39471_ & ~new_n39573_;
  assign new_n39575_ = ~pi0207 & ~new_n39558_;
  assign new_n39576_ = ~new_n39574_ & new_n39575_;
  assign new_n39577_ = pi0208 & ~new_n39576_;
  assign new_n39578_ = ~new_n39571_ & new_n39577_;
  assign new_n39579_ = ~pi0299 & new_n39442_;
  assign new_n39580_ = ~pi1157 & ~new_n39432_;
  assign new_n39581_ = ~new_n39579_ & new_n39580_;
  assign new_n39582_ = new_n39486_ & ~new_n39581_;
  assign new_n39583_ = ~pi0208 & ~new_n39561_;
  assign new_n39584_ = ~new_n39582_ & new_n39583_;
  assign new_n39585_ = ~new_n39578_ & ~new_n39584_;
  assign new_n39586_ = ~pi0211 & ~new_n39585_;
  assign new_n39587_ = ~pi1157 & ~new_n39499_;
  assign new_n39588_ = ~pi0208 & ~new_n39587_;
  assign new_n39589_ = new_n39523_ & new_n39588_;
  assign new_n39590_ = ~pi0208 & ~new_n39589_;
  assign new_n39591_ = ~new_n38763_ & new_n39590_;
  assign new_n39592_ = pi0207 & ~new_n38775_;
  assign new_n39593_ = ~pi0207 & ~new_n38761_;
  assign new_n39594_ = ~new_n39574_ & new_n39593_;
  assign new_n39595_ = pi0208 & ~new_n39594_;
  assign new_n39596_ = ~new_n39592_ & new_n39595_;
  assign new_n39597_ = ~new_n39591_ & ~new_n39596_;
  assign new_n39598_ = pi0211 & ~new_n39597_;
  assign new_n39599_ = ~new_n39586_ & ~new_n39598_;
  assign new_n39600_ = ~pi0214 & ~new_n39599_;
  assign new_n39601_ = ~new_n38731_ & new_n39590_;
  assign new_n39602_ = pi0207 & ~new_n38746_;
  assign new_n39603_ = ~pi0207 & ~new_n38729_;
  assign new_n39604_ = ~new_n39574_ & new_n39603_;
  assign new_n39605_ = pi0208 & ~new_n39604_;
  assign new_n39606_ = ~new_n39602_ & new_n39605_;
  assign new_n39607_ = ~new_n39601_ & ~new_n39606_;
  assign new_n39608_ = pi0211 & new_n39607_;
  assign new_n39609_ = ~pi0211 & new_n39597_;
  assign new_n39610_ = pi0214 & ~new_n39609_;
  assign new_n39611_ = ~new_n39608_ & new_n39610_;
  assign new_n39612_ = pi0212 & ~new_n39611_;
  assign new_n39613_ = ~new_n39600_ & new_n39612_;
  assign new_n39614_ = pi0214 & ~new_n39599_;
  assign new_n39615_ = new_n39454_ & ~new_n39614_;
  assign new_n39616_ = ~pi0219 & ~new_n39615_;
  assign new_n39617_ = ~new_n39613_ & new_n39616_;
  assign new_n39618_ = new_n38414_ & ~new_n39607_;
  assign new_n39619_ = ~new_n39534_ & ~new_n39618_;
  assign new_n39620_ = pi0219 & ~new_n39619_;
  assign new_n39621_ = ~po1038 & ~new_n39620_;
  assign new_n39622_ = ~new_n39617_ & new_n39621_;
  assign new_n39623_ = pi0213 & ~new_n39379_;
  assign new_n39624_ = ~new_n39622_ & new_n39623_;
  assign new_n39625_ = ~pi0209 & ~new_n39624_;
  assign new_n39626_ = ~new_n39557_ & new_n39625_;
  assign new_n39627_ = ~new_n39430_ & ~new_n39626_;
  assign new_n39628_ = pi0230 & ~new_n39627_;
  assign new_n39629_ = ~pi0230 & ~pi0237;
  assign po0394 = new_n39628_ | new_n39629_;
  assign new_n39631_ = ~pi0211 & ~pi1153;
  assign new_n39632_ = pi0219 & new_n39631_;
  assign new_n39633_ = new_n38416_ & ~new_n39632_;
  assign new_n39634_ = ~new_n39345_ & new_n39633_;
  assign new_n39635_ = ~new_n10624_ & new_n38548_;
  assign new_n39636_ = ~new_n38836_ & new_n39635_;
  assign new_n39637_ = new_n38533_ & new_n39060_;
  assign new_n39638_ = ~new_n39636_ & ~new_n39637_;
  assign new_n39639_ = ~new_n38962_ & ~new_n39638_;
  assign new_n39640_ = ~pi0214 & ~new_n39639_;
  assign new_n39641_ = ~pi0212 & ~new_n39640_;
  assign new_n39642_ = new_n38548_ & ~new_n38958_;
  assign new_n39643_ = ~pi1153 & ~new_n38608_;
  assign new_n39644_ = ~new_n38588_ & ~new_n39643_;
  assign new_n39645_ = pi1155 & ~new_n39644_;
  assign new_n39646_ = ~new_n39642_ & ~new_n39645_;
  assign new_n39647_ = new_n38442_ & ~new_n38533_;
  assign new_n39648_ = pi0208 & ~new_n39647_;
  assign new_n39649_ = ~new_n38614_ & ~new_n39648_;
  assign new_n39650_ = ~new_n39646_ & ~new_n39649_;
  assign new_n39651_ = ~new_n39637_ & ~new_n39650_;
  assign new_n39652_ = ~pi0299 & ~new_n39651_;
  assign new_n39653_ = pi0299 & ~new_n38489_;
  assign new_n39654_ = pi0214 & ~new_n39653_;
  assign new_n39655_ = ~new_n39652_ & new_n39654_;
  assign new_n39656_ = new_n39641_ & ~new_n39655_;
  assign new_n39657_ = new_n38668_ & new_n39651_;
  assign new_n39658_ = ~pi0299 & ~new_n39498_;
  assign new_n39659_ = ~pi0208 & ~new_n39658_;
  assign new_n39660_ = pi0200 & new_n38634_;
  assign new_n39661_ = new_n39648_ & ~new_n39660_;
  assign new_n39662_ = ~new_n39659_ & ~new_n39661_;
  assign new_n39663_ = ~new_n38589_ & ~new_n39662_;
  assign new_n39664_ = new_n10484_ & ~new_n39663_;
  assign new_n39665_ = ~new_n38512_ & new_n38717_;
  assign new_n39666_ = ~new_n39639_ & new_n39665_;
  assign new_n39667_ = pi0212 & ~new_n39666_;
  assign new_n39668_ = ~new_n39664_ & new_n39667_;
  assign new_n39669_ = ~new_n39657_ & new_n39668_;
  assign new_n39670_ = ~pi0219 & ~new_n39669_;
  assign new_n39671_ = ~new_n39656_ & new_n39670_;
  assign new_n39672_ = pi1151 & ~po1038;
  assign new_n39673_ = ~pi0211 & ~new_n39662_;
  assign new_n39674_ = pi0211 & ~new_n39638_;
  assign new_n39675_ = ~new_n39673_ & ~new_n39674_;
  assign new_n39676_ = ~new_n38589_ & ~new_n39675_;
  assign new_n39677_ = new_n38413_ & ~new_n39639_;
  assign new_n39678_ = new_n39676_ & ~new_n39677_;
  assign new_n39679_ = pi0219 & ~new_n39678_;
  assign new_n39680_ = new_n39672_ & ~new_n39679_;
  assign new_n39681_ = ~new_n39671_ & new_n39680_;
  assign new_n39682_ = new_n38837_ & new_n38955_;
  assign new_n39683_ = pi1153 & new_n39682_;
  assign new_n39684_ = ~new_n38512_ & ~new_n39683_;
  assign new_n39685_ = ~pi0211 & ~new_n39684_;
  assign new_n39686_ = new_n10817_ & new_n38837_;
  assign new_n39687_ = ~pi0299 & ~new_n39686_;
  assign new_n39688_ = new_n38828_ & ~new_n39687_;
  assign new_n39689_ = new_n10729_ & ~new_n39688_;
  assign new_n39690_ = ~new_n39685_ & new_n39689_;
  assign new_n39691_ = ~new_n38423_ & ~new_n39653_;
  assign new_n39692_ = ~new_n39683_ & new_n39691_;
  assign new_n39693_ = ~new_n39690_ & ~new_n39692_;
  assign new_n39694_ = ~pi0219 & ~new_n39693_;
  assign new_n39695_ = ~pi1151 & ~po1038;
  assign new_n39696_ = ~new_n13061_ & ~new_n39687_;
  assign new_n39697_ = ~pi0214 & ~new_n39682_;
  assign new_n39698_ = ~pi0212 & new_n39697_;
  assign new_n39699_ = new_n39696_ & ~new_n39698_;
  assign new_n39700_ = pi1153 & new_n39699_;
  assign new_n39701_ = ~new_n38794_ & ~new_n39700_;
  assign new_n39702_ = new_n39695_ & ~new_n39701_;
  assign new_n39703_ = ~new_n39694_ & new_n39702_;
  assign new_n39704_ = ~pi1152 & ~new_n39703_;
  assign new_n39705_ = ~new_n39681_ & new_n39704_;
  assign new_n39706_ = ~new_n11445_ & ~new_n39034_;
  assign new_n39707_ = pi0207 & ~new_n39706_;
  assign new_n39708_ = ~new_n38990_ & ~new_n39707_;
  assign new_n39709_ = ~pi0208 & ~new_n39708_;
  assign new_n39710_ = pi0200 & pi0207;
  assign new_n39711_ = ~pi0199 & ~new_n39710_;
  assign new_n39712_ = ~pi0299 & ~new_n39711_;
  assign new_n39713_ = pi0208 & ~new_n39712_;
  assign new_n39714_ = ~pi0207 & new_n10817_;
  assign new_n39715_ = ~pi0299 & ~new_n39714_;
  assign new_n39716_ = ~pi1153 & ~new_n39715_;
  assign new_n39717_ = new_n39713_ & ~new_n39716_;
  assign new_n39718_ = ~new_n39709_ & ~new_n39717_;
  assign new_n39719_ = pi0211 & ~new_n39718_;
  assign new_n39720_ = ~pi0207 & ~new_n38948_;
  assign new_n39721_ = ~new_n39028_ & ~new_n39720_;
  assign new_n39722_ = pi0208 & ~new_n39721_;
  assign new_n39723_ = new_n38635_ & ~new_n38948_;
  assign new_n39724_ = ~new_n39722_ & ~new_n39723_;
  assign new_n39725_ = ~pi0211 & ~new_n38677_;
  assign new_n39726_ = ~new_n39724_ & new_n39725_;
  assign new_n39727_ = ~new_n39719_ & ~new_n39726_;
  assign new_n39728_ = new_n10729_ & ~new_n39727_;
  assign new_n39729_ = pi0299 & new_n38489_;
  assign new_n39730_ = ~new_n38423_ & ~new_n39724_;
  assign new_n39731_ = ~new_n39729_ & new_n39730_;
  assign new_n39732_ = ~new_n39728_ & ~new_n39731_;
  assign new_n39733_ = ~pi0219 & ~new_n39732_;
  assign new_n39734_ = ~new_n10624_ & new_n38946_;
  assign new_n39735_ = ~new_n38837_ & ~new_n39498_;
  assign new_n39736_ = new_n11373_ & ~new_n39735_;
  assign new_n39737_ = ~new_n39734_ & new_n39736_;
  assign new_n39738_ = ~pi0211 & new_n38514_;
  assign new_n39739_ = ~new_n38413_ & new_n39738_;
  assign new_n39740_ = ~new_n39737_ & ~new_n39739_;
  assign new_n39741_ = ~new_n38794_ & ~new_n39740_;
  assign new_n39742_ = ~new_n39733_ & ~new_n39741_;
  assign new_n39743_ = new_n39695_ & ~new_n39742_;
  assign new_n39744_ = new_n38949_ & ~new_n39001_;
  assign new_n39745_ = pi0208 & ~new_n39744_;
  assign new_n39746_ = new_n38635_ & ~new_n38950_;
  assign new_n39747_ = ~new_n39745_ & ~new_n39746_;
  assign new_n39748_ = ~pi0211 & ~new_n39747_;
  assign new_n39749_ = ~new_n38658_ & new_n39748_;
  assign new_n39750_ = pi0211 & ~new_n39747_;
  assign new_n39751_ = ~new_n38677_ & new_n39750_;
  assign new_n39752_ = ~new_n39749_ & ~new_n39751_;
  assign new_n39753_ = ~new_n38423_ & ~new_n39752_;
  assign new_n39754_ = new_n38442_ & new_n38533_;
  assign new_n39755_ = pi0208 & new_n38539_;
  assign new_n39756_ = ~new_n39714_ & new_n39755_;
  assign new_n39757_ = ~new_n39754_ & ~new_n39756_;
  assign new_n39758_ = ~new_n39688_ & new_n39757_;
  assign new_n39759_ = ~new_n39726_ & new_n39758_;
  assign new_n39760_ = new_n10729_ & ~new_n39759_;
  assign new_n39761_ = ~pi0214 & new_n39757_;
  assign new_n39762_ = ~new_n39683_ & new_n39761_;
  assign new_n39763_ = ~pi0212 & ~new_n39762_;
  assign new_n39764_ = ~pi0214 & new_n39763_;
  assign new_n39765_ = ~pi0219 & ~new_n39764_;
  assign new_n39766_ = ~new_n39760_ & new_n39765_;
  assign new_n39767_ = ~new_n39753_ & new_n39766_;
  assign new_n39768_ = pi0219 & new_n39757_;
  assign new_n39769_ = ~new_n39700_ & new_n39768_;
  assign new_n39770_ = new_n39672_ & ~new_n39769_;
  assign new_n39771_ = ~new_n39767_ & new_n39770_;
  assign new_n39772_ = pi1152 & ~new_n39771_;
  assign new_n39773_ = ~new_n39743_ & new_n39772_;
  assign new_n39774_ = ~new_n39705_ & ~new_n39773_;
  assign new_n39775_ = ~pi0209 & ~new_n39774_;
  assign new_n39776_ = new_n38534_ & new_n39021_;
  assign new_n39777_ = new_n38983_ & ~new_n39776_;
  assign new_n39778_ = pi0207 & ~new_n39777_;
  assign new_n39779_ = ~new_n39324_ & ~new_n39778_;
  assign new_n39780_ = pi0208 & ~new_n39779_;
  assign new_n39781_ = ~new_n39323_ & ~new_n39780_;
  assign new_n39782_ = pi0211 & ~new_n39781_;
  assign new_n39783_ = ~new_n38539_ & new_n39084_;
  assign new_n39784_ = ~pi1154 & ~new_n39042_;
  assign new_n39785_ = ~new_n38618_ & new_n39784_;
  assign new_n39786_ = pi0207 & ~new_n39785_;
  assign new_n39787_ = new_n38983_ & new_n39786_;
  assign new_n39788_ = pi0208 & ~new_n39787_;
  assign new_n39789_ = ~new_n39783_ & new_n39788_;
  assign new_n39790_ = ~new_n39245_ & new_n39789_;
  assign new_n39791_ = ~new_n39244_ & ~new_n39790_;
  assign new_n39792_ = ~pi0211 & ~new_n39791_;
  assign new_n39793_ = new_n38421_ & ~new_n39792_;
  assign new_n39794_ = ~new_n39782_ & new_n39793_;
  assign new_n39795_ = new_n38717_ & ~new_n39781_;
  assign new_n39796_ = new_n38668_ & ~new_n39791_;
  assign new_n39797_ = pi1153 & ~new_n38618_;
  assign new_n39798_ = ~new_n38957_ & ~new_n39797_;
  assign new_n39799_ = pi0207 & ~new_n39798_;
  assign new_n39800_ = ~new_n39315_ & ~new_n39799_;
  assign new_n39801_ = pi0208 & ~new_n39800_;
  assign new_n39802_ = ~new_n39314_ & ~new_n39801_;
  assign new_n39803_ = new_n10484_ & ~new_n39802_;
  assign new_n39804_ = pi0212 & ~new_n39803_;
  assign new_n39805_ = ~new_n39796_ & new_n39804_;
  assign new_n39806_ = ~new_n39795_ & new_n39805_;
  assign new_n39807_ = ~new_n39794_ & ~new_n39806_;
  assign new_n39808_ = ~pi0219 & ~new_n39807_;
  assign new_n39809_ = new_n10624_ & ~new_n39776_;
  assign new_n39810_ = ~new_n38957_ & new_n39809_;
  assign new_n39811_ = ~new_n39226_ & ~new_n39810_;
  assign new_n39812_ = pi0211 & new_n39811_;
  assign new_n39813_ = ~pi0211 & ~new_n39802_;
  assign new_n39814_ = ~new_n39812_ & ~new_n39813_;
  assign new_n39815_ = new_n38970_ & new_n39814_;
  assign new_n39816_ = ~pi0214 & ~new_n39811_;
  assign new_n39817_ = ~pi0212 & new_n39816_;
  assign new_n39818_ = ~po1038 & ~new_n39817_;
  assign new_n39819_ = ~new_n39815_ & new_n39818_;
  assign new_n39820_ = ~new_n39808_ & new_n39819_;
  assign new_n39821_ = pi0209 & ~new_n39820_;
  assign new_n39822_ = ~new_n39775_ & ~new_n39821_;
  assign new_n39823_ = ~new_n39634_ & ~new_n39822_;
  assign new_n39824_ = pi0213 & ~new_n39823_;
  assign new_n39825_ = ~new_n10485_ & new_n38794_;
  assign new_n39826_ = po1038 & new_n39825_;
  assign new_n39827_ = ~new_n10729_ & ~new_n39631_;
  assign new_n39828_ = ~new_n38728_ & ~new_n39827_;
  assign new_n39829_ = new_n39826_ & ~new_n39828_;
  assign new_n39830_ = ~new_n10486_ & new_n38416_;
  assign new_n39831_ = pi1151 & ~new_n39830_;
  assign new_n39832_ = ~new_n39829_ & new_n39831_;
  assign new_n39833_ = ~new_n39232_ & new_n39788_;
  assign new_n39834_ = ~new_n39229_ & ~new_n39833_;
  assign new_n39835_ = ~pi0211 & ~new_n39834_;
  assign new_n39836_ = ~new_n39812_ & ~new_n39835_;
  assign new_n39837_ = ~new_n38413_ & new_n39836_;
  assign new_n39838_ = ~new_n39817_ & ~new_n39837_;
  assign new_n39839_ = pi0219 & ~new_n39838_;
  assign new_n39840_ = ~po1038 & ~new_n39839_;
  assign new_n39841_ = pi0211 & ~new_n39834_;
  assign new_n39842_ = ~new_n39813_ & ~new_n39841_;
  assign new_n39843_ = pi0214 & new_n39842_;
  assign new_n39844_ = ~pi0212 & ~new_n39816_;
  assign new_n39845_ = ~new_n39843_ & new_n39844_;
  assign new_n39846_ = ~pi0219 & ~new_n39845_;
  assign new_n39847_ = ~pi0214 & ~new_n39842_;
  assign new_n39848_ = pi0214 & ~new_n39834_;
  assign new_n39849_ = ~new_n39847_ & ~new_n39848_;
  assign new_n39850_ = pi0212 & ~new_n39849_;
  assign new_n39851_ = new_n39846_ & ~new_n39850_;
  assign new_n39852_ = new_n39840_ & ~new_n39851_;
  assign new_n39853_ = new_n39832_ & ~new_n39852_;
  assign new_n39854_ = ~pi1151 & ~new_n39829_;
  assign new_n39855_ = pi0214 & ~new_n39836_;
  assign new_n39856_ = ~new_n39847_ & ~new_n39855_;
  assign new_n39857_ = pi0212 & ~new_n39856_;
  assign new_n39858_ = new_n39846_ & ~new_n39857_;
  assign new_n39859_ = pi0219 & ~new_n39811_;
  assign new_n39860_ = ~po1038 & ~new_n39859_;
  assign new_n39861_ = ~new_n39858_ & new_n39860_;
  assign new_n39862_ = new_n39854_ & ~new_n39861_;
  assign new_n39863_ = pi1152 & ~new_n39862_;
  assign new_n39864_ = ~new_n39853_ & new_n39863_;
  assign new_n39865_ = ~pi0211 & new_n38788_;
  assign new_n39866_ = pi1153 & new_n39865_;
  assign new_n39867_ = new_n10486_ & ~new_n39866_;
  assign new_n39868_ = new_n38416_ & ~new_n39867_;
  assign new_n39869_ = pi1151 & ~new_n39868_;
  assign new_n39870_ = pi0214 & new_n39814_;
  assign new_n39871_ = ~new_n39816_ & ~new_n39870_;
  assign new_n39872_ = ~pi0212 & ~new_n39871_;
  assign new_n39873_ = ~pi0211 & new_n39811_;
  assign new_n39874_ = ~new_n39841_ & ~new_n39873_;
  assign new_n39875_ = pi0214 & ~new_n39874_;
  assign new_n39876_ = ~pi0214 & ~new_n39814_;
  assign new_n39877_ = pi0212 & ~new_n39876_;
  assign new_n39878_ = ~new_n39875_ & new_n39877_;
  assign new_n39879_ = ~new_n39872_ & ~new_n39878_;
  assign new_n39880_ = ~pi0219 & ~new_n39879_;
  assign new_n39881_ = new_n39840_ & ~new_n39880_;
  assign new_n39882_ = new_n39869_ & ~new_n39881_;
  assign new_n39883_ = new_n39405_ & new_n39866_;
  assign new_n39884_ = ~pi1151 & ~new_n39883_;
  assign new_n39885_ = ~pi0219 & new_n38788_;
  assign new_n39886_ = new_n39814_ & new_n39885_;
  assign new_n39887_ = ~new_n39811_ & ~new_n39885_;
  assign new_n39888_ = ~po1038 & ~new_n39887_;
  assign new_n39889_ = ~new_n39886_ & new_n39888_;
  assign new_n39890_ = new_n39884_ & ~new_n39889_;
  assign new_n39891_ = ~pi1152 & ~new_n39890_;
  assign new_n39892_ = ~new_n39882_ & new_n39891_;
  assign new_n39893_ = pi0209 & ~new_n39892_;
  assign new_n39894_ = ~new_n39864_ & new_n39893_;
  assign new_n39895_ = ~pi0214 & new_n39676_;
  assign new_n39896_ = ~new_n13061_ & ~new_n39683_;
  assign new_n39897_ = ~new_n39639_ & new_n39896_;
  assign new_n39898_ = pi0214 & ~new_n39897_;
  assign new_n39899_ = pi0212 & ~new_n39898_;
  assign new_n39900_ = ~new_n39895_ & new_n39899_;
  assign new_n39901_ = ~pi0212 & ~new_n39678_;
  assign new_n39902_ = ~new_n39900_ & ~new_n39901_;
  assign new_n39903_ = ~pi0219 & ~new_n39902_;
  assign new_n39904_ = ~pi0211 & pi0299;
  assign new_n39905_ = ~new_n39683_ & ~new_n39904_;
  assign new_n39906_ = ~new_n39639_ & new_n39905_;
  assign new_n39907_ = ~new_n39677_ & ~new_n39906_;
  assign new_n39908_ = pi0219 & ~new_n39907_;
  assign new_n39909_ = ~po1038 & ~new_n39908_;
  assign new_n39910_ = ~new_n39903_ & new_n39909_;
  assign new_n39911_ = new_n39869_ & ~new_n39910_;
  assign new_n39912_ = new_n39697_ & new_n39700_;
  assign new_n39913_ = pi0212 & ~new_n39697_;
  assign new_n39914_ = ~new_n39896_ & new_n39913_;
  assign new_n39915_ = ~pi0219 & ~new_n39914_;
  assign new_n39916_ = new_n38421_ & new_n39738_;
  assign new_n39917_ = ~new_n39682_ & ~new_n39916_;
  assign new_n39918_ = new_n39915_ & new_n39917_;
  assign new_n39919_ = ~new_n39912_ & new_n39918_;
  assign new_n39920_ = pi0219 & ~new_n39682_;
  assign new_n39921_ = ~po1038 & ~new_n39920_;
  assign new_n39922_ = new_n39700_ & new_n39921_;
  assign new_n39923_ = ~new_n39919_ & new_n39922_;
  assign new_n39924_ = new_n39884_ & ~new_n39923_;
  assign new_n39925_ = ~pi1152 & ~new_n39924_;
  assign new_n39926_ = ~new_n39911_ & new_n39925_;
  assign new_n39927_ = ~new_n39683_ & new_n39757_;
  assign new_n39928_ = ~new_n39748_ & new_n39927_;
  assign new_n39929_ = pi0214 & new_n39928_;
  assign new_n39930_ = ~new_n39762_ & ~new_n39929_;
  assign new_n39931_ = ~pi0212 & ~new_n39930_;
  assign new_n39932_ = ~new_n39928_ & ~new_n39931_;
  assign new_n39933_ = pi0219 & ~new_n39932_;
  assign new_n39934_ = ~po1038 & ~new_n39933_;
  assign new_n39935_ = pi1153 & ~new_n39687_;
  assign new_n39936_ = ~new_n39750_ & ~new_n39935_;
  assign new_n39937_ = new_n39761_ & new_n39936_;
  assign new_n39938_ = pi0214 & new_n39747_;
  assign new_n39939_ = pi0212 & ~new_n39938_;
  assign new_n39940_ = ~new_n39937_ & new_n39939_;
  assign new_n39941_ = pi0214 & new_n39757_;
  assign new_n39942_ = new_n39936_ & new_n39941_;
  assign new_n39943_ = new_n39763_ & ~new_n39942_;
  assign new_n39944_ = ~pi0219 & ~new_n39943_;
  assign new_n39945_ = ~new_n39940_ & new_n39944_;
  assign new_n39946_ = new_n39934_ & ~new_n39945_;
  assign new_n39947_ = new_n39832_ & ~new_n39946_;
  assign new_n39948_ = pi0219 & ~new_n39737_;
  assign new_n39949_ = ~po1038 & ~new_n39948_;
  assign new_n39950_ = ~pi0211 & new_n39718_;
  assign new_n39951_ = new_n39730_ & ~new_n39950_;
  assign new_n39952_ = ~new_n38788_ & new_n39737_;
  assign new_n39953_ = pi0299 & new_n38728_;
  assign new_n39954_ = ~pi0219 & ~new_n39953_;
  assign new_n39955_ = ~new_n39952_ & new_n39954_;
  assign new_n39956_ = ~new_n39951_ & new_n39955_;
  assign new_n39957_ = new_n39949_ & ~new_n39956_;
  assign new_n39958_ = new_n39854_ & ~new_n39957_;
  assign new_n39959_ = pi1152 & ~new_n39958_;
  assign new_n39960_ = ~new_n39947_ & new_n39959_;
  assign new_n39961_ = ~new_n39926_ & ~new_n39960_;
  assign new_n39962_ = ~pi0209 & new_n39961_;
  assign new_n39963_ = ~pi0213 & ~new_n39962_;
  assign new_n39964_ = ~new_n39894_ & new_n39963_;
  assign new_n39965_ = ~new_n39824_ & ~new_n39964_;
  assign new_n39966_ = pi0230 & ~new_n39965_;
  assign new_n39967_ = ~pi0230 & pi0238;
  assign po0395 = new_n39966_ | new_n39967_;
  assign new_n39969_ = new_n38449_ & ~new_n38566_;
  assign new_n39970_ = ~pi0214 & new_n39969_;
  assign new_n39971_ = ~pi0212 & ~new_n39970_;
  assign new_n39972_ = ~pi0219 & new_n39971_;
  assign new_n39973_ = pi0299 & pi1158;
  assign new_n39974_ = ~new_n38449_ & new_n39973_;
  assign new_n39975_ = ~pi0208 & new_n39465_;
  assign new_n39976_ = ~new_n39974_ & ~new_n39975_;
  assign new_n39977_ = ~pi0211 & ~new_n39976_;
  assign new_n39978_ = pi0208 & pi0299;
  assign new_n39979_ = pi1157 & ~new_n39978_;
  assign new_n39980_ = ~new_n38862_ & new_n39979_;
  assign new_n39981_ = ~pi1157 & ~new_n39969_;
  assign new_n39982_ = pi0211 & ~new_n39981_;
  assign new_n39983_ = ~new_n39980_ & new_n39982_;
  assign new_n39984_ = ~new_n39977_ & ~new_n39983_;
  assign new_n39985_ = pi0214 & ~new_n39984_;
  assign new_n39986_ = new_n39972_ & ~new_n39985_;
  assign new_n39987_ = pi0219 & new_n39971_;
  assign new_n39988_ = pi0211 & ~new_n39969_;
  assign new_n39989_ = pi0214 & ~new_n39988_;
  assign new_n39990_ = ~new_n38905_ & new_n39092_;
  assign new_n39991_ = new_n39989_ & ~new_n39990_;
  assign new_n39992_ = new_n39987_ & ~new_n39991_;
  assign new_n39993_ = pi0212 & ~new_n39969_;
  assign new_n39994_ = ~po1038 & ~new_n39993_;
  assign new_n39995_ = ~pi0209 & new_n39994_;
  assign new_n39996_ = ~new_n39992_ & new_n39995_;
  assign new_n39997_ = ~new_n39986_ & new_n39996_;
  assign new_n39998_ = new_n39447_ & ~new_n39539_;
  assign new_n39999_ = ~pi0214 & new_n39998_;
  assign new_n40000_ = ~pi0212 & ~new_n39999_;
  assign new_n40001_ = ~pi0219 & new_n40000_;
  assign new_n40002_ = pi0208 & ~new_n39973_;
  assign new_n40003_ = ~new_n38707_ & ~new_n40002_;
  assign new_n40004_ = ~new_n39480_ & new_n40003_;
  assign new_n40005_ = new_n39489_ & ~new_n40004_;
  assign new_n40006_ = ~new_n39456_ & new_n39979_;
  assign new_n40007_ = ~new_n39539_ & ~new_n40006_;
  assign new_n40008_ = pi0211 & ~new_n40007_;
  assign new_n40009_ = pi0214 & ~new_n40008_;
  assign new_n40010_ = ~new_n40005_ & new_n40009_;
  assign new_n40011_ = new_n40001_ & ~new_n40010_;
  assign new_n40012_ = pi0219 & new_n40000_;
  assign new_n40013_ = pi0211 & ~new_n39998_;
  assign new_n40014_ = new_n39092_ & ~new_n39998_;
  assign new_n40015_ = pi0214 & ~new_n40014_;
  assign new_n40016_ = ~new_n40013_ & new_n40015_;
  assign new_n40017_ = new_n40012_ & ~new_n40016_;
  assign new_n40018_ = pi0212 & ~new_n39998_;
  assign new_n40019_ = ~po1038 & ~new_n40018_;
  assign new_n40020_ = pi0209 & new_n40019_;
  assign new_n40021_ = ~new_n40017_ & new_n40020_;
  assign new_n40022_ = ~new_n40011_ & new_n40021_;
  assign new_n40023_ = ~pi0219 & ~new_n39403_;
  assign new_n40024_ = ~new_n39408_ & ~new_n40023_;
  assign new_n40025_ = pi0213 & ~new_n40024_;
  assign new_n40026_ = ~new_n40022_ & new_n40025_;
  assign new_n40027_ = ~new_n39997_ & new_n40026_;
  assign new_n40028_ = ~pi0211 & ~new_n38512_;
  assign new_n40029_ = ~new_n39589_ & new_n40028_;
  assign new_n40030_ = pi0214 & ~new_n40013_;
  assign new_n40031_ = ~new_n40029_ & new_n40030_;
  assign new_n40032_ = new_n40012_ & ~new_n40031_;
  assign new_n40033_ = pi0211 & ~new_n38510_;
  assign new_n40034_ = ~new_n39589_ & new_n40033_;
  assign new_n40035_ = new_n40015_ & ~new_n40034_;
  assign new_n40036_ = new_n40001_ & ~new_n40035_;
  assign new_n40037_ = new_n40019_ & ~new_n40036_;
  assign new_n40038_ = ~new_n40032_ & new_n40037_;
  assign new_n40039_ = pi0209 & ~new_n40038_;
  assign new_n40040_ = ~new_n38512_ & ~new_n38850_;
  assign new_n40041_ = new_n39989_ & ~new_n40040_;
  assign new_n40042_ = new_n39987_ & ~new_n40041_;
  assign new_n40043_ = ~new_n38911_ & new_n40033_;
  assign new_n40044_ = pi0214 & ~new_n40043_;
  assign new_n40045_ = ~new_n39990_ & new_n40044_;
  assign new_n40046_ = new_n39972_ & ~new_n40045_;
  assign new_n40047_ = new_n39994_ & ~new_n40046_;
  assign new_n40048_ = ~new_n40042_ & new_n40047_;
  assign new_n40049_ = ~pi0209 & ~new_n40048_;
  assign new_n40050_ = ~new_n40039_ & ~new_n40049_;
  assign new_n40051_ = po1038 & ~new_n39150_;
  assign new_n40052_ = new_n38421_ & ~new_n39148_;
  assign new_n40053_ = new_n40051_ & new_n40052_;
  assign new_n40054_ = ~pi0213 & ~new_n40053_;
  assign new_n40055_ = ~new_n40050_ & new_n40054_;
  assign new_n40056_ = ~new_n40027_ & ~new_n40055_;
  assign new_n40057_ = pi0230 & ~new_n40056_;
  assign new_n40058_ = ~pi0230 & ~pi0239;
  assign po0396 = ~new_n40057_ & ~new_n40058_;
  assign new_n40060_ = ~po1038 & new_n39736_;
  assign new_n40061_ = ~new_n39921_ & ~new_n40060_;
  assign new_n40062_ = ~pi0214 & ~new_n39736_;
  assign new_n40063_ = ~pi0212 & ~new_n40062_;
  assign new_n40064_ = new_n11373_ & new_n38449_;
  assign new_n40065_ = ~pi0299 & ~new_n40064_;
  assign new_n40066_ = ~new_n39713_ & new_n40065_;
  assign new_n40067_ = pi0214 & new_n40066_;
  assign new_n40068_ = new_n40063_ & ~new_n40067_;
  assign new_n40069_ = ~pi0219 & ~new_n40068_;
  assign new_n40070_ = ~pi0211 & ~new_n40066_;
  assign new_n40071_ = pi0211 & new_n39736_;
  assign new_n40072_ = pi0214 & ~new_n40071_;
  assign new_n40073_ = ~new_n40070_ & new_n40072_;
  assign new_n40074_ = pi0212 & ~new_n40073_;
  assign new_n40075_ = ~new_n40066_ & new_n40074_;
  assign new_n40076_ = new_n40069_ & ~new_n40075_;
  assign new_n40077_ = ~new_n40061_ & ~new_n40076_;
  assign new_n40078_ = ~new_n39826_ & ~new_n40077_;
  assign new_n40079_ = ~pi1147 & new_n40078_;
  assign new_n40080_ = ~pi0211 & po1038;
  assign new_n40081_ = ~new_n39405_ & ~new_n40080_;
  assign new_n40082_ = ~new_n38413_ & ~new_n40081_;
  assign new_n40083_ = pi0299 & ~new_n38413_;
  assign new_n40084_ = ~po1038 & ~new_n38415_;
  assign new_n40085_ = new_n40083_ & new_n40084_;
  assign new_n40086_ = new_n38539_ & ~new_n38836_;
  assign new_n40087_ = ~po1038 & new_n40086_;
  assign new_n40088_ = ~new_n40085_ & ~new_n40087_;
  assign new_n40089_ = ~new_n40082_ & new_n40088_;
  assign new_n40090_ = pi1147 & new_n40089_;
  assign new_n40091_ = pi1149 & ~new_n40090_;
  assign new_n40092_ = ~new_n40079_ & new_n40091_;
  assign new_n40093_ = pi0211 & new_n38421_;
  assign new_n40094_ = pi0212 & new_n38717_;
  assign new_n40095_ = ~new_n40093_ & ~new_n40094_;
  assign new_n40096_ = new_n39405_ & ~new_n40095_;
  assign new_n40097_ = ~new_n38837_ & ~new_n39028_;
  assign new_n40098_ = ~new_n10624_ & new_n38638_;
  assign new_n40099_ = ~new_n40097_ & ~new_n40098_;
  assign new_n40100_ = new_n39715_ & new_n40099_;
  assign new_n40101_ = pi0299 & new_n10484_;
  assign new_n40102_ = ~new_n40100_ & ~new_n40101_;
  assign new_n40103_ = ~pi0212 & ~new_n40102_;
  assign new_n40104_ = ~pi0219 & ~new_n40103_;
  assign new_n40105_ = ~pi0299 & ~new_n40099_;
  assign new_n40106_ = pi0214 & ~new_n40105_;
  assign new_n40107_ = ~pi0214 & new_n40100_;
  assign new_n40108_ = ~pi0212 & ~new_n40107_;
  assign new_n40109_ = ~new_n40106_ & new_n40108_;
  assign new_n40110_ = ~pi0211 & ~new_n40105_;
  assign new_n40111_ = ~new_n40100_ & ~new_n40110_;
  assign new_n40112_ = pi0214 & ~new_n40111_;
  assign new_n40113_ = pi0212 & ~new_n40112_;
  assign new_n40114_ = ~pi0214 & ~new_n40105_;
  assign new_n40115_ = new_n40113_ & ~new_n40114_;
  assign new_n40116_ = ~new_n40109_ & ~new_n40115_;
  assign new_n40117_ = ~new_n13061_ & ~new_n40100_;
  assign new_n40118_ = ~new_n40106_ & new_n40117_;
  assign new_n40119_ = pi0212 & ~new_n40118_;
  assign new_n40120_ = new_n40116_ & new_n40119_;
  assign new_n40121_ = new_n40104_ & ~new_n40120_;
  assign new_n40122_ = pi0219 & ~new_n40100_;
  assign new_n40123_ = ~po1038 & ~new_n40122_;
  assign new_n40124_ = ~new_n40121_ & new_n40123_;
  assign new_n40125_ = ~new_n40096_ & ~new_n40124_;
  assign new_n40126_ = ~pi1147 & new_n40125_;
  assign new_n40127_ = pi0212 & ~new_n38668_;
  assign new_n40128_ = ~pi0219 & ~new_n40093_;
  assign new_n40129_ = ~new_n40127_ & new_n40128_;
  assign new_n40130_ = new_n40085_ & ~new_n40129_;
  assign new_n40131_ = ~po1038 & ~new_n39757_;
  assign new_n40132_ = new_n38416_ & ~new_n40129_;
  assign new_n40133_ = ~new_n40131_ & ~new_n40132_;
  assign new_n40134_ = ~new_n40130_ & new_n40133_;
  assign new_n40135_ = pi1147 & new_n40134_;
  assign new_n40136_ = ~pi1149 & ~new_n40135_;
  assign new_n40137_ = ~new_n40126_ & new_n40136_;
  assign new_n40138_ = ~new_n40092_ & ~new_n40137_;
  assign new_n40139_ = pi1148 & ~new_n40138_;
  assign new_n40140_ = new_n10486_ & ~new_n39865_;
  assign new_n40141_ = new_n38416_ & ~new_n40140_;
  assign new_n40142_ = ~pi0211 & ~new_n39638_;
  assign new_n40143_ = pi0211 & ~new_n39662_;
  assign new_n40144_ = pi0214 & ~new_n40143_;
  assign new_n40145_ = ~new_n40142_ & new_n40144_;
  assign new_n40146_ = new_n10729_ & ~new_n40145_;
  assign new_n40147_ = ~pi0214 & new_n39638_;
  assign new_n40148_ = ~pi0212 & ~new_n40147_;
  assign new_n40149_ = pi0214 & new_n39675_;
  assign new_n40150_ = new_n40148_ & ~new_n40149_;
  assign new_n40151_ = ~pi0219 & ~new_n40150_;
  assign new_n40152_ = pi0212 & ~new_n40145_;
  assign new_n40153_ = ~new_n39675_ & new_n40152_;
  assign new_n40154_ = new_n40151_ & ~new_n40153_;
  assign new_n40155_ = ~new_n40146_ & new_n40154_;
  assign new_n40156_ = pi0212 & ~new_n39675_;
  assign new_n40157_ = pi0219 & ~new_n40156_;
  assign new_n40158_ = ~new_n40150_ & new_n40157_;
  assign new_n40159_ = ~po1038 & ~new_n40158_;
  assign new_n40160_ = ~new_n40155_ & new_n40159_;
  assign new_n40161_ = ~new_n40141_ & ~new_n40160_;
  assign new_n40162_ = pi1147 & new_n40161_;
  assign new_n40163_ = new_n16479_ & new_n39686_;
  assign new_n40164_ = ~pi0219 & ~new_n16479_;
  assign new_n40165_ = new_n39865_ & new_n40164_;
  assign new_n40166_ = ~new_n40163_ & ~new_n40165_;
  assign new_n40167_ = ~pi1147 & new_n40166_;
  assign new_n40168_ = pi1149 & ~new_n40167_;
  assign new_n40169_ = ~new_n40162_ & new_n40168_;
  assign new_n40170_ = ~pi0212 & ~new_n40101_;
  assign new_n40171_ = new_n39757_ & new_n40170_;
  assign new_n40172_ = new_n39757_ & ~new_n39904_;
  assign new_n40173_ = ~new_n39761_ & ~new_n40172_;
  assign new_n40174_ = ~pi0214 & new_n13061_;
  assign new_n40175_ = pi0212 & ~new_n40174_;
  assign new_n40176_ = ~new_n40173_ & new_n40175_;
  assign new_n40177_ = ~new_n40171_ & ~new_n40176_;
  assign new_n40178_ = ~pi0219 & ~new_n40177_;
  assign new_n40179_ = new_n38608_ & ~new_n39710_;
  assign new_n40180_ = pi0208 & ~new_n40179_;
  assign new_n40181_ = ~pi0199 & ~new_n40180_;
  assign new_n40182_ = ~new_n39757_ & ~new_n40181_;
  assign new_n40183_ = ~pi0299 & ~new_n40182_;
  assign new_n40184_ = ~pi0219 & new_n40183_;
  assign new_n40185_ = ~new_n40178_ & ~new_n40184_;
  assign new_n40186_ = ~pi0211 & ~new_n40185_;
  assign new_n40187_ = ~new_n13061_ & new_n39941_;
  assign new_n40188_ = ~pi0214 & new_n40172_;
  assign new_n40189_ = pi0212 & ~new_n40188_;
  assign new_n40190_ = ~new_n40187_ & new_n40189_;
  assign new_n40191_ = ~pi0212 & new_n40173_;
  assign new_n40192_ = ~pi0219 & ~new_n40191_;
  assign new_n40193_ = ~new_n40190_ & new_n40192_;
  assign new_n40194_ = pi0219 & ~new_n39904_;
  assign new_n40195_ = new_n40084_ & ~new_n40194_;
  assign new_n40196_ = ~new_n40131_ & ~new_n40195_;
  assign new_n40197_ = ~new_n40193_ & ~new_n40196_;
  assign new_n40198_ = ~new_n40183_ & new_n40197_;
  assign new_n40199_ = ~new_n40186_ & new_n40198_;
  assign new_n40200_ = ~new_n39830_ & ~new_n40199_;
  assign new_n40201_ = pi1147 & ~pi1149;
  assign new_n40202_ = ~new_n40200_ & new_n40201_;
  assign new_n40203_ = ~new_n40169_ & ~new_n40202_;
  assign new_n40204_ = ~pi1148 & ~new_n40203_;
  assign new_n40205_ = ~new_n40139_ & ~new_n40204_;
  assign new_n40206_ = pi0213 & ~new_n40205_;
  assign new_n40207_ = ~po1038 & new_n40100_;
  assign new_n40208_ = ~pi0211 & pi1146;
  assign new_n40209_ = pi0211 & pi1145;
  assign new_n40210_ = ~new_n40208_ & ~new_n40209_;
  assign new_n40211_ = pi0214 & ~new_n40210_;
  assign new_n40212_ = pi0211 & pi1146;
  assign new_n40213_ = ~pi0214 & new_n40212_;
  assign new_n40214_ = ~new_n40211_ & ~new_n40213_;
  assign new_n40215_ = pi0212 & ~new_n40214_;
  assign new_n40216_ = new_n38421_ & new_n40212_;
  assign new_n40217_ = ~new_n40215_ & ~new_n40216_;
  assign new_n40218_ = ~new_n38970_ & new_n40217_;
  assign new_n40219_ = po1038 & new_n39369_;
  assign new_n40220_ = ~new_n39405_ & ~new_n40219_;
  assign new_n40221_ = ~new_n40218_ & ~new_n40220_;
  assign new_n40222_ = ~pi1147 & ~new_n40221_;
  assign new_n40223_ = ~pi0211 & new_n39561_;
  assign new_n40224_ = pi0219 & ~new_n40223_;
  assign new_n40225_ = new_n40084_ & ~new_n40224_;
  assign new_n40226_ = pi0219 & new_n40225_;
  assign new_n40227_ = pi0299 & ~new_n40217_;
  assign new_n40228_ = new_n36114_ & new_n40227_;
  assign new_n40229_ = ~new_n40226_ & ~new_n40228_;
  assign new_n40230_ = new_n40222_ & new_n40229_;
  assign new_n40231_ = ~new_n40207_ & new_n40230_;
  assign new_n40232_ = new_n10732_ & new_n38794_;
  assign new_n40233_ = po1038 & new_n40232_;
  assign new_n40234_ = pi1147 & ~new_n40233_;
  assign new_n40235_ = ~new_n40221_ & new_n40234_;
  assign new_n40236_ = ~new_n40131_ & ~new_n40225_;
  assign new_n40237_ = pi0299 & pi1146;
  assign new_n40238_ = pi0211 & new_n40237_;
  assign new_n40239_ = ~new_n39904_ & ~new_n40238_;
  assign new_n40240_ = new_n39757_ & new_n40239_;
  assign new_n40241_ = new_n38788_ & ~new_n40240_;
  assign new_n40242_ = new_n38413_ & ~new_n39757_;
  assign new_n40243_ = ~pi0219 & ~new_n40242_;
  assign new_n40244_ = pi0299 & ~new_n40210_;
  assign new_n40245_ = new_n39757_ & ~new_n40244_;
  assign new_n40246_ = new_n10729_ & ~new_n40245_;
  assign new_n40247_ = new_n40243_ & ~new_n40246_;
  assign new_n40248_ = ~new_n40241_ & new_n40247_;
  assign new_n40249_ = ~new_n40236_ & ~new_n40248_;
  assign new_n40250_ = new_n40235_ & ~new_n40249_;
  assign new_n40251_ = pi1148 & ~new_n40250_;
  assign new_n40252_ = ~new_n40231_ & new_n40251_;
  assign new_n40253_ = ~pi1146 & new_n13061_;
  assign new_n40254_ = new_n38788_ & ~new_n40253_;
  assign new_n40255_ = ~new_n40246_ & ~new_n40254_;
  assign new_n40256_ = ~pi0219 & ~new_n40183_;
  assign new_n40257_ = ~new_n40255_ & new_n40256_;
  assign new_n40258_ = new_n39369_ & new_n39393_;
  assign new_n40259_ = ~new_n38794_ & new_n40182_;
  assign new_n40260_ = ~new_n40258_ & ~new_n40259_;
  assign new_n40261_ = ~new_n40257_ & new_n40260_;
  assign new_n40262_ = ~po1038 & ~new_n40261_;
  assign new_n40263_ = new_n40235_ & ~new_n40262_;
  assign new_n40264_ = ~pi1148 & ~new_n40230_;
  assign new_n40265_ = ~new_n40263_ & new_n40264_;
  assign new_n40266_ = ~new_n40252_ & ~new_n40265_;
  assign new_n40267_ = ~pi1149 & ~new_n40266_;
  assign new_n40268_ = pi0219 & new_n39638_;
  assign new_n40269_ = ~po1038 & ~new_n40268_;
  assign new_n40270_ = ~new_n40225_ & ~new_n40269_;
  assign new_n40271_ = ~pi0299 & new_n39661_;
  assign new_n40272_ = ~new_n39431_ & ~new_n40271_;
  assign new_n40273_ = ~new_n40237_ & new_n40272_;
  assign new_n40274_ = pi0211 & ~new_n40273_;
  assign new_n40275_ = ~new_n39673_ & ~new_n40274_;
  assign new_n40276_ = ~pi0214 & new_n40275_;
  assign new_n40277_ = pi0214 & ~new_n40244_;
  assign new_n40278_ = new_n40272_ & new_n40277_;
  assign new_n40279_ = pi0212 & ~new_n40278_;
  assign new_n40280_ = ~new_n40276_ & new_n40279_;
  assign new_n40281_ = pi0214 & new_n40275_;
  assign new_n40282_ = new_n40148_ & ~new_n40281_;
  assign new_n40283_ = ~pi0219 & ~new_n40282_;
  assign new_n40284_ = ~new_n40280_ & new_n40283_;
  assign new_n40285_ = ~new_n40270_ & ~new_n40284_;
  assign new_n40286_ = new_n40235_ & ~new_n40285_;
  assign new_n40287_ = ~new_n40163_ & new_n40230_;
  assign new_n40288_ = ~pi1148 & ~new_n40287_;
  assign new_n40289_ = ~new_n40286_ & new_n40288_;
  assign new_n40290_ = ~new_n38413_ & new_n40070_;
  assign new_n40291_ = ~new_n38414_ & new_n39736_;
  assign new_n40292_ = pi0219 & ~new_n40291_;
  assign new_n40293_ = ~new_n40290_ & new_n40292_;
  assign new_n40294_ = ~po1038 & ~new_n40293_;
  assign new_n40295_ = new_n11373_ & new_n40294_;
  assign new_n40296_ = ~new_n40225_ & ~new_n40295_;
  assign new_n40297_ = pi0212 & ~new_n40066_;
  assign new_n40298_ = ~new_n39736_ & new_n40214_;
  assign new_n40299_ = new_n40297_ & ~new_n40298_;
  assign new_n40300_ = ~new_n39736_ & ~new_n40238_;
  assign new_n40301_ = new_n40063_ & ~new_n40300_;
  assign new_n40302_ = ~pi0219 & ~new_n40301_;
  assign new_n40303_ = ~new_n40299_ & new_n40302_;
  assign new_n40304_ = ~new_n40296_ & ~new_n40303_;
  assign new_n40305_ = new_n40222_ & ~new_n40304_;
  assign new_n40306_ = pi0219 & ~new_n40086_;
  assign new_n40307_ = ~po1038 & ~new_n40306_;
  assign new_n40308_ = ~pi0299 & ~new_n40086_;
  assign new_n40309_ = pi0212 & ~new_n40308_;
  assign new_n40310_ = pi0299 & new_n40127_;
  assign new_n40311_ = new_n40309_ & ~new_n40310_;
  assign new_n40312_ = pi0211 & ~new_n40086_;
  assign new_n40313_ = pi0214 & pi0299;
  assign new_n40314_ = ~new_n40086_ & ~new_n40313_;
  assign new_n40315_ = ~pi0212 & ~new_n40314_;
  assign new_n40316_ = ~new_n40312_ & new_n40315_;
  assign new_n40317_ = ~pi0219 & ~new_n40316_;
  assign new_n40318_ = ~new_n40311_ & new_n40317_;
  assign new_n40319_ = new_n40307_ & ~new_n40318_;
  assign new_n40320_ = new_n40229_ & new_n40235_;
  assign new_n40321_ = ~new_n40319_ & new_n40320_;
  assign new_n40322_ = pi1148 & ~new_n40321_;
  assign new_n40323_ = ~new_n40305_ & new_n40322_;
  assign new_n40324_ = ~new_n40289_ & ~new_n40323_;
  assign new_n40325_ = pi1149 & ~new_n40324_;
  assign new_n40326_ = ~new_n40267_ & ~new_n40325_;
  assign new_n40327_ = ~pi0213 & ~new_n40326_;
  assign new_n40328_ = pi0209 & ~new_n40327_;
  assign new_n40329_ = ~new_n40206_ & new_n40328_;
  assign new_n40330_ = pi0199 & pi1145;
  assign new_n40331_ = ~pi0200 & ~new_n40330_;
  assign new_n40332_ = ~pi0199 & pi1146;
  assign new_n40333_ = new_n40331_ & ~new_n40332_;
  assign new_n40334_ = pi0200 & ~new_n39386_;
  assign new_n40335_ = new_n38442_ & ~new_n40334_;
  assign new_n40336_ = ~new_n40333_ & new_n40335_;
  assign new_n40337_ = ~new_n38837_ & ~new_n40336_;
  assign new_n40338_ = pi0200 & ~new_n40332_;
  assign new_n40339_ = ~pi0299 & ~new_n40338_;
  assign new_n40340_ = ~new_n40331_ & new_n40339_;
  assign new_n40341_ = ~new_n10624_ & ~new_n40340_;
  assign new_n40342_ = ~new_n40337_ & ~new_n40341_;
  assign new_n40343_ = ~pi1147 & ~po1038;
  assign new_n40344_ = new_n40342_ & new_n40343_;
  assign new_n40345_ = new_n38607_ & ~new_n40330_;
  assign new_n40346_ = new_n40339_ & ~new_n40345_;
  assign new_n40347_ = ~new_n10624_ & ~new_n40346_;
  assign new_n40348_ = ~new_n40337_ & ~new_n40347_;
  assign new_n40349_ = ~new_n38414_ & new_n40348_;
  assign new_n40350_ = pi0219 & ~new_n40349_;
  assign new_n40351_ = ~pi0207 & new_n40346_;
  assign new_n40352_ = ~new_n40237_ & ~new_n40336_;
  assign new_n40353_ = ~new_n40351_ & new_n40352_;
  assign new_n40354_ = pi0208 & ~new_n40353_;
  assign new_n40355_ = new_n38449_ & new_n40346_;
  assign new_n40356_ = ~new_n40354_ & ~new_n40355_;
  assign new_n40357_ = ~pi0299 & new_n40356_;
  assign new_n40358_ = ~pi0211 & ~new_n40357_;
  assign new_n40359_ = ~new_n38413_ & new_n40358_;
  assign new_n40360_ = new_n40350_ & ~new_n40359_;
  assign new_n40361_ = ~po1038 & ~new_n40360_;
  assign new_n40362_ = pi0211 & ~new_n40357_;
  assign new_n40363_ = new_n40331_ & new_n40351_;
  assign new_n40364_ = new_n40354_ & ~new_n40363_;
  assign new_n40365_ = new_n38449_ & new_n40340_;
  assign new_n40366_ = ~new_n40364_ & ~new_n40365_;
  assign new_n40367_ = ~pi0299 & new_n40366_;
  assign new_n40368_ = pi0214 & ~new_n40367_;
  assign new_n40369_ = ~new_n40362_ & ~new_n40368_;
  assign new_n40370_ = pi0212 & ~new_n40369_;
  assign new_n40371_ = new_n10484_ & ~new_n40357_;
  assign new_n40372_ = ~pi0219 & ~new_n40348_;
  assign new_n40373_ = ~new_n40371_ & new_n40372_;
  assign new_n40374_ = ~new_n40370_ & new_n40373_;
  assign new_n40375_ = new_n40361_ & ~new_n40374_;
  assign new_n40376_ = ~pi0214 & ~new_n40348_;
  assign new_n40377_ = ~new_n40358_ & new_n40376_;
  assign new_n40378_ = pi0214 & ~new_n40348_;
  assign new_n40379_ = ~new_n40362_ & new_n40378_;
  assign new_n40380_ = pi0212 & ~new_n40379_;
  assign new_n40381_ = ~new_n40377_ & new_n40380_;
  assign new_n40382_ = ~new_n40348_ & ~new_n40358_;
  assign new_n40383_ = ~pi0212 & ~new_n40376_;
  assign new_n40384_ = ~new_n40382_ & new_n40383_;
  assign new_n40385_ = ~pi0219 & ~new_n40384_;
  assign new_n40386_ = ~new_n40381_ & new_n40385_;
  assign new_n40387_ = new_n40375_ & ~new_n40386_;
  assign new_n40388_ = ~new_n39830_ & ~new_n40387_;
  assign new_n40389_ = pi1147 & ~new_n40388_;
  assign new_n40390_ = ~new_n40344_ & ~new_n40389_;
  assign new_n40391_ = ~pi1149 & ~new_n40390_;
  assign new_n40392_ = new_n40361_ & ~new_n40386_;
  assign new_n40393_ = ~new_n40141_ & ~new_n40392_;
  assign new_n40394_ = pi1147 & ~new_n40393_;
  assign new_n40395_ = ~pi1147 & new_n40232_;
  assign new_n40396_ = ~new_n40344_ & ~new_n40395_;
  assign new_n40397_ = new_n16479_ & new_n40232_;
  assign new_n40398_ = new_n40366_ & new_n40397_;
  assign new_n40399_ = ~new_n40396_ & ~new_n40398_;
  assign new_n40400_ = ~new_n40394_ & ~new_n40399_;
  assign new_n40401_ = pi1149 & ~new_n40400_;
  assign new_n40402_ = ~pi1148 & ~new_n40401_;
  assign new_n40403_ = ~new_n40391_ & new_n40402_;
  assign new_n40404_ = new_n38413_ & new_n40342_;
  assign new_n40405_ = new_n40374_ & ~new_n40404_;
  assign new_n40406_ = pi0214 & new_n40382_;
  assign new_n40407_ = ~new_n40367_ & ~new_n40406_;
  assign new_n40408_ = pi0212 & ~new_n40407_;
  assign new_n40409_ = ~pi0214 & new_n40342_;
  assign new_n40410_ = ~pi0212 & ~new_n40409_;
  assign new_n40411_ = ~new_n40368_ & new_n40410_;
  assign new_n40412_ = ~new_n40408_ & ~new_n40411_;
  assign new_n40413_ = ~pi0219 & ~new_n40412_;
  assign new_n40414_ = pi0219 & ~new_n40342_;
  assign new_n40415_ = ~po1038 & ~new_n40414_;
  assign new_n40416_ = ~new_n40413_ & new_n40415_;
  assign new_n40417_ = ~new_n40405_ & new_n40416_;
  assign new_n40418_ = ~pi1147 & ~new_n40096_;
  assign new_n40419_ = ~new_n40417_ & new_n40418_;
  assign new_n40420_ = pi1147 & ~new_n40132_;
  assign new_n40421_ = ~new_n40375_ & new_n40420_;
  assign new_n40422_ = ~pi1149 & ~new_n40421_;
  assign new_n40423_ = ~new_n40419_ & new_n40422_;
  assign new_n40424_ = ~pi1147 & ~new_n39826_;
  assign new_n40425_ = ~new_n40416_ & new_n40424_;
  assign new_n40426_ = ~new_n40083_ & new_n40372_;
  assign new_n40427_ = new_n40361_ & ~new_n40426_;
  assign new_n40428_ = pi1147 & ~new_n40082_;
  assign new_n40429_ = ~new_n40427_ & new_n40428_;
  assign new_n40430_ = pi1149 & ~new_n40429_;
  assign new_n40431_ = ~new_n40425_ & new_n40430_;
  assign new_n40432_ = pi1148 & ~new_n40431_;
  assign new_n40433_ = ~new_n40423_ & new_n40432_;
  assign new_n40434_ = pi0213 & ~new_n40433_;
  assign new_n40435_ = ~new_n40403_ & new_n40434_;
  assign new_n40436_ = ~new_n40238_ & ~new_n40342_;
  assign new_n40437_ = ~pi0214 & ~new_n40342_;
  assign new_n40438_ = ~pi0212 & ~new_n40437_;
  assign new_n40439_ = ~new_n40436_ & new_n40438_;
  assign new_n40440_ = ~pi0219 & ~new_n40439_;
  assign new_n40441_ = ~pi0299 & ~new_n40366_;
  assign new_n40442_ = new_n40277_ & ~new_n40441_;
  assign new_n40443_ = ~pi0214 & new_n40436_;
  assign new_n40444_ = pi0212 & ~new_n40443_;
  assign new_n40445_ = ~new_n40442_ & new_n40444_;
  assign new_n40446_ = new_n40440_ & ~new_n40445_;
  assign new_n40447_ = pi0219 & ~new_n40404_;
  assign new_n40448_ = ~new_n38413_ & new_n40342_;
  assign new_n40449_ = ~new_n38414_ & ~new_n40448_;
  assign new_n40450_ = ~pi0211 & ~new_n39561_;
  assign new_n40451_ = ~new_n40441_ & new_n40450_;
  assign new_n40452_ = ~new_n40449_ & ~new_n40451_;
  assign new_n40453_ = new_n40447_ & ~new_n40452_;
  assign new_n40454_ = ~po1038 & ~new_n40453_;
  assign new_n40455_ = ~new_n40446_ & new_n40454_;
  assign new_n40456_ = new_n40222_ & ~new_n40455_;
  assign new_n40457_ = ~new_n39558_ & new_n40362_;
  assign new_n40458_ = new_n40277_ & new_n40356_;
  assign new_n40459_ = ~new_n40371_ & ~new_n40458_;
  assign new_n40460_ = ~new_n40457_ & ~new_n40459_;
  assign new_n40461_ = ~pi0214 & new_n40239_;
  assign new_n40462_ = new_n40356_ & new_n40461_;
  assign new_n40463_ = pi0212 & ~new_n40462_;
  assign new_n40464_ = ~new_n40460_ & new_n40463_;
  assign new_n40465_ = ~new_n40384_ & new_n40440_;
  assign new_n40466_ = ~new_n40464_ & new_n40465_;
  assign new_n40467_ = ~new_n39558_ & new_n40358_;
  assign new_n40468_ = ~new_n38413_ & new_n40467_;
  assign new_n40469_ = new_n40350_ & ~new_n40468_;
  assign new_n40470_ = ~po1038 & ~new_n40469_;
  assign new_n40471_ = ~new_n40466_ & new_n40470_;
  assign new_n40472_ = new_n40235_ & ~new_n40471_;
  assign new_n40473_ = ~new_n40456_ & ~new_n40472_;
  assign new_n40474_ = ~pi0213 & new_n40473_;
  assign new_n40475_ = ~pi0209 & ~new_n40474_;
  assign new_n40476_ = ~new_n40435_ & new_n40475_;
  assign new_n40477_ = ~new_n40329_ & ~new_n40476_;
  assign new_n40478_ = pi0230 & ~new_n40477_;
  assign new_n40479_ = ~pi0230 & ~pi0240;
  assign po0397 = ~new_n40478_ & ~new_n40479_;
  assign new_n40481_ = po1038 & ~new_n40232_;
  assign new_n40482_ = pi1151 & ~new_n40481_;
  assign new_n40483_ = ~new_n39747_ & new_n40232_;
  assign new_n40484_ = new_n39927_ & ~new_n40483_;
  assign new_n40485_ = pi1152 & ~new_n40484_;
  assign new_n40486_ = ~po1038 & ~new_n40485_;
  assign new_n40487_ = new_n40482_ & ~new_n40486_;
  assign new_n40488_ = new_n39683_ & new_n39695_;
  assign new_n40489_ = new_n38508_ & new_n39865_;
  assign new_n40490_ = ~new_n39639_ & ~new_n40489_;
  assign new_n40491_ = new_n40482_ & ~new_n40490_;
  assign new_n40492_ = ~new_n40488_ & ~new_n40491_;
  assign new_n40493_ = ~pi1152 & ~new_n40492_;
  assign new_n40494_ = pi1152 & new_n39695_;
  assign new_n40495_ = new_n39737_ & new_n40494_;
  assign new_n40496_ = ~new_n40493_ & ~new_n40495_;
  assign new_n40497_ = ~new_n40487_ & new_n40496_;
  assign new_n40498_ = ~pi1150 & ~new_n40497_;
  assign new_n40499_ = pi1151 & ~new_n39826_;
  assign new_n40500_ = pi0219 & ~new_n39683_;
  assign new_n40501_ = ~po1038 & ~new_n40500_;
  assign new_n40502_ = ~new_n40131_ & ~new_n40501_;
  assign new_n40503_ = new_n39763_ & ~new_n39938_;
  assign new_n40504_ = ~pi0219 & ~new_n40503_;
  assign new_n40505_ = ~pi0214 & new_n39747_;
  assign new_n40506_ = pi0212 & ~new_n40505_;
  assign new_n40507_ = ~new_n39929_ & new_n40506_;
  assign new_n40508_ = new_n40504_ & ~new_n40507_;
  assign new_n40509_ = pi1152 & ~new_n40508_;
  assign new_n40510_ = ~pi0299 & ~new_n39663_;
  assign new_n40511_ = ~pi0214 & new_n39662_;
  assign new_n40512_ = pi0212 & ~new_n40511_;
  assign new_n40513_ = ~new_n40149_ & new_n40512_;
  assign new_n40514_ = ~new_n39641_ & ~new_n40513_;
  assign new_n40515_ = ~new_n40510_ & ~new_n40514_;
  assign new_n40516_ = ~pi0219 & ~new_n40515_;
  assign new_n40517_ = ~pi1152 & ~new_n40268_;
  assign new_n40518_ = ~new_n40516_ & new_n40517_;
  assign new_n40519_ = ~new_n40509_ & ~new_n40518_;
  assign new_n40520_ = ~new_n40502_ & ~new_n40519_;
  assign new_n40521_ = new_n40499_ & ~new_n40520_;
  assign new_n40522_ = ~pi1151 & ~new_n40096_;
  assign new_n40523_ = ~pi0212 & ~new_n39687_;
  assign new_n40524_ = ~new_n39697_ & new_n40523_;
  assign new_n40525_ = ~new_n39904_ & new_n40524_;
  assign new_n40526_ = ~pi0219 & ~new_n40525_;
  assign new_n40527_ = pi0214 & ~new_n39696_;
  assign new_n40528_ = ~pi0211 & new_n39697_;
  assign new_n40529_ = pi0212 & ~new_n39687_;
  assign new_n40530_ = ~new_n40528_ & new_n40529_;
  assign new_n40531_ = ~new_n40527_ & new_n40530_;
  assign new_n40532_ = new_n40526_ & ~new_n40531_;
  assign new_n40533_ = ~new_n39683_ & new_n39915_;
  assign new_n40534_ = ~pi0299 & new_n40533_;
  assign new_n40535_ = ~new_n40532_ & ~new_n40534_;
  assign new_n40536_ = new_n40501_ & new_n40535_;
  assign new_n40537_ = ~pi1152 & ~new_n40536_;
  assign new_n40538_ = ~new_n39737_ & ~new_n40535_;
  assign new_n40539_ = new_n39949_ & ~new_n40538_;
  assign new_n40540_ = pi1152 & ~new_n40539_;
  assign new_n40541_ = ~new_n40537_ & ~new_n40540_;
  assign new_n40542_ = new_n40522_ & ~new_n40541_;
  assign new_n40543_ = pi1150 & ~new_n40542_;
  assign new_n40544_ = ~new_n40521_ & new_n40543_;
  assign new_n40545_ = ~new_n40498_ & ~new_n40544_;
  assign new_n40546_ = ~pi1149 & ~new_n40545_;
  assign new_n40547_ = ~new_n38717_ & ~new_n39747_;
  assign new_n40548_ = pi0212 & new_n39927_;
  assign new_n40549_ = ~new_n40547_ & new_n40548_;
  assign new_n40550_ = ~new_n39931_ & ~new_n40549_;
  assign new_n40551_ = ~pi0219 & ~new_n40550_;
  assign new_n40552_ = pi1152 & ~new_n40551_;
  assign new_n40553_ = new_n39934_ & new_n40552_;
  assign new_n40554_ = pi1151 & ~new_n40141_;
  assign new_n40555_ = ~pi0214 & ~new_n39906_;
  assign new_n40556_ = new_n39899_ & ~new_n40555_;
  assign new_n40557_ = ~pi0212 & ~new_n39907_;
  assign new_n40558_ = ~new_n40556_ & ~new_n40557_;
  assign new_n40559_ = ~pi0219 & ~new_n40558_;
  assign new_n40560_ = ~pi1152 & new_n39909_;
  assign new_n40561_ = ~new_n40559_ & new_n40560_;
  assign new_n40562_ = new_n40554_ & ~new_n40561_;
  assign new_n40563_ = ~new_n40553_ & new_n40562_;
  assign new_n40564_ = ~new_n39737_ & new_n39915_;
  assign new_n40565_ = ~new_n40195_ & ~new_n40501_;
  assign new_n40566_ = ~new_n39949_ & new_n40565_;
  assign new_n40567_ = pi1152 & ~new_n40566_;
  assign new_n40568_ = ~new_n40564_ & new_n40567_;
  assign new_n40569_ = ~pi1151 & ~new_n39830_;
  assign new_n40570_ = ~new_n40533_ & ~new_n40565_;
  assign new_n40571_ = ~pi1152 & new_n40570_;
  assign new_n40572_ = new_n40569_ & ~new_n40571_;
  assign new_n40573_ = ~new_n40568_ & new_n40572_;
  assign new_n40574_ = ~pi1150 & ~new_n40573_;
  assign new_n40575_ = ~new_n40563_ & new_n40574_;
  assign new_n40576_ = pi0212 & ~new_n39747_;
  assign new_n40577_ = new_n40504_ & ~new_n40576_;
  assign new_n40578_ = pi1152 & ~new_n40577_;
  assign new_n40579_ = new_n39934_ & new_n40578_;
  assign new_n40580_ = pi1151 & ~new_n40082_;
  assign new_n40581_ = ~new_n39677_ & ~new_n40510_;
  assign new_n40582_ = ~pi0219 & ~new_n40581_;
  assign new_n40583_ = new_n40560_ & ~new_n40582_;
  assign new_n40584_ = new_n40580_ & ~new_n40583_;
  assign new_n40585_ = ~new_n40579_ & new_n40584_;
  assign new_n40586_ = ~pi1151 & ~new_n40132_;
  assign new_n40587_ = new_n10729_ & new_n39724_;
  assign new_n40588_ = ~new_n39698_ & ~new_n39896_;
  assign new_n40589_ = ~new_n10729_ & ~new_n39737_;
  assign new_n40590_ = ~new_n40588_ & new_n40589_;
  assign new_n40591_ = ~new_n40587_ & ~new_n40590_;
  assign new_n40592_ = ~pi0219 & ~new_n40591_;
  assign new_n40593_ = ~new_n40566_ & ~new_n40592_;
  assign new_n40594_ = pi1152 & ~new_n40593_;
  assign new_n40595_ = new_n40537_ & ~new_n40570_;
  assign new_n40596_ = ~new_n40594_ & ~new_n40595_;
  assign new_n40597_ = new_n40586_ & ~new_n40596_;
  assign new_n40598_ = pi1150 & ~new_n40597_;
  assign new_n40599_ = ~new_n40585_ & new_n40598_;
  assign new_n40600_ = ~new_n40575_ & ~new_n40599_;
  assign new_n40601_ = pi1149 & ~new_n40600_;
  assign new_n40602_ = ~new_n40546_ & ~new_n40601_;
  assign new_n40603_ = ~pi0213 & ~new_n40602_;
  assign new_n40604_ = pi0213 & ~new_n39961_;
  assign new_n40605_ = pi0209 & ~new_n40604_;
  assign new_n40606_ = ~new_n40603_ & new_n40605_;
  assign new_n40607_ = ~new_n40148_ & ~new_n40152_;
  assign new_n40608_ = ~new_n38646_ & new_n39673_;
  assign new_n40609_ = ~new_n39674_ & ~new_n40608_;
  assign new_n40610_ = ~new_n40146_ & new_n40609_;
  assign new_n40611_ = ~new_n40607_ & ~new_n40610_;
  assign new_n40612_ = ~pi0219 & ~new_n40611_;
  assign new_n40613_ = new_n40159_ & ~new_n40612_;
  assign new_n40614_ = new_n39869_ & ~new_n40613_;
  assign new_n40615_ = pi0299 & new_n39631_;
  assign new_n40616_ = ~new_n40182_ & ~new_n40489_;
  assign new_n40617_ = ~po1038 & ~new_n40616_;
  assign new_n40618_ = ~new_n40615_ & new_n40617_;
  assign new_n40619_ = new_n39884_ & ~new_n40618_;
  assign new_n40620_ = ~pi1152 & ~new_n40619_;
  assign new_n40621_ = ~new_n40614_ & new_n40620_;
  assign new_n40622_ = ~new_n40145_ & ~new_n40147_;
  assign new_n40623_ = ~pi0219 & ~new_n40310_;
  assign new_n40624_ = ~new_n39678_ & new_n40623_;
  assign new_n40625_ = ~new_n40622_ & new_n40624_;
  assign new_n40626_ = new_n40159_ & ~new_n40625_;
  assign new_n40627_ = new_n39832_ & ~new_n40626_;
  assign new_n40628_ = ~new_n40083_ & ~new_n40182_;
  assign new_n40629_ = ~new_n38534_ & new_n39828_;
  assign new_n40630_ = ~new_n40628_ & ~new_n40629_;
  assign new_n40631_ = ~pi0219 & ~new_n40630_;
  assign new_n40632_ = pi0219 & ~new_n40182_;
  assign new_n40633_ = ~po1038 & ~new_n40632_;
  assign new_n40634_ = ~new_n40631_ & new_n40633_;
  assign new_n40635_ = new_n39854_ & ~new_n40634_;
  assign new_n40636_ = pi1152 & ~new_n40635_;
  assign new_n40637_ = ~new_n40627_ & new_n40636_;
  assign new_n40638_ = ~pi1150 & ~new_n40637_;
  assign new_n40639_ = ~new_n40621_ & new_n40638_;
  assign new_n40640_ = ~pi0219 & ~new_n40086_;
  assign new_n40641_ = ~new_n40310_ & new_n40640_;
  assign new_n40642_ = ~pi1153 & new_n40641_;
  assign new_n40643_ = pi0299 & new_n10485_;
  assign new_n40644_ = ~pi0219 & ~new_n40643_;
  assign new_n40645_ = new_n40195_ & ~new_n40644_;
  assign new_n40646_ = ~new_n40319_ & ~new_n40645_;
  assign new_n40647_ = ~new_n40642_ & ~new_n40646_;
  assign new_n40648_ = ~pi0211 & new_n40641_;
  assign new_n40649_ = ~new_n40088_ & ~new_n40648_;
  assign new_n40650_ = new_n39832_ & ~new_n40649_;
  assign new_n40651_ = ~new_n40647_ & new_n40650_;
  assign new_n40652_ = ~po1038 & ~new_n39768_;
  assign new_n40653_ = ~pi0299 & new_n39757_;
  assign new_n40654_ = ~new_n38423_ & ~new_n40615_;
  assign new_n40655_ = ~new_n40653_ & new_n40654_;
  assign new_n40656_ = new_n10729_ & ~new_n40172_;
  assign new_n40657_ = new_n40243_ & ~new_n40656_;
  assign new_n40658_ = ~new_n40655_ & new_n40657_;
  assign new_n40659_ = new_n40652_ & ~new_n40658_;
  assign new_n40660_ = new_n39854_ & ~new_n40659_;
  assign new_n40661_ = pi1152 & ~new_n40660_;
  assign new_n40662_ = ~new_n40651_ & new_n40661_;
  assign new_n40663_ = new_n39869_ & ~new_n40647_;
  assign new_n40664_ = pi1153 & new_n40489_;
  assign new_n40665_ = new_n39884_ & ~new_n40664_;
  assign new_n40666_ = ~pi1152 & ~new_n40665_;
  assign new_n40667_ = ~pi1151 & ~new_n40131_;
  assign new_n40668_ = ~pi1152 & ~new_n40667_;
  assign new_n40669_ = ~new_n40666_ & ~new_n40668_;
  assign new_n40670_ = ~new_n40663_ & ~new_n40669_;
  assign new_n40671_ = pi1150 & ~new_n40670_;
  assign new_n40672_ = ~new_n40662_ & new_n40671_;
  assign new_n40673_ = pi1149 & ~new_n40672_;
  assign new_n40674_ = ~new_n40639_ & new_n40673_;
  assign new_n40675_ = ~new_n40105_ & ~new_n40615_;
  assign new_n40676_ = pi0214 & new_n40675_;
  assign new_n40677_ = new_n40108_ & ~new_n40676_;
  assign new_n40678_ = ~pi0214 & new_n40675_;
  assign new_n40679_ = new_n40113_ & ~new_n40678_;
  assign new_n40680_ = ~new_n40677_ & ~new_n40679_;
  assign new_n40681_ = ~pi0219 & ~new_n40680_;
  assign new_n40682_ = new_n40123_ & ~new_n40681_;
  assign new_n40683_ = new_n39854_ & ~new_n40682_;
  assign new_n40684_ = pi0211 & ~new_n40066_;
  assign new_n40685_ = ~new_n11383_ & new_n38635_;
  assign new_n40686_ = ~new_n39713_ & ~new_n40685_;
  assign new_n40687_ = ~pi0211 & ~new_n38646_;
  assign new_n40688_ = ~new_n40686_ & new_n40687_;
  assign new_n40689_ = ~new_n40684_ & ~new_n40688_;
  assign new_n40690_ = ~pi0214 & new_n40689_;
  assign new_n40691_ = new_n40297_ & ~new_n40690_;
  assign new_n40692_ = pi0214 & new_n40689_;
  assign new_n40693_ = new_n40063_ & ~new_n40692_;
  assign new_n40694_ = ~pi0219 & ~new_n40693_;
  assign new_n40695_ = ~new_n40691_ & new_n40694_;
  assign new_n40696_ = new_n40294_ & ~new_n40695_;
  assign new_n40697_ = new_n39832_ & ~new_n40696_;
  assign new_n40698_ = pi1152 & ~new_n40697_;
  assign new_n40699_ = ~new_n40683_ & new_n40698_;
  assign new_n40700_ = ~new_n39736_ & ~new_n40684_;
  assign new_n40701_ = pi0214 & new_n40700_;
  assign new_n40702_ = new_n40062_ & ~new_n40070_;
  assign new_n40703_ = pi0212 & ~new_n40702_;
  assign new_n40704_ = ~new_n40701_ & new_n40703_;
  assign new_n40705_ = ~new_n40689_ & new_n40704_;
  assign new_n40706_ = ~new_n40071_ & ~new_n40688_;
  assign new_n40707_ = new_n40063_ & ~new_n40706_;
  assign new_n40708_ = ~pi0219 & ~new_n40707_;
  assign new_n40709_ = ~new_n40705_ & new_n40708_;
  assign new_n40710_ = new_n40294_ & ~new_n40709_;
  assign new_n40711_ = new_n39869_ & ~new_n40710_;
  assign new_n40712_ = ~new_n39885_ & new_n40100_;
  assign new_n40713_ = ~new_n38646_ & ~new_n40105_;
  assign new_n40714_ = ~pi0211 & ~new_n40713_;
  assign new_n40715_ = new_n39885_ & ~new_n40111_;
  assign new_n40716_ = ~new_n40714_ & new_n40715_;
  assign new_n40717_ = ~new_n40712_ & ~new_n40716_;
  assign new_n40718_ = ~po1038 & ~new_n40717_;
  assign new_n40719_ = new_n39884_ & ~new_n40718_;
  assign new_n40720_ = ~pi1152 & ~new_n40719_;
  assign new_n40721_ = ~new_n40711_ & new_n40720_;
  assign new_n40722_ = pi1150 & ~new_n40721_;
  assign new_n40723_ = ~new_n40699_ & new_n40722_;
  assign new_n40724_ = pi0219 & ~new_n39699_;
  assign new_n40725_ = ~po1038 & ~new_n40724_;
  assign new_n40726_ = new_n40526_ & ~new_n40530_;
  assign new_n40727_ = new_n40725_ & ~new_n40726_;
  assign new_n40728_ = ~new_n39919_ & new_n40725_;
  assign new_n40729_ = new_n39832_ & ~new_n40728_;
  assign new_n40730_ = ~new_n40727_ & new_n40729_;
  assign new_n40731_ = pi0299 & new_n39825_;
  assign new_n40732_ = ~new_n39828_ & new_n40731_;
  assign new_n40733_ = new_n39854_ & ~new_n40732_;
  assign new_n40734_ = pi1152 & ~new_n40733_;
  assign new_n40735_ = ~new_n40730_ & new_n40734_;
  assign new_n40736_ = new_n39869_ & ~new_n40728_;
  assign new_n40737_ = new_n40666_ & ~new_n40736_;
  assign new_n40738_ = ~pi1150 & ~new_n40737_;
  assign new_n40739_ = ~new_n40735_ & new_n40738_;
  assign new_n40740_ = ~pi1149 & ~new_n40739_;
  assign new_n40741_ = ~new_n40723_ & new_n40740_;
  assign new_n40742_ = ~new_n40674_ & ~new_n40741_;
  assign new_n40743_ = pi0213 & ~new_n40742_;
  assign new_n40744_ = ~new_n40124_ & new_n40522_;
  assign new_n40745_ = ~new_n40077_ & new_n40499_;
  assign new_n40746_ = pi1150 & ~new_n40745_;
  assign new_n40747_ = ~new_n40744_ & new_n40746_;
  assign new_n40748_ = ~pi1150 & pi1151;
  assign new_n40749_ = ~new_n40166_ & new_n40748_;
  assign new_n40750_ = ~pi1149 & ~new_n40749_;
  assign new_n40751_ = ~new_n40747_ & new_n40750_;
  assign new_n40752_ = ~new_n40160_ & new_n40554_;
  assign new_n40753_ = ~new_n40199_ & new_n40569_;
  assign new_n40754_ = ~pi1150 & ~new_n40753_;
  assign new_n40755_ = ~new_n40752_ & new_n40754_;
  assign new_n40756_ = ~pi1151 & new_n40134_;
  assign new_n40757_ = new_n40088_ & new_n40580_;
  assign new_n40758_ = pi1150 & ~new_n40757_;
  assign new_n40759_ = ~new_n40756_ & new_n40758_;
  assign new_n40760_ = pi1149 & ~new_n40759_;
  assign new_n40761_ = ~new_n40755_ & new_n40760_;
  assign new_n40762_ = ~new_n40751_ & ~new_n40761_;
  assign new_n40763_ = ~pi0213 & new_n40762_;
  assign new_n40764_ = ~pi0209 & ~new_n40763_;
  assign new_n40765_ = ~new_n40743_ & new_n40764_;
  assign new_n40766_ = ~new_n40606_ & ~new_n40765_;
  assign new_n40767_ = pi0230 & ~new_n40766_;
  assign new_n40768_ = ~pi0230 & ~pi0241;
  assign po0398 = ~new_n40767_ & ~new_n40768_;
  assign new_n40770_ = ~pi0230 & ~pi0242;
  assign new_n40771_ = pi0214 & ~new_n39371_;
  assign new_n40772_ = ~pi0214 & ~new_n40210_;
  assign new_n40773_ = ~new_n40771_ & ~new_n40772_;
  assign new_n40774_ = pi0212 & ~new_n40773_;
  assign new_n40775_ = ~pi0212 & new_n40211_;
  assign new_n40776_ = ~pi0219 & ~new_n40775_;
  assign new_n40777_ = ~new_n40774_ & new_n40776_;
  assign new_n40778_ = pi0219 & ~new_n38419_;
  assign new_n40779_ = new_n38416_ & ~new_n40778_;
  assign new_n40780_ = ~new_n40777_ & new_n40779_;
  assign new_n40781_ = ~pi0299 & ~new_n39388_;
  assign new_n40782_ = pi0199 & pi1144;
  assign new_n40783_ = ~pi0200 & ~new_n40782_;
  assign new_n40784_ = ~new_n39386_ & new_n40783_;
  assign new_n40785_ = new_n40781_ & ~new_n40784_;
  assign new_n40786_ = pi0207 & ~new_n40785_;
  assign new_n40787_ = ~new_n40332_ & new_n40783_;
  assign new_n40788_ = ~pi0299 & ~new_n40334_;
  assign new_n40789_ = ~new_n40787_ & new_n40788_;
  assign new_n40790_ = ~pi0207 & ~new_n40789_;
  assign new_n40791_ = pi0208 & ~new_n40790_;
  assign new_n40792_ = ~new_n40786_ & new_n40791_;
  assign new_n40793_ = new_n38449_ & new_n40789_;
  assign new_n40794_ = ~new_n40237_ & ~new_n40793_;
  assign new_n40795_ = ~new_n40792_ & new_n40794_;
  assign new_n40796_ = ~pi0211 & ~new_n40795_;
  assign new_n40797_ = ~new_n39561_ & ~new_n40793_;
  assign new_n40798_ = ~new_n40792_ & new_n40797_;
  assign new_n40799_ = pi0211 & ~new_n40798_;
  assign new_n40800_ = ~new_n40796_ & ~new_n40799_;
  assign new_n40801_ = ~pi0214 & new_n40800_;
  assign new_n40802_ = ~new_n38763_ & ~new_n40793_;
  assign new_n40803_ = ~new_n40792_ & new_n40802_;
  assign new_n40804_ = pi0211 & ~new_n40803_;
  assign new_n40805_ = ~pi0211 & ~new_n40798_;
  assign new_n40806_ = pi0214 & ~new_n40805_;
  assign new_n40807_ = ~new_n40804_ & new_n40806_;
  assign new_n40808_ = pi0212 & ~new_n40807_;
  assign new_n40809_ = ~new_n40801_ & new_n40808_;
  assign new_n40810_ = new_n38837_ & new_n40789_;
  assign new_n40811_ = ~new_n40792_ & ~new_n40810_;
  assign new_n40812_ = ~pi0214 & new_n40811_;
  assign new_n40813_ = ~pi0212 & ~new_n40812_;
  assign new_n40814_ = pi0214 & new_n40800_;
  assign new_n40815_ = new_n40813_ & ~new_n40814_;
  assign new_n40816_ = ~pi0219 & ~new_n40815_;
  assign new_n40817_ = ~new_n40809_ & new_n40816_;
  assign new_n40818_ = ~new_n38414_ & ~new_n40811_;
  assign new_n40819_ = pi0219 & ~new_n40818_;
  assign new_n40820_ = new_n38414_ & ~new_n40803_;
  assign new_n40821_ = new_n40819_ & ~new_n40820_;
  assign new_n40822_ = ~po1038 & ~new_n40821_;
  assign new_n40823_ = ~new_n40817_ & new_n40822_;
  assign new_n40824_ = ~new_n40780_ & ~new_n40823_;
  assign new_n40825_ = pi0213 & new_n40824_;
  assign new_n40826_ = pi0211 & ~new_n40810_;
  assign new_n40827_ = new_n38414_ & ~new_n38798_;
  assign new_n40828_ = ~new_n40793_ & new_n40827_;
  assign new_n40829_ = ~new_n40826_ & ~new_n40828_;
  assign new_n40830_ = pi0219 & ~new_n40829_;
  assign new_n40831_ = new_n38413_ & ~new_n40810_;
  assign new_n40832_ = new_n10729_ & ~new_n38460_;
  assign new_n40833_ = ~new_n38431_ & new_n38788_;
  assign new_n40834_ = ~new_n40832_ & ~new_n40833_;
  assign new_n40835_ = ~pi0219 & ~new_n40793_;
  assign new_n40836_ = ~new_n40834_ & new_n40835_;
  assign new_n40837_ = ~new_n40831_ & ~new_n40836_;
  assign new_n40838_ = ~new_n40830_ & new_n40837_;
  assign new_n40839_ = ~new_n40792_ & ~new_n40838_;
  assign new_n40840_ = ~po1038 & ~new_n40839_;
  assign new_n40841_ = ~pi0213 & ~new_n38430_;
  assign new_n40842_ = ~new_n40840_ & new_n40841_;
  assign new_n40843_ = ~new_n40825_ & ~new_n40842_;
  assign new_n40844_ = pi0209 & ~new_n40843_;
  assign new_n40845_ = ~pi0213 & ~new_n38476_;
  assign new_n40846_ = pi0219 & new_n38413_;
  assign new_n40847_ = ~new_n40778_ & ~new_n40846_;
  assign new_n40848_ = ~new_n40777_ & new_n40847_;
  assign new_n40849_ = pi0299 & ~new_n40848_;
  assign new_n40850_ = ~po1038 & ~new_n40849_;
  assign new_n40851_ = ~new_n38467_ & new_n40850_;
  assign new_n40852_ = ~new_n40780_ & ~new_n40851_;
  assign new_n40853_ = pi0213 & ~new_n40852_;
  assign new_n40854_ = ~pi0209 & ~new_n40853_;
  assign new_n40855_ = ~new_n40845_ & new_n40854_;
  assign new_n40856_ = ~new_n40844_ & ~new_n40855_;
  assign new_n40857_ = pi0230 & ~new_n40856_;
  assign po0399 = ~new_n40770_ & ~new_n40857_;
  assign new_n40859_ = pi0243 & ~pi1091;
  assign new_n40860_ = ~pi0083 & ~pi0085;
  assign new_n40861_ = pi0314 & ~new_n40860_;
  assign new_n40862_ = pi0802 & new_n40861_;
  assign new_n40863_ = pi0276 & new_n40862_;
  assign new_n40864_ = ~pi1091 & ~new_n40863_;
  assign new_n40865_ = pi0271 & ~new_n40864_;
  assign new_n40866_ = ~pi1091 & ~new_n40865_;
  assign new_n40867_ = pi0273 & ~new_n40866_;
  assign new_n40868_ = ~pi1091 & ~new_n40867_;
  assign new_n40869_ = ~pi0200 & ~new_n40868_;
  assign new_n40870_ = pi0199 & ~new_n40868_;
  assign new_n40871_ = ~pi0081 & new_n40860_;
  assign new_n40872_ = pi0314 & ~new_n40871_;
  assign new_n40873_ = pi0802 & new_n40872_;
  assign new_n40874_ = pi0276 & new_n40873_;
  assign new_n40875_ = ~pi1091 & new_n40874_;
  assign new_n40876_ = pi0271 & new_n40875_;
  assign new_n40877_ = pi0273 & new_n40876_;
  assign new_n40878_ = ~new_n40867_ & ~new_n40877_;
  assign new_n40879_ = ~pi1091 & new_n40878_;
  assign new_n40880_ = ~pi0199 & ~new_n40879_;
  assign new_n40881_ = ~new_n40870_ & ~new_n40880_;
  assign new_n40882_ = new_n40875_ & ~new_n40881_;
  assign new_n40883_ = ~pi0299 & ~new_n40882_;
  assign new_n40884_ = ~new_n40870_ & new_n40883_;
  assign new_n40885_ = ~new_n40869_ & new_n40884_;
  assign new_n40886_ = pi0299 & ~new_n40877_;
  assign new_n40887_ = ~new_n40885_ & ~new_n40886_;
  assign new_n40888_ = ~new_n40859_ & ~new_n40887_;
  assign new_n40889_ = ~pi0200 & ~new_n40875_;
  assign new_n40890_ = ~new_n40881_ & ~new_n40889_;
  assign new_n40891_ = ~pi0299 & ~new_n40890_;
  assign new_n40892_ = ~new_n40870_ & new_n40891_;
  assign new_n40893_ = ~pi1091 & new_n40863_;
  assign new_n40894_ = pi0271 & new_n40893_;
  assign new_n40895_ = pi0273 & new_n40894_;
  assign new_n40896_ = pi0299 & ~new_n40895_;
  assign new_n40897_ = ~new_n40869_ & new_n40883_;
  assign new_n40898_ = ~new_n40880_ & new_n40897_;
  assign new_n40899_ = ~new_n40896_ & ~new_n40898_;
  assign new_n40900_ = ~new_n40892_ & new_n40899_;
  assign new_n40901_ = pi0299 & new_n40868_;
  assign new_n40902_ = ~new_n40897_ & ~new_n40901_;
  assign new_n40903_ = pi0243 & ~new_n40902_;
  assign new_n40904_ = ~new_n40900_ & new_n40903_;
  assign new_n40905_ = pi1155 & ~new_n40904_;
  assign new_n40906_ = ~new_n40877_ & new_n40901_;
  assign new_n40907_ = ~new_n40898_ & ~new_n40906_;
  assign new_n40908_ = pi1155 & new_n40907_;
  assign new_n40909_ = ~new_n40905_ & ~new_n40908_;
  assign new_n40910_ = ~new_n40886_ & ~new_n40891_;
  assign new_n40911_ = ~pi0243 & new_n40910_;
  assign new_n40912_ = ~new_n40885_ & new_n40911_;
  assign new_n40913_ = ~new_n40909_ & ~new_n40912_;
  assign new_n40914_ = ~new_n40880_ & new_n40891_;
  assign new_n40915_ = ~new_n40885_ & ~new_n40914_;
  assign new_n40916_ = ~new_n40906_ & new_n40915_;
  assign new_n40917_ = ~pi0243 & ~new_n40916_;
  assign new_n40918_ = ~new_n40886_ & ~new_n40892_;
  assign new_n40919_ = pi0243 & ~new_n40898_;
  assign new_n40920_ = new_n40918_ & new_n40919_;
  assign new_n40921_ = ~new_n40917_ & ~new_n40920_;
  assign new_n40922_ = ~pi1155 & ~new_n40921_;
  assign new_n40923_ = ~new_n40913_ & ~new_n40922_;
  assign new_n40924_ = ~new_n40888_ & new_n40923_;
  assign new_n40925_ = pi1156 & ~new_n40924_;
  assign new_n40926_ = ~new_n40901_ & ~new_n40914_;
  assign new_n40927_ = ~pi0243 & ~new_n40926_;
  assign new_n40928_ = ~pi1155 & ~new_n40927_;
  assign new_n40929_ = ~new_n40883_ & ~new_n40886_;
  assign new_n40930_ = ~pi1155 & new_n40929_;
  assign new_n40931_ = ~new_n40928_ & ~new_n40930_;
  assign new_n40932_ = ~new_n40886_ & ~new_n40897_;
  assign new_n40933_ = pi0243 & new_n40932_;
  assign new_n40934_ = ~new_n40884_ & new_n40933_;
  assign new_n40935_ = ~new_n40931_ & ~new_n40934_;
  assign new_n40936_ = ~pi1156 & ~new_n40935_;
  assign new_n40937_ = ~new_n40891_ & ~new_n40906_;
  assign new_n40938_ = ~pi0243 & ~new_n40937_;
  assign new_n40939_ = pi1155 & ~new_n40938_;
  assign new_n40940_ = ~new_n40933_ & new_n40939_;
  assign new_n40941_ = new_n40936_ & ~new_n40940_;
  assign new_n40942_ = pi1157 & ~new_n40941_;
  assign new_n40943_ = ~new_n40925_ & new_n40942_;
  assign new_n40944_ = pi0243 & new_n40929_;
  assign new_n40945_ = ~pi0243 & ~pi1091;
  assign new_n40946_ = ~new_n40883_ & ~new_n40896_;
  assign new_n40947_ = new_n40945_ & ~new_n40946_;
  assign new_n40948_ = ~pi1155 & ~new_n40947_;
  assign new_n40949_ = ~new_n40930_ & ~new_n40948_;
  assign new_n40950_ = ~new_n40944_ & ~new_n40949_;
  assign new_n40951_ = ~pi1156 & ~new_n40950_;
  assign new_n40952_ = pi1155 & ~new_n40859_;
  assign new_n40953_ = new_n40870_ & new_n40952_;
  assign new_n40954_ = ~new_n40940_ & ~new_n40953_;
  assign new_n40955_ = new_n40951_ & new_n40954_;
  assign new_n40956_ = ~new_n40880_ & new_n40883_;
  assign new_n40957_ = ~new_n40906_ & ~new_n40956_;
  assign new_n40958_ = pi0243 & ~new_n40957_;
  assign new_n40959_ = ~new_n40884_ & ~new_n40886_;
  assign new_n40960_ = ~pi0243 & new_n40959_;
  assign new_n40961_ = ~new_n40958_ & ~new_n40960_;
  assign new_n40962_ = ~pi1155 & new_n40932_;
  assign new_n40963_ = ~new_n40875_ & new_n40962_;
  assign new_n40964_ = pi1156 & ~new_n40963_;
  assign new_n40965_ = new_n40961_ & new_n40964_;
  assign new_n40966_ = ~pi1157 & ~new_n40965_;
  assign new_n40967_ = ~new_n40955_ & new_n40966_;
  assign new_n40968_ = pi0211 & ~new_n40967_;
  assign new_n40969_ = ~new_n40943_ & new_n40968_;
  assign new_n40970_ = pi1156 & ~new_n40923_;
  assign new_n40971_ = ~new_n40897_ & ~new_n40906_;
  assign new_n40972_ = pi0243 & ~new_n40971_;
  assign new_n40973_ = ~new_n40911_ & ~new_n40972_;
  assign new_n40974_ = new_n40936_ & new_n40973_;
  assign new_n40975_ = pi1157 & ~new_n40974_;
  assign new_n40976_ = ~new_n40970_ & new_n40975_;
  assign new_n40977_ = new_n40961_ & new_n40973_;
  assign new_n40978_ = pi1155 & ~new_n40977_;
  assign new_n40979_ = new_n40951_ & ~new_n40978_;
  assign new_n40980_ = ~pi1155 & new_n40971_;
  assign new_n40981_ = ~new_n40910_ & new_n40980_;
  assign new_n40982_ = new_n40965_ & ~new_n40981_;
  assign new_n40983_ = ~pi1157 & ~new_n40982_;
  assign new_n40984_ = ~new_n40979_ & new_n40983_;
  assign new_n40985_ = ~pi0211 & ~new_n40984_;
  assign new_n40986_ = ~new_n40976_ & new_n40985_;
  assign new_n40987_ = ~pi0219 & ~new_n40986_;
  assign new_n40988_ = ~new_n40969_ & new_n40987_;
  assign new_n40989_ = pi0253 & pi0254;
  assign new_n40990_ = pi0267 & new_n40989_;
  assign new_n40991_ = ~pi0263 & new_n40990_;
  assign new_n40992_ = ~new_n40885_ & ~new_n40901_;
  assign new_n40993_ = ~pi0243 & new_n40992_;
  assign new_n40994_ = ~new_n40891_ & ~new_n40896_;
  assign new_n40995_ = new_n40993_ & new_n40994_;
  assign new_n40996_ = new_n40905_ & ~new_n40995_;
  assign new_n40997_ = pi0243 & ~new_n40900_;
  assign new_n40998_ = ~new_n40993_ & ~new_n40997_;
  assign new_n40999_ = ~new_n40888_ & ~new_n40927_;
  assign new_n41000_ = ~new_n40998_ & new_n40999_;
  assign new_n41001_ = ~pi1155 & ~new_n41000_;
  assign new_n41002_ = ~new_n40996_ & ~new_n41001_;
  assign new_n41003_ = pi1156 & ~new_n41002_;
  assign new_n41004_ = ~new_n40896_ & ~new_n40914_;
  assign new_n41005_ = ~pi0243 & ~new_n41004_;
  assign new_n41006_ = pi0243 & ~new_n40884_;
  assign new_n41007_ = ~pi1155 & ~new_n41006_;
  assign new_n41008_ = ~new_n41005_ & new_n41007_;
  assign new_n41009_ = ~pi0243 & pi1155;
  assign new_n41010_ = new_n40994_ & new_n41009_;
  assign new_n41011_ = ~pi1156 & ~new_n41010_;
  assign new_n41012_ = ~new_n40903_ & new_n41011_;
  assign new_n41013_ = ~new_n41008_ & new_n41012_;
  assign new_n41014_ = new_n38478_ & ~new_n41013_;
  assign new_n41015_ = ~new_n41003_ & new_n41014_;
  assign new_n41016_ = pi0243 & new_n40899_;
  assign new_n41017_ = new_n40939_ & ~new_n41016_;
  assign new_n41018_ = ~new_n40928_ & ~new_n41017_;
  assign new_n41019_ = ~new_n40998_ & ~new_n41018_;
  assign new_n41020_ = pi1156 & ~new_n41019_;
  assign new_n41021_ = ~new_n40896_ & ~new_n40897_;
  assign new_n41022_ = pi0243 & new_n41021_;
  assign new_n41023_ = ~new_n40938_ & ~new_n41022_;
  assign new_n41024_ = pi1155 & ~new_n41023_;
  assign new_n41025_ = ~new_n40884_ & new_n41021_;
  assign new_n41026_ = pi0243 & new_n41025_;
  assign new_n41027_ = ~new_n40927_ & ~new_n41026_;
  assign new_n41028_ = ~new_n41024_ & new_n41027_;
  assign new_n41029_ = ~pi1156 & ~new_n41028_;
  assign new_n41030_ = new_n39400_ & ~new_n41029_;
  assign new_n41031_ = ~new_n41020_ & new_n41030_;
  assign new_n41032_ = ~new_n40896_ & ~new_n40956_;
  assign new_n41033_ = pi1155 & new_n41032_;
  assign new_n41034_ = ~new_n40891_ & new_n41032_;
  assign new_n41035_ = ~new_n41033_ & ~new_n41034_;
  assign new_n41036_ = pi0243 & ~new_n41035_;
  assign new_n41037_ = ~new_n40884_ & ~new_n40901_;
  assign new_n41038_ = ~pi0243 & ~new_n41037_;
  assign new_n41039_ = ~new_n40963_ & new_n41038_;
  assign new_n41040_ = ~new_n41036_ & ~new_n41039_;
  assign new_n41041_ = pi1156 & ~new_n41040_;
  assign new_n41042_ = ~new_n40956_ & new_n41022_;
  assign new_n41043_ = ~new_n40892_ & ~new_n40901_;
  assign new_n41044_ = ~pi0243 & ~new_n41043_;
  assign new_n41045_ = pi1155 & ~new_n41044_;
  assign new_n41046_ = ~new_n41042_ & new_n41045_;
  assign new_n41047_ = pi0243 & new_n40946_;
  assign new_n41048_ = new_n40948_ & ~new_n41047_;
  assign new_n41049_ = ~pi1156 & ~new_n41048_;
  assign new_n41050_ = ~new_n41046_ & new_n41049_;
  assign new_n41051_ = ~pi1157 & ~new_n41050_;
  assign new_n41052_ = ~new_n41041_ & new_n41051_;
  assign new_n41053_ = ~new_n41031_ & ~new_n41052_;
  assign new_n41054_ = ~new_n41015_ & new_n41053_;
  assign new_n41055_ = pi0219 & ~new_n41054_;
  assign new_n41056_ = new_n40991_ & ~new_n41055_;
  assign new_n41057_ = ~new_n40988_ & new_n41056_;
  assign new_n41058_ = ~pi0299 & pi1091;
  assign new_n41059_ = new_n38852_ & new_n41058_;
  assign new_n41060_ = ~new_n40945_ & ~new_n41059_;
  assign new_n41061_ = pi1156 & ~new_n41060_;
  assign new_n41062_ = pi1091 & ~new_n38955_;
  assign new_n41063_ = new_n39519_ & new_n41062_;
  assign new_n41064_ = ~new_n41061_ & ~new_n41063_;
  assign new_n41065_ = ~pi0299 & new_n38607_;
  assign new_n41066_ = pi1091 & ~new_n41065_;
  assign new_n41067_ = ~new_n40859_ & ~new_n41066_;
  assign new_n41068_ = ~pi1155 & ~new_n40945_;
  assign new_n41069_ = ~new_n40859_ & ~new_n41068_;
  assign new_n41070_ = new_n38548_ & new_n41069_;
  assign new_n41071_ = ~new_n41067_ & ~new_n41070_;
  assign new_n41072_ = ~pi1156 & ~new_n41071_;
  assign new_n41073_ = new_n41064_ & ~new_n41072_;
  assign new_n41074_ = pi1157 & ~new_n41073_;
  assign new_n41075_ = pi0199 & pi1091;
  assign new_n41076_ = ~pi0299 & new_n41075_;
  assign new_n41077_ = new_n40952_ & ~new_n41076_;
  assign new_n41078_ = pi1156 & ~new_n41077_;
  assign new_n41079_ = ~pi1155 & ~new_n40859_;
  assign new_n41080_ = ~new_n11444_ & new_n41058_;
  assign new_n41081_ = new_n41079_ & ~new_n41080_;
  assign new_n41082_ = new_n41078_ & ~new_n41081_;
  assign new_n41083_ = ~new_n41062_ & new_n41069_;
  assign new_n41084_ = ~pi1156 & ~new_n41083_;
  assign new_n41085_ = ~pi1157 & ~new_n41084_;
  assign new_n41086_ = ~new_n41082_ & new_n41085_;
  assign new_n41087_ = ~new_n41074_ & ~new_n41086_;
  assign new_n41088_ = pi0211 & ~new_n41087_;
  assign new_n41089_ = new_n41060_ & new_n41078_;
  assign new_n41090_ = ~pi1155 & new_n41067_;
  assign new_n41091_ = pi0200 & pi1091;
  assign new_n41092_ = ~pi0299 & new_n41091_;
  assign new_n41093_ = new_n40952_ & ~new_n41092_;
  assign new_n41094_ = ~pi1156 & ~new_n41093_;
  assign new_n41095_ = ~new_n41090_ & new_n41094_;
  assign new_n41096_ = ~new_n41089_ & ~new_n41095_;
  assign new_n41097_ = pi1157 & ~new_n41096_;
  assign new_n41098_ = pi1091 & ~new_n11445_;
  assign new_n41099_ = new_n41079_ & ~new_n41098_;
  assign new_n41100_ = ~new_n41077_ & ~new_n41099_;
  assign new_n41101_ = pi0200 & ~pi1156;
  assign new_n41102_ = new_n41058_ & new_n41101_;
  assign new_n41103_ = ~new_n41100_ & ~new_n41102_;
  assign new_n41104_ = ~pi1157 & ~new_n41103_;
  assign new_n41105_ = ~pi0211 & ~new_n41104_;
  assign new_n41106_ = ~new_n41097_ & new_n41105_;
  assign new_n41107_ = ~new_n41088_ & ~new_n41106_;
  assign new_n41108_ = ~pi0219 & ~new_n41107_;
  assign new_n41109_ = new_n39400_ & ~new_n41061_;
  assign new_n41110_ = ~new_n41072_ & new_n41109_;
  assign new_n41111_ = pi0219 & ~new_n41110_;
  assign new_n41112_ = pi0299 & pi1091;
  assign new_n41113_ = new_n41103_ & ~new_n41112_;
  assign new_n41114_ = ~pi1157 & ~new_n41113_;
  assign new_n41115_ = pi1091 & new_n38608_;
  assign new_n41116_ = new_n41079_ & ~new_n41115_;
  assign new_n41117_ = ~new_n41093_ & ~new_n41116_;
  assign new_n41118_ = ~pi1156 & ~new_n41117_;
  assign new_n41119_ = new_n38478_ & ~new_n41118_;
  assign new_n41120_ = new_n41064_ & new_n41119_;
  assign new_n41121_ = ~new_n41114_ & ~new_n41120_;
  assign new_n41122_ = new_n41111_ & new_n41121_;
  assign new_n41123_ = ~new_n41108_ & ~new_n41122_;
  assign new_n41124_ = ~new_n40991_ & ~new_n41123_;
  assign new_n41125_ = ~po1038 & ~new_n41124_;
  assign new_n41126_ = ~new_n41057_ & new_n41125_;
  assign new_n41127_ = ~pi0243 & new_n40868_;
  assign new_n41128_ = pi0243 & new_n40895_;
  assign new_n41129_ = new_n38478_ & ~new_n40859_;
  assign new_n41130_ = ~new_n40893_ & new_n41129_;
  assign new_n41131_ = ~new_n41128_ & ~new_n41130_;
  assign new_n41132_ = ~new_n41127_ & new_n41131_;
  assign new_n41133_ = pi0219 & ~new_n41132_;
  assign new_n41134_ = new_n40859_ & new_n40878_;
  assign new_n41135_ = ~pi0243 & new_n40877_;
  assign new_n41136_ = ~new_n38479_ & ~new_n38487_;
  assign new_n41137_ = pi1091 & new_n41136_;
  assign new_n41138_ = ~pi0219 & ~new_n41137_;
  assign new_n41139_ = ~new_n41135_ & new_n41138_;
  assign new_n41140_ = ~new_n41134_ & new_n41139_;
  assign new_n41141_ = ~new_n41133_ & ~new_n41140_;
  assign new_n41142_ = new_n40991_ & ~new_n41141_;
  assign new_n41143_ = ~pi0219 & ~new_n41136_;
  assign new_n41144_ = pi1157 & new_n38519_;
  assign new_n41145_ = ~new_n41143_ & ~new_n41144_;
  assign new_n41146_ = pi1091 & ~new_n41145_;
  assign new_n41147_ = ~new_n40945_ & ~new_n41146_;
  assign new_n41148_ = ~new_n40991_ & ~new_n41147_;
  assign new_n41149_ = po1038 & ~new_n41148_;
  assign new_n41150_ = ~new_n41142_ & new_n41149_;
  assign new_n41151_ = pi0272 & pi0283;
  assign new_n41152_ = pi0275 & new_n41151_;
  assign new_n41153_ = pi0268 & new_n41152_;
  assign new_n41154_ = ~new_n41150_ & new_n41153_;
  assign new_n41155_ = ~new_n41126_ & new_n41154_;
  assign new_n41156_ = ~po1038 & new_n41123_;
  assign new_n41157_ = po1038 & new_n41147_;
  assign new_n41158_ = ~new_n41153_ & ~new_n41157_;
  assign new_n41159_ = ~new_n41156_ & new_n41158_;
  assign new_n41160_ = ~pi0230 & ~new_n41159_;
  assign new_n41161_ = ~new_n41155_ & new_n41160_;
  assign new_n41162_ = pi0199 & ~new_n39572_;
  assign new_n41163_ = ~new_n38851_ & ~new_n41101_;
  assign new_n41164_ = ~new_n41162_ & new_n41163_;
  assign new_n41165_ = new_n16479_ & new_n41164_;
  assign new_n41166_ = ~new_n16479_ & ~new_n41145_;
  assign new_n41167_ = pi0230 & ~new_n41166_;
  assign new_n41168_ = ~new_n41165_ & new_n41167_;
  assign po0400 = ~new_n41161_ & ~new_n41168_;
  assign new_n41170_ = ~pi0230 & ~pi0244;
  assign new_n41171_ = pi0213 & ~new_n40473_;
  assign new_n41172_ = ~new_n38761_ & new_n40362_;
  assign new_n41173_ = ~new_n40467_ & ~new_n41172_;
  assign new_n41174_ = ~pi0214 & new_n41173_;
  assign new_n41175_ = new_n38420_ & new_n40313_;
  assign new_n41176_ = pi0212 & ~new_n41175_;
  assign new_n41177_ = ~new_n41174_ & new_n41176_;
  assign new_n41178_ = ~new_n40367_ & new_n41177_;
  assign new_n41179_ = ~new_n40367_ & ~new_n41173_;
  assign new_n41180_ = pi0214 & ~new_n41179_;
  assign new_n41181_ = new_n40438_ & ~new_n41180_;
  assign new_n41182_ = ~pi0219 & ~new_n41181_;
  assign new_n41183_ = ~new_n41178_ & new_n41182_;
  assign new_n41184_ = ~pi0211 & ~new_n38731_;
  assign new_n41185_ = ~new_n40441_ & new_n41184_;
  assign new_n41186_ = ~new_n40449_ & ~new_n41185_;
  assign new_n41187_ = new_n40447_ & ~new_n41186_;
  assign new_n41188_ = new_n40343_ & ~new_n41187_;
  assign new_n41189_ = ~new_n41183_ & new_n41188_;
  assign new_n41190_ = ~new_n40357_ & new_n41177_;
  assign new_n41191_ = pi0214 & new_n41173_;
  assign new_n41192_ = new_n40383_ & ~new_n41191_;
  assign new_n41193_ = ~pi0219 & ~new_n41192_;
  assign new_n41194_ = ~new_n41190_ & new_n41193_;
  assign new_n41195_ = pi0299 & new_n39377_;
  assign new_n41196_ = pi1147 & ~new_n41195_;
  assign new_n41197_ = new_n40361_ & new_n41196_;
  assign new_n41198_ = ~new_n41194_ & new_n41197_;
  assign new_n41199_ = ~pi0213 & ~new_n39379_;
  assign new_n41200_ = ~new_n41198_ & new_n41199_;
  assign new_n41201_ = ~new_n41189_ & new_n41200_;
  assign new_n41202_ = ~new_n41171_ & ~new_n41201_;
  assign new_n41203_ = pi0209 & ~new_n41202_;
  assign new_n41204_ = new_n40222_ & ~new_n40228_;
  assign new_n41205_ = ~new_n40235_ & ~new_n41204_;
  assign new_n41206_ = new_n40222_ & ~new_n40227_;
  assign new_n41207_ = new_n10729_ & ~new_n40244_;
  assign new_n41208_ = ~new_n10729_ & new_n40239_;
  assign new_n41209_ = new_n38794_ & ~new_n41208_;
  assign new_n41210_ = ~new_n41207_ & new_n41209_;
  assign new_n41211_ = ~new_n41206_ & new_n41210_;
  assign new_n41212_ = ~new_n39392_ & ~new_n40258_;
  assign new_n41213_ = ~new_n41211_ & new_n41212_;
  assign new_n41214_ = ~po1038 & ~new_n41213_;
  assign new_n41215_ = ~new_n41205_ & ~new_n41214_;
  assign new_n41216_ = pi0213 & ~new_n41215_;
  assign new_n41217_ = ~pi0213 & ~new_n39398_;
  assign new_n41218_ = ~pi0209 & ~new_n41217_;
  assign new_n41219_ = ~new_n41216_ & new_n41218_;
  assign new_n41220_ = ~new_n41203_ & ~new_n41219_;
  assign new_n41221_ = pi0230 & ~new_n41220_;
  assign po0401 = ~new_n41170_ & ~new_n41221_;
  assign new_n41223_ = pi1146 & new_n39830_;
  assign new_n41224_ = pi1147 & ~new_n39826_;
  assign new_n41225_ = ~new_n41223_ & new_n41224_;
  assign new_n41226_ = ~new_n38413_ & new_n40796_;
  assign new_n41227_ = new_n40819_ & ~new_n41226_;
  assign new_n41228_ = ~po1038 & ~new_n41227_;
  assign new_n41229_ = ~pi0299 & new_n40798_;
  assign new_n41230_ = ~pi0211 & ~new_n41229_;
  assign new_n41231_ = pi0211 & ~new_n40795_;
  assign new_n41232_ = ~new_n41230_ & ~new_n41231_;
  assign new_n41233_ = pi0214 & ~new_n41232_;
  assign new_n41234_ = ~pi0214 & ~new_n41229_;
  assign new_n41235_ = ~new_n41233_ & ~new_n41234_;
  assign new_n41236_ = pi0212 & ~new_n41235_;
  assign new_n41237_ = new_n40813_ & ~new_n41229_;
  assign new_n41238_ = ~pi0219 & ~new_n41237_;
  assign new_n41239_ = ~new_n41236_ & new_n41238_;
  assign new_n41240_ = new_n41228_ & ~new_n41239_;
  assign new_n41241_ = new_n41225_ & ~new_n41240_;
  assign new_n41242_ = ~pi1147 & ~new_n41223_;
  assign new_n41243_ = new_n39826_ & ~new_n40140_;
  assign new_n41244_ = new_n41242_ & ~new_n41243_;
  assign new_n41245_ = pi0214 & ~new_n40238_;
  assign new_n41246_ = ~pi0299 & ~new_n40800_;
  assign new_n41247_ = new_n41245_ & ~new_n41246_;
  assign new_n41248_ = pi0212 & ~new_n41247_;
  assign new_n41249_ = new_n40811_ & ~new_n41230_;
  assign new_n41250_ = ~pi0214 & new_n41249_;
  assign new_n41251_ = new_n41248_ & ~new_n41250_;
  assign new_n41252_ = new_n40813_ & ~new_n41249_;
  assign new_n41253_ = ~pi0219 & ~new_n41252_;
  assign new_n41254_ = ~new_n41251_ & new_n41253_;
  assign new_n41255_ = new_n41228_ & ~new_n41254_;
  assign new_n41256_ = new_n41244_ & ~new_n41255_;
  assign new_n41257_ = pi1148 & ~new_n41256_;
  assign new_n41258_ = ~new_n41241_ & new_n41257_;
  assign new_n41259_ = ~new_n40812_ & new_n41248_;
  assign new_n41260_ = ~pi0212 & ~new_n40811_;
  assign new_n41261_ = ~pi0219 & ~new_n41260_;
  assign new_n41262_ = ~new_n41259_ & new_n41261_;
  assign new_n41263_ = new_n41228_ & ~new_n41262_;
  assign new_n41264_ = new_n41242_ & ~new_n41263_;
  assign new_n41265_ = ~new_n40420_ & ~new_n41225_;
  assign new_n41266_ = ~new_n13061_ & new_n40811_;
  assign new_n41267_ = ~pi0214 & ~new_n41266_;
  assign new_n41268_ = ~new_n41233_ & ~new_n41267_;
  assign new_n41269_ = pi0212 & ~new_n41268_;
  assign new_n41270_ = new_n40813_ & ~new_n41266_;
  assign new_n41271_ = ~pi0219 & ~new_n41270_;
  assign new_n41272_ = ~new_n41269_ & new_n41271_;
  assign new_n41273_ = new_n41228_ & ~new_n41272_;
  assign new_n41274_ = ~new_n41265_ & ~new_n41273_;
  assign new_n41275_ = ~pi1148 & ~new_n41274_;
  assign new_n41276_ = ~new_n41264_ & new_n41275_;
  assign new_n41277_ = ~new_n41258_ & ~new_n41276_;
  assign new_n41278_ = pi0213 & ~new_n41277_;
  assign new_n41279_ = ~pi0213 & ~new_n40824_;
  assign new_n41280_ = ~pi0209 & ~new_n41279_;
  assign new_n41281_ = ~new_n41278_ & new_n41280_;
  assign new_n41282_ = pi0199 & pi1146;
  assign new_n41283_ = new_n38607_ & ~new_n41282_;
  assign new_n41284_ = new_n40339_ & ~new_n41283_;
  assign new_n41285_ = pi0208 & new_n41284_;
  assign new_n41286_ = ~pi0207 & ~new_n41285_;
  assign new_n41287_ = new_n39635_ & ~new_n41283_;
  assign new_n41288_ = ~new_n41286_ & new_n41287_;
  assign new_n41289_ = ~pi0208 & new_n40237_;
  assign new_n41290_ = ~pi0200 & ~new_n41282_;
  assign new_n41291_ = new_n40339_ & ~new_n41290_;
  assign new_n41292_ = pi0207 & new_n41291_;
  assign new_n41293_ = pi1146 & ~new_n38608_;
  assign new_n41294_ = ~new_n41292_ & ~new_n41293_;
  assign new_n41295_ = pi0208 & ~new_n41294_;
  assign new_n41296_ = ~new_n41289_ & ~new_n41295_;
  assign new_n41297_ = ~new_n41288_ & new_n41296_;
  assign new_n41298_ = ~pi0299 & ~new_n41297_;
  assign new_n41299_ = ~pi0214 & ~new_n41298_;
  assign new_n41300_ = ~pi0212 & ~new_n41299_;
  assign new_n41301_ = ~new_n10624_ & ~new_n39636_;
  assign new_n41302_ = new_n41291_ & ~new_n41301_;
  assign new_n41303_ = pi0211 & ~new_n41302_;
  assign new_n41304_ = ~pi0299 & ~new_n41291_;
  assign new_n41305_ = ~new_n41297_ & ~new_n41304_;
  assign new_n41306_ = ~pi0299 & ~new_n41305_;
  assign new_n41307_ = ~pi0211 & new_n41306_;
  assign new_n41308_ = ~new_n41303_ & ~new_n41307_;
  assign new_n41309_ = ~new_n41298_ & ~new_n41308_;
  assign new_n41310_ = new_n41300_ & ~new_n41309_;
  assign new_n41311_ = ~pi0219 & ~new_n41310_;
  assign new_n41312_ = new_n41245_ & ~new_n41298_;
  assign new_n41313_ = ~pi0214 & new_n41309_;
  assign new_n41314_ = pi0212 & ~new_n41313_;
  assign new_n41315_ = ~new_n41312_ & new_n41314_;
  assign new_n41316_ = new_n41311_ & ~new_n41315_;
  assign new_n41317_ = ~new_n38414_ & new_n41298_;
  assign new_n41318_ = pi0219 & ~new_n41317_;
  assign new_n41319_ = new_n38414_ & ~new_n41297_;
  assign new_n41320_ = new_n41318_ & ~new_n41319_;
  assign new_n41321_ = ~po1038 & ~new_n41320_;
  assign new_n41322_ = ~new_n41316_ & new_n41321_;
  assign new_n41323_ = new_n41244_ & ~new_n41322_;
  assign new_n41324_ = new_n38539_ & ~new_n41283_;
  assign new_n41325_ = ~new_n10624_ & ~new_n41324_;
  assign new_n41326_ = pi0207 & new_n41284_;
  assign new_n41327_ = ~new_n38837_ & ~new_n41326_;
  assign new_n41328_ = ~new_n41325_ & ~new_n41327_;
  assign new_n41329_ = ~pi0214 & ~new_n41328_;
  assign new_n41330_ = ~pi0212 & ~new_n41329_;
  assign new_n41331_ = new_n38539_ & ~new_n41290_;
  assign new_n41332_ = ~pi0207 & new_n41331_;
  assign new_n41333_ = ~new_n40237_ & ~new_n41332_;
  assign new_n41334_ = ~new_n41326_ & new_n41333_;
  assign new_n41335_ = pi0208 & ~new_n41334_;
  assign new_n41336_ = ~pi0299 & new_n41335_;
  assign new_n41337_ = new_n38449_ & new_n41324_;
  assign new_n41338_ = ~new_n41285_ & ~new_n41337_;
  assign new_n41339_ = ~new_n41336_ & new_n41338_;
  assign new_n41340_ = ~pi0299 & new_n41339_;
  assign new_n41341_ = new_n41330_ & ~new_n41340_;
  assign new_n41342_ = ~pi0219 & ~new_n41341_;
  assign new_n41343_ = pi0212 & ~new_n41340_;
  assign new_n41344_ = ~new_n40237_ & new_n41339_;
  assign new_n41345_ = new_n10484_ & new_n41344_;
  assign new_n41346_ = new_n41343_ & ~new_n41345_;
  assign new_n41347_ = new_n41342_ & ~new_n41346_;
  assign new_n41348_ = ~new_n38414_ & new_n41328_;
  assign new_n41349_ = pi0219 & ~new_n41348_;
  assign new_n41350_ = new_n38414_ & ~new_n41344_;
  assign new_n41351_ = new_n41349_ & ~new_n41350_;
  assign new_n41352_ = ~po1038 & ~new_n41351_;
  assign new_n41353_ = ~new_n41347_ & new_n41352_;
  assign new_n41354_ = new_n41225_ & ~new_n41353_;
  assign new_n41355_ = pi1148 & ~new_n41354_;
  assign new_n41356_ = ~new_n41323_ & new_n41355_;
  assign new_n41357_ = ~new_n10624_ & ~new_n41331_;
  assign new_n41358_ = ~new_n41327_ & ~new_n41357_;
  assign new_n41359_ = ~new_n13061_ & ~new_n41358_;
  assign new_n41360_ = pi0214 & ~new_n41359_;
  assign new_n41361_ = ~pi0214 & new_n41358_;
  assign new_n41362_ = ~pi0212 & ~new_n41361_;
  assign new_n41363_ = ~new_n41360_ & new_n41362_;
  assign new_n41364_ = ~pi0214 & ~new_n41359_;
  assign new_n41365_ = new_n38449_ & new_n41331_;
  assign new_n41366_ = ~new_n41289_ & ~new_n41365_;
  assign new_n41367_ = ~new_n41335_ & new_n41366_;
  assign new_n41368_ = ~pi0299 & new_n41367_;
  assign new_n41369_ = pi0214 & ~new_n41368_;
  assign new_n41370_ = ~pi0211 & ~new_n41340_;
  assign new_n41371_ = ~new_n41328_ & ~new_n41370_;
  assign new_n41372_ = new_n41369_ & ~new_n41371_;
  assign new_n41373_ = pi0212 & ~new_n41372_;
  assign new_n41374_ = ~new_n41364_ & new_n41373_;
  assign new_n41375_ = ~new_n41363_ & ~new_n41374_;
  assign new_n41376_ = ~pi0219 & ~new_n41375_;
  assign new_n41377_ = ~pi1146 & ~new_n38717_;
  assign new_n41378_ = new_n40310_ & ~new_n41377_;
  assign new_n41379_ = new_n41376_ & ~new_n41378_;
  assign new_n41380_ = ~new_n38413_ & new_n41358_;
  assign new_n41381_ = ~new_n38414_ & ~new_n41380_;
  assign new_n41382_ = ~new_n41367_ & ~new_n41381_;
  assign new_n41383_ = ~pi0212 & new_n41361_;
  assign new_n41384_ = pi0219 & ~new_n41383_;
  assign new_n41385_ = ~new_n41382_ & new_n41384_;
  assign new_n41386_ = ~po1038 & ~new_n41385_;
  assign new_n41387_ = ~new_n41379_ & new_n41386_;
  assign new_n41388_ = ~new_n41265_ & ~new_n41387_;
  assign new_n41389_ = ~new_n40643_ & ~new_n41298_;
  assign new_n41390_ = ~new_n41294_ & ~new_n41389_;
  assign new_n41391_ = ~pi0219 & ~new_n41390_;
  assign new_n41392_ = pi0219 & ~new_n41302_;
  assign new_n41393_ = ~new_n38970_ & ~new_n41392_;
  assign new_n41394_ = ~new_n38413_ & ~new_n41303_;
  assign new_n41395_ = new_n41305_ & new_n41394_;
  assign new_n41396_ = ~new_n41393_ & ~new_n41395_;
  assign new_n41397_ = ~po1038 & ~new_n41396_;
  assign new_n41398_ = ~new_n41391_ & new_n41397_;
  assign new_n41399_ = new_n41242_ & ~new_n41398_;
  assign new_n41400_ = ~pi1148 & ~new_n41399_;
  assign new_n41401_ = ~new_n41388_ & new_n41400_;
  assign new_n41402_ = ~new_n41356_ & ~new_n41401_;
  assign new_n41403_ = pi0213 & ~new_n41402_;
  assign new_n41404_ = ~pi0214 & new_n41302_;
  assign new_n41405_ = ~new_n40244_ & ~new_n41298_;
  assign new_n41406_ = pi0214 & ~new_n41306_;
  assign new_n41407_ = ~new_n41405_ & new_n41406_;
  assign new_n41408_ = ~new_n41404_ & ~new_n41407_;
  assign new_n41409_ = ~pi0212 & ~new_n41408_;
  assign new_n41410_ = pi0299 & ~new_n40773_;
  assign new_n41411_ = ~new_n41298_ & ~new_n41410_;
  assign new_n41412_ = pi0212 & ~new_n41411_;
  assign new_n41413_ = ~new_n41304_ & new_n41412_;
  assign new_n41414_ = ~pi0219 & ~new_n41413_;
  assign new_n41415_ = ~new_n41409_ & new_n41414_;
  assign new_n41416_ = ~new_n38761_ & ~new_n41306_;
  assign new_n41417_ = ~pi0211 & ~new_n41416_;
  assign new_n41418_ = new_n41394_ & ~new_n41417_;
  assign new_n41419_ = ~new_n41393_ & ~new_n41418_;
  assign new_n41420_ = new_n40343_ & ~new_n41419_;
  assign new_n41421_ = ~new_n41415_ & new_n41420_;
  assign new_n41422_ = ~new_n38763_ & new_n41339_;
  assign new_n41423_ = ~new_n41368_ & ~new_n41422_;
  assign new_n41424_ = ~pi0211 & ~new_n41423_;
  assign new_n41425_ = ~new_n41381_ & ~new_n41424_;
  assign new_n41426_ = new_n41384_ & ~new_n41425_;
  assign new_n41427_ = pi1147 & ~po1038;
  assign new_n41428_ = ~new_n40244_ & new_n41339_;
  assign new_n41429_ = new_n41369_ & ~new_n41428_;
  assign new_n41430_ = ~new_n41361_ & ~new_n41429_;
  assign new_n41431_ = ~pi0212 & ~new_n41430_;
  assign new_n41432_ = new_n41339_ & ~new_n41410_;
  assign new_n41433_ = pi0212 & ~new_n41432_;
  assign new_n41434_ = ~new_n41368_ & new_n41433_;
  assign new_n41435_ = ~pi0219 & ~new_n41434_;
  assign new_n41436_ = ~new_n41431_ & new_n41435_;
  assign new_n41437_ = new_n41427_ & ~new_n41436_;
  assign new_n41438_ = ~new_n41426_ & new_n41437_;
  assign new_n41439_ = ~pi1148 & ~new_n40780_;
  assign new_n41440_ = ~new_n41438_ & new_n41439_;
  assign new_n41441_ = ~new_n41421_ & new_n41440_;
  assign new_n41442_ = new_n41300_ & ~new_n41405_;
  assign new_n41443_ = ~pi0219 & ~new_n41412_;
  assign new_n41444_ = ~new_n41442_ & new_n41443_;
  assign new_n41445_ = ~pi0299 & new_n41297_;
  assign new_n41446_ = new_n38414_ & ~new_n41445_;
  assign new_n41447_ = ~new_n38761_ & new_n41446_;
  assign new_n41448_ = new_n41318_ & ~new_n41447_;
  assign new_n41449_ = new_n40343_ & ~new_n41448_;
  assign new_n41450_ = ~new_n41444_ & new_n41449_;
  assign new_n41451_ = pi0214 & new_n41428_;
  assign new_n41452_ = new_n41330_ & ~new_n41451_;
  assign new_n41453_ = ~pi0219 & ~new_n41433_;
  assign new_n41454_ = ~new_n41452_ & new_n41453_;
  assign new_n41455_ = new_n38414_ & ~new_n41422_;
  assign new_n41456_ = new_n41349_ & ~new_n41455_;
  assign new_n41457_ = new_n41427_ & ~new_n41456_;
  assign new_n41458_ = ~new_n41454_ & new_n41457_;
  assign new_n41459_ = pi1148 & ~new_n40780_;
  assign new_n41460_ = ~new_n41458_ & new_n41459_;
  assign new_n41461_ = ~new_n41450_ & new_n41460_;
  assign new_n41462_ = ~pi0213 & ~new_n41461_;
  assign new_n41463_ = ~new_n41441_ & new_n41462_;
  assign new_n41464_ = pi0209 & ~new_n41463_;
  assign new_n41465_ = ~new_n41403_ & new_n41464_;
  assign new_n41466_ = ~new_n41281_ & ~new_n41465_;
  assign new_n41467_ = pi0230 & ~new_n41466_;
  assign new_n41468_ = ~pi0230 & ~pi0245;
  assign po0402 = ~new_n41467_ & ~new_n41468_;
  assign new_n41470_ = ~new_n41225_ & ~new_n41244_;
  assign new_n41471_ = pi0219 & ~new_n40237_;
  assign new_n41472_ = new_n40084_ & ~new_n41471_;
  assign new_n41473_ = new_n40131_ & ~new_n40181_;
  assign new_n41474_ = ~new_n41472_ & ~new_n41473_;
  assign new_n41475_ = ~new_n40183_ & ~new_n40253_;
  assign new_n41476_ = new_n38423_ & ~new_n41475_;
  assign new_n41477_ = ~new_n40628_ & ~new_n41476_;
  assign new_n41478_ = ~pi0219 & ~new_n41477_;
  assign new_n41479_ = ~new_n41474_ & ~new_n41478_;
  assign new_n41480_ = ~new_n41470_ & ~new_n41479_;
  assign new_n41481_ = ~new_n40184_ & ~new_n40193_;
  assign new_n41482_ = new_n41244_ & ~new_n41481_;
  assign new_n41483_ = ~pi1150 & ~new_n41482_;
  assign new_n41484_ = ~new_n41480_ & new_n41483_;
  assign new_n41485_ = ~new_n40269_ & ~new_n41472_;
  assign new_n41486_ = ~new_n40281_ & new_n40512_;
  assign new_n41487_ = ~pi0212 & ~new_n39638_;
  assign new_n41488_ = ~pi0219 & ~new_n41487_;
  assign new_n41489_ = ~new_n40524_ & new_n41488_;
  assign new_n41490_ = ~new_n41486_ & new_n41489_;
  assign new_n41491_ = ~new_n41485_ & ~new_n41490_;
  assign new_n41492_ = new_n41225_ & ~new_n41491_;
  assign new_n41493_ = pi0214 & ~new_n40142_;
  assign new_n41494_ = ~new_n40274_ & new_n41493_;
  assign new_n41495_ = ~pi0214 & new_n39675_;
  assign new_n41496_ = pi0212 & ~new_n41495_;
  assign new_n41497_ = ~new_n41494_ & new_n41496_;
  assign new_n41498_ = new_n40151_ & ~new_n41497_;
  assign new_n41499_ = ~new_n41485_ & ~new_n41498_;
  assign new_n41500_ = new_n41244_ & ~new_n41499_;
  assign new_n41501_ = pi1150 & ~new_n41500_;
  assign new_n41502_ = ~new_n41492_ & new_n41501_;
  assign new_n41503_ = ~new_n41484_ & ~new_n41502_;
  assign new_n41504_ = pi1148 & ~new_n41503_;
  assign new_n41505_ = ~pi0219 & ~new_n40212_;
  assign new_n41506_ = ~new_n40644_ & ~new_n41505_;
  assign new_n41507_ = new_n41472_ & new_n41506_;
  assign new_n41508_ = new_n41242_ & ~new_n41507_;
  assign new_n41509_ = ~new_n41265_ & ~new_n41472_;
  assign new_n41510_ = ~new_n41508_ & ~new_n41509_;
  assign new_n41511_ = pi1150 & new_n40163_;
  assign new_n41512_ = ~new_n41510_ & ~new_n41511_;
  assign new_n41513_ = pi1150 & new_n39682_;
  assign new_n41514_ = pi0299 & new_n40093_;
  assign new_n41515_ = ~pi0219 & ~new_n41514_;
  assign new_n41516_ = ~new_n41378_ & new_n41515_;
  assign new_n41517_ = ~new_n41513_ & new_n41516_;
  assign new_n41518_ = ~new_n41265_ & new_n41517_;
  assign new_n41519_ = ~pi1148 & ~new_n41518_;
  assign new_n41520_ = ~new_n41512_ & new_n41519_;
  assign new_n41521_ = ~new_n41504_ & ~new_n41520_;
  assign new_n41522_ = ~pi1149 & ~new_n41521_;
  assign new_n41523_ = new_n40212_ & new_n40313_;
  assign new_n41524_ = ~new_n40100_ & ~new_n41523_;
  assign new_n41525_ = new_n40121_ & new_n41524_;
  assign new_n41526_ = ~pi1146 & new_n40122_;
  assign new_n41527_ = new_n40084_ & ~new_n40105_;
  assign new_n41528_ = ~new_n40123_ & ~new_n41527_;
  assign new_n41529_ = ~new_n41526_ & ~new_n41528_;
  assign new_n41530_ = ~new_n41525_ & new_n41529_;
  assign new_n41531_ = ~new_n41265_ & ~new_n41530_;
  assign new_n41532_ = ~new_n40102_ & ~new_n40523_;
  assign new_n41533_ = ~pi0219 & ~new_n41532_;
  assign new_n41534_ = ~new_n41528_ & ~new_n41533_;
  assign new_n41535_ = ~pi1146 & ~new_n40100_;
  assign new_n41536_ = new_n41534_ & ~new_n41535_;
  assign new_n41537_ = new_n41242_ & ~new_n41536_;
  assign new_n41538_ = ~pi1150 & ~new_n41537_;
  assign new_n41539_ = ~new_n41531_ & new_n41538_;
  assign new_n41540_ = ~pi0214 & new_n40700_;
  assign new_n41541_ = new_n40074_ & ~new_n41540_;
  assign new_n41542_ = ~pi0219 & ~new_n41541_;
  assign new_n41543_ = ~new_n40062_ & ~new_n40700_;
  assign new_n41544_ = ~pi0212 & new_n41543_;
  assign new_n41545_ = new_n41542_ & ~new_n41544_;
  assign new_n41546_ = ~pi0299 & new_n39713_;
  assign new_n41547_ = ~new_n40064_ & ~new_n40237_;
  assign new_n41548_ = ~new_n41546_ & new_n41547_;
  assign new_n41549_ = new_n41545_ & new_n41548_;
  assign new_n41550_ = ~new_n40295_ & ~new_n41472_;
  assign new_n41551_ = new_n41542_ & ~new_n41543_;
  assign new_n41552_ = ~new_n41550_ & ~new_n41551_;
  assign new_n41553_ = ~new_n41549_ & new_n41552_;
  assign new_n41554_ = ~new_n40060_ & ~new_n41553_;
  assign new_n41555_ = new_n40063_ & ~new_n40073_;
  assign new_n41556_ = ~pi0219 & ~new_n41555_;
  assign new_n41557_ = ~new_n40704_ & new_n41556_;
  assign new_n41558_ = new_n40294_ & ~new_n41557_;
  assign new_n41559_ = ~new_n41554_ & new_n41558_;
  assign new_n41560_ = new_n41242_ & ~new_n41559_;
  assign new_n41561_ = ~new_n41265_ & ~new_n41553_;
  assign new_n41562_ = pi1150 & ~new_n41561_;
  assign new_n41563_ = ~new_n41560_ & new_n41562_;
  assign new_n41564_ = ~pi1148 & ~new_n41563_;
  assign new_n41565_ = ~new_n41539_ & new_n41564_;
  assign new_n41566_ = ~new_n40131_ & ~new_n41472_;
  assign new_n41567_ = ~new_n40172_ & new_n40190_;
  assign new_n41568_ = ~new_n40177_ & ~new_n41567_;
  assign new_n41569_ = ~new_n41244_ & ~new_n41568_;
  assign new_n41570_ = new_n39757_ & new_n41245_;
  assign new_n41571_ = new_n40189_ & ~new_n41570_;
  assign new_n41572_ = new_n40192_ & ~new_n41571_;
  assign new_n41573_ = ~new_n41569_ & new_n41572_;
  assign new_n41574_ = ~new_n41566_ & ~new_n41573_;
  assign new_n41575_ = ~new_n41470_ & ~new_n41574_;
  assign new_n41576_ = ~pi1150 & ~new_n41575_;
  assign new_n41577_ = ~new_n40319_ & ~new_n41507_;
  assign new_n41578_ = new_n41244_ & new_n41577_;
  assign new_n41579_ = pi0214 & new_n40312_;
  assign new_n41580_ = new_n40309_ & ~new_n41579_;
  assign new_n41581_ = ~pi0219 & ~new_n40315_;
  assign new_n41582_ = ~new_n41580_ & new_n41581_;
  assign new_n41583_ = new_n40307_ & ~new_n41582_;
  assign new_n41584_ = pi1146 & new_n40085_;
  assign new_n41585_ = new_n41225_ & ~new_n41584_;
  assign new_n41586_ = ~new_n41583_ & new_n41585_;
  assign new_n41587_ = pi1150 & ~new_n41586_;
  assign new_n41588_ = ~new_n41578_ & new_n41587_;
  assign new_n41589_ = pi1148 & ~new_n41588_;
  assign new_n41590_ = ~new_n41576_ & new_n41589_;
  assign new_n41591_ = pi1149 & ~new_n41590_;
  assign new_n41592_ = ~new_n41565_ & new_n41591_;
  assign new_n41593_ = ~new_n41522_ & ~new_n41592_;
  assign new_n41594_ = ~pi0213 & ~new_n41593_;
  assign new_n41595_ = pi1150 & new_n40089_;
  assign new_n41596_ = ~pi1150 & new_n40134_;
  assign new_n41597_ = pi1149 & ~new_n41596_;
  assign new_n41598_ = ~new_n41595_ & new_n41597_;
  assign new_n41599_ = pi1150 & new_n40161_;
  assign new_n41600_ = ~pi1150 & new_n40200_;
  assign new_n41601_ = ~pi1149 & ~new_n41600_;
  assign new_n41602_ = ~new_n41599_ & new_n41601_;
  assign new_n41603_ = ~new_n41598_ & ~new_n41602_;
  assign new_n41604_ = pi1148 & ~new_n41603_;
  assign new_n41605_ = ~pi1150 & new_n40125_;
  assign new_n41606_ = pi1150 & new_n40078_;
  assign new_n41607_ = pi1149 & ~new_n41606_;
  assign new_n41608_ = ~new_n41605_ & new_n41607_;
  assign new_n41609_ = ~pi1149 & pi1150;
  assign new_n41610_ = ~new_n40166_ & new_n41609_;
  assign new_n41611_ = ~new_n41608_ & ~new_n41610_;
  assign new_n41612_ = ~pi1148 & ~new_n41611_;
  assign new_n41613_ = ~new_n41604_ & ~new_n41612_;
  assign new_n41614_ = pi0213 & ~new_n41613_;
  assign new_n41615_ = pi0209 & ~new_n41614_;
  assign new_n41616_ = ~new_n41594_ & new_n41615_;
  assign new_n41617_ = ~pi0212 & ~new_n41404_;
  assign new_n41618_ = ~new_n13061_ & ~new_n41302_;
  assign new_n41619_ = pi0214 & ~new_n41618_;
  assign new_n41620_ = new_n41617_ & ~new_n41619_;
  assign new_n41621_ = ~pi0214 & ~new_n41618_;
  assign new_n41622_ = pi0214 & new_n41308_;
  assign new_n41623_ = pi0212 & ~new_n41622_;
  assign new_n41624_ = ~new_n41621_ & new_n41623_;
  assign new_n41625_ = ~new_n41620_ & ~new_n41624_;
  assign new_n41626_ = ~pi0219 & ~new_n41625_;
  assign new_n41627_ = new_n40343_ & ~new_n41392_;
  assign new_n41628_ = ~new_n41626_ & new_n41627_;
  assign new_n41629_ = pi0219 & ~new_n41358_;
  assign new_n41630_ = new_n41427_ & ~new_n41629_;
  assign new_n41631_ = ~new_n41376_ & new_n41630_;
  assign new_n41632_ = ~pi1150 & ~new_n40096_;
  assign new_n41633_ = ~new_n41631_ & new_n41632_;
  assign new_n41634_ = ~new_n41628_ & new_n41633_;
  assign new_n41635_ = ~new_n41406_ & new_n41617_;
  assign new_n41636_ = ~pi0214 & ~new_n41306_;
  assign new_n41637_ = new_n41623_ & ~new_n41636_;
  assign new_n41638_ = ~new_n41635_ & ~new_n41637_;
  assign new_n41639_ = ~pi0219 & ~new_n41638_;
  assign new_n41640_ = ~new_n41392_ & ~new_n41639_;
  assign new_n41641_ = ~pi1147 & ~new_n41640_;
  assign new_n41642_ = new_n41362_ & ~new_n41369_;
  assign new_n41643_ = ~pi0214 & ~new_n41368_;
  assign new_n41644_ = new_n41373_ & ~new_n41643_;
  assign new_n41645_ = ~new_n41642_ & ~new_n41644_;
  assign new_n41646_ = ~pi0219 & ~new_n41645_;
  assign new_n41647_ = ~new_n41629_ & ~new_n41646_;
  assign new_n41648_ = pi1147 & ~new_n41647_;
  assign new_n41649_ = ~po1038 & ~new_n41648_;
  assign new_n41650_ = ~new_n41641_ & new_n41649_;
  assign new_n41651_ = pi1150 & ~new_n39826_;
  assign new_n41652_ = ~new_n41650_ & new_n41651_;
  assign new_n41653_ = ~new_n41634_ & ~new_n41652_;
  assign new_n41654_ = pi1149 & ~new_n41653_;
  assign new_n41655_ = pi1150 & new_n40232_;
  assign new_n41656_ = ~pi1147 & new_n41305_;
  assign new_n41657_ = new_n16479_ & ~new_n41656_;
  assign new_n41658_ = new_n41655_ & ~new_n41657_;
  assign new_n41659_ = pi1147 & ~new_n41358_;
  assign new_n41660_ = new_n41302_ & ~new_n41655_;
  assign new_n41661_ = ~pi1147 & ~new_n41660_;
  assign new_n41662_ = ~po1038 & ~new_n41661_;
  assign new_n41663_ = ~new_n41659_ & new_n41662_;
  assign new_n41664_ = ~pi1149 & ~new_n41663_;
  assign new_n41665_ = ~new_n41658_ & new_n41664_;
  assign new_n41666_ = ~new_n41654_ & ~new_n41665_;
  assign new_n41667_ = ~pi1148 & ~new_n41666_;
  assign new_n41668_ = new_n41318_ & ~new_n41446_;
  assign new_n41669_ = new_n40343_ & ~new_n41668_;
  assign new_n41670_ = ~new_n41298_ & new_n41618_;
  assign new_n41671_ = pi0214 & new_n41670_;
  assign new_n41672_ = new_n41314_ & ~new_n41671_;
  assign new_n41673_ = new_n41311_ & ~new_n41672_;
  assign new_n41674_ = new_n41669_ & ~new_n41673_;
  assign new_n41675_ = ~new_n38413_ & new_n41370_;
  assign new_n41676_ = new_n41349_ & ~new_n41675_;
  assign new_n41677_ = new_n41427_ & ~new_n41676_;
  assign new_n41678_ = pi0214 & ~new_n13061_;
  assign new_n41679_ = new_n41339_ & new_n41678_;
  assign new_n41680_ = pi0212 & ~new_n41679_;
  assign new_n41681_ = ~pi0214 & new_n41371_;
  assign new_n41682_ = new_n41680_ & ~new_n41681_;
  assign new_n41683_ = new_n41330_ & ~new_n41371_;
  assign new_n41684_ = ~pi0219 & ~new_n41683_;
  assign new_n41685_ = ~new_n41682_ & new_n41684_;
  assign new_n41686_ = new_n41677_ & ~new_n41685_;
  assign new_n41687_ = pi1150 & ~new_n40141_;
  assign new_n41688_ = ~new_n41686_ & new_n41687_;
  assign new_n41689_ = ~new_n41674_ & new_n41688_;
  assign new_n41690_ = ~pi0219 & new_n41389_;
  assign new_n41691_ = new_n41669_ & ~new_n41690_;
  assign new_n41692_ = ~new_n41329_ & new_n41680_;
  assign new_n41693_ = ~pi0212 & new_n41328_;
  assign new_n41694_ = ~pi0219 & ~new_n41693_;
  assign new_n41695_ = ~new_n41692_ & new_n41694_;
  assign new_n41696_ = new_n41677_ & ~new_n41695_;
  assign new_n41697_ = ~pi1150 & ~new_n39830_;
  assign new_n41698_ = ~new_n41696_ & new_n41697_;
  assign new_n41699_ = ~new_n41691_ & new_n41698_;
  assign new_n41700_ = ~pi1149 & ~new_n41699_;
  assign new_n41701_ = ~new_n41689_ & new_n41700_;
  assign new_n41702_ = new_n41342_ & ~new_n41343_;
  assign new_n41703_ = ~new_n41676_ & ~new_n41702_;
  assign new_n41704_ = new_n6305_ & new_n41703_;
  assign new_n41705_ = ~new_n6305_ & ~new_n38795_;
  assign new_n41706_ = ~pi0057 & pi1147;
  assign new_n41707_ = ~new_n41705_ & new_n41706_;
  assign new_n41708_ = ~new_n41704_ & new_n41707_;
  assign new_n41709_ = pi0057 & new_n38795_;
  assign new_n41710_ = new_n6305_ & ~new_n38794_;
  assign new_n41711_ = new_n41317_ & new_n41710_;
  assign new_n41712_ = ~new_n38795_ & ~new_n41445_;
  assign new_n41713_ = ~pi0057 & ~pi1147;
  assign new_n41714_ = ~new_n41705_ & new_n41713_;
  assign new_n41715_ = ~new_n41712_ & new_n41714_;
  assign new_n41716_ = ~new_n41711_ & new_n41715_;
  assign new_n41717_ = ~new_n41709_ & ~new_n41716_;
  assign new_n41718_ = ~new_n41708_ & new_n41717_;
  assign new_n41719_ = pi1150 & ~new_n41718_;
  assign new_n41720_ = ~new_n41406_ & new_n41670_;
  assign new_n41721_ = pi0212 & ~new_n41720_;
  assign new_n41722_ = new_n41300_ & ~new_n41671_;
  assign new_n41723_ = ~pi0219 & ~new_n41722_;
  assign new_n41724_ = ~new_n41721_ & new_n41723_;
  assign new_n41725_ = new_n41669_ & ~new_n41724_;
  assign new_n41726_ = ~new_n40648_ & new_n41427_;
  assign new_n41727_ = new_n41703_ & new_n41726_;
  assign new_n41728_ = ~pi1150 & ~new_n40132_;
  assign new_n41729_ = ~new_n41727_ & new_n41728_;
  assign new_n41730_ = ~new_n41725_ & new_n41729_;
  assign new_n41731_ = pi1149 & ~new_n41730_;
  assign new_n41732_ = ~new_n41719_ & new_n41731_;
  assign new_n41733_ = pi1148 & ~new_n41732_;
  assign new_n41734_ = ~new_n41701_ & new_n41733_;
  assign new_n41735_ = pi0213 & ~new_n41734_;
  assign new_n41736_ = ~new_n41667_ & new_n41735_;
  assign new_n41737_ = ~pi0213 & ~new_n41402_;
  assign new_n41738_ = ~pi0209 & ~new_n41737_;
  assign new_n41739_ = ~new_n41736_ & new_n41738_;
  assign new_n41740_ = ~new_n41616_ & ~new_n41739_;
  assign new_n41741_ = pi0230 & ~new_n41740_;
  assign new_n41742_ = ~pi0230 & ~pi0246;
  assign po0403 = ~new_n41741_ & ~new_n41742_;
  assign new_n41744_ = ~pi1147 & ~new_n40744_;
  assign new_n41745_ = pi1151 & ~new_n40096_;
  assign new_n41746_ = ~new_n40061_ & ~new_n41545_;
  assign new_n41747_ = new_n41745_ & ~new_n41746_;
  assign new_n41748_ = new_n41744_ & ~new_n41747_;
  assign new_n41749_ = new_n40104_ & ~new_n40119_;
  assign new_n41750_ = ~new_n41528_ & ~new_n41749_;
  assign new_n41751_ = ~new_n40132_ & ~new_n41750_;
  assign new_n41752_ = ~pi1151 & new_n41751_;
  assign new_n41753_ = pi1151 & ~new_n40132_;
  assign new_n41754_ = new_n40294_ & ~new_n41551_;
  assign new_n41755_ = new_n41753_ & ~new_n41754_;
  assign new_n41756_ = pi1147 & ~new_n41755_;
  assign new_n41757_ = ~new_n41752_ & new_n41756_;
  assign new_n41758_ = ~pi1149 & ~new_n41757_;
  assign new_n41759_ = ~new_n41748_ & new_n41758_;
  assign new_n41760_ = ~pi1151 & ~new_n39826_;
  assign new_n41761_ = new_n40192_ & ~new_n41567_;
  assign new_n41762_ = new_n40652_ & ~new_n41761_;
  assign new_n41763_ = ~new_n40178_ & new_n40652_;
  assign new_n41764_ = ~new_n41762_ & ~new_n41763_;
  assign new_n41765_ = new_n41760_ & new_n41764_;
  assign new_n41766_ = new_n40499_ & ~new_n41583_;
  assign new_n41767_ = ~pi1147 & ~new_n41766_;
  assign new_n41768_ = ~new_n41765_ & new_n41767_;
  assign new_n41769_ = pi1147 & ~new_n40757_;
  assign new_n41770_ = ~new_n40082_ & ~new_n40085_;
  assign new_n41771_ = new_n40667_ & new_n41770_;
  assign new_n41772_ = new_n41769_ & ~new_n41771_;
  assign new_n41773_ = pi1149 & ~new_n41772_;
  assign new_n41774_ = ~new_n41768_ & new_n41773_;
  assign new_n41775_ = pi1150 & ~new_n41774_;
  assign new_n41776_ = ~new_n41759_ & new_n41775_;
  assign new_n41777_ = pi0212 & ~new_n39662_;
  assign new_n41778_ = new_n41489_ & ~new_n41777_;
  assign new_n41779_ = new_n40159_ & ~new_n41778_;
  assign new_n41780_ = new_n40580_ & ~new_n41779_;
  assign new_n41781_ = pi1147 & ~new_n41780_;
  assign new_n41782_ = new_n38423_ & ~new_n40173_;
  assign new_n41783_ = ~new_n40183_ & new_n40633_;
  assign new_n41784_ = ~new_n41782_ & new_n41783_;
  assign new_n41785_ = ~pi1151 & ~new_n40082_;
  assign new_n41786_ = ~new_n41784_ & new_n41785_;
  assign new_n41787_ = ~new_n40198_ & new_n41786_;
  assign new_n41788_ = new_n41781_ & ~new_n41787_;
  assign new_n41789_ = ~new_n40513_ & new_n41489_;
  assign new_n41790_ = new_n40269_ & ~new_n41789_;
  assign new_n41791_ = ~new_n39826_ & ~new_n41790_;
  assign new_n41792_ = pi1151 & new_n41791_;
  assign new_n41793_ = new_n41760_ & ~new_n41784_;
  assign new_n41794_ = ~pi1147 & ~new_n41793_;
  assign new_n41795_ = ~new_n41792_ & new_n41794_;
  assign new_n41796_ = pi1149 & ~new_n41795_;
  assign new_n41797_ = ~new_n41788_ & new_n41796_;
  assign new_n41798_ = ~new_n40727_ & new_n41753_;
  assign new_n41799_ = ~new_n40130_ & new_n40586_;
  assign new_n41800_ = pi1147 & ~new_n41799_;
  assign new_n41801_ = ~new_n41798_ & new_n41800_;
  assign new_n41802_ = ~new_n40095_ & new_n40164_;
  assign new_n41803_ = ~pi1151 & ~new_n41802_;
  assign new_n41804_ = ~pi1147 & ~new_n41803_;
  assign new_n41805_ = new_n39921_ & ~new_n40532_;
  assign new_n41806_ = new_n41745_ & ~new_n41805_;
  assign new_n41807_ = new_n41804_ & ~new_n41806_;
  assign new_n41808_ = ~pi1149 & ~new_n41807_;
  assign new_n41809_ = ~new_n41801_ & new_n41808_;
  assign new_n41810_ = ~pi1150 & ~new_n41809_;
  assign new_n41811_ = ~new_n41797_ & new_n41810_;
  assign new_n41812_ = ~new_n41776_ & ~new_n41811_;
  assign new_n41813_ = pi1148 & ~new_n41812_;
  assign new_n41814_ = pi1147 & ~new_n40752_;
  assign new_n41815_ = ~pi1151 & ~new_n40141_;
  assign new_n41816_ = ~new_n40198_ & new_n41815_;
  assign new_n41817_ = new_n41814_ & ~new_n41816_;
  assign new_n41818_ = ~new_n40154_ & new_n40269_;
  assign new_n41819_ = ~new_n40233_ & ~new_n41818_;
  assign new_n41820_ = pi1151 & new_n41819_;
  assign new_n41821_ = ~pi1151 & ~new_n40233_;
  assign new_n41822_ = ~new_n40617_ & new_n41821_;
  assign new_n41823_ = ~pi1147 & ~new_n41822_;
  assign new_n41824_ = ~new_n41820_ & new_n41823_;
  assign new_n41825_ = ~pi1150 & ~new_n41824_;
  assign new_n41826_ = ~new_n41817_ & new_n41825_;
  assign new_n41827_ = ~new_n41762_ & new_n41821_;
  assign new_n41828_ = pi1151 & ~new_n40233_;
  assign new_n41829_ = ~new_n40319_ & new_n41828_;
  assign new_n41830_ = ~pi1147 & ~new_n41829_;
  assign new_n41831_ = ~new_n41827_ & new_n41830_;
  assign new_n41832_ = new_n40554_ & new_n40646_;
  assign new_n41833_ = pi1147 & ~new_n41832_;
  assign new_n41834_ = ~new_n40141_ & ~new_n40197_;
  assign new_n41835_ = ~pi1151 & new_n41834_;
  assign new_n41836_ = new_n41833_ & ~new_n41835_;
  assign new_n41837_ = pi1150 & ~new_n41836_;
  assign new_n41838_ = ~new_n41831_ & new_n41837_;
  assign new_n41839_ = ~new_n41826_ & ~new_n41838_;
  assign new_n41840_ = pi1149 & ~new_n41839_;
  assign new_n41841_ = ~new_n41557_ & new_n41754_;
  assign new_n41842_ = new_n39831_ & ~new_n41841_;
  assign new_n41843_ = ~new_n39830_ & ~new_n41534_;
  assign new_n41844_ = ~pi1151 & new_n41843_;
  assign new_n41845_ = pi1147 & ~new_n41844_;
  assign new_n41846_ = ~new_n41842_ & new_n41845_;
  assign new_n41847_ = ~pi1151 & ~new_n40207_;
  assign new_n41848_ = ~pi1147 & ~new_n41847_;
  assign new_n41849_ = pi1151 & ~new_n40060_;
  assign new_n41850_ = new_n41848_ & ~new_n41849_;
  assign new_n41851_ = pi1150 & ~new_n41850_;
  assign new_n41852_ = ~new_n41846_ & new_n41851_;
  assign new_n41853_ = ~new_n39682_ & new_n40644_;
  assign new_n41854_ = new_n40725_ & ~new_n41853_;
  assign new_n41855_ = new_n39831_ & ~new_n41854_;
  assign new_n41856_ = new_n40569_ & ~new_n40645_;
  assign new_n41857_ = pi1147 & ~new_n41856_;
  assign new_n41858_ = ~new_n41855_ & new_n41857_;
  assign new_n41859_ = ~pi1147 & pi1151;
  assign new_n41860_ = new_n40163_ & new_n41859_;
  assign new_n41861_ = ~pi1150 & ~new_n41860_;
  assign new_n41862_ = ~new_n41858_ & new_n41861_;
  assign new_n41863_ = ~new_n41852_ & ~new_n41862_;
  assign new_n41864_ = ~pi1149 & ~new_n41863_;
  assign new_n41865_ = ~pi1148 & ~new_n41864_;
  assign new_n41866_ = ~new_n41840_ & new_n41865_;
  assign new_n41867_ = ~new_n41813_ & ~new_n41866_;
  assign new_n41868_ = ~pi0213 & ~new_n41867_;
  assign new_n41869_ = pi0213 & new_n40762_;
  assign new_n41870_ = pi0209 & ~new_n41869_;
  assign new_n41871_ = ~new_n41868_ & new_n41870_;
  assign new_n41872_ = ~new_n41762_ & new_n41828_;
  assign new_n41873_ = pi1147 & ~new_n40667_;
  assign new_n41874_ = ~new_n41872_ & new_n41873_;
  assign new_n41875_ = ~po1038 & ~new_n40712_;
  assign new_n41876_ = ~new_n40715_ & new_n41875_;
  assign new_n41877_ = ~new_n40481_ & ~new_n41876_;
  assign new_n41878_ = new_n41848_ & new_n41877_;
  assign new_n41879_ = ~pi1150 & ~new_n41878_;
  assign new_n41880_ = ~new_n41874_ & new_n41879_;
  assign new_n41881_ = new_n40116_ & new_n40123_;
  assign new_n41882_ = new_n40499_ & ~new_n41881_;
  assign new_n41883_ = new_n41744_ & ~new_n41882_;
  assign new_n41884_ = new_n40499_ & new_n41764_;
  assign new_n41885_ = new_n40522_ & ~new_n41763_;
  assign new_n41886_ = pi1147 & ~new_n41885_;
  assign new_n41887_ = ~new_n41884_ & new_n41886_;
  assign new_n41888_ = pi1150 & ~new_n41887_;
  assign new_n41889_ = ~new_n41883_ & new_n41888_;
  assign new_n41890_ = ~new_n41880_ & ~new_n41889_;
  assign new_n41891_ = ~pi1149 & ~new_n41890_;
  assign new_n41892_ = new_n40569_ & ~new_n41841_;
  assign new_n41893_ = ~new_n40141_ & ~new_n41558_;
  assign new_n41894_ = pi1151 & new_n41893_;
  assign new_n41895_ = ~pi1147 & ~new_n41894_;
  assign new_n41896_ = ~new_n41892_ & new_n41895_;
  assign new_n41897_ = ~new_n40087_ & new_n41856_;
  assign new_n41898_ = new_n41833_ & ~new_n41897_;
  assign new_n41899_ = ~pi1150 & ~new_n41898_;
  assign new_n41900_ = ~new_n41896_ & new_n41899_;
  assign new_n41901_ = new_n40586_ & ~new_n41754_;
  assign new_n41902_ = new_n40069_ & ~new_n40297_;
  assign new_n41903_ = new_n40294_ & ~new_n41902_;
  assign new_n41904_ = new_n40580_ & ~new_n41903_;
  assign new_n41905_ = ~pi1147 & ~new_n41904_;
  assign new_n41906_ = ~new_n41901_ & new_n41905_;
  assign new_n41907_ = ~new_n40132_ & ~new_n40649_;
  assign new_n41908_ = ~pi1151 & new_n41907_;
  assign new_n41909_ = new_n41769_ & ~new_n41908_;
  assign new_n41910_ = pi1150 & ~new_n41909_;
  assign new_n41911_ = ~new_n41906_ & new_n41910_;
  assign new_n41912_ = ~new_n41900_ & ~new_n41911_;
  assign new_n41913_ = pi1149 & ~new_n41912_;
  assign new_n41914_ = pi1148 & ~new_n41913_;
  assign new_n41915_ = ~new_n41891_ & new_n41914_;
  assign new_n41916_ = ~pi0219 & ~new_n40530_;
  assign new_n41917_ = ~new_n40622_ & new_n41916_;
  assign new_n41918_ = new_n40159_ & ~new_n41917_;
  assign new_n41919_ = ~new_n40155_ & new_n41918_;
  assign new_n41920_ = new_n40569_ & ~new_n41919_;
  assign new_n41921_ = new_n41814_ & ~new_n41920_;
  assign new_n41922_ = new_n39699_ & new_n39921_;
  assign new_n41923_ = ~new_n10729_ & new_n41922_;
  assign new_n41924_ = ~new_n41854_ & ~new_n41923_;
  assign new_n41925_ = new_n40554_ & new_n41924_;
  assign new_n41926_ = new_n40569_ & ~new_n41854_;
  assign new_n41927_ = ~pi1147 & ~new_n41926_;
  assign new_n41928_ = ~new_n41925_ & new_n41927_;
  assign new_n41929_ = ~pi1150 & ~new_n41928_;
  assign new_n41930_ = ~new_n41921_ & new_n41929_;
  assign new_n41931_ = ~new_n40132_ & ~new_n41918_;
  assign new_n41932_ = ~pi1151 & new_n41931_;
  assign new_n41933_ = new_n41781_ & ~new_n41932_;
  assign new_n41934_ = new_n40586_ & ~new_n40727_;
  assign new_n41935_ = new_n40580_ & ~new_n41922_;
  assign new_n41936_ = ~new_n40727_ & new_n41935_;
  assign new_n41937_ = ~pi1147 & ~new_n41936_;
  assign new_n41938_ = ~new_n41934_ & new_n41937_;
  assign new_n41939_ = pi1150 & ~new_n41938_;
  assign new_n41940_ = ~new_n41933_ & new_n41939_;
  assign new_n41941_ = ~new_n41930_ & ~new_n41940_;
  assign new_n41942_ = pi1149 & ~new_n41941_;
  assign new_n41943_ = new_n40185_ & new_n40633_;
  assign new_n41944_ = ~new_n40096_ & ~new_n41943_;
  assign new_n41945_ = ~pi1151 & new_n41944_;
  assign new_n41946_ = new_n40499_ & ~new_n41784_;
  assign new_n41947_ = pi1147 & ~new_n41946_;
  assign new_n41948_ = ~new_n41945_ & new_n41947_;
  assign new_n41949_ = ~new_n16479_ & new_n39825_;
  assign new_n41950_ = pi1151 & ~new_n41949_;
  assign new_n41951_ = new_n41804_ & ~new_n41950_;
  assign new_n41952_ = pi1150 & ~new_n41951_;
  assign new_n41953_ = ~new_n41948_ & new_n41952_;
  assign new_n41954_ = ~new_n40233_ & ~new_n40617_;
  assign new_n41955_ = ~pi1151 & ~new_n41473_;
  assign new_n41956_ = pi1147 & ~new_n41955_;
  assign new_n41957_ = ~new_n41954_ & new_n41956_;
  assign new_n41958_ = new_n40165_ & new_n41859_;
  assign new_n41959_ = ~pi1150 & ~new_n41958_;
  assign new_n41960_ = ~new_n41957_ & new_n41959_;
  assign new_n41961_ = ~new_n41953_ & ~new_n41960_;
  assign new_n41962_ = ~pi1149 & ~new_n41961_;
  assign new_n41963_ = ~pi1148 & ~new_n41962_;
  assign new_n41964_ = ~new_n41942_ & new_n41963_;
  assign new_n41965_ = ~new_n41915_ & ~new_n41964_;
  assign new_n41966_ = pi0213 & ~new_n41965_;
  assign new_n41967_ = ~pi0213 & ~new_n40205_;
  assign new_n41968_ = ~pi0209 & ~new_n41967_;
  assign new_n41969_ = ~new_n41966_ & new_n41968_;
  assign new_n41970_ = ~new_n41871_ & ~new_n41969_;
  assign new_n41971_ = pi0230 & ~new_n41970_;
  assign new_n41972_ = ~pi0230 & ~pi0247;
  assign po0404 = ~new_n41971_ & ~new_n41972_;
  assign new_n41974_ = pi1152 & ~new_n40757_;
  assign new_n41975_ = ~new_n41779_ & new_n41785_;
  assign new_n41976_ = new_n41974_ & ~new_n41975_;
  assign new_n41977_ = pi1151 & ~new_n40131_;
  assign new_n41978_ = new_n41770_ & new_n41977_;
  assign new_n41979_ = ~pi1152 & ~new_n41978_;
  assign new_n41980_ = ~new_n41787_ & new_n41979_;
  assign new_n41981_ = pi1150 & ~new_n41980_;
  assign new_n41982_ = ~new_n41976_ & new_n41981_;
  assign new_n41983_ = pi1151 & new_n41751_;
  assign new_n41984_ = ~pi1152 & ~new_n41799_;
  assign new_n41985_ = ~new_n41983_ & new_n41984_;
  assign new_n41986_ = pi1152 & ~new_n41934_;
  assign new_n41987_ = ~new_n41755_ & new_n41986_;
  assign new_n41988_ = ~pi1150 & ~new_n41987_;
  assign new_n41989_ = ~new_n41985_ & new_n41988_;
  assign new_n41990_ = pi1148 & ~new_n41989_;
  assign new_n41991_ = ~new_n41982_ & new_n41990_;
  assign new_n41992_ = ~new_n40124_ & new_n41745_;
  assign new_n41993_ = ~pi1152 & ~new_n41992_;
  assign new_n41994_ = ~new_n41803_ & new_n41993_;
  assign new_n41995_ = new_n40522_ & ~new_n41805_;
  assign new_n41996_ = pi1152 & ~new_n41995_;
  assign new_n41997_ = ~new_n41747_ & new_n41996_;
  assign new_n41998_ = ~pi1150 & ~new_n41997_;
  assign new_n41999_ = ~new_n41994_ & new_n41998_;
  assign new_n42000_ = ~pi1152 & ~new_n41793_;
  assign new_n42001_ = ~new_n41884_ & new_n42000_;
  assign new_n42002_ = ~pi1151 & new_n41791_;
  assign new_n42003_ = pi1152 & ~new_n41766_;
  assign new_n42004_ = ~new_n42002_ & new_n42003_;
  assign new_n42005_ = pi1150 & ~new_n42004_;
  assign new_n42006_ = ~new_n42001_ & new_n42005_;
  assign new_n42007_ = ~pi1148 & ~new_n42006_;
  assign new_n42008_ = ~new_n41999_ & new_n42007_;
  assign new_n42009_ = ~new_n41991_ & ~new_n42008_;
  assign new_n42010_ = pi1149 & ~new_n42009_;
  assign new_n42011_ = ~new_n40160_ & new_n41815_;
  assign new_n42012_ = pi1152 & ~new_n42011_;
  assign new_n42013_ = ~new_n41832_ & new_n42012_;
  assign new_n42014_ = pi1151 & new_n41834_;
  assign new_n42015_ = ~pi1152 & ~new_n41816_;
  assign new_n42016_ = ~new_n42014_ & new_n42015_;
  assign new_n42017_ = ~new_n42013_ & ~new_n42016_;
  assign new_n42018_ = pi1150 & ~new_n42017_;
  assign new_n42019_ = ~new_n41842_ & ~new_n41926_;
  assign new_n42020_ = pi1152 & ~new_n42019_;
  assign new_n42021_ = pi1151 & new_n41843_;
  assign new_n42022_ = ~new_n41856_ & ~new_n42021_;
  assign new_n42023_ = ~pi1152 & ~new_n42022_;
  assign new_n42024_ = ~pi1150 & ~new_n42023_;
  assign new_n42025_ = ~new_n42020_ & new_n42024_;
  assign new_n42026_ = pi1148 & ~new_n42025_;
  assign new_n42027_ = ~new_n42018_ & new_n42026_;
  assign new_n42028_ = ~pi1151 & new_n41819_;
  assign new_n42029_ = pi1152 & ~new_n41829_;
  assign new_n42030_ = ~new_n42028_ & new_n42029_;
  assign new_n42031_ = ~pi1152 & ~new_n41822_;
  assign new_n42032_ = ~new_n41872_ & new_n42031_;
  assign new_n42033_ = pi1150 & ~new_n42032_;
  assign new_n42034_ = ~new_n42030_ & new_n42033_;
  assign new_n42035_ = ~pi1151 & ~new_n40163_;
  assign new_n42036_ = pi1152 & ~new_n41849_;
  assign new_n42037_ = ~new_n42035_ & new_n42036_;
  assign new_n42038_ = pi1151 & ~pi1152;
  assign new_n42039_ = new_n40207_ & new_n42038_;
  assign new_n42040_ = ~pi1150 & ~new_n42039_;
  assign new_n42041_ = ~new_n42037_ & new_n42040_;
  assign new_n42042_ = ~new_n42034_ & ~new_n42041_;
  assign new_n42043_ = ~pi1148 & ~new_n42042_;
  assign new_n42044_ = ~pi1149 & ~new_n42043_;
  assign new_n42045_ = ~new_n42027_ & new_n42044_;
  assign new_n42046_ = ~new_n42010_ & ~new_n42045_;
  assign new_n42047_ = ~pi0213 & ~new_n42046_;
  assign new_n42048_ = ~new_n40125_ & new_n42038_;
  assign new_n42049_ = ~pi1151 & ~new_n40165_;
  assign new_n42050_ = ~new_n40163_ & new_n42049_;
  assign new_n42051_ = pi1152 & ~new_n42050_;
  assign new_n42052_ = ~new_n40745_ & new_n42051_;
  assign new_n42053_ = ~pi1150 & ~new_n42052_;
  assign new_n42054_ = ~new_n42048_ & new_n42053_;
  assign new_n42055_ = new_n41974_ & ~new_n42011_;
  assign new_n42056_ = pi1151 & new_n40134_;
  assign new_n42057_ = ~pi1152 & ~new_n42056_;
  assign new_n42058_ = ~new_n40753_ & new_n42057_;
  assign new_n42059_ = pi1150 & ~new_n42058_;
  assign new_n42060_ = ~new_n42055_ & new_n42059_;
  assign new_n42061_ = ~new_n42054_ & ~new_n42060_;
  assign new_n42062_ = pi0213 & new_n42061_;
  assign new_n42063_ = pi0209 & ~new_n42062_;
  assign new_n42064_ = ~new_n42047_ & new_n42063_;
  assign new_n42065_ = pi1151 & new_n41931_;
  assign new_n42066_ = ~pi1152 & ~new_n41920_;
  assign new_n42067_ = ~new_n42065_ & new_n42066_;
  assign new_n42068_ = ~new_n41780_ & new_n42012_;
  assign new_n42069_ = pi1150 & ~new_n42068_;
  assign new_n42070_ = ~new_n42067_ & new_n42069_;
  assign new_n42071_ = pi1151 & new_n41944_;
  assign new_n42072_ = ~pi1152 & ~new_n41955_;
  assign new_n42073_ = ~new_n42071_ & new_n42072_;
  assign new_n42074_ = pi1152 & ~new_n41822_;
  assign new_n42075_ = ~new_n41946_ & new_n42074_;
  assign new_n42076_ = ~pi1150 & ~new_n42075_;
  assign new_n42077_ = ~new_n42073_ & new_n42076_;
  assign new_n42078_ = ~pi1149 & ~new_n42077_;
  assign new_n42079_ = ~new_n42070_ & new_n42078_;
  assign new_n42080_ = pi1152 & ~new_n41827_;
  assign new_n42081_ = ~new_n41884_ & new_n42080_;
  assign new_n42082_ = new_n41745_ & ~new_n41763_;
  assign new_n42083_ = new_n40668_ & ~new_n42082_;
  assign new_n42084_ = ~pi1150 & ~new_n42083_;
  assign new_n42085_ = ~new_n42081_ & new_n42084_;
  assign new_n42086_ = new_n40646_ & new_n41815_;
  assign new_n42087_ = new_n41974_ & ~new_n42086_;
  assign new_n42088_ = pi1151 & new_n41907_;
  assign new_n42089_ = ~pi1152 & ~new_n41897_;
  assign new_n42090_ = ~new_n42088_ & new_n42089_;
  assign new_n42091_ = pi1150 & ~new_n42090_;
  assign new_n42092_ = ~new_n42087_ & new_n42091_;
  assign new_n42093_ = pi1149 & ~new_n42092_;
  assign new_n42094_ = ~new_n42085_ & new_n42093_;
  assign new_n42095_ = pi1148 & ~new_n42094_;
  assign new_n42096_ = ~new_n42079_ & new_n42095_;
  assign new_n42097_ = ~new_n41847_ & new_n41993_;
  assign new_n42098_ = ~pi1151 & ~new_n41877_;
  assign new_n42099_ = pi1152 & ~new_n42098_;
  assign new_n42100_ = ~new_n41882_ & new_n42099_;
  assign new_n42101_ = ~pi1150 & ~new_n42100_;
  assign new_n42102_ = ~new_n42097_ & new_n42101_;
  assign new_n42103_ = ~pi1152 & ~new_n41755_;
  assign new_n42104_ = ~new_n41892_ & new_n42103_;
  assign new_n42105_ = ~pi1151 & new_n41893_;
  assign new_n42106_ = pi1152 & ~new_n41904_;
  assign new_n42107_ = ~new_n42105_ & new_n42106_;
  assign new_n42108_ = pi1150 & ~new_n42107_;
  assign new_n42109_ = ~new_n42104_ & new_n42108_;
  assign new_n42110_ = pi1149 & ~new_n42109_;
  assign new_n42111_ = ~new_n42102_ & new_n42110_;
  assign new_n42112_ = new_n41815_ & new_n41924_;
  assign new_n42113_ = pi1152 & ~new_n41936_;
  assign new_n42114_ = ~new_n42112_ & new_n42113_;
  assign new_n42115_ = ~pi1152 & ~new_n41926_;
  assign new_n42116_ = ~new_n41798_ & new_n42115_;
  assign new_n42117_ = pi1150 & ~new_n42116_;
  assign new_n42118_ = ~new_n42114_ & new_n42117_;
  assign new_n42119_ = pi1152 & ~new_n41950_;
  assign new_n42120_ = ~new_n42049_ & new_n42119_;
  assign new_n42121_ = new_n41802_ & new_n42038_;
  assign new_n42122_ = ~pi1150 & ~new_n42121_;
  assign new_n42123_ = ~new_n42120_ & new_n42122_;
  assign new_n42124_ = ~pi1149 & ~new_n42123_;
  assign new_n42125_ = ~new_n42118_ & new_n42124_;
  assign new_n42126_ = ~pi1148 & ~new_n42125_;
  assign new_n42127_ = ~new_n42111_ & new_n42126_;
  assign new_n42128_ = pi0213 & ~new_n42127_;
  assign new_n42129_ = ~new_n42096_ & new_n42128_;
  assign new_n42130_ = ~pi0213 & ~new_n41613_;
  assign new_n42131_ = ~pi0209 & ~new_n42130_;
  assign new_n42132_ = ~new_n42129_ & new_n42131_;
  assign new_n42133_ = ~new_n42064_ & ~new_n42132_;
  assign new_n42134_ = pi0230 & ~new_n42133_;
  assign new_n42135_ = ~pi0230 & ~pi0248;
  assign po0405 = ~new_n42134_ & ~new_n42135_;
  assign new_n42137_ = ~pi0213 & new_n42061_;
  assign new_n42138_ = pi0299 & new_n38829_;
  assign new_n42139_ = ~new_n40183_ & ~new_n42138_;
  assign new_n42140_ = ~new_n39761_ & new_n42139_;
  assign new_n42141_ = ~pi0212 & ~new_n42140_;
  assign new_n42142_ = ~pi0214 & new_n42139_;
  assign new_n42143_ = ~new_n39904_ & ~new_n40182_;
  assign new_n42144_ = pi0214 & ~new_n40615_;
  assign new_n42145_ = ~new_n42143_ & new_n42144_;
  assign new_n42146_ = pi0212 & ~new_n42145_;
  assign new_n42147_ = ~new_n42142_ & new_n42146_;
  assign new_n42148_ = ~new_n42141_ & ~new_n42147_;
  assign new_n42149_ = ~pi0219 & ~new_n42148_;
  assign new_n42150_ = new_n6305_ & ~new_n40632_;
  assign new_n42151_ = ~new_n42149_ & new_n42150_;
  assign new_n42152_ = ~new_n6305_ & new_n38889_;
  assign new_n42153_ = ~pi0057 & ~pi1151;
  assign new_n42154_ = ~new_n42152_ & new_n42153_;
  assign new_n42155_ = ~new_n42151_ & new_n42154_;
  assign new_n42156_ = pi0057 & ~new_n38889_;
  assign new_n42157_ = ~new_n40653_ & ~new_n42138_;
  assign new_n42158_ = pi0214 & ~new_n42157_;
  assign new_n42159_ = ~pi0212 & ~new_n39761_;
  assign new_n42160_ = ~new_n42158_ & new_n42159_;
  assign new_n42161_ = ~pi0214 & ~new_n42157_;
  assign new_n42162_ = ~new_n39738_ & new_n39941_;
  assign new_n42163_ = pi0212 & ~new_n42162_;
  assign new_n42164_ = ~new_n42161_ & new_n42163_;
  assign new_n42165_ = ~pi0219 & ~new_n42164_;
  assign new_n42166_ = ~new_n42160_ & new_n42165_;
  assign new_n42167_ = new_n6305_ & ~new_n39768_;
  assign new_n42168_ = ~new_n42166_ & new_n42167_;
  assign new_n42169_ = ~pi0057 & pi1151;
  assign new_n42170_ = ~new_n42152_ & new_n42169_;
  assign new_n42171_ = ~new_n42168_ & new_n42170_;
  assign new_n42172_ = ~new_n42156_ & ~new_n42171_;
  assign new_n42173_ = ~new_n42155_ & new_n42172_;
  assign new_n42174_ = ~pi1152 & ~new_n42173_;
  assign new_n42175_ = new_n40144_ & ~new_n40608_;
  assign new_n42176_ = ~new_n39662_ & ~new_n42138_;
  assign new_n42177_ = ~pi0214 & ~new_n42176_;
  assign new_n42178_ = pi0212 & ~new_n42177_;
  assign new_n42179_ = ~new_n42175_ & new_n42178_;
  assign new_n42180_ = new_n40524_ & ~new_n42138_;
  assign new_n42181_ = new_n41488_ & ~new_n42180_;
  assign new_n42182_ = ~new_n42179_ & new_n42181_;
  assign new_n42183_ = ~pi1151 & ~new_n42182_;
  assign new_n42184_ = new_n40159_ & new_n42183_;
  assign new_n42185_ = pi0299 & ~new_n38829_;
  assign new_n42186_ = ~new_n10729_ & new_n42185_;
  assign new_n42187_ = ~new_n38827_ & ~new_n42186_;
  assign new_n42188_ = new_n40083_ & ~new_n42187_;
  assign new_n42189_ = new_n40640_ & ~new_n42188_;
  assign new_n42190_ = ~new_n40195_ & ~new_n40307_;
  assign new_n42191_ = pi1151 & ~new_n42190_;
  assign new_n42192_ = ~new_n42189_ & new_n42191_;
  assign new_n42193_ = new_n38834_ & ~new_n42192_;
  assign new_n42194_ = ~new_n42184_ & new_n42193_;
  assign new_n42195_ = pi1150 & ~new_n42194_;
  assign new_n42196_ = ~new_n42174_ & new_n42195_;
  assign new_n42197_ = pi0211 & new_n40713_;
  assign new_n42198_ = ~new_n38677_ & new_n40110_;
  assign new_n42199_ = new_n38788_ & ~new_n42198_;
  assign new_n42200_ = ~new_n42197_ & new_n42199_;
  assign new_n42201_ = new_n10729_ & new_n40714_;
  assign new_n42202_ = new_n39066_ & ~new_n40100_;
  assign new_n42203_ = ~new_n42201_ & ~new_n42202_;
  assign new_n42204_ = ~new_n42200_ & new_n42203_;
  assign new_n42205_ = ~pi0219 & ~new_n42204_;
  assign new_n42206_ = pi1151 & new_n40123_;
  assign new_n42207_ = ~new_n42205_ & new_n42206_;
  assign new_n42208_ = ~new_n39738_ & ~new_n42186_;
  assign new_n42209_ = new_n38888_ & new_n39695_;
  assign new_n42210_ = ~new_n42208_ & new_n42209_;
  assign new_n42211_ = new_n38891_ & ~new_n42210_;
  assign new_n42212_ = ~new_n42207_ & new_n42211_;
  assign new_n42213_ = new_n40062_ & ~new_n42185_;
  assign new_n42214_ = pi0212 & ~new_n42213_;
  assign new_n42215_ = ~new_n40692_ & new_n42214_;
  assign new_n42216_ = ~pi0212 & new_n39736_;
  assign new_n42217_ = ~pi0219 & ~new_n42216_;
  assign new_n42218_ = ~new_n42180_ & new_n42217_;
  assign new_n42219_ = ~new_n42215_ & new_n42218_;
  assign new_n42220_ = new_n39672_ & ~new_n40293_;
  assign new_n42221_ = ~new_n42219_ & new_n42220_;
  assign new_n42222_ = ~pi1151 & new_n41854_;
  assign new_n42223_ = new_n38834_ & ~new_n42210_;
  assign new_n42224_ = ~new_n42222_ & new_n42223_;
  assign new_n42225_ = ~new_n42221_ & new_n42224_;
  assign new_n42226_ = ~pi1150 & ~new_n42225_;
  assign new_n42227_ = ~new_n42212_ & new_n42226_;
  assign new_n42228_ = ~new_n42196_ & ~new_n42227_;
  assign new_n42229_ = pi0213 & ~new_n42228_;
  assign new_n42230_ = ~pi0209 & ~new_n42229_;
  assign new_n42231_ = ~new_n42137_ & new_n42230_;
  assign new_n42232_ = ~new_n10484_ & ~new_n39063_;
  assign new_n42233_ = new_n38635_ & ~new_n39231_;
  assign new_n42234_ = ~pi0207 & new_n39230_;
  assign new_n42235_ = pi0207 & ~new_n38646_;
  assign new_n42236_ = ~new_n39061_ & new_n42235_;
  assign new_n42237_ = pi0208 & ~new_n42236_;
  assign new_n42238_ = ~new_n42234_ & new_n42237_;
  assign new_n42239_ = ~new_n42233_ & ~new_n42238_;
  assign new_n42240_ = pi0211 & ~new_n42239_;
  assign new_n42241_ = pi0214 & new_n42240_;
  assign new_n42242_ = ~new_n42232_ & ~new_n42241_;
  assign new_n42243_ = ~pi0212 & ~new_n42242_;
  assign new_n42244_ = ~pi0219 & ~new_n42243_;
  assign new_n42245_ = ~pi0211 & new_n42239_;
  assign new_n42246_ = ~new_n39099_ & ~new_n42245_;
  assign new_n42247_ = pi0214 & ~new_n42246_;
  assign new_n42248_ = ~pi0211 & ~new_n39063_;
  assign new_n42249_ = ~pi0214 & ~new_n42248_;
  assign new_n42250_ = ~new_n42240_ & new_n42249_;
  assign new_n42251_ = pi0212 & ~new_n42250_;
  assign new_n42252_ = ~new_n42247_ & new_n42251_;
  assign new_n42253_ = new_n42244_ & ~new_n42252_;
  assign new_n42254_ = new_n39065_ & ~new_n42253_;
  assign new_n42255_ = new_n41745_ & ~new_n42254_;
  assign new_n42256_ = ~new_n39063_ & new_n39073_;
  assign new_n42257_ = ~new_n42038_ & ~new_n42256_;
  assign new_n42258_ = ~new_n42255_ & ~new_n42257_;
  assign new_n42259_ = pi0214 & new_n38953_;
  assign new_n42260_ = new_n38976_ & ~new_n42259_;
  assign new_n42261_ = ~pi0219 & ~new_n42260_;
  assign new_n42262_ = pi0214 & ~new_n38968_;
  assign new_n42263_ = ~pi0214 & new_n38953_;
  assign new_n42264_ = pi0212 & ~new_n42263_;
  assign new_n42265_ = ~new_n42262_ & new_n42264_;
  assign new_n42266_ = new_n42261_ & ~new_n42265_;
  assign new_n42267_ = ~po1038 & ~new_n38971_;
  assign new_n42268_ = ~new_n42266_ & new_n42267_;
  assign new_n42269_ = new_n40499_ & ~new_n42268_;
  assign new_n42270_ = ~new_n38968_ & new_n39885_;
  assign new_n42271_ = ~new_n38966_ & ~new_n39885_;
  assign new_n42272_ = ~po1038 & ~new_n42271_;
  assign new_n42273_ = ~new_n42270_ & new_n42272_;
  assign new_n42274_ = new_n41821_ & ~new_n42273_;
  assign new_n42275_ = pi1152 & ~new_n42274_;
  assign new_n42276_ = ~new_n42269_ & new_n42275_;
  assign new_n42277_ = ~new_n42258_ & ~new_n42276_;
  assign new_n42278_ = ~pi1150 & ~new_n42277_;
  assign new_n42279_ = ~new_n38413_ & new_n42246_;
  assign new_n42280_ = pi0219 & ~new_n39098_;
  assign new_n42281_ = ~new_n42279_ & new_n42280_;
  assign new_n42282_ = ~po1038 & ~new_n42281_;
  assign new_n42283_ = pi0214 & new_n42239_;
  assign new_n42284_ = new_n42251_ & ~new_n42283_;
  assign new_n42285_ = new_n42244_ & ~new_n42284_;
  assign new_n42286_ = new_n42282_ & ~new_n42285_;
  assign new_n42287_ = new_n41753_ & ~new_n42286_;
  assign new_n42288_ = pi0212 & ~new_n42242_;
  assign new_n42289_ = ~pi0212 & ~new_n39063_;
  assign new_n42290_ = ~pi0219 & ~new_n42289_;
  assign new_n42291_ = ~new_n42288_ & new_n42290_;
  assign new_n42292_ = new_n42282_ & ~new_n42291_;
  assign new_n42293_ = new_n40569_ & ~new_n42292_;
  assign new_n42294_ = ~pi1152 & ~new_n42293_;
  assign new_n42295_ = ~new_n42287_ & new_n42294_;
  assign new_n42296_ = ~new_n38975_ & ~new_n42262_;
  assign new_n42297_ = ~pi0212 & ~new_n42296_;
  assign new_n42298_ = ~pi0214 & new_n38968_;
  assign new_n42299_ = ~pi0211 & new_n38966_;
  assign new_n42300_ = ~new_n39011_ & ~new_n42299_;
  assign new_n42301_ = pi0214 & ~new_n42300_;
  assign new_n42302_ = pi0212 & ~new_n42301_;
  assign new_n42303_ = ~new_n42298_ & new_n42302_;
  assign new_n42304_ = ~new_n42297_ & ~new_n42303_;
  assign new_n42305_ = ~pi0219 & ~new_n42304_;
  assign new_n42306_ = new_n38974_ & ~new_n42305_;
  assign new_n42307_ = new_n41815_ & ~new_n42306_;
  assign new_n42308_ = pi0212 & ~new_n38953_;
  assign new_n42309_ = new_n42261_ & ~new_n42308_;
  assign new_n42310_ = new_n38974_ & ~new_n42309_;
  assign new_n42311_ = new_n40580_ & ~new_n42310_;
  assign new_n42312_ = pi1152 & ~new_n42311_;
  assign new_n42313_ = ~new_n42307_ & new_n42312_;
  assign new_n42314_ = ~new_n42295_ & ~new_n42313_;
  assign new_n42315_ = pi1150 & ~new_n42314_;
  assign new_n42316_ = ~new_n42278_ & ~new_n42315_;
  assign new_n42317_ = ~pi0213 & ~new_n42316_;
  assign new_n42318_ = pi0213 & new_n39071_;
  assign new_n42319_ = pi0209 & ~new_n42318_;
  assign new_n42320_ = ~new_n42317_ & new_n42319_;
  assign new_n42321_ = ~new_n42231_ & ~new_n42320_;
  assign new_n42322_ = pi0230 & ~new_n42321_;
  assign new_n42323_ = ~pi0230 & ~pi0249;
  assign po0406 = ~new_n42322_ & ~new_n42323_;
  assign new_n42325_ = new_n3281_ & new_n11510_;
  assign new_n42326_ = ~new_n6259_ & ~new_n42325_;
  assign new_n42327_ = ~pi0075 & ~new_n42326_;
  assign new_n42328_ = new_n7333_ & new_n8966_;
  assign new_n42329_ = ~new_n42327_ & ~new_n42328_;
  assign new_n42330_ = ~pi0087 & ~pi0250;
  assign new_n42331_ = new_n8881_ & new_n42330_;
  assign po0407 = ~new_n42329_ & new_n42331_;
  assign new_n42333_ = pi0897 & new_n10817_;
  assign new_n42334_ = ~pi0476 & new_n11444_;
  assign new_n42335_ = ~new_n42333_ & ~new_n42334_;
  assign new_n42336_ = pi0200 & pi1039;
  assign new_n42337_ = ~pi0200 & pi1053;
  assign new_n42338_ = ~pi0199 & ~new_n42337_;
  assign new_n42339_ = ~new_n42336_ & new_n42338_;
  assign new_n42340_ = ~new_n42335_ & ~new_n42339_;
  assign new_n42341_ = pi0251 & new_n42335_;
  assign po0408 = new_n42340_ | new_n42341_;
  assign new_n42343_ = ~pi0979 & ~pi0984;
  assign new_n42344_ = pi1001 & new_n42343_;
  assign new_n42345_ = new_n6191_ & new_n42344_;
  assign new_n42346_ = ~new_n6194_ & new_n42345_;
  assign new_n42347_ = new_n6454_ & new_n42346_;
  assign new_n42348_ = ~pi0252 & ~new_n42347_;
  assign new_n42349_ = pi1092 & ~pi1093;
  assign new_n42350_ = ~new_n42348_ & new_n42349_;
  assign new_n42351_ = new_n6466_ & ~new_n42350_;
  assign new_n42352_ = new_n6465_ & new_n42350_;
  assign new_n42353_ = ~new_n42351_ & ~new_n42352_;
  assign new_n42354_ = ~new_n6215_ & new_n42353_;
  assign new_n42355_ = new_n6215_ & new_n11550_;
  assign new_n42356_ = ~new_n42354_ & ~new_n42355_;
  assign new_n42357_ = ~new_n6238_ & ~new_n42356_;
  assign new_n42358_ = ~new_n6221_ & new_n11550_;
  assign new_n42359_ = new_n6221_ & new_n42353_;
  assign new_n42360_ = ~new_n42358_ & ~new_n42359_;
  assign new_n42361_ = new_n6238_ & ~new_n42360_;
  assign new_n42362_ = ~pi0299 & ~new_n42361_;
  assign new_n42363_ = ~new_n42357_ & new_n42362_;
  assign new_n42364_ = ~new_n6212_ & ~new_n42356_;
  assign new_n42365_ = new_n6212_ & ~new_n42360_;
  assign new_n42366_ = pi0299 & ~new_n42365_;
  assign new_n42367_ = ~new_n42364_ & new_n42366_;
  assign new_n42368_ = new_n10983_ & ~new_n42367_;
  assign new_n42369_ = ~new_n42363_ & new_n42368_;
  assign new_n42370_ = ~new_n10983_ & new_n11550_;
  assign new_n42371_ = ~new_n8870_ & ~new_n42370_;
  assign new_n42372_ = ~new_n42369_ & new_n42371_;
  assign new_n42373_ = new_n10982_ & new_n42345_;
  assign new_n42374_ = new_n21153_ & new_n42373_;
  assign new_n42375_ = new_n6198_ & new_n42374_;
  assign new_n42376_ = ~new_n38387_ & new_n42375_;
  assign new_n42377_ = new_n6454_ & new_n42376_;
  assign new_n42378_ = ~pi0252 & ~new_n42377_;
  assign new_n42379_ = ~pi0057 & pi1092;
  assign new_n42380_ = ~new_n42378_ & new_n42379_;
  assign new_n42381_ = pi0057 & new_n11549_;
  assign new_n42382_ = new_n8870_ & ~new_n42381_;
  assign new_n42383_ = ~new_n42380_ & new_n42382_;
  assign po0409 = ~new_n42372_ & ~new_n42383_;
  assign new_n42385_ = ~new_n13061_ & ~new_n38508_;
  assign new_n42386_ = ~new_n38608_ & new_n42385_;
  assign new_n42387_ = ~po1038 & new_n42386_;
  assign new_n42388_ = pi0219 & new_n40080_;
  assign new_n42389_ = ~new_n42387_ & ~new_n42388_;
  assign new_n42390_ = pi1153 & ~new_n42389_;
  assign new_n42391_ = ~pi1151 & ~new_n42390_;
  assign new_n42392_ = new_n10730_ & new_n38590_;
  assign new_n42393_ = pi0211 & ~new_n38550_;
  assign new_n42394_ = ~new_n42392_ & ~new_n42393_;
  assign new_n42395_ = ~new_n38543_ & ~new_n38556_;
  assign new_n42396_ = new_n38519_ & ~new_n42395_;
  assign new_n42397_ = ~po1038 & ~new_n42396_;
  assign new_n42398_ = new_n42394_ & new_n42397_;
  assign new_n42399_ = ~new_n11446_ & new_n39347_;
  assign new_n42400_ = pi1151 & ~new_n42399_;
  assign new_n42401_ = ~new_n42398_ & new_n42400_;
  assign new_n42402_ = ~new_n42391_ & ~new_n42401_;
  assign new_n42403_ = ~pi1152 & ~new_n42402_;
  assign new_n42404_ = new_n38519_ & new_n39797_;
  assign new_n42405_ = ~pi1151 & ~new_n11447_;
  assign new_n42406_ = ~new_n38595_ & new_n42405_;
  assign new_n42407_ = ~new_n42404_ & new_n42406_;
  assign new_n42408_ = ~new_n38548_ & ~new_n39904_;
  assign new_n42409_ = pi1153 & ~new_n42408_;
  assign new_n42410_ = ~new_n11373_ & ~new_n38508_;
  assign new_n42411_ = pi1151 & new_n42410_;
  assign new_n42412_ = ~new_n42409_ & new_n42411_;
  assign new_n42413_ = ~po1038 & ~new_n42412_;
  assign new_n42414_ = ~new_n42407_ & new_n42413_;
  assign new_n42415_ = ~pi1151 & new_n10730_;
  assign new_n42416_ = ~new_n39346_ & ~new_n42415_;
  assign new_n42417_ = po1038 & new_n42416_;
  assign new_n42418_ = pi1152 & ~new_n42417_;
  assign new_n42419_ = ~new_n42414_ & new_n42418_;
  assign new_n42420_ = ~new_n42403_ & ~new_n42419_;
  assign new_n42421_ = pi0230 & ~new_n42420_;
  assign new_n42422_ = ~new_n40892_ & ~new_n40906_;
  assign new_n42423_ = ~pi0211 & new_n40886_;
  assign new_n42424_ = new_n42422_ & ~new_n42423_;
  assign new_n42425_ = ~new_n40885_ & new_n40926_;
  assign new_n42426_ = new_n42424_ & new_n42425_;
  assign new_n42427_ = pi1153 & ~new_n42426_;
  assign new_n42428_ = ~pi1153 & ~new_n41037_;
  assign new_n42429_ = pi0219 & ~new_n42428_;
  assign new_n42430_ = ~new_n42427_ & new_n42429_;
  assign new_n42431_ = new_n40887_ & new_n40937_;
  assign new_n42432_ = pi1153 & ~new_n42431_;
  assign new_n42433_ = ~pi1153 & ~new_n40959_;
  assign new_n42434_ = ~pi0219 & ~new_n42433_;
  assign new_n42435_ = ~new_n42432_ & new_n42434_;
  assign new_n42436_ = pi0253 & ~new_n42435_;
  assign new_n42437_ = ~new_n42430_ & new_n42436_;
  assign new_n42438_ = ~new_n40897_ & new_n41037_;
  assign new_n42439_ = ~pi0211 & new_n42438_;
  assign new_n42440_ = ~new_n40899_ & ~new_n42439_;
  assign new_n42441_ = pi1153 & ~new_n42440_;
  assign new_n42442_ = ~new_n41032_ & ~new_n42441_;
  assign new_n42443_ = pi0219 & new_n42442_;
  assign new_n42444_ = pi1153 & new_n40907_;
  assign new_n42445_ = ~pi1153 & new_n40957_;
  assign new_n42446_ = ~pi0219 & ~new_n42445_;
  assign new_n42447_ = ~new_n42444_ & new_n42446_;
  assign new_n42448_ = ~pi0253 & ~new_n42447_;
  assign new_n42449_ = ~new_n42443_ & new_n42448_;
  assign new_n42450_ = ~new_n42437_ & ~new_n42449_;
  assign new_n42451_ = ~po1038 & ~new_n42450_;
  assign new_n42452_ = ~pi0211 & ~new_n40868_;
  assign new_n42453_ = pi0211 & new_n40895_;
  assign new_n42454_ = pi0219 & ~new_n42453_;
  assign new_n42455_ = ~new_n42452_ & new_n42454_;
  assign new_n42456_ = pi0219 & pi1091;
  assign new_n42457_ = ~new_n38500_ & new_n42456_;
  assign new_n42458_ = ~pi0219 & ~new_n40877_;
  assign new_n42459_ = ~new_n42457_ & ~new_n42458_;
  assign new_n42460_ = ~new_n42455_ & new_n42459_;
  assign new_n42461_ = ~pi0253 & ~new_n42460_;
  assign new_n42462_ = ~pi0219 & ~new_n40879_;
  assign new_n42463_ = ~new_n40895_ & ~new_n42457_;
  assign new_n42464_ = ~new_n42462_ & new_n42463_;
  assign new_n42465_ = pi0253 & ~new_n42464_;
  assign new_n42466_ = po1038 & ~new_n42465_;
  assign new_n42467_ = ~new_n42461_ & new_n42466_;
  assign new_n42468_ = ~pi0211 & ~new_n40877_;
  assign new_n42469_ = new_n42462_ & ~new_n42468_;
  assign new_n42470_ = ~pi0219 & ~new_n42469_;
  assign new_n42471_ = po1038 & new_n42470_;
  assign new_n42472_ = ~new_n40868_ & new_n42471_;
  assign new_n42473_ = pi1151 & ~new_n42472_;
  assign new_n42474_ = ~new_n42467_ & new_n42473_;
  assign new_n42475_ = ~new_n42451_ & new_n42474_;
  assign new_n42476_ = ~new_n40906_ & ~new_n40914_;
  assign new_n42477_ = ~pi1153 & ~new_n42476_;
  assign new_n42478_ = ~new_n40898_ & new_n42424_;
  assign new_n42479_ = ~new_n42477_ & new_n42478_;
  assign new_n42480_ = ~pi0219 & ~new_n42479_;
  assign new_n42481_ = pi0219 & new_n40892_;
  assign new_n42482_ = ~new_n42480_ & ~new_n42481_;
  assign new_n42483_ = ~new_n42443_ & new_n42482_;
  assign new_n42484_ = ~pi0253 & ~new_n42483_;
  assign new_n42485_ = ~new_n40887_ & ~new_n42439_;
  assign new_n42486_ = new_n42462_ & ~new_n42485_;
  assign new_n42487_ = ~new_n40915_ & ~new_n42477_;
  assign new_n42488_ = new_n42486_ & ~new_n42487_;
  assign new_n42489_ = pi0219 & new_n40992_;
  assign new_n42490_ = ~new_n41004_ & new_n42427_;
  assign new_n42491_ = new_n42489_ & ~new_n42490_;
  assign new_n42492_ = ~new_n42488_ & ~new_n42491_;
  assign new_n42493_ = pi0253 & ~new_n42492_;
  assign new_n42494_ = ~po1038 & ~new_n42493_;
  assign new_n42495_ = ~new_n42484_ & new_n42494_;
  assign new_n42496_ = ~pi1151 & ~new_n42495_;
  assign new_n42497_ = ~new_n42475_ & ~new_n42496_;
  assign new_n42498_ = ~new_n42452_ & new_n42458_;
  assign new_n42499_ = new_n42462_ & ~new_n42498_;
  assign new_n42500_ = pi0219 & ~new_n40868_;
  assign new_n42501_ = po1038 & ~new_n42500_;
  assign new_n42502_ = ~new_n42499_ & new_n42501_;
  assign new_n42503_ = ~new_n40868_ & new_n42502_;
  assign new_n42504_ = ~new_n42467_ & ~new_n42503_;
  assign new_n42505_ = ~new_n42497_ & new_n42504_;
  assign new_n42506_ = pi1152 & ~new_n42505_;
  assign new_n42507_ = pi0219 & ~new_n42442_;
  assign new_n42508_ = ~new_n42447_ & new_n42486_;
  assign new_n42509_ = ~new_n42507_ & ~new_n42508_;
  assign new_n42510_ = ~new_n40897_ & ~new_n42509_;
  assign new_n42511_ = ~pi0253 & ~new_n42510_;
  assign new_n42512_ = pi1153 & ~new_n40937_;
  assign new_n42513_ = new_n42424_ & new_n42462_;
  assign new_n42514_ = ~new_n42512_ & new_n42513_;
  assign new_n42515_ = ~new_n40994_ & ~new_n42426_;
  assign new_n42516_ = pi1153 & new_n42515_;
  assign new_n42517_ = ~pi1153 & ~new_n41043_;
  assign new_n42518_ = pi0219 & ~new_n42517_;
  assign new_n42519_ = ~new_n42516_ & new_n42518_;
  assign new_n42520_ = ~new_n42514_ & ~new_n42519_;
  assign new_n42521_ = pi0253 & ~new_n42520_;
  assign new_n42522_ = ~po1038 & ~new_n42521_;
  assign new_n42523_ = ~new_n42511_ & new_n42522_;
  assign new_n42524_ = new_n42474_ & ~new_n42523_;
  assign new_n42525_ = ~new_n40884_ & new_n42507_;
  assign new_n42526_ = ~pi1153 & ~new_n40929_;
  assign new_n42527_ = ~new_n40897_ & ~new_n42526_;
  assign new_n42528_ = ~pi0219 & new_n40959_;
  assign new_n42529_ = new_n42527_ & new_n42528_;
  assign new_n42530_ = ~pi0253 & ~new_n42529_;
  assign new_n42531_ = ~new_n42525_ & new_n42530_;
  assign new_n42532_ = ~new_n41004_ & ~new_n42426_;
  assign new_n42533_ = ~pi1091 & ~new_n41032_;
  assign new_n42534_ = ~pi1153 & ~new_n42533_;
  assign new_n42535_ = ~pi0219 & new_n42476_;
  assign new_n42536_ = ~new_n42534_ & ~new_n42535_;
  assign new_n42537_ = new_n42532_ & new_n42536_;
  assign new_n42538_ = pi0253 & ~new_n42537_;
  assign new_n42539_ = ~po1038 & ~new_n42538_;
  assign new_n42540_ = ~new_n42531_ & new_n42539_;
  assign new_n42541_ = ~pi1151 & ~new_n42467_;
  assign new_n42542_ = ~new_n42540_ & new_n42541_;
  assign new_n42543_ = ~pi1152 & ~new_n42542_;
  assign new_n42544_ = ~new_n42524_ & new_n42543_;
  assign new_n42545_ = ~new_n42506_ & ~new_n42544_;
  assign new_n42546_ = new_n41153_ & ~new_n42545_;
  assign new_n42547_ = pi1091 & ~new_n42394_;
  assign new_n42548_ = ~pi1153 & ~new_n41062_;
  assign new_n42549_ = pi1153 & ~new_n41092_;
  assign new_n42550_ = new_n38519_ & ~new_n42549_;
  assign new_n42551_ = ~new_n42548_ & new_n42550_;
  assign new_n42552_ = ~new_n42547_ & ~new_n42551_;
  assign new_n42553_ = pi0253 & ~new_n42552_;
  assign new_n42554_ = ~new_n13064_ & ~new_n42409_;
  assign new_n42555_ = pi1091 & ~new_n42554_;
  assign new_n42556_ = ~pi0253 & ~new_n42555_;
  assign new_n42557_ = ~po1038 & ~new_n42556_;
  assign new_n42558_ = ~new_n42553_ & new_n42557_;
  assign new_n42559_ = ~pi0253 & ~pi1091;
  assign new_n42560_ = po1038 & ~new_n42559_;
  assign new_n42561_ = pi0211 & pi1091;
  assign new_n42562_ = pi1091 & ~pi1153;
  assign new_n42563_ = pi0219 & new_n42562_;
  assign new_n42564_ = ~new_n42561_ & ~new_n42563_;
  assign new_n42565_ = new_n42560_ & new_n42564_;
  assign new_n42566_ = pi1151 & ~new_n42565_;
  assign new_n42567_ = ~new_n42558_ & new_n42566_;
  assign new_n42568_ = ~new_n42457_ & new_n42560_;
  assign new_n42569_ = pi0219 & new_n42568_;
  assign new_n42570_ = pi1091 & pi1153;
  assign new_n42571_ = new_n42387_ & new_n42570_;
  assign new_n42572_ = pi0253 & ~pi1091;
  assign new_n42573_ = ~pi1151 & ~new_n42572_;
  assign new_n42574_ = ~new_n42571_ & new_n42573_;
  assign new_n42575_ = ~new_n42569_ & new_n42574_;
  assign new_n42576_ = ~new_n42567_ & ~new_n42575_;
  assign new_n42577_ = ~pi1152 & ~new_n42576_;
  assign new_n42578_ = ~pi1153 & ~new_n41098_;
  assign new_n42579_ = ~new_n38533_ & new_n41058_;
  assign new_n42580_ = pi1153 & ~new_n42579_;
  assign new_n42581_ = new_n38519_ & ~new_n42580_;
  assign new_n42582_ = ~new_n42578_ & new_n42581_;
  assign new_n42583_ = new_n11446_ & new_n41058_;
  assign new_n42584_ = ~new_n38595_ & new_n42583_;
  assign new_n42585_ = pi0253 & ~new_n42584_;
  assign new_n42586_ = ~new_n42582_ & new_n42585_;
  assign new_n42587_ = pi1091 & new_n38595_;
  assign new_n42588_ = pi0211 & ~new_n41112_;
  assign new_n42589_ = ~new_n42587_ & new_n42588_;
  assign new_n42590_ = pi1091 & new_n39797_;
  assign new_n42591_ = pi1091 & new_n38556_;
  assign new_n42592_ = new_n38958_ & new_n42591_;
  assign new_n42593_ = new_n38519_ & ~new_n42592_;
  assign new_n42594_ = ~new_n42590_ & new_n42593_;
  assign new_n42595_ = ~pi0253 & ~new_n42594_;
  assign new_n42596_ = ~new_n42589_ & new_n42595_;
  assign new_n42597_ = ~new_n42586_ & ~new_n42596_;
  assign new_n42598_ = ~new_n11446_ & ~new_n38519_;
  assign new_n42599_ = ~new_n42572_ & new_n42598_;
  assign new_n42600_ = ~new_n42587_ & new_n42599_;
  assign new_n42601_ = new_n39695_ & ~new_n42600_;
  assign new_n42602_ = ~new_n42597_ & new_n42601_;
  assign new_n42603_ = new_n42408_ & ~new_n42572_;
  assign new_n42604_ = ~new_n42562_ & ~new_n42603_;
  assign new_n42605_ = new_n42410_ & ~new_n42604_;
  assign new_n42606_ = ~po1038 & ~new_n42559_;
  assign new_n42607_ = ~new_n42605_ & new_n42606_;
  assign new_n42608_ = ~new_n42568_ & ~new_n42607_;
  assign new_n42609_ = pi1151 & ~new_n42608_;
  assign new_n42610_ = ~pi0211 & pi1091;
  assign new_n42611_ = ~pi0219 & new_n42610_;
  assign new_n42612_ = new_n42568_ & ~new_n42611_;
  assign new_n42613_ = pi1152 & ~new_n42612_;
  assign new_n42614_ = ~new_n42609_ & new_n42613_;
  assign new_n42615_ = ~new_n42602_ & new_n42614_;
  assign new_n42616_ = ~new_n41153_ & ~new_n42615_;
  assign new_n42617_ = ~new_n42577_ & new_n42616_;
  assign new_n42618_ = ~pi0230 & ~new_n42617_;
  assign new_n42619_ = ~new_n42546_ & new_n42618_;
  assign po0410 = ~new_n42421_ & ~new_n42619_;
  assign new_n42621_ = pi1154 & new_n38992_;
  assign new_n42622_ = ~new_n39022_ & ~new_n42621_;
  assign new_n42623_ = new_n11446_ & ~new_n42622_;
  assign new_n42624_ = pi0299 & new_n38519_;
  assign new_n42625_ = ~new_n11446_ & new_n38959_;
  assign new_n42626_ = ~new_n42624_ & ~new_n42625_;
  assign new_n42627_ = ~new_n38939_ & ~new_n42626_;
  assign new_n42628_ = ~new_n42623_ & ~new_n42627_;
  assign new_n42629_ = ~po1038 & ~new_n42628_;
  assign new_n42630_ = ~pi0219 & ~new_n38828_;
  assign new_n42631_ = ~new_n39150_ & ~new_n42630_;
  assign new_n42632_ = po1038 & new_n42631_;
  assign new_n42633_ = ~pi1152 & ~new_n42632_;
  assign new_n42634_ = ~new_n42629_ & new_n42633_;
  assign new_n42635_ = ~new_n38540_ & ~new_n38991_;
  assign new_n42636_ = new_n38488_ & ~new_n42635_;
  assign new_n42637_ = ~pi1154 & ~new_n39056_;
  assign new_n42638_ = ~new_n38941_ & ~new_n42637_;
  assign new_n42639_ = ~new_n42636_ & new_n42638_;
  assign new_n42640_ = pi0219 & ~new_n42639_;
  assign new_n42641_ = ~pi0200 & pi1154;
  assign new_n42642_ = new_n11383_ & ~new_n42641_;
  assign new_n42643_ = new_n38991_ & ~new_n39904_;
  assign new_n42644_ = ~new_n42642_ & ~new_n42643_;
  assign new_n42645_ = ~pi0219 & ~new_n42644_;
  assign new_n42646_ = ~po1038 & ~new_n42645_;
  assign new_n42647_ = ~new_n42640_ & new_n42646_;
  assign new_n42648_ = new_n11446_ & ~new_n38828_;
  assign new_n42649_ = new_n40051_ & ~new_n42648_;
  assign new_n42650_ = pi1152 & ~new_n42649_;
  assign new_n42651_ = ~new_n42647_ & new_n42650_;
  assign new_n42652_ = ~new_n42634_ & ~new_n42651_;
  assign new_n42653_ = pi0230 & ~new_n42652_;
  assign new_n42654_ = ~pi1153 & new_n42479_;
  assign new_n42655_ = ~new_n40959_ & ~new_n42654_;
  assign new_n42656_ = ~pi1154 & ~new_n42655_;
  assign new_n42657_ = pi1154 & ~new_n40891_;
  assign new_n42658_ = new_n42424_ & new_n42657_;
  assign new_n42659_ = ~new_n42432_ & new_n42658_;
  assign new_n42660_ = pi0254 & ~new_n42659_;
  assign new_n42661_ = ~new_n42656_ & new_n42660_;
  assign new_n42662_ = ~new_n40898_ & new_n41043_;
  assign new_n42663_ = pi1154 & new_n42662_;
  assign new_n42664_ = ~new_n40957_ & ~new_n42663_;
  assign new_n42665_ = pi0211 & new_n40886_;
  assign new_n42666_ = ~new_n40897_ & ~new_n42665_;
  assign new_n42667_ = ~pi1153 & ~new_n42666_;
  assign new_n42668_ = ~pi0254 & ~new_n42667_;
  assign new_n42669_ = ~new_n42664_ & new_n42668_;
  assign new_n42670_ = ~new_n42661_ & ~new_n42669_;
  assign new_n42671_ = ~pi0219 & ~new_n42670_;
  assign new_n42672_ = pi1154 & ~new_n42427_;
  assign new_n42673_ = ~new_n42515_ & new_n42672_;
  assign new_n42674_ = pi1153 & ~new_n41037_;
  assign new_n42675_ = ~pi1154 & ~new_n42517_;
  assign new_n42676_ = ~new_n42674_ & new_n42675_;
  assign new_n42677_ = pi0254 & ~new_n42676_;
  assign new_n42678_ = ~new_n42673_ & new_n42677_;
  assign new_n42679_ = ~pi1153 & ~new_n40946_;
  assign new_n42680_ = new_n41034_ & ~new_n42679_;
  assign new_n42681_ = ~pi1154 & ~new_n42680_;
  assign new_n42682_ = ~new_n40897_ & new_n41032_;
  assign new_n42683_ = new_n42681_ & ~new_n42682_;
  assign new_n42684_ = ~new_n42428_ & new_n42662_;
  assign new_n42685_ = new_n38498_ & ~new_n42684_;
  assign new_n42686_ = ~new_n40869_ & new_n42685_;
  assign new_n42687_ = pi1153 & new_n40899_;
  assign new_n42688_ = new_n38488_ & ~new_n41021_;
  assign new_n42689_ = ~new_n42687_ & new_n42688_;
  assign new_n42690_ = ~pi0254 & ~new_n42689_;
  assign new_n42691_ = ~new_n42686_ & new_n42690_;
  assign new_n42692_ = ~new_n42683_ & new_n42691_;
  assign new_n42693_ = ~new_n42678_ & ~new_n42692_;
  assign new_n42694_ = pi0219 & ~new_n42693_;
  assign new_n42695_ = pi0253 & ~new_n42694_;
  assign new_n42696_ = ~new_n42671_ & new_n42695_;
  assign new_n42697_ = ~pi0211 & new_n38589_;
  assign new_n42698_ = pi1153 & ~new_n41076_;
  assign new_n42699_ = ~pi1154 & ~new_n42698_;
  assign new_n42700_ = ~new_n42548_ & new_n42699_;
  assign new_n42701_ = ~new_n42697_ & new_n42700_;
  assign new_n42702_ = pi1091 & new_n38488_;
  assign new_n42703_ = ~new_n38548_ & new_n42702_;
  assign new_n42704_ = ~new_n39034_ & new_n42703_;
  assign new_n42705_ = ~new_n42701_ & ~new_n42704_;
  assign new_n42706_ = ~pi0219 & ~new_n42705_;
  assign new_n42707_ = pi1154 & new_n42610_;
  assign new_n42708_ = ~new_n42456_ & ~new_n42707_;
  assign new_n42709_ = ~new_n42639_ & ~new_n42708_;
  assign new_n42710_ = ~new_n42706_ & ~new_n42709_;
  assign new_n42711_ = pi0254 & ~new_n42710_;
  assign new_n42712_ = ~pi0254 & ~pi1091;
  assign new_n42713_ = pi1154 & ~new_n42408_;
  assign new_n42714_ = pi0219 & ~new_n39056_;
  assign new_n42715_ = ~new_n42713_ & new_n42714_;
  assign new_n42716_ = ~new_n42645_ & ~new_n42715_;
  assign new_n42717_ = ~pi0254 & ~new_n42716_;
  assign new_n42718_ = ~new_n42712_ & ~new_n42717_;
  assign new_n42719_ = ~new_n42711_ & new_n42718_;
  assign new_n42720_ = ~pi0253 & ~new_n42719_;
  assign new_n42721_ = ~po1038 & ~new_n42720_;
  assign new_n42722_ = ~new_n42696_ & new_n42721_;
  assign new_n42723_ = new_n42498_ & ~new_n42570_;
  assign new_n42724_ = pi1091 & new_n39150_;
  assign new_n42725_ = ~pi0254 & ~new_n42724_;
  assign new_n42726_ = ~new_n42455_ & new_n42725_;
  assign new_n42727_ = ~new_n42723_ & new_n42726_;
  assign new_n42728_ = ~pi0211 & ~new_n40893_;
  assign new_n42729_ = new_n42500_ & ~new_n42728_;
  assign new_n42730_ = ~pi0219 & new_n40877_;
  assign new_n42731_ = ~new_n42729_ & ~new_n42730_;
  assign new_n42732_ = new_n11446_ & new_n42562_;
  assign new_n42733_ = pi0254 & ~new_n42732_;
  assign new_n42734_ = ~new_n42724_ & new_n42733_;
  assign new_n42735_ = new_n42731_ & new_n42734_;
  assign new_n42736_ = pi0253 & ~new_n42735_;
  assign new_n42737_ = ~new_n42727_ & new_n42736_;
  assign new_n42738_ = pi1091 & ~new_n42631_;
  assign new_n42739_ = po1038 & ~new_n42712_;
  assign new_n42740_ = ~new_n42738_ & new_n42739_;
  assign new_n42741_ = po1038 & new_n42611_;
  assign new_n42742_ = ~new_n42740_ & ~new_n42741_;
  assign new_n42743_ = pi0253 & po1038;
  assign new_n42744_ = new_n42742_ & ~new_n42743_;
  assign new_n42745_ = ~new_n42737_ & ~new_n42744_;
  assign new_n42746_ = pi1152 & ~new_n42745_;
  assign new_n42747_ = ~new_n42722_ & new_n42746_;
  assign new_n42748_ = ~pi1154 & ~new_n41025_;
  assign new_n42749_ = ~pi1154 & ~new_n42748_;
  assign new_n42750_ = ~pi1153 & new_n40926_;
  assign new_n42751_ = ~new_n42425_ & ~new_n42750_;
  assign new_n42752_ = ~new_n42749_ & new_n42751_;
  assign new_n42753_ = new_n38498_ & ~new_n41004_;
  assign new_n42754_ = pi0219 & ~new_n42753_;
  assign new_n42755_ = ~new_n42752_ & new_n42754_;
  assign new_n42756_ = new_n42485_ & ~new_n42750_;
  assign new_n42757_ = pi1154 & new_n40914_;
  assign new_n42758_ = ~pi0219 & ~new_n42757_;
  assign new_n42759_ = ~new_n42756_ & new_n42758_;
  assign new_n42760_ = ~new_n42755_ & ~new_n42759_;
  assign new_n42761_ = pi0254 & ~new_n42760_;
  assign new_n42762_ = new_n40900_ & ~new_n42428_;
  assign new_n42763_ = new_n38488_ & ~new_n42762_;
  assign new_n42764_ = pi0219 & ~new_n42685_;
  assign new_n42765_ = ~new_n42681_ & new_n42764_;
  assign new_n42766_ = ~new_n42763_ & new_n42765_;
  assign new_n42767_ = ~new_n40891_ & new_n40957_;
  assign new_n42768_ = ~new_n42526_ & new_n42767_;
  assign new_n42769_ = ~new_n40897_ & new_n40959_;
  assign new_n42770_ = pi1154 & ~new_n42769_;
  assign new_n42771_ = ~new_n42768_ & new_n42770_;
  assign new_n42772_ = ~pi1154 & ~new_n42768_;
  assign new_n42773_ = pi1154 & new_n40892_;
  assign new_n42774_ = ~new_n40886_ & ~new_n42773_;
  assign new_n42775_ = ~pi0211 & ~new_n42774_;
  assign new_n42776_ = ~pi0219 & ~new_n42775_;
  assign new_n42777_ = ~new_n42772_ & new_n42776_;
  assign new_n42778_ = ~new_n42771_ & new_n42777_;
  assign new_n42779_ = ~pi0254 & ~new_n42778_;
  assign new_n42780_ = ~new_n42766_ & new_n42779_;
  assign new_n42781_ = ~new_n42761_ & ~new_n42780_;
  assign new_n42782_ = pi0253 & ~new_n42781_;
  assign new_n42783_ = new_n41065_ & new_n42562_;
  assign new_n42784_ = ~new_n42590_ & ~new_n42783_;
  assign new_n42785_ = pi0211 & ~new_n42699_;
  assign new_n42786_ = ~new_n42784_ & new_n42785_;
  assign new_n42787_ = pi1091 & new_n38959_;
  assign new_n42788_ = pi1154 & ~new_n42787_;
  assign new_n42789_ = new_n11445_ & new_n42570_;
  assign new_n42790_ = ~pi1154 & ~new_n42789_;
  assign new_n42791_ = ~pi0211 & ~new_n42790_;
  assign new_n42792_ = ~new_n42788_ & new_n42791_;
  assign new_n42793_ = ~new_n42786_ & ~new_n42792_;
  assign new_n42794_ = ~pi0219 & ~new_n42793_;
  assign new_n42795_ = pi0211 & new_n42788_;
  assign new_n42796_ = pi1091 & new_n39643_;
  assign new_n42797_ = new_n38498_ & ~new_n42796_;
  assign new_n42798_ = ~new_n42590_ & new_n42797_;
  assign new_n42799_ = pi0219 & ~new_n42790_;
  assign new_n42800_ = ~new_n42798_ & new_n42799_;
  assign new_n42801_ = ~new_n42795_ & new_n42800_;
  assign new_n42802_ = ~new_n42794_ & ~new_n42801_;
  assign new_n42803_ = ~pi0254 & ~new_n42802_;
  assign new_n42804_ = pi1091 & ~new_n11446_;
  assign new_n42805_ = ~new_n38938_ & new_n42804_;
  assign new_n42806_ = ~pi1154 & ~new_n42805_;
  assign new_n42807_ = ~pi1153 & ~new_n41066_;
  assign new_n42808_ = ~new_n42580_ & ~new_n42807_;
  assign new_n42809_ = pi1091 & ~new_n38534_;
  assign new_n42810_ = ~new_n42808_ & ~new_n42809_;
  assign new_n42811_ = new_n42598_ & ~new_n42810_;
  assign new_n42812_ = new_n41115_ & new_n42581_;
  assign new_n42813_ = pi1154 & ~new_n42812_;
  assign new_n42814_ = ~new_n42811_ & new_n42813_;
  assign new_n42815_ = ~new_n42806_ & ~new_n42814_;
  assign new_n42816_ = pi1091 & ~pi1154;
  assign new_n42817_ = new_n38638_ & new_n42816_;
  assign new_n42818_ = ~new_n42808_ & ~new_n42817_;
  assign new_n42819_ = new_n11446_ & ~new_n42818_;
  assign new_n42820_ = pi0254 & ~new_n42819_;
  assign new_n42821_ = ~new_n42815_ & new_n42820_;
  assign new_n42822_ = ~new_n42803_ & ~new_n42821_;
  assign new_n42823_ = ~pi0253 & new_n42822_;
  assign new_n42824_ = ~po1038 & ~new_n42823_;
  assign new_n42825_ = ~new_n42782_ & new_n42824_;
  assign new_n42826_ = ~new_n42740_ & ~new_n42743_;
  assign new_n42827_ = ~new_n42470_ & new_n42727_;
  assign new_n42828_ = ~new_n42499_ & new_n42735_;
  assign new_n42829_ = pi0253 & ~new_n42828_;
  assign new_n42830_ = ~new_n42827_ & new_n42829_;
  assign new_n42831_ = ~new_n42826_ & ~new_n42830_;
  assign new_n42832_ = ~pi1152 & ~new_n42831_;
  assign new_n42833_ = ~new_n42825_ & new_n42832_;
  assign new_n42834_ = new_n41153_ & ~new_n42833_;
  assign new_n42835_ = ~new_n42747_ & new_n42834_;
  assign new_n42836_ = ~po1038 & ~new_n42822_;
  assign new_n42837_ = ~pi1152 & ~new_n42740_;
  assign new_n42838_ = ~new_n42836_ & new_n42837_;
  assign new_n42839_ = ~po1038 & new_n42719_;
  assign new_n42840_ = pi1152 & new_n42742_;
  assign new_n42841_ = ~new_n42839_ & new_n42840_;
  assign new_n42842_ = ~new_n41153_ & ~new_n42841_;
  assign new_n42843_ = ~new_n42838_ & new_n42842_;
  assign new_n42844_ = ~pi0230 & ~new_n42843_;
  assign new_n42845_ = ~new_n42835_ & new_n42844_;
  assign po0411 = ~new_n42653_ & ~new_n42845_;
  assign new_n42847_ = ~pi0200 & pi1049;
  assign new_n42848_ = pi0200 & pi1036;
  assign new_n42849_ = ~new_n42847_ & ~new_n42848_;
  assign new_n42850_ = ~new_n42335_ & new_n42849_;
  assign new_n42851_ = ~pi0255 & new_n42335_;
  assign po0412 = ~new_n42850_ & ~new_n42851_;
  assign new_n42853_ = ~pi0200 & pi1048;
  assign new_n42854_ = pi0200 & pi1070;
  assign new_n42855_ = ~new_n42853_ & ~new_n42854_;
  assign new_n42856_ = ~new_n42335_ & new_n42855_;
  assign new_n42857_ = ~pi0256 & new_n42335_;
  assign po0413 = ~new_n42856_ & ~new_n42857_;
  assign new_n42859_ = ~pi0200 & pi1084;
  assign new_n42860_ = pi0200 & pi1065;
  assign new_n42861_ = ~new_n42859_ & ~new_n42860_;
  assign new_n42862_ = ~new_n42335_ & new_n42861_;
  assign new_n42863_ = ~pi0257 & new_n42335_;
  assign po0414 = ~new_n42862_ & ~new_n42863_;
  assign new_n42865_ = ~pi0200 & pi1072;
  assign new_n42866_ = pi0200 & pi1062;
  assign new_n42867_ = ~new_n42865_ & ~new_n42866_;
  assign new_n42868_ = ~new_n42335_ & new_n42867_;
  assign new_n42869_ = ~pi0258 & new_n42335_;
  assign po0415 = ~new_n42868_ & ~new_n42869_;
  assign new_n42871_ = ~pi0200 & pi1059;
  assign new_n42872_ = pi0200 & pi1069;
  assign new_n42873_ = ~new_n42871_ & ~new_n42872_;
  assign new_n42874_ = ~new_n42335_ & new_n42873_;
  assign new_n42875_ = ~pi0259 & new_n42335_;
  assign po0416 = ~new_n42874_ & ~new_n42875_;
  assign new_n42877_ = pi0200 & pi1067;
  assign new_n42878_ = ~pi0200 & pi1044;
  assign new_n42879_ = ~pi0199 & ~new_n42878_;
  assign new_n42880_ = ~new_n42877_ & new_n42879_;
  assign new_n42881_ = ~new_n42335_ & ~new_n42880_;
  assign new_n42882_ = pi0260 & new_n42335_;
  assign po0417 = new_n42881_ | new_n42882_;
  assign new_n42884_ = pi0200 & pi1040;
  assign new_n42885_ = ~pi0200 & pi1037;
  assign new_n42886_ = ~pi0199 & ~new_n42885_;
  assign new_n42887_ = ~new_n42884_ & new_n42886_;
  assign new_n42888_ = ~new_n42335_ & ~new_n42887_;
  assign new_n42889_ = pi0261 & new_n42335_;
  assign po0418 = new_n42888_ | new_n42889_;
  assign new_n42891_ = pi1093 & pi1142;
  assign new_n42892_ = ~pi0262 & ~pi1093;
  assign new_n42893_ = ~new_n42891_ & ~new_n42892_;
  assign new_n42894_ = ~pi0228 & ~new_n42893_;
  assign new_n42895_ = pi0123 & pi0262;
  assign new_n42896_ = ~pi0123 & ~pi1142;
  assign new_n42897_ = pi0228 & ~new_n42896_;
  assign new_n42898_ = ~new_n42895_ & new_n42897_;
  assign new_n42899_ = ~new_n42894_ & ~new_n42898_;
  assign new_n42900_ = ~pi0228 & ~pi1093;
  assign new_n42901_ = pi0123 & pi0228;
  assign new_n42902_ = ~new_n42900_ & ~new_n42901_;
  assign new_n42903_ = ~pi0262 & ~new_n42902_;
  assign new_n42904_ = ~new_n40731_ & ~new_n42903_;
  assign new_n42905_ = pi0199 & new_n42902_;
  assign new_n42906_ = new_n38442_ & ~new_n42905_;
  assign new_n42907_ = new_n42904_ & ~new_n42906_;
  assign new_n42908_ = ~new_n42899_ & ~new_n42907_;
  assign new_n42909_ = ~pi0207 & new_n42903_;
  assign new_n42910_ = ~pi0208 & ~new_n42909_;
  assign new_n42911_ = ~new_n40731_ & ~new_n42910_;
  assign new_n42912_ = ~new_n42908_ & ~new_n42911_;
  assign new_n42913_ = pi0299 & ~new_n42904_;
  assign new_n42914_ = ~new_n39711_ & new_n42902_;
  assign new_n42915_ = ~pi0299 & ~new_n42914_;
  assign new_n42916_ = ~new_n42899_ & new_n42915_;
  assign new_n42917_ = pi0208 & ~new_n42916_;
  assign new_n42918_ = ~new_n42913_ & new_n42917_;
  assign new_n42919_ = ~po1038 & ~new_n42918_;
  assign new_n42920_ = ~new_n42912_ & new_n42919_;
  assign new_n42921_ = ~new_n39825_ & new_n42902_;
  assign new_n42922_ = po1038 & ~new_n42899_;
  assign new_n42923_ = ~new_n42921_ & new_n42922_;
  assign po0419 = new_n42920_ | new_n42923_;
  assign new_n42925_ = pi1154 & ~new_n40908_;
  assign new_n42926_ = ~new_n40962_ & new_n42925_;
  assign new_n42927_ = ~pi1154 & ~new_n40930_;
  assign new_n42928_ = pi1155 & new_n42767_;
  assign new_n42929_ = new_n42927_ & ~new_n42928_;
  assign new_n42930_ = ~new_n40980_ & new_n42925_;
  assign new_n42931_ = ~pi1156 & ~new_n42757_;
  assign new_n42932_ = ~new_n42930_ & new_n42931_;
  assign new_n42933_ = ~pi1156 & ~new_n42932_;
  assign new_n42934_ = ~new_n42929_ & ~new_n42933_;
  assign new_n42935_ = pi1156 & new_n42769_;
  assign new_n42936_ = ~new_n42934_ & ~new_n42935_;
  assign new_n42937_ = ~new_n42926_ & ~new_n42936_;
  assign new_n42938_ = pi0211 & ~new_n42937_;
  assign new_n42939_ = new_n40910_ & ~new_n40956_;
  assign new_n42940_ = pi1155 & new_n42939_;
  assign new_n42941_ = new_n42927_ & ~new_n42940_;
  assign new_n42942_ = new_n42932_ & ~new_n42941_;
  assign new_n42943_ = ~new_n42769_ & new_n42941_;
  assign new_n42944_ = pi1156 & ~new_n42943_;
  assign new_n42945_ = ~new_n42930_ & new_n42944_;
  assign new_n42946_ = ~pi0211 & ~new_n42945_;
  assign new_n42947_ = ~new_n42942_ & new_n42946_;
  assign new_n42948_ = ~pi0219 & ~new_n42947_;
  assign new_n42949_ = ~new_n42938_ & new_n42948_;
  assign new_n42950_ = ~new_n40902_ & ~new_n41033_;
  assign new_n42951_ = ~new_n40900_ & ~new_n42773_;
  assign new_n42952_ = ~new_n42950_ & ~new_n42951_;
  assign new_n42953_ = ~new_n40956_ & new_n42952_;
  assign new_n42954_ = ~pi1156 & ~new_n42953_;
  assign new_n42955_ = new_n38479_ & ~new_n42952_;
  assign new_n42956_ = ~pi1155 & ~new_n42438_;
  assign new_n42957_ = pi1155 & ~new_n42662_;
  assign new_n42958_ = ~pi1154 & ~new_n42957_;
  assign new_n42959_ = ~new_n42956_ & new_n42958_;
  assign new_n42960_ = pi1154 & ~new_n42950_;
  assign new_n42961_ = new_n38483_ & ~new_n42960_;
  assign new_n42962_ = ~new_n42959_ & new_n42961_;
  assign new_n42963_ = pi0219 & ~new_n42962_;
  assign new_n42964_ = ~new_n42955_ & new_n42963_;
  assign new_n42965_ = ~new_n42954_ & new_n42964_;
  assign new_n42966_ = pi0263 & ~new_n42965_;
  assign new_n42967_ = ~new_n42949_ & new_n42966_;
  assign new_n42968_ = ~pi1155 & new_n42533_;
  assign new_n42969_ = ~new_n40957_ & new_n42968_;
  assign new_n42970_ = pi1155 & ~new_n40887_;
  assign new_n42971_ = ~pi1154 & ~new_n42970_;
  assign new_n42972_ = ~new_n42969_ & new_n42971_;
  assign new_n42973_ = ~pi1156 & ~new_n42972_;
  assign new_n42974_ = pi1155 & ~new_n40959_;
  assign new_n42975_ = pi1154 & ~new_n42974_;
  assign new_n42976_ = new_n42422_ & new_n42975_;
  assign new_n42977_ = new_n42973_ & ~new_n42976_;
  assign new_n42978_ = ~pi1155 & new_n40926_;
  assign new_n42979_ = ~new_n40886_ & new_n40915_;
  assign new_n42980_ = ~new_n42978_ & ~new_n42979_;
  assign new_n42981_ = ~pi1154 & ~new_n42980_;
  assign new_n42982_ = pi1156 & ~new_n42981_;
  assign new_n42983_ = new_n40937_ & new_n42975_;
  assign new_n42984_ = new_n42982_ & ~new_n42983_;
  assign new_n42985_ = pi0211 & ~new_n42984_;
  assign new_n42986_ = ~new_n42977_ & new_n42985_;
  assign new_n42987_ = pi1155 & ~new_n40992_;
  assign new_n42988_ = ~pi1154 & ~new_n42987_;
  assign new_n42989_ = new_n40926_ & new_n42988_;
  assign new_n42990_ = new_n40918_ & new_n42975_;
  assign new_n42991_ = ~new_n40889_ & new_n42990_;
  assign new_n42992_ = ~new_n42989_ & ~new_n42991_;
  assign new_n42993_ = new_n42982_ & new_n42992_;
  assign new_n42994_ = ~new_n42968_ & new_n42988_;
  assign new_n42995_ = ~new_n42990_ & ~new_n42994_;
  assign new_n42996_ = new_n42973_ & new_n42995_;
  assign new_n42997_ = ~pi0211 & ~new_n42996_;
  assign new_n42998_ = ~new_n42993_ & new_n42997_;
  assign new_n42999_ = ~pi0219 & ~new_n42998_;
  assign new_n43000_ = ~new_n42986_ & new_n42999_;
  assign new_n43001_ = pi1155 & new_n40885_;
  assign new_n43002_ = pi1154 & new_n41043_;
  assign new_n43003_ = ~new_n43001_ & new_n43002_;
  assign new_n43004_ = ~new_n42994_ & ~new_n43003_;
  assign new_n43005_ = ~pi1156 & ~new_n43004_;
  assign new_n43006_ = ~new_n40891_ & new_n43003_;
  assign new_n43007_ = ~new_n42989_ & ~new_n43006_;
  assign new_n43008_ = new_n38479_ & ~new_n43007_;
  assign new_n43009_ = ~pi1154 & new_n41032_;
  assign new_n43010_ = ~new_n40994_ & ~new_n43009_;
  assign new_n43011_ = new_n38483_ & ~new_n43001_;
  assign new_n43012_ = ~new_n43010_ & new_n43011_;
  assign new_n43013_ = pi0219 & ~new_n43012_;
  assign new_n43014_ = ~new_n43008_ & new_n43013_;
  assign new_n43015_ = ~new_n43005_ & new_n43014_;
  assign new_n43016_ = ~pi0263 & ~new_n43015_;
  assign new_n43017_ = ~new_n43000_ & new_n43016_;
  assign new_n43018_ = new_n40990_ & ~new_n43017_;
  assign new_n43019_ = ~new_n42967_ & new_n43018_;
  assign new_n43020_ = pi1155 & ~new_n39000_;
  assign new_n43021_ = new_n41092_ & ~new_n43020_;
  assign new_n43022_ = ~pi1154 & new_n42809_;
  assign new_n43023_ = ~new_n43021_ & ~new_n43022_;
  assign new_n43024_ = ~new_n41112_ & new_n43023_;
  assign new_n43025_ = new_n38479_ & ~new_n43024_;
  assign new_n43026_ = ~pi1154 & ~new_n38655_;
  assign new_n43027_ = new_n38556_ & ~new_n38557_;
  assign new_n43028_ = pi1154 & ~new_n43027_;
  assign new_n43029_ = pi1091 & new_n38483_;
  assign new_n43030_ = ~new_n43028_ & new_n43029_;
  assign new_n43031_ = ~new_n43026_ & new_n43030_;
  assign new_n43032_ = ~new_n41062_ & ~new_n42816_;
  assign new_n43033_ = ~pi1156 & ~new_n38558_;
  assign new_n43034_ = ~new_n43032_ & new_n43033_;
  assign new_n43035_ = pi0219 & ~new_n43034_;
  assign new_n43036_ = ~new_n43031_ & new_n43035_;
  assign new_n43037_ = ~new_n43025_ & new_n43036_;
  assign new_n43038_ = ~pi0211 & ~new_n43023_;
  assign new_n43039_ = new_n38548_ & ~new_n39112_;
  assign new_n43040_ = new_n42561_ & ~new_n43039_;
  assign new_n43041_ = ~new_n38659_ & new_n43040_;
  assign new_n43042_ = ~new_n43038_ & ~new_n43041_;
  assign new_n43043_ = pi1156 & ~new_n43042_;
  assign new_n43044_ = ~new_n38659_ & ~new_n43032_;
  assign new_n43045_ = pi0211 & new_n43044_;
  assign new_n43046_ = ~new_n38558_ & ~new_n38982_;
  assign new_n43047_ = new_n42610_ & new_n43046_;
  assign new_n43048_ = ~new_n43045_ & ~new_n43047_;
  assign new_n43049_ = ~pi1156 & ~new_n43048_;
  assign new_n43050_ = ~pi0219 & ~new_n43049_;
  assign new_n43051_ = ~new_n43043_ & new_n43050_;
  assign new_n43052_ = ~new_n43037_ & ~new_n43051_;
  assign new_n43053_ = ~pi0263 & ~new_n43052_;
  assign new_n43054_ = ~new_n38627_ & new_n43026_;
  assign new_n43055_ = ~new_n38548_ & ~new_n38594_;
  assign new_n43056_ = pi1154 & ~new_n43055_;
  assign new_n43057_ = pi1156 & ~new_n43056_;
  assign new_n43058_ = ~new_n43054_ & new_n43057_;
  assign new_n43059_ = ~pi1156 & new_n43044_;
  assign new_n43060_ = pi0211 & ~new_n43059_;
  assign new_n43061_ = ~new_n43058_ & new_n43060_;
  assign new_n43062_ = ~new_n38563_ & new_n39483_;
  assign new_n43063_ = ~new_n38982_ & ~new_n43062_;
  assign new_n43064_ = ~pi0211 & ~new_n43063_;
  assign new_n43065_ = ~pi0219 & ~new_n43064_;
  assign new_n43066_ = ~new_n43061_ & new_n43065_;
  assign new_n43067_ = pi1154 & ~new_n38560_;
  assign new_n43068_ = pi1156 & ~new_n43067_;
  assign new_n43069_ = ~pi0299 & ~new_n43068_;
  assign new_n43070_ = ~pi1154 & new_n38561_;
  assign new_n43071_ = ~new_n39904_ & ~new_n43070_;
  assign new_n43072_ = ~new_n43069_ & new_n43071_;
  assign new_n43073_ = pi1156 & ~new_n43072_;
  assign new_n43074_ = ~new_n43046_ & new_n43069_;
  assign new_n43075_ = pi0219 & ~new_n43074_;
  assign new_n43076_ = ~new_n43073_ & new_n43075_;
  assign new_n43077_ = pi0263 & pi1091;
  assign new_n43078_ = ~new_n43076_ & new_n43077_;
  assign new_n43079_ = ~new_n43066_ & new_n43078_;
  assign new_n43080_ = ~new_n43053_ & ~new_n43079_;
  assign new_n43081_ = ~new_n40990_ & ~new_n43080_;
  assign new_n43082_ = ~po1038 & ~new_n43081_;
  assign new_n43083_ = ~new_n43019_ & new_n43082_;
  assign new_n43084_ = pi0211 & new_n40868_;
  assign new_n43085_ = ~pi0211 & ~new_n42816_;
  assign new_n43086_ = ~new_n38484_ & ~new_n43085_;
  assign new_n43087_ = ~new_n43084_ & new_n43086_;
  assign new_n43088_ = ~new_n40877_ & ~new_n43087_;
  assign new_n43089_ = ~pi0219 & ~new_n43088_;
  assign new_n43090_ = ~pi0263 & ~new_n42729_;
  assign new_n43091_ = ~new_n43089_ & new_n43090_;
  assign new_n43092_ = ~new_n38484_ & ~new_n42707_;
  assign new_n43093_ = ~new_n43084_ & ~new_n43092_;
  assign new_n43094_ = new_n42458_ & ~new_n43093_;
  assign new_n43095_ = pi0263 & ~new_n42455_;
  assign new_n43096_ = ~new_n43094_ & new_n43095_;
  assign new_n43097_ = ~new_n43091_ & ~new_n43096_;
  assign new_n43098_ = pi0219 & ~new_n38483_;
  assign new_n43099_ = pi1091 & new_n43098_;
  assign new_n43100_ = new_n40990_ & ~new_n43099_;
  assign new_n43101_ = ~new_n43097_ & new_n43100_;
  assign new_n43102_ = ~pi0219 & ~new_n38484_;
  assign new_n43103_ = ~new_n38498_ & new_n43102_;
  assign new_n43104_ = ~new_n43098_ & ~new_n43103_;
  assign new_n43105_ = pi1091 & ~new_n43104_;
  assign new_n43106_ = pi0263 & ~pi1091;
  assign new_n43107_ = ~new_n43105_ & ~new_n43106_;
  assign new_n43108_ = ~new_n40990_ & new_n43107_;
  assign new_n43109_ = po1038 & ~new_n43108_;
  assign new_n43110_ = ~new_n43101_ & new_n43109_;
  assign new_n43111_ = new_n41153_ & ~new_n43110_;
  assign new_n43112_ = ~new_n43083_ & new_n43111_;
  assign new_n43113_ = ~po1038 & new_n43080_;
  assign new_n43114_ = po1038 & ~new_n43107_;
  assign new_n43115_ = ~new_n41153_ & ~new_n43114_;
  assign new_n43116_ = ~new_n43113_ & new_n43115_;
  assign new_n43117_ = ~pi0230 & ~new_n43116_;
  assign new_n43118_ = ~new_n43112_ & new_n43117_;
  assign new_n43119_ = ~new_n38559_ & new_n38564_;
  assign new_n43120_ = ~pi1156 & ~new_n43119_;
  assign new_n43121_ = new_n38741_ & ~new_n39113_;
  assign new_n43122_ = ~new_n43120_ & new_n43121_;
  assign new_n43123_ = ~new_n38510_ & ~new_n43122_;
  assign new_n43124_ = pi0211 & ~new_n43123_;
  assign new_n43125_ = new_n43065_ & ~new_n43124_;
  assign new_n43126_ = pi1156 & new_n39904_;
  assign new_n43127_ = pi0219 & ~new_n43126_;
  assign new_n43128_ = ~new_n43122_ & new_n43127_;
  assign new_n43129_ = ~po1038 & ~new_n43128_;
  assign new_n43130_ = ~new_n43125_ & new_n43129_;
  assign new_n43131_ = po1038 & new_n43104_;
  assign new_n43132_ = pi0230 & ~new_n43131_;
  assign new_n43133_ = ~new_n43130_ & new_n43132_;
  assign po0420 = ~new_n43118_ & ~new_n43133_;
  assign new_n43135_ = pi0264 & ~new_n40872_;
  assign new_n43136_ = ~pi0796 & new_n40872_;
  assign new_n43137_ = ~pi1091 & ~new_n43136_;
  assign new_n43138_ = ~new_n43135_ & new_n43137_;
  assign new_n43139_ = pi1091 & pi1142;
  assign new_n43140_ = ~new_n43138_ & ~new_n43139_;
  assign new_n43141_ = pi0200 & ~new_n43140_;
  assign new_n43142_ = pi1091 & pi1141;
  assign new_n43143_ = ~new_n43138_ & ~new_n43142_;
  assign new_n43144_ = ~pi0200 & ~new_n43143_;
  assign new_n43145_ = ~pi0199 & ~new_n43144_;
  assign new_n43146_ = ~new_n43141_ & new_n43145_;
  assign new_n43147_ = pi0264 & ~new_n40861_;
  assign new_n43148_ = ~pi0796 & new_n40861_;
  assign new_n43149_ = ~pi1091 & ~new_n43148_;
  assign new_n43150_ = ~new_n43147_ & new_n43149_;
  assign new_n43151_ = pi1091 & pi1143;
  assign new_n43152_ = ~pi0200 & new_n43151_;
  assign new_n43153_ = pi0199 & ~new_n43152_;
  assign new_n43154_ = ~new_n43150_ & new_n43153_;
  assign new_n43155_ = new_n16479_ & ~new_n43154_;
  assign new_n43156_ = ~new_n43146_ & new_n43155_;
  assign new_n43157_ = pi0211 & ~new_n43140_;
  assign new_n43158_ = ~pi0211 & ~new_n43143_;
  assign new_n43159_ = ~pi0219 & ~new_n43158_;
  assign new_n43160_ = ~new_n43157_ & new_n43159_;
  assign new_n43161_ = pi0219 & ~new_n42610_;
  assign new_n43162_ = ~new_n39377_ & ~new_n43161_;
  assign new_n43163_ = ~new_n43150_ & ~new_n43162_;
  assign new_n43164_ = ~new_n16479_ & ~new_n43163_;
  assign new_n43165_ = ~new_n43160_ & new_n43164_;
  assign new_n43166_ = ~new_n43156_ & ~new_n43165_;
  assign new_n43167_ = ~pi0230 & ~new_n43166_;
  assign new_n43168_ = ~pi0199 & pi1141;
  assign new_n43169_ = new_n39382_ & ~new_n43168_;
  assign new_n43170_ = ~new_n38444_ & ~new_n43169_;
  assign new_n43171_ = new_n16479_ & ~new_n43170_;
  assign new_n43172_ = ~pi0211 & pi1141;
  assign new_n43173_ = ~pi0219 & ~new_n38458_;
  assign new_n43174_ = ~new_n43172_ & new_n43173_;
  assign new_n43175_ = ~new_n39377_ & ~new_n43174_;
  assign new_n43176_ = ~new_n16479_ & ~new_n43175_;
  assign new_n43177_ = pi0230 & ~new_n43176_;
  assign new_n43178_ = ~new_n43171_ & new_n43177_;
  assign po0421 = new_n43167_ | new_n43178_;
  assign new_n43180_ = pi0265 & ~new_n40872_;
  assign new_n43181_ = ~pi0819 & new_n40872_;
  assign new_n43182_ = ~pi1091 & ~new_n43181_;
  assign new_n43183_ = ~new_n43180_ & new_n43182_;
  assign new_n43184_ = ~new_n43151_ & ~new_n43183_;
  assign new_n43185_ = pi0200 & ~new_n43184_;
  assign new_n43186_ = ~new_n43139_ & ~new_n43183_;
  assign new_n43187_ = ~pi0200 & ~new_n43186_;
  assign new_n43188_ = ~pi0199 & ~new_n43187_;
  assign new_n43189_ = ~new_n43185_ & new_n43188_;
  assign new_n43190_ = pi0265 & ~new_n40861_;
  assign new_n43191_ = ~pi0819 & new_n40861_;
  assign new_n43192_ = ~pi1091 & ~new_n43191_;
  assign new_n43193_ = ~new_n43190_ & new_n43192_;
  assign new_n43194_ = pi1091 & pi1144;
  assign new_n43195_ = ~pi0200 & new_n43194_;
  assign new_n43196_ = pi0199 & ~new_n43195_;
  assign new_n43197_ = ~new_n43193_ & new_n43196_;
  assign new_n43198_ = new_n16479_ & ~new_n43197_;
  assign new_n43199_ = ~new_n43189_ & new_n43198_;
  assign new_n43200_ = pi0211 & ~new_n43184_;
  assign new_n43201_ = ~pi0211 & ~new_n43186_;
  assign new_n43202_ = ~pi0219 & ~new_n43201_;
  assign new_n43203_ = ~new_n43200_ & new_n43202_;
  assign new_n43204_ = ~new_n40778_ & ~new_n43161_;
  assign new_n43205_ = ~new_n43193_ & ~new_n43204_;
  assign new_n43206_ = ~new_n16479_ & ~new_n43205_;
  assign new_n43207_ = ~new_n43203_ & new_n43206_;
  assign new_n43208_ = ~new_n43199_ & ~new_n43207_;
  assign new_n43209_ = ~pi0230 & ~new_n43208_;
  assign new_n43210_ = ~new_n38443_ & new_n40783_;
  assign new_n43211_ = ~new_n38437_ & ~new_n43210_;
  assign new_n43212_ = new_n16479_ & ~new_n43211_;
  assign new_n43213_ = ~pi0211 & pi1142;
  assign new_n43214_ = ~pi0219 & ~new_n38418_;
  assign new_n43215_ = ~new_n43213_ & new_n43214_;
  assign new_n43216_ = ~new_n40778_ & ~new_n43215_;
  assign new_n43217_ = ~new_n16479_ & ~new_n43216_;
  assign new_n43218_ = pi0230 & ~new_n43217_;
  assign new_n43219_ = ~new_n43212_ & new_n43218_;
  assign po0422 = new_n43209_ | new_n43219_;
  assign new_n43221_ = ~pi0211 & pi1136;
  assign new_n43222_ = pi0219 & ~new_n43221_;
  assign new_n43223_ = pi0211 & ~pi1135;
  assign new_n43224_ = ~new_n43222_ & ~new_n43223_;
  assign new_n43225_ = ~new_n10730_ & new_n43224_;
  assign new_n43226_ = pi0299 & new_n43225_;
  assign new_n43227_ = pi0199 & pi1136;
  assign new_n43228_ = ~pi0200 & ~new_n43227_;
  assign new_n43229_ = ~pi0199 & pi1135;
  assign new_n43230_ = pi0200 & ~new_n43229_;
  assign new_n43231_ = ~pi0299 & ~new_n43230_;
  assign new_n43232_ = ~new_n43228_ & new_n43231_;
  assign new_n43233_ = ~new_n43226_ & ~new_n43232_;
  assign new_n43234_ = ~po1038 & ~new_n43233_;
  assign new_n43235_ = po1038 & new_n43225_;
  assign new_n43236_ = pi0230 & ~new_n43235_;
  assign new_n43237_ = ~new_n43234_ & new_n43236_;
  assign new_n43238_ = ~pi0948 & new_n40872_;
  assign new_n43239_ = ~pi0266 & ~new_n40872_;
  assign new_n43240_ = ~pi1091 & ~new_n43239_;
  assign new_n43241_ = ~new_n43238_ & new_n43240_;
  assign new_n43242_ = ~pi0199 & ~new_n43241_;
  assign new_n43243_ = pi1091 & pi1136;
  assign new_n43244_ = ~pi0948 & new_n40861_;
  assign new_n43245_ = ~pi0266 & ~new_n40861_;
  assign new_n43246_ = ~pi1091 & ~new_n43245_;
  assign new_n43247_ = ~new_n43244_ & new_n43246_;
  assign new_n43248_ = pi0199 & ~new_n43247_;
  assign new_n43249_ = ~new_n43243_ & new_n43248_;
  assign new_n43250_ = ~new_n43242_ & ~new_n43249_;
  assign new_n43251_ = ~pi0200 & new_n43250_;
  assign new_n43252_ = pi1091 & pi1135;
  assign new_n43253_ = new_n43242_ & ~new_n43252_;
  assign new_n43254_ = pi0200 & ~new_n43248_;
  assign new_n43255_ = ~new_n43253_ & new_n43254_;
  assign new_n43256_ = ~new_n43251_ & ~new_n43255_;
  assign new_n43257_ = new_n16479_ & ~new_n43256_;
  assign new_n43258_ = ~new_n43161_ & ~new_n43222_;
  assign new_n43259_ = ~new_n43247_ & ~new_n43258_;
  assign new_n43260_ = ~new_n16479_ & ~new_n43259_;
  assign new_n43261_ = ~pi0219 & ~new_n43241_;
  assign new_n43262_ = pi1135 & new_n42561_;
  assign new_n43263_ = new_n43261_ & ~new_n43262_;
  assign new_n43264_ = new_n43260_ & ~new_n43263_;
  assign new_n43265_ = ~pi0230 & ~new_n43264_;
  assign new_n43266_ = ~new_n43257_ & new_n43265_;
  assign new_n43267_ = ~new_n43237_ & ~new_n43266_;
  assign new_n43268_ = ~pi1134 & ~new_n43267_;
  assign new_n43269_ = ~new_n16479_ & new_n43224_;
  assign new_n43270_ = new_n38607_ & ~new_n43227_;
  assign new_n43271_ = ~new_n43230_ & ~new_n43270_;
  assign new_n43272_ = new_n16479_ & new_n43271_;
  assign new_n43273_ = pi0230 & ~new_n43272_;
  assign new_n43274_ = ~new_n43269_ & new_n43273_;
  assign new_n43275_ = ~pi0199 & pi1091;
  assign new_n43276_ = ~new_n43250_ & ~new_n43275_;
  assign new_n43277_ = ~pi0200 & ~new_n43276_;
  assign new_n43278_ = ~new_n43255_ & ~new_n43277_;
  assign new_n43279_ = new_n16479_ & ~new_n43278_;
  assign new_n43280_ = pi1091 & ~new_n43223_;
  assign new_n43281_ = new_n43261_ & ~new_n43280_;
  assign new_n43282_ = new_n43260_ & ~new_n43281_;
  assign new_n43283_ = ~pi0230 & ~new_n43282_;
  assign new_n43284_ = ~new_n43279_ & new_n43283_;
  assign new_n43285_ = ~new_n43274_ & ~new_n43284_;
  assign new_n43286_ = pi1134 & ~new_n43285_;
  assign po0423 = ~new_n43268_ & ~new_n43286_;
  assign new_n43288_ = ~new_n42679_ & new_n42682_;
  assign new_n43289_ = new_n42748_ & ~new_n43288_;
  assign new_n43290_ = pi1154 & pi1155;
  assign new_n43291_ = ~new_n40900_ & new_n43290_;
  assign new_n43292_ = ~new_n42687_ & new_n43291_;
  assign new_n43293_ = ~new_n43289_ & ~new_n43292_;
  assign new_n43294_ = pi0211 & ~new_n43293_;
  assign new_n43295_ = pi1153 & new_n40902_;
  assign new_n43296_ = new_n38487_ & ~new_n42438_;
  assign new_n43297_ = ~new_n43295_ & new_n43296_;
  assign new_n43298_ = ~new_n42663_ & new_n43297_;
  assign new_n43299_ = new_n41032_ & new_n42657_;
  assign new_n43300_ = ~pi1155 & ~new_n43299_;
  assign new_n43301_ = ~new_n43288_ & new_n43300_;
  assign new_n43302_ = ~pi0267 & ~new_n43301_;
  assign new_n43303_ = ~new_n43298_ & new_n43302_;
  assign new_n43304_ = ~new_n43294_ & new_n43303_;
  assign new_n43305_ = ~new_n42422_ & ~new_n42445_;
  assign new_n43306_ = new_n40992_ & ~new_n43305_;
  assign new_n43307_ = pi1154 & ~new_n43306_;
  assign new_n43308_ = ~pi1154 & ~new_n41043_;
  assign new_n43309_ = ~new_n42534_ & new_n43308_;
  assign new_n43310_ = ~pi1155 & ~new_n43309_;
  assign new_n43311_ = ~new_n43307_ & new_n43310_;
  assign new_n43312_ = pi1155 & ~new_n42512_;
  assign new_n43313_ = new_n40885_ & ~new_n43009_;
  assign new_n43314_ = new_n43312_ & ~new_n43313_;
  assign new_n43315_ = ~new_n42532_ & new_n43314_;
  assign new_n43316_ = pi0267 & ~new_n43315_;
  assign new_n43317_ = ~new_n43311_ & new_n43316_;
  assign new_n43318_ = ~new_n43304_ & ~new_n43317_;
  assign new_n43319_ = pi0219 & ~new_n43318_;
  assign new_n43320_ = new_n40887_ & ~new_n43306_;
  assign new_n43321_ = new_n42957_ & ~new_n43320_;
  assign new_n43322_ = pi1154 & ~new_n43321_;
  assign new_n43323_ = ~pi1154 & ~new_n42433_;
  assign new_n43324_ = pi1155 & ~new_n43323_;
  assign new_n43325_ = new_n40932_ & ~new_n43324_;
  assign new_n43326_ = ~new_n43322_ & ~new_n43325_;
  assign new_n43327_ = ~pi1155 & ~new_n42767_;
  assign new_n43328_ = ~new_n43288_ & new_n43327_;
  assign new_n43329_ = pi0211 & ~new_n43328_;
  assign new_n43330_ = ~new_n43326_ & new_n43329_;
  assign new_n43331_ = pi1153 & ~new_n40957_;
  assign new_n43332_ = ~pi1155 & ~new_n43331_;
  assign new_n43333_ = ~pi1153 & ~new_n42939_;
  assign new_n43334_ = new_n43332_ & ~new_n43333_;
  assign new_n43335_ = ~new_n42769_ & ~new_n43295_;
  assign new_n43336_ = pi1155 & ~new_n43335_;
  assign new_n43337_ = pi1154 & ~new_n42940_;
  assign new_n43338_ = ~new_n43336_ & new_n43337_;
  assign new_n43339_ = ~new_n43334_ & new_n43338_;
  assign new_n43340_ = new_n42527_ & new_n43332_;
  assign new_n43341_ = ~pi1154 & ~new_n43336_;
  assign new_n43342_ = ~new_n43340_ & new_n43341_;
  assign new_n43343_ = ~pi0211 & ~new_n43342_;
  assign new_n43344_ = ~new_n43339_ & new_n43343_;
  assign new_n43345_ = ~pi0267 & ~new_n43344_;
  assign new_n43346_ = ~new_n43330_ & new_n43345_;
  assign new_n43347_ = new_n42979_ & new_n43312_;
  assign new_n43348_ = ~pi1153 & new_n40971_;
  assign new_n43349_ = ~new_n40959_ & ~new_n43348_;
  assign new_n43350_ = ~pi1155 & new_n40887_;
  assign new_n43351_ = ~new_n43349_ & new_n43350_;
  assign new_n43352_ = pi1154 & ~new_n43351_;
  assign new_n43353_ = ~new_n43347_ & new_n43352_;
  assign new_n43354_ = ~pi1154 & ~new_n42445_;
  assign new_n43355_ = ~new_n40918_ & new_n43354_;
  assign new_n43356_ = ~pi1155 & ~new_n43355_;
  assign new_n43357_ = ~new_n40937_ & new_n43354_;
  assign new_n43358_ = ~new_n43356_ & new_n43357_;
  assign new_n43359_ = ~new_n43353_ & ~new_n43358_;
  assign new_n43360_ = pi0211 & ~new_n43359_;
  assign new_n43361_ = pi1154 & new_n43349_;
  assign new_n43362_ = new_n43356_ & ~new_n43361_;
  assign new_n43363_ = ~new_n40910_ & ~new_n42750_;
  assign new_n43364_ = pi1154 & new_n40885_;
  assign new_n43365_ = pi1155 & ~new_n43364_;
  assign new_n43366_ = ~new_n43363_ & new_n43365_;
  assign new_n43367_ = ~pi0211 & ~new_n43366_;
  assign new_n43368_ = ~new_n43362_ & new_n43367_;
  assign new_n43369_ = pi0267 & ~new_n43368_;
  assign new_n43370_ = ~new_n43360_ & new_n43369_;
  assign new_n43371_ = ~pi0219 & ~new_n43370_;
  assign new_n43372_ = ~new_n43346_ & new_n43371_;
  assign new_n43373_ = ~new_n43319_ & ~new_n43372_;
  assign new_n43374_ = new_n40989_ & ~new_n43373_;
  assign new_n43375_ = pi1155 & ~new_n42549_;
  assign new_n43376_ = new_n42809_ & new_n43375_;
  assign new_n43377_ = ~pi1155 & ~new_n42698_;
  assign new_n43378_ = ~new_n42578_ & new_n43377_;
  assign new_n43379_ = ~new_n43376_ & ~new_n43378_;
  assign new_n43380_ = pi1154 & ~new_n43379_;
  assign new_n43381_ = ~new_n42807_ & new_n43375_;
  assign new_n43382_ = ~pi1155 & ~new_n39061_;
  assign new_n43383_ = pi1091 & new_n43382_;
  assign new_n43384_ = ~new_n43381_ & ~new_n43383_;
  assign new_n43385_ = ~pi1154 & ~new_n43384_;
  assign new_n43386_ = ~pi0219 & ~new_n43385_;
  assign new_n43387_ = ~new_n43380_ & new_n43386_;
  assign new_n43388_ = pi1091 & new_n43020_;
  assign new_n43389_ = ~new_n42548_ & new_n43388_;
  assign new_n43390_ = pi1154 & ~new_n43389_;
  assign new_n43391_ = ~pi0299 & new_n38947_;
  assign new_n43392_ = pi1091 & ~new_n43391_;
  assign new_n43393_ = new_n43390_ & new_n43392_;
  assign new_n43394_ = pi1153 & new_n38955_;
  assign new_n43395_ = new_n42816_ & ~new_n43394_;
  assign new_n43396_ = ~new_n39645_ & new_n43395_;
  assign new_n43397_ = pi0219 & ~new_n43396_;
  assign new_n43398_ = ~new_n43393_ & new_n43397_;
  assign new_n43399_ = ~new_n43387_ & ~new_n43398_;
  assign new_n43400_ = ~pi0211 & ~new_n43399_;
  assign new_n43401_ = ~pi1155 & ~new_n38948_;
  assign new_n43402_ = ~new_n38654_ & ~new_n43401_;
  assign new_n43403_ = ~new_n13062_ & ~new_n43402_;
  assign new_n43404_ = pi1155 & new_n38963_;
  assign new_n43405_ = pi1154 & ~new_n43404_;
  assign new_n43406_ = pi1091 & new_n43405_;
  assign new_n43407_ = ~new_n43403_ & new_n43406_;
  assign new_n43408_ = ~new_n38609_ & ~new_n41066_;
  assign new_n43409_ = new_n43395_ & ~new_n43408_;
  assign new_n43410_ = pi0211 & ~new_n43409_;
  assign new_n43411_ = ~new_n43407_ & new_n43410_;
  assign new_n43412_ = ~new_n43400_ & ~new_n43411_;
  assign new_n43413_ = pi0267 & ~new_n43412_;
  assign new_n43414_ = ~pi1154 & new_n38556_;
  assign new_n43415_ = ~new_n38630_ & ~new_n43414_;
  assign new_n43416_ = ~new_n38589_ & new_n43415_;
  assign new_n43417_ = pi1091 & new_n43416_;
  assign new_n43418_ = ~pi0211 & ~new_n43417_;
  assign new_n43419_ = pi1091 & ~pi1155;
  assign new_n43420_ = ~new_n38948_ & new_n43419_;
  assign new_n43421_ = new_n38488_ & ~new_n43420_;
  assign new_n43422_ = ~new_n43389_ & new_n43421_;
  assign new_n43423_ = ~pi0219 & ~new_n43422_;
  assign new_n43424_ = ~new_n43418_ & new_n43423_;
  assign new_n43425_ = new_n43391_ & new_n43419_;
  assign new_n43426_ = new_n43390_ & ~new_n43425_;
  assign new_n43427_ = pi1154 & ~new_n43426_;
  assign new_n43428_ = ~new_n38609_ & new_n42816_;
  assign new_n43429_ = ~new_n39644_ & new_n43428_;
  assign new_n43430_ = ~pi0211 & ~new_n43429_;
  assign new_n43431_ = ~new_n43427_ & new_n43430_;
  assign new_n43432_ = new_n43020_ & new_n43405_;
  assign new_n43433_ = ~new_n43426_ & ~new_n43432_;
  assign new_n43434_ = pi0211 & ~new_n43433_;
  assign new_n43435_ = pi0219 & ~new_n43434_;
  assign new_n43436_ = ~new_n43431_ & new_n43435_;
  assign new_n43437_ = ~new_n43424_ & ~new_n43436_;
  assign new_n43438_ = new_n38548_ & new_n42570_;
  assign new_n43439_ = ~new_n42783_ & ~new_n43438_;
  assign new_n43440_ = ~new_n43382_ & ~new_n43439_;
  assign new_n43441_ = pi0211 & ~pi1154;
  assign new_n43442_ = ~new_n43440_ & new_n43441_;
  assign new_n43443_ = ~pi0267 & ~new_n43442_;
  assign new_n43444_ = ~new_n43437_ & new_n43443_;
  assign new_n43445_ = ~new_n43413_ & ~new_n43444_;
  assign new_n43446_ = ~new_n40989_ & ~new_n43445_;
  assign new_n43447_ = ~po1038 & ~new_n43446_;
  assign new_n43448_ = ~new_n43374_ & new_n43447_;
  assign new_n43449_ = pi0267 & new_n42731_;
  assign new_n43450_ = ~pi0267 & ~new_n40879_;
  assign new_n43451_ = ~new_n42455_ & new_n43450_;
  assign new_n43452_ = new_n40989_ & ~new_n43451_;
  assign new_n43453_ = ~new_n43449_ & new_n43452_;
  assign new_n43454_ = ~pi0219 & ~new_n38488_;
  assign new_n43455_ = ~new_n38500_ & new_n43454_;
  assign new_n43456_ = ~new_n39273_ & ~new_n43455_;
  assign new_n43457_ = pi1091 & ~new_n43456_;
  assign new_n43458_ = ~pi0267 & ~pi1091;
  assign new_n43459_ = ~new_n40989_ & new_n43458_;
  assign new_n43460_ = ~new_n43457_ & ~new_n43459_;
  assign new_n43461_ = ~new_n43453_ & new_n43460_;
  assign new_n43462_ = po1038 & ~new_n43461_;
  assign new_n43463_ = new_n41153_ & ~new_n43462_;
  assign new_n43464_ = ~new_n43448_ & new_n43463_;
  assign new_n43465_ = ~po1038 & new_n43445_;
  assign new_n43466_ = ~new_n43457_ & ~new_n43458_;
  assign new_n43467_ = po1038 & ~new_n43466_;
  assign new_n43468_ = ~new_n41153_ & ~new_n43467_;
  assign new_n43469_ = ~new_n43465_ & new_n43468_;
  assign new_n43470_ = ~pi0230 & ~new_n43469_;
  assign new_n43471_ = ~new_n43464_ & new_n43470_;
  assign new_n43472_ = pi0219 & ~new_n38963_;
  assign new_n43473_ = ~pi1155 & new_n43394_;
  assign new_n43474_ = ~pi1154 & ~new_n43473_;
  assign new_n43475_ = ~new_n38948_ & ~new_n43474_;
  assign new_n43476_ = pi1155 & new_n39642_;
  assign new_n43477_ = ~new_n43475_ & ~new_n43476_;
  assign new_n43478_ = ~new_n43472_ & ~new_n43477_;
  assign new_n43479_ = pi0211 & ~new_n43478_;
  assign new_n43480_ = ~pi0199 & pi1154;
  assign new_n43481_ = pi0200 & ~new_n43480_;
  assign new_n43482_ = ~new_n38619_ & ~new_n38962_;
  assign new_n43483_ = ~new_n43481_ & new_n43482_;
  assign new_n43484_ = ~new_n38510_ & ~new_n43483_;
  assign new_n43485_ = pi0219 & ~new_n43484_;
  assign new_n43486_ = ~pi0219 & new_n43416_;
  assign new_n43487_ = ~pi0211 & ~new_n43486_;
  assign new_n43488_ = ~new_n43485_ & new_n43487_;
  assign new_n43489_ = ~po1038 & ~new_n43488_;
  assign new_n43490_ = ~new_n43479_ & new_n43489_;
  assign new_n43491_ = po1038 & new_n43456_;
  assign new_n43492_ = pi0230 & ~new_n43491_;
  assign new_n43493_ = ~new_n43490_ & new_n43492_;
  assign po0424 = ~new_n43471_ & ~new_n43493_;
  assign new_n43495_ = ~new_n42469_ & new_n42501_;
  assign new_n43496_ = ~new_n40898_ & new_n42513_;
  assign new_n43497_ = pi0219 & ~new_n42440_;
  assign new_n43498_ = ~new_n40892_ & new_n43497_;
  assign new_n43499_ = ~new_n43496_ & ~new_n43498_;
  assign new_n43500_ = ~po1038 & ~new_n42426_;
  assign new_n43501_ = new_n43499_ & new_n43500_;
  assign new_n43502_ = ~new_n43495_ & ~new_n43501_;
  assign new_n43503_ = ~pi1151 & ~new_n43502_;
  assign new_n43504_ = ~po1038 & ~new_n42528_;
  assign new_n43505_ = pi0219 & new_n41037_;
  assign new_n43506_ = new_n43504_ & ~new_n43505_;
  assign new_n43507_ = new_n42501_ & ~new_n42730_;
  assign new_n43508_ = ~new_n43506_ & ~new_n43507_;
  assign new_n43509_ = pi1151 & ~new_n43508_;
  assign new_n43510_ = ~new_n43503_ & ~new_n43509_;
  assign new_n43511_ = pi0268 & ~new_n43510_;
  assign new_n43512_ = po1038 & ~new_n42455_;
  assign new_n43513_ = ~new_n42498_ & new_n43512_;
  assign new_n43514_ = po1038 & ~new_n42729_;
  assign new_n43515_ = ~new_n42462_ & new_n43514_;
  assign new_n43516_ = new_n43513_ & ~new_n43515_;
  assign new_n43517_ = pi0219 & ~new_n40896_;
  assign new_n43518_ = ~new_n42486_ & ~new_n43517_;
  assign new_n43519_ = ~new_n40897_ & ~new_n43518_;
  assign new_n43520_ = ~po1038 & ~new_n40956_;
  assign new_n43521_ = new_n43519_ & new_n43520_;
  assign new_n43522_ = ~new_n43516_ & ~new_n43521_;
  assign new_n43523_ = ~pi1151 & new_n43522_;
  assign new_n43524_ = ~new_n40868_ & ~new_n43508_;
  assign new_n43525_ = ~new_n40946_ & new_n43504_;
  assign new_n43526_ = pi0219 & po1038;
  assign new_n43527_ = ~new_n40895_ & new_n43526_;
  assign new_n43528_ = ~new_n42458_ & ~new_n43527_;
  assign new_n43529_ = ~new_n43525_ & new_n43528_;
  assign new_n43530_ = ~new_n43524_ & ~new_n43529_;
  assign new_n43531_ = pi1151 & new_n43530_;
  assign new_n43532_ = ~pi0268 & ~new_n43531_;
  assign new_n43533_ = ~new_n43523_ & new_n43532_;
  assign new_n43534_ = ~new_n43511_ & ~new_n43533_;
  assign new_n43535_ = ~pi1152 & ~new_n43534_;
  assign new_n43536_ = ~new_n42469_ & new_n43514_;
  assign new_n43537_ = ~new_n40994_ & ~new_n42535_;
  assign new_n43538_ = ~new_n43499_ & ~new_n43537_;
  assign new_n43539_ = ~po1038 & ~new_n43538_;
  assign new_n43540_ = ~new_n40895_ & ~new_n42515_;
  assign new_n43541_ = new_n43539_ & ~new_n43540_;
  assign new_n43542_ = ~new_n43536_ & ~new_n43541_;
  assign new_n43543_ = ~pi1151 & ~new_n43542_;
  assign new_n43544_ = ~new_n40864_ & new_n43500_;
  assign new_n43545_ = ~new_n42730_ & new_n43514_;
  assign new_n43546_ = ~new_n43506_ & ~new_n43545_;
  assign new_n43547_ = ~new_n43544_ & new_n43546_;
  assign new_n43548_ = pi1151 & ~new_n43547_;
  assign new_n43549_ = pi0268 & ~new_n43548_;
  assign new_n43550_ = ~new_n43543_ & new_n43549_;
  assign new_n43551_ = ~new_n42439_ & ~new_n43519_;
  assign new_n43552_ = ~po1038 & ~new_n43551_;
  assign new_n43553_ = ~new_n43513_ & ~new_n43552_;
  assign new_n43554_ = ~pi1151 & ~new_n43553_;
  assign new_n43555_ = ~pi0219 & new_n40907_;
  assign new_n43556_ = ~new_n43497_ & ~new_n43555_;
  assign new_n43557_ = ~po1038 & ~new_n43556_;
  assign new_n43558_ = ~new_n42470_ & new_n43512_;
  assign new_n43559_ = ~new_n43516_ & ~new_n43558_;
  assign new_n43560_ = ~new_n43557_ & new_n43559_;
  assign new_n43561_ = pi1151 & ~new_n43560_;
  assign new_n43562_ = ~pi0268 & ~new_n43561_;
  assign new_n43563_ = ~new_n43554_ & new_n43562_;
  assign new_n43564_ = pi1152 & ~new_n43563_;
  assign new_n43565_ = ~new_n43550_ & new_n43564_;
  assign new_n43566_ = ~new_n43535_ & ~new_n43565_;
  assign new_n43567_ = pi1150 & ~new_n43566_;
  assign new_n43568_ = ~po1038 & ~new_n43499_;
  assign new_n43569_ = ~new_n43558_ & ~new_n43568_;
  assign new_n43570_ = pi1151 & ~new_n43569_;
  assign new_n43571_ = ~new_n42458_ & new_n43512_;
  assign new_n43572_ = ~pi0219 & ~new_n40932_;
  assign new_n43573_ = ~new_n40884_ & ~new_n43572_;
  assign new_n43574_ = new_n43557_ & new_n43573_;
  assign new_n43575_ = ~new_n43571_ & ~new_n43574_;
  assign new_n43576_ = ~pi1151 & ~new_n43575_;
  assign new_n43577_ = pi1152 & ~new_n43576_;
  assign new_n43578_ = ~new_n43570_ & new_n43577_;
  assign new_n43579_ = ~new_n42471_ & ~new_n43527_;
  assign new_n43580_ = ~new_n43539_ & new_n43579_;
  assign new_n43581_ = pi1151 & new_n43580_;
  assign new_n43582_ = ~pi1151 & new_n43529_;
  assign new_n43583_ = ~pi1152 & ~new_n43582_;
  assign new_n43584_ = ~new_n43581_ & new_n43583_;
  assign new_n43585_ = ~new_n43578_ & ~new_n43584_;
  assign new_n43586_ = ~pi0268 & ~new_n43585_;
  assign new_n43587_ = ~new_n42499_ & new_n43514_;
  assign new_n43588_ = pi0219 & ~new_n42532_;
  assign new_n43589_ = ~new_n42486_ & ~new_n43588_;
  assign new_n43590_ = new_n40915_ & ~new_n43589_;
  assign new_n43591_ = ~po1038 & ~new_n43590_;
  assign new_n43592_ = ~new_n43587_ & ~new_n43591_;
  assign new_n43593_ = pi1151 & new_n43592_;
  assign new_n43594_ = ~po1038 & ~new_n42535_;
  assign new_n43595_ = ~new_n43588_ & new_n43594_;
  assign new_n43596_ = ~new_n43515_ & ~new_n43595_;
  assign new_n43597_ = ~pi1151 & new_n43596_;
  assign new_n43598_ = pi1152 & ~new_n43597_;
  assign new_n43599_ = ~new_n43593_ & new_n43598_;
  assign new_n43600_ = ~po1038 & ~new_n42489_;
  assign new_n43601_ = ~new_n42486_ & new_n43600_;
  assign new_n43602_ = ~new_n42502_ & ~new_n43601_;
  assign new_n43603_ = pi1151 & new_n43602_;
  assign new_n43604_ = new_n40868_ & ~new_n43508_;
  assign new_n43605_ = ~pi1151 & ~new_n43604_;
  assign new_n43606_ = ~pi1152 & ~new_n43605_;
  assign new_n43607_ = ~new_n43603_ & new_n43606_;
  assign new_n43608_ = pi0268 & ~new_n43607_;
  assign new_n43609_ = ~new_n43599_ & new_n43608_;
  assign new_n43610_ = ~pi1150 & ~new_n43609_;
  assign new_n43611_ = ~new_n43586_ & new_n43610_;
  assign new_n43612_ = ~new_n43567_ & ~new_n43611_;
  assign new_n43613_ = new_n41152_ & ~new_n43612_;
  assign new_n43614_ = pi0268 & pi1152;
  assign new_n43615_ = ~pi0199 & new_n16479_;
  assign new_n43616_ = ~new_n40164_ & ~new_n43615_;
  assign new_n43617_ = ~pi0211 & ~new_n16479_;
  assign new_n43618_ = ~po1038 & new_n38548_;
  assign new_n43619_ = ~new_n43617_ & ~new_n43618_;
  assign new_n43620_ = pi1152 & ~new_n43619_;
  assign new_n43621_ = new_n43616_ & ~new_n43620_;
  assign new_n43622_ = ~pi1151 & new_n43619_;
  assign new_n43623_ = pi1150 & ~new_n43622_;
  assign new_n43624_ = ~new_n43621_ & new_n43623_;
  assign new_n43625_ = ~new_n43614_ & new_n43624_;
  assign new_n43626_ = ~new_n16479_ & new_n42598_;
  assign new_n43627_ = ~po1038 & new_n38618_;
  assign new_n43628_ = ~new_n43626_ & ~new_n43627_;
  assign new_n43629_ = pi1151 & ~new_n43628_;
  assign new_n43630_ = pi1152 & new_n43629_;
  assign new_n43631_ = ~po1038 & ~new_n11448_;
  assign new_n43632_ = po1038 & new_n11446_;
  assign new_n43633_ = ~new_n43631_ & ~new_n43632_;
  assign new_n43634_ = pi1151 & ~new_n43633_;
  assign new_n43635_ = ~pi1152 & ~new_n43634_;
  assign new_n43636_ = ~pi1151 & new_n42389_;
  assign new_n43637_ = ~pi1150 & ~new_n43636_;
  assign new_n43638_ = ~new_n43635_ & new_n43637_;
  assign new_n43639_ = ~new_n43630_ & new_n43638_;
  assign new_n43640_ = ~new_n43625_ & ~new_n43639_;
  assign new_n43641_ = pi1091 & ~new_n43640_;
  assign new_n43642_ = pi1152 & new_n43624_;
  assign new_n43643_ = pi1091 & ~new_n43642_;
  assign new_n43644_ = pi0268 & ~new_n43643_;
  assign new_n43645_ = ~new_n43641_ & ~new_n43644_;
  assign new_n43646_ = ~new_n41152_ & ~new_n43645_;
  assign new_n43647_ = ~pi0230 & ~new_n43646_;
  assign new_n43648_ = ~new_n43613_ & new_n43647_;
  assign new_n43649_ = pi0230 & ~new_n43624_;
  assign new_n43650_ = ~new_n43639_ & new_n43649_;
  assign po0425 = ~new_n43648_ & ~new_n43650_;
  assign new_n43652_ = ~pi0199 & pi1137;
  assign new_n43653_ = pi0200 & ~new_n43652_;
  assign new_n43654_ = ~pi0199 & pi1136;
  assign new_n43655_ = pi0199 & pi1138;
  assign new_n43656_ = ~pi0200 & ~new_n43655_;
  assign new_n43657_ = ~new_n43654_ & new_n43656_;
  assign new_n43658_ = ~new_n43653_ & ~new_n43657_;
  assign new_n43659_ = new_n16479_ & ~new_n43658_;
  assign new_n43660_ = ~pi0211 & pi1138;
  assign new_n43661_ = pi0219 & new_n43660_;
  assign new_n43662_ = pi0211 & pi1137;
  assign new_n43663_ = ~new_n43221_ & ~new_n43662_;
  assign new_n43664_ = ~pi0219 & ~new_n43663_;
  assign new_n43665_ = ~new_n43661_ & ~new_n43664_;
  assign new_n43666_ = ~new_n16479_ & new_n43665_;
  assign new_n43667_ = ~new_n43659_ & ~new_n43666_;
  assign new_n43668_ = pi0230 & ~new_n43667_;
  assign new_n43669_ = ~pi0200 & new_n43243_;
  assign new_n43670_ = pi1137 & new_n41091_;
  assign new_n43671_ = ~new_n43669_ & ~new_n43670_;
  assign new_n43672_ = new_n43615_ & new_n43671_;
  assign new_n43673_ = pi1091 & ~new_n43663_;
  assign new_n43674_ = new_n40164_ & ~new_n43673_;
  assign new_n43675_ = ~new_n43672_ & ~new_n43674_;
  assign new_n43676_ = pi0269 & ~new_n40872_;
  assign new_n43677_ = ~pi0817 & new_n40872_;
  assign new_n43678_ = ~pi1091 & ~new_n43677_;
  assign new_n43679_ = ~new_n43676_ & new_n43678_;
  assign new_n43680_ = ~new_n43675_ & ~new_n43679_;
  assign new_n43681_ = pi0269 & ~new_n40861_;
  assign new_n43682_ = ~pi0817 & new_n40861_;
  assign new_n43683_ = ~pi1091 & ~new_n43682_;
  assign new_n43684_ = ~new_n43681_ & new_n43683_;
  assign new_n43685_ = pi1138 & new_n42610_;
  assign new_n43686_ = pi0219 & ~new_n16479_;
  assign new_n43687_ = ~new_n43685_ & new_n43686_;
  assign new_n43688_ = ~pi0200 & pi1091;
  assign new_n43689_ = pi1138 & new_n43688_;
  assign new_n43690_ = pi0199 & ~new_n43689_;
  assign new_n43691_ = new_n16479_ & new_n43690_;
  assign new_n43692_ = ~new_n43687_ & ~new_n43691_;
  assign new_n43693_ = ~new_n43684_ & ~new_n43692_;
  assign new_n43694_ = ~new_n43680_ & ~new_n43693_;
  assign new_n43695_ = ~pi0230 & ~new_n43694_;
  assign po0426 = ~new_n43668_ & ~new_n43695_;
  assign new_n43697_ = pi0270 & ~new_n40872_;
  assign new_n43698_ = ~pi0805 & new_n40872_;
  assign new_n43699_ = ~pi1091 & ~new_n43698_;
  assign new_n43700_ = ~new_n43697_ & new_n43699_;
  assign new_n43701_ = ~pi0211 & pi1139;
  assign new_n43702_ = pi0211 & pi1140;
  assign new_n43703_ = ~new_n43701_ & ~new_n43702_;
  assign new_n43704_ = pi1091 & ~new_n43703_;
  assign new_n43705_ = new_n40164_ & ~new_n43704_;
  assign new_n43706_ = pi1091 & pi1140;
  assign new_n43707_ = pi0200 & new_n43706_;
  assign new_n43708_ = pi1139 & new_n43688_;
  assign new_n43709_ = ~new_n43707_ & ~new_n43708_;
  assign new_n43710_ = new_n43615_ & new_n43709_;
  assign new_n43711_ = ~new_n43705_ & ~new_n43710_;
  assign new_n43712_ = ~new_n43700_ & ~new_n43711_;
  assign new_n43713_ = pi0270 & ~new_n40861_;
  assign new_n43714_ = ~pi0805 & new_n40861_;
  assign new_n43715_ = ~pi1091 & ~new_n43714_;
  assign new_n43716_ = ~new_n43713_ & new_n43715_;
  assign new_n43717_ = new_n42610_ & new_n43172_;
  assign new_n43718_ = new_n43686_ & ~new_n43717_;
  assign new_n43719_ = ~pi0200 & new_n43142_;
  assign new_n43720_ = pi0199 & ~new_n43719_;
  assign new_n43721_ = new_n16479_ & new_n43720_;
  assign new_n43722_ = ~new_n43718_ & ~new_n43721_;
  assign new_n43723_ = ~new_n43716_ & ~new_n43722_;
  assign new_n43724_ = ~pi0230 & ~new_n43723_;
  assign new_n43725_ = ~new_n43712_ & new_n43724_;
  assign new_n43726_ = ~pi0199 & pi1140;
  assign new_n43727_ = pi0200 & ~new_n43726_;
  assign new_n43728_ = ~pi0199 & pi1139;
  assign new_n43729_ = pi0199 & pi1141;
  assign new_n43730_ = ~pi0200 & ~new_n43729_;
  assign new_n43731_ = ~new_n43728_ & new_n43730_;
  assign new_n43732_ = ~new_n43727_ & ~new_n43731_;
  assign new_n43733_ = new_n16479_ & ~new_n43732_;
  assign new_n43734_ = pi0219 & ~new_n43172_;
  assign new_n43735_ = ~pi0219 & new_n43703_;
  assign new_n43736_ = ~new_n43734_ & ~new_n43735_;
  assign new_n43737_ = ~new_n16479_ & ~new_n43736_;
  assign new_n43738_ = pi0230 & ~new_n43737_;
  assign new_n43739_ = ~new_n43733_ & new_n43738_;
  assign po0427 = new_n43725_ | new_n43739_;
  assign new_n43741_ = ~pi0271 & ~new_n40893_;
  assign new_n43742_ = ~new_n40865_ & ~new_n43741_;
  assign new_n43743_ = pi0219 & ~new_n43742_;
  assign new_n43744_ = ~pi1091 & ~new_n40874_;
  assign new_n43745_ = pi0271 & ~new_n43744_;
  assign new_n43746_ = ~pi0271 & ~new_n40875_;
  assign new_n43747_ = ~new_n43745_ & ~new_n43746_;
  assign new_n43748_ = pi1091 & pi1146;
  assign new_n43749_ = ~new_n43747_ & ~new_n43748_;
  assign new_n43750_ = ~pi0211 & new_n43748_;
  assign new_n43751_ = ~new_n43749_ & ~new_n43750_;
  assign new_n43752_ = pi1091 & new_n39369_;
  assign new_n43753_ = ~pi0219 & ~new_n43752_;
  assign new_n43754_ = ~new_n43751_ & new_n43753_;
  assign new_n43755_ = ~new_n43743_ & ~new_n43754_;
  assign new_n43756_ = ~pi0211 & pi1147;
  assign new_n43757_ = new_n42456_ & new_n43756_;
  assign new_n43758_ = ~new_n16479_ & ~new_n43757_;
  assign new_n43759_ = ~new_n43755_ & new_n43758_;
  assign new_n43760_ = pi0199 & ~new_n43742_;
  assign new_n43761_ = ~pi0199 & new_n43749_;
  assign new_n43762_ = ~new_n43760_ & ~new_n43761_;
  assign new_n43763_ = pi0200 & ~new_n43762_;
  assign new_n43764_ = pi1091 & pi1145;
  assign new_n43765_ = ~pi0199 & ~new_n43764_;
  assign new_n43766_ = ~new_n43747_ & new_n43765_;
  assign new_n43767_ = ~new_n43760_ & ~new_n43766_;
  assign new_n43768_ = pi1147 & new_n41075_;
  assign new_n43769_ = ~pi0200 & ~new_n43768_;
  assign new_n43770_ = ~new_n43767_ & new_n43769_;
  assign new_n43771_ = ~new_n43763_ & ~new_n43770_;
  assign new_n43772_ = new_n16479_ & ~new_n43771_;
  assign new_n43773_ = ~new_n43759_ & ~new_n43772_;
  assign new_n43774_ = ~pi0230 & ~new_n43773_;
  assign new_n43775_ = ~pi0200 & ~new_n39386_;
  assign new_n43776_ = new_n40339_ & ~new_n43775_;
  assign new_n43777_ = pi1147 & new_n42386_;
  assign new_n43778_ = ~new_n40223_ & ~new_n40238_;
  assign new_n43779_ = ~pi0219 & ~new_n43778_;
  assign new_n43780_ = ~new_n43777_ & ~new_n43779_;
  assign new_n43781_ = ~new_n43776_ & new_n43780_;
  assign new_n43782_ = ~po1038 & ~new_n43781_;
  assign new_n43783_ = pi0219 & ~new_n43756_;
  assign new_n43784_ = ~new_n39369_ & new_n41505_;
  assign new_n43785_ = ~new_n43783_ & ~new_n43784_;
  assign new_n43786_ = po1038 & new_n43785_;
  assign new_n43787_ = pi0230 & ~new_n43786_;
  assign new_n43788_ = ~new_n43782_ & new_n43787_;
  assign po0428 = ~new_n43774_ & ~new_n43788_;
  assign new_n43790_ = pi1150 & ~new_n43560_;
  assign new_n43791_ = ~pi1150 & ~new_n43530_;
  assign new_n43792_ = pi1149 & ~new_n43791_;
  assign new_n43793_ = ~new_n43790_ & new_n43792_;
  assign new_n43794_ = pi1150 & ~new_n43553_;
  assign new_n43795_ = ~pi1150 & ~new_n43522_;
  assign new_n43796_ = ~pi1149 & ~new_n43795_;
  assign new_n43797_ = ~new_n43794_ & new_n43796_;
  assign new_n43798_ = ~new_n43793_ & ~new_n43797_;
  assign new_n43799_ = pi1148 & ~new_n43798_;
  assign new_n43800_ = ~pi1150 & ~new_n43580_;
  assign new_n43801_ = pi1150 & new_n43569_;
  assign new_n43802_ = pi1149 & ~new_n43801_;
  assign new_n43803_ = ~new_n43800_ & new_n43802_;
  assign new_n43804_ = pi1150 & new_n43575_;
  assign new_n43805_ = ~pi1150 & ~new_n43529_;
  assign new_n43806_ = ~pi1149 & ~new_n43805_;
  assign new_n43807_ = ~new_n43804_ & new_n43806_;
  assign new_n43808_ = ~pi1148 & ~new_n43807_;
  assign new_n43809_ = ~new_n43803_ & new_n43808_;
  assign new_n43810_ = ~new_n43799_ & ~new_n43809_;
  assign new_n43811_ = pi0283 & ~new_n43810_;
  assign new_n43812_ = ~po1038 & new_n38539_;
  assign new_n43813_ = ~new_n40164_ & ~new_n43812_;
  assign new_n43814_ = ~new_n43617_ & new_n43813_;
  assign new_n43815_ = pi1150 & ~new_n43814_;
  assign new_n43816_ = pi1149 & ~new_n43815_;
  assign new_n43817_ = new_n43616_ & new_n43816_;
  assign new_n43818_ = po1038 & new_n10730_;
  assign new_n43819_ = ~new_n13065_ & ~new_n43818_;
  assign new_n43820_ = ~pi1150 & new_n43819_;
  assign new_n43821_ = ~new_n43619_ & ~new_n43820_;
  assign new_n43822_ = ~pi1149 & ~new_n43821_;
  assign new_n43823_ = pi1148 & ~new_n43822_;
  assign new_n43824_ = ~new_n43817_ & new_n43823_;
  assign new_n43825_ = pi1091 & new_n43824_;
  assign new_n43826_ = pi1150 & ~new_n42389_;
  assign new_n43827_ = ~pi1149 & ~new_n43826_;
  assign new_n43828_ = ~pi1148 & ~new_n43827_;
  assign new_n43829_ = pi1150 & new_n43628_;
  assign new_n43830_ = ~pi1150 & ~new_n43633_;
  assign new_n43831_ = pi1149 & ~new_n43830_;
  assign new_n43832_ = ~new_n43829_ & new_n43831_;
  assign new_n43833_ = pi1091 & ~new_n43832_;
  assign new_n43834_ = new_n43828_ & new_n43833_;
  assign new_n43835_ = ~pi0283 & ~new_n43834_;
  assign new_n43836_ = ~new_n43825_ & new_n43835_;
  assign new_n43837_ = ~pi0272 & ~new_n43836_;
  assign new_n43838_ = ~new_n43811_ & new_n43837_;
  assign new_n43839_ = pi1150 & new_n43547_;
  assign new_n43840_ = ~pi1150 & new_n43508_;
  assign new_n43841_ = pi1149 & ~new_n43840_;
  assign new_n43842_ = ~new_n43839_ & new_n43841_;
  assign new_n43843_ = pi1150 & new_n43542_;
  assign new_n43844_ = ~pi1150 & new_n43502_;
  assign new_n43845_ = ~pi1149 & ~new_n43844_;
  assign new_n43846_ = ~new_n43843_ & new_n43845_;
  assign new_n43847_ = ~new_n43842_ & ~new_n43846_;
  assign new_n43848_ = pi1148 & ~new_n43847_;
  assign new_n43849_ = pi1150 & new_n43596_;
  assign new_n43850_ = ~pi1150 & ~new_n43604_;
  assign new_n43851_ = ~pi1149 & ~new_n43850_;
  assign new_n43852_ = ~new_n43849_ & new_n43851_;
  assign new_n43853_ = pi1150 & new_n43592_;
  assign new_n43854_ = ~pi1150 & new_n43602_;
  assign new_n43855_ = pi1149 & ~new_n43854_;
  assign new_n43856_ = ~new_n43853_ & new_n43855_;
  assign new_n43857_ = ~new_n43852_ & ~new_n43856_;
  assign new_n43858_ = ~pi1148 & ~new_n43857_;
  assign new_n43859_ = pi0283 & ~new_n43858_;
  assign new_n43860_ = ~new_n43848_ & new_n43859_;
  assign new_n43861_ = pi1091 & ~new_n43628_;
  assign new_n43862_ = pi1150 & ~new_n43861_;
  assign new_n43863_ = ~new_n16479_ & new_n42804_;
  assign new_n43864_ = ~po1038 & new_n41080_;
  assign new_n43865_ = ~new_n43863_ & ~new_n43864_;
  assign new_n43866_ = ~pi1150 & new_n43865_;
  assign new_n43867_ = pi1149 & ~new_n43866_;
  assign new_n43868_ = ~new_n43862_ & new_n43867_;
  assign new_n43869_ = pi1091 & new_n43827_;
  assign new_n43870_ = ~pi1148 & ~new_n43869_;
  assign new_n43871_ = ~new_n43868_ & new_n43870_;
  assign new_n43872_ = pi1149 & ~pi1150;
  assign new_n43873_ = ~new_n43619_ & ~new_n43872_;
  assign new_n43874_ = new_n43616_ & ~new_n43873_;
  assign new_n43875_ = ~new_n43822_ & ~new_n43874_;
  assign new_n43876_ = pi1091 & ~new_n43875_;
  assign new_n43877_ = pi1148 & ~new_n43876_;
  assign new_n43878_ = ~pi0283 & ~new_n43877_;
  assign new_n43879_ = ~new_n43871_ & new_n43878_;
  assign new_n43880_ = pi0272 & ~new_n43879_;
  assign new_n43881_ = ~new_n43860_ & new_n43880_;
  assign new_n43882_ = ~pi0230 & ~new_n43881_;
  assign new_n43883_ = ~new_n43838_ & new_n43882_;
  assign new_n43884_ = pi1149 & ~new_n43628_;
  assign new_n43885_ = ~new_n43816_ & ~new_n43884_;
  assign new_n43886_ = ~new_n43830_ & ~new_n43885_;
  assign new_n43887_ = new_n43828_ & ~new_n43886_;
  assign new_n43888_ = pi0230 & ~new_n43824_;
  assign new_n43889_ = ~new_n43887_ & new_n43888_;
  assign po0429 = ~new_n43883_ & ~new_n43889_;
  assign new_n43891_ = ~pi0273 & ~new_n40894_;
  assign new_n43892_ = ~new_n40867_ & ~new_n43891_;
  assign new_n43893_ = pi0219 & ~new_n43892_;
  assign new_n43894_ = ~pi0273 & ~new_n40876_;
  assign new_n43895_ = new_n40878_ & ~new_n43894_;
  assign new_n43896_ = ~pi0219 & ~new_n43750_;
  assign new_n43897_ = ~new_n43895_ & new_n43896_;
  assign new_n43898_ = ~new_n43893_ & ~new_n43897_;
  assign new_n43899_ = pi0299 & new_n43898_;
  assign new_n43900_ = ~pi0200 & new_n43748_;
  assign new_n43901_ = ~pi0199 & ~new_n43900_;
  assign new_n43902_ = ~new_n43895_ & new_n43901_;
  assign new_n43903_ = pi0199 & ~new_n43892_;
  assign new_n43904_ = ~pi0299 & ~new_n43903_;
  assign new_n43905_ = ~new_n43902_ & new_n43904_;
  assign new_n43906_ = ~new_n43899_ & ~new_n43905_;
  assign new_n43907_ = ~new_n11447_ & ~new_n41034_;
  assign new_n43908_ = pi1091 & ~new_n43907_;
  assign new_n43909_ = new_n43906_ & ~new_n43908_;
  assign new_n43910_ = ~po1038 & ~new_n43909_;
  assign new_n43911_ = pi1091 & new_n42502_;
  assign new_n43912_ = ~new_n43910_ & ~new_n43911_;
  assign new_n43913_ = pi1147 & ~new_n43912_;
  assign new_n43914_ = po1038 & new_n43898_;
  assign new_n43915_ = new_n40343_ & ~new_n43906_;
  assign new_n43916_ = ~pi1148 & ~new_n43915_;
  assign new_n43917_ = pi1091 & new_n38519_;
  assign new_n43918_ = ~new_n43898_ & ~new_n43917_;
  assign new_n43919_ = pi0299 & ~new_n43918_;
  assign new_n43920_ = new_n41076_ & ~new_n43763_;
  assign new_n43921_ = ~new_n43905_ & ~new_n43920_;
  assign new_n43922_ = ~new_n43919_ & new_n43921_;
  assign new_n43923_ = ~po1038 & ~new_n43922_;
  assign new_n43924_ = new_n40080_ & new_n42456_;
  assign new_n43925_ = pi1148 & ~new_n43924_;
  assign new_n43926_ = ~new_n43923_ & new_n43925_;
  assign new_n43927_ = ~new_n43916_ & ~new_n43926_;
  assign new_n43928_ = ~new_n43914_ & ~new_n43927_;
  assign new_n43929_ = ~new_n43913_ & new_n43928_;
  assign new_n43930_ = ~pi0230 & ~new_n43929_;
  assign new_n43931_ = ~pi1146 & new_n10730_;
  assign new_n43932_ = pi1147 & new_n40164_;
  assign new_n43933_ = ~new_n43617_ & ~new_n43932_;
  assign new_n43934_ = ~new_n43931_ & ~new_n43933_;
  assign new_n43935_ = ~pi1146 & new_n10817_;
  assign new_n43936_ = ~pi0199 & pi1147;
  assign new_n43937_ = pi0200 & ~new_n43936_;
  assign new_n43938_ = ~new_n43935_ & ~new_n43937_;
  assign new_n43939_ = new_n16479_ & new_n43938_;
  assign new_n43940_ = pi1148 & ~new_n43939_;
  assign new_n43941_ = ~new_n43934_ & new_n43940_;
  assign new_n43942_ = ~pi0211 & ~new_n40237_;
  assign new_n43943_ = new_n40164_ & ~new_n43942_;
  assign new_n43944_ = new_n43615_ & ~new_n43935_;
  assign new_n43945_ = ~new_n43943_ & ~new_n43944_;
  assign new_n43946_ = pi1147 & ~new_n43945_;
  assign new_n43947_ = pi1146 & ~new_n41427_;
  assign new_n43948_ = ~new_n43819_ & new_n43947_;
  assign new_n43949_ = ~pi1148 & ~new_n43948_;
  assign new_n43950_ = ~new_n43946_ & new_n43949_;
  assign new_n43951_ = pi0230 & ~new_n43950_;
  assign new_n43952_ = ~new_n43941_ & new_n43951_;
  assign po0430 = new_n43930_ | new_n43952_;
  assign new_n43954_ = pi0274 & ~new_n40872_;
  assign new_n43955_ = ~pi0659 & new_n40872_;
  assign new_n43956_ = ~pi1091 & ~new_n43955_;
  assign new_n43957_ = ~new_n43954_ & new_n43956_;
  assign new_n43958_ = ~new_n43151_ & ~new_n43957_;
  assign new_n43959_ = ~pi0211 & ~new_n43958_;
  assign new_n43960_ = ~new_n43194_ & ~new_n43957_;
  assign new_n43961_ = pi0211 & ~new_n43960_;
  assign new_n43962_ = ~pi0219 & ~new_n43961_;
  assign new_n43963_ = ~new_n43959_ & new_n43962_;
  assign new_n43964_ = pi0274 & ~new_n40861_;
  assign new_n43965_ = ~pi0659 & new_n40861_;
  assign new_n43966_ = ~pi1091 & ~new_n43965_;
  assign new_n43967_ = ~new_n43964_ & new_n43966_;
  assign new_n43968_ = pi0219 & ~new_n43752_;
  assign new_n43969_ = ~new_n43967_ & new_n43968_;
  assign new_n43970_ = ~new_n16479_ & ~new_n43969_;
  assign new_n43971_ = ~new_n43963_ & new_n43970_;
  assign new_n43972_ = ~pi0200 & ~new_n43958_;
  assign new_n43973_ = pi0200 & ~new_n43960_;
  assign new_n43974_ = ~pi0199 & ~new_n43973_;
  assign new_n43975_ = ~new_n43972_ & new_n43974_;
  assign new_n43976_ = ~pi0200 & new_n43764_;
  assign new_n43977_ = pi0199 & ~new_n43976_;
  assign new_n43978_ = ~new_n43967_ & new_n43977_;
  assign new_n43979_ = new_n16479_ & ~new_n43978_;
  assign new_n43980_ = ~new_n43975_ & new_n43979_;
  assign new_n43981_ = ~pi0230 & ~new_n43980_;
  assign new_n43982_ = ~new_n43971_ & new_n43981_;
  assign new_n43983_ = ~pi0219 & ~new_n38425_;
  assign new_n43984_ = ~new_n39370_ & new_n43983_;
  assign new_n43985_ = ~new_n40220_ & ~new_n43984_;
  assign new_n43986_ = ~new_n38508_ & ~new_n40223_;
  assign new_n43987_ = ~new_n43984_ & ~new_n43986_;
  assign new_n43988_ = ~new_n38436_ & new_n40331_;
  assign new_n43989_ = new_n40781_ & ~new_n43988_;
  assign new_n43990_ = ~new_n43987_ & ~new_n43989_;
  assign new_n43991_ = ~po1038 & ~new_n43990_;
  assign new_n43992_ = pi0230 & ~new_n43991_;
  assign new_n43993_ = ~new_n43985_ & new_n43992_;
  assign po0431 = ~new_n43982_ & ~new_n43993_;
  assign new_n43995_ = pi1151 & ~new_n43619_;
  assign new_n43996_ = pi1149 & new_n43616_;
  assign new_n43997_ = ~new_n43995_ & new_n43996_;
  assign new_n43998_ = ~pi1149 & new_n43629_;
  assign new_n43999_ = ~new_n43997_ & ~new_n43998_;
  assign new_n44000_ = pi1150 & ~new_n43999_;
  assign new_n44001_ = ~pi1151 & new_n43819_;
  assign new_n44002_ = pi1149 & ~new_n43619_;
  assign new_n44003_ = ~new_n44001_ & new_n44002_;
  assign new_n44004_ = ~pi1149 & pi1151;
  assign new_n44005_ = ~new_n42389_ & new_n44004_;
  assign new_n44006_ = ~pi1150 & ~new_n44005_;
  assign new_n44007_ = ~new_n44003_ & new_n44006_;
  assign new_n44008_ = ~new_n44000_ & ~new_n44007_;
  assign new_n44009_ = pi1091 & ~new_n44008_;
  assign new_n44010_ = ~pi1151 & new_n41609_;
  assign new_n44011_ = ~new_n43865_ & new_n44010_;
  assign new_n44012_ = ~new_n44009_ & ~new_n44011_;
  assign new_n44013_ = pi0275 & ~new_n44012_;
  assign new_n44014_ = ~pi1151 & new_n43633_;
  assign new_n44015_ = pi1150 & ~new_n44014_;
  assign new_n44016_ = ~new_n43629_ & new_n44015_;
  assign new_n44017_ = new_n40748_ & ~new_n42389_;
  assign new_n44018_ = ~pi1149 & ~new_n44017_;
  assign new_n44019_ = ~new_n44016_ & new_n44018_;
  assign new_n44020_ = new_n43619_ & new_n43872_;
  assign new_n44021_ = ~new_n43997_ & ~new_n44020_;
  assign new_n44022_ = ~new_n44019_ & new_n44021_;
  assign new_n44023_ = pi1091 & new_n44022_;
  assign new_n44024_ = ~pi0275 & ~new_n44023_;
  assign new_n44025_ = ~new_n41151_ & ~new_n44024_;
  assign new_n44026_ = ~new_n44013_ & new_n44025_;
  assign new_n44027_ = pi1151 & ~new_n43542_;
  assign new_n44028_ = ~pi1150 & ~new_n43503_;
  assign new_n44029_ = ~new_n44027_ & new_n44028_;
  assign new_n44030_ = ~pi1151 & ~new_n43508_;
  assign new_n44031_ = pi1150 & ~new_n44030_;
  assign new_n44032_ = ~new_n43548_ & new_n44031_;
  assign new_n44033_ = pi0275 & ~new_n44032_;
  assign new_n44034_ = ~new_n44029_ & new_n44033_;
  assign new_n44035_ = ~pi1150 & ~new_n43553_;
  assign new_n44036_ = pi1151 & ~new_n43790_;
  assign new_n44037_ = ~new_n44035_ & new_n44036_;
  assign new_n44038_ = pi1150 & ~new_n43530_;
  assign new_n44039_ = ~pi1151 & ~new_n44038_;
  assign new_n44040_ = ~new_n43795_ & new_n44039_;
  assign new_n44041_ = ~pi0275 & ~new_n44040_;
  assign new_n44042_ = ~new_n44037_ & new_n44041_;
  assign new_n44043_ = pi1149 & ~new_n44042_;
  assign new_n44044_ = ~new_n44034_ & new_n44043_;
  assign new_n44045_ = ~pi1150 & new_n43575_;
  assign new_n44046_ = pi1151 & ~new_n43801_;
  assign new_n44047_ = ~new_n44045_ & new_n44046_;
  assign new_n44048_ = pi1150 & ~new_n43580_;
  assign new_n44049_ = ~pi1151 & ~new_n43805_;
  assign new_n44050_ = ~new_n44048_ & new_n44049_;
  assign new_n44051_ = ~new_n44047_ & ~new_n44050_;
  assign new_n44052_ = ~pi0275 & ~new_n44051_;
  assign new_n44053_ = ~pi1150 & new_n43596_;
  assign new_n44054_ = ~new_n43853_ & ~new_n44053_;
  assign new_n44055_ = pi1151 & ~new_n44054_;
  assign new_n44056_ = pi1150 & new_n43602_;
  assign new_n44057_ = ~new_n43850_ & ~new_n44056_;
  assign new_n44058_ = ~pi1151 & ~new_n44057_;
  assign new_n44059_ = pi0275 & ~new_n44058_;
  assign new_n44060_ = ~new_n44055_ & new_n44059_;
  assign new_n44061_ = ~pi1149 & ~new_n44060_;
  assign new_n44062_ = ~new_n44052_ & new_n44061_;
  assign new_n44063_ = new_n41151_ & ~new_n44062_;
  assign new_n44064_ = ~new_n44044_ & new_n44063_;
  assign new_n44065_ = ~new_n44026_ & ~new_n44064_;
  assign new_n44066_ = ~pi0230 & ~new_n44065_;
  assign new_n44067_ = pi0230 & new_n44022_;
  assign po0432 = new_n44066_ | new_n44067_;
  assign new_n44069_ = ~pi0276 & ~new_n40862_;
  assign new_n44070_ = new_n40864_ & ~new_n44069_;
  assign new_n44071_ = new_n43686_ & ~new_n43750_;
  assign new_n44072_ = pi0199 & ~new_n43900_;
  assign new_n44073_ = new_n16479_ & new_n44072_;
  assign new_n44074_ = ~new_n44071_ & ~new_n44073_;
  assign new_n44075_ = ~new_n44070_ & ~new_n44074_;
  assign new_n44076_ = ~pi0276 & ~new_n40873_;
  assign new_n44077_ = new_n43744_ & ~new_n44076_;
  assign new_n44078_ = ~new_n38419_ & ~new_n40209_;
  assign new_n44079_ = pi1091 & ~new_n44078_;
  assign new_n44080_ = new_n40164_ & ~new_n44079_;
  assign new_n44081_ = pi1145 & new_n41091_;
  assign new_n44082_ = ~new_n43195_ & ~new_n44081_;
  assign new_n44083_ = new_n43615_ & new_n44082_;
  assign new_n44084_ = ~new_n44080_ & ~new_n44083_;
  assign new_n44085_ = ~new_n44077_ & ~new_n44084_;
  assign new_n44086_ = ~pi0230 & ~new_n44085_;
  assign new_n44087_ = ~new_n44075_ & new_n44086_;
  assign new_n44088_ = ~pi0219 & ~new_n44078_;
  assign new_n44089_ = pi1146 & new_n38519_;
  assign new_n44090_ = ~new_n44088_ & ~new_n44089_;
  assign new_n44091_ = ~new_n16479_ & new_n44090_;
  assign new_n44092_ = ~new_n38434_ & new_n41290_;
  assign new_n44093_ = ~new_n40334_ & ~new_n44092_;
  assign new_n44094_ = new_n16479_ & ~new_n44093_;
  assign new_n44095_ = pi0230 & ~new_n44094_;
  assign new_n44096_ = ~new_n44091_ & new_n44095_;
  assign po0433 = new_n44087_ | new_n44096_;
  assign new_n44098_ = pi0277 & ~new_n40872_;
  assign new_n44099_ = ~pi0820 & new_n40872_;
  assign new_n44100_ = ~pi1091 & ~new_n44099_;
  assign new_n44101_ = ~new_n44098_ & new_n44100_;
  assign new_n44102_ = ~new_n43142_ & ~new_n44101_;
  assign new_n44103_ = pi0200 & ~new_n44102_;
  assign new_n44104_ = ~new_n43706_ & ~new_n44101_;
  assign new_n44105_ = ~pi0200 & ~new_n44104_;
  assign new_n44106_ = ~pi0199 & ~new_n44105_;
  assign new_n44107_ = ~new_n44103_ & new_n44106_;
  assign new_n44108_ = pi0277 & ~new_n40861_;
  assign new_n44109_ = ~pi0820 & new_n40861_;
  assign new_n44110_ = ~pi1091 & ~new_n44109_;
  assign new_n44111_ = ~new_n44108_ & new_n44110_;
  assign new_n44112_ = ~pi0200 & new_n43139_;
  assign new_n44113_ = pi0199 & ~new_n44112_;
  assign new_n44114_ = ~new_n44111_ & new_n44113_;
  assign new_n44115_ = new_n16479_ & ~new_n44114_;
  assign new_n44116_ = ~new_n44107_ & new_n44115_;
  assign new_n44117_ = pi0211 & ~new_n44102_;
  assign new_n44118_ = ~pi0211 & ~new_n44104_;
  assign new_n44119_ = ~pi0219 & ~new_n44118_;
  assign new_n44120_ = ~new_n44117_ & new_n44119_;
  assign new_n44121_ = pi0219 & ~new_n43213_;
  assign new_n44122_ = ~new_n43161_ & ~new_n44121_;
  assign new_n44123_ = ~new_n44111_ & ~new_n44122_;
  assign new_n44124_ = ~new_n16479_ & ~new_n44123_;
  assign new_n44125_ = ~new_n44120_ & new_n44124_;
  assign new_n44126_ = ~new_n44116_ & ~new_n44125_;
  assign new_n44127_ = ~pi0230 & ~new_n44126_;
  assign new_n44128_ = new_n38433_ & ~new_n43726_;
  assign new_n44129_ = pi0200 & ~new_n43168_;
  assign new_n44130_ = ~new_n44128_ & ~new_n44129_;
  assign new_n44131_ = new_n16479_ & ~new_n44130_;
  assign new_n44132_ = ~pi0211 & pi1140;
  assign new_n44133_ = pi0211 & pi1141;
  assign new_n44134_ = ~pi0219 & ~new_n44133_;
  assign new_n44135_ = ~new_n44132_ & new_n44134_;
  assign new_n44136_ = ~new_n44121_ & ~new_n44135_;
  assign new_n44137_ = ~new_n16479_ & ~new_n44136_;
  assign new_n44138_ = pi0230 & ~new_n44137_;
  assign new_n44139_ = ~new_n44131_ & new_n44138_;
  assign po0434 = new_n44127_ | new_n44139_;
  assign new_n44141_ = ~pi0976 & new_n40861_;
  assign new_n44142_ = ~pi0278 & ~new_n40861_;
  assign new_n44143_ = ~pi1091 & ~new_n44142_;
  assign new_n44144_ = ~new_n44141_ & new_n44143_;
  assign new_n44145_ = pi0199 & ~new_n44144_;
  assign new_n44146_ = pi1091 & ~pi1132;
  assign new_n44147_ = pi0278 & ~new_n40872_;
  assign new_n44148_ = pi0976 & new_n40872_;
  assign new_n44149_ = ~pi1091 & ~new_n44148_;
  assign new_n44150_ = ~new_n44147_ & new_n44149_;
  assign new_n44151_ = ~new_n44146_ & ~new_n44150_;
  assign new_n44152_ = ~pi0199 & ~new_n44151_;
  assign new_n44153_ = ~new_n44145_ & ~new_n44152_;
  assign new_n44154_ = ~pi0200 & ~new_n44153_;
  assign new_n44155_ = pi1091 & ~pi1133;
  assign new_n44156_ = ~new_n44150_ & ~new_n44155_;
  assign new_n44157_ = ~pi0199 & ~new_n44156_;
  assign new_n44158_ = ~new_n44145_ & ~new_n44157_;
  assign new_n44159_ = pi0200 & ~new_n44158_;
  assign new_n44160_ = ~pi0299 & ~new_n44159_;
  assign new_n44161_ = ~new_n44154_ & new_n44160_;
  assign new_n44162_ = pi0219 & ~new_n44144_;
  assign new_n44163_ = pi0211 & ~pi1133;
  assign new_n44164_ = ~pi0211 & ~pi1132;
  assign new_n44165_ = ~new_n44163_ & ~new_n44164_;
  assign new_n44166_ = pi1091 & ~new_n44165_;
  assign new_n44167_ = ~new_n44150_ & ~new_n44166_;
  assign new_n44168_ = ~pi0219 & ~new_n44167_;
  assign new_n44169_ = ~new_n44162_ & ~new_n44168_;
  assign new_n44170_ = pi0299 & new_n44169_;
  assign new_n44171_ = ~new_n44161_ & ~new_n44170_;
  assign new_n44172_ = ~po1038 & ~new_n44171_;
  assign new_n44173_ = po1038 & new_n44169_;
  assign new_n44174_ = ~pi0230 & ~new_n44173_;
  assign new_n44175_ = ~new_n44172_ & new_n44174_;
  assign new_n44176_ = ~pi0199 & pi1132;
  assign new_n44177_ = ~pi0200 & ~new_n44176_;
  assign new_n44178_ = ~pi0199 & pi1133;
  assign new_n44179_ = pi0200 & ~new_n44178_;
  assign new_n44180_ = ~pi0299 & ~new_n44179_;
  assign new_n44181_ = ~new_n44177_ & new_n44180_;
  assign new_n44182_ = new_n38508_ & new_n44165_;
  assign new_n44183_ = ~new_n44181_ & ~new_n44182_;
  assign new_n44184_ = ~po1038 & ~new_n44183_;
  assign new_n44185_ = new_n39405_ & new_n44165_;
  assign new_n44186_ = pi0230 & ~new_n44185_;
  assign new_n44187_ = ~new_n44184_ & new_n44186_;
  assign new_n44188_ = ~new_n44175_ & ~new_n44187_;
  assign new_n44189_ = ~pi1134 & ~new_n44188_;
  assign new_n44190_ = ~pi0219 & ~new_n44165_;
  assign new_n44191_ = ~new_n40081_ & ~new_n44190_;
  assign new_n44192_ = new_n10817_ & ~new_n44176_;
  assign new_n44193_ = new_n44180_ & ~new_n44192_;
  assign new_n44194_ = ~new_n42624_ & ~new_n44182_;
  assign new_n44195_ = ~new_n44193_ & new_n44194_;
  assign new_n44196_ = ~po1038 & ~new_n44195_;
  assign new_n44197_ = pi0230 & ~new_n44196_;
  assign new_n44198_ = ~new_n44191_ & new_n44197_;
  assign new_n44199_ = ~new_n41075_ & new_n44154_;
  assign new_n44200_ = new_n44160_ & ~new_n44199_;
  assign new_n44201_ = new_n13062_ & new_n42610_;
  assign new_n44202_ = ~new_n44170_ & ~new_n44201_;
  assign new_n44203_ = ~new_n44200_ & new_n44202_;
  assign new_n44204_ = ~po1038 & ~new_n44203_;
  assign new_n44205_ = ~new_n43924_ & new_n44174_;
  assign new_n44206_ = ~new_n44204_ & new_n44205_;
  assign new_n44207_ = ~new_n44198_ & ~new_n44206_;
  assign new_n44208_ = pi1134 & ~new_n44207_;
  assign po0435 = ~new_n44189_ & ~new_n44208_;
  assign new_n44210_ = ~pi0958 & new_n40861_;
  assign new_n44211_ = ~pi0279 & ~new_n40861_;
  assign new_n44212_ = ~pi1091 & ~new_n44211_;
  assign new_n44213_ = ~new_n44210_ & new_n44212_;
  assign new_n44214_ = pi1135 & new_n43688_;
  assign new_n44215_ = ~new_n44213_ & ~new_n44214_;
  assign new_n44216_ = pi0199 & ~new_n44215_;
  assign new_n44217_ = pi0279 & ~new_n40872_;
  assign new_n44218_ = pi0958 & new_n40872_;
  assign new_n44219_ = ~pi1091 & ~new_n44218_;
  assign new_n44220_ = ~new_n44217_ & new_n44219_;
  assign new_n44221_ = ~pi1133 & new_n43688_;
  assign new_n44222_ = ~pi0199 & ~new_n44221_;
  assign new_n44223_ = ~new_n44220_ & new_n44222_;
  assign new_n44224_ = ~new_n44216_ & ~new_n44223_;
  assign new_n44225_ = new_n16479_ & ~new_n44224_;
  assign new_n44226_ = ~new_n41091_ & new_n44225_;
  assign new_n44227_ = ~new_n42561_ & ~new_n44155_;
  assign new_n44228_ = ~new_n44220_ & new_n44227_;
  assign new_n44229_ = ~pi0219 & ~new_n44228_;
  assign new_n44230_ = pi1135 & new_n42610_;
  assign new_n44231_ = pi0219 & ~new_n44230_;
  assign new_n44232_ = ~new_n44213_ & new_n44231_;
  assign new_n44233_ = ~new_n16479_ & ~new_n44232_;
  assign new_n44234_ = ~new_n44229_ & new_n44233_;
  assign new_n44235_ = ~pi0230 & ~new_n44234_;
  assign new_n44236_ = ~new_n44226_ & new_n44235_;
  assign new_n44237_ = pi0199 & pi1135;
  assign new_n44238_ = ~new_n44178_ & ~new_n44237_;
  assign new_n44239_ = new_n38548_ & ~new_n44238_;
  assign new_n44240_ = pi1135 & new_n38519_;
  assign new_n44241_ = ~pi0211 & ~pi1133;
  assign new_n44242_ = ~pi0219 & ~new_n44241_;
  assign new_n44243_ = ~pi0211 & new_n44242_;
  assign new_n44244_ = ~new_n44240_ & ~new_n44243_;
  assign new_n44245_ = pi0299 & ~new_n44244_;
  assign new_n44246_ = ~new_n44239_ & ~new_n44245_;
  assign new_n44247_ = ~po1038 & ~new_n44246_;
  assign new_n44248_ = po1038 & ~new_n44244_;
  assign new_n44249_ = pi0230 & ~new_n44248_;
  assign new_n44250_ = ~new_n44247_ & new_n44249_;
  assign new_n44251_ = ~new_n44236_ & ~new_n44250_;
  assign new_n44252_ = ~pi1134 & ~new_n44251_;
  assign new_n44253_ = ~pi1133 & new_n10817_;
  assign new_n44254_ = ~pi0200 & pi1135;
  assign new_n44255_ = pi0199 & ~new_n44254_;
  assign new_n44256_ = ~new_n44253_ & ~new_n44255_;
  assign new_n44257_ = new_n16479_ & ~new_n44256_;
  assign new_n44258_ = ~new_n44240_ & ~new_n44242_;
  assign new_n44259_ = ~new_n16479_ & new_n44258_;
  assign new_n44260_ = ~new_n44257_ & ~new_n44259_;
  assign new_n44261_ = pi0230 & ~new_n44260_;
  assign new_n44262_ = pi1091 & ~new_n44241_;
  assign new_n44263_ = new_n40164_ & new_n44262_;
  assign new_n44264_ = ~new_n44225_ & ~new_n44263_;
  assign new_n44265_ = new_n44235_ & new_n44264_;
  assign new_n44266_ = ~new_n44261_ & ~new_n44265_;
  assign new_n44267_ = pi1134 & ~new_n44266_;
  assign po0436 = ~new_n44252_ & ~new_n44267_;
  assign new_n44269_ = ~pi0211 & pi1135;
  assign new_n44270_ = pi0211 & pi1136;
  assign new_n44271_ = ~new_n44269_ & ~new_n44270_;
  assign new_n44272_ = pi1091 & new_n44271_;
  assign new_n44273_ = pi0914 & new_n40872_;
  assign new_n44274_ = ~pi0280 & ~new_n40872_;
  assign new_n44275_ = ~pi1091 & ~new_n44274_;
  assign new_n44276_ = ~new_n44273_ & new_n44275_;
  assign new_n44277_ = ~new_n44272_ & ~new_n44276_;
  assign new_n44278_ = ~pi0219 & ~new_n44277_;
  assign new_n44279_ = ~pi0211 & pi1137;
  assign new_n44280_ = pi0219 & ~new_n44279_;
  assign new_n44281_ = ~new_n43161_ & ~new_n44280_;
  assign new_n44282_ = pi0280 & ~new_n40861_;
  assign new_n44283_ = ~pi0914 & new_n40861_;
  assign new_n44284_ = ~pi1091 & ~new_n44283_;
  assign new_n44285_ = ~new_n44282_ & new_n44284_;
  assign new_n44286_ = ~new_n44281_ & ~new_n44285_;
  assign new_n44287_ = ~new_n44278_ & ~new_n44286_;
  assign new_n44288_ = ~new_n16479_ & ~new_n44287_;
  assign new_n44289_ = pi0200 & pi1136;
  assign new_n44290_ = pi1091 & ~new_n44254_;
  assign new_n44291_ = ~new_n44289_ & new_n44290_;
  assign new_n44292_ = ~pi0199 & ~new_n44291_;
  assign new_n44293_ = ~new_n44276_ & new_n44292_;
  assign new_n44294_ = pi1137 & new_n43688_;
  assign new_n44295_ = ~new_n44285_ & ~new_n44294_;
  assign new_n44296_ = pi0199 & ~new_n44295_;
  assign new_n44297_ = new_n16479_ & ~new_n44296_;
  assign new_n44298_ = ~new_n44293_ & new_n44297_;
  assign new_n44299_ = ~new_n44288_ & ~new_n44298_;
  assign new_n44300_ = ~pi0230 & ~new_n44299_;
  assign new_n44301_ = ~pi0219 & new_n44271_;
  assign new_n44302_ = ~new_n44280_ & ~new_n44301_;
  assign new_n44303_ = ~new_n16479_ & new_n44302_;
  assign new_n44304_ = pi0200 & ~new_n43654_;
  assign new_n44305_ = pi0199 & pi1137;
  assign new_n44306_ = ~pi0200 & ~new_n43229_;
  assign new_n44307_ = ~new_n44305_ & new_n44306_;
  assign new_n44308_ = ~new_n44304_ & ~new_n44307_;
  assign new_n44309_ = new_n16479_ & new_n44308_;
  assign new_n44310_ = pi0230 & ~new_n44309_;
  assign new_n44311_ = ~new_n44303_ & new_n44310_;
  assign po0437 = ~new_n44300_ & ~new_n44311_;
  assign new_n44313_ = ~pi0199 & pi1138;
  assign new_n44314_ = pi0200 & ~new_n44313_;
  assign new_n44315_ = pi0199 & pi1139;
  assign new_n44316_ = ~pi0200 & ~new_n43652_;
  assign new_n44317_ = ~new_n44315_ & new_n44316_;
  assign new_n44318_ = ~new_n44314_ & ~new_n44317_;
  assign new_n44319_ = new_n16479_ & ~new_n44318_;
  assign new_n44320_ = pi0219 & new_n43701_;
  assign new_n44321_ = pi0211 & pi1138;
  assign new_n44322_ = ~new_n44279_ & ~new_n44321_;
  assign new_n44323_ = ~pi0219 & ~new_n44322_;
  assign new_n44324_ = ~new_n44320_ & ~new_n44323_;
  assign new_n44325_ = ~new_n16479_ & new_n44324_;
  assign new_n44326_ = ~new_n44319_ & ~new_n44325_;
  assign new_n44327_ = pi0230 & ~new_n44326_;
  assign new_n44328_ = pi0281 & ~new_n40872_;
  assign new_n44329_ = ~pi0830 & new_n40872_;
  assign new_n44330_ = ~pi1091 & ~new_n44329_;
  assign new_n44331_ = ~new_n44328_ & new_n44330_;
  assign new_n44332_ = pi1091 & ~new_n44322_;
  assign new_n44333_ = new_n40164_ & ~new_n44332_;
  assign new_n44334_ = pi1138 & new_n41091_;
  assign new_n44335_ = ~new_n44294_ & ~new_n44334_;
  assign new_n44336_ = new_n43615_ & new_n44335_;
  assign new_n44337_ = ~new_n44333_ & ~new_n44336_;
  assign new_n44338_ = ~new_n44331_ & ~new_n44337_;
  assign new_n44339_ = pi0281 & ~new_n40861_;
  assign new_n44340_ = ~pi0830 & new_n40861_;
  assign new_n44341_ = ~pi1091 & ~new_n44340_;
  assign new_n44342_ = ~new_n44339_ & new_n44341_;
  assign new_n44343_ = pi1139 & new_n42610_;
  assign new_n44344_ = new_n43686_ & ~new_n44343_;
  assign new_n44345_ = pi0199 & ~new_n43708_;
  assign new_n44346_ = new_n16479_ & new_n44345_;
  assign new_n44347_ = ~new_n44344_ & ~new_n44346_;
  assign new_n44348_ = ~new_n44342_ & ~new_n44347_;
  assign new_n44349_ = ~new_n44338_ & ~new_n44348_;
  assign new_n44350_ = ~pi0230 & ~new_n44349_;
  assign po0438 = ~new_n44327_ & ~new_n44350_;
  assign new_n44352_ = pi0200 & ~new_n43728_;
  assign new_n44353_ = pi0199 & pi1140;
  assign new_n44354_ = ~pi0200 & ~new_n44313_;
  assign new_n44355_ = ~new_n44353_ & new_n44354_;
  assign new_n44356_ = ~new_n44352_ & ~new_n44355_;
  assign new_n44357_ = new_n16479_ & ~new_n44356_;
  assign new_n44358_ = pi0219 & new_n44132_;
  assign new_n44359_ = pi0211 & pi1139;
  assign new_n44360_ = ~new_n43660_ & ~new_n44359_;
  assign new_n44361_ = ~pi0219 & ~new_n44360_;
  assign new_n44362_ = ~new_n44358_ & ~new_n44361_;
  assign new_n44363_ = ~new_n16479_ & new_n44362_;
  assign new_n44364_ = ~new_n44357_ & ~new_n44363_;
  assign new_n44365_ = pi0230 & ~new_n44364_;
  assign new_n44366_ = pi0282 & ~new_n40872_;
  assign new_n44367_ = ~pi0836 & new_n40872_;
  assign new_n44368_ = ~pi1091 & ~new_n44367_;
  assign new_n44369_ = ~new_n44366_ & new_n44368_;
  assign new_n44370_ = pi1091 & ~new_n44360_;
  assign new_n44371_ = new_n40164_ & ~new_n44370_;
  assign new_n44372_ = pi1139 & new_n41091_;
  assign new_n44373_ = ~new_n43689_ & ~new_n44372_;
  assign new_n44374_ = new_n43615_ & new_n44373_;
  assign new_n44375_ = ~new_n44371_ & ~new_n44374_;
  assign new_n44376_ = ~new_n44369_ & ~new_n44375_;
  assign new_n44377_ = pi0282 & ~new_n40861_;
  assign new_n44378_ = ~pi0836 & new_n40861_;
  assign new_n44379_ = ~pi1091 & ~new_n44378_;
  assign new_n44380_ = ~new_n44377_ & new_n44379_;
  assign new_n44381_ = pi1140 & new_n42610_;
  assign new_n44382_ = new_n43686_ & ~new_n44381_;
  assign new_n44383_ = ~pi0200 & new_n43706_;
  assign new_n44384_ = pi0199 & ~new_n44383_;
  assign new_n44385_ = new_n16479_ & new_n44384_;
  assign new_n44386_ = ~new_n44382_ & ~new_n44385_;
  assign new_n44387_ = ~new_n44380_ & ~new_n44386_;
  assign new_n44388_ = ~new_n44376_ & ~new_n44387_;
  assign new_n44389_ = ~pi0230 & ~new_n44388_;
  assign po0439 = ~new_n44365_ & ~new_n44389_;
  assign new_n44391_ = pi1147 & ~new_n43616_;
  assign new_n44392_ = ~pi1149 & new_n43633_;
  assign new_n44393_ = ~new_n44391_ & new_n44392_;
  assign new_n44394_ = pi1147 & ~new_n43819_;
  assign new_n44395_ = new_n43884_ & ~new_n44394_;
  assign new_n44396_ = pi1148 & ~new_n44395_;
  assign new_n44397_ = ~new_n44393_ & new_n44396_;
  assign new_n44398_ = pi1149 & ~new_n42389_;
  assign new_n44399_ = ~new_n44394_ & ~new_n44398_;
  assign new_n44400_ = ~pi1148 & ~new_n44399_;
  assign new_n44401_ = pi0230 & ~new_n44400_;
  assign new_n44402_ = ~new_n44397_ & new_n44401_;
  assign new_n44403_ = ~pi1147 & ~new_n43580_;
  assign new_n44404_ = pi1147 & new_n43530_;
  assign new_n44405_ = ~pi1149 & ~new_n44404_;
  assign new_n44406_ = ~new_n44403_ & new_n44405_;
  assign new_n44407_ = ~pi1147 & new_n43569_;
  assign new_n44408_ = pi1147 & new_n43560_;
  assign new_n44409_ = pi1149 & ~new_n44408_;
  assign new_n44410_ = ~new_n44407_ & new_n44409_;
  assign new_n44411_ = pi1148 & ~new_n44410_;
  assign new_n44412_ = ~new_n44406_ & new_n44411_;
  assign new_n44413_ = pi1147 & new_n43553_;
  assign new_n44414_ = ~pi1147 & new_n43575_;
  assign new_n44415_ = pi1149 & ~new_n44414_;
  assign new_n44416_ = ~new_n44413_ & new_n44415_;
  assign new_n44417_ = pi1147 & new_n43522_;
  assign new_n44418_ = ~pi1147 & ~new_n43529_;
  assign new_n44419_ = ~pi1149 & ~new_n44418_;
  assign new_n44420_ = ~new_n44417_ & new_n44419_;
  assign new_n44421_ = ~pi1148 & ~new_n44420_;
  assign new_n44422_ = ~new_n44416_ & new_n44421_;
  assign new_n44423_ = ~pi0283 & ~new_n44422_;
  assign new_n44424_ = ~new_n44412_ & new_n44423_;
  assign new_n44425_ = pi1147 & new_n43542_;
  assign new_n44426_ = ~pi1147 & new_n43596_;
  assign new_n44427_ = ~pi1148 & ~new_n44426_;
  assign new_n44428_ = ~new_n44425_ & new_n44427_;
  assign new_n44429_ = ~pi1147 & new_n43592_;
  assign new_n44430_ = pi1147 & new_n43547_;
  assign new_n44431_ = pi1148 & ~new_n44430_;
  assign new_n44432_ = ~new_n44429_ & new_n44431_;
  assign new_n44433_ = pi1149 & ~new_n44432_;
  assign new_n44434_ = ~new_n44428_ & new_n44433_;
  assign new_n44435_ = pi1147 & new_n43502_;
  assign new_n44436_ = ~pi1147 & ~new_n43604_;
  assign new_n44437_ = ~pi1148 & ~new_n44436_;
  assign new_n44438_ = ~new_n44435_ & new_n44437_;
  assign new_n44439_ = ~pi1147 & new_n43602_;
  assign new_n44440_ = pi1147 & new_n43508_;
  assign new_n44441_ = pi1148 & ~new_n44440_;
  assign new_n44442_ = ~new_n44439_ & new_n44441_;
  assign new_n44443_ = ~pi1149 & ~new_n44442_;
  assign new_n44444_ = ~new_n44438_ & new_n44443_;
  assign new_n44445_ = pi0283 & ~new_n44444_;
  assign new_n44446_ = ~new_n44434_ & new_n44445_;
  assign new_n44447_ = ~pi0230 & ~new_n44446_;
  assign new_n44448_ = ~new_n44424_ & new_n44447_;
  assign po0440 = ~new_n44402_ & ~new_n44448_;
  assign new_n44450_ = ~pi0284 & ~new_n42902_;
  assign new_n44451_ = pi1143 & new_n42902_;
  assign new_n44452_ = ~new_n40166_ & new_n44451_;
  assign po0441 = new_n44450_ | new_n44452_;
  assign new_n44454_ = new_n3273_ & ~new_n10418_;
  assign new_n44455_ = ~new_n8057_ & new_n44454_;
  assign new_n44456_ = pi0286 & new_n44455_;
  assign new_n44457_ = pi0288 & pi0289;
  assign new_n44458_ = new_n44456_ & new_n44457_;
  assign new_n44459_ = pi0285 & new_n44454_;
  assign new_n44460_ = ~new_n44458_ & ~new_n44459_;
  assign new_n44461_ = pi0285 & new_n44458_;
  assign new_n44462_ = ~po1038 & ~new_n44461_;
  assign new_n44463_ = ~new_n44460_ & new_n44462_;
  assign new_n44464_ = ~po1038 & new_n44458_;
  assign new_n44465_ = ~pi0286 & new_n8057_;
  assign new_n44466_ = ~pi0288 & new_n44465_;
  assign new_n44467_ = ~pi0289 & new_n44466_;
  assign new_n44468_ = pi0285 & ~new_n44467_;
  assign new_n44469_ = ~new_n44464_ & new_n44468_;
  assign new_n44470_ = ~new_n44463_ & ~new_n44469_;
  assign po0442 = ~pi0793 & ~new_n44470_;
  assign new_n44472_ = ~pi0286 & ~new_n44455_;
  assign new_n44473_ = pi0288 & ~new_n44456_;
  assign new_n44474_ = ~new_n44472_ & new_n44473_;
  assign new_n44475_ = ~pi0288 & ~new_n7732_;
  assign new_n44476_ = new_n8057_ & ~new_n44454_;
  assign new_n44477_ = pi0286 & ~new_n44476_;
  assign new_n44478_ = ~new_n44454_ & new_n44465_;
  assign new_n44479_ = ~new_n44477_ & ~new_n44478_;
  assign new_n44480_ = new_n44475_ & ~new_n44479_;
  assign new_n44481_ = ~po1038 & ~new_n44480_;
  assign new_n44482_ = ~new_n44474_ & new_n44481_;
  assign new_n44483_ = new_n8057_ & new_n44475_;
  assign new_n44484_ = ~pi0286 & new_n44483_;
  assign new_n44485_ = pi0286 & ~new_n44483_;
  assign new_n44486_ = po1038 & ~new_n44485_;
  assign new_n44487_ = ~new_n44484_ & new_n44486_;
  assign new_n44488_ = ~pi0793 & ~new_n44487_;
  assign po0443 = ~new_n44482_ & new_n44488_;
  assign new_n44490_ = ~pi0287 & pi0457;
  assign po0444 = ~pi0332 & ~new_n44490_;
  assign new_n44492_ = pi0288 & ~new_n8057_;
  assign new_n44493_ = ~new_n44483_ & ~new_n44492_;
  assign po0637 = ~po1038 & new_n44454_;
  assign new_n44495_ = new_n44493_ & ~po0637;
  assign new_n44496_ = ~new_n44493_ & po0637;
  assign new_n44497_ = ~pi0793 & ~new_n44496_;
  assign po0445 = ~new_n44495_ & new_n44497_;
  assign new_n44499_ = pi0289 & ~new_n44478_;
  assign new_n44500_ = pi0285 & ~pi0289;
  assign new_n44501_ = new_n44478_ & new_n44500_;
  assign new_n44502_ = ~pi0288 & ~new_n44501_;
  assign new_n44503_ = ~new_n44499_ & new_n44502_;
  assign new_n44504_ = ~pi0289 & new_n44473_;
  assign new_n44505_ = ~new_n44458_ & ~new_n44504_;
  assign new_n44506_ = ~new_n44503_ & new_n44505_;
  assign new_n44507_ = ~po1038 & ~new_n44506_;
  assign new_n44508_ = new_n44466_ & new_n44500_;
  assign new_n44509_ = pi0289 & ~new_n44466_;
  assign new_n44510_ = po1038 & ~new_n44509_;
  assign new_n44511_ = ~new_n44508_ & new_n44510_;
  assign new_n44512_ = ~pi0793 & ~new_n44511_;
  assign po0446 = ~new_n44507_ & new_n44512_;
  assign new_n44514_ = ~pi0290 & pi0476;
  assign new_n44515_ = ~pi0476 & ~pi1048;
  assign po0447 = ~new_n44514_ & ~new_n44515_;
  assign new_n44517_ = ~pi0291 & pi0476;
  assign new_n44518_ = ~pi0476 & ~pi1049;
  assign po0448 = ~new_n44517_ & ~new_n44518_;
  assign new_n44520_ = ~pi0292 & pi0476;
  assign new_n44521_ = ~pi0476 & ~pi1084;
  assign po0449 = ~new_n44520_ & ~new_n44521_;
  assign new_n44523_ = ~pi0293 & pi0476;
  assign new_n44524_ = ~pi0476 & ~pi1059;
  assign po0450 = ~new_n44523_ & ~new_n44524_;
  assign new_n44526_ = ~pi0294 & pi0476;
  assign new_n44527_ = ~pi0476 & ~pi1072;
  assign po0451 = ~new_n44526_ & ~new_n44527_;
  assign new_n44529_ = ~pi0295 & pi0476;
  assign new_n44530_ = ~pi0476 & ~pi1053;
  assign po0452 = ~new_n44529_ & ~new_n44530_;
  assign new_n44532_ = ~pi0296 & pi0476;
  assign new_n44533_ = ~pi0476 & ~pi1037;
  assign po0453 = ~new_n44532_ & ~new_n44533_;
  assign new_n44535_ = ~pi0297 & pi0476;
  assign new_n44536_ = ~pi0476 & ~pi1044;
  assign po0454 = ~new_n44535_ & ~new_n44536_;
  assign new_n44538_ = ~pi0478 & pi1044;
  assign new_n44539_ = pi0298 & pi0478;
  assign po0455 = new_n44538_ | new_n44539_;
  assign new_n44541_ = pi0054 & new_n3100_;
  assign new_n44542_ = ~pi0054 & new_n13152_;
  assign new_n44543_ = new_n13411_ & new_n44542_;
  assign new_n44544_ = ~new_n44541_ & ~new_n44543_;
  assign new_n44545_ = new_n3247_ & new_n8880_;
  assign new_n44546_ = ~new_n44544_ & new_n44545_;
  assign new_n44547_ = ~pi0039 & ~new_n44546_;
  assign po0456 = ~new_n11269_ & ~new_n44547_;
  assign new_n44549_ = pi0057 & ~pi0059;
  assign new_n44550_ = new_n10142_ & new_n44549_;
  assign new_n44551_ = ~pi0312 & new_n44550_;
  assign new_n44552_ = pi0300 & ~new_n44551_;
  assign new_n44553_ = ~pi0300 & new_n44551_;
  assign new_n44554_ = ~pi0055 & ~new_n44553_;
  assign po0457 = new_n44552_ | ~new_n44554_;
  assign new_n44556_ = ~pi0301 & new_n44554_;
  assign new_n44557_ = ~pi0055 & pi0301;
  assign new_n44558_ = new_n44553_ & new_n44557_;
  assign po0458 = new_n44556_ | new_n44558_;
  assign new_n44560_ = new_n5798_ & ~po1038;
  assign new_n44561_ = new_n5809_ & ~new_n16479_;
  assign new_n44562_ = ~new_n44560_ & ~new_n44561_;
  assign new_n44563_ = ~pi1148 & new_n44562_;
  assign new_n44564_ = ~pi0222 & ~pi0223;
  assign new_n44565_ = pi0937 & ~new_n44564_;
  assign new_n44566_ = pi0273 & new_n3313_;
  assign new_n44567_ = ~new_n44565_ & ~new_n44566_;
  assign new_n44568_ = new_n44560_ & new_n44567_;
  assign new_n44569_ = new_n3468_ & ~new_n16479_;
  assign new_n44570_ = ~new_n44568_ & ~new_n44569_;
  assign new_n44571_ = pi0237 & ~new_n44570_;
  assign new_n44572_ = ~new_n3057_ & new_n44568_;
  assign new_n44573_ = ~pi0215 & new_n3329_;
  assign new_n44574_ = ~pi0273 & new_n44573_;
  assign new_n44575_ = pi0833 & new_n8075_;
  assign new_n44576_ = ~pi0937 & new_n44575_;
  assign new_n44577_ = ~new_n44574_ & ~new_n44576_;
  assign new_n44578_ = ~new_n16479_ & ~new_n44577_;
  assign new_n44579_ = ~new_n44572_ & ~new_n44578_;
  assign new_n44580_ = ~new_n44571_ & new_n44579_;
  assign po0459 = ~new_n44563_ & new_n44580_;
  assign new_n44582_ = ~pi0478 & pi1049;
  assign new_n44583_ = pi0303 & pi0478;
  assign po0460 = new_n44582_ | new_n44583_;
  assign new_n44585_ = ~pi0478 & pi1048;
  assign new_n44586_ = pi0304 & pi0478;
  assign po0461 = new_n44585_ | new_n44586_;
  assign new_n44588_ = ~pi0478 & pi1084;
  assign new_n44589_ = pi0305 & pi0478;
  assign po0462 = new_n44588_ | new_n44589_;
  assign new_n44591_ = ~pi0478 & pi1059;
  assign new_n44592_ = pi0306 & pi0478;
  assign po0463 = new_n44591_ | new_n44592_;
  assign new_n44594_ = ~pi0478 & pi1053;
  assign new_n44595_ = pi0307 & pi0478;
  assign po0464 = new_n44594_ | new_n44595_;
  assign new_n44597_ = ~pi0478 & pi1037;
  assign new_n44598_ = pi0308 & pi0478;
  assign po0465 = new_n44597_ | new_n44598_;
  assign new_n44600_ = ~pi0478 & pi1072;
  assign new_n44601_ = pi0309 & pi0478;
  assign po0466 = new_n44600_ | new_n44601_;
  assign new_n44603_ = pi1147 & new_n44562_;
  assign new_n44604_ = ~new_n3467_ & new_n44561_;
  assign new_n44605_ = pi0934 & ~new_n3141_;
  assign new_n44606_ = pi0271 & new_n3329_;
  assign new_n44607_ = ~new_n44605_ & ~new_n44606_;
  assign new_n44608_ = new_n44604_ & ~new_n44607_;
  assign new_n44609_ = pi0222 & ~pi0934;
  assign new_n44610_ = ~pi0271 & new_n3313_;
  assign new_n44611_ = ~new_n44609_ & ~new_n44610_;
  assign new_n44612_ = new_n44560_ & new_n44611_;
  assign new_n44613_ = ~new_n44569_ & ~new_n44612_;
  assign new_n44614_ = ~new_n44608_ & new_n44613_;
  assign new_n44615_ = ~new_n44603_ & new_n44614_;
  assign new_n44616_ = ~pi0233 & ~new_n44615_;
  assign new_n44617_ = new_n44561_ & new_n44607_;
  assign new_n44618_ = new_n44560_ & ~new_n44611_;
  assign new_n44619_ = new_n3105_ & new_n16479_;
  assign new_n44620_ = pi1147 & ~new_n44619_;
  assign new_n44621_ = ~new_n44618_ & new_n44620_;
  assign new_n44622_ = ~new_n44617_ & new_n44621_;
  assign new_n44623_ = ~new_n3057_ & new_n44560_;
  assign new_n44624_ = ~new_n44604_ & ~new_n44623_;
  assign new_n44625_ = ~pi1147 & ~new_n44624_;
  assign new_n44626_ = ~new_n44614_ & new_n44625_;
  assign new_n44627_ = ~new_n44622_ & ~new_n44626_;
  assign new_n44628_ = pi0233 & ~new_n44627_;
  assign po0467 = new_n44616_ | new_n44628_;
  assign new_n44630_ = ~pi0055 & ~pi0311;
  assign new_n44631_ = ~new_n44558_ & ~new_n44630_;
  assign new_n44632_ = ~pi0311 & new_n44558_;
  assign po0468 = ~new_n44631_ & ~new_n44632_;
  assign new_n44634_ = pi0312 & ~new_n44550_;
  assign new_n44635_ = ~new_n44551_ & ~new_n44634_;
  assign po0469 = ~pi0055 & ~new_n44635_;
  assign new_n44637_ = ~new_n10407_ & ~new_n13446_;
  assign new_n44638_ = po0740 & ~new_n13453_;
  assign new_n44639_ = new_n10166_ & ~new_n44638_;
  assign po0634 = new_n44637_ | ~new_n44639_;
  assign new_n44641_ = ~pi0954 & po0634;
  assign new_n44642_ = pi0313 & pi0954;
  assign po0470 = ~new_n44641_ & ~new_n44642_;
  assign new_n44644_ = new_n6554_ & new_n8880_;
  assign new_n44645_ = new_n14451_ & ~new_n44644_;
  assign new_n44646_ = ~pi0039 & ~new_n14520_;
  assign new_n44647_ = pi0039 & ~new_n15296_;
  assign new_n44648_ = new_n3211_ & ~new_n44647_;
  assign new_n44649_ = ~new_n44646_ & new_n44648_;
  assign new_n44650_ = ~new_n15592_ & ~new_n44649_;
  assign new_n44651_ = new_n3282_ & new_n10163_;
  assign new_n44652_ = ~new_n44650_ & new_n44651_;
  assign new_n44653_ = ~new_n44645_ & ~new_n44652_;
  assign new_n44654_ = new_n14445_ & new_n14446_;
  assign po0471 = ~new_n44653_ & new_n44654_;
  assign new_n44656_ = ~pi0340 & new_n44454_;
  assign new_n44657_ = ~po1038 & new_n44656_;
  assign new_n44658_ = pi0315 & ~new_n44657_;
  assign new_n44659_ = pi1080 & new_n44657_;
  assign po0472 = new_n44658_ | new_n44659_;
  assign new_n44661_ = pi0316 & ~new_n44657_;
  assign new_n44662_ = pi1047 & new_n44657_;
  assign po0473 = new_n44661_ | new_n44662_;
  assign new_n44664_ = ~pi0330 & po0637;
  assign new_n44665_ = pi0317 & ~new_n44664_;
  assign new_n44666_ = pi1078 & new_n44664_;
  assign po0474 = new_n44665_ | new_n44666_;
  assign new_n44668_ = ~pi0341 & new_n44454_;
  assign new_n44669_ = ~po1038 & new_n44668_;
  assign new_n44670_ = pi0318 & ~new_n44669_;
  assign new_n44671_ = pi1074 & new_n44669_;
  assign po0475 = new_n44670_ | new_n44671_;
  assign new_n44673_ = pi0319 & ~new_n44669_;
  assign new_n44674_ = pi1072 & new_n44669_;
  assign po0476 = new_n44673_ | new_n44674_;
  assign new_n44676_ = pi0320 & ~new_n44657_;
  assign new_n44677_ = pi1048 & new_n44657_;
  assign po0477 = new_n44676_ | new_n44677_;
  assign new_n44679_ = pi0321 & ~new_n44657_;
  assign new_n44680_ = pi1058 & new_n44657_;
  assign po0478 = new_n44679_ | new_n44680_;
  assign new_n44682_ = pi0322 & ~new_n44657_;
  assign new_n44683_ = pi1051 & new_n44657_;
  assign po0479 = new_n44682_ | new_n44683_;
  assign new_n44685_ = pi0323 & ~new_n44657_;
  assign new_n44686_ = pi1065 & new_n44657_;
  assign po0480 = new_n44685_ | new_n44686_;
  assign new_n44688_ = pi0324 & ~new_n44669_;
  assign new_n44689_ = pi1086 & new_n44669_;
  assign po0481 = new_n44688_ | new_n44689_;
  assign new_n44691_ = pi0325 & ~new_n44669_;
  assign new_n44692_ = pi1063 & new_n44669_;
  assign po0482 = new_n44691_ | new_n44692_;
  assign new_n44694_ = pi0326 & ~new_n44669_;
  assign new_n44695_ = pi1057 & new_n44669_;
  assign po0483 = new_n44694_ | new_n44695_;
  assign new_n44697_ = pi0327 & ~new_n44657_;
  assign new_n44698_ = pi1040 & new_n44657_;
  assign po0484 = new_n44697_ | new_n44698_;
  assign new_n44700_ = pi0328 & ~new_n44669_;
  assign new_n44701_ = pi1058 & new_n44669_;
  assign po0485 = new_n44700_ | new_n44701_;
  assign new_n44703_ = pi0329 & ~new_n44669_;
  assign new_n44704_ = pi1043 & new_n44669_;
  assign po0486 = new_n44703_ | new_n44704_;
  assign new_n44706_ = pi1092 & ~new_n2797_;
  assign new_n44707_ = po1038 & new_n44706_;
  assign new_n44708_ = ~pi0330 & new_n44707_;
  assign new_n44709_ = ~po1038 & new_n44706_;
  assign new_n44710_ = ~pi0330 & ~new_n44454_;
  assign new_n44711_ = ~new_n44656_ & ~new_n44710_;
  assign new_n44712_ = new_n44709_ & ~new_n44711_;
  assign po0487 = new_n44708_ | new_n44712_;
  assign new_n44714_ = ~pi0331 & new_n44707_;
  assign new_n44715_ = ~pi0331 & ~new_n44454_;
  assign new_n44716_ = ~new_n44668_ & ~new_n44715_;
  assign new_n44717_ = new_n44709_ & ~new_n44716_;
  assign po0488 = new_n44714_ | new_n44717_;
  assign new_n44719_ = new_n11002_ & new_n13173_;
  assign new_n44720_ = ~new_n11002_ & ~new_n13103_;
  assign new_n44721_ = new_n7471_ & ~new_n44720_;
  assign new_n44722_ = ~pi0070 & ~new_n44721_;
  assign new_n44723_ = pi0332 & new_n9569_;
  assign new_n44724_ = ~new_n44722_ & new_n44723_;
  assign new_n44725_ = ~new_n44719_ & ~new_n44724_;
  assign new_n44726_ = ~pi0039 & ~new_n44725_;
  assign new_n44727_ = pi0039 & new_n10434_;
  assign new_n44728_ = ~pi0038 & ~new_n44727_;
  assign new_n44729_ = ~new_n44726_ & new_n44728_;
  assign po0489 = new_n38269_ & ~new_n44729_;
  assign new_n44731_ = pi0333 & ~new_n44669_;
  assign new_n44732_ = pi1040 & new_n44669_;
  assign po0490 = new_n44731_ | new_n44732_;
  assign new_n44734_ = pi0334 & ~new_n44669_;
  assign new_n44735_ = pi1065 & new_n44669_;
  assign po0491 = new_n44734_ | new_n44735_;
  assign new_n44737_ = pi0335 & ~new_n44669_;
  assign new_n44738_ = pi1069 & new_n44669_;
  assign po0492 = new_n44737_ | new_n44738_;
  assign new_n44740_ = pi0336 & ~new_n44664_;
  assign new_n44741_ = pi1070 & new_n44664_;
  assign po0493 = new_n44740_ | new_n44741_;
  assign new_n44743_ = pi0337 & ~new_n44664_;
  assign new_n44744_ = pi1044 & new_n44664_;
  assign po0494 = new_n44743_ | new_n44744_;
  assign new_n44746_ = pi0338 & ~new_n44664_;
  assign new_n44747_ = pi1072 & new_n44664_;
  assign po0495 = new_n44746_ | new_n44747_;
  assign new_n44749_ = pi0339 & ~new_n44664_;
  assign new_n44750_ = pi1086 & new_n44664_;
  assign po0496 = new_n44749_ | new_n44750_;
  assign new_n44752_ = pi0340 & new_n44707_;
  assign new_n44753_ = ~pi0331 & new_n44454_;
  assign new_n44754_ = ~pi0340 & ~new_n44454_;
  assign new_n44755_ = new_n44709_ & ~new_n44754_;
  assign new_n44756_ = ~new_n44753_ & new_n44755_;
  assign po0497 = ~new_n44752_ & ~new_n44756_;
  assign new_n44758_ = ~pi0341 & ~po0637;
  assign new_n44759_ = ~new_n44664_ & ~new_n44758_;
  assign po0498 = new_n44706_ & ~new_n44759_;
  assign new_n44761_ = pi0342 & ~new_n44657_;
  assign new_n44762_ = pi1049 & new_n44657_;
  assign po0499 = new_n44761_ | new_n44762_;
  assign new_n44764_ = pi0343 & ~new_n44657_;
  assign new_n44765_ = pi1062 & new_n44657_;
  assign po0500 = new_n44764_ | new_n44765_;
  assign new_n44767_ = pi0344 & ~new_n44657_;
  assign new_n44768_ = pi1069 & new_n44657_;
  assign po0501 = new_n44767_ | new_n44768_;
  assign new_n44770_ = pi0345 & ~new_n44657_;
  assign new_n44771_ = pi1039 & new_n44657_;
  assign po0502 = new_n44770_ | new_n44771_;
  assign new_n44773_ = pi0346 & ~new_n44657_;
  assign new_n44774_ = pi1067 & new_n44657_;
  assign po0503 = new_n44773_ | new_n44774_;
  assign new_n44776_ = pi0347 & ~new_n44657_;
  assign new_n44777_ = pi1055 & new_n44657_;
  assign po0504 = new_n44776_ | new_n44777_;
  assign new_n44779_ = pi0348 & ~new_n44657_;
  assign new_n44780_ = pi1087 & new_n44657_;
  assign po0505 = new_n44779_ | new_n44780_;
  assign new_n44782_ = pi0349 & ~new_n44657_;
  assign new_n44783_ = pi1043 & new_n44657_;
  assign po0506 = new_n44782_ | new_n44783_;
  assign new_n44785_ = pi0350 & ~new_n44657_;
  assign new_n44786_ = pi1035 & new_n44657_;
  assign po0507 = new_n44785_ | new_n44786_;
  assign new_n44788_ = pi0351 & ~new_n44657_;
  assign new_n44789_ = pi1079 & new_n44657_;
  assign po0508 = new_n44788_ | new_n44789_;
  assign new_n44791_ = pi0352 & ~new_n44657_;
  assign new_n44792_ = pi1078 & new_n44657_;
  assign po0509 = new_n44791_ | new_n44792_;
  assign new_n44794_ = pi0353 & ~new_n44657_;
  assign new_n44795_ = pi1063 & new_n44657_;
  assign po0510 = new_n44794_ | new_n44795_;
  assign new_n44797_ = pi0354 & ~new_n44657_;
  assign new_n44798_ = pi1045 & new_n44657_;
  assign po0511 = new_n44797_ | new_n44798_;
  assign new_n44800_ = pi0355 & ~new_n44657_;
  assign new_n44801_ = pi1084 & new_n44657_;
  assign po0512 = new_n44800_ | new_n44801_;
  assign new_n44803_ = pi0356 & ~new_n44657_;
  assign new_n44804_ = pi1081 & new_n44657_;
  assign po0513 = new_n44803_ | new_n44804_;
  assign new_n44806_ = pi0357 & ~new_n44657_;
  assign new_n44807_ = pi1076 & new_n44657_;
  assign po0514 = new_n44806_ | new_n44807_;
  assign new_n44809_ = pi0358 & ~new_n44657_;
  assign new_n44810_ = pi1071 & new_n44657_;
  assign po0515 = new_n44809_ | new_n44810_;
  assign new_n44812_ = pi0359 & ~new_n44657_;
  assign new_n44813_ = pi1068 & new_n44657_;
  assign po0516 = new_n44812_ | new_n44813_;
  assign new_n44815_ = pi0360 & ~new_n44657_;
  assign new_n44816_ = pi1042 & new_n44657_;
  assign po0517 = new_n44815_ | new_n44816_;
  assign new_n44818_ = pi0361 & ~new_n44657_;
  assign new_n44819_ = pi1059 & new_n44657_;
  assign po0518 = new_n44818_ | new_n44819_;
  assign new_n44821_ = pi0362 & ~new_n44657_;
  assign new_n44822_ = pi1070 & new_n44657_;
  assign po0519 = new_n44821_ | new_n44822_;
  assign new_n44824_ = pi0363 & ~new_n44664_;
  assign new_n44825_ = pi1049 & new_n44664_;
  assign po0520 = new_n44824_ | new_n44825_;
  assign new_n44827_ = pi0364 & ~new_n44664_;
  assign new_n44828_ = pi1062 & new_n44664_;
  assign po0521 = new_n44827_ | new_n44828_;
  assign new_n44830_ = pi0365 & ~new_n44664_;
  assign new_n44831_ = pi1065 & new_n44664_;
  assign po0522 = new_n44830_ | new_n44831_;
  assign new_n44833_ = pi0366 & ~new_n44664_;
  assign new_n44834_ = pi1069 & new_n44664_;
  assign po0523 = new_n44833_ | new_n44834_;
  assign new_n44836_ = pi0367 & ~new_n44664_;
  assign new_n44837_ = pi1039 & new_n44664_;
  assign po0524 = new_n44836_ | new_n44837_;
  assign new_n44839_ = pi0368 & ~new_n44664_;
  assign new_n44840_ = pi1067 & new_n44664_;
  assign po0525 = new_n44839_ | new_n44840_;
  assign new_n44842_ = pi0369 & ~new_n44664_;
  assign new_n44843_ = pi1080 & new_n44664_;
  assign po0526 = new_n44842_ | new_n44843_;
  assign new_n44845_ = pi0370 & ~new_n44664_;
  assign new_n44846_ = pi1055 & new_n44664_;
  assign po0527 = new_n44845_ | new_n44846_;
  assign new_n44848_ = pi0371 & ~new_n44664_;
  assign new_n44849_ = pi1051 & new_n44664_;
  assign po0528 = new_n44848_ | new_n44849_;
  assign new_n44851_ = pi0372 & ~new_n44664_;
  assign new_n44852_ = pi1048 & new_n44664_;
  assign po0529 = new_n44851_ | new_n44852_;
  assign new_n44854_ = pi0373 & ~new_n44664_;
  assign new_n44855_ = pi1087 & new_n44664_;
  assign po0530 = new_n44854_ | new_n44855_;
  assign new_n44857_ = pi0374 & ~new_n44664_;
  assign new_n44858_ = pi1035 & new_n44664_;
  assign po0531 = new_n44857_ | new_n44858_;
  assign new_n44860_ = pi0375 & ~new_n44664_;
  assign new_n44861_ = pi1047 & new_n44664_;
  assign po0532 = new_n44860_ | new_n44861_;
  assign new_n44863_ = pi0376 & ~new_n44664_;
  assign new_n44864_ = pi1079 & new_n44664_;
  assign po0533 = new_n44863_ | new_n44864_;
  assign new_n44866_ = pi0377 & ~new_n44664_;
  assign new_n44867_ = pi1074 & new_n44664_;
  assign po0534 = new_n44866_ | new_n44867_;
  assign new_n44869_ = pi0378 & ~new_n44664_;
  assign new_n44870_ = pi1063 & new_n44664_;
  assign po0535 = new_n44869_ | new_n44870_;
  assign new_n44872_ = pi0379 & ~new_n44664_;
  assign new_n44873_ = pi1045 & new_n44664_;
  assign po0536 = new_n44872_ | new_n44873_;
  assign new_n44875_ = pi0380 & ~new_n44664_;
  assign new_n44876_ = pi1084 & new_n44664_;
  assign po0537 = new_n44875_ | new_n44876_;
  assign new_n44878_ = pi0381 & ~new_n44664_;
  assign new_n44879_ = pi1081 & new_n44664_;
  assign po0538 = new_n44878_ | new_n44879_;
  assign new_n44881_ = pi0382 & ~new_n44664_;
  assign new_n44882_ = pi1076 & new_n44664_;
  assign po0539 = new_n44881_ | new_n44882_;
  assign new_n44884_ = pi0383 & ~new_n44664_;
  assign new_n44885_ = pi1071 & new_n44664_;
  assign po0540 = new_n44884_ | new_n44885_;
  assign new_n44887_ = pi0384 & ~new_n44664_;
  assign new_n44888_ = pi1068 & new_n44664_;
  assign po0541 = new_n44887_ | new_n44888_;
  assign new_n44890_ = pi0385 & ~new_n44664_;
  assign new_n44891_ = pi1042 & new_n44664_;
  assign po0542 = new_n44890_ | new_n44891_;
  assign new_n44893_ = pi0386 & ~new_n44664_;
  assign new_n44894_ = pi1059 & new_n44664_;
  assign po0543 = new_n44893_ | new_n44894_;
  assign new_n44896_ = pi0387 & ~new_n44664_;
  assign new_n44897_ = pi1053 & new_n44664_;
  assign po0544 = new_n44896_ | new_n44897_;
  assign new_n44899_ = pi0388 & ~new_n44664_;
  assign new_n44900_ = pi1037 & new_n44664_;
  assign po0545 = new_n44899_ | new_n44900_;
  assign new_n44902_ = pi0389 & ~new_n44664_;
  assign new_n44903_ = pi1036 & new_n44664_;
  assign po0546 = new_n44902_ | new_n44903_;
  assign new_n44905_ = pi0390 & ~new_n44669_;
  assign new_n44906_ = pi1049 & new_n44669_;
  assign po0547 = new_n44905_ | new_n44906_;
  assign new_n44908_ = pi0391 & ~new_n44669_;
  assign new_n44909_ = pi1062 & new_n44669_;
  assign po0548 = new_n44908_ | new_n44909_;
  assign new_n44911_ = pi0392 & ~new_n44669_;
  assign new_n44912_ = pi1039 & new_n44669_;
  assign po0549 = new_n44911_ | new_n44912_;
  assign new_n44914_ = pi0393 & ~new_n44669_;
  assign new_n44915_ = pi1067 & new_n44669_;
  assign po0550 = new_n44914_ | new_n44915_;
  assign new_n44917_ = pi0394 & ~new_n44669_;
  assign new_n44918_ = pi1080 & new_n44669_;
  assign po0551 = new_n44917_ | new_n44918_;
  assign new_n44920_ = pi0395 & ~new_n44669_;
  assign new_n44921_ = pi1055 & new_n44669_;
  assign po0552 = new_n44920_ | new_n44921_;
  assign new_n44923_ = pi0396 & ~new_n44669_;
  assign new_n44924_ = pi1051 & new_n44669_;
  assign po0553 = new_n44923_ | new_n44924_;
  assign new_n44926_ = pi0397 & ~new_n44669_;
  assign new_n44927_ = pi1048 & new_n44669_;
  assign po0554 = new_n44926_ | new_n44927_;
  assign new_n44929_ = pi0398 & ~new_n44669_;
  assign new_n44930_ = pi1087 & new_n44669_;
  assign po0555 = new_n44929_ | new_n44930_;
  assign new_n44932_ = pi0399 & ~new_n44669_;
  assign new_n44933_ = pi1047 & new_n44669_;
  assign po0556 = new_n44932_ | new_n44933_;
  assign new_n44935_ = pi0400 & ~new_n44669_;
  assign new_n44936_ = pi1035 & new_n44669_;
  assign po0557 = new_n44935_ | new_n44936_;
  assign new_n44938_ = pi0401 & ~new_n44669_;
  assign new_n44939_ = pi1079 & new_n44669_;
  assign po0558 = new_n44938_ | new_n44939_;
  assign new_n44941_ = pi0402 & ~new_n44669_;
  assign new_n44942_ = pi1078 & new_n44669_;
  assign po0559 = new_n44941_ | new_n44942_;
  assign new_n44944_ = pi0403 & ~new_n44669_;
  assign new_n44945_ = pi1045 & new_n44669_;
  assign po0560 = new_n44944_ | new_n44945_;
  assign new_n44947_ = pi0404 & ~new_n44669_;
  assign new_n44948_ = pi1084 & new_n44669_;
  assign po0561 = new_n44947_ | new_n44948_;
  assign new_n44950_ = pi0405 & ~new_n44669_;
  assign new_n44951_ = pi1081 & new_n44669_;
  assign po0562 = new_n44950_ | new_n44951_;
  assign new_n44953_ = pi0406 & ~new_n44669_;
  assign new_n44954_ = pi1076 & new_n44669_;
  assign po0563 = new_n44953_ | new_n44954_;
  assign new_n44956_ = pi0407 & ~new_n44669_;
  assign new_n44957_ = pi1071 & new_n44669_;
  assign po0564 = new_n44956_ | new_n44957_;
  assign new_n44959_ = pi0408 & ~new_n44669_;
  assign new_n44960_ = pi1068 & new_n44669_;
  assign po0565 = new_n44959_ | new_n44960_;
  assign new_n44962_ = pi0409 & ~new_n44669_;
  assign new_n44963_ = pi1042 & new_n44669_;
  assign po0566 = new_n44962_ | new_n44963_;
  assign new_n44965_ = pi0410 & ~new_n44669_;
  assign new_n44966_ = pi1059 & new_n44669_;
  assign po0567 = new_n44965_ | new_n44966_;
  assign new_n44968_ = pi0411 & ~new_n44669_;
  assign new_n44969_ = pi1053 & new_n44669_;
  assign po0568 = new_n44968_ | new_n44969_;
  assign new_n44971_ = pi0412 & ~new_n44669_;
  assign new_n44972_ = pi1037 & new_n44669_;
  assign po0569 = new_n44971_ | new_n44972_;
  assign new_n44974_ = pi0413 & ~new_n44669_;
  assign new_n44975_ = pi1036 & new_n44669_;
  assign po0570 = new_n44974_ | new_n44975_;
  assign new_n44977_ = ~po1038 & new_n44753_;
  assign new_n44978_ = pi0414 & ~new_n44977_;
  assign new_n44979_ = pi1049 & new_n44977_;
  assign po0571 = new_n44978_ | new_n44979_;
  assign new_n44981_ = pi0415 & ~new_n44977_;
  assign new_n44982_ = pi1062 & new_n44977_;
  assign po0572 = new_n44981_ | new_n44982_;
  assign new_n44984_ = pi0416 & ~new_n44977_;
  assign new_n44985_ = pi1069 & new_n44977_;
  assign po0573 = new_n44984_ | new_n44985_;
  assign new_n44987_ = pi0417 & ~new_n44977_;
  assign new_n44988_ = pi1039 & new_n44977_;
  assign po0574 = new_n44987_ | new_n44988_;
  assign new_n44990_ = pi0418 & ~new_n44977_;
  assign new_n44991_ = pi1067 & new_n44977_;
  assign po0575 = new_n44990_ | new_n44991_;
  assign new_n44993_ = pi0419 & ~new_n44977_;
  assign new_n44994_ = pi1080 & new_n44977_;
  assign po0576 = new_n44993_ | new_n44994_;
  assign new_n44996_ = pi0420 & ~new_n44977_;
  assign new_n44997_ = pi1055 & new_n44977_;
  assign po0577 = new_n44996_ | new_n44997_;
  assign new_n44999_ = pi0421 & ~new_n44977_;
  assign new_n45000_ = pi1051 & new_n44977_;
  assign po0578 = new_n44999_ | new_n45000_;
  assign new_n45002_ = pi0422 & ~new_n44977_;
  assign new_n45003_ = pi1048 & new_n44977_;
  assign po0579 = new_n45002_ | new_n45003_;
  assign new_n45005_ = pi0423 & ~new_n44977_;
  assign new_n45006_ = pi1087 & new_n44977_;
  assign po0580 = new_n45005_ | new_n45006_;
  assign new_n45008_ = pi0424 & ~new_n44977_;
  assign new_n45009_ = pi1047 & new_n44977_;
  assign po0581 = new_n45008_ | new_n45009_;
  assign new_n45011_ = pi0425 & ~new_n44977_;
  assign new_n45012_ = pi1035 & new_n44977_;
  assign po0582 = new_n45011_ | new_n45012_;
  assign new_n45014_ = pi0426 & ~new_n44977_;
  assign new_n45015_ = pi1079 & new_n44977_;
  assign po0583 = new_n45014_ | new_n45015_;
  assign new_n45017_ = pi0427 & ~new_n44977_;
  assign new_n45018_ = pi1078 & new_n44977_;
  assign po0584 = new_n45017_ | new_n45018_;
  assign new_n45020_ = pi0428 & ~new_n44977_;
  assign new_n45021_ = pi1045 & new_n44977_;
  assign po0585 = new_n45020_ | new_n45021_;
  assign new_n45023_ = pi0429 & ~new_n44977_;
  assign new_n45024_ = pi1084 & new_n44977_;
  assign po0586 = new_n45023_ | new_n45024_;
  assign new_n45026_ = pi0430 & ~new_n44977_;
  assign new_n45027_ = pi1076 & new_n44977_;
  assign po0587 = new_n45026_ | new_n45027_;
  assign new_n45029_ = pi0431 & ~new_n44977_;
  assign new_n45030_ = pi1071 & new_n44977_;
  assign po0588 = new_n45029_ | new_n45030_;
  assign new_n45032_ = pi0432 & ~new_n44977_;
  assign new_n45033_ = pi1068 & new_n44977_;
  assign po0589 = new_n45032_ | new_n45033_;
  assign new_n45035_ = pi0433 & ~new_n44977_;
  assign new_n45036_ = pi1042 & new_n44977_;
  assign po0590 = new_n45035_ | new_n45036_;
  assign new_n45038_ = pi0434 & ~new_n44977_;
  assign new_n45039_ = pi1059 & new_n44977_;
  assign po0591 = new_n45038_ | new_n45039_;
  assign new_n45041_ = pi0435 & ~new_n44977_;
  assign new_n45042_ = pi1053 & new_n44977_;
  assign po0592 = new_n45041_ | new_n45042_;
  assign new_n45044_ = pi0436 & ~new_n44977_;
  assign new_n45045_ = pi1037 & new_n44977_;
  assign po0593 = new_n45044_ | new_n45045_;
  assign new_n45047_ = pi0437 & ~new_n44977_;
  assign new_n45048_ = pi1070 & new_n44977_;
  assign po0594 = new_n45047_ | new_n45048_;
  assign new_n45050_ = pi0438 & ~new_n44977_;
  assign new_n45051_ = pi1036 & new_n44977_;
  assign po0595 = new_n45050_ | new_n45051_;
  assign new_n45053_ = pi0439 & ~new_n44664_;
  assign new_n45054_ = pi1057 & new_n44664_;
  assign po0596 = new_n45053_ | new_n45054_;
  assign new_n45056_ = pi0440 & ~new_n44664_;
  assign new_n45057_ = pi1043 & new_n44664_;
  assign po0597 = new_n45056_ | new_n45057_;
  assign new_n45059_ = pi0441 & ~new_n44657_;
  assign new_n45060_ = pi1044 & new_n44657_;
  assign po0598 = new_n45059_ | new_n45060_;
  assign new_n45062_ = pi0442 & ~new_n44664_;
  assign new_n45063_ = pi1058 & new_n44664_;
  assign po0599 = new_n45062_ | new_n45063_;
  assign new_n45065_ = pi0443 & ~new_n44977_;
  assign new_n45066_ = pi1044 & new_n44977_;
  assign po0600 = new_n45065_ | new_n45066_;
  assign new_n45068_ = pi0444 & ~new_n44977_;
  assign new_n45069_ = pi1072 & new_n44977_;
  assign po0601 = new_n45068_ | new_n45069_;
  assign new_n45071_ = pi0445 & ~new_n44977_;
  assign new_n45072_ = pi1081 & new_n44977_;
  assign po0602 = new_n45071_ | new_n45072_;
  assign new_n45074_ = pi0446 & ~new_n44977_;
  assign new_n45075_ = pi1086 & new_n44977_;
  assign po0603 = new_n45074_ | new_n45075_;
  assign new_n45077_ = pi0447 & ~new_n44664_;
  assign new_n45078_ = pi1040 & new_n44664_;
  assign po0604 = new_n45077_ | new_n45078_;
  assign new_n45080_ = pi0448 & ~new_n44977_;
  assign new_n45081_ = pi1074 & new_n44977_;
  assign po0605 = new_n45080_ | new_n45081_;
  assign new_n45083_ = pi0449 & ~new_n44977_;
  assign new_n45084_ = pi1057 & new_n44977_;
  assign po0606 = new_n45083_ | new_n45084_;
  assign new_n45086_ = pi0450 & ~new_n44657_;
  assign new_n45087_ = pi1036 & new_n44657_;
  assign po0607 = new_n45086_ | new_n45087_;
  assign new_n45089_ = pi0451 & ~new_n44977_;
  assign new_n45090_ = pi1063 & new_n44977_;
  assign po0608 = new_n45089_ | new_n45090_;
  assign new_n45092_ = pi0452 & ~new_n44657_;
  assign new_n45093_ = pi1053 & new_n44657_;
  assign po0609 = new_n45092_ | new_n45093_;
  assign new_n45095_ = pi0453 & ~new_n44977_;
  assign new_n45096_ = pi1040 & new_n44977_;
  assign po0610 = new_n45095_ | new_n45096_;
  assign new_n45098_ = pi0454 & ~new_n44977_;
  assign new_n45099_ = pi1043 & new_n44977_;
  assign po0611 = new_n45098_ | new_n45099_;
  assign new_n45101_ = pi0455 & ~new_n44657_;
  assign new_n45102_ = pi1037 & new_n44657_;
  assign po0612 = new_n45101_ | new_n45102_;
  assign new_n45104_ = pi0456 & ~new_n44669_;
  assign new_n45105_ = pi1044 & new_n44669_;
  assign po0613 = new_n45104_ | new_n45105_;
  assign new_n45107_ = pi0594 & pi0600;
  assign new_n45108_ = pi0597 & new_n45107_;
  assign new_n45109_ = pi0601 & new_n45108_;
  assign new_n45110_ = ~pi0804 & ~pi0810;
  assign new_n45111_ = ~pi0595 & new_n45110_;
  assign new_n45112_ = ~pi0599 & pi0810;
  assign new_n45113_ = pi0596 & ~new_n45112_;
  assign new_n45114_ = pi0804 & ~new_n45113_;
  assign new_n45115_ = pi0595 & pi0815;
  assign new_n45116_ = ~new_n45114_ & new_n45115_;
  assign new_n45117_ = ~new_n45111_ & ~new_n45116_;
  assign new_n45118_ = new_n45109_ & ~new_n45117_;
  assign new_n45119_ = ~pi0601 & ~new_n45110_;
  assign new_n45120_ = pi0600 & ~pi0810;
  assign new_n45121_ = pi0804 & ~new_n45120_;
  assign new_n45122_ = ~pi0815 & ~new_n45121_;
  assign new_n45123_ = ~new_n45119_ & new_n45122_;
  assign new_n45124_ = ~new_n45118_ & ~new_n45123_;
  assign new_n45125_ = pi0605 & ~new_n45124_;
  assign new_n45126_ = pi0990 & new_n45107_;
  assign new_n45127_ = ~pi0815 & new_n45121_;
  assign new_n45128_ = new_n45126_ & new_n45127_;
  assign new_n45129_ = ~new_n45125_ & ~new_n45128_;
  assign po0614 = pi0821 & ~new_n45129_;
  assign new_n45131_ = pi0458 & ~new_n44657_;
  assign new_n45132_ = pi1072 & new_n44657_;
  assign po0615 = new_n45131_ | new_n45132_;
  assign new_n45134_ = pi0459 & ~new_n44977_;
  assign new_n45135_ = pi1058 & new_n44977_;
  assign po0616 = new_n45134_ | new_n45135_;
  assign new_n45137_ = pi0460 & ~new_n44657_;
  assign new_n45138_ = pi1086 & new_n44657_;
  assign po0617 = new_n45137_ | new_n45138_;
  assign new_n45140_ = pi0461 & ~new_n44657_;
  assign new_n45141_ = pi1057 & new_n44657_;
  assign po0618 = new_n45140_ | new_n45141_;
  assign new_n45143_ = pi0462 & ~new_n44657_;
  assign new_n45144_ = pi1074 & new_n44657_;
  assign po0619 = new_n45143_ | new_n45144_;
  assign new_n45146_ = pi0463 & ~new_n44669_;
  assign new_n45147_ = pi1070 & new_n44669_;
  assign po0620 = new_n45146_ | new_n45147_;
  assign new_n45149_ = pi0464 & ~new_n44977_;
  assign new_n45150_ = pi1065 & new_n44977_;
  assign po0621 = new_n45149_ | new_n45150_;
  assign new_n45152_ = ~new_n5789_ & ~new_n5798_;
  assign new_n45153_ = pi1157 & new_n45152_;
  assign new_n45154_ = ~new_n11396_ & ~new_n11399_;
  assign new_n45155_ = ~pi0243 & ~new_n45154_;
  assign new_n45156_ = pi0926 & ~new_n45152_;
  assign new_n45157_ = ~new_n45155_ & ~new_n45156_;
  assign new_n45158_ = ~new_n45153_ & new_n45157_;
  assign new_n45159_ = ~pi0299 & new_n44564_;
  assign new_n45160_ = ~new_n11423_ & ~new_n45159_;
  assign new_n45161_ = ~pi0243 & pi1157;
  assign new_n45162_ = ~new_n45160_ & ~new_n45161_;
  assign new_n45163_ = ~new_n45155_ & new_n45162_;
  assign new_n45164_ = ~new_n3490_ & ~new_n11424_;
  assign new_n45165_ = pi0926 & new_n45161_;
  assign new_n45166_ = ~new_n45164_ & new_n45165_;
  assign new_n45167_ = ~new_n45163_ & ~new_n45166_;
  assign new_n45168_ = ~new_n45158_ & new_n45167_;
  assign new_n45169_ = ~po1038 & ~new_n45168_;
  assign new_n45170_ = ~pi0243 & new_n44573_;
  assign new_n45171_ = po1038 & ~new_n45170_;
  assign new_n45172_ = pi0926 & new_n44575_;
  assign new_n45173_ = pi1157 & ~new_n5809_;
  assign new_n45174_ = ~new_n45172_ & ~new_n45173_;
  assign new_n45175_ = new_n45171_ & new_n45174_;
  assign po0622 = ~new_n45169_ & ~new_n45175_;
  assign new_n45177_ = po1038 & ~new_n44573_;
  assign new_n45178_ = ~po1038 & new_n45154_;
  assign new_n45179_ = ~new_n45177_ & ~new_n45178_;
  assign new_n45180_ = ~pi0943 & ~new_n45179_;
  assign new_n45181_ = pi0943 & new_n44624_;
  assign new_n45182_ = ~new_n45180_ & ~new_n45181_;
  assign new_n45183_ = ~pi1151 & ~new_n45182_;
  assign new_n45184_ = ~new_n44569_ & ~new_n44619_;
  assign new_n45185_ = pi0943 & pi1151;
  assign new_n45186_ = ~new_n45184_ & new_n45185_;
  assign new_n45187_ = ~new_n44562_ & new_n45180_;
  assign new_n45188_ = ~po1038 & ~new_n45160_;
  assign new_n45189_ = new_n3141_ & po1038;
  assign new_n45190_ = ~new_n45188_ & ~new_n45189_;
  assign new_n45191_ = ~pi0275 & ~new_n45190_;
  assign new_n45192_ = ~new_n45187_ & ~new_n45191_;
  assign new_n45193_ = ~new_n45186_ & new_n45192_;
  assign po0623 = ~new_n45183_ & new_n45193_;
  assign new_n45195_ = pi0040 & ~pi0287;
  assign new_n45196_ = new_n42344_ & new_n45195_;
  assign new_n45197_ = po0950 & new_n45196_;
  assign new_n45198_ = ~new_n10165_ & ~new_n45197_;
  assign new_n45199_ = ~pi0102 & ~new_n13381_;
  assign new_n45200_ = new_n8899_ & new_n10162_;
  assign new_n45201_ = new_n17083_ & new_n45200_;
  assign new_n45202_ = ~new_n45199_ & new_n45201_;
  assign new_n45203_ = new_n17081_ & new_n45202_;
  assign new_n45204_ = new_n45196_ & ~new_n45203_;
  assign new_n45205_ = ~new_n45196_ & new_n45203_;
  assign new_n45206_ = ~new_n45204_ & ~new_n45205_;
  assign new_n45207_ = ~new_n6277_ & ~new_n45206_;
  assign new_n45208_ = new_n6277_ & new_n45203_;
  assign new_n45209_ = ~new_n45207_ & ~new_n45208_;
  assign new_n45210_ = ~new_n7574_ & ~new_n45209_;
  assign new_n45211_ = new_n7574_ & ~new_n45206_;
  assign new_n45212_ = pi1091 & ~new_n45211_;
  assign new_n45213_ = ~new_n45210_ & new_n45212_;
  assign new_n45214_ = ~new_n7511_ & ~new_n45206_;
  assign new_n45215_ = new_n7511_ & new_n45203_;
  assign new_n45216_ = ~new_n45214_ & ~new_n45215_;
  assign new_n45217_ = pi1093 & ~new_n45216_;
  assign new_n45218_ = ~pi1093 & ~new_n45209_;
  assign new_n45219_ = ~pi1091 & ~new_n45218_;
  assign new_n45220_ = ~new_n45217_ & new_n45219_;
  assign new_n45221_ = ~new_n45213_ & ~new_n45220_;
  assign new_n45222_ = new_n3227_ & new_n44644_;
  assign new_n45223_ = ~new_n45221_ & new_n45222_;
  assign po0624 = ~new_n45198_ & ~new_n45223_;
  assign new_n45225_ = new_n10200_ & new_n11337_;
  assign new_n45226_ = pi0038 & ~pi0039;
  assign new_n45227_ = new_n10197_ & new_n45226_;
  assign new_n45228_ = new_n8962_ & new_n45227_;
  assign new_n45229_ = pi0468 & ~new_n45228_;
  assign po0625 = new_n45225_ | new_n45229_;
  assign new_n45231_ = pi1156 & new_n45152_;
  assign new_n45232_ = ~pi0263 & ~new_n45154_;
  assign new_n45233_ = pi0942 & ~new_n45152_;
  assign new_n45234_ = ~new_n45232_ & ~new_n45233_;
  assign new_n45235_ = ~new_n45231_ & new_n45234_;
  assign new_n45236_ = ~pi0263 & pi1156;
  assign new_n45237_ = ~new_n45160_ & ~new_n45236_;
  assign new_n45238_ = ~new_n45232_ & new_n45237_;
  assign new_n45239_ = pi0942 & new_n45236_;
  assign new_n45240_ = ~new_n45164_ & new_n45239_;
  assign new_n45241_ = ~new_n45238_ & ~new_n45240_;
  assign new_n45242_ = ~new_n45235_ & new_n45241_;
  assign new_n45243_ = ~po1038 & ~new_n45242_;
  assign new_n45244_ = ~pi0263 & new_n44573_;
  assign new_n45245_ = po1038 & ~new_n45244_;
  assign new_n45246_ = pi1156 & ~new_n5809_;
  assign new_n45247_ = pi0942 & new_n44575_;
  assign new_n45248_ = ~new_n45246_ & ~new_n45247_;
  assign new_n45249_ = new_n45245_ & new_n45248_;
  assign po0626 = ~new_n45243_ & ~new_n45249_;
  assign new_n45251_ = pi1155 & new_n45152_;
  assign new_n45252_ = pi0267 & ~new_n45154_;
  assign new_n45253_ = pi0925 & ~new_n45152_;
  assign new_n45254_ = ~new_n45252_ & ~new_n45253_;
  assign new_n45255_ = ~new_n45251_ & new_n45254_;
  assign new_n45256_ = pi0267 & pi1155;
  assign new_n45257_ = ~new_n45160_ & ~new_n45256_;
  assign new_n45258_ = ~new_n45252_ & new_n45257_;
  assign new_n45259_ = pi0925 & new_n45256_;
  assign new_n45260_ = ~new_n45164_ & new_n45259_;
  assign new_n45261_ = ~new_n45258_ & ~new_n45260_;
  assign new_n45262_ = ~new_n45255_ & new_n45261_;
  assign new_n45263_ = ~po1038 & ~new_n45262_;
  assign new_n45264_ = pi0267 & new_n44573_;
  assign new_n45265_ = po1038 & ~new_n45264_;
  assign new_n45266_ = pi1155 & ~new_n5809_;
  assign new_n45267_ = pi0925 & new_n44575_;
  assign new_n45268_ = ~new_n45266_ & ~new_n45267_;
  assign new_n45269_ = new_n45265_ & new_n45268_;
  assign po0627 = ~new_n45263_ & ~new_n45269_;
  assign new_n45271_ = pi1153 & new_n45152_;
  assign new_n45272_ = pi0253 & ~new_n45154_;
  assign new_n45273_ = pi0941 & ~new_n45152_;
  assign new_n45274_ = ~new_n45272_ & ~new_n45273_;
  assign new_n45275_ = ~new_n45271_ & new_n45274_;
  assign new_n45276_ = pi0253 & pi1153;
  assign new_n45277_ = ~new_n45160_ & ~new_n45276_;
  assign new_n45278_ = ~new_n45272_ & new_n45277_;
  assign new_n45279_ = pi0941 & new_n45276_;
  assign new_n45280_ = ~new_n45164_ & new_n45279_;
  assign new_n45281_ = ~new_n45278_ & ~new_n45280_;
  assign new_n45282_ = ~new_n45275_ & new_n45281_;
  assign new_n45283_ = ~po1038 & ~new_n45282_;
  assign new_n45284_ = pi0253 & new_n44573_;
  assign new_n45285_ = po1038 & ~new_n45284_;
  assign new_n45286_ = pi1153 & ~new_n5809_;
  assign new_n45287_ = pi0941 & new_n44575_;
  assign new_n45288_ = ~new_n45286_ & ~new_n45287_;
  assign new_n45289_ = new_n45285_ & new_n45288_;
  assign po0628 = ~new_n45283_ & ~new_n45289_;
  assign new_n45291_ = pi1154 & new_n45152_;
  assign new_n45292_ = pi0254 & ~new_n45154_;
  assign new_n45293_ = pi0923 & ~new_n45152_;
  assign new_n45294_ = ~new_n45292_ & ~new_n45293_;
  assign new_n45295_ = ~new_n45291_ & new_n45294_;
  assign new_n45296_ = pi0254 & pi1154;
  assign new_n45297_ = ~new_n45160_ & ~new_n45296_;
  assign new_n45298_ = ~new_n45292_ & new_n45297_;
  assign new_n45299_ = pi0923 & new_n45296_;
  assign new_n45300_ = ~new_n45164_ & new_n45299_;
  assign new_n45301_ = ~new_n45298_ & ~new_n45300_;
  assign new_n45302_ = ~new_n45295_ & new_n45301_;
  assign new_n45303_ = ~po1038 & ~new_n45302_;
  assign new_n45304_ = pi0254 & new_n44573_;
  assign new_n45305_ = po1038 & ~new_n45304_;
  assign new_n45306_ = pi1154 & ~new_n5809_;
  assign new_n45307_ = pi0923 & new_n44575_;
  assign new_n45308_ = ~new_n45306_ & ~new_n45307_;
  assign new_n45309_ = new_n45305_ & new_n45308_;
  assign po0629 = ~new_n45303_ & ~new_n45309_;
  assign new_n45311_ = ~pi0922 & ~new_n45179_;
  assign new_n45312_ = pi0922 & new_n44624_;
  assign new_n45313_ = ~new_n45311_ & ~new_n45312_;
  assign new_n45314_ = ~pi1152 & ~new_n45313_;
  assign new_n45315_ = pi0922 & pi1152;
  assign new_n45316_ = ~new_n45184_ & new_n45315_;
  assign new_n45317_ = ~new_n44562_ & new_n45311_;
  assign new_n45318_ = ~pi0268 & ~new_n45190_;
  assign new_n45319_ = ~new_n45317_ & ~new_n45318_;
  assign new_n45320_ = ~new_n45316_ & new_n45319_;
  assign po0630 = ~new_n45314_ & new_n45320_;
  assign new_n45322_ = ~pi0931 & ~new_n45179_;
  assign new_n45323_ = pi0931 & new_n44624_;
  assign new_n45324_ = ~new_n45322_ & ~new_n45323_;
  assign new_n45325_ = ~pi1150 & ~new_n45324_;
  assign new_n45326_ = pi0931 & pi1150;
  assign new_n45327_ = ~new_n45184_ & new_n45326_;
  assign new_n45328_ = ~new_n44562_ & new_n45322_;
  assign new_n45329_ = ~pi0272 & ~new_n45190_;
  assign new_n45330_ = ~new_n45328_ & ~new_n45329_;
  assign new_n45331_ = ~new_n45327_ & new_n45330_;
  assign po0631 = ~new_n45325_ & new_n45331_;
  assign new_n45333_ = ~pi0936 & ~new_n45179_;
  assign new_n45334_ = pi0936 & new_n44624_;
  assign new_n45335_ = ~new_n45333_ & ~new_n45334_;
  assign new_n45336_ = ~pi1149 & ~new_n45335_;
  assign new_n45337_ = pi0936 & pi1149;
  assign new_n45338_ = ~new_n45184_ & new_n45337_;
  assign new_n45339_ = ~new_n44562_ & new_n45333_;
  assign new_n45340_ = ~pi0283 & ~new_n45190_;
  assign new_n45341_ = ~new_n45339_ & ~new_n45340_;
  assign new_n45342_ = ~new_n45338_ & new_n45341_;
  assign po0632 = ~new_n45336_ & new_n45342_;
  assign new_n45344_ = pi0071 & new_n43632_;
  assign new_n45345_ = pi0071 & ~new_n11448_;
  assign new_n45346_ = new_n11448_ & new_n13048_;
  assign new_n45347_ = new_n10151_ & ~new_n11448_;
  assign new_n45348_ = new_n10147_ & new_n45347_;
  assign new_n45349_ = ~new_n45346_ & ~new_n45348_;
  assign new_n45350_ = new_n3273_ & new_n10162_;
  assign new_n45351_ = ~new_n45349_ & new_n45350_;
  assign new_n45352_ = new_n13056_ & new_n45351_;
  assign new_n45353_ = ~new_n45345_ & ~new_n45352_;
  assign new_n45354_ = ~po1038 & ~new_n45353_;
  assign po0633 = new_n45344_ | new_n45354_;
  assign po0635 = pi0071 & ~new_n43819_;
  assign new_n45357_ = pi0481 & ~new_n34775_;
  assign new_n45358_ = pi0248 & new_n34775_;
  assign po0638 = new_n45357_ | new_n45358_;
  assign new_n45360_ = pi0482 & ~new_n34791_;
  assign new_n45361_ = pi0249 & new_n34791_;
  assign po0639 = new_n45360_ | new_n45361_;
  assign new_n45363_ = pi0483 & ~new_n34915_;
  assign new_n45364_ = pi0242 & new_n34915_;
  assign po0640 = new_n45363_ | new_n45364_;
  assign new_n45366_ = pi0484 & ~new_n34915_;
  assign new_n45367_ = pi0249 & new_n34915_;
  assign po0641 = new_n45366_ | new_n45367_;
  assign new_n45369_ = pi0485 & ~new_n36111_;
  assign new_n45370_ = pi0234 & new_n36111_;
  assign po0642 = new_n45369_ | new_n45370_;
  assign new_n45372_ = pi0486 & ~new_n36111_;
  assign new_n45373_ = pi0244 & new_n36111_;
  assign po0643 = new_n45372_ | new_n45373_;
  assign new_n45375_ = pi0487 & ~new_n34775_;
  assign new_n45376_ = pi0246 & new_n34775_;
  assign po0644 = new_n45375_ | new_n45376_;
  assign new_n45378_ = pi0488 & ~new_n34775_;
  assign new_n45379_ = ~pi0239 & new_n34775_;
  assign po0645 = ~new_n45378_ & ~new_n45379_;
  assign new_n45381_ = pi0489 & ~new_n36111_;
  assign new_n45382_ = pi0242 & new_n36111_;
  assign po0646 = new_n45381_ | new_n45382_;
  assign new_n45384_ = pi0490 & ~new_n34915_;
  assign new_n45385_ = pi0241 & new_n34915_;
  assign po0647 = new_n45384_ | new_n45385_;
  assign new_n45387_ = pi0491 & ~new_n34915_;
  assign new_n45388_ = pi0238 & new_n34915_;
  assign po0648 = new_n45387_ | new_n45388_;
  assign new_n45390_ = pi0492 & ~new_n34915_;
  assign new_n45391_ = pi0240 & new_n34915_;
  assign po0649 = new_n45390_ | new_n45391_;
  assign new_n45393_ = pi0493 & ~new_n34915_;
  assign new_n45394_ = pi0244 & new_n34915_;
  assign po0650 = new_n45393_ | new_n45394_;
  assign new_n45396_ = pi0494 & ~new_n34915_;
  assign new_n45397_ = ~pi0239 & new_n34915_;
  assign po0651 = ~new_n45396_ & ~new_n45397_;
  assign new_n45399_ = pi0495 & ~new_n34915_;
  assign new_n45400_ = pi0235 & new_n34915_;
  assign po0652 = new_n45399_ | new_n45400_;
  assign new_n45402_ = pi0496 & ~new_n34907_;
  assign new_n45403_ = pi0249 & new_n34907_;
  assign po0653 = new_n45402_ | new_n45403_;
  assign new_n45405_ = pi0497 & ~new_n34907_;
  assign new_n45406_ = ~pi0239 & new_n34907_;
  assign po0654 = ~new_n45405_ & ~new_n45406_;
  assign new_n45408_ = pi0498 & ~new_n34791_;
  assign new_n45409_ = pi0238 & new_n34791_;
  assign po0655 = new_n45408_ | new_n45409_;
  assign new_n45411_ = pi0499 & ~new_n34907_;
  assign new_n45412_ = pi0246 & new_n34907_;
  assign po0656 = new_n45411_ | new_n45412_;
  assign new_n45414_ = pi0500 & ~new_n34907_;
  assign new_n45415_ = pi0241 & new_n34907_;
  assign po0657 = new_n45414_ | new_n45415_;
  assign new_n45417_ = pi0501 & ~new_n34907_;
  assign new_n45418_ = pi0248 & new_n34907_;
  assign po0658 = new_n45417_ | new_n45418_;
  assign new_n45420_ = pi0502 & ~new_n34907_;
  assign new_n45421_ = pi0247 & new_n34907_;
  assign po0659 = new_n45420_ | new_n45421_;
  assign new_n45423_ = pi0503 & ~new_n34907_;
  assign new_n45424_ = pi0245 & new_n34907_;
  assign po0660 = new_n45423_ | new_n45424_;
  assign new_n45426_ = pi0504 & ~new_n34900_;
  assign new_n45427_ = pi0242 & new_n34900_;
  assign po0661 = new_n45426_ | new_n45427_;
  assign new_n45429_ = ~new_n6318_ & new_n16479_;
  assign new_n45430_ = ~new_n34897_ & ~new_n45429_;
  assign new_n45431_ = ~pi0234 & new_n45430_;
  assign new_n45432_ = new_n34907_ & new_n45431_;
  assign new_n45433_ = pi0505 & ~new_n45432_;
  assign new_n45434_ = pi0234 & new_n34899_;
  assign new_n45435_ = ~pi0505 & new_n34778_;
  assign new_n45436_ = new_n45434_ & new_n45435_;
  assign po0662 = new_n45433_ | new_n45436_;
  assign new_n45438_ = pi0506 & ~new_n34900_;
  assign new_n45439_ = pi0241 & new_n34900_;
  assign po0663 = new_n45438_ | new_n45439_;
  assign new_n45441_ = pi0507 & ~new_n34900_;
  assign new_n45442_ = pi0238 & new_n34900_;
  assign po0664 = new_n45441_ | new_n45442_;
  assign new_n45444_ = pi0508 & ~new_n34900_;
  assign new_n45445_ = pi0247 & new_n34900_;
  assign po0665 = new_n45444_ | new_n45445_;
  assign new_n45447_ = pi0509 & ~new_n34900_;
  assign new_n45448_ = pi0245 & new_n34900_;
  assign po0666 = new_n45447_ | new_n45448_;
  assign new_n45450_ = pi0510 & ~new_n34775_;
  assign new_n45451_ = pi0242 & new_n34775_;
  assign po0667 = new_n45450_ | new_n45451_;
  assign new_n45453_ = new_n6616_ & ~po1038;
  assign new_n45454_ = ~new_n34770_ & ~new_n45453_;
  assign new_n45455_ = ~pi0234 & new_n45454_;
  assign new_n45456_ = new_n34775_ & ~new_n45455_;
  assign new_n45457_ = pi0511 & ~new_n34775_;
  assign po0668 = new_n45456_ | new_n45457_;
  assign new_n45459_ = pi0512 & ~new_n34775_;
  assign new_n45460_ = pi0235 & new_n34775_;
  assign po0669 = new_n45459_ | new_n45460_;
  assign new_n45462_ = pi0513 & ~new_n34775_;
  assign new_n45463_ = pi0244 & new_n34775_;
  assign po0670 = new_n45462_ | new_n45463_;
  assign new_n45465_ = pi0514 & ~new_n34775_;
  assign new_n45466_ = pi0245 & new_n34775_;
  assign po0671 = new_n45465_ | new_n45466_;
  assign new_n45468_ = pi0515 & ~new_n34775_;
  assign new_n45469_ = pi0240 & new_n34775_;
  assign po0672 = new_n45468_ | new_n45469_;
  assign new_n45471_ = pi0516 & ~new_n34775_;
  assign new_n45472_ = pi0247 & new_n34775_;
  assign po0673 = new_n45471_ | new_n45472_;
  assign new_n45474_ = pi0517 & ~new_n34775_;
  assign new_n45475_ = pi0238 & new_n34775_;
  assign po0674 = new_n45474_ | new_n45475_;
  assign new_n45477_ = new_n34783_ & new_n45455_;
  assign new_n45478_ = pi0518 & ~new_n45477_;
  assign new_n45479_ = pi0234 & new_n34774_;
  assign new_n45480_ = ~pi0518 & new_n34778_;
  assign new_n45481_ = new_n45479_ & new_n45480_;
  assign po0675 = new_n45478_ | new_n45481_;
  assign new_n45483_ = pi0519 & ~new_n34783_;
  assign new_n45484_ = ~pi0239 & new_n34783_;
  assign po0676 = ~new_n45483_ & ~new_n45484_;
  assign new_n45486_ = pi0520 & ~new_n34783_;
  assign new_n45487_ = pi0246 & new_n34783_;
  assign po0677 = new_n45486_ | new_n45487_;
  assign new_n45489_ = pi0521 & ~new_n34783_;
  assign new_n45490_ = pi0248 & new_n34783_;
  assign po0678 = new_n45489_ | new_n45490_;
  assign new_n45492_ = pi0522 & ~new_n34783_;
  assign new_n45493_ = pi0238 & new_n34783_;
  assign po0679 = new_n45492_ | new_n45493_;
  assign new_n45495_ = new_n36139_ & new_n45455_;
  assign new_n45496_ = pi0523 & ~new_n45495_;
  assign new_n45497_ = ~pi0523 & new_n34910_;
  assign new_n45498_ = new_n45479_ & new_n45497_;
  assign po0680 = new_n45496_ | new_n45498_;
  assign new_n45500_ = pi0524 & ~new_n36139_;
  assign new_n45501_ = ~pi0239 & new_n36139_;
  assign po0681 = ~new_n45500_ & ~new_n45501_;
  assign new_n45503_ = pi0525 & ~new_n36139_;
  assign new_n45504_ = pi0245 & new_n36139_;
  assign po0682 = new_n45503_ | new_n45504_;
  assign new_n45506_ = pi0526 & ~new_n36139_;
  assign new_n45507_ = pi0246 & new_n36139_;
  assign po0683 = new_n45506_ | new_n45507_;
  assign new_n45509_ = pi0527 & ~new_n36139_;
  assign new_n45510_ = pi0247 & new_n36139_;
  assign po0684 = new_n45509_ | new_n45510_;
  assign new_n45512_ = pi0528 & ~new_n36139_;
  assign new_n45513_ = pi0249 & new_n36139_;
  assign po0685 = new_n45512_ | new_n45513_;
  assign new_n45515_ = pi0529 & ~new_n36139_;
  assign new_n45516_ = pi0238 & new_n36139_;
  assign po0686 = new_n45515_ | new_n45516_;
  assign new_n45518_ = pi0530 & ~new_n36139_;
  assign new_n45519_ = pi0240 & new_n36139_;
  assign po0687 = new_n45518_ | new_n45519_;
  assign new_n45521_ = pi0531 & ~new_n34791_;
  assign new_n45522_ = pi0235 & new_n34791_;
  assign po0688 = new_n45521_ | new_n45522_;
  assign new_n45524_ = pi0532 & ~new_n34791_;
  assign new_n45525_ = pi0247 & new_n34791_;
  assign po0689 = new_n45524_ | new_n45525_;
  assign new_n45527_ = pi0533 & ~new_n34900_;
  assign new_n45528_ = pi0235 & new_n34900_;
  assign po0690 = new_n45527_ | new_n45528_;
  assign new_n45530_ = pi0534 & ~new_n34900_;
  assign new_n45531_ = ~pi0239 & new_n34900_;
  assign po0691 = ~new_n45530_ & ~new_n45531_;
  assign new_n45533_ = pi0535 & ~new_n34900_;
  assign new_n45534_ = pi0240 & new_n34900_;
  assign po0692 = new_n45533_ | new_n45534_;
  assign new_n45536_ = pi0536 & ~new_n34900_;
  assign new_n45537_ = pi0246 & new_n34900_;
  assign po0693 = new_n45536_ | new_n45537_;
  assign new_n45539_ = pi0537 & ~new_n34900_;
  assign new_n45540_ = pi0248 & new_n34900_;
  assign po0694 = new_n45539_ | new_n45540_;
  assign new_n45542_ = pi0538 & ~new_n34900_;
  assign new_n45543_ = pi0249 & new_n34900_;
  assign po0695 = new_n45542_ | new_n45543_;
  assign new_n45545_ = pi0539 & ~new_n34907_;
  assign new_n45546_ = pi0242 & new_n34907_;
  assign po0696 = new_n45545_ | new_n45546_;
  assign new_n45548_ = pi0540 & ~new_n34907_;
  assign new_n45549_ = pi0235 & new_n34907_;
  assign po0697 = new_n45548_ | new_n45549_;
  assign new_n45551_ = pi0541 & ~new_n34907_;
  assign new_n45552_ = pi0244 & new_n34907_;
  assign po0698 = new_n45551_ | new_n45552_;
  assign new_n45554_ = pi0542 & ~new_n34907_;
  assign new_n45555_ = pi0240 & new_n34907_;
  assign po0699 = new_n45554_ | new_n45555_;
  assign new_n45557_ = pi0543 & ~new_n34907_;
  assign new_n45558_ = pi0238 & new_n34907_;
  assign po0700 = new_n45557_ | new_n45558_;
  assign new_n45560_ = new_n34915_ & new_n45431_;
  assign new_n45561_ = pi0544 & ~new_n45560_;
  assign new_n45562_ = ~pi0544 & new_n34910_;
  assign new_n45563_ = new_n45434_ & new_n45562_;
  assign po0701 = new_n45561_ | new_n45563_;
  assign new_n45565_ = pi0545 & ~new_n34915_;
  assign new_n45566_ = pi0245 & new_n34915_;
  assign po0702 = new_n45565_ | new_n45566_;
  assign new_n45568_ = pi0546 & ~new_n34915_;
  assign new_n45569_ = pi0246 & new_n34915_;
  assign po0703 = new_n45568_ | new_n45569_;
  assign new_n45571_ = pi0547 & ~new_n34915_;
  assign new_n45572_ = pi0247 & new_n34915_;
  assign po0704 = new_n45571_ | new_n45572_;
  assign new_n45574_ = pi0548 & ~new_n34915_;
  assign new_n45575_ = pi0248 & new_n34915_;
  assign po0705 = new_n45574_ | new_n45575_;
  assign new_n45577_ = pi0549 & ~new_n36111_;
  assign new_n45578_ = pi0235 & new_n36111_;
  assign po0706 = new_n45577_ | new_n45578_;
  assign new_n45580_ = pi0550 & ~new_n36111_;
  assign new_n45581_ = ~pi0239 & new_n36111_;
  assign po0707 = ~new_n45580_ & ~new_n45581_;
  assign new_n45583_ = pi0551 & ~new_n36111_;
  assign new_n45584_ = pi0240 & new_n36111_;
  assign po0708 = new_n45583_ | new_n45584_;
  assign new_n45586_ = pi0552 & ~new_n36111_;
  assign new_n45587_ = pi0247 & new_n36111_;
  assign po0709 = new_n45586_ | new_n45587_;
  assign new_n45589_ = pi0553 & ~new_n36111_;
  assign new_n45590_ = pi0241 & new_n36111_;
  assign po0710 = new_n45589_ | new_n45590_;
  assign new_n45592_ = pi0554 & ~new_n36111_;
  assign new_n45593_ = pi0248 & new_n36111_;
  assign po0711 = new_n45592_ | new_n45593_;
  assign new_n45595_ = pi0555 & ~new_n36111_;
  assign new_n45596_ = pi0249 & new_n36111_;
  assign po0712 = new_n45595_ | new_n45596_;
  assign new_n45598_ = pi0556 & ~new_n34791_;
  assign new_n45599_ = pi0242 & new_n34791_;
  assign po0713 = new_n45598_ | new_n45599_;
  assign new_n45601_ = new_n34900_ & new_n45431_;
  assign new_n45602_ = pi0557 & ~new_n45601_;
  assign new_n45603_ = ~pi0557 & new_n34583_;
  assign new_n45604_ = new_n45434_ & new_n45603_;
  assign po0714 = new_n45602_ | new_n45604_;
  assign new_n45606_ = pi0558 & ~new_n34900_;
  assign new_n45607_ = pi0244 & new_n34900_;
  assign po0715 = new_n45606_ | new_n45607_;
  assign new_n45609_ = pi0559 & ~new_n34775_;
  assign new_n45610_ = pi0241 & new_n34775_;
  assign po0716 = new_n45609_ | new_n45610_;
  assign new_n45612_ = pi0560 & ~new_n34791_;
  assign new_n45613_ = pi0240 & new_n34791_;
  assign po0717 = new_n45612_ | new_n45613_;
  assign new_n45615_ = pi0561 & ~new_n34783_;
  assign new_n45616_ = pi0247 & new_n34783_;
  assign po0718 = new_n45615_ | new_n45616_;
  assign new_n45618_ = pi0562 & ~new_n34791_;
  assign new_n45619_ = pi0241 & new_n34791_;
  assign po0719 = new_n45618_ | new_n45619_;
  assign new_n45621_ = pi0563 & ~new_n36111_;
  assign new_n45622_ = pi0246 & new_n36111_;
  assign po0720 = new_n45621_ | new_n45622_;
  assign new_n45624_ = pi0564 & ~new_n34791_;
  assign new_n45625_ = pi0246 & new_n34791_;
  assign po0721 = new_n45624_ | new_n45625_;
  assign new_n45627_ = pi0565 & ~new_n34791_;
  assign new_n45628_ = pi0248 & new_n34791_;
  assign po0722 = new_n45627_ | new_n45628_;
  assign new_n45630_ = pi0566 & ~new_n34791_;
  assign new_n45631_ = pi0244 & new_n34791_;
  assign po0723 = new_n45630_ | new_n45631_;
  assign new_n45633_ = pi0603 & ~new_n17590_;
  assign new_n45634_ = new_n16869_ & ~new_n20223_;
  assign new_n45635_ = ~new_n20229_ & new_n45634_;
  assign new_n45636_ = new_n45633_ & new_n45635_;
  assign new_n45637_ = ~pi0567 & pi1092;
  assign new_n45638_ = ~pi1093 & new_n45637_;
  assign new_n45639_ = ~pi0789 & ~new_n45638_;
  assign new_n45640_ = ~new_n45636_ & new_n45639_;
  assign new_n45641_ = pi0619 & new_n45636_;
  assign new_n45642_ = ~new_n45638_ & ~new_n45641_;
  assign new_n45643_ = pi1159 & ~new_n45642_;
  assign new_n45644_ = ~pi0619 & new_n45636_;
  assign new_n45645_ = ~new_n45638_ & ~new_n45644_;
  assign new_n45646_ = ~pi1159 & ~new_n45645_;
  assign new_n45647_ = pi0789 & ~new_n45646_;
  assign new_n45648_ = ~new_n45643_ & new_n45647_;
  assign new_n45649_ = ~new_n45640_ & ~new_n45648_;
  assign new_n45650_ = pi0680 & new_n17523_;
  assign new_n45651_ = ~new_n19188_ & new_n45650_;
  assign new_n45652_ = ~new_n45638_ & ~new_n45651_;
  assign new_n45653_ = new_n19280_ & ~new_n45652_;
  assign new_n45654_ = ~new_n17690_ & new_n45648_;
  assign new_n45655_ = new_n45653_ & ~new_n45654_;
  assign new_n45656_ = ~new_n45649_ & ~new_n45655_;
  assign new_n45657_ = new_n17969_ & ~new_n45656_;
  assign new_n45658_ = new_n35259_ & new_n45649_;
  assign new_n45659_ = ~new_n17691_ & new_n45653_;
  assign new_n45660_ = pi0641 & new_n45659_;
  assign new_n45661_ = ~new_n45638_ & ~new_n45660_;
  assign new_n45662_ = new_n17850_ & ~new_n45661_;
  assign new_n45663_ = ~pi0641 & new_n45659_;
  assign new_n45664_ = ~new_n45638_ & ~new_n45663_;
  assign new_n45665_ = new_n17851_ & ~new_n45664_;
  assign new_n45666_ = ~new_n45662_ & ~new_n45665_;
  assign new_n45667_ = ~new_n45658_ & new_n45666_;
  assign new_n45668_ = pi0788 & ~new_n45667_;
  assign new_n45669_ = ~new_n45657_ & ~new_n45668_;
  assign new_n45670_ = ~new_n20364_ & ~new_n45669_;
  assign new_n45671_ = ~new_n17968_ & new_n45649_;
  assign new_n45672_ = new_n17968_ & new_n45638_;
  assign new_n45673_ = ~new_n45671_ & ~new_n45672_;
  assign new_n45674_ = new_n18007_ & ~new_n45673_;
  assign new_n45675_ = new_n19281_ & ~new_n45652_;
  assign new_n45676_ = ~pi0628 & new_n45675_;
  assign new_n45677_ = ~new_n45638_ & ~new_n45676_;
  assign new_n45678_ = ~pi1156 & ~new_n45677_;
  assign new_n45679_ = pi0629 & ~new_n45678_;
  assign new_n45680_ = ~new_n45674_ & new_n45679_;
  assign new_n45681_ = new_n18008_ & ~new_n45673_;
  assign new_n45682_ = pi0628 & new_n45675_;
  assign new_n45683_ = ~new_n45638_ & ~new_n45682_;
  assign new_n45684_ = pi1156 & ~new_n45683_;
  assign new_n45685_ = ~pi0629 & ~new_n45684_;
  assign new_n45686_ = ~new_n45681_ & new_n45685_;
  assign new_n45687_ = pi0792 & ~new_n45686_;
  assign new_n45688_ = ~new_n45680_ & new_n45687_;
  assign new_n45689_ = ~new_n45670_ & ~new_n45688_;
  assign new_n45690_ = ~pi0647 & ~new_n45689_;
  assign new_n45691_ = ~new_n17762_ & ~new_n45673_;
  assign new_n45692_ = new_n17762_ & new_n45638_;
  assign new_n45693_ = ~new_n45691_ & ~new_n45692_;
  assign new_n45694_ = pi0647 & ~new_n45693_;
  assign new_n45695_ = ~pi1157 & ~new_n45694_;
  assign new_n45696_ = ~new_n45690_ & new_n45695_;
  assign new_n45697_ = ~new_n19311_ & new_n45675_;
  assign new_n45698_ = pi0647 & new_n45697_;
  assign new_n45699_ = pi1157 & ~new_n45638_;
  assign new_n45700_ = ~new_n45698_ & new_n45699_;
  assign new_n45701_ = ~pi0630 & ~new_n45700_;
  assign new_n45702_ = ~new_n45696_ & new_n45701_;
  assign new_n45703_ = pi0647 & ~new_n45689_;
  assign new_n45704_ = ~pi0647 & ~new_n45693_;
  assign new_n45705_ = pi1157 & ~new_n45704_;
  assign new_n45706_ = ~new_n45703_ & new_n45705_;
  assign new_n45707_ = ~pi0647 & new_n45697_;
  assign new_n45708_ = ~pi1157 & ~new_n45638_;
  assign new_n45709_ = ~new_n45707_ & new_n45708_;
  assign new_n45710_ = pi0630 & ~new_n45709_;
  assign new_n45711_ = ~new_n45706_ & new_n45710_;
  assign new_n45712_ = ~new_n45702_ & ~new_n45711_;
  assign new_n45713_ = pi0787 & ~new_n45712_;
  assign new_n45714_ = ~pi0787 & ~new_n45689_;
  assign new_n45715_ = ~new_n45713_ & ~new_n45714_;
  assign new_n45716_ = ~pi0790 & ~new_n45715_;
  assign new_n45717_ = ~pi0644 & ~new_n45715_;
  assign new_n45718_ = ~new_n19335_ & new_n45697_;
  assign new_n45719_ = ~new_n45638_ & ~new_n45718_;
  assign new_n45720_ = pi0644 & ~new_n45719_;
  assign new_n45721_ = ~pi0715 & ~new_n45720_;
  assign new_n45722_ = ~new_n45717_ & new_n45721_;
  assign new_n45723_ = ~new_n17804_ & new_n45691_;
  assign new_n45724_ = ~pi0644 & new_n45723_;
  assign new_n45725_ = pi0715 & ~new_n45638_;
  assign new_n45726_ = ~new_n45724_ & new_n45725_;
  assign new_n45727_ = ~new_n45722_ & ~new_n45726_;
  assign new_n45728_ = ~pi1160 & ~new_n45727_;
  assign new_n45729_ = pi0644 & new_n45715_;
  assign new_n45730_ = ~pi0644 & new_n45719_;
  assign new_n45731_ = pi0715 & ~new_n45730_;
  assign new_n45732_ = ~new_n45729_ & new_n45731_;
  assign new_n45733_ = pi0644 & new_n45723_;
  assign new_n45734_ = ~new_n45638_ & ~new_n45733_;
  assign new_n45735_ = ~pi0715 & ~new_n45734_;
  assign new_n45736_ = pi1160 & ~new_n45735_;
  assign new_n45737_ = ~new_n45732_ & new_n45736_;
  assign new_n45738_ = pi0790 & ~new_n45737_;
  assign new_n45739_ = ~new_n45728_ & new_n45738_;
  assign new_n45740_ = ~new_n45716_ & ~new_n45739_;
  assign new_n45741_ = pi0230 & ~new_n45740_;
  assign new_n45742_ = ~pi0230 & new_n45637_;
  assign po0724 = new_n45741_ | new_n45742_;
  assign new_n45744_ = pi0568 & ~new_n34791_;
  assign new_n45745_ = pi0245 & new_n34791_;
  assign po0725 = new_n45744_ | new_n45745_;
  assign new_n45747_ = pi0569 & ~new_n34791_;
  assign new_n45748_ = ~pi0239 & new_n34791_;
  assign po0726 = ~new_n45747_ & ~new_n45748_;
  assign new_n45750_ = new_n34791_ & new_n45455_;
  assign new_n45751_ = pi0570 & ~new_n45750_;
  assign new_n45752_ = ~pi0570 & new_n34786_;
  assign new_n45753_ = new_n45479_ & new_n45752_;
  assign po0727 = new_n45751_ | new_n45753_;
  assign new_n45755_ = pi0571 & ~new_n36139_;
  assign new_n45756_ = pi0241 & new_n36139_;
  assign po0728 = new_n45755_ | new_n45756_;
  assign new_n45758_ = pi0572 & ~new_n36139_;
  assign new_n45759_ = pi0244 & new_n36139_;
  assign po0729 = new_n45758_ | new_n45759_;
  assign new_n45761_ = pi0573 & ~new_n36139_;
  assign new_n45762_ = pi0242 & new_n36139_;
  assign po0730 = new_n45761_ | new_n45762_;
  assign new_n45764_ = pi0574 & ~new_n34783_;
  assign new_n45765_ = pi0241 & new_n34783_;
  assign po0731 = new_n45764_ | new_n45765_;
  assign new_n45767_ = pi0575 & ~new_n36139_;
  assign new_n45768_ = pi0235 & new_n36139_;
  assign po0732 = new_n45767_ | new_n45768_;
  assign new_n45770_ = pi0576 & ~new_n36139_;
  assign new_n45771_ = pi0248 & new_n36139_;
  assign po0733 = new_n45770_ | new_n45771_;
  assign new_n45773_ = pi0577 & ~new_n36111_;
  assign new_n45774_ = pi0238 & new_n36111_;
  assign po0734 = new_n45773_ | new_n45774_;
  assign new_n45776_ = pi0578 & ~new_n34783_;
  assign new_n45777_ = pi0249 & new_n34783_;
  assign po0735 = new_n45776_ | new_n45777_;
  assign new_n45779_ = pi0579 & ~new_n34775_;
  assign new_n45780_ = pi0249 & new_n34775_;
  assign po0736 = new_n45779_ | new_n45780_;
  assign new_n45782_ = pi0580 & ~new_n36111_;
  assign new_n45783_ = pi0245 & new_n36111_;
  assign po0737 = new_n45782_ | new_n45783_;
  assign new_n45785_ = pi0581 & ~new_n34783_;
  assign new_n45786_ = pi0235 & new_n34783_;
  assign po0738 = new_n45785_ | new_n45786_;
  assign new_n45788_ = pi0582 & ~new_n34783_;
  assign new_n45789_ = pi0240 & new_n34783_;
  assign po0739 = new_n45788_ | new_n45789_;
  assign new_n45791_ = pi0584 & ~new_n34783_;
  assign new_n45792_ = pi0245 & new_n34783_;
  assign po0741 = new_n45791_ | new_n45792_;
  assign new_n45794_ = pi0585 & ~new_n34783_;
  assign new_n45795_ = pi0244 & new_n34783_;
  assign po0742 = new_n45794_ | new_n45795_;
  assign new_n45797_ = pi0586 & ~new_n34783_;
  assign new_n45798_ = pi0242 & new_n34783_;
  assign po0743 = new_n45797_ | new_n45798_;
  assign new_n45800_ = ~pi0230 & pi0587;
  assign new_n45801_ = pi0230 & new_n16639_;
  assign new_n45802_ = ~new_n20223_ & new_n45801_;
  assign new_n45803_ = ~new_n35636_ & new_n45802_;
  assign new_n45804_ = new_n20235_ & new_n45803_;
  assign new_n45805_ = new_n30802_ & new_n45804_;
  assign po0744 = new_n45800_ | new_n45805_;
  assign new_n45807_ = ~pi0123 & new_n12202_;
  assign new_n45808_ = ~pi0591 & new_n45807_;
  assign new_n45809_ = ~pi0588 & ~new_n45807_;
  assign new_n45810_ = new_n44706_ & ~new_n45809_;
  assign po0745 = ~new_n45808_ & new_n45810_;
  assign new_n45812_ = ~pi0201 & new_n45454_;
  assign new_n45813_ = ~pi0204 & new_n45430_;
  assign new_n45814_ = pi0233 & ~new_n45813_;
  assign new_n45815_ = ~new_n45812_ & new_n45814_;
  assign new_n45816_ = ~pi0202 & new_n45454_;
  assign new_n45817_ = ~pi0205 & new_n45430_;
  assign new_n45818_ = ~pi0233 & ~new_n45817_;
  assign new_n45819_ = ~new_n45816_ & new_n45818_;
  assign new_n45820_ = ~new_n45815_ & ~new_n45819_;
  assign new_n45821_ = pi0237 & ~new_n45820_;
  assign new_n45822_ = ~pi0220 & new_n45454_;
  assign new_n45823_ = ~pi0206 & new_n45430_;
  assign new_n45824_ = pi0233 & ~new_n45823_;
  assign new_n45825_ = ~new_n45822_ & new_n45824_;
  assign new_n45826_ = ~pi0203 & new_n45454_;
  assign new_n45827_ = ~pi0218 & new_n45430_;
  assign new_n45828_ = ~pi0233 & ~new_n45827_;
  assign new_n45829_ = ~new_n45826_ & new_n45828_;
  assign new_n45830_ = ~new_n45825_ & ~new_n45829_;
  assign new_n45831_ = ~pi0237 & ~new_n45830_;
  assign po0746 = ~new_n45821_ & ~new_n45831_;
  assign new_n45833_ = pi0590 & ~new_n45807_;
  assign new_n45834_ = pi0588 & new_n45807_;
  assign new_n45835_ = new_n44706_ & ~new_n45834_;
  assign po0747 = new_n45833_ | ~new_n45835_;
  assign new_n45837_ = ~pi0592 & new_n45807_;
  assign new_n45838_ = ~pi0591 & ~new_n45807_;
  assign new_n45839_ = new_n44706_ & ~new_n45838_;
  assign po0748 = ~new_n45837_ & new_n45839_;
  assign new_n45841_ = ~pi0590 & new_n45807_;
  assign new_n45842_ = ~pi0592 & ~new_n45807_;
  assign new_n45843_ = new_n44706_ & ~new_n45842_;
  assign po0749 = ~new_n45841_ & new_n45843_;
  assign new_n45845_ = pi0234 & new_n45430_;
  assign new_n45846_ = pi0557 & ~new_n45845_;
  assign new_n45847_ = pi0246 & pi0536;
  assign new_n45848_ = ~pi0246 & ~pi0536;
  assign new_n45849_ = ~new_n45847_ & ~new_n45848_;
  assign new_n45850_ = ~pi0557 & ~new_n45431_;
  assign new_n45851_ = ~new_n45849_ & ~new_n45850_;
  assign new_n45852_ = ~new_n45846_ & new_n45851_;
  assign new_n45853_ = ~pi0538 & new_n45852_;
  assign new_n45854_ = ~pi0249 & ~new_n45853_;
  assign new_n45855_ = pi0538 & new_n45852_;
  assign new_n45856_ = pi0249 & ~new_n45855_;
  assign new_n45857_ = ~new_n45854_ & ~new_n45856_;
  assign new_n45858_ = ~pi0537 & new_n45857_;
  assign new_n45859_ = ~pi0248 & ~new_n45858_;
  assign new_n45860_ = pi0537 & new_n45857_;
  assign new_n45861_ = pi0248 & ~new_n45860_;
  assign new_n45862_ = ~new_n45859_ & ~new_n45861_;
  assign new_n45863_ = pi0241 & pi0506;
  assign new_n45864_ = ~pi0241 & ~pi0506;
  assign new_n45865_ = ~new_n45863_ & ~new_n45864_;
  assign new_n45866_ = new_n45862_ & ~new_n45865_;
  assign new_n45867_ = pi0240 & pi0535;
  assign new_n45868_ = ~pi0240 & ~pi0535;
  assign new_n45869_ = ~new_n45867_ & ~new_n45868_;
  assign new_n45870_ = new_n45866_ & ~new_n45869_;
  assign new_n45871_ = pi0534 & new_n45870_;
  assign new_n45872_ = ~pi0239 & ~new_n45871_;
  assign new_n45873_ = ~pi0534 & new_n45870_;
  assign new_n45874_ = pi0239 & ~new_n45873_;
  assign new_n45875_ = ~new_n45872_ & ~new_n45874_;
  assign new_n45876_ = pi0504 & new_n45875_;
  assign new_n45877_ = pi0242 & ~new_n45876_;
  assign new_n45878_ = ~pi0504 & new_n45875_;
  assign new_n45879_ = ~pi0242 & ~new_n45878_;
  assign new_n45880_ = ~new_n45877_ & ~new_n45879_;
  assign new_n45881_ = pi0533 & new_n45880_;
  assign new_n45882_ = pi0235 & ~new_n45881_;
  assign new_n45883_ = ~pi0533 & new_n45880_;
  assign new_n45884_ = ~pi0235 & ~new_n45883_;
  assign new_n45885_ = ~new_n45882_ & ~new_n45884_;
  assign new_n45886_ = pi0558 & new_n45885_;
  assign new_n45887_ = pi0244 & ~new_n45886_;
  assign new_n45888_ = ~pi0558 & new_n45885_;
  assign new_n45889_ = ~pi0244 & ~new_n45888_;
  assign new_n45890_ = ~new_n45887_ & ~new_n45889_;
  assign new_n45891_ = pi0509 & new_n45890_;
  assign new_n45892_ = pi0245 & ~new_n45891_;
  assign new_n45893_ = ~pi0509 & new_n45890_;
  assign new_n45894_ = ~pi0245 & ~new_n45893_;
  assign new_n45895_ = ~new_n45892_ & ~new_n45894_;
  assign new_n45896_ = pi0508 & new_n45895_;
  assign new_n45897_ = pi0247 & ~new_n45896_;
  assign new_n45898_ = pi0248 & pi0481;
  assign new_n45899_ = ~pi0248 & ~pi0481;
  assign new_n45900_ = ~new_n45898_ & ~new_n45899_;
  assign new_n45901_ = pi0234 & new_n45454_;
  assign new_n45902_ = pi0511 & ~new_n45901_;
  assign new_n45903_ = pi0246 & pi0487;
  assign new_n45904_ = ~pi0246 & ~pi0487;
  assign new_n45905_ = ~new_n45903_ & ~new_n45904_;
  assign new_n45906_ = ~pi0511 & ~new_n45455_;
  assign new_n45907_ = ~new_n45905_ & ~new_n45906_;
  assign new_n45908_ = ~new_n45902_ & new_n45907_;
  assign new_n45909_ = ~pi0249 & ~pi0579;
  assign new_n45910_ = pi0249 & pi0579;
  assign new_n45911_ = ~new_n45909_ & ~new_n45910_;
  assign new_n45912_ = new_n45908_ & ~new_n45911_;
  assign new_n45913_ = ~new_n45900_ & new_n45912_;
  assign new_n45914_ = pi0559 & new_n45913_;
  assign new_n45915_ = pi0241 & ~new_n45914_;
  assign new_n45916_ = ~pi0559 & new_n45913_;
  assign new_n45917_ = ~pi0241 & ~new_n45916_;
  assign new_n45918_ = ~new_n45915_ & ~new_n45917_;
  assign new_n45919_ = pi0515 & new_n45918_;
  assign new_n45920_ = pi0240 & ~new_n45919_;
  assign new_n45921_ = ~pi0579 & ~new_n45912_;
  assign new_n45922_ = ~new_n45854_ & new_n45908_;
  assign new_n45923_ = pi0579 & ~new_n45922_;
  assign new_n45924_ = ~new_n45921_ & ~new_n45923_;
  assign new_n45925_ = ~new_n45857_ & ~new_n45924_;
  assign new_n45926_ = ~pi0537 & ~new_n45925_;
  assign new_n45927_ = pi0537 & new_n45912_;
  assign new_n45928_ = ~pi0248 & ~new_n45927_;
  assign new_n45929_ = ~new_n45926_ & new_n45928_;
  assign new_n45930_ = ~new_n45861_ & ~new_n45929_;
  assign new_n45931_ = ~pi0481 & ~new_n45930_;
  assign new_n45932_ = pi0537 & ~new_n45925_;
  assign new_n45933_ = ~pi0537 & new_n45912_;
  assign new_n45934_ = pi0248 & ~new_n45933_;
  assign new_n45935_ = ~new_n45932_ & new_n45934_;
  assign new_n45936_ = ~new_n45859_ & ~new_n45935_;
  assign new_n45937_ = pi0481 & ~new_n45936_;
  assign new_n45938_ = ~new_n45931_ & ~new_n45937_;
  assign new_n45939_ = ~pi0559 & new_n45938_;
  assign new_n45940_ = pi0559 & new_n45862_;
  assign new_n45941_ = ~pi0241 & ~new_n45940_;
  assign new_n45942_ = ~new_n45939_ & new_n45941_;
  assign new_n45943_ = ~new_n45915_ & ~new_n45942_;
  assign new_n45944_ = ~pi0506 & ~new_n45943_;
  assign new_n45945_ = pi0559 & new_n45938_;
  assign new_n45946_ = ~pi0559 & new_n45862_;
  assign new_n45947_ = pi0241 & ~new_n45946_;
  assign new_n45948_ = ~new_n45945_ & new_n45947_;
  assign new_n45949_ = ~new_n45917_ & ~new_n45948_;
  assign new_n45950_ = pi0506 & ~new_n45949_;
  assign new_n45951_ = ~new_n45944_ & ~new_n45950_;
  assign new_n45952_ = ~pi0515 & new_n45951_;
  assign new_n45953_ = pi0515 & new_n45866_;
  assign new_n45954_ = ~pi0240 & ~new_n45953_;
  assign new_n45955_ = ~new_n45952_ & new_n45954_;
  assign new_n45956_ = ~new_n45920_ & ~new_n45955_;
  assign new_n45957_ = ~pi0535 & ~new_n45956_;
  assign new_n45958_ = ~pi0515 & new_n45918_;
  assign new_n45959_ = ~pi0240 & ~new_n45958_;
  assign new_n45960_ = pi0515 & new_n45951_;
  assign new_n45961_ = ~pi0515 & new_n45866_;
  assign new_n45962_ = pi0240 & ~new_n45961_;
  assign new_n45963_ = ~new_n45960_ & new_n45962_;
  assign new_n45964_ = ~new_n45959_ & ~new_n45963_;
  assign new_n45965_ = pi0535 & ~new_n45964_;
  assign new_n45966_ = ~new_n45957_ & ~new_n45965_;
  assign new_n45967_ = ~pi0534 & new_n45966_;
  assign new_n45968_ = ~new_n45920_ & ~new_n45959_;
  assign new_n45969_ = pi0534 & new_n45968_;
  assign new_n45970_ = pi0239 & ~new_n45969_;
  assign new_n45971_ = ~new_n45967_ & new_n45970_;
  assign new_n45972_ = ~new_n45872_ & ~new_n45971_;
  assign new_n45973_ = ~pi0488 & ~new_n45972_;
  assign new_n45974_ = pi0534 & new_n45966_;
  assign new_n45975_ = ~pi0534 & new_n45968_;
  assign new_n45976_ = ~pi0239 & ~new_n45975_;
  assign new_n45977_ = ~new_n45974_ & new_n45976_;
  assign new_n45978_ = ~new_n45874_ & ~new_n45977_;
  assign new_n45979_ = pi0488 & ~new_n45978_;
  assign new_n45980_ = ~new_n45973_ & ~new_n45979_;
  assign new_n45981_ = ~pi0504 & new_n45980_;
  assign new_n45982_ = ~pi0239 & pi0488;
  assign new_n45983_ = pi0239 & ~pi0488;
  assign new_n45984_ = ~new_n45982_ & ~new_n45983_;
  assign new_n45985_ = new_n45968_ & ~new_n45984_;
  assign new_n45986_ = pi0504 & new_n45985_;
  assign new_n45987_ = ~pi0242 & ~new_n45986_;
  assign new_n45988_ = ~new_n45981_ & new_n45987_;
  assign new_n45989_ = ~new_n45877_ & ~new_n45988_;
  assign new_n45990_ = ~pi0510 & ~new_n45989_;
  assign new_n45991_ = pi0504 & new_n45980_;
  assign new_n45992_ = ~pi0504 & new_n45985_;
  assign new_n45993_ = pi0242 & ~new_n45992_;
  assign new_n45994_ = ~new_n45991_ & new_n45993_;
  assign new_n45995_ = ~new_n45879_ & ~new_n45994_;
  assign new_n45996_ = pi0510 & ~new_n45995_;
  assign new_n45997_ = ~new_n45990_ & ~new_n45996_;
  assign new_n45998_ = ~pi0533 & new_n45997_;
  assign new_n45999_ = pi0242 & pi0510;
  assign new_n46000_ = ~pi0242 & ~pi0510;
  assign new_n46001_ = ~new_n45999_ & ~new_n46000_;
  assign new_n46002_ = new_n45985_ & ~new_n46001_;
  assign new_n46003_ = pi0533 & new_n46002_;
  assign new_n46004_ = ~pi0235 & ~new_n46003_;
  assign new_n46005_ = ~new_n45998_ & new_n46004_;
  assign new_n46006_ = ~new_n45882_ & ~new_n46005_;
  assign new_n46007_ = ~pi0512 & ~new_n46006_;
  assign new_n46008_ = pi0533 & new_n45997_;
  assign new_n46009_ = ~pi0533 & new_n46002_;
  assign new_n46010_ = pi0235 & ~new_n46009_;
  assign new_n46011_ = ~new_n46008_ & new_n46010_;
  assign new_n46012_ = ~new_n45884_ & ~new_n46011_;
  assign new_n46013_ = pi0512 & ~new_n46012_;
  assign new_n46014_ = ~new_n46007_ & ~new_n46013_;
  assign new_n46015_ = ~pi0558 & new_n46014_;
  assign new_n46016_ = pi0235 & pi0512;
  assign new_n46017_ = ~pi0235 & ~pi0512;
  assign new_n46018_ = ~new_n46016_ & ~new_n46017_;
  assign new_n46019_ = new_n46002_ & ~new_n46018_;
  assign new_n46020_ = pi0558 & new_n46019_;
  assign new_n46021_ = ~pi0244 & ~new_n46020_;
  assign new_n46022_ = ~new_n46015_ & new_n46021_;
  assign new_n46023_ = ~new_n45887_ & ~new_n46022_;
  assign new_n46024_ = ~pi0513 & ~new_n46023_;
  assign new_n46025_ = pi0558 & new_n46014_;
  assign new_n46026_ = ~pi0558 & new_n46019_;
  assign new_n46027_ = pi0244 & ~new_n46026_;
  assign new_n46028_ = ~new_n46025_ & new_n46027_;
  assign new_n46029_ = ~new_n45889_ & ~new_n46028_;
  assign new_n46030_ = pi0513 & ~new_n46029_;
  assign new_n46031_ = ~new_n46024_ & ~new_n46030_;
  assign new_n46032_ = ~pi0509 & new_n46031_;
  assign new_n46033_ = pi0244 & pi0513;
  assign new_n46034_ = ~pi0244 & ~pi0513;
  assign new_n46035_ = ~new_n46033_ & ~new_n46034_;
  assign new_n46036_ = new_n46019_ & ~new_n46035_;
  assign new_n46037_ = pi0509 & new_n46036_;
  assign new_n46038_ = ~pi0245 & ~new_n46037_;
  assign new_n46039_ = ~new_n46032_ & new_n46038_;
  assign new_n46040_ = ~new_n45892_ & ~new_n46039_;
  assign new_n46041_ = ~pi0514 & ~new_n46040_;
  assign new_n46042_ = pi0509 & new_n46031_;
  assign new_n46043_ = ~pi0509 & new_n46036_;
  assign new_n46044_ = pi0245 & ~new_n46043_;
  assign new_n46045_ = ~new_n46042_ & new_n46044_;
  assign new_n46046_ = ~new_n45894_ & ~new_n46045_;
  assign new_n46047_ = pi0514 & ~new_n46046_;
  assign new_n46048_ = ~new_n46041_ & ~new_n46047_;
  assign new_n46049_ = ~pi0508 & new_n46048_;
  assign new_n46050_ = pi0245 & pi0514;
  assign new_n46051_ = ~pi0245 & ~pi0514;
  assign new_n46052_ = ~new_n46050_ & ~new_n46051_;
  assign new_n46053_ = new_n46036_ & ~new_n46052_;
  assign new_n46054_ = pi0508 & new_n46053_;
  assign new_n46055_ = ~pi0247 & ~new_n46054_;
  assign new_n46056_ = ~new_n46049_ & new_n46055_;
  assign new_n46057_ = ~new_n45897_ & ~new_n46056_;
  assign new_n46058_ = ~pi0516 & ~new_n46057_;
  assign new_n46059_ = ~pi0508 & new_n45895_;
  assign new_n46060_ = ~pi0247 & ~new_n46059_;
  assign new_n46061_ = pi0508 & new_n46048_;
  assign new_n46062_ = ~pi0508 & new_n46053_;
  assign new_n46063_ = pi0247 & ~new_n46062_;
  assign new_n46064_ = ~new_n46061_ & new_n46063_;
  assign new_n46065_ = ~new_n46060_ & ~new_n46064_;
  assign new_n46066_ = pi0516 & ~new_n46065_;
  assign new_n46067_ = ~new_n46058_ & ~new_n46066_;
  assign new_n46068_ = ~pi0238 & new_n46067_;
  assign new_n46069_ = ~pi0517 & ~new_n46068_;
  assign new_n46070_ = ~new_n45897_ & ~new_n46060_;
  assign new_n46071_ = ~pi0238 & new_n46070_;
  assign new_n46072_ = pi0247 & pi0516;
  assign new_n46073_ = ~pi0247 & ~pi0516;
  assign new_n46074_ = ~new_n46072_ & ~new_n46073_;
  assign new_n46075_ = new_n46053_ & ~new_n46074_;
  assign new_n46076_ = pi0238 & new_n46075_;
  assign new_n46077_ = pi0517 & ~new_n46076_;
  assign new_n46078_ = ~new_n46071_ & new_n46077_;
  assign new_n46079_ = ~pi0507 & ~new_n46078_;
  assign new_n46080_ = ~new_n46069_ & new_n46079_;
  assign new_n46081_ = pi0238 & new_n46067_;
  assign new_n46082_ = pi0517 & ~new_n46081_;
  assign new_n46083_ = pi0238 & new_n46070_;
  assign new_n46084_ = ~pi0238 & new_n46075_;
  assign new_n46085_ = ~pi0517 & ~new_n46084_;
  assign new_n46086_ = ~new_n46083_ & new_n46085_;
  assign new_n46087_ = pi0507 & ~new_n46086_;
  assign new_n46088_ = ~new_n46082_ & new_n46087_;
  assign new_n46089_ = ~new_n46080_ & ~new_n46088_;
  assign new_n46090_ = pi0233 & ~new_n46089_;
  assign new_n46091_ = ~pi0247 & ~pi0561;
  assign new_n46092_ = pi0240 & pi0542;
  assign new_n46093_ = ~pi0240 & ~pi0542;
  assign new_n46094_ = ~new_n46092_ & ~new_n46093_;
  assign new_n46095_ = ~pi0505 & ~new_n45431_;
  assign new_n46096_ = pi0505 & ~new_n45845_;
  assign new_n46097_ = ~pi0246 & ~pi0499;
  assign new_n46098_ = pi0246 & pi0499;
  assign new_n46099_ = ~new_n46097_ & ~new_n46098_;
  assign new_n46100_ = ~pi0248 & ~pi0501;
  assign new_n46101_ = pi0248 & pi0501;
  assign new_n46102_ = ~new_n46100_ & ~new_n46101_;
  assign new_n46103_ = pi0249 & ~pi0496;
  assign new_n46104_ = ~pi0249 & pi0496;
  assign new_n46105_ = ~new_n46103_ & ~new_n46104_;
  assign new_n46106_ = ~new_n46102_ & new_n46105_;
  assign new_n46107_ = ~new_n46099_ & new_n46106_;
  assign new_n46108_ = ~new_n46096_ & new_n46107_;
  assign new_n46109_ = ~new_n46095_ & new_n46108_;
  assign new_n46110_ = ~pi0241 & ~pi0500;
  assign new_n46111_ = pi0241 & pi0500;
  assign new_n46112_ = ~new_n46110_ & ~new_n46111_;
  assign new_n46113_ = new_n46109_ & ~new_n46112_;
  assign new_n46114_ = ~new_n46094_ & new_n46113_;
  assign new_n46115_ = pi0497 & new_n46114_;
  assign new_n46116_ = ~pi0239 & ~new_n46115_;
  assign new_n46117_ = ~pi0497 & new_n46114_;
  assign new_n46118_ = pi0239 & ~new_n46117_;
  assign new_n46119_ = ~new_n46116_ & ~new_n46118_;
  assign new_n46120_ = pi0539 & new_n46119_;
  assign new_n46121_ = pi0242 & ~new_n46120_;
  assign new_n46122_ = ~pi0539 & new_n46119_;
  assign new_n46123_ = ~pi0242 & ~new_n46122_;
  assign new_n46124_ = ~new_n46121_ & ~new_n46123_;
  assign new_n46125_ = pi0540 & new_n46124_;
  assign new_n46126_ = pi0235 & ~new_n46125_;
  assign new_n46127_ = ~pi0540 & new_n46124_;
  assign new_n46128_ = ~pi0235 & ~new_n46127_;
  assign new_n46129_ = ~new_n46126_ & ~new_n46128_;
  assign new_n46130_ = pi0244 & pi0541;
  assign new_n46131_ = ~pi0244 & ~pi0541;
  assign new_n46132_ = ~new_n46130_ & ~new_n46131_;
  assign new_n46133_ = new_n46129_ & ~new_n46132_;
  assign new_n46134_ = pi0245 & pi0503;
  assign new_n46135_ = ~pi0245 & ~pi0503;
  assign new_n46136_ = ~new_n46134_ & ~new_n46135_;
  assign new_n46137_ = new_n46133_ & ~new_n46136_;
  assign new_n46138_ = ~pi0502 & new_n46137_;
  assign new_n46139_ = ~pi0247 & ~new_n46138_;
  assign new_n46140_ = ~new_n46091_ & ~new_n46139_;
  assign new_n46141_ = ~pi0518 & ~new_n45455_;
  assign new_n46142_ = pi0518 & ~new_n45901_;
  assign new_n46143_ = pi0249 & ~pi0578;
  assign new_n46144_ = ~pi0249 & pi0578;
  assign new_n46145_ = ~new_n46143_ & ~new_n46144_;
  assign new_n46146_ = pi0248 & ~pi0521;
  assign new_n46147_ = ~pi0248 & pi0521;
  assign new_n46148_ = ~new_n46146_ & ~new_n46147_;
  assign new_n46149_ = new_n46145_ & new_n46148_;
  assign new_n46150_ = pi0241 & pi0574;
  assign new_n46151_ = ~pi0241 & ~pi0574;
  assign new_n46152_ = ~new_n46150_ & ~new_n46151_;
  assign new_n46153_ = pi0246 & ~pi0520;
  assign new_n46154_ = ~pi0246 & pi0520;
  assign new_n46155_ = ~new_n46153_ & ~new_n46154_;
  assign new_n46156_ = ~new_n46152_ & new_n46155_;
  assign new_n46157_ = new_n46149_ & new_n46156_;
  assign new_n46158_ = ~new_n46142_ & new_n46157_;
  assign new_n46159_ = ~new_n46141_ & new_n46158_;
  assign new_n46160_ = pi0582 & new_n46159_;
  assign new_n46161_ = pi0240 & ~new_n46160_;
  assign new_n46162_ = ~pi0582 & new_n46159_;
  assign new_n46163_ = ~pi0240 & ~new_n46162_;
  assign new_n46164_ = ~new_n46161_ & ~new_n46163_;
  assign new_n46165_ = ~pi0239 & pi0519;
  assign new_n46166_ = pi0239 & ~pi0519;
  assign new_n46167_ = ~new_n46165_ & ~new_n46166_;
  assign new_n46168_ = new_n46164_ & ~new_n46167_;
  assign new_n46169_ = pi0242 & pi0586;
  assign new_n46170_ = ~pi0242 & ~pi0586;
  assign new_n46171_ = ~new_n46169_ & ~new_n46170_;
  assign new_n46172_ = new_n46168_ & ~new_n46171_;
  assign new_n46173_ = pi0235 & pi0581;
  assign new_n46174_ = ~pi0235 & ~pi0581;
  assign new_n46175_ = ~new_n46173_ & ~new_n46174_;
  assign new_n46176_ = new_n46172_ & ~new_n46175_;
  assign new_n46177_ = pi0585 & new_n46176_;
  assign new_n46178_ = pi0244 & ~new_n46177_;
  assign new_n46179_ = ~pi0585 & new_n46176_;
  assign new_n46180_ = ~pi0244 & ~new_n46179_;
  assign new_n46181_ = ~new_n46178_ & ~new_n46180_;
  assign new_n46182_ = pi0584 & new_n46181_;
  assign new_n46183_ = pi0245 & ~new_n46182_;
  assign new_n46184_ = ~pi0500 & new_n46113_;
  assign new_n46185_ = new_n46109_ & new_n46111_;
  assign new_n46186_ = ~new_n46159_ & ~new_n46185_;
  assign new_n46187_ = ~new_n46184_ & new_n46186_;
  assign new_n46188_ = ~pi0582 & ~new_n46187_;
  assign new_n46189_ = pi0582 & new_n46113_;
  assign new_n46190_ = ~pi0240 & ~new_n46189_;
  assign new_n46191_ = ~new_n46188_ & new_n46190_;
  assign new_n46192_ = ~new_n46161_ & ~new_n46191_;
  assign new_n46193_ = ~pi0542 & ~new_n46192_;
  assign new_n46194_ = pi0582 & ~new_n46187_;
  assign new_n46195_ = ~pi0582 & new_n46113_;
  assign new_n46196_ = pi0240 & ~new_n46195_;
  assign new_n46197_ = ~new_n46194_ & new_n46196_;
  assign new_n46198_ = ~new_n46163_ & ~new_n46197_;
  assign new_n46199_ = pi0542 & ~new_n46198_;
  assign new_n46200_ = ~new_n46193_ & ~new_n46199_;
  assign new_n46201_ = ~pi0497 & new_n46200_;
  assign new_n46202_ = pi0497 & new_n46164_;
  assign new_n46203_ = pi0239 & ~new_n46202_;
  assign new_n46204_ = ~new_n46201_ & new_n46203_;
  assign new_n46205_ = ~new_n46116_ & ~new_n46204_;
  assign new_n46206_ = ~pi0519 & ~new_n46205_;
  assign new_n46207_ = pi0497 & new_n46200_;
  assign new_n46208_ = ~pi0497 & new_n46164_;
  assign new_n46209_ = ~pi0239 & ~new_n46208_;
  assign new_n46210_ = ~new_n46207_ & new_n46209_;
  assign new_n46211_ = ~new_n46118_ & ~new_n46210_;
  assign new_n46212_ = pi0519 & ~new_n46211_;
  assign new_n46213_ = ~new_n46206_ & ~new_n46212_;
  assign new_n46214_ = ~pi0539 & new_n46213_;
  assign new_n46215_ = pi0539 & new_n46168_;
  assign new_n46216_ = ~pi0242 & ~new_n46215_;
  assign new_n46217_ = ~new_n46214_ & new_n46216_;
  assign new_n46218_ = ~new_n46121_ & ~new_n46217_;
  assign new_n46219_ = ~pi0586 & ~new_n46218_;
  assign new_n46220_ = pi0539 & new_n46213_;
  assign new_n46221_ = ~pi0539 & new_n46168_;
  assign new_n46222_ = pi0242 & ~new_n46221_;
  assign new_n46223_ = ~new_n46220_ & new_n46222_;
  assign new_n46224_ = ~new_n46123_ & ~new_n46223_;
  assign new_n46225_ = pi0586 & ~new_n46224_;
  assign new_n46226_ = ~new_n46219_ & ~new_n46225_;
  assign new_n46227_ = ~pi0540 & new_n46226_;
  assign new_n46228_ = pi0540 & new_n46172_;
  assign new_n46229_ = ~pi0235 & ~new_n46228_;
  assign new_n46230_ = ~new_n46227_ & new_n46229_;
  assign new_n46231_ = ~new_n46126_ & ~new_n46230_;
  assign new_n46232_ = ~pi0581 & ~new_n46231_;
  assign new_n46233_ = pi0540 & new_n46226_;
  assign new_n46234_ = ~pi0540 & new_n46172_;
  assign new_n46235_ = pi0235 & ~new_n46234_;
  assign new_n46236_ = ~new_n46233_ & new_n46235_;
  assign new_n46237_ = ~new_n46128_ & ~new_n46236_;
  assign new_n46238_ = pi0581 & ~new_n46237_;
  assign new_n46239_ = ~new_n46232_ & ~new_n46238_;
  assign new_n46240_ = ~pi0585 & new_n46239_;
  assign new_n46241_ = pi0585 & new_n46129_;
  assign new_n46242_ = ~pi0244 & ~new_n46241_;
  assign new_n46243_ = ~new_n46240_ & new_n46242_;
  assign new_n46244_ = ~new_n46178_ & ~new_n46243_;
  assign new_n46245_ = ~pi0541 & ~new_n46244_;
  assign new_n46246_ = pi0585 & new_n46239_;
  assign new_n46247_ = ~pi0585 & new_n46129_;
  assign new_n46248_ = pi0244 & ~new_n46247_;
  assign new_n46249_ = ~new_n46246_ & new_n46248_;
  assign new_n46250_ = ~new_n46180_ & ~new_n46249_;
  assign new_n46251_ = pi0541 & ~new_n46250_;
  assign new_n46252_ = ~new_n46245_ & ~new_n46251_;
  assign new_n46253_ = ~pi0584 & new_n46252_;
  assign new_n46254_ = pi0584 & new_n46133_;
  assign new_n46255_ = ~pi0245 & ~new_n46254_;
  assign new_n46256_ = ~new_n46253_ & new_n46255_;
  assign new_n46257_ = ~new_n46183_ & ~new_n46256_;
  assign new_n46258_ = ~pi0503 & ~new_n46257_;
  assign new_n46259_ = ~pi0584 & new_n46181_;
  assign new_n46260_ = ~pi0245 & ~new_n46259_;
  assign new_n46261_ = pi0584 & new_n46252_;
  assign new_n46262_ = ~pi0584 & new_n46133_;
  assign new_n46263_ = pi0245 & ~new_n46262_;
  assign new_n46264_ = ~new_n46261_ & new_n46263_;
  assign new_n46265_ = ~new_n46260_ & ~new_n46264_;
  assign new_n46266_ = pi0503 & ~new_n46265_;
  assign new_n46267_ = ~new_n46258_ & ~new_n46266_;
  assign new_n46268_ = ~pi0502 & ~new_n46267_;
  assign new_n46269_ = ~new_n46183_ & ~new_n46260_;
  assign new_n46270_ = pi0502 & ~new_n46269_;
  assign new_n46271_ = ~pi0561 & ~new_n46270_;
  assign new_n46272_ = ~new_n46268_ & new_n46271_;
  assign new_n46273_ = ~new_n46140_ & ~new_n46272_;
  assign new_n46274_ = pi0247 & pi0561;
  assign new_n46275_ = pi0502 & new_n46137_;
  assign new_n46276_ = pi0247 & ~new_n46275_;
  assign new_n46277_ = ~new_n46274_ & ~new_n46276_;
  assign new_n46278_ = pi0502 & ~new_n46267_;
  assign new_n46279_ = ~pi0502 & ~new_n46269_;
  assign new_n46280_ = pi0561 & ~new_n46279_;
  assign new_n46281_ = ~new_n46278_ & new_n46280_;
  assign new_n46282_ = ~new_n46277_ & ~new_n46281_;
  assign new_n46283_ = ~new_n46273_ & ~new_n46282_;
  assign new_n46284_ = ~pi0238 & new_n46283_;
  assign new_n46285_ = ~pi0522 & ~new_n46284_;
  assign new_n46286_ = ~new_n46139_ & ~new_n46276_;
  assign new_n46287_ = ~pi0238 & new_n46286_;
  assign new_n46288_ = ~new_n46091_ & ~new_n46274_;
  assign new_n46289_ = new_n46269_ & ~new_n46288_;
  assign new_n46290_ = pi0238 & new_n46289_;
  assign new_n46291_ = pi0522 & ~new_n46290_;
  assign new_n46292_ = ~new_n46287_ & new_n46291_;
  assign new_n46293_ = ~pi0543 & ~new_n46292_;
  assign new_n46294_ = ~new_n46285_ & new_n46293_;
  assign new_n46295_ = pi0238 & new_n46283_;
  assign new_n46296_ = pi0522 & ~new_n46295_;
  assign new_n46297_ = pi0238 & new_n46286_;
  assign new_n46298_ = ~pi0238 & new_n46289_;
  assign new_n46299_ = ~pi0522 & ~new_n46298_;
  assign new_n46300_ = ~new_n46297_ & new_n46299_;
  assign new_n46301_ = pi0543 & ~new_n46300_;
  assign new_n46302_ = ~new_n46296_ & new_n46301_;
  assign new_n46303_ = ~new_n46294_ & ~new_n46302_;
  assign new_n46304_ = ~pi0233 & ~new_n46303_;
  assign new_n46305_ = pi0237 & ~new_n46304_;
  assign new_n46306_ = ~new_n46090_ & new_n46305_;
  assign new_n46307_ = ~pi0240 & ~pi0492;
  assign new_n46308_ = pi0240 & pi0492;
  assign new_n46309_ = ~new_n46307_ & ~new_n46308_;
  assign new_n46310_ = pi0241 & pi0490;
  assign new_n46311_ = ~pi0241 & ~pi0490;
  assign new_n46312_ = ~new_n46310_ & ~new_n46311_;
  assign new_n46313_ = pi0544 & ~new_n45845_;
  assign new_n46314_ = ~pi0544 & ~new_n45431_;
  assign new_n46315_ = pi0246 & pi0546;
  assign new_n46316_ = ~pi0246 & ~pi0546;
  assign new_n46317_ = ~new_n46315_ & ~new_n46316_;
  assign new_n46318_ = pi0248 & pi0548;
  assign new_n46319_ = ~pi0248 & ~pi0548;
  assign new_n46320_ = ~new_n46318_ & ~new_n46319_;
  assign new_n46321_ = pi0249 & pi0484;
  assign new_n46322_ = ~pi0249 & ~pi0484;
  assign new_n46323_ = ~new_n46321_ & ~new_n46322_;
  assign new_n46324_ = ~new_n46320_ & ~new_n46323_;
  assign new_n46325_ = ~new_n46317_ & new_n46324_;
  assign new_n46326_ = ~new_n46314_ & new_n46325_;
  assign new_n46327_ = ~new_n46313_ & new_n46326_;
  assign new_n46328_ = ~new_n46312_ & new_n46327_;
  assign new_n46329_ = ~new_n46309_ & new_n46328_;
  assign new_n46330_ = pi0494 & new_n46329_;
  assign new_n46331_ = ~pi0239 & ~new_n46330_;
  assign new_n46332_ = ~pi0494 & new_n46329_;
  assign new_n46333_ = pi0239 & ~new_n46332_;
  assign new_n46334_ = ~new_n46331_ & ~new_n46333_;
  assign new_n46335_ = pi0483 & new_n46334_;
  assign new_n46336_ = pi0242 & ~new_n46335_;
  assign new_n46337_ = ~pi0483 & new_n46334_;
  assign new_n46338_ = ~pi0242 & ~new_n46337_;
  assign new_n46339_ = ~new_n46336_ & ~new_n46338_;
  assign new_n46340_ = pi0495 & new_n46339_;
  assign new_n46341_ = pi0235 & ~new_n46340_;
  assign new_n46342_ = ~pi0495 & new_n46339_;
  assign new_n46343_ = ~pi0235 & ~new_n46342_;
  assign new_n46344_ = ~new_n46341_ & ~new_n46343_;
  assign new_n46345_ = pi0244 & pi0493;
  assign new_n46346_ = ~pi0244 & ~pi0493;
  assign new_n46347_ = ~new_n46345_ & ~new_n46346_;
  assign new_n46348_ = new_n46344_ & ~new_n46347_;
  assign new_n46349_ = pi0545 & new_n46348_;
  assign new_n46350_ = pi0245 & ~new_n46349_;
  assign new_n46351_ = ~pi0545 & new_n46348_;
  assign new_n46352_ = ~pi0245 & ~new_n46351_;
  assign new_n46353_ = ~new_n46350_ & ~new_n46352_;
  assign new_n46354_ = pi0547 & new_n46353_;
  assign new_n46355_ = pi0247 & ~new_n46354_;
  assign new_n46356_ = ~pi0523 & ~new_n45455_;
  assign new_n46357_ = pi0523 & ~new_n45901_;
  assign new_n46358_ = pi0246 & pi0526;
  assign new_n46359_ = ~pi0246 & ~pi0526;
  assign new_n46360_ = ~new_n46358_ & ~new_n46359_;
  assign new_n46361_ = pi0248 & pi0576;
  assign new_n46362_ = ~pi0248 & ~pi0576;
  assign new_n46363_ = ~new_n46361_ & ~new_n46362_;
  assign new_n46364_ = pi0249 & pi0528;
  assign new_n46365_ = ~pi0249 & ~pi0528;
  assign new_n46366_ = ~new_n46364_ & ~new_n46365_;
  assign new_n46367_ = ~new_n46363_ & ~new_n46366_;
  assign new_n46368_ = ~new_n46360_ & new_n46367_;
  assign new_n46369_ = ~new_n46357_ & new_n46368_;
  assign new_n46370_ = ~new_n46356_ & new_n46369_;
  assign new_n46371_ = pi0571 & new_n46370_;
  assign new_n46372_ = pi0241 & ~new_n46371_;
  assign new_n46373_ = ~pi0571 & new_n46370_;
  assign new_n46374_ = ~pi0241 & ~new_n46373_;
  assign new_n46375_ = ~new_n46372_ & ~new_n46374_;
  assign new_n46376_ = ~pi0530 & new_n46375_;
  assign new_n46377_ = ~pi0240 & ~new_n46376_;
  assign new_n46378_ = pi0530 & new_n46375_;
  assign new_n46379_ = pi0240 & ~new_n46378_;
  assign new_n46380_ = ~new_n46377_ & ~new_n46379_;
  assign new_n46381_ = ~pi0239 & pi0524;
  assign new_n46382_ = pi0239 & ~pi0524;
  assign new_n46383_ = ~new_n46381_ & ~new_n46382_;
  assign new_n46384_ = new_n46380_ & ~new_n46383_;
  assign new_n46385_ = pi0242 & pi0573;
  assign new_n46386_ = ~pi0242 & ~pi0573;
  assign new_n46387_ = ~new_n46385_ & ~new_n46386_;
  assign new_n46388_ = new_n46384_ & ~new_n46387_;
  assign new_n46389_ = pi0235 & pi0575;
  assign new_n46390_ = ~pi0235 & ~pi0575;
  assign new_n46391_ = ~new_n46389_ & ~new_n46390_;
  assign new_n46392_ = new_n46388_ & ~new_n46391_;
  assign new_n46393_ = pi0572 & new_n46392_;
  assign new_n46394_ = pi0244 & ~new_n46393_;
  assign new_n46395_ = ~new_n46307_ & ~new_n46377_;
  assign new_n46396_ = ~pi0241 & ~new_n46327_;
  assign new_n46397_ = ~new_n46373_ & new_n46396_;
  assign new_n46398_ = ~new_n46372_ & ~new_n46397_;
  assign new_n46399_ = ~pi0490 & ~new_n46398_;
  assign new_n46400_ = pi0241 & ~new_n46327_;
  assign new_n46401_ = ~new_n46371_ & new_n46400_;
  assign new_n46402_ = ~new_n46374_ & ~new_n46401_;
  assign new_n46403_ = pi0490 & ~new_n46402_;
  assign new_n46404_ = ~new_n46399_ & ~new_n46403_;
  assign new_n46405_ = ~pi0530 & ~new_n46404_;
  assign new_n46406_ = pi0530 & ~new_n46328_;
  assign new_n46407_ = ~pi0492 & ~new_n46406_;
  assign new_n46408_ = ~new_n46405_ & new_n46407_;
  assign new_n46409_ = ~new_n46395_ & ~new_n46408_;
  assign new_n46410_ = ~new_n46308_ & ~new_n46379_;
  assign new_n46411_ = pi0530 & ~new_n46404_;
  assign new_n46412_ = ~pi0530 & ~new_n46328_;
  assign new_n46413_ = pi0492 & ~new_n46412_;
  assign new_n46414_ = ~new_n46411_ & new_n46413_;
  assign new_n46415_ = ~new_n46410_ & ~new_n46414_;
  assign new_n46416_ = ~new_n46409_ & ~new_n46415_;
  assign new_n46417_ = ~pi0494 & new_n46416_;
  assign new_n46418_ = pi0494 & new_n46380_;
  assign new_n46419_ = pi0239 & ~new_n46418_;
  assign new_n46420_ = ~new_n46417_ & new_n46419_;
  assign new_n46421_ = ~new_n46331_ & ~new_n46420_;
  assign new_n46422_ = ~pi0524 & ~new_n46421_;
  assign new_n46423_ = pi0494 & new_n46416_;
  assign new_n46424_ = ~pi0494 & new_n46380_;
  assign new_n46425_ = ~pi0239 & ~new_n46424_;
  assign new_n46426_ = ~new_n46423_ & new_n46425_;
  assign new_n46427_ = ~new_n46333_ & ~new_n46426_;
  assign new_n46428_ = pi0524 & ~new_n46427_;
  assign new_n46429_ = ~new_n46422_ & ~new_n46428_;
  assign new_n46430_ = ~pi0483 & new_n46429_;
  assign new_n46431_ = pi0483 & new_n46384_;
  assign new_n46432_ = ~pi0242 & ~new_n46431_;
  assign new_n46433_ = ~new_n46430_ & new_n46432_;
  assign new_n46434_ = ~new_n46336_ & ~new_n46433_;
  assign new_n46435_ = ~pi0573 & ~new_n46434_;
  assign new_n46436_ = pi0483 & new_n46429_;
  assign new_n46437_ = ~pi0483 & new_n46384_;
  assign new_n46438_ = pi0242 & ~new_n46437_;
  assign new_n46439_ = ~new_n46436_ & new_n46438_;
  assign new_n46440_ = ~new_n46338_ & ~new_n46439_;
  assign new_n46441_ = pi0573 & ~new_n46440_;
  assign new_n46442_ = ~new_n46435_ & ~new_n46441_;
  assign new_n46443_ = ~pi0495 & new_n46442_;
  assign new_n46444_ = pi0495 & new_n46388_;
  assign new_n46445_ = ~pi0235 & ~new_n46444_;
  assign new_n46446_ = ~new_n46443_ & new_n46445_;
  assign new_n46447_ = ~new_n46341_ & ~new_n46446_;
  assign new_n46448_ = ~pi0575 & ~new_n46447_;
  assign new_n46449_ = pi0495 & new_n46442_;
  assign new_n46450_ = ~pi0495 & new_n46388_;
  assign new_n46451_ = pi0235 & ~new_n46450_;
  assign new_n46452_ = ~new_n46449_ & new_n46451_;
  assign new_n46453_ = ~new_n46343_ & ~new_n46452_;
  assign new_n46454_ = pi0575 & ~new_n46453_;
  assign new_n46455_ = ~new_n46448_ & ~new_n46454_;
  assign new_n46456_ = ~pi0572 & new_n46455_;
  assign new_n46457_ = pi0572 & new_n46344_;
  assign new_n46458_ = ~pi0244 & ~new_n46457_;
  assign new_n46459_ = ~new_n46456_ & new_n46458_;
  assign new_n46460_ = ~new_n46394_ & ~new_n46459_;
  assign new_n46461_ = ~pi0493 & ~new_n46460_;
  assign new_n46462_ = ~pi0572 & new_n46392_;
  assign new_n46463_ = ~pi0244 & ~new_n46462_;
  assign new_n46464_ = pi0572 & new_n46455_;
  assign new_n46465_ = ~pi0572 & new_n46344_;
  assign new_n46466_ = pi0244 & ~new_n46465_;
  assign new_n46467_ = ~new_n46464_ & new_n46466_;
  assign new_n46468_ = ~new_n46463_ & ~new_n46467_;
  assign new_n46469_ = pi0493 & ~new_n46468_;
  assign new_n46470_ = ~new_n46461_ & ~new_n46469_;
  assign new_n46471_ = ~pi0545 & new_n46470_;
  assign new_n46472_ = ~new_n46394_ & ~new_n46463_;
  assign new_n46473_ = pi0545 & new_n46472_;
  assign new_n46474_ = ~pi0245 & ~new_n46473_;
  assign new_n46475_ = ~new_n46471_ & new_n46474_;
  assign new_n46476_ = ~new_n46350_ & ~new_n46475_;
  assign new_n46477_ = ~pi0525 & ~new_n46476_;
  assign new_n46478_ = pi0545 & new_n46470_;
  assign new_n46479_ = ~pi0545 & new_n46472_;
  assign new_n46480_ = pi0245 & ~new_n46479_;
  assign new_n46481_ = ~new_n46478_ & new_n46480_;
  assign new_n46482_ = ~new_n46352_ & ~new_n46481_;
  assign new_n46483_ = pi0525 & ~new_n46482_;
  assign new_n46484_ = ~new_n46477_ & ~new_n46483_;
  assign new_n46485_ = ~pi0547 & new_n46484_;
  assign new_n46486_ = pi0245 & pi0525;
  assign new_n46487_ = ~pi0245 & ~pi0525;
  assign new_n46488_ = ~new_n46486_ & ~new_n46487_;
  assign new_n46489_ = new_n46472_ & ~new_n46488_;
  assign new_n46490_ = pi0547 & new_n46489_;
  assign new_n46491_ = ~pi0247 & ~new_n46490_;
  assign new_n46492_ = ~new_n46485_ & new_n46491_;
  assign new_n46493_ = ~new_n46355_ & ~new_n46492_;
  assign new_n46494_ = ~pi0527 & ~new_n46493_;
  assign new_n46495_ = ~pi0547 & new_n46353_;
  assign new_n46496_ = ~pi0247 & ~new_n46495_;
  assign new_n46497_ = pi0547 & new_n46484_;
  assign new_n46498_ = ~pi0547 & new_n46489_;
  assign new_n46499_ = pi0247 & ~new_n46498_;
  assign new_n46500_ = ~new_n46497_ & new_n46499_;
  assign new_n46501_ = ~new_n46496_ & ~new_n46500_;
  assign new_n46502_ = pi0527 & ~new_n46501_;
  assign new_n46503_ = ~new_n46494_ & ~new_n46502_;
  assign new_n46504_ = ~pi0238 & new_n46503_;
  assign new_n46505_ = ~pi0529 & ~new_n46504_;
  assign new_n46506_ = ~new_n46355_ & ~new_n46496_;
  assign new_n46507_ = ~pi0238 & new_n46506_;
  assign new_n46508_ = pi0247 & pi0527;
  assign new_n46509_ = ~pi0247 & ~pi0527;
  assign new_n46510_ = ~new_n46508_ & ~new_n46509_;
  assign new_n46511_ = new_n46489_ & ~new_n46510_;
  assign new_n46512_ = pi0238 & new_n46511_;
  assign new_n46513_ = pi0529 & ~new_n46512_;
  assign new_n46514_ = ~new_n46507_ & new_n46513_;
  assign new_n46515_ = ~pi0491 & ~new_n46514_;
  assign new_n46516_ = ~new_n46505_ & new_n46515_;
  assign new_n46517_ = pi0238 & new_n46503_;
  assign new_n46518_ = pi0529 & ~new_n46517_;
  assign new_n46519_ = pi0238 & new_n46506_;
  assign new_n46520_ = ~pi0238 & new_n46511_;
  assign new_n46521_ = ~pi0529 & ~new_n46520_;
  assign new_n46522_ = ~new_n46519_ & new_n46521_;
  assign new_n46523_ = pi0491 & ~new_n46522_;
  assign new_n46524_ = ~new_n46518_ & new_n46523_;
  assign new_n46525_ = ~new_n46516_ & ~new_n46524_;
  assign new_n46526_ = pi0233 & ~new_n46525_;
  assign new_n46527_ = ~pi0485 & ~new_n45431_;
  assign new_n46528_ = pi0485 & ~new_n45845_;
  assign new_n46529_ = pi0248 & ~pi0554;
  assign new_n46530_ = ~pi0248 & pi0554;
  assign new_n46531_ = ~new_n46529_ & ~new_n46530_;
  assign new_n46532_ = ~pi0246 & pi0563;
  assign new_n46533_ = pi0246 & ~pi0563;
  assign new_n46534_ = ~new_n46532_ & ~new_n46533_;
  assign new_n46535_ = new_n46531_ & new_n46534_;
  assign new_n46536_ = pi0240 & pi0551;
  assign new_n46537_ = ~pi0240 & ~pi0551;
  assign new_n46538_ = ~new_n46536_ & ~new_n46537_;
  assign new_n46539_ = pi0249 & ~pi0555;
  assign new_n46540_ = ~pi0249 & pi0555;
  assign new_n46541_ = ~new_n46539_ & ~new_n46540_;
  assign new_n46542_ = pi0241 & ~pi0553;
  assign new_n46543_ = ~pi0241 & pi0553;
  assign new_n46544_ = ~new_n46542_ & ~new_n46543_;
  assign new_n46545_ = new_n46541_ & new_n46544_;
  assign new_n46546_ = ~new_n46538_ & new_n46545_;
  assign new_n46547_ = new_n46535_ & new_n46546_;
  assign new_n46548_ = ~new_n46528_ & new_n46547_;
  assign new_n46549_ = ~new_n46527_ & new_n46548_;
  assign new_n46550_ = pi0550 & new_n46549_;
  assign new_n46551_ = ~pi0239 & ~new_n46550_;
  assign new_n46552_ = ~pi0550 & new_n46549_;
  assign new_n46553_ = pi0239 & ~new_n46552_;
  assign new_n46554_ = ~new_n46551_ & ~new_n46553_;
  assign new_n46555_ = ~pi0489 & new_n46554_;
  assign new_n46556_ = ~pi0242 & ~new_n46555_;
  assign new_n46557_ = pi0489 & new_n46554_;
  assign new_n46558_ = pi0242 & ~new_n46557_;
  assign new_n46559_ = ~new_n46556_ & ~new_n46558_;
  assign new_n46560_ = pi0549 & new_n46559_;
  assign new_n46561_ = pi0235 & ~new_n46560_;
  assign new_n46562_ = ~pi0549 & new_n46559_;
  assign new_n46563_ = ~pi0235 & ~new_n46562_;
  assign new_n46564_ = ~new_n46561_ & ~new_n46563_;
  assign new_n46565_ = pi0486 & new_n46564_;
  assign new_n46566_ = pi0244 & ~new_n46565_;
  assign new_n46567_ = ~pi0486 & new_n46564_;
  assign new_n46568_ = ~pi0244 & ~new_n46567_;
  assign new_n46569_ = ~new_n46566_ & ~new_n46568_;
  assign new_n46570_ = pi0245 & pi0580;
  assign new_n46571_ = ~pi0245 & ~pi0580;
  assign new_n46572_ = ~new_n46570_ & ~new_n46571_;
  assign new_n46573_ = new_n46569_ & ~new_n46572_;
  assign new_n46574_ = pi0552 & new_n46573_;
  assign new_n46575_ = pi0247 & ~new_n46574_;
  assign new_n46576_ = ~pi0242 & ~pi0556;
  assign new_n46577_ = pi0242 & pi0556;
  assign new_n46578_ = ~new_n46576_ & ~new_n46577_;
  assign new_n46579_ = ~pi0570 & ~new_n45455_;
  assign new_n46580_ = pi0570 & ~new_n45901_;
  assign new_n46581_ = pi0241 & pi0562;
  assign new_n46582_ = ~pi0241 & ~pi0562;
  assign new_n46583_ = ~new_n46581_ & ~new_n46582_;
  assign new_n46584_ = ~pi0249 & pi0482;
  assign new_n46585_ = ~pi0246 & pi0564;
  assign new_n46586_ = pi0249 & ~pi0482;
  assign new_n46587_ = ~new_n46585_ & ~new_n46586_;
  assign new_n46588_ = ~new_n46584_ & new_n46587_;
  assign new_n46589_ = ~new_n46583_ & new_n46588_;
  assign new_n46590_ = ~new_n46580_ & new_n46589_;
  assign new_n46591_ = ~new_n46579_ & new_n46590_;
  assign new_n46592_ = pi0240 & pi0560;
  assign new_n46593_ = ~pi0240 & ~pi0560;
  assign new_n46594_ = ~new_n46592_ & ~new_n46593_;
  assign new_n46595_ = pi0246 & ~pi0564;
  assign new_n46596_ = pi0248 & ~pi0565;
  assign new_n46597_ = ~pi0248 & pi0565;
  assign new_n46598_ = ~new_n46596_ & ~new_n46597_;
  assign new_n46599_ = ~new_n46595_ & new_n46598_;
  assign new_n46600_ = ~new_n46594_ & new_n46599_;
  assign new_n46601_ = new_n46591_ & new_n46600_;
  assign new_n46602_ = ~pi0240 & ~new_n46601_;
  assign new_n46603_ = pi0560 & ~new_n46595_;
  assign new_n46604_ = new_n46598_ & new_n46603_;
  assign new_n46605_ = new_n46591_ & new_n46604_;
  assign new_n46606_ = pi0240 & ~new_n46605_;
  assign new_n46607_ = ~new_n46602_ & ~new_n46606_;
  assign new_n46608_ = ~pi0239 & pi0569;
  assign new_n46609_ = pi0239 & ~pi0569;
  assign new_n46610_ = ~new_n46608_ & ~new_n46609_;
  assign new_n46611_ = new_n46607_ & ~new_n46610_;
  assign new_n46612_ = ~new_n46578_ & new_n46611_;
  assign new_n46613_ = pi0235 & pi0531;
  assign new_n46614_ = ~pi0235 & ~pi0531;
  assign new_n46615_ = ~new_n46613_ & ~new_n46614_;
  assign new_n46616_ = new_n46612_ & ~new_n46615_;
  assign new_n46617_ = pi0244 & pi0566;
  assign new_n46618_ = ~pi0244 & ~pi0566;
  assign new_n46619_ = ~new_n46617_ & ~new_n46618_;
  assign new_n46620_ = new_n46616_ & ~new_n46619_;
  assign new_n46621_ = pi0568 & new_n46620_;
  assign new_n46622_ = pi0245 & ~new_n46621_;
  assign new_n46623_ = ~new_n46556_ & ~new_n46576_;
  assign new_n46624_ = pi0569 & ~new_n46553_;
  assign new_n46625_ = new_n46607_ & new_n46624_;
  assign new_n46626_ = new_n46601_ & new_n46609_;
  assign new_n46627_ = ~new_n46554_ & ~new_n46626_;
  assign new_n46628_ = ~new_n46625_ & new_n46627_;
  assign new_n46629_ = ~pi0489 & new_n46628_;
  assign new_n46630_ = pi0489 & ~new_n46611_;
  assign new_n46631_ = ~pi0556 & ~new_n46630_;
  assign new_n46632_ = ~new_n46629_ & new_n46631_;
  assign new_n46633_ = ~new_n46623_ & ~new_n46632_;
  assign new_n46634_ = ~new_n46558_ & ~new_n46577_;
  assign new_n46635_ = pi0489 & new_n46628_;
  assign new_n46636_ = ~pi0489 & ~new_n46611_;
  assign new_n46637_ = pi0556 & ~new_n46636_;
  assign new_n46638_ = ~new_n46635_ & new_n46637_;
  assign new_n46639_ = ~new_n46634_ & ~new_n46638_;
  assign new_n46640_ = ~new_n46633_ & ~new_n46639_;
  assign new_n46641_ = ~pi0549 & new_n46640_;
  assign new_n46642_ = pi0549 & new_n46612_;
  assign new_n46643_ = ~pi0235 & ~new_n46642_;
  assign new_n46644_ = ~new_n46641_ & new_n46643_;
  assign new_n46645_ = ~new_n46561_ & ~new_n46644_;
  assign new_n46646_ = ~pi0531 & ~new_n46645_;
  assign new_n46647_ = pi0549 & new_n46640_;
  assign new_n46648_ = ~pi0549 & new_n46612_;
  assign new_n46649_ = pi0235 & ~new_n46648_;
  assign new_n46650_ = ~new_n46647_ & new_n46649_;
  assign new_n46651_ = ~new_n46563_ & ~new_n46650_;
  assign new_n46652_ = pi0531 & ~new_n46651_;
  assign new_n46653_ = ~new_n46646_ & ~new_n46652_;
  assign new_n46654_ = ~pi0486 & new_n46653_;
  assign new_n46655_ = pi0486 & new_n46616_;
  assign new_n46656_ = ~pi0244 & ~new_n46655_;
  assign new_n46657_ = ~new_n46654_ & new_n46656_;
  assign new_n46658_ = ~new_n46566_ & ~new_n46657_;
  assign new_n46659_ = ~pi0566 & ~new_n46658_;
  assign new_n46660_ = pi0486 & new_n46653_;
  assign new_n46661_ = ~pi0486 & new_n46616_;
  assign new_n46662_ = pi0244 & ~new_n46661_;
  assign new_n46663_ = ~new_n46660_ & new_n46662_;
  assign new_n46664_ = ~new_n46568_ & ~new_n46663_;
  assign new_n46665_ = pi0566 & ~new_n46664_;
  assign new_n46666_ = ~new_n46659_ & ~new_n46665_;
  assign new_n46667_ = ~pi0568 & new_n46666_;
  assign new_n46668_ = pi0568 & new_n46569_;
  assign new_n46669_ = ~pi0245 & ~new_n46668_;
  assign new_n46670_ = ~new_n46667_ & new_n46669_;
  assign new_n46671_ = ~new_n46622_ & ~new_n46670_;
  assign new_n46672_ = ~pi0580 & ~new_n46671_;
  assign new_n46673_ = ~pi0568 & new_n46620_;
  assign new_n46674_ = ~pi0245 & ~new_n46673_;
  assign new_n46675_ = pi0568 & new_n46666_;
  assign new_n46676_ = ~pi0568 & new_n46569_;
  assign new_n46677_ = pi0245 & ~new_n46676_;
  assign new_n46678_ = ~new_n46675_ & new_n46677_;
  assign new_n46679_ = ~new_n46674_ & ~new_n46678_;
  assign new_n46680_ = pi0580 & ~new_n46679_;
  assign new_n46681_ = ~new_n46672_ & ~new_n46680_;
  assign new_n46682_ = ~pi0552 & new_n46681_;
  assign new_n46683_ = ~new_n46622_ & ~new_n46674_;
  assign new_n46684_ = pi0552 & new_n46683_;
  assign new_n46685_ = ~pi0247 & ~new_n46684_;
  assign new_n46686_ = ~new_n46682_ & new_n46685_;
  assign new_n46687_ = ~new_n46575_ & ~new_n46686_;
  assign new_n46688_ = ~pi0532 & ~new_n46687_;
  assign new_n46689_ = ~pi0552 & new_n46573_;
  assign new_n46690_ = ~pi0247 & ~new_n46689_;
  assign new_n46691_ = pi0552 & new_n46681_;
  assign new_n46692_ = ~pi0552 & new_n46683_;
  assign new_n46693_ = pi0247 & ~new_n46692_;
  assign new_n46694_ = ~new_n46691_ & new_n46693_;
  assign new_n46695_ = ~new_n46690_ & ~new_n46694_;
  assign new_n46696_ = pi0532 & ~new_n46695_;
  assign new_n46697_ = ~new_n46688_ & ~new_n46696_;
  assign new_n46698_ = ~pi0238 & new_n46697_;
  assign new_n46699_ = ~pi0577 & ~new_n46698_;
  assign new_n46700_ = ~new_n46575_ & ~new_n46690_;
  assign new_n46701_ = pi0238 & new_n46700_;
  assign new_n46702_ = pi0247 & pi0532;
  assign new_n46703_ = ~pi0247 & ~pi0532;
  assign new_n46704_ = ~new_n46702_ & ~new_n46703_;
  assign new_n46705_ = new_n46683_ & ~new_n46704_;
  assign new_n46706_ = ~pi0238 & new_n46705_;
  assign new_n46707_ = pi0577 & ~new_n46706_;
  assign new_n46708_ = ~new_n46701_ & new_n46707_;
  assign new_n46709_ = ~pi0498 & ~new_n46708_;
  assign new_n46710_ = ~new_n46699_ & new_n46709_;
  assign new_n46711_ = pi0238 & new_n46697_;
  assign new_n46712_ = pi0577 & ~new_n46711_;
  assign new_n46713_ = ~pi0238 & new_n46700_;
  assign new_n46714_ = pi0238 & new_n46705_;
  assign new_n46715_ = ~pi0577 & ~new_n46714_;
  assign new_n46716_ = ~new_n46713_ & new_n46715_;
  assign new_n46717_ = pi0498 & ~new_n46716_;
  assign new_n46718_ = ~new_n46712_ & new_n46717_;
  assign new_n46719_ = ~new_n46710_ & ~new_n46718_;
  assign new_n46720_ = ~pi0233 & ~new_n46719_;
  assign new_n46721_ = ~pi0237 & ~new_n46720_;
  assign new_n46722_ = ~new_n46526_ & new_n46721_;
  assign po0750 = ~new_n46306_ & ~new_n46722_;
  assign new_n46724_ = ~pi0806 & new_n45126_;
  assign new_n46725_ = ~pi0332 & ~pi0806;
  assign new_n46726_ = pi0990 & new_n46725_;
  assign new_n46727_ = pi0600 & new_n46726_;
  assign new_n46728_ = ~pi0332 & pi0594;
  assign new_n46729_ = ~new_n46727_ & ~new_n46728_;
  assign po0751 = ~new_n46724_ & ~new_n46729_;
  assign new_n46731_ = pi0605 & ~pi0806;
  assign new_n46732_ = new_n45109_ & new_n46731_;
  assign new_n46733_ = pi0595 & new_n46732_;
  assign new_n46734_ = ~pi0595 & ~new_n46732_;
  assign new_n46735_ = ~pi0332 & ~new_n46734_;
  assign po0752 = ~new_n46733_ & new_n46735_;
  assign new_n46737_ = ~pi0332 & pi0596;
  assign new_n46738_ = pi0595 & new_n45108_;
  assign new_n46739_ = new_n46726_ & new_n46738_;
  assign new_n46740_ = ~new_n46737_ & ~new_n46739_;
  assign new_n46741_ = pi0596 & new_n46739_;
  assign po0753 = ~new_n46740_ & ~new_n46741_;
  assign new_n46743_ = pi0597 & new_n46724_;
  assign new_n46744_ = ~pi0597 & ~new_n46724_;
  assign new_n46745_ = ~pi0332 & ~new_n46744_;
  assign po0754 = ~new_n46743_ & new_n46745_;
  assign new_n46747_ = ~pi0882 & ~po1038;
  assign new_n46748_ = pi0947 & new_n46747_;
  assign new_n46749_ = pi0598 & ~new_n46748_;
  assign new_n46750_ = pi0740 & pi0780;
  assign new_n46751_ = new_n6180_ & new_n46750_;
  assign po0755 = new_n46749_ | new_n46751_;
  assign new_n46753_ = ~pi0332 & pi0599;
  assign new_n46754_ = ~new_n46741_ & ~new_n46753_;
  assign new_n46755_ = pi0599 & new_n46741_;
  assign po0756 = ~new_n46754_ & ~new_n46755_;
  assign new_n46757_ = ~pi0332 & pi0600;
  assign new_n46758_ = ~new_n46726_ & ~new_n46757_;
  assign po0757 = ~new_n46727_ & ~new_n46758_;
  assign new_n46760_ = ~pi0601 & pi0806;
  assign new_n46761_ = ~pi0806 & ~pi0989;
  assign new_n46762_ = ~pi0332 & ~new_n46761_;
  assign po0758 = ~new_n46760_ & new_n46762_;
  assign new_n46764_ = ~pi0230 & pi0602;
  assign new_n46765_ = pi0230 & new_n16914_;
  assign new_n46766_ = ~new_n18010_ & new_n46765_;
  assign new_n46767_ = pi0715 & pi1160;
  assign new_n46768_ = ~pi0715 & ~pi1160;
  assign new_n46769_ = pi0790 & ~new_n46768_;
  assign new_n46770_ = ~new_n46767_ & new_n46769_;
  assign new_n46771_ = ~new_n19188_ & ~new_n19335_;
  assign new_n46772_ = ~new_n46770_ & new_n46771_;
  assign new_n46773_ = new_n46766_ & new_n46772_;
  assign new_n46774_ = new_n19281_ & new_n46773_;
  assign po0759 = new_n46764_ | new_n46774_;
  assign new_n46776_ = ~pi0980 & pi1038;
  assign new_n46777_ = pi1060 & new_n46776_;
  assign new_n46778_ = pi0952 & ~pi1061;
  assign new_n46779_ = new_n46777_ & new_n46778_;
  assign po0897 = pi0832 & new_n46779_;
  assign new_n46781_ = ~pi0603 & ~po0897;
  assign new_n46782_ = pi0832 & ~pi1100;
  assign new_n46783_ = new_n46779_ & new_n46782_;
  assign new_n46784_ = ~pi0966 & ~new_n46783_;
  assign new_n46785_ = ~new_n46781_ & new_n46784_;
  assign new_n46786_ = pi0871 & pi0966;
  assign new_n46787_ = pi0872 & pi0966;
  assign new_n46788_ = ~new_n46786_ & ~new_n46787_;
  assign po0760 = new_n46785_ | ~new_n46788_;
  assign new_n46790_ = pi0823 & new_n16630_;
  assign new_n46791_ = ~pi0779 & new_n46790_;
  assign new_n46792_ = ~pi0299 & pi0983;
  assign new_n46793_ = pi0907 & new_n46792_;
  assign new_n46794_ = pi0604 & ~new_n46793_;
  assign new_n46795_ = ~new_n46790_ & new_n46794_;
  assign po0761 = new_n46791_ | new_n46795_;
  assign new_n46797_ = ~pi0605 & ~new_n46725_;
  assign new_n46798_ = ~pi0332 & ~new_n46731_;
  assign po0762 = ~new_n46797_ & new_n46798_;
  assign new_n46800_ = ~pi0606 & ~po0897;
  assign new_n46801_ = ~pi1104 & po0897;
  assign new_n46802_ = ~new_n46800_ & ~new_n46801_;
  assign new_n46803_ = ~pi0966 & ~new_n46802_;
  assign new_n46804_ = ~pi0837 & pi0966;
  assign po0763 = ~new_n46803_ & ~new_n46804_;
  assign new_n46806_ = ~pi1107 & po0897;
  assign new_n46807_ = ~pi0607 & ~po0897;
  assign new_n46808_ = ~pi0966 & ~new_n46807_;
  assign po0764 = ~new_n46806_ & new_n46808_;
  assign new_n46810_ = ~pi1116 & po0897;
  assign new_n46811_ = ~pi0608 & ~po0897;
  assign new_n46812_ = ~pi0966 & ~new_n46811_;
  assign po0765 = ~new_n46810_ & new_n46812_;
  assign new_n46814_ = ~pi1118 & po0897;
  assign new_n46815_ = ~pi0609 & ~po0897;
  assign new_n46816_ = ~pi0966 & ~new_n46815_;
  assign po0766 = ~new_n46814_ & new_n46816_;
  assign new_n46818_ = ~pi1113 & po0897;
  assign new_n46819_ = ~pi0610 & ~po0897;
  assign new_n46820_ = ~pi0966 & ~new_n46819_;
  assign po0767 = ~new_n46818_ & new_n46820_;
  assign new_n46822_ = ~pi1114 & po0897;
  assign new_n46823_ = ~pi0611 & ~po0897;
  assign new_n46824_ = ~pi0966 & ~new_n46823_;
  assign po0768 = ~new_n46822_ & new_n46824_;
  assign new_n46826_ = ~pi1111 & po0897;
  assign new_n46827_ = ~pi0612 & ~po0897;
  assign new_n46828_ = ~pi0966 & ~new_n46827_;
  assign po0769 = ~new_n46826_ & new_n46828_;
  assign new_n46830_ = ~pi1115 & po0897;
  assign new_n46831_ = ~pi0613 & ~po0897;
  assign new_n46832_ = ~pi0966 & ~new_n46831_;
  assign po0770 = ~new_n46830_ & new_n46832_;
  assign new_n46834_ = ~pi1102 & po0897;
  assign new_n46835_ = ~pi0614 & ~po0897;
  assign new_n46836_ = ~pi0966 & ~new_n46835_;
  assign new_n46837_ = ~new_n46834_ & new_n46836_;
  assign po0771 = new_n46786_ | new_n46837_;
  assign new_n46839_ = pi0907 & new_n46747_;
  assign new_n46840_ = ~pi0615 & ~new_n46839_;
  assign new_n46841_ = pi0779 & pi0797;
  assign new_n46842_ = new_n6183_ & new_n46841_;
  assign po0772 = new_n46840_ | new_n46842_;
  assign new_n46844_ = ~pi1101 & po0897;
  assign new_n46845_ = ~pi0616 & ~po0897;
  assign new_n46846_ = ~pi0966 & ~new_n46845_;
  assign new_n46847_ = ~new_n46844_ & new_n46846_;
  assign po0773 = new_n46787_ | new_n46847_;
  assign new_n46849_ = ~pi0617 & ~po0897;
  assign new_n46850_ = ~pi1105 & po0897;
  assign new_n46851_ = ~new_n46849_ & ~new_n46850_;
  assign new_n46852_ = ~pi0966 & ~new_n46851_;
  assign new_n46853_ = ~pi0850 & pi0966;
  assign po0774 = ~new_n46852_ & ~new_n46853_;
  assign new_n46855_ = ~pi1117 & po0897;
  assign new_n46856_ = ~pi0618 & ~po0897;
  assign new_n46857_ = ~pi0966 & ~new_n46856_;
  assign po0775 = ~new_n46855_ & new_n46857_;
  assign new_n46859_ = ~pi1122 & po0897;
  assign new_n46860_ = ~pi0619 & ~po0897;
  assign new_n46861_ = ~pi0966 & ~new_n46860_;
  assign po0776 = ~new_n46859_ & new_n46861_;
  assign new_n46863_ = ~pi1112 & po0897;
  assign new_n46864_ = ~pi0620 & ~po0897;
  assign new_n46865_ = ~pi0966 & ~new_n46864_;
  assign po0777 = ~new_n46863_ & new_n46865_;
  assign new_n46867_ = ~pi1108 & po0897;
  assign new_n46868_ = ~pi0621 & ~po0897;
  assign new_n46869_ = ~pi0966 & ~new_n46868_;
  assign po0778 = ~new_n46867_ & new_n46869_;
  assign new_n46871_ = ~pi1109 & po0897;
  assign new_n46872_ = ~pi0622 & ~po0897;
  assign new_n46873_ = ~pi0966 & ~new_n46872_;
  assign po0779 = ~new_n46871_ & new_n46873_;
  assign new_n46875_ = ~pi1106 & po0897;
  assign new_n46876_ = ~pi0623 & ~po0897;
  assign new_n46877_ = ~pi0966 & ~new_n46876_;
  assign po0780 = ~new_n46875_ & new_n46877_;
  assign new_n46879_ = pi0831 & new_n16707_;
  assign new_n46880_ = ~pi0780 & new_n46879_;
  assign new_n46881_ = pi0947 & new_n46792_;
  assign new_n46882_ = pi0624 & ~new_n46881_;
  assign new_n46883_ = ~new_n46879_ & new_n46882_;
  assign po0781 = new_n46880_ | new_n46883_;
  assign new_n46885_ = pi0832 & ~pi0973;
  assign new_n46886_ = ~pi1054 & pi1066;
  assign new_n46887_ = pi1088 & new_n46886_;
  assign new_n46888_ = new_n46885_ & new_n46887_;
  assign po0954 = ~pi0953 & new_n46888_;
  assign new_n46890_ = ~pi1116 & po0954;
  assign new_n46891_ = ~pi0625 & ~po0954;
  assign new_n46892_ = ~pi0962 & ~new_n46891_;
  assign po0782 = ~new_n46890_ & new_n46892_;
  assign new_n46894_ = ~pi1121 & po0897;
  assign new_n46895_ = ~pi0626 & ~po0897;
  assign new_n46896_ = ~pi0966 & ~new_n46895_;
  assign po0783 = ~new_n46894_ & new_n46896_;
  assign new_n46898_ = ~pi1117 & po0954;
  assign new_n46899_ = ~pi0627 & ~po0954;
  assign new_n46900_ = ~pi0962 & ~new_n46899_;
  assign po0784 = ~new_n46898_ & new_n46900_;
  assign new_n46902_ = ~pi1119 & po0954;
  assign new_n46903_ = ~pi0628 & ~po0954;
  assign new_n46904_ = ~pi0962 & ~new_n46903_;
  assign po0785 = ~new_n46902_ & new_n46904_;
  assign new_n46906_ = ~pi1119 & po0897;
  assign new_n46907_ = ~pi0629 & ~po0897;
  assign new_n46908_ = ~pi0966 & ~new_n46907_;
  assign po0786 = ~new_n46906_ & new_n46908_;
  assign new_n46910_ = ~pi1120 & po0897;
  assign new_n46911_ = ~pi0630 & ~po0897;
  assign new_n46912_ = ~pi0966 & ~new_n46911_;
  assign po0787 = ~new_n46910_ & new_n46912_;
  assign new_n46914_ = pi0631 & ~po0954;
  assign new_n46915_ = ~pi1113 & po0954;
  assign new_n46916_ = ~pi0962 & ~new_n46915_;
  assign po0788 = ~new_n46914_ & new_n46916_;
  assign new_n46918_ = pi0632 & ~po0954;
  assign new_n46919_ = ~pi1115 & po0954;
  assign new_n46920_ = ~pi0962 & ~new_n46919_;
  assign po0789 = ~new_n46918_ & new_n46920_;
  assign new_n46922_ = ~pi1110 & po0897;
  assign new_n46923_ = ~pi0633 & ~po0897;
  assign new_n46924_ = ~pi0966 & ~new_n46923_;
  assign po0790 = ~new_n46922_ & new_n46924_;
  assign new_n46926_ = ~pi1110 & po0954;
  assign new_n46927_ = ~pi0634 & ~po0954;
  assign new_n46928_ = ~pi0962 & ~new_n46927_;
  assign po0791 = ~new_n46926_ & new_n46928_;
  assign new_n46930_ = pi0635 & ~po0954;
  assign new_n46931_ = ~pi1112 & po0954;
  assign new_n46932_ = ~pi0962 & ~new_n46931_;
  assign po0792 = ~new_n46930_ & new_n46932_;
  assign new_n46934_ = ~pi1127 & po0897;
  assign new_n46935_ = ~pi0636 & ~po0897;
  assign new_n46936_ = ~pi0966 & ~new_n46935_;
  assign po0793 = ~new_n46934_ & new_n46936_;
  assign new_n46938_ = ~pi1105 & po0954;
  assign new_n46939_ = ~pi0637 & ~po0954;
  assign new_n46940_ = ~pi0962 & ~new_n46939_;
  assign po0794 = ~new_n46938_ & new_n46940_;
  assign new_n46942_ = ~pi1107 & po0954;
  assign new_n46943_ = ~pi0638 & ~po0954;
  assign new_n46944_ = ~pi0962 & ~new_n46943_;
  assign po0795 = ~new_n46942_ & new_n46944_;
  assign new_n46946_ = ~pi1109 & po0954;
  assign new_n46947_ = ~pi0639 & ~po0954;
  assign new_n46948_ = ~pi0962 & ~new_n46947_;
  assign po0796 = ~new_n46946_ & new_n46948_;
  assign new_n46950_ = ~pi1128 & po0897;
  assign new_n46951_ = ~pi0640 & ~po0897;
  assign new_n46952_ = ~pi0966 & ~new_n46951_;
  assign po0797 = ~new_n46950_ & new_n46952_;
  assign new_n46954_ = ~pi1121 & po0954;
  assign new_n46955_ = ~pi0641 & ~po0954;
  assign new_n46956_ = ~pi0962 & ~new_n46955_;
  assign po0798 = ~new_n46954_ & new_n46956_;
  assign new_n46958_ = ~pi1103 & po0897;
  assign new_n46959_ = ~pi0642 & ~po0897;
  assign new_n46960_ = ~pi0966 & ~new_n46959_;
  assign po0799 = ~new_n46958_ & new_n46960_;
  assign new_n46962_ = ~pi1104 & po0954;
  assign new_n46963_ = ~pi0643 & ~po0954;
  assign new_n46964_ = ~pi0962 & ~new_n46963_;
  assign po0800 = ~new_n46962_ & new_n46964_;
  assign new_n46966_ = ~pi1123 & po0897;
  assign new_n46967_ = ~pi0644 & ~po0897;
  assign new_n46968_ = ~pi0966 & ~new_n46967_;
  assign po0801 = ~new_n46966_ & new_n46968_;
  assign new_n46970_ = ~pi1125 & po0897;
  assign new_n46971_ = ~pi0645 & ~po0897;
  assign new_n46972_ = ~pi0966 & ~new_n46971_;
  assign po0802 = ~new_n46970_ & new_n46972_;
  assign new_n46974_ = pi0646 & ~po0954;
  assign new_n46975_ = ~pi1114 & po0954;
  assign new_n46976_ = ~pi0962 & ~new_n46975_;
  assign po0803 = ~new_n46974_ & new_n46976_;
  assign new_n46978_ = ~pi1120 & po0954;
  assign new_n46979_ = ~pi0647 & ~po0954;
  assign new_n46980_ = ~pi0962 & ~new_n46979_;
  assign po0804 = ~new_n46978_ & new_n46980_;
  assign new_n46982_ = ~pi1122 & po0954;
  assign new_n46983_ = ~pi0648 & ~po0954;
  assign new_n46984_ = ~pi0962 & ~new_n46983_;
  assign po0805 = ~new_n46982_ & new_n46984_;
  assign new_n46986_ = pi0649 & ~po0954;
  assign new_n46987_ = ~pi1126 & po0954;
  assign new_n46988_ = ~pi0962 & ~new_n46987_;
  assign po0806 = ~new_n46986_ & new_n46988_;
  assign new_n46990_ = pi0650 & ~po0954;
  assign new_n46991_ = ~pi1127 & po0954;
  assign new_n46992_ = ~pi0962 & ~new_n46991_;
  assign po0807 = ~new_n46990_ & new_n46992_;
  assign new_n46994_ = ~pi1130 & po0897;
  assign new_n46995_ = ~pi0651 & ~po0897;
  assign new_n46996_ = ~pi0966 & ~new_n46995_;
  assign po0808 = ~new_n46994_ & new_n46996_;
  assign new_n46998_ = ~pi1131 & po0897;
  assign new_n46999_ = ~pi0652 & ~po0897;
  assign new_n47000_ = ~pi0966 & ~new_n46999_;
  assign po0809 = ~new_n46998_ & new_n47000_;
  assign new_n47002_ = ~pi1129 & po0897;
  assign new_n47003_ = ~pi0653 & ~po0897;
  assign new_n47004_ = ~pi0966 & ~new_n47003_;
  assign po0810 = ~new_n47002_ & new_n47004_;
  assign new_n47006_ = pi0654 & ~po0954;
  assign new_n47007_ = ~pi1130 & po0954;
  assign new_n47008_ = ~pi0962 & ~new_n47007_;
  assign po0811 = ~new_n47006_ & new_n47008_;
  assign new_n47010_ = pi0655 & ~po0954;
  assign new_n47011_ = ~pi1124 & po0954;
  assign new_n47012_ = ~pi0962 & ~new_n47011_;
  assign po0812 = ~new_n47010_ & new_n47012_;
  assign new_n47014_ = ~pi1126 & po0897;
  assign new_n47015_ = ~pi0656 & ~po0897;
  assign new_n47016_ = ~pi0966 & ~new_n47015_;
  assign po0813 = ~new_n47014_ & new_n47016_;
  assign new_n47018_ = pi0657 & ~po0954;
  assign new_n47019_ = ~pi1131 & po0954;
  assign new_n47020_ = ~pi0962 & ~new_n47019_;
  assign po0814 = ~new_n47018_ & new_n47020_;
  assign new_n47022_ = ~pi1124 & po0897;
  assign new_n47023_ = ~pi0658 & ~po0897;
  assign new_n47024_ = ~pi0966 & ~new_n47023_;
  assign po0815 = ~new_n47022_ & new_n47024_;
  assign new_n47026_ = pi0266 & pi0992;
  assign new_n47027_ = ~pi0280 & new_n47026_;
  assign new_n47028_ = ~pi0269 & new_n47027_;
  assign new_n47029_ = ~pi0281 & new_n47028_;
  assign new_n47030_ = ~pi0270 & ~pi0277;
  assign new_n47031_ = ~pi0282 & new_n47030_;
  assign new_n47032_ = new_n47029_ & new_n47031_;
  assign new_n47033_ = ~pi0264 & new_n47032_;
  assign new_n47034_ = ~pi0265 & new_n47033_;
  assign po0959 = ~pi0274 & new_n47034_;
  assign new_n47036_ = pi0274 & ~new_n47034_;
  assign po0816 = ~po0959 & ~new_n47036_;
  assign new_n47038_ = ~pi1118 & po0954;
  assign new_n47039_ = ~pi0660 & ~po0954;
  assign new_n47040_ = ~pi0962 & ~new_n47039_;
  assign po0817 = ~new_n47038_ & new_n47040_;
  assign new_n47042_ = ~pi1101 & po0954;
  assign new_n47043_ = ~pi0661 & ~po0954;
  assign new_n47044_ = ~pi0962 & ~new_n47043_;
  assign po0818 = ~new_n47042_ & new_n47044_;
  assign new_n47046_ = ~pi1102 & po0954;
  assign new_n47047_ = ~pi0662 & ~po0954;
  assign new_n47048_ = ~pi0962 & ~new_n47047_;
  assign po0819 = ~new_n47046_ & new_n47048_;
  assign new_n47050_ = pi0199 & ~pi1065;
  assign new_n47051_ = ~pi0223 & ~pi0224;
  assign new_n47052_ = ~pi0199 & ~pi0257;
  assign new_n47053_ = ~new_n47051_ & ~new_n47052_;
  assign new_n47054_ = ~new_n47050_ & new_n47053_;
  assign new_n47055_ = ~pi0591 & pi0592;
  assign new_n47056_ = pi0365 & new_n47055_;
  assign new_n47057_ = pi0334 & pi0591;
  assign new_n47058_ = ~pi0592 & new_n47057_;
  assign new_n47059_ = ~new_n47056_ & ~new_n47058_;
  assign new_n47060_ = ~pi0590 & ~new_n47059_;
  assign new_n47061_ = pi0590 & ~pi0591;
  assign new_n47062_ = ~pi0592 & new_n47061_;
  assign new_n47063_ = pi0323 & new_n47062_;
  assign new_n47064_ = ~pi0588 & ~new_n47063_;
  assign new_n47065_ = ~new_n47060_ & new_n47064_;
  assign new_n47066_ = ~pi0592 & new_n8598_;
  assign new_n47067_ = pi0464 & new_n47066_;
  assign new_n47068_ = pi0588 & ~new_n47067_;
  assign new_n47069_ = new_n47051_ & ~new_n47068_;
  assign new_n47070_ = ~new_n47065_ & new_n47069_;
  assign new_n47071_ = ~new_n47054_ & ~new_n47070_;
  assign new_n47072_ = new_n8870_ & ~new_n47071_;
  assign new_n47073_ = ~pi1137 & ~pi1138;
  assign new_n47074_ = ~pi1134 & new_n47073_;
  assign new_n47075_ = ~pi0634 & pi1136;
  assign new_n47076_ = ~pi0784 & ~pi1136;
  assign new_n47077_ = pi1135 & ~new_n47076_;
  assign new_n47078_ = ~new_n47075_ & new_n47077_;
  assign new_n47079_ = ~pi0633 & pi1136;
  assign new_n47080_ = ~pi0815 & ~pi1136;
  assign new_n47081_ = ~pi1135 & ~new_n47080_;
  assign new_n47082_ = ~new_n47079_ & new_n47081_;
  assign new_n47083_ = ~new_n47078_ & ~new_n47082_;
  assign new_n47084_ = new_n47074_ & ~new_n47083_;
  assign new_n47085_ = pi1135 & new_n47073_;
  assign new_n47086_ = pi1136 & ~new_n47085_;
  assign new_n47087_ = ~pi0766 & new_n47086_;
  assign new_n47088_ = pi1135 & ~pi1136;
  assign new_n47089_ = pi1134 & new_n47073_;
  assign new_n47090_ = ~new_n47088_ & new_n47089_;
  assign new_n47091_ = ~pi0855 & ~pi1136;
  assign new_n47092_ = ~pi0700 & pi1135;
  assign new_n47093_ = ~new_n47091_ & ~new_n47092_;
  assign new_n47094_ = new_n47090_ & new_n47093_;
  assign new_n47095_ = ~new_n47087_ & new_n47094_;
  assign new_n47096_ = ~new_n47084_ & ~new_n47095_;
  assign new_n47097_ = ~new_n8870_ & ~new_n47096_;
  assign po0820 = new_n47072_ | new_n47097_;
  assign new_n47099_ = ~pi0590 & pi0591;
  assign new_n47100_ = pi0404 & new_n47099_;
  assign new_n47101_ = ~pi0590 & pi0592;
  assign new_n47102_ = ~pi0588 & ~new_n47101_;
  assign new_n47103_ = ~new_n47100_ & new_n47102_;
  assign new_n47104_ = pi0380 & ~pi0591;
  assign new_n47105_ = pi0592 & ~new_n47104_;
  assign new_n47106_ = ~new_n47103_ & ~new_n47105_;
  assign new_n47107_ = pi0355 & new_n47062_;
  assign new_n47108_ = ~new_n47106_ & ~new_n47107_;
  assign new_n47109_ = pi0429 & new_n47066_;
  assign new_n47110_ = pi0588 & ~new_n47109_;
  assign new_n47111_ = new_n47051_ & ~new_n47110_;
  assign new_n47112_ = ~new_n47108_ & new_n47111_;
  assign new_n47113_ = pi0199 & ~pi1084;
  assign new_n47114_ = ~pi0199 & ~pi0292;
  assign new_n47115_ = ~new_n47051_ & ~new_n47114_;
  assign new_n47116_ = ~new_n47113_ & new_n47115_;
  assign new_n47117_ = ~new_n47112_ & ~new_n47116_;
  assign new_n47118_ = new_n8870_ & ~new_n47117_;
  assign new_n47119_ = pi0662 & pi1135;
  assign new_n47120_ = pi0614 & ~pi1135;
  assign new_n47121_ = pi1136 & ~new_n47120_;
  assign new_n47122_ = ~new_n47119_ & new_n47121_;
  assign new_n47123_ = pi0785 & pi1135;
  assign new_n47124_ = pi0811 & ~pi1135;
  assign new_n47125_ = ~pi1136 & ~new_n47124_;
  assign new_n47126_ = ~new_n47123_ & new_n47125_;
  assign new_n47127_ = ~new_n47122_ & ~new_n47126_;
  assign new_n47128_ = ~pi1134 & ~new_n47127_;
  assign new_n47129_ = ~pi0727 & pi1135;
  assign new_n47130_ = ~pi0772 & ~pi1135;
  assign new_n47131_ = pi1136 & ~new_n47130_;
  assign new_n47132_ = ~new_n47129_ & new_n47131_;
  assign new_n47133_ = ~pi1135 & ~pi1136;
  assign new_n47134_ = pi0872 & new_n47133_;
  assign new_n47135_ = pi1134 & ~new_n47134_;
  assign new_n47136_ = ~new_n47132_ & new_n47135_;
  assign new_n47137_ = ~new_n8870_ & new_n47073_;
  assign new_n47138_ = ~new_n47136_ & new_n47137_;
  assign new_n47139_ = ~new_n47128_ & new_n47138_;
  assign po0821 = new_n47118_ | new_n47139_;
  assign new_n47141_ = ~pi1108 & po0954;
  assign new_n47142_ = ~pi0665 & ~po0954;
  assign new_n47143_ = ~pi0962 & ~new_n47142_;
  assign po0822 = ~new_n47141_ & new_n47143_;
  assign new_n47145_ = ~pi0638 & pi1135;
  assign new_n47146_ = ~pi0607 & ~pi1135;
  assign new_n47147_ = pi1136 & ~new_n47146_;
  assign new_n47148_ = ~new_n47145_ & new_n47147_;
  assign new_n47149_ = pi0799 & ~pi1135;
  assign new_n47150_ = ~pi0790 & pi1135;
  assign new_n47151_ = ~pi1136 & ~new_n47150_;
  assign new_n47152_ = ~new_n47149_ & new_n47151_;
  assign new_n47153_ = ~new_n47148_ & ~new_n47152_;
  assign new_n47154_ = new_n47074_ & ~new_n47153_;
  assign new_n47155_ = ~pi0764 & new_n47086_;
  assign new_n47156_ = ~pi0691 & pi1135;
  assign new_n47157_ = ~pi0873 & ~pi1136;
  assign new_n47158_ = ~new_n47156_ & ~new_n47157_;
  assign new_n47159_ = new_n47090_ & new_n47158_;
  assign new_n47160_ = ~new_n47155_ & new_n47159_;
  assign new_n47161_ = ~new_n47154_ & ~new_n47160_;
  assign new_n47162_ = ~new_n8870_ & ~new_n47161_;
  assign new_n47163_ = pi0199 & ~pi1044;
  assign new_n47164_ = ~pi0199 & ~pi0297;
  assign new_n47165_ = ~new_n47051_ & ~new_n47164_;
  assign new_n47166_ = ~new_n47163_ & new_n47165_;
  assign new_n47167_ = pi0456 & new_n47099_;
  assign new_n47168_ = new_n47102_ & ~new_n47167_;
  assign new_n47169_ = pi0337 & ~pi0591;
  assign new_n47170_ = pi0592 & ~new_n47169_;
  assign new_n47171_ = ~new_n47168_ & ~new_n47170_;
  assign new_n47172_ = pi0441 & new_n47062_;
  assign new_n47173_ = ~new_n47171_ & ~new_n47172_;
  assign new_n47174_ = pi0443 & new_n47066_;
  assign new_n47175_ = pi0588 & ~new_n47174_;
  assign new_n47176_ = new_n47051_ & ~new_n47175_;
  assign new_n47177_ = ~new_n47173_ & new_n47176_;
  assign new_n47178_ = ~new_n47166_ & ~new_n47177_;
  assign new_n47179_ = new_n8870_ & ~new_n47178_;
  assign po0823 = new_n47162_ | new_n47179_;
  assign new_n47181_ = pi0319 & new_n47099_;
  assign new_n47182_ = new_n47102_ & ~new_n47181_;
  assign new_n47183_ = pi0338 & ~pi0591;
  assign new_n47184_ = pi0592 & ~new_n47183_;
  assign new_n47185_ = ~new_n47182_ & ~new_n47184_;
  assign new_n47186_ = pi0458 & new_n47062_;
  assign new_n47187_ = ~new_n47185_ & ~new_n47186_;
  assign new_n47188_ = pi0444 & new_n47066_;
  assign new_n47189_ = pi0588 & ~new_n47188_;
  assign new_n47190_ = new_n47051_ & ~new_n47189_;
  assign new_n47191_ = ~new_n47187_ & new_n47190_;
  assign new_n47192_ = pi0199 & ~pi1072;
  assign new_n47193_ = ~pi0199 & ~pi0294;
  assign new_n47194_ = ~new_n47051_ & ~new_n47193_;
  assign new_n47195_ = ~new_n47192_ & new_n47194_;
  assign new_n47196_ = ~new_n47191_ & ~new_n47195_;
  assign new_n47197_ = new_n8870_ & ~new_n47196_;
  assign new_n47198_ = pi0681 & pi1136;
  assign new_n47199_ = pi0792 & ~pi1136;
  assign new_n47200_ = pi1135 & ~new_n47199_;
  assign new_n47201_ = ~new_n47198_ & new_n47200_;
  assign new_n47202_ = pi0642 & pi1136;
  assign new_n47203_ = ~pi0809 & ~pi1136;
  assign new_n47204_ = ~pi1135 & ~new_n47203_;
  assign new_n47205_ = ~new_n47202_ & new_n47204_;
  assign new_n47206_ = ~new_n47201_ & ~new_n47205_;
  assign new_n47207_ = ~pi1134 & ~new_n47206_;
  assign new_n47208_ = ~pi0699 & pi1135;
  assign new_n47209_ = ~pi0763 & ~pi1135;
  assign new_n47210_ = pi1136 & ~new_n47209_;
  assign new_n47211_ = ~new_n47208_ & new_n47210_;
  assign new_n47212_ = pi0871 & new_n47133_;
  assign new_n47213_ = pi1134 & ~new_n47212_;
  assign new_n47214_ = ~new_n47211_ & new_n47213_;
  assign new_n47215_ = new_n47137_ & ~new_n47214_;
  assign new_n47216_ = ~new_n47207_ & new_n47215_;
  assign po0824 = new_n47197_ | new_n47216_;
  assign new_n47218_ = ~pi0680 & pi1135;
  assign new_n47219_ = ~pi0603 & ~pi1135;
  assign new_n47220_ = pi1136 & ~new_n47219_;
  assign new_n47221_ = ~new_n47218_ & new_n47220_;
  assign new_n47222_ = ~pi0778 & pi1135;
  assign new_n47223_ = ~pi0981 & ~pi1135;
  assign new_n47224_ = ~pi1136 & ~new_n47223_;
  assign new_n47225_ = ~new_n47222_ & new_n47224_;
  assign new_n47226_ = ~new_n47221_ & ~new_n47225_;
  assign new_n47227_ = new_n47074_ & ~new_n47226_;
  assign new_n47228_ = ~pi0759 & new_n47086_;
  assign new_n47229_ = ~pi0696 & pi1135;
  assign new_n47230_ = ~pi0837 & ~pi1136;
  assign new_n47231_ = ~new_n47229_ & ~new_n47230_;
  assign new_n47232_ = new_n47090_ & new_n47231_;
  assign new_n47233_ = ~new_n47228_ & new_n47232_;
  assign new_n47234_ = ~new_n47227_ & ~new_n47233_;
  assign new_n47235_ = ~new_n8870_ & ~new_n47234_;
  assign new_n47236_ = pi0199 & ~pi1049;
  assign new_n47237_ = ~pi0199 & ~pi0291;
  assign new_n47238_ = ~new_n47051_ & ~new_n47237_;
  assign new_n47239_ = ~new_n47236_ & new_n47238_;
  assign new_n47240_ = pi0390 & new_n47099_;
  assign new_n47241_ = new_n47102_ & ~new_n47240_;
  assign new_n47242_ = pi0363 & ~pi0591;
  assign new_n47243_ = pi0592 & ~new_n47242_;
  assign new_n47244_ = ~new_n47241_ & ~new_n47243_;
  assign new_n47245_ = pi0342 & new_n47062_;
  assign new_n47246_ = ~new_n47244_ & ~new_n47245_;
  assign new_n47247_ = pi0414 & new_n47066_;
  assign new_n47248_ = pi0588 & ~new_n47247_;
  assign new_n47249_ = new_n47051_ & ~new_n47248_;
  assign new_n47250_ = ~new_n47246_ & new_n47249_;
  assign new_n47251_ = ~new_n47239_ & ~new_n47250_;
  assign new_n47252_ = new_n8870_ & ~new_n47251_;
  assign po0825 = new_n47235_ | new_n47252_;
  assign new_n47254_ = pi0669 & ~po0954;
  assign new_n47255_ = ~pi1125 & po0954;
  assign new_n47256_ = ~pi0962 & ~new_n47255_;
  assign po0826 = ~new_n47254_ & new_n47256_;
  assign new_n47258_ = pi0199 & ~pi1062;
  assign new_n47259_ = ~pi0199 & ~pi0258;
  assign new_n47260_ = ~new_n47051_ & ~new_n47259_;
  assign new_n47261_ = ~new_n47258_ & new_n47260_;
  assign new_n47262_ = pi0364 & new_n47055_;
  assign new_n47263_ = pi0391 & pi0591;
  assign new_n47264_ = ~pi0592 & new_n47263_;
  assign new_n47265_ = ~new_n47262_ & ~new_n47264_;
  assign new_n47266_ = ~pi0590 & ~new_n47265_;
  assign new_n47267_ = pi0343 & new_n47062_;
  assign new_n47268_ = ~pi0588 & ~new_n47267_;
  assign new_n47269_ = ~new_n47266_ & new_n47268_;
  assign new_n47270_ = pi0415 & new_n47066_;
  assign new_n47271_ = pi0588 & ~new_n47270_;
  assign new_n47272_ = new_n47051_ & ~new_n47271_;
  assign new_n47273_ = ~new_n47269_ & new_n47272_;
  assign new_n47274_ = ~new_n47261_ & ~new_n47273_;
  assign new_n47275_ = new_n8870_ & ~new_n47274_;
  assign new_n47276_ = pi0745 & new_n47086_;
  assign new_n47277_ = pi0723 & pi1135;
  assign new_n47278_ = ~pi0852 & ~pi1136;
  assign new_n47279_ = ~new_n47277_ & ~new_n47278_;
  assign new_n47280_ = new_n47090_ & new_n47279_;
  assign new_n47281_ = ~new_n47276_ & new_n47280_;
  assign new_n47282_ = pi1136 & new_n47073_;
  assign new_n47283_ = ~pi0612 & ~pi1135;
  assign new_n47284_ = pi0695 & pi1135;
  assign new_n47285_ = ~pi1134 & ~new_n47284_;
  assign new_n47286_ = ~new_n47283_ & new_n47285_;
  assign new_n47287_ = new_n47282_ & new_n47286_;
  assign new_n47288_ = ~new_n47281_ & ~new_n47287_;
  assign new_n47289_ = ~new_n8870_ & ~new_n47288_;
  assign po0827 = new_n47275_ | new_n47289_;
  assign new_n47291_ = pi0199 & ~pi1040;
  assign new_n47292_ = ~pi0199 & ~pi0261;
  assign new_n47293_ = ~new_n47051_ & ~new_n47292_;
  assign new_n47294_ = ~new_n47291_ & new_n47293_;
  assign new_n47295_ = pi0447 & new_n47055_;
  assign new_n47296_ = pi0333 & pi0591;
  assign new_n47297_ = ~pi0592 & new_n47296_;
  assign new_n47298_ = ~new_n47295_ & ~new_n47297_;
  assign new_n47299_ = ~pi0590 & ~new_n47298_;
  assign new_n47300_ = pi0327 & new_n47062_;
  assign new_n47301_ = ~pi0588 & ~new_n47300_;
  assign new_n47302_ = ~new_n47299_ & new_n47301_;
  assign new_n47303_ = pi0453 & new_n47066_;
  assign new_n47304_ = pi0588 & ~new_n47303_;
  assign new_n47305_ = new_n47051_ & ~new_n47304_;
  assign new_n47306_ = ~new_n47302_ & new_n47305_;
  assign new_n47307_ = ~new_n47294_ & ~new_n47306_;
  assign new_n47308_ = new_n8870_ & ~new_n47307_;
  assign new_n47309_ = pi0741 & new_n47086_;
  assign new_n47310_ = pi0724 & pi1135;
  assign new_n47311_ = ~pi0865 & ~pi1136;
  assign new_n47312_ = ~new_n47310_ & ~new_n47311_;
  assign new_n47313_ = new_n47090_ & new_n47312_;
  assign new_n47314_ = ~new_n47309_ & new_n47313_;
  assign new_n47315_ = ~pi0611 & ~pi1135;
  assign new_n47316_ = pi0646 & pi1135;
  assign new_n47317_ = ~pi1134 & ~new_n47316_;
  assign new_n47318_ = ~new_n47315_ & new_n47317_;
  assign new_n47319_ = new_n47282_ & new_n47318_;
  assign new_n47320_ = ~new_n47314_ & ~new_n47319_;
  assign new_n47321_ = ~new_n8870_ & ~new_n47320_;
  assign po0828 = new_n47308_ | new_n47321_;
  assign new_n47323_ = ~pi0661 & pi1135;
  assign new_n47324_ = ~pi0616 & ~pi1135;
  assign new_n47325_ = pi1136 & ~new_n47324_;
  assign new_n47326_ = ~new_n47323_ & new_n47325_;
  assign new_n47327_ = ~pi0781 & pi1135;
  assign new_n47328_ = ~pi0808 & ~pi1135;
  assign new_n47329_ = ~pi1136 & ~new_n47328_;
  assign new_n47330_ = ~new_n47327_ & new_n47329_;
  assign new_n47331_ = ~new_n47326_ & ~new_n47330_;
  assign new_n47332_ = new_n47074_ & ~new_n47331_;
  assign new_n47333_ = ~pi0758 & new_n47086_;
  assign new_n47334_ = ~pi0736 & pi1135;
  assign new_n47335_ = ~pi0850 & ~pi1136;
  assign new_n47336_ = ~new_n47334_ & ~new_n47335_;
  assign new_n47337_ = new_n47090_ & new_n47336_;
  assign new_n47338_ = ~new_n47333_ & new_n47337_;
  assign new_n47339_ = ~new_n47332_ & ~new_n47338_;
  assign new_n47340_ = ~new_n8870_ & ~new_n47339_;
  assign new_n47341_ = pi0199 & ~pi1048;
  assign new_n47342_ = ~pi0199 & ~pi0290;
  assign new_n47343_ = ~new_n47051_ & ~new_n47342_;
  assign new_n47344_ = ~new_n47341_ & new_n47343_;
  assign new_n47345_ = pi0397 & new_n47099_;
  assign new_n47346_ = new_n47102_ & ~new_n47345_;
  assign new_n47347_ = pi0372 & ~pi0591;
  assign new_n47348_ = pi0592 & ~new_n47347_;
  assign new_n47349_ = ~new_n47346_ & ~new_n47348_;
  assign new_n47350_ = pi0320 & new_n47062_;
  assign new_n47351_ = ~new_n47349_ & ~new_n47350_;
  assign new_n47352_ = pi0422 & new_n47066_;
  assign new_n47353_ = pi0588 & ~new_n47352_;
  assign new_n47354_ = new_n47051_ & ~new_n47353_;
  assign new_n47355_ = ~new_n47351_ & new_n47354_;
  assign new_n47356_ = ~new_n47344_ & ~new_n47355_;
  assign new_n47357_ = new_n8870_ & ~new_n47356_;
  assign po0829 = new_n47340_ | new_n47357_;
  assign new_n47359_ = ~pi0637 & pi1135;
  assign new_n47360_ = ~pi0617 & ~pi1135;
  assign new_n47361_ = pi1136 & ~new_n47360_;
  assign new_n47362_ = ~new_n47359_ & new_n47361_;
  assign new_n47363_ = pi0814 & ~pi1135;
  assign new_n47364_ = ~pi0788 & pi1135;
  assign new_n47365_ = ~pi1136 & ~new_n47364_;
  assign new_n47366_ = ~new_n47363_ & new_n47365_;
  assign new_n47367_ = ~new_n47362_ & ~new_n47366_;
  assign new_n47368_ = new_n47074_ & ~new_n47367_;
  assign new_n47369_ = ~pi0749 & new_n47086_;
  assign new_n47370_ = ~pi0706 & pi1135;
  assign new_n47371_ = ~pi0866 & ~pi1136;
  assign new_n47372_ = ~new_n47370_ & ~new_n47371_;
  assign new_n47373_ = new_n47090_ & new_n47372_;
  assign new_n47374_ = ~new_n47369_ & new_n47373_;
  assign new_n47375_ = ~new_n47368_ & ~new_n47374_;
  assign new_n47376_ = ~new_n8870_ & ~new_n47375_;
  assign new_n47377_ = pi0199 & ~pi1053;
  assign new_n47378_ = ~pi0199 & ~pi0295;
  assign new_n47379_ = ~new_n47051_ & ~new_n47378_;
  assign new_n47380_ = ~new_n47377_ & new_n47379_;
  assign new_n47381_ = pi0411 & new_n47099_;
  assign new_n47382_ = new_n47102_ & ~new_n47381_;
  assign new_n47383_ = pi0387 & ~pi0591;
  assign new_n47384_ = pi0592 & ~new_n47383_;
  assign new_n47385_ = ~new_n47382_ & ~new_n47384_;
  assign new_n47386_ = pi0452 & new_n47062_;
  assign new_n47387_ = ~new_n47385_ & ~new_n47386_;
  assign new_n47388_ = pi0435 & new_n47066_;
  assign new_n47389_ = pi0588 & ~new_n47388_;
  assign new_n47390_ = new_n47051_ & ~new_n47389_;
  assign new_n47391_ = ~new_n47387_ & new_n47390_;
  assign new_n47392_ = ~new_n47380_ & ~new_n47391_;
  assign new_n47393_ = new_n8870_ & ~new_n47392_;
  assign po0830 = new_n47376_ | new_n47393_;
  assign new_n47395_ = pi0199 & ~pi1070;
  assign new_n47396_ = ~pi0199 & ~pi0256;
  assign new_n47397_ = ~new_n47051_ & ~new_n47396_;
  assign new_n47398_ = ~new_n47395_ & new_n47397_;
  assign new_n47399_ = pi0336 & new_n47055_;
  assign new_n47400_ = pi0463 & pi0591;
  assign new_n47401_ = ~pi0592 & new_n47400_;
  assign new_n47402_ = ~new_n47399_ & ~new_n47401_;
  assign new_n47403_ = ~pi0590 & ~new_n47402_;
  assign new_n47404_ = pi0362 & new_n47062_;
  assign new_n47405_ = ~pi0588 & ~new_n47404_;
  assign new_n47406_ = ~new_n47403_ & new_n47405_;
  assign new_n47407_ = pi0437 & new_n47066_;
  assign new_n47408_ = pi0588 & ~new_n47407_;
  assign new_n47409_ = new_n47051_ & ~new_n47408_;
  assign new_n47410_ = ~new_n47406_ & new_n47409_;
  assign new_n47411_ = ~new_n47398_ & ~new_n47410_;
  assign new_n47412_ = new_n8870_ & ~new_n47411_;
  assign new_n47413_ = pi0639 & pi1135;
  assign new_n47414_ = pi0622 & ~pi1135;
  assign new_n47415_ = pi1136 & ~new_n47414_;
  assign new_n47416_ = ~new_n47413_ & new_n47415_;
  assign new_n47417_ = pi0783 & pi1135;
  assign new_n47418_ = pi0804 & ~pi1135;
  assign new_n47419_ = ~pi1136 & ~new_n47418_;
  assign new_n47420_ = ~new_n47417_ & new_n47419_;
  assign new_n47421_ = ~new_n47416_ & ~new_n47420_;
  assign new_n47422_ = ~pi1134 & ~new_n47421_;
  assign new_n47423_ = ~pi0735 & pi1135;
  assign new_n47424_ = ~pi0743 & ~pi1135;
  assign new_n47425_ = pi1136 & ~new_n47424_;
  assign new_n47426_ = ~new_n47423_ & new_n47425_;
  assign new_n47427_ = pi0859 & new_n47133_;
  assign new_n47428_ = pi1134 & ~new_n47427_;
  assign new_n47429_ = ~new_n47426_ & new_n47428_;
  assign new_n47430_ = new_n47137_ & ~new_n47429_;
  assign new_n47431_ = ~new_n47422_ & new_n47430_;
  assign po0831 = new_n47412_ | new_n47431_;
  assign new_n47433_ = pi0876 & new_n47133_;
  assign new_n47434_ = ~pi0730 & pi1135;
  assign new_n47435_ = ~pi0748 & ~pi1135;
  assign new_n47436_ = pi1136 & ~new_n47435_;
  assign new_n47437_ = ~new_n47434_ & new_n47436_;
  assign new_n47438_ = ~new_n47433_ & ~new_n47437_;
  assign new_n47439_ = new_n47089_ & ~new_n47438_;
  assign new_n47440_ = ~pi0710 & pi1135;
  assign new_n47441_ = pi1136 & ~new_n47440_;
  assign new_n47442_ = pi0789 & new_n47088_;
  assign new_n47443_ = ~pi0803 & ~pi1135;
  assign new_n47444_ = ~new_n47442_ & ~new_n47443_;
  assign new_n47445_ = ~new_n47441_ & new_n47444_;
  assign new_n47446_ = ~pi0623 & new_n47086_;
  assign new_n47447_ = new_n47074_ & ~new_n47446_;
  assign new_n47448_ = ~new_n47445_ & new_n47447_;
  assign new_n47449_ = ~new_n47439_ & ~new_n47448_;
  assign new_n47450_ = ~new_n8870_ & ~new_n47449_;
  assign new_n47451_ = pi0199 & ~pi1037;
  assign new_n47452_ = ~pi0199 & ~pi0296;
  assign new_n47453_ = ~new_n47051_ & ~new_n47452_;
  assign new_n47454_ = ~new_n47451_ & new_n47453_;
  assign new_n47455_ = pi0412 & new_n47099_;
  assign new_n47456_ = new_n47102_ & ~new_n47455_;
  assign new_n47457_ = pi0388 & ~pi0591;
  assign new_n47458_ = pi0592 & ~new_n47457_;
  assign new_n47459_ = ~new_n47456_ & ~new_n47458_;
  assign new_n47460_ = pi0455 & new_n47062_;
  assign new_n47461_ = ~new_n47459_ & ~new_n47460_;
  assign new_n47462_ = pi0436 & new_n47066_;
  assign new_n47463_ = pi0588 & ~new_n47462_;
  assign new_n47464_ = new_n47051_ & ~new_n47463_;
  assign new_n47465_ = ~new_n47461_ & new_n47464_;
  assign new_n47466_ = ~new_n47454_ & ~new_n47465_;
  assign new_n47467_ = new_n8870_ & ~new_n47466_;
  assign po0832 = new_n47450_ | new_n47467_;
  assign new_n47469_ = ~pi0643 & pi1135;
  assign new_n47470_ = ~pi0606 & ~pi1135;
  assign new_n47471_ = pi1136 & ~new_n47470_;
  assign new_n47472_ = ~new_n47469_ & new_n47471_;
  assign new_n47473_ = pi0812 & ~pi1135;
  assign new_n47474_ = ~pi0787 & pi1135;
  assign new_n47475_ = ~pi1136 & ~new_n47474_;
  assign new_n47476_ = ~new_n47473_ & new_n47475_;
  assign new_n47477_ = ~new_n47472_ & ~new_n47476_;
  assign new_n47478_ = new_n47074_ & ~new_n47477_;
  assign new_n47479_ = ~pi0746 & new_n47086_;
  assign new_n47480_ = ~pi0729 & pi1135;
  assign new_n47481_ = ~pi0881 & ~pi1136;
  assign new_n47482_ = ~new_n47480_ & ~new_n47481_;
  assign new_n47483_ = new_n47090_ & new_n47482_;
  assign new_n47484_ = ~new_n47479_ & new_n47483_;
  assign new_n47485_ = ~new_n47478_ & ~new_n47484_;
  assign new_n47486_ = ~new_n8870_ & ~new_n47485_;
  assign new_n47487_ = pi0199 & ~pi1059;
  assign new_n47488_ = ~pi0199 & ~pi0293;
  assign new_n47489_ = ~new_n47051_ & ~new_n47488_;
  assign new_n47490_ = ~new_n47487_ & new_n47489_;
  assign new_n47491_ = pi0410 & new_n47099_;
  assign new_n47492_ = new_n47102_ & ~new_n47491_;
  assign new_n47493_ = pi0386 & ~pi0591;
  assign new_n47494_ = pi0592 & ~new_n47493_;
  assign new_n47495_ = ~new_n47492_ & ~new_n47494_;
  assign new_n47496_ = pi0361 & new_n47062_;
  assign new_n47497_ = ~new_n47495_ & ~new_n47496_;
  assign new_n47498_ = pi0434 & new_n47066_;
  assign new_n47499_ = pi0588 & ~new_n47498_;
  assign new_n47500_ = new_n47051_ & ~new_n47499_;
  assign new_n47501_ = ~new_n47497_ & new_n47500_;
  assign new_n47502_ = ~new_n47490_ & ~new_n47501_;
  assign new_n47503_ = new_n8870_ & ~new_n47502_;
  assign po0833 = new_n47486_ | new_n47503_;
  assign new_n47505_ = pi0199 & ~pi1069;
  assign new_n47506_ = ~pi0199 & ~pi0259;
  assign new_n47507_ = ~new_n47051_ & ~new_n47506_;
  assign new_n47508_ = ~new_n47505_ & new_n47507_;
  assign new_n47509_ = pi0366 & new_n47055_;
  assign new_n47510_ = pi0335 & pi0591;
  assign new_n47511_ = ~pi0592 & new_n47510_;
  assign new_n47512_ = ~new_n47509_ & ~new_n47511_;
  assign new_n47513_ = ~pi0590 & ~new_n47512_;
  assign new_n47514_ = pi0344 & new_n47062_;
  assign new_n47515_ = ~pi0588 & ~new_n47514_;
  assign new_n47516_ = ~new_n47513_ & new_n47515_;
  assign new_n47517_ = pi0416 & new_n47066_;
  assign new_n47518_ = pi0588 & ~new_n47517_;
  assign new_n47519_ = new_n47051_ & ~new_n47518_;
  assign new_n47520_ = ~new_n47516_ & new_n47519_;
  assign new_n47521_ = ~new_n47508_ & ~new_n47520_;
  assign new_n47522_ = new_n8870_ & ~new_n47521_;
  assign new_n47523_ = pi0742 & new_n47086_;
  assign new_n47524_ = pi0704 & pi1135;
  assign new_n47525_ = ~pi0870 & ~pi1136;
  assign new_n47526_ = ~new_n47524_ & ~new_n47525_;
  assign new_n47527_ = new_n47090_ & new_n47526_;
  assign new_n47528_ = ~new_n47523_ & new_n47527_;
  assign new_n47529_ = ~pi0620 & ~pi1135;
  assign new_n47530_ = pi0635 & pi1135;
  assign new_n47531_ = ~pi1134 & ~new_n47530_;
  assign new_n47532_ = ~new_n47529_ & new_n47531_;
  assign new_n47533_ = new_n47282_ & new_n47532_;
  assign new_n47534_ = ~new_n47528_ & ~new_n47533_;
  assign new_n47535_ = ~new_n8870_ & ~new_n47534_;
  assign po0834 = new_n47522_ | new_n47535_;
  assign new_n47537_ = pi0199 & ~pi1067;
  assign new_n47538_ = ~pi0199 & ~pi0260;
  assign new_n47539_ = ~new_n47051_ & ~new_n47538_;
  assign new_n47540_ = ~new_n47537_ & new_n47539_;
  assign new_n47541_ = pi0368 & new_n47055_;
  assign new_n47542_ = pi0393 & pi0591;
  assign new_n47543_ = ~pi0592 & new_n47542_;
  assign new_n47544_ = ~new_n47541_ & ~new_n47543_;
  assign new_n47545_ = ~pi0590 & ~new_n47544_;
  assign new_n47546_ = pi0346 & new_n47062_;
  assign new_n47547_ = ~pi0588 & ~new_n47546_;
  assign new_n47548_ = ~new_n47545_ & new_n47547_;
  assign new_n47549_ = pi0418 & new_n47066_;
  assign new_n47550_ = pi0588 & ~new_n47549_;
  assign new_n47551_ = new_n47051_ & ~new_n47550_;
  assign new_n47552_ = ~new_n47548_ & new_n47551_;
  assign new_n47553_ = ~new_n47540_ & ~new_n47552_;
  assign new_n47554_ = new_n8870_ & ~new_n47553_;
  assign new_n47555_ = pi0760 & new_n47086_;
  assign new_n47556_ = pi0688 & pi1135;
  assign new_n47557_ = ~pi0856 & ~pi1136;
  assign new_n47558_ = ~new_n47556_ & ~new_n47557_;
  assign new_n47559_ = new_n47090_ & new_n47558_;
  assign new_n47560_ = ~new_n47555_ & new_n47559_;
  assign new_n47561_ = ~pi0613 & ~pi1135;
  assign new_n47562_ = pi0632 & pi1135;
  assign new_n47563_ = ~pi1134 & ~new_n47562_;
  assign new_n47564_ = ~new_n47561_ & new_n47563_;
  assign new_n47565_ = new_n47282_ & new_n47564_;
  assign new_n47566_ = ~new_n47560_ & ~new_n47565_;
  assign new_n47567_ = ~new_n8870_ & ~new_n47566_;
  assign po0835 = new_n47554_ | new_n47567_;
  assign new_n47569_ = pi0199 & ~pi1036;
  assign new_n47570_ = ~pi0199 & ~pi0255;
  assign new_n47571_ = ~new_n47051_ & ~new_n47570_;
  assign new_n47572_ = ~new_n47569_ & new_n47571_;
  assign new_n47573_ = pi0389 & new_n47055_;
  assign new_n47574_ = pi0413 & pi0591;
  assign new_n47575_ = ~pi0592 & new_n47574_;
  assign new_n47576_ = ~new_n47573_ & ~new_n47575_;
  assign new_n47577_ = ~pi0590 & ~new_n47576_;
  assign new_n47578_ = pi0450 & new_n47062_;
  assign new_n47579_ = ~pi0588 & ~new_n47578_;
  assign new_n47580_ = ~new_n47577_ & new_n47579_;
  assign new_n47581_ = pi0438 & new_n47066_;
  assign new_n47582_ = pi0588 & ~new_n47581_;
  assign new_n47583_ = new_n47051_ & ~new_n47582_;
  assign new_n47584_ = ~new_n47580_ & new_n47583_;
  assign new_n47585_ = ~new_n47572_ & ~new_n47584_;
  assign new_n47586_ = new_n8870_ & ~new_n47585_;
  assign new_n47587_ = ~pi0665 & pi1136;
  assign new_n47588_ = ~pi0791 & ~pi1136;
  assign new_n47589_ = pi1135 & ~new_n47588_;
  assign new_n47590_ = ~new_n47587_ & new_n47589_;
  assign new_n47591_ = ~pi0621 & pi1136;
  assign new_n47592_ = ~pi0810 & ~pi1136;
  assign new_n47593_ = ~pi1135 & ~new_n47592_;
  assign new_n47594_ = ~new_n47591_ & new_n47593_;
  assign new_n47595_ = ~new_n47590_ & ~new_n47594_;
  assign new_n47596_ = new_n47074_ & ~new_n47595_;
  assign new_n47597_ = ~pi0739 & new_n47086_;
  assign new_n47598_ = ~pi0874 & ~pi1136;
  assign new_n47599_ = ~pi0690 & pi1135;
  assign new_n47600_ = ~new_n47598_ & ~new_n47599_;
  assign new_n47601_ = new_n47090_ & new_n47600_;
  assign new_n47602_ = ~new_n47597_ & new_n47601_;
  assign new_n47603_ = ~new_n47596_ & ~new_n47602_;
  assign new_n47604_ = ~new_n8870_ & ~new_n47603_;
  assign po0836 = new_n47586_ | new_n47604_;
  assign new_n47606_ = ~pi1100 & po0954;
  assign new_n47607_ = ~pi0680 & ~po0954;
  assign new_n47608_ = ~pi0962 & ~new_n47607_;
  assign po0837 = ~new_n47606_ & new_n47608_;
  assign new_n47610_ = ~pi1103 & po0954;
  assign new_n47611_ = ~pi0681 & ~po0954;
  assign new_n47612_ = ~pi0962 & ~new_n47611_;
  assign po0838 = ~new_n47610_ & new_n47612_;
  assign new_n47614_ = pi0199 & ~pi1039;
  assign new_n47615_ = ~pi0199 & ~pi0251;
  assign new_n47616_ = ~new_n47051_ & ~new_n47615_;
  assign new_n47617_ = ~new_n47614_ & new_n47616_;
  assign new_n47618_ = pi0367 & new_n47055_;
  assign new_n47619_ = pi0392 & pi0591;
  assign new_n47620_ = ~pi0592 & new_n47619_;
  assign new_n47621_ = ~new_n47618_ & ~new_n47620_;
  assign new_n47622_ = ~pi0590 & ~new_n47621_;
  assign new_n47623_ = pi0345 & new_n47062_;
  assign new_n47624_ = ~pi0588 & ~new_n47623_;
  assign new_n47625_ = ~new_n47622_ & new_n47624_;
  assign new_n47626_ = pi0417 & new_n47066_;
  assign new_n47627_ = pi0588 & ~new_n47626_;
  assign new_n47628_ = new_n47051_ & ~new_n47627_;
  assign new_n47629_ = ~new_n47625_ & new_n47628_;
  assign new_n47630_ = ~new_n47617_ & ~new_n47629_;
  assign new_n47631_ = new_n8870_ & ~new_n47630_;
  assign new_n47632_ = pi0757 & new_n47086_;
  assign new_n47633_ = pi0686 & pi1135;
  assign new_n47634_ = ~pi0848 & ~pi1136;
  assign new_n47635_ = ~new_n47633_ & ~new_n47634_;
  assign new_n47636_ = new_n47090_ & new_n47635_;
  assign new_n47637_ = ~new_n47632_ & new_n47636_;
  assign new_n47638_ = ~pi0610 & ~pi1135;
  assign new_n47639_ = pi0631 & pi1135;
  assign new_n47640_ = ~pi1134 & ~new_n47639_;
  assign new_n47641_ = ~new_n47638_ & new_n47640_;
  assign new_n47642_ = new_n47282_ & new_n47641_;
  assign new_n47643_ = ~new_n47637_ & ~new_n47642_;
  assign new_n47644_ = ~new_n8870_ & ~new_n47643_;
  assign po0839 = new_n47631_ | new_n47644_;
  assign po0980 = pi0953 & new_n46888_;
  assign new_n47647_ = pi0684 & ~po0980;
  assign new_n47648_ = ~pi1130 & po0980;
  assign new_n47649_ = ~pi0962 & ~new_n47648_;
  assign po0841 = ~new_n47647_ & new_n47649_;
  assign new_n47651_ = pi0590 & ~pi0592;
  assign new_n47652_ = pi0357 & new_n47651_;
  assign new_n47653_ = pi0382 & new_n47101_;
  assign new_n47654_ = ~new_n47652_ & ~new_n47653_;
  assign new_n47655_ = ~pi0591 & ~new_n47654_;
  assign new_n47656_ = pi0406 & ~pi0592;
  assign new_n47657_ = new_n47099_ & new_n47656_;
  assign new_n47658_ = ~new_n47655_ & ~new_n47657_;
  assign new_n47659_ = ~pi0588 & ~new_n47658_;
  assign new_n47660_ = pi0588 & ~pi0590;
  assign new_n47661_ = ~pi0591 & ~pi0592;
  assign new_n47662_ = pi0430 & new_n47661_;
  assign new_n47663_ = new_n47660_ & new_n47662_;
  assign new_n47664_ = ~new_n47659_ & ~new_n47663_;
  assign new_n47665_ = new_n47051_ & ~new_n47664_;
  assign new_n47666_ = pi0199 & ~pi1076;
  assign new_n47667_ = ~new_n47051_ & ~new_n47666_;
  assign new_n47668_ = ~new_n42880_ & new_n47667_;
  assign new_n47669_ = ~new_n47665_ & ~new_n47668_;
  assign new_n47670_ = new_n8870_ & ~new_n47669_;
  assign new_n47671_ = pi0860 & new_n47133_;
  assign new_n47672_ = pi0728 & pi1135;
  assign new_n47673_ = pi0744 & ~pi1135;
  assign new_n47674_ = pi1136 & ~new_n47673_;
  assign new_n47675_ = ~new_n47672_ & new_n47674_;
  assign new_n47676_ = ~new_n47671_ & ~new_n47675_;
  assign new_n47677_ = new_n47089_ & ~new_n47676_;
  assign new_n47678_ = pi1136 & ~new_n47073_;
  assign new_n47679_ = ~pi1134 & ~new_n47678_;
  assign new_n47680_ = pi0657 & pi1135;
  assign new_n47681_ = ~pi0652 & ~pi1135;
  assign new_n47682_ = pi1136 & ~new_n47681_;
  assign new_n47683_ = ~new_n47680_ & new_n47682_;
  assign new_n47684_ = pi0813 & new_n47073_;
  assign new_n47685_ = new_n47133_ & new_n47684_;
  assign new_n47686_ = ~new_n47683_ & ~new_n47685_;
  assign new_n47687_ = new_n47679_ & ~new_n47686_;
  assign new_n47688_ = ~new_n47677_ & ~new_n47687_;
  assign new_n47689_ = ~new_n8870_ & ~new_n47688_;
  assign po0842 = new_n47670_ | new_n47689_;
  assign new_n47691_ = pi0686 & ~po0980;
  assign new_n47692_ = ~pi1113 & po0980;
  assign new_n47693_ = ~pi0962 & ~new_n47692_;
  assign po0843 = ~new_n47691_ & new_n47693_;
  assign new_n47695_ = ~pi1127 & po0980;
  assign new_n47696_ = ~pi0687 & ~po0980;
  assign new_n47697_ = ~pi0962 & ~new_n47696_;
  assign po0844 = ~new_n47695_ & new_n47697_;
  assign new_n47699_ = pi0688 & ~po0980;
  assign new_n47700_ = ~pi1115 & po0980;
  assign new_n47701_ = ~pi0962 & ~new_n47700_;
  assign po0845 = ~new_n47699_ & new_n47701_;
  assign new_n47703_ = pi0351 & new_n47651_;
  assign new_n47704_ = pi0376 & new_n47101_;
  assign new_n47705_ = ~new_n47703_ & ~new_n47704_;
  assign new_n47706_ = ~pi0591 & ~new_n47705_;
  assign new_n47707_ = pi0401 & ~pi0592;
  assign new_n47708_ = new_n47099_ & new_n47707_;
  assign new_n47709_ = ~new_n47706_ & ~new_n47708_;
  assign new_n47710_ = ~pi0588 & ~new_n47709_;
  assign new_n47711_ = pi0426 & new_n47661_;
  assign new_n47712_ = new_n47660_ & new_n47711_;
  assign new_n47713_ = ~new_n47710_ & ~new_n47712_;
  assign new_n47714_ = new_n47051_ & ~new_n47713_;
  assign new_n47715_ = ~pi0199 & new_n42849_;
  assign new_n47716_ = pi0199 & ~pi1079;
  assign new_n47717_ = ~new_n47051_ & ~new_n47716_;
  assign new_n47718_ = ~new_n47715_ & new_n47717_;
  assign new_n47719_ = ~new_n47714_ & ~new_n47718_;
  assign new_n47720_ = new_n8870_ & ~new_n47719_;
  assign new_n47721_ = pi0798 & new_n47133_;
  assign new_n47722_ = pi0655 & pi1135;
  assign new_n47723_ = ~pi0658 & ~pi1135;
  assign new_n47724_ = pi1136 & ~new_n47723_;
  assign new_n47725_ = ~new_n47722_ & new_n47724_;
  assign new_n47726_ = ~new_n47721_ & ~new_n47725_;
  assign new_n47727_ = new_n47074_ & ~new_n47726_;
  assign new_n47728_ = pi0752 & new_n47086_;
  assign new_n47729_ = ~pi0703 & pi1135;
  assign new_n47730_ = ~pi0843 & ~pi1136;
  assign new_n47731_ = ~new_n47729_ & ~new_n47730_;
  assign new_n47732_ = new_n47090_ & new_n47731_;
  assign new_n47733_ = ~new_n47728_ & new_n47732_;
  assign new_n47734_ = ~new_n47727_ & ~new_n47733_;
  assign new_n47735_ = ~new_n8870_ & ~new_n47734_;
  assign po0846 = new_n47720_ | new_n47735_;
  assign new_n47737_ = ~pi1108 & po0980;
  assign new_n47738_ = ~pi0690 & ~po0980;
  assign new_n47739_ = ~pi0962 & ~new_n47738_;
  assign po0847 = ~new_n47737_ & new_n47739_;
  assign new_n47741_ = ~pi1107 & po0980;
  assign new_n47742_ = ~pi0691 & ~po0980;
  assign new_n47743_ = ~pi0962 & ~new_n47742_;
  assign po0848 = ~new_n47741_ & new_n47743_;
  assign new_n47745_ = pi0352 & new_n47651_;
  assign new_n47746_ = pi0317 & new_n47101_;
  assign new_n47747_ = ~new_n47745_ & ~new_n47746_;
  assign new_n47748_ = ~pi0591 & ~new_n47747_;
  assign new_n47749_ = pi0402 & ~pi0592;
  assign new_n47750_ = new_n47099_ & new_n47749_;
  assign new_n47751_ = ~new_n47748_ & ~new_n47750_;
  assign new_n47752_ = ~pi0588 & ~new_n47751_;
  assign new_n47753_ = pi0427 & new_n47661_;
  assign new_n47754_ = new_n47660_ & new_n47753_;
  assign new_n47755_ = ~new_n47752_ & ~new_n47754_;
  assign new_n47756_ = new_n47051_ & ~new_n47755_;
  assign new_n47757_ = ~pi0199 & new_n42861_;
  assign new_n47758_ = pi0199 & ~pi1078;
  assign new_n47759_ = ~new_n47051_ & ~new_n47758_;
  assign new_n47760_ = ~new_n47757_ & new_n47759_;
  assign new_n47761_ = ~new_n47756_ & ~new_n47760_;
  assign new_n47762_ = new_n8870_ & ~new_n47761_;
  assign new_n47763_ = pi0649 & pi1135;
  assign new_n47764_ = ~pi0656 & ~pi1135;
  assign new_n47765_ = pi1136 & ~new_n47764_;
  assign new_n47766_ = ~new_n47763_ & new_n47765_;
  assign new_n47767_ = pi0801 & new_n47133_;
  assign new_n47768_ = ~pi1134 & ~new_n47767_;
  assign new_n47769_ = ~new_n47766_ & new_n47768_;
  assign new_n47770_ = pi0770 & ~pi1135;
  assign new_n47771_ = ~pi0726 & pi1135;
  assign new_n47772_ = pi1136 & ~new_n47771_;
  assign new_n47773_ = ~new_n47770_ & new_n47772_;
  assign new_n47774_ = pi0844 & new_n47133_;
  assign new_n47775_ = pi1134 & ~new_n47774_;
  assign new_n47776_ = ~new_n47773_ & new_n47775_;
  assign new_n47777_ = new_n47137_ & ~new_n47776_;
  assign new_n47778_ = ~new_n47769_ & new_n47777_;
  assign po0849 = new_n47762_ | new_n47778_;
  assign new_n47780_ = pi0693 & ~po0954;
  assign new_n47781_ = ~pi1129 & po0954;
  assign new_n47782_ = ~pi0962 & ~new_n47781_;
  assign po0850 = ~new_n47780_ & new_n47782_;
  assign new_n47784_ = pi0694 & ~po0980;
  assign new_n47785_ = ~pi1128 & po0980;
  assign new_n47786_ = ~pi0962 & ~new_n47785_;
  assign po0851 = ~new_n47784_ & new_n47786_;
  assign new_n47788_ = pi0695 & ~po0954;
  assign new_n47789_ = ~pi1111 & po0954;
  assign new_n47790_ = ~pi0962 & ~new_n47789_;
  assign po0852 = ~new_n47788_ & new_n47790_;
  assign new_n47792_ = ~pi1100 & po0980;
  assign new_n47793_ = ~pi0696 & ~po0980;
  assign new_n47794_ = ~pi0962 & ~new_n47793_;
  assign po0853 = ~new_n47792_ & new_n47794_;
  assign new_n47796_ = pi0697 & ~po0980;
  assign new_n47797_ = ~pi1129 & po0980;
  assign new_n47798_ = ~pi0962 & ~new_n47797_;
  assign po0854 = ~new_n47796_ & new_n47798_;
  assign new_n47800_ = pi0698 & ~po0980;
  assign new_n47801_ = ~pi1116 & po0980;
  assign new_n47802_ = ~pi0962 & ~new_n47801_;
  assign po0855 = ~new_n47800_ & new_n47802_;
  assign new_n47804_ = ~pi1103 & po0980;
  assign new_n47805_ = ~pi0699 & ~po0980;
  assign new_n47806_ = ~pi0962 & ~new_n47805_;
  assign po0856 = ~new_n47804_ & new_n47806_;
  assign new_n47808_ = ~pi1110 & po0980;
  assign new_n47809_ = ~pi0700 & ~po0980;
  assign new_n47810_ = ~pi0962 & ~new_n47809_;
  assign po0857 = ~new_n47808_ & new_n47810_;
  assign new_n47812_ = pi0701 & ~po0980;
  assign new_n47813_ = ~pi1123 & po0980;
  assign new_n47814_ = ~pi0962 & ~new_n47813_;
  assign po0858 = ~new_n47812_ & new_n47814_;
  assign new_n47816_ = pi0702 & ~po0980;
  assign new_n47817_ = ~pi1117 & po0980;
  assign new_n47818_ = ~pi0962 & ~new_n47817_;
  assign po0859 = ~new_n47816_ & new_n47818_;
  assign new_n47820_ = ~pi1124 & po0980;
  assign new_n47821_ = ~pi0703 & ~po0980;
  assign new_n47822_ = ~pi0962 & ~new_n47821_;
  assign po0860 = ~new_n47820_ & new_n47822_;
  assign new_n47824_ = pi0704 & ~po0980;
  assign new_n47825_ = ~pi1112 & po0980;
  assign new_n47826_ = ~pi0962 & ~new_n47825_;
  assign po0861 = ~new_n47824_ & new_n47826_;
  assign new_n47828_ = ~pi1125 & po0980;
  assign new_n47829_ = ~pi0705 & ~po0980;
  assign new_n47830_ = ~pi0962 & ~new_n47829_;
  assign po0862 = ~new_n47828_ & new_n47830_;
  assign new_n47832_ = ~pi1105 & po0980;
  assign new_n47833_ = ~pi0706 & ~po0980;
  assign new_n47834_ = ~pi0962 & ~new_n47833_;
  assign po0863 = ~new_n47832_ & new_n47834_;
  assign new_n47836_ = pi0370 & new_n47055_;
  assign new_n47837_ = pi0395 & pi0591;
  assign new_n47838_ = ~pi0592 & new_n47837_;
  assign new_n47839_ = ~new_n47836_ & ~new_n47838_;
  assign new_n47840_ = ~pi0590 & ~new_n47839_;
  assign new_n47841_ = pi0347 & new_n47062_;
  assign new_n47842_ = ~new_n47840_ & ~new_n47841_;
  assign new_n47843_ = ~pi0588 & new_n47051_;
  assign new_n47844_ = ~new_n47842_ & new_n47843_;
  assign new_n47845_ = ~pi0200 & ~pi0304;
  assign new_n47846_ = pi0200 & ~pi1048;
  assign new_n47847_ = ~new_n47845_ & ~new_n47846_;
  assign new_n47848_ = ~pi0199 & ~new_n47847_;
  assign new_n47849_ = pi0199 & ~pi1055;
  assign new_n47850_ = ~new_n47051_ & ~new_n47849_;
  assign new_n47851_ = ~new_n47848_ & new_n47850_;
  assign new_n47852_ = new_n47051_ & new_n47066_;
  assign new_n47853_ = pi0420 & pi0588;
  assign new_n47854_ = new_n47852_ & new_n47853_;
  assign new_n47855_ = ~new_n47851_ & ~new_n47854_;
  assign new_n47856_ = ~new_n47844_ & new_n47855_;
  assign new_n47857_ = new_n8870_ & ~new_n47856_;
  assign new_n47858_ = ~pi0618 & ~pi1135;
  assign new_n47859_ = ~pi0627 & pi1135;
  assign new_n47860_ = ~pi1134 & ~new_n47859_;
  assign new_n47861_ = ~new_n47858_ & new_n47860_;
  assign new_n47862_ = new_n47282_ & new_n47861_;
  assign new_n47863_ = pi0753 & new_n47086_;
  assign new_n47864_ = pi0702 & pi1135;
  assign new_n47865_ = ~pi0847 & ~pi1136;
  assign new_n47866_ = ~new_n47864_ & ~new_n47865_;
  assign new_n47867_ = new_n47090_ & new_n47866_;
  assign new_n47868_ = ~new_n47863_ & new_n47867_;
  assign new_n47869_ = ~new_n47862_ & ~new_n47868_;
  assign new_n47870_ = ~new_n8870_ & ~new_n47869_;
  assign po0864 = new_n47857_ | new_n47870_;
  assign new_n47872_ = new_n47051_ & new_n47055_;
  assign new_n47873_ = pi0442 & new_n47872_;
  assign new_n47874_ = ~pi0592 & new_n47051_;
  assign new_n47875_ = pi0328 & pi0591;
  assign new_n47876_ = new_n47874_ & new_n47875_;
  assign new_n47877_ = ~new_n47873_ & ~new_n47876_;
  assign new_n47878_ = ~pi0590 & ~new_n47877_;
  assign new_n47879_ = pi0321 & new_n47051_;
  assign new_n47880_ = new_n47062_ & new_n47879_;
  assign new_n47881_ = ~new_n47878_ & ~new_n47880_;
  assign new_n47882_ = ~pi0588 & ~new_n47881_;
  assign new_n47883_ = ~pi0200 & ~pi0305;
  assign new_n47884_ = pi0200 & ~pi1084;
  assign new_n47885_ = ~new_n47883_ & ~new_n47884_;
  assign new_n47886_ = ~pi0199 & ~new_n47885_;
  assign new_n47887_ = pi0199 & ~pi1058;
  assign new_n47888_ = ~new_n47051_ & ~new_n47887_;
  assign new_n47889_ = ~new_n47886_ & new_n47888_;
  assign new_n47890_ = new_n47051_ & new_n47661_;
  assign new_n47891_ = pi0459 & new_n47660_;
  assign new_n47892_ = new_n47890_ & new_n47891_;
  assign new_n47893_ = new_n8870_ & ~new_n47892_;
  assign new_n47894_ = ~new_n47889_ & new_n47893_;
  assign new_n47895_ = ~new_n47882_ & new_n47894_;
  assign new_n47896_ = pi0754 & new_n47086_;
  assign new_n47897_ = new_n47073_ & ~new_n47088_;
  assign new_n47898_ = ~pi0857 & ~pi1136;
  assign new_n47899_ = pi0709 & pi1135;
  assign new_n47900_ = pi1134 & ~new_n47899_;
  assign new_n47901_ = ~new_n47898_ & new_n47900_;
  assign new_n47902_ = new_n47897_ & new_n47901_;
  assign new_n47903_ = ~new_n47896_ & new_n47902_;
  assign new_n47904_ = ~pi0660 & pi1135;
  assign new_n47905_ = ~pi0609 & ~pi1135;
  assign new_n47906_ = ~pi1134 & ~new_n47905_;
  assign new_n47907_ = ~new_n47904_ & new_n47906_;
  assign new_n47908_ = new_n47282_ & new_n47907_;
  assign new_n47909_ = ~new_n8870_ & ~new_n47908_;
  assign new_n47910_ = ~new_n47903_ & new_n47909_;
  assign po0865 = ~new_n47895_ & ~new_n47910_;
  assign new_n47912_ = pi0709 & ~po0980;
  assign new_n47913_ = ~pi1118 & po0980;
  assign new_n47914_ = ~pi0962 & ~new_n47913_;
  assign po0866 = ~new_n47912_ & new_n47914_;
  assign new_n47916_ = ~pi1106 & po0954;
  assign new_n47917_ = ~pi0710 & ~po0954;
  assign new_n47918_ = ~pi0962 & ~new_n47917_;
  assign po0867 = ~new_n47916_ & new_n47918_;
  assign new_n47920_ = pi0373 & new_n47055_;
  assign new_n47921_ = pi0398 & pi0591;
  assign new_n47922_ = ~pi0592 & new_n47921_;
  assign new_n47923_ = ~new_n47920_ & ~new_n47922_;
  assign new_n47924_ = ~pi0590 & ~new_n47923_;
  assign new_n47925_ = pi0348 & new_n47062_;
  assign new_n47926_ = ~new_n47924_ & ~new_n47925_;
  assign new_n47927_ = new_n47843_ & ~new_n47926_;
  assign new_n47928_ = ~pi0200 & ~pi0306;
  assign new_n47929_ = pi0200 & ~pi1059;
  assign new_n47930_ = ~new_n47928_ & ~new_n47929_;
  assign new_n47931_ = ~pi0199 & ~new_n47930_;
  assign new_n47932_ = pi0199 & ~pi1087;
  assign new_n47933_ = ~new_n47051_ & ~new_n47932_;
  assign new_n47934_ = ~new_n47931_ & new_n47933_;
  assign new_n47935_ = pi0423 & pi0588;
  assign new_n47936_ = new_n47852_ & new_n47935_;
  assign new_n47937_ = ~new_n47934_ & ~new_n47936_;
  assign new_n47938_ = ~new_n47927_ & new_n47937_;
  assign new_n47939_ = new_n8870_ & ~new_n47938_;
  assign new_n47940_ = ~pi0630 & ~pi1135;
  assign new_n47941_ = ~pi0647 & pi1135;
  assign new_n47942_ = ~pi1134 & ~new_n47941_;
  assign new_n47943_ = ~new_n47940_ & new_n47942_;
  assign new_n47944_ = new_n47282_ & new_n47943_;
  assign new_n47945_ = pi0755 & new_n47086_;
  assign new_n47946_ = pi0725 & pi1135;
  assign new_n47947_ = ~pi0858 & ~pi1136;
  assign new_n47948_ = ~new_n47946_ & ~new_n47947_;
  assign new_n47949_ = new_n47090_ & new_n47948_;
  assign new_n47950_ = ~new_n47945_ & new_n47949_;
  assign new_n47951_ = ~new_n47944_ & ~new_n47950_;
  assign new_n47952_ = ~new_n8870_ & ~new_n47951_;
  assign po0868 = new_n47939_ | new_n47952_;
  assign new_n47954_ = pi0751 & new_n47086_;
  assign new_n47955_ = ~pi0842 & ~pi1136;
  assign new_n47956_ = pi0701 & pi1135;
  assign new_n47957_ = pi1134 & ~new_n47956_;
  assign new_n47958_ = ~new_n47955_ & new_n47957_;
  assign new_n47959_ = new_n47897_ & new_n47958_;
  assign new_n47960_ = ~new_n47954_ & new_n47959_;
  assign new_n47961_ = ~pi0644 & ~pi1135;
  assign new_n47962_ = ~pi0715 & pi1135;
  assign new_n47963_ = ~pi1134 & ~new_n47962_;
  assign new_n47964_ = ~new_n47961_ & new_n47963_;
  assign new_n47965_ = new_n47282_ & new_n47964_;
  assign new_n47966_ = ~new_n47960_ & ~new_n47965_;
  assign new_n47967_ = ~new_n8870_ & ~new_n47966_;
  assign new_n47968_ = pi0374 & new_n47055_;
  assign new_n47969_ = pi0400 & pi0591;
  assign new_n47970_ = ~pi0592 & new_n47969_;
  assign new_n47971_ = ~new_n47968_ & ~new_n47970_;
  assign new_n47972_ = ~pi0590 & ~new_n47971_;
  assign new_n47973_ = pi0350 & new_n47062_;
  assign new_n47974_ = ~new_n47972_ & ~new_n47973_;
  assign new_n47975_ = ~pi0588 & ~new_n47974_;
  assign new_n47976_ = pi0425 & new_n47661_;
  assign new_n47977_ = new_n47660_ & new_n47976_;
  assign new_n47978_ = new_n47051_ & ~new_n47977_;
  assign new_n47979_ = ~new_n47975_ & new_n47978_;
  assign new_n47980_ = pi1044 & new_n11444_;
  assign new_n47981_ = pi0298 & new_n10817_;
  assign new_n47982_ = pi0199 & pi1035;
  assign new_n47983_ = ~new_n47051_ & ~new_n47982_;
  assign new_n47984_ = ~new_n47981_ & new_n47983_;
  assign new_n47985_ = ~new_n47980_ & new_n47984_;
  assign new_n47986_ = new_n8870_ & ~new_n47985_;
  assign new_n47987_ = ~new_n47979_ & new_n47986_;
  assign po0869 = new_n47967_ | new_n47987_;
  assign new_n47989_ = pi0371 & new_n47055_;
  assign new_n47990_ = pi0396 & pi0591;
  assign new_n47991_ = ~pi0592 & new_n47990_;
  assign new_n47992_ = ~new_n47989_ & ~new_n47991_;
  assign new_n47993_ = ~pi0590 & ~new_n47992_;
  assign new_n47994_ = pi0322 & new_n47062_;
  assign new_n47995_ = ~new_n47993_ & ~new_n47994_;
  assign new_n47996_ = new_n47843_ & ~new_n47995_;
  assign new_n47997_ = ~pi0200 & ~pi0309;
  assign new_n47998_ = pi0200 & ~pi1072;
  assign new_n47999_ = ~new_n47997_ & ~new_n47998_;
  assign new_n48000_ = ~pi0199 & ~new_n47999_;
  assign new_n48001_ = pi0199 & ~pi1051;
  assign new_n48002_ = ~new_n47051_ & ~new_n48001_;
  assign new_n48003_ = ~new_n48000_ & new_n48002_;
  assign new_n48004_ = pi0421 & pi0588;
  assign new_n48005_ = new_n47852_ & new_n48004_;
  assign new_n48006_ = ~new_n48003_ & ~new_n48005_;
  assign new_n48007_ = ~new_n47996_ & new_n48006_;
  assign new_n48008_ = new_n8870_ & ~new_n48007_;
  assign new_n48009_ = ~pi0629 & ~pi1135;
  assign new_n48010_ = ~pi0628 & pi1135;
  assign new_n48011_ = ~pi1134 & ~new_n48010_;
  assign new_n48012_ = ~new_n48009_ & new_n48011_;
  assign new_n48013_ = new_n47282_ & new_n48012_;
  assign new_n48014_ = pi0756 & new_n47086_;
  assign new_n48015_ = pi0734 & pi1135;
  assign new_n48016_ = ~pi0854 & ~pi1136;
  assign new_n48017_ = ~new_n48015_ & ~new_n48016_;
  assign new_n48018_ = new_n47090_ & new_n48017_;
  assign new_n48019_ = ~new_n48014_ & new_n48018_;
  assign new_n48020_ = ~new_n48013_ & ~new_n48019_;
  assign new_n48021_ = ~new_n8870_ & ~new_n48020_;
  assign po0870 = new_n48008_ | new_n48021_;
  assign new_n48023_ = pi0461 & new_n47651_;
  assign new_n48024_ = pi0439 & new_n47101_;
  assign new_n48025_ = ~new_n48023_ & ~new_n48024_;
  assign new_n48026_ = ~pi0591 & ~new_n48025_;
  assign new_n48027_ = pi0326 & ~pi0592;
  assign new_n48028_ = new_n47099_ & new_n48027_;
  assign new_n48029_ = ~new_n48026_ & ~new_n48028_;
  assign new_n48030_ = ~pi0588 & ~new_n48029_;
  assign new_n48031_ = pi0449 & new_n47661_;
  assign new_n48032_ = new_n47660_ & new_n48031_;
  assign new_n48033_ = ~new_n48030_ & ~new_n48032_;
  assign new_n48034_ = new_n47051_ & ~new_n48033_;
  assign new_n48035_ = pi0199 & ~pi1057;
  assign new_n48036_ = ~new_n47051_ & ~new_n48035_;
  assign new_n48037_ = ~new_n42339_ & new_n48036_;
  assign new_n48038_ = ~new_n48034_ & ~new_n48037_;
  assign new_n48039_ = new_n8870_ & ~new_n48038_;
  assign new_n48040_ = pi0867 & new_n47133_;
  assign new_n48041_ = pi0697 & pi1135;
  assign new_n48042_ = pi0762 & ~pi1135;
  assign new_n48043_ = pi1136 & ~new_n48042_;
  assign new_n48044_ = ~new_n48041_ & new_n48043_;
  assign new_n48045_ = ~new_n48040_ & ~new_n48044_;
  assign new_n48046_ = new_n47089_ & ~new_n48045_;
  assign new_n48047_ = pi0693 & pi1135;
  assign new_n48048_ = ~pi0653 & ~pi1135;
  assign new_n48049_ = pi1136 & ~new_n48048_;
  assign new_n48050_ = ~new_n48047_ & new_n48049_;
  assign new_n48051_ = pi0816 & new_n47073_;
  assign new_n48052_ = new_n47133_ & new_n48051_;
  assign new_n48053_ = ~new_n48050_ & ~new_n48052_;
  assign new_n48054_ = new_n47679_ & ~new_n48053_;
  assign new_n48055_ = ~new_n48046_ & ~new_n48054_;
  assign new_n48056_ = ~new_n8870_ & ~new_n48055_;
  assign po0871 = new_n48039_ | new_n48056_;
  assign new_n48058_ = ~pi1123 & po0954;
  assign new_n48059_ = ~pi0715 & ~po0954;
  assign new_n48060_ = ~pi0962 & ~new_n48059_;
  assign po0872 = ~new_n48058_ & new_n48060_;
  assign new_n48062_ = pi0440 & new_n47872_;
  assign new_n48063_ = pi0329 & pi0591;
  assign new_n48064_ = new_n47874_ & new_n48063_;
  assign new_n48065_ = ~new_n48062_ & ~new_n48064_;
  assign new_n48066_ = ~pi0590 & ~new_n48065_;
  assign new_n48067_ = pi0349 & new_n47051_;
  assign new_n48068_ = new_n47062_ & new_n48067_;
  assign new_n48069_ = ~new_n48066_ & ~new_n48068_;
  assign new_n48070_ = ~pi0588 & ~new_n48069_;
  assign new_n48071_ = ~pi0200 & ~pi0307;
  assign new_n48072_ = pi0200 & ~pi1053;
  assign new_n48073_ = ~new_n48071_ & ~new_n48072_;
  assign new_n48074_ = ~pi0199 & ~new_n48073_;
  assign new_n48075_ = pi0199 & ~pi1043;
  assign new_n48076_ = ~new_n47051_ & ~new_n48075_;
  assign new_n48077_ = ~new_n48074_ & new_n48076_;
  assign new_n48078_ = pi0454 & new_n47660_;
  assign new_n48079_ = new_n47890_ & new_n48078_;
  assign new_n48080_ = new_n8870_ & ~new_n48079_;
  assign new_n48081_ = ~new_n48077_ & new_n48080_;
  assign new_n48082_ = ~new_n48070_ & new_n48081_;
  assign new_n48083_ = pi0761 & new_n47086_;
  assign new_n48084_ = ~pi0845 & ~pi1136;
  assign new_n48085_ = pi0738 & pi1135;
  assign new_n48086_ = pi1134 & ~new_n48085_;
  assign new_n48087_ = ~new_n48084_ & new_n48086_;
  assign new_n48088_ = new_n47897_ & new_n48087_;
  assign new_n48089_ = ~new_n48083_ & new_n48088_;
  assign new_n48090_ = ~pi0641 & pi1135;
  assign new_n48091_ = ~pi0626 & ~pi1135;
  assign new_n48092_ = ~pi1134 & ~new_n48091_;
  assign new_n48093_ = ~new_n48090_ & new_n48092_;
  assign new_n48094_ = new_n47282_ & new_n48093_;
  assign new_n48095_ = ~new_n8870_ & ~new_n48094_;
  assign new_n48096_ = ~new_n48089_ & new_n48095_;
  assign po0873 = ~new_n48082_ & ~new_n48096_;
  assign new_n48098_ = pi0318 & pi0591;
  assign new_n48099_ = ~pi0592 & new_n48098_;
  assign new_n48100_ = ~pi0591 & new_n7785_;
  assign new_n48101_ = ~new_n48099_ & ~new_n48100_;
  assign new_n48102_ = ~pi0590 & ~new_n48101_;
  assign new_n48103_ = pi0462 & new_n47062_;
  assign new_n48104_ = ~new_n48102_ & ~new_n48103_;
  assign new_n48105_ = new_n47843_ & ~new_n48104_;
  assign new_n48106_ = ~pi0199 & new_n42855_;
  assign new_n48107_ = pi0199 & ~pi1074;
  assign new_n48108_ = ~new_n47051_ & ~new_n48107_;
  assign new_n48109_ = ~new_n48106_ & new_n48108_;
  assign new_n48110_ = pi0448 & pi0588;
  assign new_n48111_ = new_n47852_ & new_n48110_;
  assign new_n48112_ = ~new_n48109_ & ~new_n48111_;
  assign new_n48113_ = ~new_n48105_ & new_n48112_;
  assign new_n48114_ = new_n8870_ & ~new_n48113_;
  assign new_n48115_ = pi0768 & new_n47086_;
  assign new_n48116_ = ~pi0839 & ~pi1136;
  assign new_n48117_ = ~pi0705 & pi1135;
  assign new_n48118_ = pi1134 & ~new_n48117_;
  assign new_n48119_ = ~new_n48116_ & new_n48118_;
  assign new_n48120_ = new_n47897_ & new_n48119_;
  assign new_n48121_ = ~new_n48115_ & new_n48120_;
  assign new_n48122_ = pi0800 & new_n47133_;
  assign new_n48123_ = pi0669 & pi1135;
  assign new_n48124_ = ~pi0645 & ~pi1135;
  assign new_n48125_ = pi1136 & ~new_n48124_;
  assign new_n48126_ = ~new_n48123_ & new_n48125_;
  assign new_n48127_ = ~new_n48122_ & ~new_n48126_;
  assign new_n48128_ = new_n47074_ & ~new_n48127_;
  assign new_n48129_ = ~new_n48121_ & ~new_n48128_;
  assign new_n48130_ = ~new_n8870_ & ~new_n48129_;
  assign po0874 = new_n48114_ | new_n48130_;
  assign new_n48132_ = pi0369 & new_n47872_;
  assign new_n48133_ = pi0394 & pi0591;
  assign new_n48134_ = new_n47874_ & new_n48133_;
  assign new_n48135_ = ~new_n48132_ & ~new_n48134_;
  assign new_n48136_ = ~pi0590 & ~new_n48135_;
  assign new_n48137_ = pi0315 & new_n47051_;
  assign new_n48138_ = new_n47062_ & new_n48137_;
  assign new_n48139_ = ~new_n48136_ & ~new_n48138_;
  assign new_n48140_ = ~pi0588 & ~new_n48139_;
  assign new_n48141_ = ~pi0200 & ~pi0303;
  assign new_n48142_ = pi0200 & ~pi1049;
  assign new_n48143_ = ~new_n48141_ & ~new_n48142_;
  assign new_n48144_ = ~pi0199 & ~new_n48143_;
  assign new_n48145_ = pi0199 & ~pi1080;
  assign new_n48146_ = ~new_n47051_ & ~new_n48145_;
  assign new_n48147_ = ~new_n48144_ & new_n48146_;
  assign new_n48148_ = pi0419 & new_n47660_;
  assign new_n48149_ = new_n47890_ & new_n48148_;
  assign new_n48150_ = new_n8870_ & ~new_n48149_;
  assign new_n48151_ = ~new_n48147_ & new_n48150_;
  assign new_n48152_ = ~new_n48140_ & new_n48151_;
  assign new_n48153_ = pi0767 & new_n47086_;
  assign new_n48154_ = ~pi0853 & ~pi1136;
  assign new_n48155_ = pi0698 & pi1135;
  assign new_n48156_ = pi1134 & ~new_n48155_;
  assign new_n48157_ = ~new_n48154_ & new_n48156_;
  assign new_n48158_ = new_n47897_ & new_n48157_;
  assign new_n48159_ = ~new_n48153_ & new_n48158_;
  assign new_n48160_ = ~pi0625 & pi1135;
  assign new_n48161_ = ~pi0608 & ~pi1135;
  assign new_n48162_ = ~pi1134 & ~new_n48161_;
  assign new_n48163_ = ~new_n48160_ & new_n48162_;
  assign new_n48164_ = new_n47282_ & new_n48163_;
  assign new_n48165_ = ~new_n8870_ & ~new_n48164_;
  assign new_n48166_ = ~new_n48159_ & new_n48165_;
  assign po0875 = ~new_n48152_ & ~new_n48166_;
  assign new_n48168_ = pi0378 & new_n47055_;
  assign new_n48169_ = pi0325 & pi0591;
  assign new_n48170_ = ~pi0592 & new_n48169_;
  assign new_n48171_ = ~new_n48168_ & ~new_n48170_;
  assign new_n48172_ = ~pi0590 & ~new_n48171_;
  assign new_n48173_ = pi0353 & new_n47062_;
  assign new_n48174_ = ~new_n48172_ & ~new_n48173_;
  assign new_n48175_ = new_n47843_ & ~new_n48174_;
  assign new_n48176_ = ~pi0199 & new_n42867_;
  assign new_n48177_ = pi0199 & ~pi1063;
  assign new_n48178_ = ~new_n47051_ & ~new_n48177_;
  assign new_n48179_ = ~new_n48176_ & new_n48178_;
  assign new_n48180_ = pi0451 & pi0588;
  assign new_n48181_ = new_n47852_ & new_n48180_;
  assign new_n48182_ = ~new_n48179_ & ~new_n48181_;
  assign new_n48183_ = ~new_n48175_ & new_n48182_;
  assign new_n48184_ = new_n8870_ & ~new_n48183_;
  assign new_n48185_ = pi0774 & new_n47086_;
  assign new_n48186_ = ~pi0868 & ~pi1136;
  assign new_n48187_ = ~pi0687 & pi1135;
  assign new_n48188_ = pi1134 & ~new_n48187_;
  assign new_n48189_ = ~new_n48186_ & new_n48188_;
  assign new_n48190_ = new_n47897_ & new_n48189_;
  assign new_n48191_ = ~new_n48185_ & new_n48190_;
  assign new_n48192_ = pi0807 & new_n47133_;
  assign new_n48193_ = pi0650 & pi1135;
  assign new_n48194_ = ~pi0636 & ~pi1135;
  assign new_n48195_ = pi1136 & ~new_n48194_;
  assign new_n48196_ = ~new_n48193_ & new_n48195_;
  assign new_n48197_ = ~new_n48192_ & ~new_n48196_;
  assign new_n48198_ = new_n47074_ & ~new_n48197_;
  assign new_n48199_ = ~new_n48191_ & ~new_n48198_;
  assign new_n48200_ = ~new_n8870_ & ~new_n48199_;
  assign po0876 = new_n48184_ | new_n48200_;
  assign new_n48202_ = pi0356 & new_n47651_;
  assign new_n48203_ = pi0381 & new_n47101_;
  assign new_n48204_ = ~new_n48202_ & ~new_n48203_;
  assign new_n48205_ = ~pi0591 & ~new_n48204_;
  assign new_n48206_ = pi0405 & ~pi0592;
  assign new_n48207_ = new_n47099_ & new_n48206_;
  assign new_n48208_ = ~new_n48205_ & ~new_n48207_;
  assign new_n48209_ = ~pi0588 & ~new_n48208_;
  assign new_n48210_ = pi0445 & new_n47661_;
  assign new_n48211_ = new_n47660_ & new_n48210_;
  assign new_n48212_ = ~new_n48209_ & ~new_n48211_;
  assign new_n48213_ = new_n47051_ & ~new_n48212_;
  assign new_n48214_ = pi0199 & ~pi1081;
  assign new_n48215_ = ~new_n47051_ & ~new_n48214_;
  assign new_n48216_ = ~new_n42887_ & new_n48215_;
  assign new_n48217_ = ~new_n48213_ & ~new_n48216_;
  assign new_n48218_ = new_n8870_ & ~new_n48217_;
  assign new_n48219_ = pi0880 & new_n47133_;
  assign new_n48220_ = pi0684 & pi1135;
  assign new_n48221_ = pi0750 & ~pi1135;
  assign new_n48222_ = pi1136 & ~new_n48221_;
  assign new_n48223_ = ~new_n48220_ & new_n48222_;
  assign new_n48224_ = ~new_n48219_ & ~new_n48223_;
  assign new_n48225_ = new_n47089_ & ~new_n48224_;
  assign new_n48226_ = pi0654 & pi1135;
  assign new_n48227_ = ~pi0651 & ~pi1135;
  assign new_n48228_ = pi1136 & ~new_n48227_;
  assign new_n48229_ = ~new_n48226_ & new_n48228_;
  assign new_n48230_ = pi0794 & new_n47073_;
  assign new_n48231_ = new_n47133_ & new_n48230_;
  assign new_n48232_ = ~new_n48229_ & ~new_n48231_;
  assign new_n48233_ = new_n47679_ & ~new_n48232_;
  assign new_n48234_ = ~new_n48225_ & ~new_n48233_;
  assign new_n48235_ = ~new_n8870_ & ~new_n48234_;
  assign po0877 = new_n48218_ | new_n48235_;
  assign new_n48237_ = pi0747 & pi0773;
  assign new_n48238_ = pi0769 & new_n48237_;
  assign new_n48239_ = ~pi0721 & ~new_n48238_;
  assign new_n48240_ = pi0721 & new_n48238_;
  assign new_n48241_ = pi0775 & ~new_n48240_;
  assign new_n48242_ = ~new_n48239_ & new_n48241_;
  assign new_n48243_ = pi0721 & pi0813;
  assign new_n48244_ = ~pi0773 & ~pi0801;
  assign new_n48245_ = pi0773 & pi0801;
  assign new_n48246_ = ~new_n48244_ & ~new_n48245_;
  assign new_n48247_ = ~pi0771 & ~pi0800;
  assign new_n48248_ = pi0771 & pi0800;
  assign new_n48249_ = ~new_n48247_ & ~new_n48248_;
  assign new_n48250_ = ~pi0769 & ~pi0794;
  assign new_n48251_ = pi0769 & pi0794;
  assign new_n48252_ = ~new_n48250_ & ~new_n48251_;
  assign new_n48253_ = ~pi0765 & ~pi0798;
  assign new_n48254_ = pi0765 & pi0798;
  assign new_n48255_ = ~new_n48253_ & ~new_n48254_;
  assign new_n48256_ = pi0807 & ~new_n48255_;
  assign new_n48257_ = pi0747 & new_n48256_;
  assign new_n48258_ = ~pi0747 & ~pi0807;
  assign new_n48259_ = ~new_n48255_ & new_n48258_;
  assign new_n48260_ = ~new_n48257_ & ~new_n48259_;
  assign new_n48261_ = ~new_n48252_ & ~new_n48260_;
  assign new_n48262_ = ~new_n48249_ & new_n48261_;
  assign new_n48263_ = ~new_n48246_ & new_n48262_;
  assign new_n48264_ = new_n48243_ & new_n48263_;
  assign new_n48265_ = ~new_n48249_ & new_n48256_;
  assign new_n48266_ = ~pi0721 & ~pi0813;
  assign new_n48267_ = pi0794 & pi0801;
  assign new_n48268_ = new_n48266_ & new_n48267_;
  assign new_n48269_ = new_n48265_ & new_n48268_;
  assign new_n48270_ = ~new_n48264_ & ~new_n48269_;
  assign new_n48271_ = pi0816 & ~new_n48270_;
  assign new_n48272_ = new_n48242_ & ~new_n48271_;
  assign new_n48273_ = pi0795 & ~new_n48272_;
  assign new_n48274_ = ~pi0945 & pi0988;
  assign new_n48275_ = pi0731 & new_n48274_;
  assign new_n48276_ = pi0721 & ~pi0775;
  assign new_n48277_ = ~new_n48242_ & ~new_n48276_;
  assign new_n48278_ = new_n48275_ & ~new_n48277_;
  assign new_n48279_ = ~new_n48273_ & new_n48278_;
  assign new_n48280_ = ~pi0775 & ~pi0816;
  assign new_n48281_ = pi0775 & pi0816;
  assign new_n48282_ = ~new_n48280_ & ~new_n48281_;
  assign new_n48283_ = new_n48264_ & ~new_n48282_;
  assign new_n48284_ = new_n48276_ & ~new_n48283_;
  assign new_n48285_ = ~pi0731 & ~pi0795;
  assign new_n48286_ = pi0731 & pi0795;
  assign new_n48287_ = ~new_n48285_ & ~new_n48286_;
  assign new_n48288_ = new_n48283_ & ~new_n48287_;
  assign new_n48289_ = pi0721 & ~new_n48275_;
  assign new_n48290_ = ~new_n48288_ & new_n48289_;
  assign new_n48291_ = ~new_n48284_ & ~new_n48290_;
  assign po0878 = new_n48279_ | ~new_n48291_;
  assign new_n48293_ = pi0379 & new_n47055_;
  assign new_n48294_ = pi0403 & pi0591;
  assign new_n48295_ = ~pi0592 & new_n48294_;
  assign new_n48296_ = ~new_n48293_ & ~new_n48295_;
  assign new_n48297_ = ~pi0590 & ~new_n48296_;
  assign new_n48298_ = pi0354 & new_n47062_;
  assign new_n48299_ = ~new_n48297_ & ~new_n48298_;
  assign new_n48300_ = new_n47843_ & ~new_n48299_;
  assign new_n48301_ = ~pi0199 & new_n42873_;
  assign new_n48302_ = pi0199 & ~pi1045;
  assign new_n48303_ = ~new_n47051_ & ~new_n48302_;
  assign new_n48304_ = ~new_n48301_ & new_n48303_;
  assign new_n48305_ = pi0428 & pi0588;
  assign new_n48306_ = new_n47852_ & new_n48305_;
  assign new_n48307_ = ~new_n48304_ & ~new_n48306_;
  assign new_n48308_ = ~new_n48300_ & new_n48307_;
  assign new_n48309_ = new_n8870_ & ~new_n48308_;
  assign new_n48310_ = ~pi0851 & pi1134;
  assign new_n48311_ = ~pi0795 & ~pi1134;
  assign new_n48312_ = ~pi1136 & ~new_n48311_;
  assign new_n48313_ = ~new_n48310_ & new_n48312_;
  assign new_n48314_ = pi0776 & pi1134;
  assign new_n48315_ = ~pi0640 & ~pi1134;
  assign new_n48316_ = pi1136 & ~new_n48315_;
  assign new_n48317_ = ~new_n48314_ & new_n48316_;
  assign new_n48318_ = ~new_n48313_ & ~new_n48317_;
  assign new_n48319_ = ~pi1135 & ~new_n48318_;
  assign new_n48320_ = pi0732 & ~pi1134;
  assign new_n48321_ = pi0694 & pi1134;
  assign new_n48322_ = pi1135 & pi1136;
  assign new_n48323_ = ~new_n48321_ & new_n48322_;
  assign new_n48324_ = ~new_n48320_ & new_n48323_;
  assign new_n48325_ = ~new_n48319_ & ~new_n48324_;
  assign new_n48326_ = new_n47137_ & ~new_n48325_;
  assign po0879 = new_n48309_ | new_n48326_;
  assign new_n48328_ = pi0723 & ~po0980;
  assign new_n48329_ = ~pi1111 & po0980;
  assign new_n48330_ = ~pi0962 & ~new_n48329_;
  assign po0880 = ~new_n48328_ & new_n48330_;
  assign new_n48332_ = pi0724 & ~po0980;
  assign new_n48333_ = ~pi1114 & po0980;
  assign new_n48334_ = ~pi0962 & ~new_n48333_;
  assign po0881 = ~new_n48332_ & new_n48334_;
  assign new_n48336_ = pi0725 & ~po0980;
  assign new_n48337_ = ~pi1120 & po0980;
  assign new_n48338_ = ~pi0962 & ~new_n48337_;
  assign po0882 = ~new_n48336_ & new_n48338_;
  assign new_n48340_ = ~pi1126 & po0980;
  assign new_n48341_ = ~pi0726 & ~po0980;
  assign new_n48342_ = ~pi0962 & ~new_n48341_;
  assign po0883 = ~new_n48340_ & new_n48342_;
  assign new_n48344_ = ~pi1102 & po0980;
  assign new_n48345_ = ~pi0727 & ~po0980;
  assign new_n48346_ = ~pi0962 & ~new_n48345_;
  assign po0884 = ~new_n48344_ & new_n48346_;
  assign new_n48348_ = pi0728 & ~po0980;
  assign new_n48349_ = ~pi1131 & po0980;
  assign new_n48350_ = ~pi0962 & ~new_n48349_;
  assign po0885 = ~new_n48348_ & new_n48350_;
  assign new_n48352_ = ~pi1104 & po0980;
  assign new_n48353_ = ~pi0729 & ~po0980;
  assign new_n48354_ = ~pi0962 & ~new_n48353_;
  assign po0886 = ~new_n48352_ & new_n48354_;
  assign new_n48356_ = ~pi1106 & po0980;
  assign new_n48357_ = ~pi0730 & ~po0980;
  assign new_n48358_ = ~pi0962 & ~new_n48357_;
  assign po0887 = ~new_n48356_ & new_n48358_;
  assign new_n48360_ = ~new_n48243_ & ~new_n48266_;
  assign new_n48361_ = new_n48263_ & ~new_n48360_;
  assign new_n48362_ = pi0795 & ~new_n48282_;
  assign new_n48363_ = new_n48361_ & new_n48362_;
  assign new_n48364_ = ~new_n48237_ & ~new_n48363_;
  assign new_n48365_ = new_n48275_ & ~new_n48364_;
  assign new_n48366_ = pi0731 & ~new_n48363_;
  assign new_n48367_ = ~new_n48282_ & ~new_n48360_;
  assign new_n48368_ = ~pi0795 & pi0801;
  assign new_n48369_ = ~new_n48252_ & new_n48368_;
  assign new_n48370_ = new_n48367_ & new_n48369_;
  assign new_n48371_ = new_n48265_ & new_n48370_;
  assign new_n48372_ = new_n48237_ & ~new_n48371_;
  assign new_n48373_ = ~pi0731 & ~new_n48372_;
  assign new_n48374_ = new_n48274_ & ~new_n48373_;
  assign new_n48375_ = ~new_n48366_ & ~new_n48374_;
  assign po0888 = ~new_n48365_ & ~new_n48375_;
  assign new_n48377_ = pi0732 & ~po0954;
  assign new_n48378_ = ~pi1128 & po0954;
  assign new_n48379_ = ~pi0962 & ~new_n48378_;
  assign po0889 = ~new_n48377_ & new_n48379_;
  assign new_n48381_ = pi0375 & new_n47872_;
  assign new_n48382_ = pi0399 & pi0591;
  assign new_n48383_ = new_n47874_ & new_n48382_;
  assign new_n48384_ = ~new_n48381_ & ~new_n48383_;
  assign new_n48385_ = ~pi0590 & ~new_n48384_;
  assign new_n48386_ = pi0316 & new_n47051_;
  assign new_n48387_ = new_n47062_ & new_n48386_;
  assign new_n48388_ = ~new_n48385_ & ~new_n48387_;
  assign new_n48389_ = ~pi0588 & ~new_n48388_;
  assign new_n48390_ = ~pi0200 & ~pi0308;
  assign new_n48391_ = pi0200 & ~pi1037;
  assign new_n48392_ = ~new_n48390_ & ~new_n48391_;
  assign new_n48393_ = ~pi0199 & ~new_n48392_;
  assign new_n48394_ = pi0199 & ~pi1047;
  assign new_n48395_ = ~new_n47051_ & ~new_n48394_;
  assign new_n48396_ = ~new_n48393_ & new_n48395_;
  assign new_n48397_ = pi0424 & new_n47660_;
  assign new_n48398_ = new_n47890_ & new_n48397_;
  assign new_n48399_ = new_n8870_ & ~new_n48398_;
  assign new_n48400_ = ~new_n48396_ & new_n48399_;
  assign new_n48401_ = ~new_n48389_ & new_n48400_;
  assign new_n48402_ = pi0777 & new_n47086_;
  assign new_n48403_ = ~pi0838 & ~pi1136;
  assign new_n48404_ = pi0737 & pi1135;
  assign new_n48405_ = pi1134 & ~new_n48404_;
  assign new_n48406_ = ~new_n48403_ & new_n48405_;
  assign new_n48407_ = new_n47897_ & new_n48406_;
  assign new_n48408_ = ~new_n48402_ & new_n48407_;
  assign new_n48409_ = ~pi0648 & pi1135;
  assign new_n48410_ = ~pi0619 & ~pi1135;
  assign new_n48411_ = ~pi1134 & ~new_n48410_;
  assign new_n48412_ = ~new_n48409_ & new_n48411_;
  assign new_n48413_ = new_n47282_ & new_n48412_;
  assign new_n48414_ = ~new_n8870_ & ~new_n48413_;
  assign new_n48415_ = ~new_n48408_ & new_n48414_;
  assign po0890 = ~new_n48401_ & ~new_n48415_;
  assign new_n48417_ = pi0734 & ~po0980;
  assign new_n48418_ = ~pi1119 & po0980;
  assign new_n48419_ = ~pi0962 & ~new_n48418_;
  assign po0891 = ~new_n48417_ & new_n48419_;
  assign new_n48421_ = ~pi1109 & po0980;
  assign new_n48422_ = ~pi0735 & ~po0980;
  assign new_n48423_ = ~pi0962 & ~new_n48422_;
  assign po0892 = ~new_n48421_ & new_n48423_;
  assign new_n48425_ = ~pi1101 & po0980;
  assign new_n48426_ = ~pi0736 & ~po0980;
  assign new_n48427_ = ~pi0962 & ~new_n48426_;
  assign po0893 = ~new_n48425_ & new_n48427_;
  assign new_n48429_ = pi0737 & ~po0980;
  assign new_n48430_ = ~pi1122 & po0980;
  assign new_n48431_ = ~pi0962 & ~new_n48430_;
  assign po0894 = ~new_n48429_ & new_n48431_;
  assign new_n48433_ = pi0738 & ~po0980;
  assign new_n48434_ = ~pi1121 & po0980;
  assign new_n48435_ = ~pi0962 & ~new_n48434_;
  assign po0895 = ~new_n48433_ & new_n48435_;
  assign new_n48437_ = ~pi0952 & ~pi1061;
  assign new_n48438_ = new_n46777_ & new_n48437_;
  assign po0988 = pi0832 & new_n48438_;
  assign new_n48440_ = pi0739 & ~po0988;
  assign new_n48441_ = pi1108 & po0988;
  assign new_n48442_ = ~pi0966 & ~new_n48441_;
  assign po0896 = new_n48440_ | ~new_n48442_;
  assign new_n48444_ = pi1114 & po0988;
  assign new_n48445_ = ~pi0741 & ~po0988;
  assign new_n48446_ = ~pi0966 & ~new_n48445_;
  assign po0898 = new_n48444_ | ~new_n48446_;
  assign new_n48448_ = pi1112 & po0988;
  assign new_n48449_ = ~pi0742 & ~po0988;
  assign new_n48450_ = ~pi0966 & ~new_n48449_;
  assign po0899 = new_n48448_ | ~new_n48450_;
  assign new_n48452_ = pi0743 & ~po0988;
  assign new_n48453_ = pi1109 & po0988;
  assign new_n48454_ = ~pi0966 & ~new_n48453_;
  assign po0900 = new_n48452_ | ~new_n48454_;
  assign new_n48456_ = pi1131 & po0988;
  assign new_n48457_ = ~pi0744 & ~po0988;
  assign new_n48458_ = ~pi0966 & ~new_n48457_;
  assign po0901 = new_n48456_ | ~new_n48458_;
  assign new_n48460_ = pi1111 & po0988;
  assign new_n48461_ = ~pi0745 & ~po0988;
  assign new_n48462_ = ~pi0966 & ~new_n48461_;
  assign po0902 = new_n48460_ | ~new_n48462_;
  assign new_n48464_ = pi0746 & ~po0988;
  assign new_n48465_ = pi1104 & po0988;
  assign new_n48466_ = ~pi0966 & ~new_n48465_;
  assign po0903 = new_n48464_ | ~new_n48466_;
  assign new_n48468_ = pi0801 & new_n48259_;
  assign new_n48469_ = pi0773 & new_n48274_;
  assign new_n48470_ = ~new_n48246_ & ~new_n48469_;
  assign new_n48471_ = new_n48256_ & new_n48470_;
  assign new_n48472_ = ~new_n48468_ & ~new_n48471_;
  assign new_n48473_ = ~new_n48287_ & new_n48367_;
  assign new_n48474_ = ~new_n48249_ & ~new_n48252_;
  assign new_n48475_ = new_n48473_ & new_n48474_;
  assign new_n48476_ = ~new_n48472_ & new_n48475_;
  assign new_n48477_ = ~pi0747 & ~new_n48469_;
  assign new_n48478_ = new_n48237_ & new_n48274_;
  assign new_n48479_ = ~new_n48477_ & ~new_n48478_;
  assign po0904 = ~new_n48476_ & new_n48479_;
  assign new_n48481_ = pi0748 & ~po0988;
  assign new_n48482_ = pi1106 & po0988;
  assign new_n48483_ = ~pi0966 & ~new_n48482_;
  assign po0905 = new_n48481_ | ~new_n48483_;
  assign new_n48485_ = pi0749 & ~po0988;
  assign new_n48486_ = pi1105 & po0988;
  assign new_n48487_ = ~pi0966 & ~new_n48486_;
  assign po0906 = new_n48485_ | ~new_n48487_;
  assign new_n48489_ = pi1130 & po0988;
  assign new_n48490_ = ~pi0750 & ~po0988;
  assign new_n48491_ = ~pi0966 & ~new_n48490_;
  assign po0907 = new_n48489_ | ~new_n48491_;
  assign new_n48493_ = pi1123 & po0988;
  assign new_n48494_ = ~pi0751 & ~po0988;
  assign new_n48495_ = ~pi0966 & ~new_n48494_;
  assign po0908 = new_n48493_ | ~new_n48495_;
  assign new_n48497_ = pi1124 & po0988;
  assign new_n48498_ = ~pi0752 & ~po0988;
  assign new_n48499_ = ~pi0966 & ~new_n48498_;
  assign po0909 = new_n48497_ | ~new_n48499_;
  assign new_n48501_ = pi1117 & po0988;
  assign new_n48502_ = ~pi0753 & ~po0988;
  assign new_n48503_ = ~pi0966 & ~new_n48502_;
  assign po0910 = new_n48501_ | ~new_n48503_;
  assign new_n48505_ = pi1118 & po0988;
  assign new_n48506_ = ~pi0754 & ~po0988;
  assign new_n48507_ = ~pi0966 & ~new_n48506_;
  assign po0911 = new_n48505_ | ~new_n48507_;
  assign new_n48509_ = pi1120 & po0988;
  assign new_n48510_ = ~pi0755 & ~po0988;
  assign new_n48511_ = ~pi0966 & ~new_n48510_;
  assign po0912 = new_n48509_ | ~new_n48511_;
  assign new_n48513_ = pi1119 & po0988;
  assign new_n48514_ = ~pi0756 & ~po0988;
  assign new_n48515_ = ~pi0966 & ~new_n48514_;
  assign po0913 = new_n48513_ | ~new_n48515_;
  assign new_n48517_ = pi1113 & po0988;
  assign new_n48518_ = ~pi0757 & ~po0988;
  assign new_n48519_ = ~pi0966 & ~new_n48518_;
  assign po0914 = new_n48517_ | ~new_n48519_;
  assign new_n48521_ = pi0758 & ~po0988;
  assign new_n48522_ = pi1101 & po0988;
  assign new_n48523_ = ~pi0966 & ~new_n48522_;
  assign po0915 = new_n48521_ | ~new_n48523_;
  assign new_n48525_ = ~pi0759 & ~po0988;
  assign new_n48526_ = new_n46782_ & new_n48438_;
  assign new_n48527_ = ~new_n48525_ & ~new_n48526_;
  assign po0916 = pi0966 | new_n48527_;
  assign new_n48529_ = pi1115 & po0988;
  assign new_n48530_ = ~pi0760 & ~po0988;
  assign new_n48531_ = ~pi0966 & ~new_n48530_;
  assign po0917 = new_n48529_ | ~new_n48531_;
  assign new_n48533_ = pi1121 & po0988;
  assign new_n48534_ = ~pi0761 & ~po0988;
  assign new_n48535_ = ~pi0966 & ~new_n48534_;
  assign po0918 = new_n48533_ | ~new_n48535_;
  assign new_n48537_ = pi1129 & po0988;
  assign new_n48538_ = ~pi0762 & ~po0988;
  assign new_n48539_ = ~pi0966 & ~new_n48538_;
  assign po0919 = new_n48537_ | ~new_n48539_;
  assign new_n48541_ = pi0763 & ~po0988;
  assign new_n48542_ = pi1103 & po0988;
  assign new_n48543_ = ~pi0966 & ~new_n48542_;
  assign po0920 = new_n48541_ | ~new_n48543_;
  assign new_n48545_ = pi0764 & ~po0988;
  assign new_n48546_ = pi1107 & po0988;
  assign new_n48547_ = ~pi0966 & ~new_n48546_;
  assign po0921 = new_n48545_ | ~new_n48547_;
  assign po0978 = new_n48263_ & new_n48473_;
  assign new_n48550_ = pi0765 & ~po0978;
  assign new_n48551_ = pi0945 & ~new_n48550_;
  assign new_n48552_ = ~new_n48264_ & ~new_n48266_;
  assign new_n48553_ = ~pi0765 & ~new_n48248_;
  assign new_n48554_ = ~new_n48251_ & new_n48553_;
  assign new_n48555_ = ~new_n48257_ & new_n48554_;
  assign new_n48556_ = new_n48244_ & ~new_n48555_;
  assign new_n48557_ = ~new_n48245_ & ~new_n48556_;
  assign new_n48558_ = new_n48262_ & ~new_n48557_;
  assign new_n48559_ = ~pi0721 & ~new_n48558_;
  assign new_n48560_ = new_n48280_ & ~new_n48559_;
  assign new_n48561_ = ~new_n48552_ & new_n48560_;
  assign new_n48562_ = new_n48281_ & new_n48361_;
  assign new_n48563_ = ~pi0765 & ~new_n48562_;
  assign new_n48564_ = ~new_n48561_ & new_n48563_;
  assign new_n48565_ = ~pi0795 & ~new_n48564_;
  assign new_n48566_ = ~pi0731 & ~new_n48565_;
  assign new_n48567_ = ~pi0795 & new_n48566_;
  assign new_n48568_ = pi0765 & ~new_n48567_;
  assign new_n48569_ = ~new_n48366_ & ~new_n48566_;
  assign new_n48570_ = ~new_n48568_ & ~new_n48569_;
  assign new_n48571_ = ~pi0945 & ~new_n48570_;
  assign po0922 = ~new_n48551_ & ~new_n48571_;
  assign new_n48573_ = pi0766 & ~po0988;
  assign new_n48574_ = pi1110 & po0988;
  assign new_n48575_ = ~pi0966 & ~new_n48574_;
  assign po0923 = new_n48573_ | ~new_n48575_;
  assign new_n48577_ = pi1116 & po0988;
  assign new_n48578_ = ~pi0767 & ~po0988;
  assign new_n48579_ = ~pi0966 & ~new_n48578_;
  assign po0924 = new_n48577_ | ~new_n48579_;
  assign new_n48581_ = pi1125 & po0988;
  assign new_n48582_ = ~pi0768 & ~po0988;
  assign new_n48583_ = ~pi0966 & ~new_n48582_;
  assign po0925 = new_n48581_ | ~new_n48583_;
  assign new_n48585_ = pi0794 & ~new_n48246_;
  assign new_n48586_ = ~new_n48249_ & new_n48585_;
  assign new_n48587_ = new_n48367_ & new_n48586_;
  assign new_n48588_ = ~new_n48260_ & new_n48587_;
  assign new_n48589_ = ~pi0775 & new_n48588_;
  assign new_n48590_ = ~new_n48562_ & ~new_n48589_;
  assign new_n48591_ = pi0795 & ~new_n48590_;
  assign new_n48592_ = pi0775 & new_n48237_;
  assign new_n48593_ = pi0769 & ~new_n48592_;
  assign new_n48594_ = ~pi0769 & new_n48592_;
  assign new_n48595_ = ~new_n48593_ & ~new_n48594_;
  assign new_n48596_ = new_n48275_ & ~new_n48595_;
  assign new_n48597_ = ~new_n48591_ & new_n48596_;
  assign new_n48598_ = ~new_n48287_ & new_n48588_;
  assign new_n48599_ = pi0769 & ~new_n48275_;
  assign new_n48600_ = ~new_n48598_ & new_n48599_;
  assign po0926 = new_n48597_ | new_n48600_;
  assign new_n48602_ = pi1126 & po0988;
  assign new_n48603_ = ~pi0770 & ~po0988;
  assign new_n48604_ = ~pi0966 & ~new_n48603_;
  assign po0927 = new_n48602_ | ~new_n48604_;
  assign new_n48606_ = ~new_n48281_ & ~new_n48560_;
  assign new_n48607_ = new_n48285_ & ~new_n48606_;
  assign new_n48608_ = ~new_n48282_ & new_n48286_;
  assign new_n48609_ = ~new_n48607_ & ~new_n48608_;
  assign po0963 = new_n48361_ & ~new_n48609_;
  assign new_n48611_ = ~pi0945 & pi0987;
  assign new_n48612_ = ~po0963 & new_n48611_;
  assign new_n48613_ = pi0771 & pi0945;
  assign new_n48614_ = ~po0978 & new_n48613_;
  assign po0928 = new_n48612_ | new_n48614_;
  assign new_n48616_ = pi0772 & ~po0988;
  assign new_n48617_ = pi1102 & po0988;
  assign new_n48618_ = ~pi0966 & ~new_n48617_;
  assign po0929 = new_n48616_ | ~new_n48618_;
  assign new_n48620_ = ~pi0801 & new_n48262_;
  assign new_n48621_ = po0963 & new_n48620_;
  assign new_n48622_ = new_n48274_ & ~new_n48621_;
  assign new_n48623_ = pi0801 & ~new_n48473_;
  assign new_n48624_ = new_n48263_ & ~new_n48623_;
  assign new_n48625_ = pi0773 & ~new_n48624_;
  assign new_n48626_ = ~new_n48622_ & ~new_n48625_;
  assign po0930 = ~new_n48469_ & ~new_n48626_;
  assign new_n48628_ = pi1127 & po0988;
  assign new_n48629_ = ~pi0774 & ~po0988;
  assign new_n48630_ = ~pi0966 & ~new_n48629_;
  assign po0931 = new_n48628_ | ~new_n48630_;
  assign new_n48632_ = pi0775 & ~po0978;
  assign new_n48633_ = pi0731 & ~pi0945;
  assign new_n48634_ = pi0765 & pi0771;
  assign new_n48635_ = new_n48237_ & new_n48634_;
  assign new_n48636_ = pi0795 & pi0800;
  assign new_n48637_ = pi0801 & ~pi0816;
  assign new_n48638_ = new_n48636_ & new_n48637_;
  assign new_n48639_ = ~new_n48360_ & new_n48638_;
  assign new_n48640_ = new_n48261_ & new_n48639_;
  assign new_n48641_ = new_n48635_ & ~new_n48640_;
  assign new_n48642_ = ~pi0775 & ~new_n48641_;
  assign new_n48643_ = new_n48633_ & ~new_n48642_;
  assign new_n48644_ = ~new_n48632_ & ~new_n48643_;
  assign new_n48645_ = ~new_n48363_ & ~new_n48635_;
  assign new_n48646_ = pi0775 & new_n48633_;
  assign new_n48647_ = ~new_n48645_ & new_n48646_;
  assign po0932 = ~new_n48644_ & ~new_n48647_;
  assign new_n48649_ = pi1128 & po0988;
  assign new_n48650_ = ~pi0776 & ~po0988;
  assign new_n48651_ = ~pi0966 & ~new_n48650_;
  assign po0933 = new_n48649_ | ~new_n48651_;
  assign new_n48653_ = pi1122 & po0988;
  assign new_n48654_ = ~pi0777 & ~po0988;
  assign new_n48655_ = ~pi0966 & ~new_n48654_;
  assign po0934 = new_n48653_ | ~new_n48655_;
  assign new_n48657_ = pi0832 & pi0956;
  assign new_n48658_ = ~pi1046 & ~pi1083;
  assign new_n48659_ = pi1085 & new_n48658_;
  assign new_n48660_ = new_n48657_ & new_n48659_;
  assign new_n48661_ = ~pi0968 & new_n48660_;
  assign new_n48662_ = pi0778 & ~new_n48661_;
  assign new_n48663_ = pi1100 & new_n48661_;
  assign po0935 = new_n48662_ | new_n48663_;
  assign po0936 = ~pi0779 | new_n46839_;
  assign po0937 = ~pi0780 | new_n46748_;
  assign new_n48667_ = pi0781 & ~new_n48661_;
  assign new_n48668_ = pi1101 & new_n48661_;
  assign po0938 = new_n48667_ | new_n48668_;
  assign new_n48670_ = ~new_n42343_ & ~new_n46792_;
  assign po0939 = new_n46747_ | ~new_n48670_;
  assign new_n48672_ = pi0783 & ~new_n48661_;
  assign new_n48673_ = pi1109 & new_n48661_;
  assign po0940 = new_n48672_ | new_n48673_;
  assign new_n48675_ = pi0784 & ~new_n48661_;
  assign new_n48676_ = pi1110 & new_n48661_;
  assign po0941 = new_n48675_ | new_n48676_;
  assign new_n48678_ = pi0785 & ~new_n48661_;
  assign new_n48679_ = pi1102 & new_n48661_;
  assign po0942 = new_n48678_ | new_n48679_;
  assign new_n48681_ = pi0024 & ~pi0954;
  assign new_n48682_ = pi0786 & pi0954;
  assign po0943 = ~new_n48681_ & ~new_n48682_;
  assign new_n48684_ = pi0787 & ~new_n48661_;
  assign new_n48685_ = pi1104 & new_n48661_;
  assign po0944 = new_n48684_ | new_n48685_;
  assign new_n48687_ = pi0788 & ~new_n48661_;
  assign new_n48688_ = pi1105 & new_n48661_;
  assign po0945 = new_n48687_ | new_n48688_;
  assign new_n48690_ = pi0789 & ~new_n48661_;
  assign new_n48691_ = pi1106 & new_n48661_;
  assign po0946 = new_n48690_ | new_n48691_;
  assign new_n48693_ = pi0790 & ~new_n48661_;
  assign new_n48694_ = pi1107 & new_n48661_;
  assign po0947 = new_n48693_ | new_n48694_;
  assign new_n48696_ = pi0791 & ~new_n48661_;
  assign new_n48697_ = pi1108 & new_n48661_;
  assign po0948 = new_n48696_ | new_n48697_;
  assign new_n48699_ = pi0792 & ~new_n48661_;
  assign new_n48700_ = pi1103 & new_n48661_;
  assign po0949 = new_n48699_ | new_n48700_;
  assign new_n48702_ = pi0968 & new_n48660_;
  assign new_n48703_ = pi0794 & ~new_n48702_;
  assign new_n48704_ = pi1130 & new_n48702_;
  assign po0951 = new_n48703_ | new_n48704_;
  assign new_n48706_ = pi0795 & ~new_n48702_;
  assign new_n48707_ = pi1128 & new_n48702_;
  assign po0952 = new_n48706_ | new_n48707_;
  assign new_n48709_ = pi0266 & ~pi0269;
  assign new_n48710_ = pi0278 & pi0279;
  assign new_n48711_ = ~pi0280 & new_n48710_;
  assign new_n48712_ = new_n48709_ & new_n48711_;
  assign new_n48713_ = ~pi0281 & new_n48712_;
  assign new_n48714_ = new_n47031_ & new_n48713_;
  assign new_n48715_ = pi0264 & ~new_n48714_;
  assign new_n48716_ = ~pi0264 & new_n48714_;
  assign po0953 = ~new_n48715_ & ~new_n48716_;
  assign new_n48718_ = pi0798 & ~new_n48702_;
  assign new_n48719_ = pi1124 & new_n48702_;
  assign po0955 = new_n48718_ | new_n48719_;
  assign new_n48721_ = pi0799 & ~new_n48702_;
  assign new_n48722_ = ~pi1107 & new_n48702_;
  assign po0956 = ~new_n48721_ & ~new_n48722_;
  assign new_n48724_ = pi0800 & ~new_n48702_;
  assign new_n48725_ = pi1125 & new_n48702_;
  assign po0957 = new_n48724_ | new_n48725_;
  assign new_n48727_ = pi0801 & ~new_n48702_;
  assign new_n48728_ = pi1126 & new_n48702_;
  assign po0958 = new_n48727_ | new_n48728_;
  assign new_n48730_ = pi0803 & ~new_n48702_;
  assign new_n48731_ = ~pi1106 & new_n48702_;
  assign po0960 = ~new_n48730_ & ~new_n48731_;
  assign new_n48733_ = pi0804 & ~new_n48702_;
  assign new_n48734_ = pi1109 & new_n48702_;
  assign po0961 = new_n48733_ | new_n48734_;
  assign new_n48736_ = ~pi0282 & new_n47029_;
  assign new_n48737_ = ~pi0270 & new_n48736_;
  assign new_n48738_ = pi0270 & ~new_n48736_;
  assign po0962 = ~new_n48737_ & ~new_n48738_;
  assign new_n48740_ = pi0807 & ~new_n48702_;
  assign new_n48741_ = pi1127 & new_n48702_;
  assign po0964 = new_n48740_ | new_n48741_;
  assign new_n48743_ = pi0808 & ~new_n48702_;
  assign new_n48744_ = pi1101 & new_n48702_;
  assign po0965 = new_n48743_ | new_n48744_;
  assign new_n48746_ = pi0809 & ~new_n48702_;
  assign new_n48747_ = ~pi1103 & new_n48702_;
  assign po0966 = ~new_n48746_ & ~new_n48747_;
  assign new_n48749_ = pi0810 & ~new_n48702_;
  assign new_n48750_ = pi1108 & new_n48702_;
  assign po0967 = new_n48749_ | new_n48750_;
  assign new_n48752_ = pi0811 & ~new_n48702_;
  assign new_n48753_ = pi1102 & new_n48702_;
  assign po0968 = new_n48752_ | new_n48753_;
  assign new_n48755_ = pi0812 & ~new_n48702_;
  assign new_n48756_ = ~pi1104 & new_n48702_;
  assign po0969 = ~new_n48755_ & ~new_n48756_;
  assign new_n48758_ = pi0813 & ~new_n48702_;
  assign new_n48759_ = pi1131 & new_n48702_;
  assign po0970 = new_n48758_ | new_n48759_;
  assign new_n48761_ = pi0814 & ~new_n48702_;
  assign new_n48762_ = ~pi1105 & new_n48702_;
  assign po0971 = ~new_n48761_ & ~new_n48762_;
  assign new_n48764_ = pi0815 & ~new_n48702_;
  assign new_n48765_ = pi1110 & new_n48702_;
  assign po0972 = new_n48764_ | new_n48765_;
  assign new_n48767_ = pi0816 & ~new_n48702_;
  assign new_n48768_ = pi1129 & new_n48702_;
  assign po0973 = new_n48767_ | new_n48768_;
  assign new_n48770_ = pi0269 & ~new_n47027_;
  assign po0974 = ~new_n47028_ & ~new_n48770_;
  assign new_n48772_ = new_n8870_ & new_n14172_;
  assign po0975 = new_n14025_ | new_n48772_;
  assign new_n48774_ = pi0265 & ~new_n47033_;
  assign po0976 = ~new_n47034_ & ~new_n48774_;
  assign new_n48776_ = pi0277 & ~new_n48737_;
  assign po0977 = ~new_n47032_ & ~new_n48776_;
  assign po0979 = ~pi0811 & ~pi0893;
  assign new_n48779_ = ~pi0982 & ~new_n10068_;
  assign new_n48780_ = new_n7572_ & new_n8870_;
  assign new_n48781_ = ~new_n48779_ & ~new_n48780_;
  assign po0981 = new_n2799_ & ~new_n48781_;
  assign new_n48783_ = pi0123 & new_n3105_;
  assign new_n48784_ = pi1131 & ~new_n48783_;
  assign new_n48785_ = pi1127 & ~new_n48783_;
  assign new_n48786_ = ~new_n48784_ & ~new_n48785_;
  assign new_n48787_ = ~pi0825 & new_n48783_;
  assign new_n48788_ = new_n48786_ & ~new_n48787_;
  assign new_n48789_ = pi1131 & new_n48785_;
  assign new_n48790_ = ~new_n48788_ & ~new_n48789_;
  assign new_n48791_ = pi1124 & ~pi1130;
  assign new_n48792_ = ~pi1124 & pi1130;
  assign new_n48793_ = ~new_n48791_ & ~new_n48792_;
  assign new_n48794_ = ~pi1128 & ~pi1129;
  assign new_n48795_ = pi1128 & pi1129;
  assign new_n48796_ = ~new_n48794_ & ~new_n48795_;
  assign new_n48797_ = ~pi1125 & ~pi1126;
  assign new_n48798_ = pi1125 & pi1126;
  assign new_n48799_ = ~new_n48797_ & ~new_n48798_;
  assign new_n48800_ = new_n48796_ & ~new_n48799_;
  assign new_n48801_ = ~new_n48796_ & new_n48799_;
  assign new_n48802_ = ~new_n48800_ & ~new_n48801_;
  assign new_n48803_ = new_n48793_ & new_n48802_;
  assign new_n48804_ = ~new_n48793_ & ~new_n48802_;
  assign new_n48805_ = ~new_n48803_ & ~new_n48804_;
  assign new_n48806_ = ~new_n48790_ & ~new_n48805_;
  assign new_n48807_ = pi0825 & new_n48783_;
  assign new_n48808_ = new_n48786_ & ~new_n48807_;
  assign new_n48809_ = ~new_n48789_ & new_n48805_;
  assign new_n48810_ = ~new_n48808_ & new_n48809_;
  assign po0982 = ~new_n48806_ & ~new_n48810_;
  assign new_n48812_ = pi1123 & ~new_n48783_;
  assign new_n48813_ = pi1122 & ~new_n48783_;
  assign new_n48814_ = ~new_n48812_ & ~new_n48813_;
  assign new_n48815_ = ~pi0826 & new_n48783_;
  assign new_n48816_ = new_n48814_ & ~new_n48815_;
  assign new_n48817_ = pi1123 & new_n48813_;
  assign new_n48818_ = ~new_n48816_ & ~new_n48817_;
  assign new_n48819_ = pi1118 & ~pi1119;
  assign new_n48820_ = ~pi1118 & pi1119;
  assign new_n48821_ = ~new_n48819_ & ~new_n48820_;
  assign new_n48822_ = ~pi1120 & ~pi1121;
  assign new_n48823_ = pi1120 & pi1121;
  assign new_n48824_ = ~new_n48822_ & ~new_n48823_;
  assign new_n48825_ = ~pi1116 & ~pi1117;
  assign new_n48826_ = pi1116 & pi1117;
  assign new_n48827_ = ~new_n48825_ & ~new_n48826_;
  assign new_n48828_ = new_n48824_ & ~new_n48827_;
  assign new_n48829_ = ~new_n48824_ & new_n48827_;
  assign new_n48830_ = ~new_n48828_ & ~new_n48829_;
  assign new_n48831_ = new_n48821_ & new_n48830_;
  assign new_n48832_ = ~new_n48821_ & ~new_n48830_;
  assign new_n48833_ = ~new_n48831_ & ~new_n48832_;
  assign new_n48834_ = ~new_n48818_ & ~new_n48833_;
  assign new_n48835_ = pi0826 & new_n48783_;
  assign new_n48836_ = new_n48814_ & ~new_n48835_;
  assign new_n48837_ = ~new_n48817_ & new_n48833_;
  assign new_n48838_ = ~new_n48836_ & new_n48837_;
  assign po0983 = ~new_n48834_ & ~new_n48838_;
  assign new_n48840_ = pi1100 & ~new_n48783_;
  assign new_n48841_ = pi1107 & ~new_n48783_;
  assign new_n48842_ = ~new_n48840_ & ~new_n48841_;
  assign new_n48843_ = ~pi0827 & new_n48783_;
  assign new_n48844_ = new_n48842_ & ~new_n48843_;
  assign new_n48845_ = pi1100 & new_n48841_;
  assign new_n48846_ = ~new_n48844_ & ~new_n48845_;
  assign new_n48847_ = pi1103 & ~pi1105;
  assign new_n48848_ = ~pi1103 & pi1105;
  assign new_n48849_ = ~new_n48847_ & ~new_n48848_;
  assign new_n48850_ = ~pi1101 & ~pi1102;
  assign new_n48851_ = pi1101 & pi1102;
  assign new_n48852_ = ~new_n48850_ & ~new_n48851_;
  assign new_n48853_ = ~pi1104 & ~pi1106;
  assign new_n48854_ = pi1104 & pi1106;
  assign new_n48855_ = ~new_n48853_ & ~new_n48854_;
  assign new_n48856_ = new_n48852_ & ~new_n48855_;
  assign new_n48857_ = ~new_n48852_ & new_n48855_;
  assign new_n48858_ = ~new_n48856_ & ~new_n48857_;
  assign new_n48859_ = new_n48849_ & new_n48858_;
  assign new_n48860_ = ~new_n48849_ & ~new_n48858_;
  assign new_n48861_ = ~new_n48859_ & ~new_n48860_;
  assign new_n48862_ = ~new_n48846_ & ~new_n48861_;
  assign new_n48863_ = pi0827 & new_n48783_;
  assign new_n48864_ = new_n48842_ & ~new_n48863_;
  assign new_n48865_ = ~new_n48845_ & new_n48861_;
  assign new_n48866_ = ~new_n48864_ & new_n48865_;
  assign po0984 = ~new_n48862_ & ~new_n48866_;
  assign new_n48868_ = pi1115 & ~new_n48783_;
  assign new_n48869_ = pi1114 & ~new_n48783_;
  assign new_n48870_ = ~new_n48868_ & ~new_n48869_;
  assign new_n48871_ = ~pi0828 & new_n48783_;
  assign new_n48872_ = new_n48870_ & ~new_n48871_;
  assign new_n48873_ = pi1115 & new_n48869_;
  assign new_n48874_ = ~new_n48872_ & ~new_n48873_;
  assign new_n48875_ = pi1110 & ~pi1111;
  assign new_n48876_ = ~pi1110 & pi1111;
  assign new_n48877_ = ~new_n48875_ & ~new_n48876_;
  assign new_n48878_ = ~pi1112 & ~pi1113;
  assign new_n48879_ = pi1112 & pi1113;
  assign new_n48880_ = ~new_n48878_ & ~new_n48879_;
  assign new_n48881_ = ~pi1108 & ~pi1109;
  assign new_n48882_ = pi1108 & pi1109;
  assign new_n48883_ = ~new_n48881_ & ~new_n48882_;
  assign new_n48884_ = new_n48880_ & ~new_n48883_;
  assign new_n48885_ = ~new_n48880_ & new_n48883_;
  assign new_n48886_ = ~new_n48884_ & ~new_n48885_;
  assign new_n48887_ = new_n48877_ & new_n48886_;
  assign new_n48888_ = ~new_n48877_ & ~new_n48886_;
  assign new_n48889_ = ~new_n48887_ & ~new_n48888_;
  assign new_n48890_ = ~new_n48874_ & ~new_n48889_;
  assign new_n48891_ = pi0828 & new_n48783_;
  assign new_n48892_ = new_n48870_ & ~new_n48891_;
  assign new_n48893_ = ~new_n48873_ & new_n48889_;
  assign new_n48894_ = ~new_n48892_ & new_n48893_;
  assign po0985 = ~new_n48890_ & ~new_n48894_;
  assign new_n48896_ = new_n2797_ & new_n8870_;
  assign new_n48897_ = pi0951 & ~new_n48896_;
  assign po0986 = pi1092 & ~new_n48897_;
  assign new_n48899_ = pi0281 & ~new_n48712_;
  assign po0987 = ~new_n48713_ & ~new_n48899_;
  assign new_n48901_ = ~pi0832 & pi1091;
  assign new_n48902_ = pi1162 & new_n48901_;
  assign po0989 = new_n8874_ & new_n48902_;
  assign new_n48904_ = pi0833 & ~new_n2754_;
  assign po0990 = new_n17123_ | new_n48904_;
  assign po0991 = pi0946 & new_n2754_;
  assign new_n48907_ = pi0282 & ~new_n47029_;
  assign po0992 = ~new_n48736_ & ~new_n48907_;
  assign new_n48909_ = ~pi0955 & pi1049;
  assign new_n48910_ = pi0837 & pi0955;
  assign po0993 = new_n48909_ | new_n48910_;
  assign new_n48912_ = ~pi0955 & pi1047;
  assign new_n48913_ = pi0838 & pi0955;
  assign po0994 = new_n48912_ | new_n48913_;
  assign new_n48915_ = ~pi0955 & pi1074;
  assign new_n48916_ = pi0839 & pi0955;
  assign po0995 = new_n48915_ | new_n48916_;
  assign new_n48918_ = pi0840 & ~new_n2754_;
  assign new_n48919_ = pi1196 & new_n2754_;
  assign po0996 = new_n48918_ | new_n48919_;
  assign po0997 = ~pi0033 & new_n8979_;
  assign new_n48922_ = ~pi0955 & pi1035;
  assign new_n48923_ = pi0842 & pi0955;
  assign po0998 = new_n48922_ | new_n48923_;
  assign new_n48925_ = ~pi0955 & pi1079;
  assign new_n48926_ = pi0843 & pi0955;
  assign po0999 = new_n48925_ | new_n48926_;
  assign new_n48928_ = ~pi0955 & pi1078;
  assign new_n48929_ = pi0844 & pi0955;
  assign po1000 = new_n48928_ | new_n48929_;
  assign new_n48931_ = ~pi0955 & pi1043;
  assign new_n48932_ = pi0845 & pi0955;
  assign po1001 = new_n48931_ | new_n48932_;
  assign new_n48934_ = pi0846 & ~new_n42902_;
  assign new_n48935_ = pi1134 & new_n42902_;
  assign po1002 = new_n48934_ | new_n48935_;
  assign new_n48937_ = ~pi0955 & pi1055;
  assign new_n48938_ = pi0847 & pi0955;
  assign po1003 = new_n48937_ | new_n48938_;
  assign new_n48940_ = ~pi0955 & pi1039;
  assign new_n48941_ = pi0848 & pi0955;
  assign po1004 = new_n48940_ | new_n48941_;
  assign new_n48943_ = pi0849 & ~new_n2754_;
  assign new_n48944_ = pi1198 & new_n2754_;
  assign po1005 = new_n48943_ | new_n48944_;
  assign new_n48946_ = ~pi0955 & pi1048;
  assign new_n48947_ = pi0850 & pi0955;
  assign po1006 = new_n48946_ | new_n48947_;
  assign new_n48949_ = ~pi0955 & pi1045;
  assign new_n48950_ = pi0851 & pi0955;
  assign po1007 = new_n48949_ | new_n48950_;
  assign new_n48952_ = ~pi0955 & pi1062;
  assign new_n48953_ = pi0852 & pi0955;
  assign po1008 = new_n48952_ | new_n48953_;
  assign new_n48955_ = ~pi0955 & pi1080;
  assign new_n48956_ = pi0853 & pi0955;
  assign po1009 = new_n48955_ | new_n48956_;
  assign new_n48958_ = ~pi0955 & pi1051;
  assign new_n48959_ = pi0854 & pi0955;
  assign po1010 = new_n48958_ | new_n48959_;
  assign new_n48961_ = ~pi0955 & pi1065;
  assign new_n48962_ = pi0855 & pi0955;
  assign po1011 = new_n48961_ | new_n48962_;
  assign new_n48964_ = ~pi0955 & pi1067;
  assign new_n48965_ = pi0856 & pi0955;
  assign po1012 = new_n48964_ | new_n48965_;
  assign new_n48967_ = ~pi0955 & pi1058;
  assign new_n48968_ = pi0857 & pi0955;
  assign po1013 = new_n48967_ | new_n48968_;
  assign new_n48970_ = ~pi0955 & pi1087;
  assign new_n48971_ = pi0858 & pi0955;
  assign po1014 = new_n48970_ | new_n48971_;
  assign new_n48973_ = ~pi0955 & pi1070;
  assign new_n48974_ = pi0859 & pi0955;
  assign po1015 = new_n48973_ | new_n48974_;
  assign new_n48976_ = ~pi0955 & pi1076;
  assign new_n48977_ = pi0860 & pi0955;
  assign po1016 = new_n48976_ | new_n48977_;
  assign new_n48979_ = pi1093 & pi1141;
  assign new_n48980_ = pi0861 & ~pi1093;
  assign new_n48981_ = ~new_n48979_ & ~new_n48980_;
  assign new_n48982_ = ~pi0228 & ~new_n48981_;
  assign new_n48983_ = pi0123 & ~pi0861;
  assign new_n48984_ = ~pi0123 & ~pi1141;
  assign new_n48985_ = pi0228 & ~new_n48984_;
  assign new_n48986_ = ~new_n48983_ & new_n48985_;
  assign po1017 = new_n48982_ | new_n48986_;
  assign new_n48988_ = pi0862 & ~new_n42902_;
  assign new_n48989_ = pi1139 & new_n42902_;
  assign po1018 = new_n48988_ | new_n48989_;
  assign new_n48991_ = pi0863 & ~new_n2754_;
  assign new_n48992_ = pi1199 & new_n2754_;
  assign po1019 = new_n48991_ | new_n48992_;
  assign new_n48994_ = pi0864 & ~new_n2754_;
  assign new_n48995_ = pi1197 & new_n2754_;
  assign po1020 = new_n48994_ | new_n48995_;
  assign new_n48997_ = ~pi0955 & pi1040;
  assign new_n48998_ = pi0865 & pi0955;
  assign po1021 = new_n48997_ | new_n48998_;
  assign new_n49000_ = ~pi0955 & pi1053;
  assign new_n49001_ = pi0866 & pi0955;
  assign po1022 = new_n49000_ | new_n49001_;
  assign new_n49003_ = ~pi0955 & pi1057;
  assign new_n49004_ = pi0867 & pi0955;
  assign po1023 = new_n49003_ | new_n49004_;
  assign new_n49006_ = ~pi0955 & pi1063;
  assign new_n49007_ = pi0868 & pi0955;
  assign po1024 = new_n49006_ | new_n49007_;
  assign new_n49009_ = pi1093 & pi1140;
  assign new_n49010_ = pi0869 & ~pi1093;
  assign new_n49011_ = ~new_n49009_ & ~new_n49010_;
  assign new_n49012_ = ~pi0228 & ~new_n49011_;
  assign new_n49013_ = pi0123 & ~pi0869;
  assign new_n49014_ = ~pi0123 & ~pi1140;
  assign new_n49015_ = pi0228 & ~new_n49014_;
  assign new_n49016_ = ~new_n49013_ & new_n49015_;
  assign po1025 = new_n49012_ | new_n49016_;
  assign new_n49018_ = ~pi0955 & pi1069;
  assign new_n49019_ = pi0870 & pi0955;
  assign po1026 = new_n49018_ | new_n49019_;
  assign new_n49021_ = ~pi0955 & pi1072;
  assign new_n49022_ = pi0871 & pi0955;
  assign po1027 = new_n49021_ | new_n49022_;
  assign new_n49024_ = ~pi0955 & pi1084;
  assign new_n49025_ = pi0872 & pi0955;
  assign po1028 = new_n49024_ | new_n49025_;
  assign new_n49027_ = ~pi0955 & pi1044;
  assign new_n49028_ = pi0873 & pi0955;
  assign po1029 = new_n49027_ | new_n49028_;
  assign new_n49030_ = ~pi0955 & pi1036;
  assign new_n49031_ = pi0874 & pi0955;
  assign po1030 = new_n49030_ | new_n49031_;
  assign new_n49033_ = pi1093 & ~pi1136;
  assign new_n49034_ = ~pi0875 & ~pi1093;
  assign new_n49035_ = ~new_n49033_ & ~new_n49034_;
  assign new_n49036_ = ~pi0228 & ~new_n49035_;
  assign new_n49037_ = pi0123 & pi0875;
  assign new_n49038_ = ~pi0123 & pi1136;
  assign new_n49039_ = pi0228 & ~new_n49038_;
  assign new_n49040_ = ~new_n49037_ & new_n49039_;
  assign po1031 = ~new_n49036_ & ~new_n49040_;
  assign new_n49042_ = ~pi0955 & pi1037;
  assign new_n49043_ = pi0876 & pi0955;
  assign po1032 = new_n49042_ | new_n49043_;
  assign new_n49045_ = pi1093 & pi1138;
  assign new_n49046_ = pi0877 & ~pi1093;
  assign new_n49047_ = ~new_n49045_ & ~new_n49046_;
  assign new_n49048_ = ~pi0228 & ~new_n49047_;
  assign new_n49049_ = pi0123 & ~pi0877;
  assign new_n49050_ = ~pi0123 & ~pi1138;
  assign new_n49051_ = pi0228 & ~new_n49050_;
  assign new_n49052_ = ~new_n49049_ & new_n49051_;
  assign po1033 = new_n49048_ | new_n49052_;
  assign new_n49054_ = pi1093 & pi1137;
  assign new_n49055_ = pi0878 & ~pi1093;
  assign new_n49056_ = ~new_n49054_ & ~new_n49055_;
  assign new_n49057_ = ~pi0228 & ~new_n49056_;
  assign new_n49058_ = pi0123 & ~pi0878;
  assign new_n49059_ = ~pi0123 & ~pi1137;
  assign new_n49060_ = pi0228 & ~new_n49059_;
  assign new_n49061_ = ~new_n49058_ & new_n49060_;
  assign po1034 = new_n49057_ | new_n49061_;
  assign new_n49063_ = pi1093 & pi1135;
  assign new_n49064_ = pi0879 & ~pi1093;
  assign new_n49065_ = ~new_n49063_ & ~new_n49064_;
  assign new_n49066_ = ~pi0228 & ~new_n49065_;
  assign new_n49067_ = pi0123 & ~pi0879;
  assign new_n49068_ = ~pi0123 & ~pi1135;
  assign new_n49069_ = pi0228 & ~new_n49068_;
  assign new_n49070_ = ~new_n49067_ & new_n49069_;
  assign po1035 = new_n49066_ | new_n49070_;
  assign new_n49072_ = ~pi0955 & pi1081;
  assign new_n49073_ = pi0880 & pi0955;
  assign po1036 = new_n49072_ | new_n49073_;
  assign new_n49075_ = ~pi0955 & pi1059;
  assign new_n49076_ = pi0881 & pi0955;
  assign po1037 = new_n49075_ | new_n49076_;
  assign new_n49078_ = ~pi0883 & new_n48783_;
  assign po1039 = new_n48841_ | new_n49078_;
  assign new_n49080_ = pi1124 & ~new_n48783_;
  assign new_n49081_ = ~pi0884 & new_n48783_;
  assign po1040 = new_n49080_ | new_n49081_;
  assign new_n49083_ = pi1125 & ~new_n48783_;
  assign new_n49084_ = ~pi0885 & new_n48783_;
  assign po1041 = new_n49083_ | new_n49084_;
  assign new_n49086_ = pi1109 & ~new_n48783_;
  assign new_n49087_ = ~pi0886 & new_n48783_;
  assign po1042 = new_n49086_ | new_n49087_;
  assign new_n49089_ = ~pi0887 & new_n48783_;
  assign po1043 = new_n48840_ | new_n49089_;
  assign new_n49091_ = pi1120 & ~new_n48783_;
  assign new_n49092_ = ~pi0888 & new_n48783_;
  assign po1044 = new_n49091_ | new_n49092_;
  assign new_n49094_ = pi1103 & ~new_n48783_;
  assign new_n49095_ = ~pi0889 & new_n48783_;
  assign po1045 = new_n49094_ | new_n49095_;
  assign new_n49097_ = pi1126 & ~new_n48783_;
  assign new_n49098_ = ~pi0890 & new_n48783_;
  assign po1046 = new_n49097_ | new_n49098_;
  assign new_n49100_ = pi1116 & ~new_n48783_;
  assign new_n49101_ = ~pi0891 & new_n48783_;
  assign po1047 = new_n49100_ | new_n49101_;
  assign new_n49103_ = pi1101 & ~new_n48783_;
  assign new_n49104_ = ~pi0892 & new_n48783_;
  assign po1048 = new_n49103_ | new_n49104_;
  assign new_n49106_ = pi1119 & ~new_n48783_;
  assign new_n49107_ = ~pi0894 & new_n48783_;
  assign po1050 = new_n49106_ | new_n49107_;
  assign new_n49109_ = pi1113 & ~new_n48783_;
  assign new_n49110_ = ~pi0895 & new_n48783_;
  assign po1051 = new_n49109_ | new_n49110_;
  assign new_n49112_ = pi1118 & ~new_n48783_;
  assign new_n49113_ = ~pi0896 & new_n48783_;
  assign po1052 = new_n49112_ | new_n49113_;
  assign new_n49115_ = pi1129 & ~new_n48783_;
  assign new_n49116_ = ~pi0898 & new_n48783_;
  assign po1054 = new_n49115_ | new_n49116_;
  assign new_n49118_ = ~pi0899 & new_n48783_;
  assign po1055 = new_n48868_ | new_n49118_;
  assign new_n49120_ = pi1110 & ~new_n48783_;
  assign new_n49121_ = ~pi0900 & new_n48783_;
  assign po1056 = new_n49120_ | new_n49121_;
  assign new_n49123_ = pi1111 & ~new_n48783_;
  assign new_n49124_ = ~pi0902 & new_n48783_;
  assign po1058 = new_n49123_ | new_n49124_;
  assign new_n49126_ = pi1121 & ~new_n48783_;
  assign new_n49127_ = ~pi0903 & new_n48783_;
  assign po1059 = new_n49126_ | new_n49127_;
  assign new_n49129_ = ~pi0904 & new_n48783_;
  assign po1060 = new_n48785_ | new_n49129_;
  assign new_n49131_ = ~pi0905 & new_n48783_;
  assign po1061 = new_n48784_ | new_n49131_;
  assign new_n49133_ = pi1128 & ~new_n48783_;
  assign new_n49134_ = ~pi0906 & new_n48783_;
  assign po1062 = new_n49133_ | new_n49134_;
  assign new_n49136_ = ~pi0604 & ~pi0979;
  assign new_n49137_ = pi0615 & pi0979;
  assign new_n49138_ = ~new_n49136_ & ~new_n49137_;
  assign new_n49139_ = pi0782 & ~new_n49138_;
  assign new_n49140_ = ~pi0782 & ~pi0907;
  assign new_n49141_ = ~pi0598 & pi0979;
  assign new_n49142_ = ~pi0624 & ~pi0979;
  assign new_n49143_ = pi0782 & ~new_n49142_;
  assign new_n49144_ = ~new_n49141_ & new_n49143_;
  assign new_n49145_ = ~new_n49140_ & ~new_n49144_;
  assign po1063 = ~new_n49139_ & new_n49145_;
  assign new_n49147_ = ~pi0908 & new_n48783_;
  assign po1064 = new_n48813_ | new_n49147_;
  assign new_n49149_ = pi1105 & ~new_n48783_;
  assign new_n49150_ = ~pi0909 & new_n48783_;
  assign po1065 = new_n49149_ | new_n49150_;
  assign new_n49152_ = pi1117 & ~new_n48783_;
  assign new_n49153_ = ~pi0910 & new_n48783_;
  assign po1066 = new_n49152_ | new_n49153_;
  assign new_n49155_ = pi1130 & ~new_n48783_;
  assign new_n49156_ = ~pi0911 & new_n48783_;
  assign po1067 = new_n49155_ | new_n49156_;
  assign new_n49158_ = ~pi0912 & new_n48783_;
  assign po1068 = new_n48869_ | new_n49158_;
  assign new_n49160_ = pi1106 & ~new_n48783_;
  assign new_n49161_ = ~pi0913 & new_n48783_;
  assign po1069 = new_n49160_ | new_n49161_;
  assign new_n49163_ = pi0280 & ~new_n47026_;
  assign po1070 = ~new_n47027_ & ~new_n49163_;
  assign new_n49165_ = pi1108 & ~new_n48783_;
  assign new_n49166_ = ~pi0915 & new_n48783_;
  assign po1071 = new_n49165_ | new_n49166_;
  assign new_n49168_ = ~pi0916 & new_n48783_;
  assign po1072 = new_n48812_ | new_n49168_;
  assign new_n49170_ = pi1112 & ~new_n48783_;
  assign new_n49171_ = ~pi0917 & new_n48783_;
  assign po1073 = new_n49170_ | new_n49171_;
  assign new_n49173_ = pi1104 & ~new_n48783_;
  assign new_n49174_ = ~pi0918 & new_n48783_;
  assign po1074 = new_n49173_ | new_n49174_;
  assign new_n49176_ = pi1102 & ~new_n48783_;
  assign new_n49177_ = ~pi0919 & new_n48783_;
  assign po1075 = new_n49176_ | new_n49177_;
  assign new_n49179_ = pi1093 & pi1139;
  assign new_n49180_ = pi0920 & ~pi1093;
  assign po1076 = new_n49179_ | new_n49180_;
  assign new_n49182_ = pi0921 & ~pi1093;
  assign po1077 = new_n49009_ | new_n49182_;
  assign new_n49184_ = ~pi0922 & ~pi1093;
  assign new_n49185_ = pi1093 & ~pi1152;
  assign po1078 = ~new_n49184_ & ~new_n49185_;
  assign new_n49187_ = ~pi0923 & ~pi1093;
  assign new_n49188_ = pi1093 & ~pi1154;
  assign po1079 = ~new_n49187_ & ~new_n49188_;
  assign new_n49190_ = ~pi0300 & pi0301;
  assign new_n49191_ = pi0311 & ~pi0312;
  assign po1080 = new_n49190_ & new_n49191_;
  assign new_n49193_ = ~pi0925 & ~pi1093;
  assign new_n49194_ = pi1093 & ~pi1155;
  assign po1081 = ~new_n49193_ & ~new_n49194_;
  assign new_n49196_ = ~pi0926 & ~pi1093;
  assign new_n49197_ = pi1093 & ~pi1157;
  assign po1082 = ~new_n49196_ & ~new_n49197_;
  assign new_n49199_ = ~pi0927 & ~pi1093;
  assign new_n49200_ = pi1093 & ~pi1145;
  assign po1083 = ~new_n49199_ & ~new_n49200_;
  assign new_n49202_ = ~pi0928 & ~pi1093;
  assign po1084 = ~new_n49033_ & ~new_n49202_;
  assign new_n49204_ = ~pi0929 & ~pi1093;
  assign new_n49205_ = pi1093 & ~pi1144;
  assign po1085 = ~new_n49204_ & ~new_n49205_;
  assign new_n49207_ = ~pi0930 & ~pi1093;
  assign new_n49208_ = pi1093 & ~pi1134;
  assign po1086 = ~new_n49207_ & ~new_n49208_;
  assign new_n49210_ = ~pi0931 & ~pi1093;
  assign new_n49211_ = pi1093 & ~pi1150;
  assign po1087 = ~new_n49210_ & ~new_n49211_;
  assign new_n49213_ = pi0932 & ~pi1093;
  assign po1088 = new_n42891_ | new_n49213_;
  assign new_n49215_ = pi0933 & ~pi1093;
  assign po1089 = new_n49054_ | new_n49215_;
  assign new_n49217_ = ~pi0934 & ~pi1093;
  assign new_n49218_ = pi1093 & ~pi1147;
  assign po1090 = ~new_n49217_ & ~new_n49218_;
  assign new_n49220_ = pi0935 & ~pi1093;
  assign po1091 = new_n48979_ | new_n49220_;
  assign new_n49222_ = ~pi0936 & ~pi1093;
  assign new_n49223_ = pi1093 & ~pi1149;
  assign po1092 = ~new_n49222_ & ~new_n49223_;
  assign new_n49225_ = ~pi0937 & ~pi1093;
  assign new_n49226_ = pi1093 & ~pi1148;
  assign po1093 = ~new_n49225_ & ~new_n49226_;
  assign new_n49228_ = pi0938 & ~pi1093;
  assign po1094 = new_n49063_ | new_n49228_;
  assign new_n49230_ = ~pi0939 & ~pi1093;
  assign new_n49231_ = pi1093 & ~pi1146;
  assign po1095 = ~new_n49230_ & ~new_n49231_;
  assign new_n49233_ = pi0940 & ~pi1093;
  assign po1096 = new_n49045_ | new_n49233_;
  assign new_n49235_ = ~pi0941 & ~pi1093;
  assign new_n49236_ = pi1093 & ~pi1153;
  assign po1097 = ~new_n49235_ & ~new_n49236_;
  assign new_n49238_ = ~pi0942 & ~pi1093;
  assign new_n49239_ = pi1093 & ~pi1156;
  assign po1098 = ~new_n49238_ & ~new_n49239_;
  assign new_n49241_ = ~pi0943 & ~pi1093;
  assign new_n49242_ = pi1093 & ~pi1151;
  assign po1099 = ~new_n49241_ & ~new_n49242_;
  assign new_n49244_ = pi1093 & pi1143;
  assign new_n49245_ = pi0944 & ~pi1093;
  assign po1100 = new_n49244_ | new_n49245_;
  assign po1102 = pi0230 & new_n2754_;
  assign new_n49248_ = ~pi0782 & pi0947;
  assign po1103 = new_n49144_ | new_n49248_;
  assign new_n49250_ = ~pi0266 & ~pi0992;
  assign po1104 = ~new_n47026_ & ~new_n49250_;
  assign new_n49252_ = ~pi0313 & ~pi0954;
  assign new_n49253_ = pi0949 & pi0954;
  assign po1105 = new_n49252_ | new_n49253_;
  assign po1107 = ~new_n7572_ & new_n14258_;
  assign new_n49256_ = pi0957 & pi1092;
  assign po1112 = pi0031 | new_n49256_;
  assign po1115 = ~pi0782 & pi0960;
  assign po1116 = ~pi0230 & pi0961;
  assign po1118 = ~pi0782 & pi0963;
  assign po1122 = ~pi0230 & pi0967;
  assign po1124 = ~pi0230 & pi0969;
  assign po1125 = ~pi0782 & pi0970;
  assign po1126 = ~pi0230 & pi0971;
  assign po1127 = ~pi0782 & pi0972;
  assign po1128 = ~pi0230 & pi0974;
  assign po1129 = ~pi0782 & pi0975;
  assign po1131 = ~pi0230 & pi0977;
  assign po1132 = ~pi0782 & pi0978;
  assign po1133 = pi0598 | ~pi0615;
  assign po1135 = pi0824 & pi1092;
  assign po1137 = pi0604 | pi0624;
  assign po0166 = 1'b1;
  assign po0170 = ~pi1090;
  assign po1110 = ~pi0954;
  assign po1130 = ~pi0278;
  assign po1146 = ~pi0915;
  assign po1147 = ~pi0825;
  assign po1148 = ~pi0826;
  assign po1149 = ~pi0913;
  assign po1150 = ~pi0894;
  assign po1151 = ~pi0905;
  assign po1153 = ~pi0890;
  assign po1155 = ~pi0906;
  assign po1156 = ~pi0896;
  assign po1157 = ~pi0909;
  assign po1158 = ~pi0911;
  assign po1159 = ~pi0908;
  assign po1160 = ~pi0891;
  assign po1161 = ~pi0902;
  assign po1162 = ~pi0903;
  assign po1163 = ~pi0883;
  assign po1164 = ~pi0888;
  assign po1165 = ~pi0919;
  assign po1166 = ~pi0886;
  assign po1167 = ~pi0912;
  assign po1168 = ~pi0895;
  assign po1169 = ~pi0916;
  assign po1170 = ~pi0889;
  assign po1171 = ~pi0900;
  assign po1172 = ~pi0885;
  assign po1173 = ~pi0904;
  assign po1174 = ~pi0899;
  assign po1175 = ~pi0918;
  assign po1176 = ~pi0898;
  assign po1177 = ~pi0917;
  assign po1178 = ~pi0827;
  assign po1179 = ~pi0887;
  assign po1180 = ~pi0884;
  assign po1181 = ~pi0910;
  assign po1182 = ~pi0828;
  assign po1183 = ~pi0892;
  assign po0000 = pi0668;
  assign po0001 = pi0672;
  assign po0002 = pi0664;
  assign po0003 = pi0667;
  assign po0004 = pi0676;
  assign po0005 = pi0673;
  assign po0006 = pi0675;
  assign po0007 = pi0666;
  assign po0008 = pi0679;
  assign po0009 = pi0674;
  assign po0010 = pi0663;
  assign po0011 = pi0670;
  assign po0012 = pi0677;
  assign po0013 = pi0682;
  assign po0014 = pi0671;
  assign po0015 = pi0678;
  assign po0016 = pi0718;
  assign po0017 = pi0707;
  assign po0018 = pi0708;
  assign po0019 = pi0713;
  assign po0020 = pi0711;
  assign po0021 = pi0716;
  assign po0022 = pi0733;
  assign po0023 = pi0712;
  assign po0024 = pi0689;
  assign po0025 = pi0717;
  assign po0026 = pi0692;
  assign po0027 = pi0719;
  assign po0028 = pi0722;
  assign po0029 = pi0714;
  assign po0030 = pi0720;
  assign po0031 = pi0685;
  assign po0032 = pi0837;
  assign po0033 = pi0850;
  assign po0034 = pi0872;
  assign po0035 = pi0871;
  assign po0036 = pi0881;
  assign po0037 = pi0866;
  assign po0038 = pi0876;
  assign po0039 = pi0873;
  assign po0040 = pi0874;
  assign po0041 = pi0859;
  assign po0042 = pi0855;
  assign po0043 = pi0852;
  assign po0044 = pi0870;
  assign po0045 = pi0848;
  assign po0046 = pi0865;
  assign po0047 = pi0856;
  assign po0048 = pi0853;
  assign po0049 = pi0847;
  assign po0050 = pi0857;
  assign po0051 = pi0854;
  assign po0052 = pi0858;
  assign po0053 = pi0845;
  assign po0054 = pi0838;
  assign po0055 = pi0842;
  assign po0056 = pi0843;
  assign po0057 = pi0839;
  assign po0058 = pi0844;
  assign po0059 = pi0868;
  assign po0060 = pi0851;
  assign po0061 = pi0867;
  assign po0062 = pi0880;
  assign po0063 = pi0860;
  assign po0064 = pi1030;
  assign po0065 = pi1034;
  assign po0066 = pi1015;
  assign po0067 = pi1020;
  assign po0068 = pi1025;
  assign po0069 = pi1005;
  assign po0070 = pi0996;
  assign po0071 = pi1012;
  assign po0072 = pi0993;
  assign po0073 = pi1016;
  assign po0074 = pi1021;
  assign po0075 = pi1010;
  assign po0076 = pi1027;
  assign po0077 = pi1018;
  assign po0078 = pi1017;
  assign po0079 = pi1024;
  assign po0080 = pi1009;
  assign po0081 = pi1032;
  assign po0082 = pi1003;
  assign po0083 = pi0997;
  assign po0084 = pi1013;
  assign po0085 = pi1011;
  assign po0086 = pi1008;
  assign po0087 = pi1019;
  assign po0088 = pi1031;
  assign po0089 = pi1022;
  assign po0090 = pi1000;
  assign po0091 = pi1023;
  assign po0092 = pi1002;
  assign po0093 = pi1026;
  assign po0094 = pi1006;
  assign po0095 = pi0998;
  assign po0096 = pi0031;
  assign po0097 = pi0080;
  assign po0098 = pi0893;
  assign po0099 = pi0467;
  assign po0100 = pi0078;
  assign po0101 = pi0112;
  assign po0102 = pi0013;
  assign po0103 = pi0025;
  assign po0104 = pi0226;
  assign po0105 = pi0127;
  assign po0106 = pi0822;
  assign po0107 = pi0808;
  assign po0108 = pi0227;
  assign po0109 = pi0477;
  assign po0110 = pi0834;
  assign po0111 = pi0229;
  assign po0112 = pi0012;
  assign po0113 = pi0011;
  assign po0114 = pi0010;
  assign po0115 = pi0009;
  assign po0116 = pi0008;
  assign po0117 = pi0007;
  assign po0118 = pi0006;
  assign po0119 = pi0005;
  assign po0120 = pi0004;
  assign po0121 = pi0003;
  assign po0122 = pi0000;
  assign po0123 = pi0002;
  assign po0124 = pi0001;
  assign po0125 = pi0310;
  assign po0126 = pi0302;
  assign po0127 = pi0475;
  assign po0128 = pi0474;
  assign po0129 = pi0466;
  assign po0130 = pi0473;
  assign po0131 = pi0471;
  assign po0132 = pi0472;
  assign po0133 = pi0470;
  assign po0134 = pi0469;
  assign po0135 = pi0465;
  assign po0136 = pi1028;
  assign po0137 = pi1033;
  assign po0138 = pi0995;
  assign po0139 = pi0994;
  assign po0140 = pi0028;
  assign po0141 = pi0027;
  assign po0142 = pi0026;
  assign po0143 = pi0029;
  assign po0144 = pi0015;
  assign po0145 = pi0014;
  assign po0146 = pi0021;
  assign po0147 = pi0020;
  assign po0148 = pi0019;
  assign po0149 = pi0018;
  assign po0150 = pi0017;
  assign po0151 = pi0016;
  assign po0152 = pi1096;
  assign po0168 = pi0228;
  assign po0169 = pi0022;
  assign po0179 = pi1089;
  assign po0180 = pi0023;
  assign po0181 = po0167;
  assign po0188 = pi0037;
  assign po0263 = pi0117;
  assign po0285 = pi0131;
  assign po0386 = pi0232;
  assign po0388 = pi0236;
  assign po0636 = pi0583;
  assign po1053 = pi0067;
  assign po1108 = pi1134;
  assign po1109 = pi0964;
  assign po1111 = pi0965;
  assign po1113 = pi0991;
  assign po1114 = pi0985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi0299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi0771;
  assign po1141 = pi0765;
  assign po1142 = pi0605;
  assign po1143 = pi0601;
  assign po1144 = pi0278;
  assign po1145 = pi0279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi0863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi0230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi0849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi0840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi0864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule


