module top(a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_, a_31_, a_32_, a_33_, a_34_, a_35_, a_36_, a_37_, a_38_, a_39_, a_40_, a_41_, a_42_, a_43_, a_44_, a_45_, a_46_, a_47_, a_48_, a_49_, a_50_, a_51_, a_52_, a_53_, a_54_, a_55_, a_56_, a_57_, a_58_, a_59_, a_60_, a_61_, a_62_, a_63_, a_64_, a_65_, a_66_, a_67_, a_68_, a_69_, a_70_, a_71_, a_72_, a_73_, a_74_, a_75_, a_76_, a_77_, a_78_, a_79_, a_80_, a_81_, a_82_, a_83_, a_84_, a_85_, a_86_, a_87_, a_88_, a_89_, a_90_, a_91_, a_92_, a_93_, a_94_, a_95_, a_96_, a_97_, a_98_, a_99_, a_100_, a_101_, a_102_, a_103_, a_104_, a_105_, a_106_, a_107_, a_108_, a_109_, a_110_, a_111_, a_112_, a_113_, a_114_, a_115_, a_116_, a_117_, a_118_, a_119_, a_120_, a_121_, a_122_, a_123_, a_124_, a_125_, a_126_, a_127_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, b_32_, b_33_, b_34_, b_35_, b_36_, b_37_, b_38_, b_39_, b_40_, b_41_, b_42_, b_43_, b_44_, b_45_, b_46_, b_47_, b_48_, b_49_, b_50_, b_51_, b_52_, b_53_, b_54_, b_55_, b_56_, b_57_, b_58_, b_59_, b_60_, b_61_, b_62_, b_63_, b_64_, b_65_, b_66_, b_67_, b_68_, b_69_, b_70_, b_71_, b_72_, b_73_, b_74_, b_75_, b_76_, b_77_, b_78_, b_79_, b_80_, b_81_, b_82_, b_83_, b_84_, b_85_, b_86_, b_87_, b_88_, b_89_, b_90_, b_91_, b_92_, b_93_, b_94_, b_95_, b_96_, b_97_, b_98_, b_99_, b_100_, b_101_, b_102_, b_103_, b_104_, b_105_, b_106_, b_107_, b_108_, b_109_, b_110_, b_111_, b_112_, b_113_, b_114_, b_115_, b_116_, b_117_, b_118_, b_119_, b_120_, b_121_, b_122_, b_123_, b_124_, b_125_, b_126_, b_127_, f_0_, f_1_, f_2_, f_3_, f_4_, f_5_, f_6_, f_7_, f_8_, f_9_, f_10_, f_11_, f_12_, f_13_, f_14_, f_15_, f_16_, f_17_, f_18_, f_19_, f_20_, f_21_, f_22_, f_23_, f_24_, f_25_, f_26_, f_27_, f_28_, f_29_, f_30_, f_31_, f_32_, f_33_, f_34_, f_35_, f_36_, f_37_, f_38_, f_39_, f_40_, f_41_, f_42_, f_43_, f_44_, f_45_, f_46_, f_47_, f_48_, f_49_, f_50_, f_51_, f_52_, f_53_, f_54_, f_55_, f_56_, f_57_, f_58_, f_59_, f_60_, f_61_, f_62_, f_63_, f_64_, f_65_, f_66_, f_67_, f_68_, f_69_, f_70_, f_71_, f_72_, f_73_, f_74_, f_75_, f_76_, f_77_, f_78_, f_79_, f_80_, f_81_, f_82_, f_83_, f_84_, f_85_, f_86_, f_87_, f_88_, f_89_, f_90_, f_91_, f_92_, f_93_, f_94_, f_95_, f_96_, f_97_, f_98_, f_99_, f_100_, f_101_, f_102_, f_103_, f_104_, f_105_, f_106_, f_107_, f_108_, f_109_, f_110_, f_111_, f_112_, f_113_, f_114_, f_115_, f_116_, f_117_, f_118_, f_119_, f_120_, f_121_, f_122_, f_123_, f_124_, f_125_, f_126_, f_127_, cOut);
  wire n392;
  wire n391;
  wire n396;
  wire n400;
  wire n399;
  wire n404;
  wire n408;
  wire n407;
  wire n412;
  wire n416;
  wire n415;
  wire n420;
  wire n424;
  wire n423;
  wire n428;
  wire n432;
  wire n431;
  wire n436;
  wire n440;
  wire n439;
  wire n444;
  wire n448;
  wire n447;
  wire n452;
  wire n456;
  wire n455;
  wire n460;
  wire n464;
  wire n463;
  wire n468;
  wire n472;
  wire n471;
  wire n476;
  wire n480;
  wire n479;
  wire n484;
  wire n488;
  wire n487;
  wire n492;
  wire n496;
  wire n495;
  wire n500;
  wire n504;
  wire n503;
  wire n508;
  wire n512;
  wire n511;
  wire n516;
  wire n520;
  wire n519;
  wire n524;
  wire n528;
  wire n527;
  wire n532;
  wire n536;
  wire n535;
  wire n540;
  wire n544;
  wire n543;
  wire n548;
  wire n552;
  wire n551;
  wire n556;
  wire n560;
  wire n559;
  wire n564;
  wire n568;
  wire n567;
  wire n572;
  wire n576;
  wire n575;
  wire n580;
  wire n584;
  wire n583;
  wire n588;
  wire n592;
  wire n591;
  wire n596;
  wire n600;
  wire n599;
  wire n604;
  wire n608;
  wire n607;
  wire n612;
  wire n616;
  wire n615;
  wire n620;
  wire n624;
  wire n623;
  wire n628;
  wire n632;
  wire n631;
  wire n636;
  wire n640;
  wire n639;
  wire n644;
  wire n648;
  wire n647;
  wire n652;
  wire n656;
  wire n655;
  wire n660;
  wire n664;
  wire n663;
  wire n668;
  wire n672;
  wire n671;
  wire n676;
  wire n680;
  wire n679;
  wire n684;
  wire n688;
  wire n687;
  wire n692;
  wire n696;
  wire n695;
  wire n700;
  wire n704;
  wire n703;
  wire n708;
  wire n712;
  wire n711;
  wire n716;
  wire n720;
  wire n719;
  wire n724;
  wire n728;
  wire n727;
  wire n732;
  wire n736;
  wire n735;
  wire n740;
  wire n744;
  wire n743;
  wire n748;
  wire n752;
  wire n751;
  wire n756;
  wire n760;
  wire n759;
  wire n764;
  wire n768;
  wire n767;
  wire n772;
  wire n776;
  wire n775;
  wire n780;
  wire n784;
  wire n783;
  wire n788;
  wire n792;
  wire n791;
  wire n796;
  wire n800;
  wire n799;
  wire n804;
  wire n808;
  wire n807;
  wire n812;
  wire n816;
  wire n815;
  wire n820;
  wire n824;
  wire n823;
  wire n828;
  wire n832;
  wire n831;
  wire n836;
  wire n840;
  wire n839;
  wire n844;
  wire n848;
  wire n847;
  wire n852;
  wire n856;
  wire n855;
  wire n860;
  wire n864;
  wire n863;
  wire n868;
  wire n872;
  wire n871;
  wire n876;
  wire n880;
  wire n879;
  wire n884;
  wire n888;
  wire n887;
  wire n892;
  wire n896;
  wire n895;
  wire n900;
  wire n904;
  wire n903;
  wire n908;
  wire n912;
  wire n911;
  wire n916;
  wire n920;
  wire n919;
  wire n924;
  wire n928;
  wire n927;
  wire n932;
  wire n936;
  wire n935;
  wire n940;
  wire n944;
  wire n943;
  wire n948;
  wire n952;
  wire n951;
  wire n956;
  wire n960;
  wire n959;
  wire n964;
  wire n968;
  wire n967;
  wire n972;
  wire n976;
  wire n975;
  wire n980;
  wire n984;
  wire n983;
  wire n988;
  wire n992;
  wire n1000;
  wire n991;
  wire n996;
  wire n1004;
  wire n1008;
  wire n999;
  wire n1007;
  wire n1012;
  wire n1016;
  wire n1015;
  wire n1020;
  wire n1024;
  wire n1023;
  wire n1028;
  wire n1032;
  wire n1031;
  wire n1036;
  wire n1040;
  wire n1039;
  wire n1044;
  wire n1048;
  wire n1047;
  wire n1052;
  wire n1056;
  wire n1055;
  wire n1060;
  wire n1064;
  wire n1063;
  wire n1068;
  wire n1072;
  wire n1071;
  wire n1076;
  wire n1080;
  wire n1079;
  wire n1084;
  wire n1088;
  wire n1087;
  wire n1092;
  wire n1096;
  wire n1095;
  wire n1100;
  wire n1104;
  wire n1103;
  wire n1108;
  wire n1112;
  wire n1111;
  wire n1116;
  wire n1120;
  wire n1119;
  wire n1124;
  wire n1128;
  wire n1127;
  wire n1132;
  wire n1136;
  wire n1135;
  wire n1140;
  wire n1144;
  wire n1143;
  wire n1148;
  wire n1152;
  wire n1151;
  wire n1156;
  wire n1160;
  wire n1159;
  wire n1164;
  wire n1168;
  wire n1167;
  wire n1172;
  wire n1176;
  wire n1175;
  wire n1180;
  wire n1184;
  wire n1183;
  wire n1188;
  wire n1192;
  wire n1191;
  wire n1196;
  wire n1200;
  wire n1199;
  wire n1204;
  wire n1208;
  wire n1207;
  wire n1212;
  wire n1216;
  wire n1215;
  wire n1220;
  wire n1224;
  wire n1223;
  wire n1228;
  wire n1232;
  wire n1231;
  wire n1236;
  wire n1240;
  wire n1239;
  wire n1244;
  wire n1248;
  wire n1247;
  wire n1252;
  wire n1256;
  wire n1255;
  wire n1260;
  wire n1264;
  wire n1263;
  wire n1268;
  wire n1272;
  wire n1271;
  wire n1276;
  wire n1280;
  wire n1279;
  wire n1284;
  wire n1288;
  wire n1287;
  wire n1292;
  wire n1296;
  wire n1295;
  wire n1300;
  wire n1304;
  wire n1303;
  wire n1308;
  wire n1312;
  wire n1311;
  wire n1316;
  wire n1320;
  wire n1319;
  wire n1324;
  wire n1328;
  wire n1327;
  wire n1332;
  wire n1336;
  wire n1335;
  wire n1340;
  wire n1344;
  wire n1343;
  wire n1348;
  wire n1352;
  wire n1351;
  wire n1356;
  wire n1360;
  wire n1359;
  wire n1364;
  wire n1368;
  wire n1367;
  wire n1372;
  wire n1376;
  wire n1375;
  wire n1380;
  wire n1384;
  wire n1383;
  wire n1388;
  wire n1392;
  wire n1391;
  wire n1396;
  wire n1400;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n390;
  wire n1389;
  wire n1390;
  wire n1381;
  wire n1382;
  wire n1373;
  wire n1374;
  wire n1365;
  wire n1366;
  wire n1357;
  wire n1358;
  wire n1349;
  wire n1350;
  wire n1341;
  wire n1342;
  wire n1333;
  wire n1334;
  wire n1325;
  wire n1326;
  wire n1317;
  wire n1318;
  wire n1309;
  wire n1310;
  wire n1301;
  wire n1302;
  wire n1293;
  wire n1294;
  wire n1285;
  wire n1286;
  wire n1277;
  wire n1278;
  wire n1269;
  wire n1270;
  wire n1261;
  wire n1262;
  wire n1253;
  wire n1254;
  wire n1245;
  wire n1246;
  wire n1237;
  wire n1238;
  wire n1229;
  wire n1230;
  wire n1221;
  wire n1222;
  wire n1213;
  wire n1214;
  wire n1205;
  wire n1206;
  wire n1197;
  wire n1198;
  wire n1189;
  wire n1190;
  wire n1181;
  wire n1182;
  wire n1173;
  wire n1174;
  wire n1165;
  wire n1166;
  wire n1157;
  wire n1158;
  wire n1149;
  wire n1150;
  wire n1141;
  wire n1142;
  wire n1133;
  wire n1134;
  wire n1125;
  wire n1126;
  wire n1117;
  wire n1118;
  wire n1109;
  wire n1110;
  wire n1101;
  wire n1102;
  wire n1093;
  wire n1094;
  wire n1085;
  wire n1086;
  wire n1077;
  wire n1078;
  wire n1069;
  wire n1070;
  wire n1061;
  wire n1062;
  wire n1053;
  wire n1054;
  wire n1045;
  wire n1046;
  wire n1037;
  wire n1038;
  wire n1029;
  wire n1030;
  wire n1021;
  wire n1022;
  wire n1013;
  wire n1014;
  wire n1005;
  wire n1006;
  wire n997;
  wire n998;
  wire n989;
  wire n990;
  wire n981;
  wire n982;
  wire n973;
  wire n974;
  wire n965;
  wire n966;
  wire n957;
  wire n958;
  wire n949;
  wire n950;
  wire n941;
  wire n942;
  wire n933;
  wire n934;
  wire n925;
  wire n926;
  wire n917;
  wire n918;
  wire n909;
  wire n910;
  wire n901;
  wire n902;
  wire n893;
  wire n894;
  wire n885;
  wire n886;
  wire n877;
  wire n878;
  wire n869;
  wire n870;
  wire n861;
  wire n862;
  wire n853;
  wire n854;
  wire n845;
  wire n846;
  wire n837;
  wire n838;
  wire n829;
  wire n830;
  wire n821;
  wire n822;
  wire n813;
  wire n814;
  wire n805;
  wire n806;
  wire n797;
  wire n798;
  wire n789;
  wire n790;
  wire n781;
  wire n782;
  wire n773;
  wire n774;
  wire n765;
  wire n766;
  wire n757;
  wire n758;
  wire n749;
  wire n750;
  wire n741;
  wire n742;
  wire n733;
  wire n734;
  wire n725;
  wire n726;
  wire n717;
  wire n718;
  wire n709;
  wire n710;
  wire n701;
  wire n702;
  wire n693;
  wire n694;
  wire n685;
  wire n686;
  wire n677;
  wire n678;
  wire n669;
  wire n670;
  wire n661;
  wire n662;
  wire n653;
  wire n654;
  wire n645;
  wire n646;
  wire n637;
  wire n638;
  wire n629;
  wire n630;
  wire n621;
  wire n622;
  wire n613;
  wire n614;
  wire n605;
  wire n606;
  wire n597;
  wire n598;
  wire n589;
  wire n590;
  wire n581;
  wire n582;
  wire n573;
  wire n574;
  wire n565;
  wire n566;
  wire n557;
  wire n558;
  wire n549;
  wire n550;
  wire n541;
  wire n542;
  wire n533;
  wire n534;
  wire n525;
  wire n526;
  wire n517;
  wire n518;
  wire n509;
  wire n510;
  wire n501;
  wire n502;
  wire n493;
  wire n494;
  wire n485;
  wire n486;
  wire n477;
  wire n478;
  wire n469;
  wire n470;
  wire n461;
  wire n462;
  wire n453;
  wire n454;
  wire n445;
  wire n446;
  wire n437;
  wire n438;
  wire n429;
  wire n430;
  wire n421;
  wire n422;
  wire n413;
  wire n414;
  wire n405;
  wire n406;
  wire n397;
  wire n398;
  wire n389;
  input a_0_;
  input a_1_;
  input a_2_;
  input a_3_;
  input a_4_;
  input a_5_;
  input a_6_;
  input a_7_;
  input a_8_;
  input a_9_;
  input a_10_;
  input a_11_;
  input a_12_;
  input a_13_;
  input a_14_;
  input a_15_;
  input a_16_;
  input a_17_;
  input a_18_;
  input a_19_;
  input a_20_;
  input a_21_;
  input a_22_;
  input a_23_;
  input a_24_;
  input a_25_;
  input a_26_;
  input a_27_;
  input a_28_;
  input a_29_;
  input a_30_;
  input a_31_;
  input a_32_;
  input a_33_;
  input a_34_;
  input a_35_;
  input a_36_;
  input a_37_;
  input a_38_;
  input a_39_;
  input a_40_;
  input a_41_;
  input a_42_;
  input a_43_;
  input a_44_;
  input a_45_;
  input a_46_;
  input a_47_;
  input a_48_;
  input a_49_;
  input a_50_;
  input a_51_;
  input a_52_;
  input a_53_;
  input a_54_;
  input a_55_;
  input a_56_;
  input a_57_;
  input a_58_;
  input a_59_;
  input a_60_;
  input a_61_;
  input a_62_;
  input a_63_;
  input a_64_;
  input a_65_;
  input a_66_;
  input a_67_;
  input a_68_;
  input a_69_;
  input a_70_;
  input a_71_;
  input a_72_;
  input a_73_;
  input a_74_;
  input a_75_;
  input a_76_;
  input a_77_;
  input a_78_;
  input a_79_;
  input a_80_;
  input a_81_;
  input a_82_;
  input a_83_;
  input a_84_;
  input a_85_;
  input a_86_;
  input a_87_;
  input a_88_;
  input a_89_;
  input a_90_;
  input a_91_;
  input a_92_;
  input a_93_;
  input a_94_;
  input a_95_;
  input a_96_;
  input a_97_;
  input a_98_;
  input a_99_;
  input a_100_;
  input a_101_;
  input a_102_;
  input a_103_;
  input a_104_;
  input a_105_;
  input a_106_;
  input a_107_;
  input a_108_;
  input a_109_;
  input a_110_;
  input a_111_;
  input a_112_;
  input a_113_;
  input a_114_;
  input a_115_;
  input a_116_;
  input a_117_;
  input a_118_;
  input a_119_;
  input a_120_;
  input a_121_;
  input a_122_;
  input a_123_;
  input a_124_;
  input a_125_;
  input a_126_;
  input a_127_;
  input b_0_;
  input b_1_;
  input b_2_;
  input b_3_;
  input b_4_;
  input b_5_;
  input b_6_;
  input b_7_;
  input b_8_;
  input b_9_;
  input b_10_;
  input b_11_;
  input b_12_;
  input b_13_;
  input b_14_;
  input b_15_;
  input b_16_;
  input b_17_;
  input b_18_;
  input b_19_;
  input b_20_;
  input b_21_;
  input b_22_;
  input b_23_;
  input b_24_;
  input b_25_;
  input b_26_;
  input b_27_;
  input b_28_;
  input b_29_;
  input b_30_;
  input b_31_;
  input b_32_;
  input b_33_;
  input b_34_;
  input b_35_;
  input b_36_;
  input b_37_;
  input b_38_;
  input b_39_;
  input b_40_;
  input b_41_;
  input b_42_;
  input b_43_;
  input b_44_;
  input b_45_;
  input b_46_;
  input b_47_;
  input b_48_;
  input b_49_;
  input b_50_;
  input b_51_;
  input b_52_;
  input b_53_;
  input b_54_;
  input b_55_;
  input b_56_;
  input b_57_;
  input b_58_;
  input b_59_;
  input b_60_;
  input b_61_;
  input b_62_;
  input b_63_;
  input b_64_;
  input b_65_;
  input b_66_;
  input b_67_;
  input b_68_;
  input b_69_;
  input b_70_;
  input b_71_;
  input b_72_;
  input b_73_;
  input b_74_;
  input b_75_;
  input b_76_;
  input b_77_;
  input b_78_;
  input b_79_;
  input b_80_;
  input b_81_;
  input b_82_;
  input b_83_;
  input b_84_;
  input b_85_;
  input b_86_;
  input b_87_;
  input b_88_;
  input b_89_;
  input b_90_;
  input b_91_;
  input b_92_;
  input b_93_;
  input b_94_;
  input b_95_;
  input b_96_;
  input b_97_;
  input b_98_;
  input b_99_;
  input b_100_;
  input b_101_;
  input b_102_;
  input b_103_;
  input b_104_;
  input b_105_;
  input b_106_;
  input b_107_;
  input b_108_;
  input b_109_;
  input b_110_;
  input b_111_;
  input b_112_;
  input b_113_;
  input b_114_;
  input b_115_;
  input b_116_;
  input b_117_;
  input b_118_;
  input b_119_;
  input b_120_;
  input b_121_;
  input b_122_;
  input b_123_;
  input b_124_;
  input b_125_;
  input b_126_;
  input b_127_;
  output f_0_;
  output f_1_;
  output f_2_;
  output f_3_;
  output f_4_;
  output f_5_;
  output f_6_;
  output f_7_;
  output f_8_;
  output f_9_;
  output f_10_;
  output f_11_;
  output f_12_;
  output f_13_;
  output f_14_;
  output f_15_;
  output f_16_;
  output f_17_;
  output f_18_;
  output f_19_;
  output f_20_;
  output f_21_;
  output f_22_;
  output f_23_;
  output f_24_;
  output f_25_;
  output f_26_;
  output f_27_;
  output f_28_;
  output f_29_;
  output f_30_;
  output f_31_;
  output f_32_;
  output f_33_;
  output f_34_;
  output f_35_;
  output f_36_;
  output f_37_;
  output f_38_;
  output f_39_;
  output f_40_;
  output f_41_;
  output f_42_;
  output f_43_;
  output f_44_;
  output f_45_;
  output f_46_;
  output f_47_;
  output f_48_;
  output f_49_;
  output f_50_;
  output f_51_;
  output f_52_;
  output f_53_;
  output f_54_;
  output f_55_;
  output f_56_;
  output f_57_;
  output f_58_;
  output f_59_;
  output f_60_;
  output f_61_;
  output f_62_;
  output f_63_;
  output f_64_;
  output f_65_;
  output f_66_;
  output f_67_;
  output f_68_;
  output f_69_;
  output f_70_;
  output f_71_;
  output f_72_;
  output f_73_;
  output f_74_;
  output f_75_;
  output f_76_;
  output f_77_;
  output f_78_;
  output f_79_;
  output f_80_;
  output f_81_;
  output f_82_;
  output f_83_;
  output f_84_;
  output f_85_;
  output f_86_;
  output f_87_;
  output f_88_;
  output f_89_;
  output f_90_;
  output f_91_;
  output f_92_;
  output f_93_;
  output f_94_;
  output f_95_;
  output f_96_;
  output f_97_;
  output f_98_;
  output f_99_;
  output f_100_;
  output f_101_;
  output f_102_;
  output f_103_;
  output f_104_;
  output f_105_;
  output f_106_;
  output f_107_;
  output f_108_;
  output f_109_;
  output f_110_;
  output f_111_;
  output f_112_;
  output f_113_;
  output f_114_;
  output f_115_;
  output f_116_;
  output f_117_;
  output f_118_;
  output f_119_;
  output f_120_;
  output f_121_;
  output f_122_;
  output f_123_;
  output f_124_;
  output f_125_;
  output f_126_;
  output f_127_;
  output cOut;
  AND2X2 n_n0 (
    .A1(a_0_),
    .A2(b_0_),
    .Z(f_0_)
  );
  OAI21X1 n_n1 (
    .A1(a_0_),
    .A2(b_0_),
    .A3(n392),
    .Z(f_1_)
  );
  AOI21X1 n_n2 (
    .A1(n391),
    .A2(n396),
    .A3(n400),
    .Z(f_2_)
  );
  AOI21X1 n_n3 (
    .A1(n399),
    .A2(n404),
    .A3(n408),
    .Z(f_3_)
  );
  AOI21X1 n_n4 (
    .A1(n407),
    .A2(n412),
    .A3(n416),
    .Z(f_4_)
  );
  AOI21X1 n_n5 (
    .A1(n415),
    .A2(n420),
    .A3(n424),
    .Z(f_5_)
  );
  AOI21X1 n_n6 (
    .A1(n423),
    .A2(n428),
    .A3(n432),
    .Z(f_6_)
  );
  AOI21X1 n_n7 (
    .A1(n431),
    .A2(n436),
    .A3(n440),
    .Z(f_7_)
  );
  AOI21X1 n_n8 (
    .A1(n439),
    .A2(n444),
    .A3(n448),
    .Z(f_8_)
  );
  AOI21X1 n_n9 (
    .A1(n447),
    .A2(n452),
    .A3(n456),
    .Z(f_9_)
  );
  AOI21X1 n_n10 (
    .A1(n455),
    .A2(n460),
    .A3(n464),
    .Z(f_10_)
  );
  AOI21X1 n_n11 (
    .A1(n463),
    .A2(n468),
    .A3(n472),
    .Z(f_11_)
  );
  AOI21X1 n_n12 (
    .A1(n471),
    .A2(n476),
    .A3(n480),
    .Z(f_12_)
  );
  AOI21X1 n_n13 (
    .A1(n479),
    .A2(n484),
    .A3(n488),
    .Z(f_13_)
  );
  AOI21X1 n_n14 (
    .A1(n487),
    .A2(n492),
    .A3(n496),
    .Z(f_14_)
  );
  AOI21X1 n_n15 (
    .A1(n495),
    .A2(n500),
    .A3(n504),
    .Z(f_15_)
  );
  AOI21X1 n_n16 (
    .A1(n503),
    .A2(n508),
    .A3(n512),
    .Z(f_16_)
  );
  AOI21X1 n_n17 (
    .A1(n511),
    .A2(n516),
    .A3(n520),
    .Z(f_17_)
  );
  AOI21X1 n_n18 (
    .A1(n519),
    .A2(n524),
    .A3(n528),
    .Z(f_18_)
  );
  AOI21X1 n_n19 (
    .A1(n527),
    .A2(n532),
    .A3(n536),
    .Z(f_19_)
  );
  AOI21X1 n_n20 (
    .A1(n535),
    .A2(n540),
    .A3(n544),
    .Z(f_20_)
  );
  AOI21X1 n_n21 (
    .A1(n543),
    .A2(n548),
    .A3(n552),
    .Z(f_21_)
  );
  AOI21X1 n_n22 (
    .A1(n551),
    .A2(n556),
    .A3(n560),
    .Z(f_22_)
  );
  AOI21X1 n_n23 (
    .A1(n559),
    .A2(n564),
    .A3(n568),
    .Z(f_23_)
  );
  AOI21X1 n_n24 (
    .A1(n567),
    .A2(n572),
    .A3(n576),
    .Z(f_24_)
  );
  AOI21X1 n_n25 (
    .A1(n575),
    .A2(n580),
    .A3(n584),
    .Z(f_25_)
  );
  AOI21X1 n_n26 (
    .A1(n583),
    .A2(n588),
    .A3(n592),
    .Z(f_26_)
  );
  AOI21X1 n_n27 (
    .A1(n591),
    .A2(n596),
    .A3(n600),
    .Z(f_27_)
  );
  AOI21X1 n_n28 (
    .A1(n599),
    .A2(n604),
    .A3(n608),
    .Z(f_28_)
  );
  AOI21X1 n_n29 (
    .A1(n607),
    .A2(n612),
    .A3(n616),
    .Z(f_29_)
  );
  AOI21X1 n_n30 (
    .A1(n615),
    .A2(n620),
    .A3(n624),
    .Z(f_30_)
  );
  AOI21X1 n_n31 (
    .A1(n623),
    .A2(n628),
    .A3(n632),
    .Z(f_31_)
  );
  AOI21X1 n_n32 (
    .A1(n631),
    .A2(n636),
    .A3(n640),
    .Z(f_32_)
  );
  AOI21X1 n_n33 (
    .A1(n639),
    .A2(n644),
    .A3(n648),
    .Z(f_33_)
  );
  AOI21X1 n_n34 (
    .A1(n647),
    .A2(n652),
    .A3(n656),
    .Z(f_34_)
  );
  AOI21X1 n_n35 (
    .A1(n655),
    .A2(n660),
    .A3(n664),
    .Z(f_35_)
  );
  AOI21X1 n_n36 (
    .A1(n663),
    .A2(n668),
    .A3(n672),
    .Z(f_36_)
  );
  AOI21X1 n_n37 (
    .A1(n671),
    .A2(n676),
    .A3(n680),
    .Z(f_37_)
  );
  AOI21X1 n_n38 (
    .A1(n679),
    .A2(n684),
    .A3(n688),
    .Z(f_38_)
  );
  AOI21X1 n_n39 (
    .A1(n687),
    .A2(n692),
    .A3(n696),
    .Z(f_39_)
  );
  AOI21X1 n_n40 (
    .A1(n695),
    .A2(n700),
    .A3(n704),
    .Z(f_40_)
  );
  AOI21X1 n_n41 (
    .A1(n703),
    .A2(n708),
    .A3(n712),
    .Z(f_41_)
  );
  AOI21X1 n_n42 (
    .A1(n711),
    .A2(n716),
    .A3(n720),
    .Z(f_42_)
  );
  AOI21X1 n_n43 (
    .A1(n719),
    .A2(n724),
    .A3(n728),
    .Z(f_43_)
  );
  AOI21X1 n_n44 (
    .A1(n727),
    .A2(n732),
    .A3(n736),
    .Z(f_44_)
  );
  AOI21X1 n_n45 (
    .A1(n735),
    .A2(n740),
    .A3(n744),
    .Z(f_45_)
  );
  AOI21X1 n_n46 (
    .A1(n743),
    .A2(n748),
    .A3(n752),
    .Z(f_46_)
  );
  AOI21X1 n_n47 (
    .A1(n751),
    .A2(n756),
    .A3(n760),
    .Z(f_47_)
  );
  AOI21X1 n_n48 (
    .A1(n759),
    .A2(n764),
    .A3(n768),
    .Z(f_48_)
  );
  AOI21X1 n_n49 (
    .A1(n767),
    .A2(n772),
    .A3(n776),
    .Z(f_49_)
  );
  AOI21X1 n_n50 (
    .A1(n775),
    .A2(n780),
    .A3(n784),
    .Z(f_50_)
  );
  AOI21X1 n_n51 (
    .A1(n783),
    .A2(n788),
    .A3(n792),
    .Z(f_51_)
  );
  AOI21X1 n_n52 (
    .A1(n791),
    .A2(n796),
    .A3(n800),
    .Z(f_52_)
  );
  AOI21X1 n_n53 (
    .A1(n799),
    .A2(n804),
    .A3(n808),
    .Z(f_53_)
  );
  AOI21X1 n_n54 (
    .A1(n807),
    .A2(n812),
    .A3(n816),
    .Z(f_54_)
  );
  AOI21X1 n_n55 (
    .A1(n815),
    .A2(n820),
    .A3(n824),
    .Z(f_55_)
  );
  AOI21X1 n_n56 (
    .A1(n823),
    .A2(n828),
    .A3(n832),
    .Z(f_56_)
  );
  AOI21X1 n_n57 (
    .A1(n831),
    .A2(n836),
    .A3(n840),
    .Z(f_57_)
  );
  AOI21X1 n_n58 (
    .A1(n839),
    .A2(n844),
    .A3(n848),
    .Z(f_58_)
  );
  AOI21X1 n_n59 (
    .A1(n847),
    .A2(n852),
    .A3(n856),
    .Z(f_59_)
  );
  AOI21X1 n_n60 (
    .A1(n855),
    .A2(n860),
    .A3(n864),
    .Z(f_60_)
  );
  AOI21X1 n_n61 (
    .A1(n863),
    .A2(n868),
    .A3(n872),
    .Z(f_61_)
  );
  AOI21X1 n_n62 (
    .A1(n871),
    .A2(n876),
    .A3(n880),
    .Z(f_62_)
  );
  AOI21X1 n_n63 (
    .A1(n879),
    .A2(n884),
    .A3(n888),
    .Z(f_63_)
  );
  AOI21X1 n_n64 (
    .A1(n887),
    .A2(n892),
    .A3(n896),
    .Z(f_64_)
  );
  AOI21X1 n_n65 (
    .A1(n895),
    .A2(n900),
    .A3(n904),
    .Z(f_65_)
  );
  AOI21X1 n_n66 (
    .A1(n903),
    .A2(n908),
    .A3(n912),
    .Z(f_66_)
  );
  AOI21X1 n_n67 (
    .A1(n911),
    .A2(n916),
    .A3(n920),
    .Z(f_67_)
  );
  AOI21X1 n_n68 (
    .A1(n919),
    .A2(n924),
    .A3(n928),
    .Z(f_68_)
  );
  AOI21X1 n_n69 (
    .A1(n927),
    .A2(n932),
    .A3(n936),
    .Z(f_69_)
  );
  AOI21X1 n_n70 (
    .A1(n935),
    .A2(n940),
    .A3(n944),
    .Z(f_70_)
  );
  AOI21X1 n_n71 (
    .A1(n943),
    .A2(n948),
    .A3(n952),
    .Z(f_71_)
  );
  AOI21X1 n_n72 (
    .A1(n951),
    .A2(n956),
    .A3(n960),
    .Z(f_72_)
  );
  AOI21X1 n_n73 (
    .A1(n959),
    .A2(n964),
    .A3(n968),
    .Z(f_73_)
  );
  AOI21X1 n_n74 (
    .A1(n967),
    .A2(n972),
    .A3(n976),
    .Z(f_74_)
  );
  AOI21X1 n_n75 (
    .A1(n975),
    .A2(n980),
    .A3(n984),
    .Z(f_75_)
  );
  AOI21X1 n_n76 (
    .A1(n983),
    .A2(n988),
    .A3(n992),
    .Z(f_76_)
  );
  OAI21X1 n_n77 (
    .A1(n1000),
    .A2(n991),
    .A3(n996),
    .Z(f_77_)
  );
  OAI21X1 n_n78 (
    .A1(n1004),
    .A2(n1008),
    .A3(n999),
    .Z(f_78_)
  );
  AOI21X1 n_n79 (
    .A1(n1007),
    .A2(n1012),
    .A3(n1016),
    .Z(f_79_)
  );
  AOI21X1 n_n80 (
    .A1(n1015),
    .A2(n1020),
    .A3(n1024),
    .Z(f_80_)
  );
  AOI21X1 n_n81 (
    .A1(n1023),
    .A2(n1028),
    .A3(n1032),
    .Z(f_81_)
  );
  AOI21X1 n_n82 (
    .A1(n1031),
    .A2(n1036),
    .A3(n1040),
    .Z(f_82_)
  );
  AOI21X1 n_n83 (
    .A1(n1039),
    .A2(n1044),
    .A3(n1048),
    .Z(f_83_)
  );
  AOI21X1 n_n84 (
    .A1(n1047),
    .A2(n1052),
    .A3(n1056),
    .Z(f_84_)
  );
  AOI21X1 n_n85 (
    .A1(n1055),
    .A2(n1060),
    .A3(n1064),
    .Z(f_85_)
  );
  AOI21X1 n_n86 (
    .A1(n1063),
    .A2(n1068),
    .A3(n1072),
    .Z(f_86_)
  );
  AOI21X1 n_n87 (
    .A1(n1071),
    .A2(n1076),
    .A3(n1080),
    .Z(f_87_)
  );
  AOI21X1 n_n88 (
    .A1(n1079),
    .A2(n1084),
    .A3(n1088),
    .Z(f_88_)
  );
  AOI21X1 n_n89 (
    .A1(n1087),
    .A2(n1092),
    .A3(n1096),
    .Z(f_89_)
  );
  AOI21X1 n_n90 (
    .A1(n1095),
    .A2(n1100),
    .A3(n1104),
    .Z(f_90_)
  );
  AOI21X1 n_n91 (
    .A1(n1103),
    .A2(n1108),
    .A3(n1112),
    .Z(f_91_)
  );
  AOI21X1 n_n92 (
    .A1(n1111),
    .A2(n1116),
    .A3(n1120),
    .Z(f_92_)
  );
  AOI21X1 n_n93 (
    .A1(n1119),
    .A2(n1124),
    .A3(n1128),
    .Z(f_93_)
  );
  AOI21X1 n_n94 (
    .A1(n1127),
    .A2(n1132),
    .A3(n1136),
    .Z(f_94_)
  );
  AOI21X1 n_n95 (
    .A1(n1135),
    .A2(n1140),
    .A3(n1144),
    .Z(f_95_)
  );
  AOI21X1 n_n96 (
    .A1(n1143),
    .A2(n1148),
    .A3(n1152),
    .Z(f_96_)
  );
  AOI21X1 n_n97 (
    .A1(n1151),
    .A2(n1156),
    .A3(n1160),
    .Z(f_97_)
  );
  AOI21X1 n_n98 (
    .A1(n1159),
    .A2(n1164),
    .A3(n1168),
    .Z(f_98_)
  );
  AOI21X1 n_n99 (
    .A1(n1167),
    .A2(n1172),
    .A3(n1176),
    .Z(f_99_)
  );
  AOI21X1 n_n100 (
    .A1(n1175),
    .A2(n1180),
    .A3(n1184),
    .Z(f_100_)
  );
  AOI21X1 n_n101 (
    .A1(n1183),
    .A2(n1188),
    .A3(n1192),
    .Z(f_101_)
  );
  AOI21X1 n_n102 (
    .A1(n1191),
    .A2(n1196),
    .A3(n1200),
    .Z(f_102_)
  );
  AOI21X1 n_n103 (
    .A1(n1199),
    .A2(n1204),
    .A3(n1208),
    .Z(f_103_)
  );
  AOI21X1 n_n104 (
    .A1(n1207),
    .A2(n1212),
    .A3(n1216),
    .Z(f_104_)
  );
  AOI21X1 n_n105 (
    .A1(n1215),
    .A2(n1220),
    .A3(n1224),
    .Z(f_105_)
  );
  AOI21X1 n_n106 (
    .A1(n1223),
    .A2(n1228),
    .A3(n1232),
    .Z(f_106_)
  );
  AOI21X1 n_n107 (
    .A1(n1231),
    .A2(n1236),
    .A3(n1240),
    .Z(f_107_)
  );
  AOI21X1 n_n108 (
    .A1(n1239),
    .A2(n1244),
    .A3(n1248),
    .Z(f_108_)
  );
  AOI21X1 n_n109 (
    .A1(n1247),
    .A2(n1252),
    .A3(n1256),
    .Z(f_109_)
  );
  AOI21X1 n_n110 (
    .A1(n1255),
    .A2(n1260),
    .A3(n1264),
    .Z(f_110_)
  );
  AOI21X1 n_n111 (
    .A1(n1263),
    .A2(n1268),
    .A3(n1272),
    .Z(f_111_)
  );
  AOI21X1 n_n112 (
    .A1(n1271),
    .A2(n1276),
    .A3(n1280),
    .Z(f_112_)
  );
  AOI21X1 n_n113 (
    .A1(n1279),
    .A2(n1284),
    .A3(n1288),
    .Z(f_113_)
  );
  AOI21X1 n_n114 (
    .A1(n1287),
    .A2(n1292),
    .A3(n1296),
    .Z(f_114_)
  );
  AOI21X1 n_n115 (
    .A1(n1295),
    .A2(n1300),
    .A3(n1304),
    .Z(f_115_)
  );
  AOI21X1 n_n116 (
    .A1(n1303),
    .A2(n1308),
    .A3(n1312),
    .Z(f_116_)
  );
  AOI21X1 n_n117 (
    .A1(n1311),
    .A2(n1316),
    .A3(n1320),
    .Z(f_117_)
  );
  AOI21X1 n_n118 (
    .A1(n1319),
    .A2(n1324),
    .A3(n1328),
    .Z(f_118_)
  );
  AOI21X1 n_n119 (
    .A1(n1327),
    .A2(n1332),
    .A3(n1336),
    .Z(f_119_)
  );
  AOI21X1 n_n120 (
    .A1(n1335),
    .A2(n1340),
    .A3(n1344),
    .Z(f_120_)
  );
  AOI21X1 n_n121 (
    .A1(n1343),
    .A2(n1348),
    .A3(n1352),
    .Z(f_121_)
  );
  AOI21X1 n_n122 (
    .A1(n1351),
    .A2(n1356),
    .A3(n1360),
    .Z(f_122_)
  );
  AOI21X1 n_n123 (
    .A1(n1359),
    .A2(n1364),
    .A3(n1368),
    .Z(f_123_)
  );
  AOI21X1 n_n124 (
    .A1(n1367),
    .A2(n1372),
    .A3(n1376),
    .Z(f_124_)
  );
  AOI21X1 n_n125 (
    .A1(n1375),
    .A2(n1380),
    .A3(n1384),
    .Z(f_125_)
  );
  AOI21X1 n_n126 (
    .A1(n1383),
    .A2(n1388),
    .A3(n1392),
    .Z(f_126_)
  );
  AOI21X1 n_n127 (
    .A1(n1391),
    .A2(n1396),
    .A3(n1400),
    .Z(f_127_)
  );
  AOI21X1 n_n128 (
    .A1(n1397),
    .A2(n1398),
    .A3(n1399),
    .Z(cOut)
  );
  XOR2X1 n_n129 (
    .A1(a_1_),
    .A2(b_1_),
    .Z(n392)
  );
  AND2X2 n_n130 (
    .A1(a_1_),
    .A2(b_1_),
    .Z(n391)
  );
  OAI21X1 n_n131 (
    .A1(a_0_),
    .A2(b_0_),
    .A3(n390),
    .Z(n396)
  );
  XOR2X1 n_n132 (
    .A1(a_2_),
    .A2(b_2_),
    .Z(n400)
  );
  AND2X2 n_n133 (
    .A1(a_2_),
    .A2(b_2_),
    .Z(n399)
  );
  AOI22X1 n_n134 (
    .A1(a_2_),
    .A2(b_2_),
    .A3(n391),
    .A4(n396),
    .Z(n404)
  );
  XOR2X1 n_n135 (
    .A1(a_3_),
    .A2(b_3_),
    .Z(n408)
  );
  AND2X2 n_n136 (
    .A1(a_3_),
    .A2(b_3_),
    .Z(n407)
  );
  AOI22X1 n_n137 (
    .A1(a_3_),
    .A2(b_3_),
    .A3(n399),
    .A4(n404),
    .Z(n412)
  );
  XOR2X1 n_n138 (
    .A1(a_4_),
    .A2(b_4_),
    .Z(n416)
  );
  AND2X2 n_n139 (
    .A1(a_4_),
    .A2(b_4_),
    .Z(n415)
  );
  AOI22X1 n_n140 (
    .A1(a_4_),
    .A2(b_4_),
    .A3(n407),
    .A4(n412),
    .Z(n420)
  );
  XOR2X1 n_n141 (
    .A1(a_5_),
    .A2(b_5_),
    .Z(n424)
  );
  AND2X2 n_n142 (
    .A1(a_5_),
    .A2(b_5_),
    .Z(n423)
  );
  AOI22X1 n_n143 (
    .A1(a_5_),
    .A2(b_5_),
    .A3(n415),
    .A4(n420),
    .Z(n428)
  );
  XOR2X1 n_n144 (
    .A1(a_6_),
    .A2(b_6_),
    .Z(n432)
  );
  AND2X2 n_n145 (
    .A1(a_6_),
    .A2(b_6_),
    .Z(n431)
  );
  AOI22X1 n_n146 (
    .A1(a_6_),
    .A2(b_6_),
    .A3(n423),
    .A4(n428),
    .Z(n436)
  );
  XOR2X1 n_n147 (
    .A1(a_7_),
    .A2(b_7_),
    .Z(n440)
  );
  AND2X2 n_n148 (
    .A1(a_7_),
    .A2(b_7_),
    .Z(n439)
  );
  AOI22X1 n_n149 (
    .A1(a_7_),
    .A2(b_7_),
    .A3(n431),
    .A4(n436),
    .Z(n444)
  );
  XOR2X1 n_n150 (
    .A1(a_8_),
    .A2(b_8_),
    .Z(n448)
  );
  AND2X2 n_n151 (
    .A1(a_8_),
    .A2(b_8_),
    .Z(n447)
  );
  AOI22X1 n_n152 (
    .A1(a_8_),
    .A2(b_8_),
    .A3(n439),
    .A4(n444),
    .Z(n452)
  );
  XOR2X1 n_n153 (
    .A1(a_9_),
    .A2(b_9_),
    .Z(n456)
  );
  AND2X2 n_n154 (
    .A1(a_9_),
    .A2(b_9_),
    .Z(n455)
  );
  AOI22X1 n_n155 (
    .A1(a_9_),
    .A2(b_9_),
    .A3(n447),
    .A4(n452),
    .Z(n460)
  );
  XOR2X1 n_n156 (
    .A1(a_10_),
    .A2(b_10_),
    .Z(n464)
  );
  AND2X2 n_n157 (
    .A1(a_10_),
    .A2(b_10_),
    .Z(n463)
  );
  AOI22X1 n_n158 (
    .A1(a_10_),
    .A2(b_10_),
    .A3(n455),
    .A4(n460),
    .Z(n468)
  );
  XOR2X1 n_n159 (
    .A1(a_11_),
    .A2(b_11_),
    .Z(n472)
  );
  AND2X2 n_n160 (
    .A1(a_11_),
    .A2(b_11_),
    .Z(n471)
  );
  AOI22X1 n_n161 (
    .A1(a_11_),
    .A2(b_11_),
    .A3(n463),
    .A4(n468),
    .Z(n476)
  );
  XOR2X1 n_n162 (
    .A1(a_12_),
    .A2(b_12_),
    .Z(n480)
  );
  AND2X2 n_n163 (
    .A1(a_12_),
    .A2(b_12_),
    .Z(n479)
  );
  AOI22X1 n_n164 (
    .A1(a_12_),
    .A2(b_12_),
    .A3(n471),
    .A4(n476),
    .Z(n484)
  );
  XOR2X1 n_n165 (
    .A1(a_13_),
    .A2(b_13_),
    .Z(n488)
  );
  AND2X2 n_n166 (
    .A1(a_13_),
    .A2(b_13_),
    .Z(n487)
  );
  AOI22X1 n_n167 (
    .A1(a_13_),
    .A2(b_13_),
    .A3(n479),
    .A4(n484),
    .Z(n492)
  );
  XOR2X1 n_n168 (
    .A1(a_14_),
    .A2(b_14_),
    .Z(n496)
  );
  AND2X2 n_n169 (
    .A1(a_14_),
    .A2(b_14_),
    .Z(n495)
  );
  AOI22X1 n_n170 (
    .A1(a_14_),
    .A2(b_14_),
    .A3(n487),
    .A4(n492),
    .Z(n500)
  );
  XOR2X1 n_n171 (
    .A1(a_15_),
    .A2(b_15_),
    .Z(n504)
  );
  AND2X2 n_n172 (
    .A1(a_15_),
    .A2(b_15_),
    .Z(n503)
  );
  AOI22X1 n_n173 (
    .A1(a_15_),
    .A2(b_15_),
    .A3(n495),
    .A4(n500),
    .Z(n508)
  );
  XOR2X1 n_n174 (
    .A1(a_16_),
    .A2(b_16_),
    .Z(n512)
  );
  AND2X2 n_n175 (
    .A1(a_16_),
    .A2(b_16_),
    .Z(n511)
  );
  AOI22X1 n_n176 (
    .A1(a_16_),
    .A2(b_16_),
    .A3(n503),
    .A4(n508),
    .Z(n516)
  );
  XOR2X1 n_n177 (
    .A1(a_17_),
    .A2(b_17_),
    .Z(n520)
  );
  AND2X2 n_n178 (
    .A1(a_17_),
    .A2(b_17_),
    .Z(n519)
  );
  AOI22X1 n_n179 (
    .A1(a_17_),
    .A2(b_17_),
    .A3(n511),
    .A4(n516),
    .Z(n524)
  );
  XOR2X1 n_n180 (
    .A1(a_18_),
    .A2(b_18_),
    .Z(n528)
  );
  AND2X2 n_n181 (
    .A1(a_18_),
    .A2(b_18_),
    .Z(n527)
  );
  AOI22X1 n_n182 (
    .A1(a_18_),
    .A2(b_18_),
    .A3(n519),
    .A4(n524),
    .Z(n532)
  );
  XOR2X1 n_n183 (
    .A1(a_19_),
    .A2(b_19_),
    .Z(n536)
  );
  AND2X2 n_n184 (
    .A1(a_19_),
    .A2(b_19_),
    .Z(n535)
  );
  AOI22X1 n_n185 (
    .A1(a_19_),
    .A2(b_19_),
    .A3(n527),
    .A4(n532),
    .Z(n540)
  );
  XOR2X1 n_n186 (
    .A1(a_20_),
    .A2(b_20_),
    .Z(n544)
  );
  AND2X2 n_n187 (
    .A1(a_20_),
    .A2(b_20_),
    .Z(n543)
  );
  AOI22X1 n_n188 (
    .A1(a_20_),
    .A2(b_20_),
    .A3(n535),
    .A4(n540),
    .Z(n548)
  );
  XOR2X1 n_n189 (
    .A1(a_21_),
    .A2(b_21_),
    .Z(n552)
  );
  AND2X2 n_n190 (
    .A1(a_21_),
    .A2(b_21_),
    .Z(n551)
  );
  AOI22X1 n_n191 (
    .A1(a_21_),
    .A2(b_21_),
    .A3(n543),
    .A4(n548),
    .Z(n556)
  );
  XOR2X1 n_n192 (
    .A1(a_22_),
    .A2(b_22_),
    .Z(n560)
  );
  AND2X2 n_n193 (
    .A1(a_22_),
    .A2(b_22_),
    .Z(n559)
  );
  AOI22X1 n_n194 (
    .A1(a_22_),
    .A2(b_22_),
    .A3(n551),
    .A4(n556),
    .Z(n564)
  );
  XOR2X1 n_n195 (
    .A1(a_23_),
    .A2(b_23_),
    .Z(n568)
  );
  AND2X2 n_n196 (
    .A1(a_23_),
    .A2(b_23_),
    .Z(n567)
  );
  AOI22X1 n_n197 (
    .A1(a_23_),
    .A2(b_23_),
    .A3(n559),
    .A4(n564),
    .Z(n572)
  );
  XOR2X1 n_n198 (
    .A1(a_24_),
    .A2(b_24_),
    .Z(n576)
  );
  AND2X2 n_n199 (
    .A1(a_24_),
    .A2(b_24_),
    .Z(n575)
  );
  AOI22X1 n_n200 (
    .A1(a_24_),
    .A2(b_24_),
    .A3(n567),
    .A4(n572),
    .Z(n580)
  );
  XOR2X1 n_n201 (
    .A1(a_25_),
    .A2(b_25_),
    .Z(n584)
  );
  AND2X2 n_n202 (
    .A1(a_25_),
    .A2(b_25_),
    .Z(n583)
  );
  AOI22X1 n_n203 (
    .A1(a_25_),
    .A2(b_25_),
    .A3(n575),
    .A4(n580),
    .Z(n588)
  );
  XOR2X1 n_n204 (
    .A1(a_26_),
    .A2(b_26_),
    .Z(n592)
  );
  AND2X2 n_n205 (
    .A1(a_26_),
    .A2(b_26_),
    .Z(n591)
  );
  AOI22X1 n_n206 (
    .A1(a_26_),
    .A2(b_26_),
    .A3(n583),
    .A4(n588),
    .Z(n596)
  );
  XOR2X1 n_n207 (
    .A1(a_27_),
    .A2(b_27_),
    .Z(n600)
  );
  AND2X2 n_n208 (
    .A1(a_27_),
    .A2(b_27_),
    .Z(n599)
  );
  AOI22X1 n_n209 (
    .A1(a_27_),
    .A2(b_27_),
    .A3(n591),
    .A4(n596),
    .Z(n604)
  );
  XOR2X1 n_n210 (
    .A1(a_28_),
    .A2(b_28_),
    .Z(n608)
  );
  AND2X2 n_n211 (
    .A1(a_28_),
    .A2(b_28_),
    .Z(n607)
  );
  AOI22X1 n_n212 (
    .A1(a_28_),
    .A2(b_28_),
    .A3(n599),
    .A4(n604),
    .Z(n612)
  );
  XOR2X1 n_n213 (
    .A1(a_29_),
    .A2(b_29_),
    .Z(n616)
  );
  AND2X2 n_n214 (
    .A1(a_29_),
    .A2(b_29_),
    .Z(n615)
  );
  AOI22X1 n_n215 (
    .A1(a_29_),
    .A2(b_29_),
    .A3(n607),
    .A4(n612),
    .Z(n620)
  );
  XOR2X1 n_n216 (
    .A1(a_30_),
    .A2(b_30_),
    .Z(n624)
  );
  AND2X2 n_n217 (
    .A1(a_30_),
    .A2(b_30_),
    .Z(n623)
  );
  AOI22X1 n_n218 (
    .A1(a_30_),
    .A2(b_30_),
    .A3(n615),
    .A4(n620),
    .Z(n628)
  );
  XOR2X1 n_n219 (
    .A1(a_31_),
    .A2(b_31_),
    .Z(n632)
  );
  AND2X2 n_n220 (
    .A1(a_31_),
    .A2(b_31_),
    .Z(n631)
  );
  AOI22X1 n_n221 (
    .A1(a_31_),
    .A2(b_31_),
    .A3(n623),
    .A4(n628),
    .Z(n636)
  );
  XOR2X1 n_n222 (
    .A1(a_32_),
    .A2(b_32_),
    .Z(n640)
  );
  AND2X2 n_n223 (
    .A1(a_32_),
    .A2(b_32_),
    .Z(n639)
  );
  AOI22X1 n_n224 (
    .A1(a_32_),
    .A2(b_32_),
    .A3(n631),
    .A4(n636),
    .Z(n644)
  );
  XOR2X1 n_n225 (
    .A1(a_33_),
    .A2(b_33_),
    .Z(n648)
  );
  AND2X2 n_n226 (
    .A1(a_33_),
    .A2(b_33_),
    .Z(n647)
  );
  AOI22X1 n_n227 (
    .A1(a_33_),
    .A2(b_33_),
    .A3(n639),
    .A4(n644),
    .Z(n652)
  );
  XOR2X1 n_n228 (
    .A1(a_34_),
    .A2(b_34_),
    .Z(n656)
  );
  AND2X2 n_n229 (
    .A1(a_34_),
    .A2(b_34_),
    .Z(n655)
  );
  AOI22X1 n_n230 (
    .A1(a_34_),
    .A2(b_34_),
    .A3(n647),
    .A4(n652),
    .Z(n660)
  );
  XOR2X1 n_n231 (
    .A1(a_35_),
    .A2(b_35_),
    .Z(n664)
  );
  AND2X2 n_n232 (
    .A1(a_35_),
    .A2(b_35_),
    .Z(n663)
  );
  AOI22X1 n_n233 (
    .A1(a_35_),
    .A2(b_35_),
    .A3(n655),
    .A4(n660),
    .Z(n668)
  );
  XOR2X1 n_n234 (
    .A1(a_36_),
    .A2(b_36_),
    .Z(n672)
  );
  AND2X2 n_n235 (
    .A1(a_36_),
    .A2(b_36_),
    .Z(n671)
  );
  AOI22X1 n_n236 (
    .A1(a_36_),
    .A2(b_36_),
    .A3(n663),
    .A4(n668),
    .Z(n676)
  );
  XOR2X1 n_n237 (
    .A1(a_37_),
    .A2(b_37_),
    .Z(n680)
  );
  AND2X2 n_n238 (
    .A1(a_37_),
    .A2(b_37_),
    .Z(n679)
  );
  AOI22X1 n_n239 (
    .A1(a_37_),
    .A2(b_37_),
    .A3(n671),
    .A4(n676),
    .Z(n684)
  );
  XOR2X1 n_n240 (
    .A1(a_38_),
    .A2(b_38_),
    .Z(n688)
  );
  AND2X2 n_n241 (
    .A1(a_38_),
    .A2(b_38_),
    .Z(n687)
  );
  AOI22X1 n_n242 (
    .A1(a_38_),
    .A2(b_38_),
    .A3(n679),
    .A4(n684),
    .Z(n692)
  );
  XOR2X1 n_n243 (
    .A1(a_39_),
    .A2(b_39_),
    .Z(n696)
  );
  AND2X2 n_n244 (
    .A1(a_39_),
    .A2(b_39_),
    .Z(n695)
  );
  AOI22X1 n_n245 (
    .A1(a_39_),
    .A2(b_39_),
    .A3(n687),
    .A4(n692),
    .Z(n700)
  );
  XOR2X1 n_n246 (
    .A1(a_40_),
    .A2(b_40_),
    .Z(n704)
  );
  AND2X2 n_n247 (
    .A1(a_40_),
    .A2(b_40_),
    .Z(n703)
  );
  AOI22X1 n_n248 (
    .A1(a_40_),
    .A2(b_40_),
    .A3(n695),
    .A4(n700),
    .Z(n708)
  );
  XOR2X1 n_n249 (
    .A1(a_41_),
    .A2(b_41_),
    .Z(n712)
  );
  AND2X2 n_n250 (
    .A1(a_41_),
    .A2(b_41_),
    .Z(n711)
  );
  AOI22X1 n_n251 (
    .A1(a_41_),
    .A2(b_41_),
    .A3(n703),
    .A4(n708),
    .Z(n716)
  );
  XOR2X1 n_n252 (
    .A1(a_42_),
    .A2(b_42_),
    .Z(n720)
  );
  AND2X2 n_n253 (
    .A1(a_42_),
    .A2(b_42_),
    .Z(n719)
  );
  AOI22X1 n_n254 (
    .A1(a_42_),
    .A2(b_42_),
    .A3(n711),
    .A4(n716),
    .Z(n724)
  );
  XOR2X1 n_n255 (
    .A1(a_43_),
    .A2(b_43_),
    .Z(n728)
  );
  AND2X2 n_n256 (
    .A1(a_43_),
    .A2(b_43_),
    .Z(n727)
  );
  AOI22X1 n_n257 (
    .A1(a_43_),
    .A2(b_43_),
    .A3(n719),
    .A4(n724),
    .Z(n732)
  );
  XOR2X1 n_n258 (
    .A1(a_44_),
    .A2(b_44_),
    .Z(n736)
  );
  AND2X2 n_n259 (
    .A1(a_44_),
    .A2(b_44_),
    .Z(n735)
  );
  AOI22X1 n_n260 (
    .A1(a_44_),
    .A2(b_44_),
    .A3(n727),
    .A4(n732),
    .Z(n740)
  );
  XOR2X1 n_n261 (
    .A1(a_45_),
    .A2(b_45_),
    .Z(n744)
  );
  AND2X2 n_n262 (
    .A1(a_45_),
    .A2(b_45_),
    .Z(n743)
  );
  AOI22X1 n_n263 (
    .A1(a_45_),
    .A2(b_45_),
    .A3(n735),
    .A4(n740),
    .Z(n748)
  );
  XOR2X1 n_n264 (
    .A1(a_46_),
    .A2(b_46_),
    .Z(n752)
  );
  AND2X2 n_n265 (
    .A1(a_46_),
    .A2(b_46_),
    .Z(n751)
  );
  AOI22X1 n_n266 (
    .A1(a_46_),
    .A2(b_46_),
    .A3(n743),
    .A4(n748),
    .Z(n756)
  );
  XOR2X1 n_n267 (
    .A1(a_47_),
    .A2(b_47_),
    .Z(n760)
  );
  AND2X2 n_n268 (
    .A1(a_47_),
    .A2(b_47_),
    .Z(n759)
  );
  AOI22X1 n_n269 (
    .A1(a_47_),
    .A2(b_47_),
    .A3(n751),
    .A4(n756),
    .Z(n764)
  );
  XOR2X1 n_n270 (
    .A1(a_48_),
    .A2(b_48_),
    .Z(n768)
  );
  AND2X2 n_n271 (
    .A1(a_48_),
    .A2(b_48_),
    .Z(n767)
  );
  AOI22X1 n_n272 (
    .A1(a_48_),
    .A2(b_48_),
    .A3(n759),
    .A4(n764),
    .Z(n772)
  );
  XOR2X1 n_n273 (
    .A1(a_49_),
    .A2(b_49_),
    .Z(n776)
  );
  AND2X2 n_n274 (
    .A1(a_49_),
    .A2(b_49_),
    .Z(n775)
  );
  AOI22X1 n_n275 (
    .A1(a_49_),
    .A2(b_49_),
    .A3(n767),
    .A4(n772),
    .Z(n780)
  );
  XOR2X1 n_n276 (
    .A1(a_50_),
    .A2(b_50_),
    .Z(n784)
  );
  AND2X2 n_n277 (
    .A1(a_50_),
    .A2(b_50_),
    .Z(n783)
  );
  AOI22X1 n_n278 (
    .A1(a_50_),
    .A2(b_50_),
    .A3(n775),
    .A4(n780),
    .Z(n788)
  );
  XOR2X1 n_n279 (
    .A1(a_51_),
    .A2(b_51_),
    .Z(n792)
  );
  AND2X2 n_n280 (
    .A1(a_51_),
    .A2(b_51_),
    .Z(n791)
  );
  AOI22X1 n_n281 (
    .A1(a_51_),
    .A2(b_51_),
    .A3(n783),
    .A4(n788),
    .Z(n796)
  );
  XOR2X1 n_n282 (
    .A1(a_52_),
    .A2(b_52_),
    .Z(n800)
  );
  AND2X2 n_n283 (
    .A1(a_52_),
    .A2(b_52_),
    .Z(n799)
  );
  AOI22X1 n_n284 (
    .A1(a_52_),
    .A2(b_52_),
    .A3(n791),
    .A4(n796),
    .Z(n804)
  );
  XOR2X1 n_n285 (
    .A1(a_53_),
    .A2(b_53_),
    .Z(n808)
  );
  AND2X2 n_n286 (
    .A1(a_53_),
    .A2(b_53_),
    .Z(n807)
  );
  AOI22X1 n_n287 (
    .A1(a_53_),
    .A2(b_53_),
    .A3(n799),
    .A4(n804),
    .Z(n812)
  );
  XOR2X1 n_n288 (
    .A1(a_54_),
    .A2(b_54_),
    .Z(n816)
  );
  AND2X2 n_n289 (
    .A1(a_54_),
    .A2(b_54_),
    .Z(n815)
  );
  AOI22X1 n_n290 (
    .A1(a_54_),
    .A2(b_54_),
    .A3(n807),
    .A4(n812),
    .Z(n820)
  );
  XOR2X1 n_n291 (
    .A1(a_55_),
    .A2(b_55_),
    .Z(n824)
  );
  AND2X2 n_n292 (
    .A1(a_55_),
    .A2(b_55_),
    .Z(n823)
  );
  AOI22X1 n_n293 (
    .A1(a_55_),
    .A2(b_55_),
    .A3(n815),
    .A4(n820),
    .Z(n828)
  );
  XOR2X1 n_n294 (
    .A1(a_56_),
    .A2(b_56_),
    .Z(n832)
  );
  AND2X2 n_n295 (
    .A1(a_56_),
    .A2(b_56_),
    .Z(n831)
  );
  AOI22X1 n_n296 (
    .A1(a_56_),
    .A2(b_56_),
    .A3(n823),
    .A4(n828),
    .Z(n836)
  );
  XOR2X1 n_n297 (
    .A1(a_57_),
    .A2(b_57_),
    .Z(n840)
  );
  AND2X2 n_n298 (
    .A1(a_57_),
    .A2(b_57_),
    .Z(n839)
  );
  AOI22X1 n_n299 (
    .A1(a_57_),
    .A2(b_57_),
    .A3(n831),
    .A4(n836),
    .Z(n844)
  );
  XOR2X1 n_n300 (
    .A1(a_58_),
    .A2(b_58_),
    .Z(n848)
  );
  AND2X2 n_n301 (
    .A1(a_58_),
    .A2(b_58_),
    .Z(n847)
  );
  AOI22X1 n_n302 (
    .A1(a_58_),
    .A2(b_58_),
    .A3(n839),
    .A4(n844),
    .Z(n852)
  );
  XOR2X1 n_n303 (
    .A1(a_59_),
    .A2(b_59_),
    .Z(n856)
  );
  AND2X2 n_n304 (
    .A1(a_59_),
    .A2(b_59_),
    .Z(n855)
  );
  AOI22X1 n_n305 (
    .A1(a_59_),
    .A2(b_59_),
    .A3(n847),
    .A4(n852),
    .Z(n860)
  );
  XOR2X1 n_n306 (
    .A1(a_60_),
    .A2(b_60_),
    .Z(n864)
  );
  AND2X2 n_n307 (
    .A1(a_60_),
    .A2(b_60_),
    .Z(n863)
  );
  AOI22X1 n_n308 (
    .A1(a_60_),
    .A2(b_60_),
    .A3(n855),
    .A4(n860),
    .Z(n868)
  );
  XOR2X1 n_n309 (
    .A1(a_61_),
    .A2(b_61_),
    .Z(n872)
  );
  AND2X2 n_n310 (
    .A1(a_61_),
    .A2(b_61_),
    .Z(n871)
  );
  AOI22X1 n_n311 (
    .A1(a_61_),
    .A2(b_61_),
    .A3(n863),
    .A4(n868),
    .Z(n876)
  );
  XOR2X1 n_n312 (
    .A1(a_62_),
    .A2(b_62_),
    .Z(n880)
  );
  AND2X2 n_n313 (
    .A1(a_62_),
    .A2(b_62_),
    .Z(n879)
  );
  AOI22X1 n_n314 (
    .A1(a_62_),
    .A2(b_62_),
    .A3(n871),
    .A4(n876),
    .Z(n884)
  );
  XOR2X1 n_n315 (
    .A1(a_63_),
    .A2(b_63_),
    .Z(n888)
  );
  AND2X2 n_n316 (
    .A1(a_63_),
    .A2(b_63_),
    .Z(n887)
  );
  AOI22X1 n_n317 (
    .A1(a_63_),
    .A2(b_63_),
    .A3(n879),
    .A4(n884),
    .Z(n892)
  );
  XOR2X1 n_n318 (
    .A1(a_64_),
    .A2(b_64_),
    .Z(n896)
  );
  AND2X2 n_n319 (
    .A1(a_64_),
    .A2(b_64_),
    .Z(n895)
  );
  AOI22X1 n_n320 (
    .A1(a_64_),
    .A2(b_64_),
    .A3(n887),
    .A4(n892),
    .Z(n900)
  );
  XOR2X1 n_n321 (
    .A1(a_65_),
    .A2(b_65_),
    .Z(n904)
  );
  AND2X2 n_n322 (
    .A1(a_65_),
    .A2(b_65_),
    .Z(n903)
  );
  AOI22X1 n_n323 (
    .A1(a_65_),
    .A2(b_65_),
    .A3(n895),
    .A4(n900),
    .Z(n908)
  );
  XOR2X1 n_n324 (
    .A1(a_66_),
    .A2(b_66_),
    .Z(n912)
  );
  AND2X2 n_n325 (
    .A1(a_66_),
    .A2(b_66_),
    .Z(n911)
  );
  AOI22X1 n_n326 (
    .A1(a_66_),
    .A2(b_66_),
    .A3(n903),
    .A4(n908),
    .Z(n916)
  );
  XOR2X1 n_n327 (
    .A1(a_67_),
    .A2(b_67_),
    .Z(n920)
  );
  AND2X2 n_n328 (
    .A1(a_67_),
    .A2(b_67_),
    .Z(n919)
  );
  AOI22X1 n_n329 (
    .A1(a_67_),
    .A2(b_67_),
    .A3(n911),
    .A4(n916),
    .Z(n924)
  );
  XOR2X1 n_n330 (
    .A1(a_68_),
    .A2(b_68_),
    .Z(n928)
  );
  AND2X2 n_n331 (
    .A1(a_68_),
    .A2(b_68_),
    .Z(n927)
  );
  AOI22X1 n_n332 (
    .A1(a_68_),
    .A2(b_68_),
    .A3(n919),
    .A4(n924),
    .Z(n932)
  );
  XOR2X1 n_n333 (
    .A1(a_69_),
    .A2(b_69_),
    .Z(n936)
  );
  AND2X2 n_n334 (
    .A1(a_69_),
    .A2(b_69_),
    .Z(n935)
  );
  AOI22X1 n_n335 (
    .A1(a_69_),
    .A2(b_69_),
    .A3(n927),
    .A4(n932),
    .Z(n940)
  );
  XOR2X1 n_n336 (
    .A1(a_70_),
    .A2(b_70_),
    .Z(n944)
  );
  AND2X2 n_n337 (
    .A1(a_70_),
    .A2(b_70_),
    .Z(n943)
  );
  AOI22X1 n_n338 (
    .A1(a_70_),
    .A2(b_70_),
    .A3(n935),
    .A4(n940),
    .Z(n948)
  );
  XOR2X1 n_n339 (
    .A1(a_71_),
    .A2(b_71_),
    .Z(n952)
  );
  AND2X2 n_n340 (
    .A1(a_71_),
    .A2(b_71_),
    .Z(n951)
  );
  AOI22X1 n_n341 (
    .A1(a_71_),
    .A2(b_71_),
    .A3(n943),
    .A4(n948),
    .Z(n956)
  );
  XOR2X1 n_n342 (
    .A1(a_72_),
    .A2(b_72_),
    .Z(n960)
  );
  AND2X2 n_n343 (
    .A1(a_72_),
    .A2(b_72_),
    .Z(n959)
  );
  AOI22X1 n_n344 (
    .A1(a_72_),
    .A2(b_72_),
    .A3(n951),
    .A4(n956),
    .Z(n964)
  );
  XOR2X1 n_n345 (
    .A1(a_73_),
    .A2(b_73_),
    .Z(n968)
  );
  AND2X2 n_n346 (
    .A1(a_73_),
    .A2(b_73_),
    .Z(n967)
  );
  AOI22X1 n_n347 (
    .A1(a_73_),
    .A2(b_73_),
    .A3(n959),
    .A4(n964),
    .Z(n972)
  );
  XOR2X1 n_n348 (
    .A1(a_74_),
    .A2(b_74_),
    .Z(n976)
  );
  AND2X2 n_n349 (
    .A1(a_74_),
    .A2(b_74_),
    .Z(n975)
  );
  AOI22X1 n_n350 (
    .A1(a_74_),
    .A2(b_74_),
    .A3(n967),
    .A4(n972),
    .Z(n980)
  );
  XOR2X1 n_n351 (
    .A1(a_75_),
    .A2(b_75_),
    .Z(n984)
  );
  AND2X2 n_n352 (
    .A1(a_75_),
    .A2(b_75_),
    .Z(n983)
  );
  AOI22X1 n_n353 (
    .A1(a_75_),
    .A2(b_75_),
    .A3(n975),
    .A4(n980),
    .Z(n988)
  );
  XOR2X1 n_n354 (
    .A1(a_76_),
    .A2(b_76_),
    .Z(n992)
  );
  XOR2X1 n_n355 (
    .A1(a_77_),
    .A2(b_77_),
    .Z(n1000)
  );
  AND2X2 n_n356 (
    .A1(a_76_),
    .A2(b_76_),
    .Z(n991)
  );
  AOI22X1 n_n357 (
    .A1(a_76_),
    .A2(b_76_),
    .A3(n983),
    .A4(n988),
    .Z(n996)
  );
  AOI22X1 n_n358 (
    .A1(a_77_),
    .A2(b_77_),
    .A3(n991),
    .A4(n996),
    .Z(n1004)
  );
  XOR2X1 n_n359 (
    .A1(a_78_),
    .A2(b_78_),
    .Z(n1008)
  );
  AND2X2 n_n360 (
    .A1(a_77_),
    .A2(b_77_),
    .Z(n999)
  );
  AND2X2 n_n361 (
    .A1(a_78_),
    .A2(b_78_),
    .Z(n1007)
  );
  AOI22X1 n_n362 (
    .A1(a_78_),
    .A2(b_78_),
    .A3(n1004),
    .A4(n999),
    .Z(n1012)
  );
  XOR2X1 n_n363 (
    .A1(a_79_),
    .A2(b_79_),
    .Z(n1016)
  );
  AND2X2 n_n364 (
    .A1(a_79_),
    .A2(b_79_),
    .Z(n1015)
  );
  AOI22X1 n_n365 (
    .A1(a_79_),
    .A2(b_79_),
    .A3(n1007),
    .A4(n1012),
    .Z(n1020)
  );
  XOR2X1 n_n366 (
    .A1(a_80_),
    .A2(b_80_),
    .Z(n1024)
  );
  AND2X2 n_n367 (
    .A1(a_80_),
    .A2(b_80_),
    .Z(n1023)
  );
  AOI22X1 n_n368 (
    .A1(a_80_),
    .A2(b_80_),
    .A3(n1015),
    .A4(n1020),
    .Z(n1028)
  );
  XOR2X1 n_n369 (
    .A1(a_81_),
    .A2(b_81_),
    .Z(n1032)
  );
  AND2X2 n_n370 (
    .A1(a_81_),
    .A2(b_81_),
    .Z(n1031)
  );
  AOI22X1 n_n371 (
    .A1(a_81_),
    .A2(b_81_),
    .A3(n1023),
    .A4(n1028),
    .Z(n1036)
  );
  XOR2X1 n_n372 (
    .A1(a_82_),
    .A2(b_82_),
    .Z(n1040)
  );
  AND2X2 n_n373 (
    .A1(a_82_),
    .A2(b_82_),
    .Z(n1039)
  );
  AOI22X1 n_n374 (
    .A1(a_82_),
    .A2(b_82_),
    .A3(n1031),
    .A4(n1036),
    .Z(n1044)
  );
  XOR2X1 n_n375 (
    .A1(a_83_),
    .A2(b_83_),
    .Z(n1048)
  );
  AND2X2 n_n376 (
    .A1(a_83_),
    .A2(b_83_),
    .Z(n1047)
  );
  AOI22X1 n_n377 (
    .A1(a_83_),
    .A2(b_83_),
    .A3(n1039),
    .A4(n1044),
    .Z(n1052)
  );
  XOR2X1 n_n378 (
    .A1(a_84_),
    .A2(b_84_),
    .Z(n1056)
  );
  AND2X2 n_n379 (
    .A1(a_84_),
    .A2(b_84_),
    .Z(n1055)
  );
  AOI22X1 n_n380 (
    .A1(a_84_),
    .A2(b_84_),
    .A3(n1047),
    .A4(n1052),
    .Z(n1060)
  );
  XOR2X1 n_n381 (
    .A1(a_85_),
    .A2(b_85_),
    .Z(n1064)
  );
  AND2X2 n_n382 (
    .A1(a_85_),
    .A2(b_85_),
    .Z(n1063)
  );
  AOI22X1 n_n383 (
    .A1(a_85_),
    .A2(b_85_),
    .A3(n1055),
    .A4(n1060),
    .Z(n1068)
  );
  XOR2X1 n_n384 (
    .A1(a_86_),
    .A2(b_86_),
    .Z(n1072)
  );
  AND2X2 n_n385 (
    .A1(a_86_),
    .A2(b_86_),
    .Z(n1071)
  );
  AOI22X1 n_n386 (
    .A1(a_86_),
    .A2(b_86_),
    .A3(n1063),
    .A4(n1068),
    .Z(n1076)
  );
  XOR2X1 n_n387 (
    .A1(a_87_),
    .A2(b_87_),
    .Z(n1080)
  );
  AND2X2 n_n388 (
    .A1(a_87_),
    .A2(b_87_),
    .Z(n1079)
  );
  AOI22X1 n_n389 (
    .A1(a_87_),
    .A2(b_87_),
    .A3(n1071),
    .A4(n1076),
    .Z(n1084)
  );
  XOR2X1 n_n390 (
    .A1(a_88_),
    .A2(b_88_),
    .Z(n1088)
  );
  AND2X2 n_n391 (
    .A1(a_88_),
    .A2(b_88_),
    .Z(n1087)
  );
  AOI22X1 n_n392 (
    .A1(a_88_),
    .A2(b_88_),
    .A3(n1079),
    .A4(n1084),
    .Z(n1092)
  );
  XOR2X1 n_n393 (
    .A1(a_89_),
    .A2(b_89_),
    .Z(n1096)
  );
  AND2X2 n_n394 (
    .A1(a_89_),
    .A2(b_89_),
    .Z(n1095)
  );
  AOI22X1 n_n395 (
    .A1(a_89_),
    .A2(b_89_),
    .A3(n1087),
    .A4(n1092),
    .Z(n1100)
  );
  XOR2X1 n_n396 (
    .A1(a_90_),
    .A2(b_90_),
    .Z(n1104)
  );
  AND2X2 n_n397 (
    .A1(a_90_),
    .A2(b_90_),
    .Z(n1103)
  );
  AOI22X1 n_n398 (
    .A1(a_90_),
    .A2(b_90_),
    .A3(n1095),
    .A4(n1100),
    .Z(n1108)
  );
  XOR2X1 n_n399 (
    .A1(a_91_),
    .A2(b_91_),
    .Z(n1112)
  );
  AND2X2 n_n400 (
    .A1(a_91_),
    .A2(b_91_),
    .Z(n1111)
  );
  AOI22X1 n_n401 (
    .A1(a_91_),
    .A2(b_91_),
    .A3(n1103),
    .A4(n1108),
    .Z(n1116)
  );
  XOR2X1 n_n402 (
    .A1(a_92_),
    .A2(b_92_),
    .Z(n1120)
  );
  AND2X2 n_n403 (
    .A1(a_92_),
    .A2(b_92_),
    .Z(n1119)
  );
  AOI22X1 n_n404 (
    .A1(a_92_),
    .A2(b_92_),
    .A3(n1111),
    .A4(n1116),
    .Z(n1124)
  );
  XOR2X1 n_n405 (
    .A1(a_93_),
    .A2(b_93_),
    .Z(n1128)
  );
  AND2X2 n_n406 (
    .A1(a_93_),
    .A2(b_93_),
    .Z(n1127)
  );
  AOI22X1 n_n407 (
    .A1(a_93_),
    .A2(b_93_),
    .A3(n1119),
    .A4(n1124),
    .Z(n1132)
  );
  XOR2X1 n_n408 (
    .A1(a_94_),
    .A2(b_94_),
    .Z(n1136)
  );
  AND2X2 n_n409 (
    .A1(a_94_),
    .A2(b_94_),
    .Z(n1135)
  );
  AOI22X1 n_n410 (
    .A1(a_94_),
    .A2(b_94_),
    .A3(n1127),
    .A4(n1132),
    .Z(n1140)
  );
  XOR2X1 n_n411 (
    .A1(a_95_),
    .A2(b_95_),
    .Z(n1144)
  );
  AND2X2 n_n412 (
    .A1(a_95_),
    .A2(b_95_),
    .Z(n1143)
  );
  AOI22X1 n_n413 (
    .A1(a_95_),
    .A2(b_95_),
    .A3(n1135),
    .A4(n1140),
    .Z(n1148)
  );
  XOR2X1 n_n414 (
    .A1(a_96_),
    .A2(b_96_),
    .Z(n1152)
  );
  AND2X2 n_n415 (
    .A1(a_96_),
    .A2(b_96_),
    .Z(n1151)
  );
  AOI22X1 n_n416 (
    .A1(a_96_),
    .A2(b_96_),
    .A3(n1143),
    .A4(n1148),
    .Z(n1156)
  );
  XOR2X1 n_n417 (
    .A1(a_97_),
    .A2(b_97_),
    .Z(n1160)
  );
  AND2X2 n_n418 (
    .A1(a_97_),
    .A2(b_97_),
    .Z(n1159)
  );
  AOI22X1 n_n419 (
    .A1(a_97_),
    .A2(b_97_),
    .A3(n1151),
    .A4(n1156),
    .Z(n1164)
  );
  XOR2X1 n_n420 (
    .A1(a_98_),
    .A2(b_98_),
    .Z(n1168)
  );
  AND2X2 n_n421 (
    .A1(a_98_),
    .A2(b_98_),
    .Z(n1167)
  );
  AOI22X1 n_n422 (
    .A1(a_98_),
    .A2(b_98_),
    .A3(n1159),
    .A4(n1164),
    .Z(n1172)
  );
  XOR2X1 n_n423 (
    .A1(a_99_),
    .A2(b_99_),
    .Z(n1176)
  );
  AND2X2 n_n424 (
    .A1(a_99_),
    .A2(b_99_),
    .Z(n1175)
  );
  AOI22X1 n_n425 (
    .A1(a_99_),
    .A2(b_99_),
    .A3(n1167),
    .A4(n1172),
    .Z(n1180)
  );
  XOR2X1 n_n426 (
    .A1(a_100_),
    .A2(b_100_),
    .Z(n1184)
  );
  AND2X2 n_n427 (
    .A1(a_100_),
    .A2(b_100_),
    .Z(n1183)
  );
  AOI22X1 n_n428 (
    .A1(a_100_),
    .A2(b_100_),
    .A3(n1175),
    .A4(n1180),
    .Z(n1188)
  );
  XOR2X1 n_n429 (
    .A1(a_101_),
    .A2(b_101_),
    .Z(n1192)
  );
  AND2X2 n_n430 (
    .A1(a_101_),
    .A2(b_101_),
    .Z(n1191)
  );
  AOI22X1 n_n431 (
    .A1(a_101_),
    .A2(b_101_),
    .A3(n1183),
    .A4(n1188),
    .Z(n1196)
  );
  XOR2X1 n_n432 (
    .A1(a_102_),
    .A2(b_102_),
    .Z(n1200)
  );
  AND2X2 n_n433 (
    .A1(a_102_),
    .A2(b_102_),
    .Z(n1199)
  );
  AOI22X1 n_n434 (
    .A1(a_102_),
    .A2(b_102_),
    .A3(n1191),
    .A4(n1196),
    .Z(n1204)
  );
  XOR2X1 n_n435 (
    .A1(a_103_),
    .A2(b_103_),
    .Z(n1208)
  );
  AND2X2 n_n436 (
    .A1(a_103_),
    .A2(b_103_),
    .Z(n1207)
  );
  AOI22X1 n_n437 (
    .A1(a_103_),
    .A2(b_103_),
    .A3(n1199),
    .A4(n1204),
    .Z(n1212)
  );
  XOR2X1 n_n438 (
    .A1(a_104_),
    .A2(b_104_),
    .Z(n1216)
  );
  AND2X2 n_n439 (
    .A1(a_104_),
    .A2(b_104_),
    .Z(n1215)
  );
  AOI22X1 n_n440 (
    .A1(a_104_),
    .A2(b_104_),
    .A3(n1207),
    .A4(n1212),
    .Z(n1220)
  );
  XOR2X1 n_n441 (
    .A1(a_105_),
    .A2(b_105_),
    .Z(n1224)
  );
  AND2X2 n_n442 (
    .A1(a_105_),
    .A2(b_105_),
    .Z(n1223)
  );
  AOI22X1 n_n443 (
    .A1(a_105_),
    .A2(b_105_),
    .A3(n1215),
    .A4(n1220),
    .Z(n1228)
  );
  XOR2X1 n_n444 (
    .A1(a_106_),
    .A2(b_106_),
    .Z(n1232)
  );
  AND2X2 n_n445 (
    .A1(a_106_),
    .A2(b_106_),
    .Z(n1231)
  );
  AOI22X1 n_n446 (
    .A1(a_106_),
    .A2(b_106_),
    .A3(n1223),
    .A4(n1228),
    .Z(n1236)
  );
  XOR2X1 n_n447 (
    .A1(a_107_),
    .A2(b_107_),
    .Z(n1240)
  );
  AND2X2 n_n448 (
    .A1(a_107_),
    .A2(b_107_),
    .Z(n1239)
  );
  AOI22X1 n_n449 (
    .A1(a_107_),
    .A2(b_107_),
    .A3(n1231),
    .A4(n1236),
    .Z(n1244)
  );
  XOR2X1 n_n450 (
    .A1(a_108_),
    .A2(b_108_),
    .Z(n1248)
  );
  AND2X2 n_n451 (
    .A1(a_108_),
    .A2(b_108_),
    .Z(n1247)
  );
  AOI22X1 n_n452 (
    .A1(a_108_),
    .A2(b_108_),
    .A3(n1239),
    .A4(n1244),
    .Z(n1252)
  );
  XOR2X1 n_n453 (
    .A1(a_109_),
    .A2(b_109_),
    .Z(n1256)
  );
  AND2X2 n_n454 (
    .A1(a_109_),
    .A2(b_109_),
    .Z(n1255)
  );
  AOI22X1 n_n455 (
    .A1(a_109_),
    .A2(b_109_),
    .A3(n1247),
    .A4(n1252),
    .Z(n1260)
  );
  XOR2X1 n_n456 (
    .A1(a_110_),
    .A2(b_110_),
    .Z(n1264)
  );
  AND2X2 n_n457 (
    .A1(a_110_),
    .A2(b_110_),
    .Z(n1263)
  );
  AOI22X1 n_n458 (
    .A1(a_110_),
    .A2(b_110_),
    .A3(n1255),
    .A4(n1260),
    .Z(n1268)
  );
  XOR2X1 n_n459 (
    .A1(a_111_),
    .A2(b_111_),
    .Z(n1272)
  );
  AND2X2 n_n460 (
    .A1(a_111_),
    .A2(b_111_),
    .Z(n1271)
  );
  AOI22X1 n_n461 (
    .A1(a_111_),
    .A2(b_111_),
    .A3(n1263),
    .A4(n1268),
    .Z(n1276)
  );
  XOR2X1 n_n462 (
    .A1(a_112_),
    .A2(b_112_),
    .Z(n1280)
  );
  AND2X2 n_n463 (
    .A1(a_112_),
    .A2(b_112_),
    .Z(n1279)
  );
  AOI22X1 n_n464 (
    .A1(a_112_),
    .A2(b_112_),
    .A3(n1271),
    .A4(n1276),
    .Z(n1284)
  );
  XOR2X1 n_n465 (
    .A1(a_113_),
    .A2(b_113_),
    .Z(n1288)
  );
  AND2X2 n_n466 (
    .A1(a_113_),
    .A2(b_113_),
    .Z(n1287)
  );
  AOI22X1 n_n467 (
    .A1(a_113_),
    .A2(b_113_),
    .A3(n1279),
    .A4(n1284),
    .Z(n1292)
  );
  XOR2X1 n_n468 (
    .A1(a_114_),
    .A2(b_114_),
    .Z(n1296)
  );
  AND2X2 n_n469 (
    .A1(a_114_),
    .A2(b_114_),
    .Z(n1295)
  );
  AOI22X1 n_n470 (
    .A1(a_114_),
    .A2(b_114_),
    .A3(n1287),
    .A4(n1292),
    .Z(n1300)
  );
  XOR2X1 n_n471 (
    .A1(a_115_),
    .A2(b_115_),
    .Z(n1304)
  );
  AND2X2 n_n472 (
    .A1(a_115_),
    .A2(b_115_),
    .Z(n1303)
  );
  AOI22X1 n_n473 (
    .A1(a_115_),
    .A2(b_115_),
    .A3(n1295),
    .A4(n1300),
    .Z(n1308)
  );
  XOR2X1 n_n474 (
    .A1(a_116_),
    .A2(b_116_),
    .Z(n1312)
  );
  AND2X2 n_n475 (
    .A1(a_116_),
    .A2(b_116_),
    .Z(n1311)
  );
  AOI22X1 n_n476 (
    .A1(a_116_),
    .A2(b_116_),
    .A3(n1303),
    .A4(n1308),
    .Z(n1316)
  );
  XOR2X1 n_n477 (
    .A1(a_117_),
    .A2(b_117_),
    .Z(n1320)
  );
  AND2X2 n_n478 (
    .A1(a_117_),
    .A2(b_117_),
    .Z(n1319)
  );
  AOI22X1 n_n479 (
    .A1(a_117_),
    .A2(b_117_),
    .A3(n1311),
    .A4(n1316),
    .Z(n1324)
  );
  XOR2X1 n_n480 (
    .A1(a_118_),
    .A2(b_118_),
    .Z(n1328)
  );
  AND2X2 n_n481 (
    .A1(a_118_),
    .A2(b_118_),
    .Z(n1327)
  );
  AOI22X1 n_n482 (
    .A1(a_118_),
    .A2(b_118_),
    .A3(n1319),
    .A4(n1324),
    .Z(n1332)
  );
  XOR2X1 n_n483 (
    .A1(a_119_),
    .A2(b_119_),
    .Z(n1336)
  );
  AND2X2 n_n484 (
    .A1(a_119_),
    .A2(b_119_),
    .Z(n1335)
  );
  AOI22X1 n_n485 (
    .A1(a_119_),
    .A2(b_119_),
    .A3(n1327),
    .A4(n1332),
    .Z(n1340)
  );
  XOR2X1 n_n486 (
    .A1(a_120_),
    .A2(b_120_),
    .Z(n1344)
  );
  AND2X2 n_n487 (
    .A1(a_120_),
    .A2(b_120_),
    .Z(n1343)
  );
  AOI22X1 n_n488 (
    .A1(a_120_),
    .A2(b_120_),
    .A3(n1335),
    .A4(n1340),
    .Z(n1348)
  );
  XOR2X1 n_n489 (
    .A1(a_121_),
    .A2(b_121_),
    .Z(n1352)
  );
  AND2X2 n_n490 (
    .A1(a_121_),
    .A2(b_121_),
    .Z(n1351)
  );
  AOI22X1 n_n491 (
    .A1(a_121_),
    .A2(b_121_),
    .A3(n1343),
    .A4(n1348),
    .Z(n1356)
  );
  XOR2X1 n_n492 (
    .A1(a_122_),
    .A2(b_122_),
    .Z(n1360)
  );
  AND2X2 n_n493 (
    .A1(a_122_),
    .A2(b_122_),
    .Z(n1359)
  );
  AOI22X1 n_n494 (
    .A1(a_122_),
    .A2(b_122_),
    .A3(n1351),
    .A4(n1356),
    .Z(n1364)
  );
  XOR2X1 n_n495 (
    .A1(a_123_),
    .A2(b_123_),
    .Z(n1368)
  );
  AND2X2 n_n496 (
    .A1(a_123_),
    .A2(b_123_),
    .Z(n1367)
  );
  AOI22X1 n_n497 (
    .A1(a_123_),
    .A2(b_123_),
    .A3(n1359),
    .A4(n1364),
    .Z(n1372)
  );
  XOR2X1 n_n498 (
    .A1(a_124_),
    .A2(b_124_),
    .Z(n1376)
  );
  AND2X2 n_n499 (
    .A1(a_124_),
    .A2(b_124_),
    .Z(n1375)
  );
  AOI22X1 n_n500 (
    .A1(a_124_),
    .A2(b_124_),
    .A3(n1367),
    .A4(n1372),
    .Z(n1380)
  );
  XOR2X1 n_n501 (
    .A1(a_125_),
    .A2(b_125_),
    .Z(n1384)
  );
  AND2X2 n_n502 (
    .A1(a_125_),
    .A2(b_125_),
    .Z(n1383)
  );
  AOI22X1 n_n503 (
    .A1(a_125_),
    .A2(b_125_),
    .A3(n1375),
    .A4(n1380),
    .Z(n1388)
  );
  XOR2X1 n_n504 (
    .A1(a_126_),
    .A2(b_126_),
    .Z(n1392)
  );
  AND2X2 n_n505 (
    .A1(a_126_),
    .A2(b_126_),
    .Z(n1391)
  );
  AOI22X1 n_n506 (
    .A1(a_126_),
    .A2(b_126_),
    .A3(n1383),
    .A4(n1388),
    .Z(n1396)
  );
  XOR2X1 n_n507 (
    .A1(a_127_),
    .A2(b_127_),
    .Z(n1400)
  );
  AOI21X1 n_n508 (
    .A1(n1389),
    .A2(n1390),
    .A3(n1391),
    .Z(n1397)
  );
  AND2X2 n_n509 (
    .A1(a_127_),
    .A2(b_127_),
    .Z(n1398)
  );
  AND2X2 n_n510 (
    .A1(a_127_),
    .A2(b_127_),
    .Z(n1399)
  );
  AND2X2 n_n511 (
    .A1(a_1_),
    .A2(b_1_),
    .Z(n390)
  );
  AOI21X1 n_n512 (
    .A1(n1381),
    .A2(n1382),
    .A3(n1383),
    .Z(n1389)
  );
  AND2X2 n_n513 (
    .A1(a_126_),
    .A2(b_126_),
    .Z(n1390)
  );
  AOI21X1 n_n514 (
    .A1(n1373),
    .A2(n1374),
    .A3(n1375),
    .Z(n1381)
  );
  AND2X2 n_n515 (
    .A1(a_125_),
    .A2(b_125_),
    .Z(n1382)
  );
  AOI21X1 n_n516 (
    .A1(n1365),
    .A2(n1366),
    .A3(n1367),
    .Z(n1373)
  );
  AND2X2 n_n517 (
    .A1(a_124_),
    .A2(b_124_),
    .Z(n1374)
  );
  AOI21X1 n_n518 (
    .A1(n1357),
    .A2(n1358),
    .A3(n1359),
    .Z(n1365)
  );
  AND2X2 n_n519 (
    .A1(a_123_),
    .A2(b_123_),
    .Z(n1366)
  );
  AOI21X1 n_n520 (
    .A1(n1349),
    .A2(n1350),
    .A3(n1351),
    .Z(n1357)
  );
  AND2X2 n_n521 (
    .A1(a_122_),
    .A2(b_122_),
    .Z(n1358)
  );
  AOI21X1 n_n522 (
    .A1(n1341),
    .A2(n1342),
    .A3(n1343),
    .Z(n1349)
  );
  AND2X2 n_n523 (
    .A1(a_121_),
    .A2(b_121_),
    .Z(n1350)
  );
  AOI21X1 n_n524 (
    .A1(n1333),
    .A2(n1334),
    .A3(n1335),
    .Z(n1341)
  );
  AND2X2 n_n525 (
    .A1(a_120_),
    .A2(b_120_),
    .Z(n1342)
  );
  AOI21X1 n_n526 (
    .A1(n1325),
    .A2(n1326),
    .A3(n1327),
    .Z(n1333)
  );
  AND2X2 n_n527 (
    .A1(a_119_),
    .A2(b_119_),
    .Z(n1334)
  );
  AOI21X1 n_n528 (
    .A1(n1317),
    .A2(n1318),
    .A3(n1319),
    .Z(n1325)
  );
  AND2X2 n_n529 (
    .A1(a_118_),
    .A2(b_118_),
    .Z(n1326)
  );
  AOI21X1 n_n530 (
    .A1(n1309),
    .A2(n1310),
    .A3(n1311),
    .Z(n1317)
  );
  AND2X2 n_n531 (
    .A1(a_117_),
    .A2(b_117_),
    .Z(n1318)
  );
  AOI21X1 n_n532 (
    .A1(n1301),
    .A2(n1302),
    .A3(n1303),
    .Z(n1309)
  );
  AND2X2 n_n533 (
    .A1(a_116_),
    .A2(b_116_),
    .Z(n1310)
  );
  AOI21X1 n_n534 (
    .A1(n1293),
    .A2(n1294),
    .A3(n1295),
    .Z(n1301)
  );
  AND2X2 n_n535 (
    .A1(a_115_),
    .A2(b_115_),
    .Z(n1302)
  );
  AOI21X1 n_n536 (
    .A1(n1285),
    .A2(n1286),
    .A3(n1287),
    .Z(n1293)
  );
  AND2X2 n_n537 (
    .A1(a_114_),
    .A2(b_114_),
    .Z(n1294)
  );
  AOI21X1 n_n538 (
    .A1(n1277),
    .A2(n1278),
    .A3(n1279),
    .Z(n1285)
  );
  AND2X2 n_n539 (
    .A1(a_113_),
    .A2(b_113_),
    .Z(n1286)
  );
  AOI21X1 n_n540 (
    .A1(n1269),
    .A2(n1270),
    .A3(n1271),
    .Z(n1277)
  );
  AND2X2 n_n541 (
    .A1(a_112_),
    .A2(b_112_),
    .Z(n1278)
  );
  AOI21X1 n_n542 (
    .A1(n1261),
    .A2(n1262),
    .A3(n1263),
    .Z(n1269)
  );
  AND2X2 n_n543 (
    .A1(a_111_),
    .A2(b_111_),
    .Z(n1270)
  );
  AOI21X1 n_n544 (
    .A1(n1253),
    .A2(n1254),
    .A3(n1255),
    .Z(n1261)
  );
  AND2X2 n_n545 (
    .A1(a_110_),
    .A2(b_110_),
    .Z(n1262)
  );
  AOI21X1 n_n546 (
    .A1(n1245),
    .A2(n1246),
    .A3(n1247),
    .Z(n1253)
  );
  AND2X2 n_n547 (
    .A1(a_109_),
    .A2(b_109_),
    .Z(n1254)
  );
  AOI21X1 n_n548 (
    .A1(n1237),
    .A2(n1238),
    .A3(n1239),
    .Z(n1245)
  );
  AND2X2 n_n549 (
    .A1(a_108_),
    .A2(b_108_),
    .Z(n1246)
  );
  AOI21X1 n_n550 (
    .A1(n1229),
    .A2(n1230),
    .A3(n1231),
    .Z(n1237)
  );
  AND2X2 n_n551 (
    .A1(a_107_),
    .A2(b_107_),
    .Z(n1238)
  );
  AOI21X1 n_n552 (
    .A1(n1221),
    .A2(n1222),
    .A3(n1223),
    .Z(n1229)
  );
  AND2X2 n_n553 (
    .A1(a_106_),
    .A2(b_106_),
    .Z(n1230)
  );
  AOI21X1 n_n554 (
    .A1(n1213),
    .A2(n1214),
    .A3(n1215),
    .Z(n1221)
  );
  AND2X2 n_n555 (
    .A1(a_105_),
    .A2(b_105_),
    .Z(n1222)
  );
  AOI21X1 n_n556 (
    .A1(n1205),
    .A2(n1206),
    .A3(n1207),
    .Z(n1213)
  );
  AND2X2 n_n557 (
    .A1(a_104_),
    .A2(b_104_),
    .Z(n1214)
  );
  AOI21X1 n_n558 (
    .A1(n1197),
    .A2(n1198),
    .A3(n1199),
    .Z(n1205)
  );
  AND2X2 n_n559 (
    .A1(a_103_),
    .A2(b_103_),
    .Z(n1206)
  );
  AOI21X1 n_n560 (
    .A1(n1189),
    .A2(n1190),
    .A3(n1191),
    .Z(n1197)
  );
  AND2X2 n_n561 (
    .A1(a_102_),
    .A2(b_102_),
    .Z(n1198)
  );
  AOI21X1 n_n562 (
    .A1(n1181),
    .A2(n1182),
    .A3(n1183),
    .Z(n1189)
  );
  AND2X2 n_n563 (
    .A1(a_101_),
    .A2(b_101_),
    .Z(n1190)
  );
  AOI21X1 n_n564 (
    .A1(n1173),
    .A2(n1174),
    .A3(n1175),
    .Z(n1181)
  );
  AND2X2 n_n565 (
    .A1(a_100_),
    .A2(b_100_),
    .Z(n1182)
  );
  AOI21X1 n_n566 (
    .A1(n1165),
    .A2(n1166),
    .A3(n1167),
    .Z(n1173)
  );
  AND2X2 n_n567 (
    .A1(a_99_),
    .A2(b_99_),
    .Z(n1174)
  );
  AOI21X1 n_n568 (
    .A1(n1157),
    .A2(n1158),
    .A3(n1159),
    .Z(n1165)
  );
  AND2X2 n_n569 (
    .A1(a_98_),
    .A2(b_98_),
    .Z(n1166)
  );
  AOI21X1 n_n570 (
    .A1(n1149),
    .A2(n1150),
    .A3(n1151),
    .Z(n1157)
  );
  AND2X2 n_n571 (
    .A1(a_97_),
    .A2(b_97_),
    .Z(n1158)
  );
  AOI21X1 n_n572 (
    .A1(n1141),
    .A2(n1142),
    .A3(n1143),
    .Z(n1149)
  );
  AND2X2 n_n573 (
    .A1(a_96_),
    .A2(b_96_),
    .Z(n1150)
  );
  AOI21X1 n_n574 (
    .A1(n1133),
    .A2(n1134),
    .A3(n1135),
    .Z(n1141)
  );
  AND2X2 n_n575 (
    .A1(a_95_),
    .A2(b_95_),
    .Z(n1142)
  );
  AOI21X1 n_n576 (
    .A1(n1125),
    .A2(n1126),
    .A3(n1127),
    .Z(n1133)
  );
  AND2X2 n_n577 (
    .A1(a_94_),
    .A2(b_94_),
    .Z(n1134)
  );
  AOI21X1 n_n578 (
    .A1(n1117),
    .A2(n1118),
    .A3(n1119),
    .Z(n1125)
  );
  AND2X2 n_n579 (
    .A1(a_93_),
    .A2(b_93_),
    .Z(n1126)
  );
  AOI21X1 n_n580 (
    .A1(n1109),
    .A2(n1110),
    .A3(n1111),
    .Z(n1117)
  );
  AND2X2 n_n581 (
    .A1(a_92_),
    .A2(b_92_),
    .Z(n1118)
  );
  AOI21X1 n_n582 (
    .A1(n1101),
    .A2(n1102),
    .A3(n1103),
    .Z(n1109)
  );
  AND2X2 n_n583 (
    .A1(a_91_),
    .A2(b_91_),
    .Z(n1110)
  );
  AOI21X1 n_n584 (
    .A1(n1093),
    .A2(n1094),
    .A3(n1095),
    .Z(n1101)
  );
  AND2X2 n_n585 (
    .A1(a_90_),
    .A2(b_90_),
    .Z(n1102)
  );
  AOI21X1 n_n586 (
    .A1(n1085),
    .A2(n1086),
    .A3(n1087),
    .Z(n1093)
  );
  AND2X2 n_n587 (
    .A1(a_89_),
    .A2(b_89_),
    .Z(n1094)
  );
  AOI21X1 n_n588 (
    .A1(n1077),
    .A2(n1078),
    .A3(n1079),
    .Z(n1085)
  );
  AND2X2 n_n589 (
    .A1(a_88_),
    .A2(b_88_),
    .Z(n1086)
  );
  AOI21X1 n_n590 (
    .A1(n1069),
    .A2(n1070),
    .A3(n1071),
    .Z(n1077)
  );
  AND2X2 n_n591 (
    .A1(a_87_),
    .A2(b_87_),
    .Z(n1078)
  );
  AOI21X1 n_n592 (
    .A1(n1061),
    .A2(n1062),
    .A3(n1063),
    .Z(n1069)
  );
  AND2X2 n_n593 (
    .A1(a_86_),
    .A2(b_86_),
    .Z(n1070)
  );
  AOI21X1 n_n594 (
    .A1(n1053),
    .A2(n1054),
    .A3(n1055),
    .Z(n1061)
  );
  AND2X2 n_n595 (
    .A1(a_85_),
    .A2(b_85_),
    .Z(n1062)
  );
  AOI21X1 n_n596 (
    .A1(n1045),
    .A2(n1046),
    .A3(n1047),
    .Z(n1053)
  );
  AND2X2 n_n597 (
    .A1(a_84_),
    .A2(b_84_),
    .Z(n1054)
  );
  AOI21X1 n_n598 (
    .A1(n1037),
    .A2(n1038),
    .A3(n1039),
    .Z(n1045)
  );
  AND2X2 n_n599 (
    .A1(a_83_),
    .A2(b_83_),
    .Z(n1046)
  );
  AOI21X1 n_n600 (
    .A1(n1029),
    .A2(n1030),
    .A3(n1031),
    .Z(n1037)
  );
  AND2X2 n_n601 (
    .A1(a_82_),
    .A2(b_82_),
    .Z(n1038)
  );
  AOI21X1 n_n602 (
    .A1(n1021),
    .A2(n1022),
    .A3(n1023),
    .Z(n1029)
  );
  AND2X2 n_n603 (
    .A1(a_81_),
    .A2(b_81_),
    .Z(n1030)
  );
  AOI21X1 n_n604 (
    .A1(n1013),
    .A2(n1014),
    .A3(n1015),
    .Z(n1021)
  );
  AND2X2 n_n605 (
    .A1(a_80_),
    .A2(b_80_),
    .Z(n1022)
  );
  AOI21X1 n_n606 (
    .A1(n1005),
    .A2(n1006),
    .A3(n1007),
    .Z(n1013)
  );
  AND2X2 n_n607 (
    .A1(a_79_),
    .A2(b_79_),
    .Z(n1014)
  );
  AOI21X1 n_n608 (
    .A1(n997),
    .A2(n998),
    .A3(n999),
    .Z(n1005)
  );
  AND2X2 n_n609 (
    .A1(a_78_),
    .A2(b_78_),
    .Z(n1006)
  );
  AOI21X1 n_n610 (
    .A1(n989),
    .A2(n990),
    .A3(n991),
    .Z(n997)
  );
  AND2X2 n_n611 (
    .A1(a_77_),
    .A2(b_77_),
    .Z(n998)
  );
  AOI21X1 n_n612 (
    .A1(n981),
    .A2(n982),
    .A3(n983),
    .Z(n989)
  );
  AND2X2 n_n613 (
    .A1(a_76_),
    .A2(b_76_),
    .Z(n990)
  );
  AOI21X1 n_n614 (
    .A1(n973),
    .A2(n974),
    .A3(n975),
    .Z(n981)
  );
  AND2X2 n_n615 (
    .A1(a_75_),
    .A2(b_75_),
    .Z(n982)
  );
  AOI21X1 n_n616 (
    .A1(n965),
    .A2(n966),
    .A3(n967),
    .Z(n973)
  );
  AND2X2 n_n617 (
    .A1(a_74_),
    .A2(b_74_),
    .Z(n974)
  );
  AOI21X1 n_n618 (
    .A1(n957),
    .A2(n958),
    .A3(n959),
    .Z(n965)
  );
  AND2X2 n_n619 (
    .A1(a_73_),
    .A2(b_73_),
    .Z(n966)
  );
  AOI21X1 n_n620 (
    .A1(n949),
    .A2(n950),
    .A3(n951),
    .Z(n957)
  );
  AND2X2 n_n621 (
    .A1(a_72_),
    .A2(b_72_),
    .Z(n958)
  );
  AOI21X1 n_n622 (
    .A1(n941),
    .A2(n942),
    .A3(n943),
    .Z(n949)
  );
  AND2X2 n_n623 (
    .A1(a_71_),
    .A2(b_71_),
    .Z(n950)
  );
  AOI21X1 n_n624 (
    .A1(n933),
    .A2(n934),
    .A3(n935),
    .Z(n941)
  );
  AND2X2 n_n625 (
    .A1(a_70_),
    .A2(b_70_),
    .Z(n942)
  );
  AOI21X1 n_n626 (
    .A1(n925),
    .A2(n926),
    .A3(n927),
    .Z(n933)
  );
  AND2X2 n_n627 (
    .A1(a_69_),
    .A2(b_69_),
    .Z(n934)
  );
  AOI21X1 n_n628 (
    .A1(n917),
    .A2(n918),
    .A3(n919),
    .Z(n925)
  );
  AND2X2 n_n629 (
    .A1(a_68_),
    .A2(b_68_),
    .Z(n926)
  );
  AOI21X1 n_n630 (
    .A1(n909),
    .A2(n910),
    .A3(n911),
    .Z(n917)
  );
  AND2X2 n_n631 (
    .A1(a_67_),
    .A2(b_67_),
    .Z(n918)
  );
  AOI21X1 n_n632 (
    .A1(n901),
    .A2(n902),
    .A3(n903),
    .Z(n909)
  );
  AND2X2 n_n633 (
    .A1(a_66_),
    .A2(b_66_),
    .Z(n910)
  );
  AOI21X1 n_n634 (
    .A1(n893),
    .A2(n894),
    .A3(n895),
    .Z(n901)
  );
  AND2X2 n_n635 (
    .A1(a_65_),
    .A2(b_65_),
    .Z(n902)
  );
  AOI21X1 n_n636 (
    .A1(n885),
    .A2(n886),
    .A3(n887),
    .Z(n893)
  );
  AND2X2 n_n637 (
    .A1(a_64_),
    .A2(b_64_),
    .Z(n894)
  );
  AOI21X1 n_n638 (
    .A1(n877),
    .A2(n878),
    .A3(n879),
    .Z(n885)
  );
  AND2X2 n_n639 (
    .A1(a_63_),
    .A2(b_63_),
    .Z(n886)
  );
  AOI21X1 n_n640 (
    .A1(n869),
    .A2(n870),
    .A3(n871),
    .Z(n877)
  );
  AND2X2 n_n641 (
    .A1(a_62_),
    .A2(b_62_),
    .Z(n878)
  );
  AOI21X1 n_n642 (
    .A1(n861),
    .A2(n862),
    .A3(n863),
    .Z(n869)
  );
  AND2X2 n_n643 (
    .A1(a_61_),
    .A2(b_61_),
    .Z(n870)
  );
  AOI21X1 n_n644 (
    .A1(n853),
    .A2(n854),
    .A3(n855),
    .Z(n861)
  );
  AND2X2 n_n645 (
    .A1(a_60_),
    .A2(b_60_),
    .Z(n862)
  );
  AOI21X1 n_n646 (
    .A1(n845),
    .A2(n846),
    .A3(n847),
    .Z(n853)
  );
  AND2X2 n_n647 (
    .A1(a_59_),
    .A2(b_59_),
    .Z(n854)
  );
  AOI21X1 n_n648 (
    .A1(n837),
    .A2(n838),
    .A3(n839),
    .Z(n845)
  );
  AND2X2 n_n649 (
    .A1(a_58_),
    .A2(b_58_),
    .Z(n846)
  );
  AOI21X1 n_n650 (
    .A1(n829),
    .A2(n830),
    .A3(n831),
    .Z(n837)
  );
  AND2X2 n_n651 (
    .A1(a_57_),
    .A2(b_57_),
    .Z(n838)
  );
  AOI21X1 n_n652 (
    .A1(n821),
    .A2(n822),
    .A3(n823),
    .Z(n829)
  );
  AND2X2 n_n653 (
    .A1(a_56_),
    .A2(b_56_),
    .Z(n830)
  );
  AOI21X1 n_n654 (
    .A1(n813),
    .A2(n814),
    .A3(n815),
    .Z(n821)
  );
  AND2X2 n_n655 (
    .A1(a_55_),
    .A2(b_55_),
    .Z(n822)
  );
  AOI21X1 n_n656 (
    .A1(n805),
    .A2(n806),
    .A3(n807),
    .Z(n813)
  );
  AND2X2 n_n657 (
    .A1(a_54_),
    .A2(b_54_),
    .Z(n814)
  );
  AOI21X1 n_n658 (
    .A1(n797),
    .A2(n798),
    .A3(n799),
    .Z(n805)
  );
  AND2X2 n_n659 (
    .A1(a_53_),
    .A2(b_53_),
    .Z(n806)
  );
  AOI21X1 n_n660 (
    .A1(n789),
    .A2(n790),
    .A3(n791),
    .Z(n797)
  );
  AND2X2 n_n661 (
    .A1(a_52_),
    .A2(b_52_),
    .Z(n798)
  );
  AOI21X1 n_n662 (
    .A1(n781),
    .A2(n782),
    .A3(n783),
    .Z(n789)
  );
  AND2X2 n_n663 (
    .A1(a_51_),
    .A2(b_51_),
    .Z(n790)
  );
  AOI21X1 n_n664 (
    .A1(n773),
    .A2(n774),
    .A3(n775),
    .Z(n781)
  );
  AND2X2 n_n665 (
    .A1(a_50_),
    .A2(b_50_),
    .Z(n782)
  );
  AOI21X1 n_n666 (
    .A1(n765),
    .A2(n766),
    .A3(n767),
    .Z(n773)
  );
  AND2X2 n_n667 (
    .A1(a_49_),
    .A2(b_49_),
    .Z(n774)
  );
  AOI21X1 n_n668 (
    .A1(n757),
    .A2(n758),
    .A3(n759),
    .Z(n765)
  );
  AND2X2 n_n669 (
    .A1(a_48_),
    .A2(b_48_),
    .Z(n766)
  );
  AOI21X1 n_n670 (
    .A1(n749),
    .A2(n750),
    .A3(n751),
    .Z(n757)
  );
  AND2X2 n_n671 (
    .A1(a_47_),
    .A2(b_47_),
    .Z(n758)
  );
  AOI21X1 n_n672 (
    .A1(n741),
    .A2(n742),
    .A3(n743),
    .Z(n749)
  );
  AND2X2 n_n673 (
    .A1(a_46_),
    .A2(b_46_),
    .Z(n750)
  );
  AOI21X1 n_n674 (
    .A1(n733),
    .A2(n734),
    .A3(n735),
    .Z(n741)
  );
  AND2X2 n_n675 (
    .A1(a_45_),
    .A2(b_45_),
    .Z(n742)
  );
  AOI21X1 n_n676 (
    .A1(n725),
    .A2(n726),
    .A3(n727),
    .Z(n733)
  );
  AND2X2 n_n677 (
    .A1(a_44_),
    .A2(b_44_),
    .Z(n734)
  );
  AOI21X1 n_n678 (
    .A1(n717),
    .A2(n718),
    .A3(n719),
    .Z(n725)
  );
  AND2X2 n_n679 (
    .A1(a_43_),
    .A2(b_43_),
    .Z(n726)
  );
  AOI21X1 n_n680 (
    .A1(n709),
    .A2(n710),
    .A3(n711),
    .Z(n717)
  );
  AND2X2 n_n681 (
    .A1(a_42_),
    .A2(b_42_),
    .Z(n718)
  );
  AOI21X1 n_n682 (
    .A1(n701),
    .A2(n702),
    .A3(n703),
    .Z(n709)
  );
  AND2X2 n_n683 (
    .A1(a_41_),
    .A2(b_41_),
    .Z(n710)
  );
  AOI21X1 n_n684 (
    .A1(n693),
    .A2(n694),
    .A3(n695),
    .Z(n701)
  );
  AND2X2 n_n685 (
    .A1(a_40_),
    .A2(b_40_),
    .Z(n702)
  );
  AOI21X1 n_n686 (
    .A1(n685),
    .A2(n686),
    .A3(n687),
    .Z(n693)
  );
  AND2X2 n_n687 (
    .A1(a_39_),
    .A2(b_39_),
    .Z(n694)
  );
  AOI21X1 n_n688 (
    .A1(n677),
    .A2(n678),
    .A3(n679),
    .Z(n685)
  );
  AND2X2 n_n689 (
    .A1(a_38_),
    .A2(b_38_),
    .Z(n686)
  );
  AOI21X1 n_n690 (
    .A1(n669),
    .A2(n670),
    .A3(n671),
    .Z(n677)
  );
  AND2X2 n_n691 (
    .A1(a_37_),
    .A2(b_37_),
    .Z(n678)
  );
  AOI21X1 n_n692 (
    .A1(n661),
    .A2(n662),
    .A3(n663),
    .Z(n669)
  );
  AND2X2 n_n693 (
    .A1(a_36_),
    .A2(b_36_),
    .Z(n670)
  );
  AOI21X1 n_n694 (
    .A1(n653),
    .A2(n654),
    .A3(n655),
    .Z(n661)
  );
  AND2X2 n_n695 (
    .A1(a_35_),
    .A2(b_35_),
    .Z(n662)
  );
  AOI21X1 n_n696 (
    .A1(n645),
    .A2(n646),
    .A3(n647),
    .Z(n653)
  );
  AND2X2 n_n697 (
    .A1(a_34_),
    .A2(b_34_),
    .Z(n654)
  );
  AOI21X1 n_n698 (
    .A1(n637),
    .A2(n638),
    .A3(n639),
    .Z(n645)
  );
  AND2X2 n_n699 (
    .A1(a_33_),
    .A2(b_33_),
    .Z(n646)
  );
  AOI21X1 n_n700 (
    .A1(n629),
    .A2(n630),
    .A3(n631),
    .Z(n637)
  );
  AND2X2 n_n701 (
    .A1(a_32_),
    .A2(b_32_),
    .Z(n638)
  );
  AOI21X1 n_n702 (
    .A1(n621),
    .A2(n622),
    .A3(n623),
    .Z(n629)
  );
  AND2X2 n_n703 (
    .A1(a_31_),
    .A2(b_31_),
    .Z(n630)
  );
  AOI21X1 n_n704 (
    .A1(n613),
    .A2(n614),
    .A3(n615),
    .Z(n621)
  );
  AND2X2 n_n705 (
    .A1(a_30_),
    .A2(b_30_),
    .Z(n622)
  );
  AOI21X1 n_n706 (
    .A1(n605),
    .A2(n606),
    .A3(n607),
    .Z(n613)
  );
  AND2X2 n_n707 (
    .A1(a_29_),
    .A2(b_29_),
    .Z(n614)
  );
  AOI21X1 n_n708 (
    .A1(n597),
    .A2(n598),
    .A3(n599),
    .Z(n605)
  );
  AND2X2 n_n709 (
    .A1(a_28_),
    .A2(b_28_),
    .Z(n606)
  );
  AOI21X1 n_n710 (
    .A1(n589),
    .A2(n590),
    .A3(n591),
    .Z(n597)
  );
  AND2X2 n_n711 (
    .A1(a_27_),
    .A2(b_27_),
    .Z(n598)
  );
  AOI21X1 n_n712 (
    .A1(n581),
    .A2(n582),
    .A3(n583),
    .Z(n589)
  );
  AND2X2 n_n713 (
    .A1(a_26_),
    .A2(b_26_),
    .Z(n590)
  );
  AOI21X1 n_n714 (
    .A1(n573),
    .A2(n574),
    .A3(n575),
    .Z(n581)
  );
  AND2X2 n_n715 (
    .A1(a_25_),
    .A2(b_25_),
    .Z(n582)
  );
  AOI21X1 n_n716 (
    .A1(n565),
    .A2(n566),
    .A3(n567),
    .Z(n573)
  );
  AND2X2 n_n717 (
    .A1(a_24_),
    .A2(b_24_),
    .Z(n574)
  );
  AOI21X1 n_n718 (
    .A1(n557),
    .A2(n558),
    .A3(n559),
    .Z(n565)
  );
  AND2X2 n_n719 (
    .A1(a_23_),
    .A2(b_23_),
    .Z(n566)
  );
  AOI21X1 n_n720 (
    .A1(n549),
    .A2(n550),
    .A3(n551),
    .Z(n557)
  );
  AND2X2 n_n721 (
    .A1(a_22_),
    .A2(b_22_),
    .Z(n558)
  );
  AOI21X1 n_n722 (
    .A1(n541),
    .A2(n542),
    .A3(n543),
    .Z(n549)
  );
  AND2X2 n_n723 (
    .A1(a_21_),
    .A2(b_21_),
    .Z(n550)
  );
  AOI21X1 n_n724 (
    .A1(n533),
    .A2(n534),
    .A3(n535),
    .Z(n541)
  );
  AND2X2 n_n725 (
    .A1(a_20_),
    .A2(b_20_),
    .Z(n542)
  );
  AOI21X1 n_n726 (
    .A1(n525),
    .A2(n526),
    .A3(n527),
    .Z(n533)
  );
  AND2X2 n_n727 (
    .A1(a_19_),
    .A2(b_19_),
    .Z(n534)
  );
  AOI21X1 n_n728 (
    .A1(n517),
    .A2(n518),
    .A3(n519),
    .Z(n525)
  );
  AND2X2 n_n729 (
    .A1(a_18_),
    .A2(b_18_),
    .Z(n526)
  );
  AOI21X1 n_n730 (
    .A1(n509),
    .A2(n510),
    .A3(n511),
    .Z(n517)
  );
  AND2X2 n_n731 (
    .A1(a_17_),
    .A2(b_17_),
    .Z(n518)
  );
  AOI21X1 n_n732 (
    .A1(n501),
    .A2(n502),
    .A3(n503),
    .Z(n509)
  );
  AND2X2 n_n733 (
    .A1(a_16_),
    .A2(b_16_),
    .Z(n510)
  );
  AOI21X1 n_n734 (
    .A1(n493),
    .A2(n494),
    .A3(n495),
    .Z(n501)
  );
  AND2X2 n_n735 (
    .A1(a_15_),
    .A2(b_15_),
    .Z(n502)
  );
  AOI21X1 n_n736 (
    .A1(n485),
    .A2(n486),
    .A3(n487),
    .Z(n493)
  );
  AND2X2 n_n737 (
    .A1(a_14_),
    .A2(b_14_),
    .Z(n494)
  );
  AOI21X1 n_n738 (
    .A1(n477),
    .A2(n478),
    .A3(n479),
    .Z(n485)
  );
  AND2X2 n_n739 (
    .A1(a_13_),
    .A2(b_13_),
    .Z(n486)
  );
  AOI21X1 n_n740 (
    .A1(n469),
    .A2(n470),
    .A3(n471),
    .Z(n477)
  );
  AND2X2 n_n741 (
    .A1(a_12_),
    .A2(b_12_),
    .Z(n478)
  );
  AOI21X1 n_n742 (
    .A1(n461),
    .A2(n462),
    .A3(n463),
    .Z(n469)
  );
  AND2X2 n_n743 (
    .A1(a_11_),
    .A2(b_11_),
    .Z(n470)
  );
  AOI21X1 n_n744 (
    .A1(n453),
    .A2(n454),
    .A3(n455),
    .Z(n461)
  );
  AND2X2 n_n745 (
    .A1(a_10_),
    .A2(b_10_),
    .Z(n462)
  );
  AOI21X1 n_n746 (
    .A1(n445),
    .A2(n446),
    .A3(n447),
    .Z(n453)
  );
  AND2X2 n_n747 (
    .A1(a_9_),
    .A2(b_9_),
    .Z(n454)
  );
  AOI21X1 n_n748 (
    .A1(n437),
    .A2(n438),
    .A3(n439),
    .Z(n445)
  );
  AND2X2 n_n749 (
    .A1(a_8_),
    .A2(b_8_),
    .Z(n446)
  );
  AOI21X1 n_n750 (
    .A1(n429),
    .A2(n430),
    .A3(n431),
    .Z(n437)
  );
  AND2X2 n_n751 (
    .A1(a_7_),
    .A2(b_7_),
    .Z(n438)
  );
  AOI21X1 n_n752 (
    .A1(n421),
    .A2(n422),
    .A3(n423),
    .Z(n429)
  );
  AND2X2 n_n753 (
    .A1(a_6_),
    .A2(b_6_),
    .Z(n430)
  );
  AOI21X1 n_n754 (
    .A1(n413),
    .A2(n414),
    .A3(n415),
    .Z(n421)
  );
  AND2X2 n_n755 (
    .A1(a_5_),
    .A2(b_5_),
    .Z(n422)
  );
  AOI21X1 n_n756 (
    .A1(n405),
    .A2(n406),
    .A3(n407),
    .Z(n413)
  );
  AND2X2 n_n757 (
    .A1(a_4_),
    .A2(b_4_),
    .Z(n414)
  );
  AOI21X1 n_n758 (
    .A1(n397),
    .A2(n398),
    .A3(n399),
    .Z(n405)
  );
  AND2X2 n_n759 (
    .A1(a_3_),
    .A2(b_3_),
    .Z(n406)
  );
  AOI21X1 n_n760 (
    .A1(n389),
    .A2(n390),
    .A3(n391),
    .Z(n397)
  );
  AND2X2 n_n761 (
    .A1(a_2_),
    .A2(b_2_),
    .Z(n398)
  );
  AND2X2 n_n762 (
    .A1(a_0_),
    .A2(b_0_),
    .Z(n389)
  );
endmodule
