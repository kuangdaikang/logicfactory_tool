// Benchmark "testing" written by ABC on Fri Feb 25 15:13:05 2022

module 25_25 ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A10  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A10;
  wire new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_,
    new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_,
    new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_,
    new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_,
    new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_,
    new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_,
    new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_,
    new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_,
    new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_,
    new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_,
    new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_,
    new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_,
    new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_,
    new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_,
    new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_,
    new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_,
    new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_,
    new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_,
    new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_,
    new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_,
    new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_,
    new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_,
    new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_,
    new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_,
    new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_,
    new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_,
    new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_,
    new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_,
    new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_,
    new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_,
    new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_,
    new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_,
    new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_,
    new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_,
    new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_,
    new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_,
    new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_,
    new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_,
    new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_,
    new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_,
    new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_,
    new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_,
    new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_,
    new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_,
    new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_,
    new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_,
    new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_,
    new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_,
    new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_,
    new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_,
    new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_,
    new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_,
    new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_,
    new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_,
    new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_,
    new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_,
    new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_,
    new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_,
    new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_,
    new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_,
    new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_,
    new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_,
    new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_,
    new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_,
    new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_,
    new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_,
    new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_,
    new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_,
    new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_,
    new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_,
    new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_,
    new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_,
    new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_,
    new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_,
    new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_,
    new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_,
    new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_,
    new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_,
    new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_,
    new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_,
    new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_,
    new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_,
    new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_,
    new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_,
    new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_,
    new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_,
    new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_,
    new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_,
    new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_,
    new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_,
    new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_,
    new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_,
    new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_,
    new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_,
    new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_,
    new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_,
    new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_,
    new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_,
    new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_,
    new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_,
    new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_,
    new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_,
    new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_,
    new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_,
    new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_,
    new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_,
    new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_,
    new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_,
    new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_,
    new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_,
    new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_,
    new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_,
    new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_,
    new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_,
    new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_,
    new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_,
    new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_,
    new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_,
    new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_,
    new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_,
    new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_,
    new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_,
    new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_,
    new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_,
    new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_,
    new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_,
    new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_,
    new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_,
    new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_,
    new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_,
    new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_,
    new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_,
    new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_,
    new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_,
    new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_,
    new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_,
    new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_,
    new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_,
    new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_,
    new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_,
    new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_,
    new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_,
    new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_,
    new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_,
    new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_,
    new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_,
    new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_,
    new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_,
    new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_,
    new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_,
    new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_,
    new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_,
    new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_,
    new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_,
    new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_,
    new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_,
    new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_,
    new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_,
    new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_,
    new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_,
    new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_,
    new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_,
    new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_,
    new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_,
    new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_,
    new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_,
    new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_,
    new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_,
    new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_,
    new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_,
    new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_,
    new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_,
    new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_,
    new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_,
    new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_,
    new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_,
    new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_,
    new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_,
    new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_,
    new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_,
    new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_,
    new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_,
    new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_,
    new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_,
    new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_,
    new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_,
    new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_,
    new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_,
    new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_,
    new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_,
    new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_,
    new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_,
    new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_,
    new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_,
    new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_,
    new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_,
    new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_,
    new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_,
    new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_,
    new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_,
    new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_,
    new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_,
    new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_,
    new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_,
    new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_,
    new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_,
    new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_,
    new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_,
    new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_,
    new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_,
    new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_,
    new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_,
    new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_,
    new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_,
    new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_,
    new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_,
    new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_,
    new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_,
    new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_,
    new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_,
    new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_,
    new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_,
    new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_,
    new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_,
    new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_,
    new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_,
    new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_,
    new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_,
    new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_,
    new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_,
    new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_,
    new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_,
    new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_,
    new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_,
    new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_,
    new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_,
    new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_,
    new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_,
    new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_,
    new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_,
    new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_,
    new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_,
    new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_,
    new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_,
    new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_,
    new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_,
    new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_,
    new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_,
    new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_,
    new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_,
    new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_,
    new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_,
    new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_,
    new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_,
    new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_,
    new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_,
    new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_,
    new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_,
    new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_,
    new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_,
    new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_,
    new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_,
    new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_,
    new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_,
    new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_,
    new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_,
    new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_,
    new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_,
    new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_,
    new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_,
    new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_,
    new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_,
    new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_,
    new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_,
    new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_,
    new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_,
    new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_,
    new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_,
    new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_,
    new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_,
    new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_,
    new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_,
    new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_,
    new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_,
    new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_,
    new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_,
    new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_,
    new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_,
    new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_,
    new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_,
    new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_,
    new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_,
    new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_,
    new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_,
    new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_,
    new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_,
    new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_,
    new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_,
    new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_,
    new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_,
    new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_,
    new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_,
    new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_,
    new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_,
    new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_,
    new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_,
    new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_,
    new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_,
    new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_,
    new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_,
    new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_,
    new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_,
    new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_,
    new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_,
    new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_,
    new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_,
    new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_,
    new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_,
    new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_,
    new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_,
    new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_,
    new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_,
    new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_,
    new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_,
    new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_,
    new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_,
    new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_,
    new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_,
    new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_,
    new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_,
    new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_,
    new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_,
    new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_,
    new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_,
    new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_,
    new_n9997_, new_n9998_, new_n9999_, new_n10000_, new_n10001_,
    new_n10002_, new_n10003_, new_n10004_, new_n10005_, new_n10006_,
    new_n10007_, new_n10008_, new_n10009_, new_n10010_, new_n10011_,
    new_n10012_, new_n10013_, new_n10014_, new_n10015_, new_n10016_,
    new_n10017_, new_n10018_, new_n10019_, new_n10020_, new_n10021_,
    new_n10022_, new_n10023_, new_n10024_, new_n10025_, new_n10026_,
    new_n10027_, new_n10028_, new_n10029_, new_n10030_, new_n10031_,
    new_n10032_, new_n10033_, new_n10034_, new_n10035_, new_n10036_,
    new_n10037_, new_n10038_, new_n10039_, new_n10040_, new_n10041_,
    new_n10042_, new_n10043_, new_n10044_, new_n10045_, new_n10046_,
    new_n10047_, new_n10048_, new_n10049_, new_n10050_, new_n10051_,
    new_n10052_, new_n10053_, new_n10054_, new_n10055_, new_n10056_,
    new_n10057_, new_n10058_, new_n10059_, new_n10060_, new_n10061_,
    new_n10062_, new_n10063_, new_n10064_, new_n10065_, new_n10066_,
    new_n10067_, new_n10068_, new_n10069_, new_n10070_, new_n10071_,
    new_n10072_, new_n10073_, new_n10074_, new_n10075_, new_n10076_,
    new_n10077_, new_n10078_, new_n10079_, new_n10080_, new_n10081_,
    new_n10082_, new_n10083_, new_n10084_, new_n10085_, new_n10086_,
    new_n10087_, new_n10088_, new_n10089_, new_n10090_, new_n10091_,
    new_n10092_, new_n10093_, new_n10094_, new_n10095_, new_n10096_,
    new_n10097_, new_n10098_, new_n10099_, new_n10100_, new_n10101_,
    new_n10102_, new_n10103_, new_n10104_, new_n10105_, new_n10106_,
    new_n10107_, new_n10108_, new_n10109_, new_n10110_, new_n10111_,
    new_n10112_, new_n10113_, new_n10114_, new_n10115_, new_n10116_,
    new_n10117_, new_n10118_, new_n10119_, new_n10120_, new_n10121_,
    new_n10122_, new_n10123_, new_n10124_, new_n10125_, new_n10126_,
    new_n10127_, new_n10128_, new_n10129_, new_n10130_, new_n10131_,
    new_n10132_, new_n10133_, new_n10134_, new_n10135_, new_n10136_,
    new_n10137_, new_n10138_, new_n10139_, new_n10140_, new_n10141_,
    new_n10142_, new_n10143_, new_n10144_, new_n10145_, new_n10146_,
    new_n10147_, new_n10148_, new_n10149_, new_n10150_, new_n10151_,
    new_n10152_, new_n10153_, new_n10154_, new_n10155_, new_n10156_,
    new_n10157_, new_n10158_, new_n10159_, new_n10160_, new_n10161_,
    new_n10162_, new_n10163_, new_n10164_, new_n10165_, new_n10166_,
    new_n10167_, new_n10168_, new_n10169_, new_n10170_, new_n10171_,
    new_n10172_, new_n10173_, new_n10174_, new_n10175_, new_n10176_,
    new_n10177_, new_n10178_, new_n10179_, new_n10180_, new_n10181_,
    new_n10182_, new_n10183_, new_n10184_, new_n10185_, new_n10186_,
    new_n10187_, new_n10188_, new_n10189_, new_n10190_, new_n10191_,
    new_n10192_, new_n10193_, new_n10194_, new_n10195_, new_n10196_,
    new_n10197_, new_n10198_, new_n10199_, new_n10200_, new_n10201_,
    new_n10202_, new_n10203_, new_n10204_, new_n10205_, new_n10206_,
    new_n10207_, new_n10208_, new_n10209_, new_n10210_, new_n10211_,
    new_n10212_, new_n10213_, new_n10214_, new_n10215_, new_n10216_,
    new_n10217_, new_n10218_, new_n10219_, new_n10220_, new_n10221_,
    new_n10222_, new_n10223_, new_n10224_, new_n10225_, new_n10226_,
    new_n10227_, new_n10228_, new_n10229_, new_n10230_, new_n10231_,
    new_n10232_, new_n10233_, new_n10234_, new_n10235_, new_n10236_,
    new_n10237_, new_n10238_, new_n10239_, new_n10240_, new_n10241_,
    new_n10242_, new_n10243_, new_n10244_, new_n10245_, new_n10246_,
    new_n10247_, new_n10248_, new_n10249_, new_n10250_, new_n10251_,
    new_n10252_, new_n10253_, new_n10254_, new_n10255_, new_n10256_,
    new_n10257_, new_n10258_, new_n10259_, new_n10260_, new_n10261_,
    new_n10262_, new_n10263_, new_n10264_, new_n10265_, new_n10266_,
    new_n10267_, new_n10268_, new_n10269_, new_n10270_, new_n10271_,
    new_n10272_, new_n10273_, new_n10274_, new_n10275_, new_n10276_,
    new_n10277_, new_n10278_, new_n10279_, new_n10280_, new_n10281_,
    new_n10282_, new_n10283_, new_n10284_, new_n10285_, new_n10286_,
    new_n10287_, new_n10288_, new_n10289_, new_n10290_, new_n10291_,
    new_n10292_, new_n10293_, new_n10294_, new_n10295_, new_n10296_,
    new_n10297_, new_n10298_, new_n10299_, new_n10300_, new_n10301_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10311_,
    new_n10312_, new_n10313_, new_n10314_, new_n10315_, new_n10316_,
    new_n10317_, new_n10318_, new_n10319_, new_n10320_, new_n10321_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10330_, new_n10331_,
    new_n10332_, new_n10333_, new_n10334_, new_n10335_, new_n10336_,
    new_n10337_, new_n10338_, new_n10339_, new_n10340_, new_n10341_,
    new_n10342_, new_n10343_, new_n10344_, new_n10345_, new_n10346_,
    new_n10347_, new_n10348_, new_n10349_, new_n10350_, new_n10351_,
    new_n10352_, new_n10353_, new_n10354_, new_n10355_, new_n10356_,
    new_n10357_, new_n10358_, new_n10359_, new_n10360_, new_n10361_,
    new_n10362_, new_n10363_, new_n10364_, new_n10365_, new_n10366_,
    new_n10367_, new_n10368_, new_n10369_, new_n10370_, new_n10371_,
    new_n10372_, new_n10373_, new_n10374_, new_n10375_, new_n10376_,
    new_n10377_, new_n10378_, new_n10379_, new_n10380_, new_n10381_,
    new_n10382_, new_n10383_, new_n10384_, new_n10385_, new_n10386_,
    new_n10387_, new_n10388_, new_n10389_, new_n10390_, new_n10391_,
    new_n10392_, new_n10393_, new_n10394_, new_n10395_, new_n10396_,
    new_n10397_, new_n10398_, new_n10399_, new_n10400_, new_n10401_,
    new_n10402_, new_n10403_, new_n10404_, new_n10405_, new_n10406_,
    new_n10407_, new_n10408_, new_n10409_, new_n10410_, new_n10411_,
    new_n10412_, new_n10413_, new_n10414_, new_n10415_, new_n10416_,
    new_n10417_, new_n10418_, new_n10419_, new_n10420_, new_n10421_,
    new_n10422_, new_n10423_, new_n10424_, new_n10425_, new_n10426_,
    new_n10427_, new_n10428_, new_n10429_, new_n10430_, new_n10431_,
    new_n10432_, new_n10433_, new_n10434_, new_n10435_, new_n10436_,
    new_n10437_, new_n10438_, new_n10439_, new_n10440_, new_n10441_,
    new_n10442_, new_n10443_, new_n10444_, new_n10445_, new_n10446_,
    new_n10447_, new_n10448_, new_n10449_, new_n10450_, new_n10451_,
    new_n10452_, new_n10453_, new_n10454_, new_n10455_, new_n10456_,
    new_n10457_, new_n10458_, new_n10459_, new_n10460_, new_n10461_,
    new_n10462_, new_n10463_, new_n10464_, new_n10465_, new_n10466_,
    new_n10467_, new_n10468_, new_n10469_, new_n10470_, new_n10471_,
    new_n10472_, new_n10473_, new_n10474_, new_n10475_, new_n10476_,
    new_n10477_, new_n10478_, new_n10479_, new_n10480_, new_n10481_,
    new_n10482_, new_n10483_, new_n10484_, new_n10485_, new_n10486_,
    new_n10487_, new_n10488_, new_n10489_, new_n10490_, new_n10491_,
    new_n10492_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10621_,
    new_n10622_, new_n10623_, new_n10624_, new_n10625_, new_n10626_,
    new_n10627_, new_n10628_, new_n10629_, new_n10630_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10730_, new_n10731_,
    new_n10732_, new_n10733_, new_n10734_, new_n10735_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10751_,
    new_n10752_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10764_, new_n10765_, new_n10766_,
    new_n10767_, new_n10768_, new_n10769_, new_n10770_, new_n10771_,
    new_n10772_, new_n10773_, new_n10774_, new_n10775_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10794_, new_n10795_, new_n10796_,
    new_n10797_, new_n10798_, new_n10799_, new_n10800_, new_n10801_,
    new_n10802_, new_n10803_, new_n10804_, new_n10805_, new_n10806_,
    new_n10807_, new_n10808_, new_n10809_, new_n10810_, new_n10811_,
    new_n10812_, new_n10813_, new_n10814_, new_n10815_, new_n10816_,
    new_n10817_, new_n10818_, new_n10819_, new_n10820_, new_n10821_,
    new_n10822_, new_n10823_, new_n10824_, new_n10825_, new_n10826_,
    new_n10827_, new_n10828_, new_n10829_, new_n10830_, new_n10831_,
    new_n10832_, new_n10833_, new_n10834_, new_n10835_, new_n10836_,
    new_n10837_, new_n10838_, new_n10839_, new_n10840_, new_n10841_,
    new_n10842_, new_n10843_, new_n10844_, new_n10845_, new_n10846_,
    new_n10847_, new_n10848_, new_n10849_, new_n10850_, new_n10851_,
    new_n10852_, new_n10853_, new_n10854_, new_n10855_, new_n10856_,
    new_n10857_, new_n10858_, new_n10859_, new_n10860_, new_n10861_,
    new_n10862_, new_n10863_, new_n10864_, new_n10865_, new_n10866_,
    new_n10867_, new_n10868_, new_n10869_, new_n10870_, new_n10871_,
    new_n10872_, new_n10873_, new_n10874_, new_n10875_, new_n10876_,
    new_n10877_, new_n10878_, new_n10879_, new_n10880_, new_n10881_,
    new_n10882_, new_n10883_, new_n10884_, new_n10885_, new_n10886_,
    new_n10887_, new_n10888_, new_n10889_, new_n10890_, new_n10891_,
    new_n10892_, new_n10893_, new_n10894_, new_n10895_, new_n10896_,
    new_n10897_, new_n10898_, new_n10899_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11221_,
    new_n11222_, new_n11223_, new_n11224_, new_n11225_, new_n11226_,
    new_n11227_, new_n11228_, new_n11229_, new_n11230_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11371_,
    new_n11372_, new_n11373_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11392_, new_n11393_, new_n11394_, new_n11395_, new_n11396_,
    new_n11397_, new_n11398_, new_n11399_, new_n11400_, new_n11401_,
    new_n11402_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11415_, new_n11416_,
    new_n11417_, new_n11418_, new_n11419_, new_n11420_, new_n11421_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11440_, new_n11441_,
    new_n11442_, new_n11443_, new_n11444_, new_n11445_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11460_, new_n11461_,
    new_n11462_, new_n11463_, new_n11464_, new_n11465_, new_n11466_,
    new_n11467_, new_n11468_, new_n11469_, new_n11470_, new_n11471_,
    new_n11472_, new_n11473_, new_n11474_, new_n11475_, new_n11476_,
    new_n11477_, new_n11478_, new_n11479_, new_n11480_, new_n11481_,
    new_n11482_, new_n11483_, new_n11484_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11499_, new_n11500_, new_n11501_,
    new_n11502_, new_n11503_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11510_, new_n11511_,
    new_n11512_, new_n11513_, new_n11514_, new_n11515_, new_n11516_,
    new_n11517_, new_n11518_, new_n11519_, new_n11520_, new_n11521_,
    new_n11522_, new_n11523_, new_n11524_, new_n11525_, new_n11526_,
    new_n11527_, new_n11528_, new_n11529_, new_n11530_, new_n11531_,
    new_n11532_, new_n11533_, new_n11534_, new_n11535_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11543_, new_n11544_, new_n11545_, new_n11546_,
    new_n11547_, new_n11548_, new_n11549_, new_n11550_, new_n11551_,
    new_n11552_, new_n11553_, new_n11554_, new_n11555_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12100_, new_n12101_,
    new_n12102_, new_n12103_, new_n12104_, new_n12105_, new_n12106_,
    new_n12107_, new_n12108_, new_n12109_, new_n12110_, new_n12111_,
    new_n12112_, new_n12113_, new_n12114_, new_n12115_, new_n12116_,
    new_n12117_, new_n12118_, new_n12119_, new_n12120_, new_n12121_,
    new_n12122_, new_n12123_, new_n12124_, new_n12125_, new_n12126_,
    new_n12127_, new_n12128_, new_n12129_, new_n12130_, new_n12131_,
    new_n12132_, new_n12133_, new_n12134_, new_n12135_, new_n12136_,
    new_n12137_, new_n12138_, new_n12139_, new_n12140_, new_n12141_,
    new_n12142_, new_n12143_, new_n12144_, new_n12145_, new_n12146_,
    new_n12147_, new_n12148_, new_n12149_, new_n12150_, new_n12151_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12158_, new_n12159_, new_n12160_, new_n12161_,
    new_n12162_, new_n12163_, new_n12164_, new_n12165_, new_n12166_,
    new_n12167_, new_n12168_, new_n12169_, new_n12170_, new_n12171_,
    new_n12172_, new_n12173_, new_n12174_, new_n12175_, new_n12176_,
    new_n12177_, new_n12178_, new_n12179_, new_n12180_, new_n12181_,
    new_n12182_, new_n12183_, new_n12184_, new_n12185_, new_n12186_,
    new_n12187_, new_n12188_, new_n12189_, new_n12190_, new_n12191_,
    new_n12192_, new_n12193_, new_n12194_, new_n12195_, new_n12196_,
    new_n12197_, new_n12198_, new_n12199_, new_n12200_, new_n12201_,
    new_n12202_, new_n12203_, new_n12204_, new_n12205_, new_n12206_,
    new_n12207_, new_n12208_, new_n12209_, new_n12210_, new_n12211_,
    new_n12212_, new_n12213_, new_n12214_, new_n12215_, new_n12216_,
    new_n12217_, new_n12218_, new_n12219_, new_n12220_, new_n12221_,
    new_n12222_, new_n12223_, new_n12224_, new_n12225_, new_n12226_,
    new_n12227_, new_n12228_, new_n12229_, new_n12230_, new_n12231_,
    new_n12232_, new_n12233_, new_n12234_, new_n12235_, new_n12236_,
    new_n12237_, new_n12238_, new_n12239_, new_n12240_, new_n12241_,
    new_n12242_, new_n12243_, new_n12244_, new_n12245_, new_n12246_,
    new_n12247_, new_n12248_, new_n12249_, new_n12250_, new_n12251_,
    new_n12252_, new_n12253_, new_n12254_, new_n12255_, new_n12256_,
    new_n12257_, new_n12258_, new_n12259_, new_n12260_, new_n12261_,
    new_n12262_, new_n12263_, new_n12264_, new_n12265_, new_n12266_,
    new_n12267_, new_n12268_, new_n12269_, new_n12270_, new_n12271_,
    new_n12272_, new_n12273_, new_n12274_, new_n12275_, new_n12276_,
    new_n12277_, new_n12278_, new_n12279_, new_n12280_, new_n12281_,
    new_n12282_, new_n12283_, new_n12284_, new_n12285_, new_n12286_,
    new_n12287_, new_n12288_, new_n12289_, new_n12290_, new_n12291_,
    new_n12292_, new_n12293_, new_n12294_, new_n12295_, new_n12296_,
    new_n12297_, new_n12298_, new_n12299_, new_n12300_, new_n12301_,
    new_n12302_, new_n12303_, new_n12304_, new_n12305_, new_n12306_,
    new_n12307_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12327_, new_n12328_, new_n12329_, new_n12330_, new_n12331_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12353_, new_n12354_, new_n12355_, new_n12356_,
    new_n12357_, new_n12358_, new_n12359_, new_n12360_, new_n12361_,
    new_n12362_, new_n12363_, new_n12364_, new_n12365_, new_n12366_,
    new_n12367_, new_n12368_, new_n12369_, new_n12370_, new_n12371_,
    new_n12372_, new_n12373_, new_n12374_, new_n12375_, new_n12376_,
    new_n12377_, new_n12378_, new_n12379_, new_n12380_, new_n12381_,
    new_n12382_, new_n12383_, new_n12384_, new_n12385_, new_n12386_,
    new_n12387_, new_n12388_, new_n12389_, new_n12390_, new_n12391_,
    new_n12392_, new_n12393_, new_n12394_, new_n12395_, new_n12396_,
    new_n12397_, new_n12398_, new_n12399_, new_n12400_, new_n12401_,
    new_n12402_, new_n12403_, new_n12404_, new_n12405_, new_n12406_,
    new_n12407_, new_n12408_, new_n12409_, new_n12410_, new_n12411_,
    new_n12412_, new_n12413_, new_n12414_, new_n12415_, new_n12416_,
    new_n12417_, new_n12418_, new_n12419_, new_n12420_, new_n12421_,
    new_n12422_, new_n12423_, new_n12424_, new_n12425_, new_n12426_,
    new_n12427_, new_n12428_, new_n12429_, new_n12430_, new_n12431_,
    new_n12432_, new_n12433_, new_n12434_, new_n12435_, new_n12436_,
    new_n12437_, new_n12438_, new_n12439_, new_n12440_, new_n12441_,
    new_n12442_, new_n12443_, new_n12444_, new_n12445_, new_n12446_,
    new_n12447_, new_n12448_, new_n12449_, new_n12450_, new_n12451_,
    new_n12452_, new_n12453_, new_n12454_, new_n12455_, new_n12456_,
    new_n12457_, new_n12458_, new_n12459_, new_n12460_, new_n12461_,
    new_n12462_, new_n12463_, new_n12464_, new_n12465_, new_n12466_,
    new_n12467_, new_n12468_, new_n12469_, new_n12470_, new_n12471_,
    new_n12472_, new_n12473_, new_n12474_, new_n12475_, new_n12476_,
    new_n12477_, new_n12478_, new_n12479_, new_n12480_, new_n12481_,
    new_n12482_, new_n12483_, new_n12484_, new_n12485_, new_n12486_,
    new_n12487_, new_n12488_, new_n12489_, new_n12490_, new_n12491_,
    new_n12492_, new_n12493_, new_n12494_, new_n12495_, new_n12496_,
    new_n12497_, new_n12498_, new_n12499_, new_n12500_, new_n12501_,
    new_n12502_, new_n12503_, new_n12504_, new_n12505_, new_n12506_,
    new_n12507_, new_n12508_, new_n12509_, new_n12510_, new_n12511_,
    new_n12512_, new_n12513_, new_n12514_, new_n12515_, new_n12516_,
    new_n12517_, new_n12518_, new_n12519_, new_n12520_, new_n12521_,
    new_n12522_, new_n12523_, new_n12524_, new_n12525_, new_n12526_,
    new_n12527_, new_n12528_, new_n12529_, new_n12530_, new_n12531_,
    new_n12532_, new_n12533_, new_n12534_, new_n12535_, new_n12536_,
    new_n12537_, new_n12538_, new_n12539_, new_n12540_, new_n12541_,
    new_n12542_, new_n12543_, new_n12544_, new_n12545_, new_n12546_,
    new_n12547_, new_n12548_, new_n12549_, new_n12550_, new_n12551_,
    new_n12552_, new_n12553_, new_n12554_, new_n12555_, new_n12556_,
    new_n12557_, new_n12558_, new_n12559_, new_n12560_, new_n12561_,
    new_n12562_, new_n12563_, new_n12564_, new_n12565_, new_n12566_,
    new_n12567_, new_n12568_, new_n12569_, new_n12570_, new_n12571_,
    new_n12572_, new_n12573_, new_n12574_, new_n12575_, new_n12576_,
    new_n12577_, new_n12578_, new_n12579_, new_n12580_, new_n12581_,
    new_n12582_, new_n12583_, new_n12584_, new_n12585_, new_n12586_,
    new_n12587_, new_n12588_, new_n12589_, new_n12590_, new_n12591_,
    new_n12592_, new_n12593_, new_n12594_, new_n12595_, new_n12596_,
    new_n12597_, new_n12598_, new_n12599_, new_n12600_, new_n12601_,
    new_n12602_, new_n12603_, new_n12604_, new_n12605_, new_n12606_,
    new_n12607_, new_n12608_, new_n12609_, new_n12610_, new_n12611_,
    new_n12612_, new_n12613_, new_n12614_, new_n12615_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12629_, new_n12630_, new_n12631_,
    new_n12632_, new_n12633_, new_n12634_, new_n12635_, new_n12636_,
    new_n12637_, new_n12638_, new_n12639_, new_n12640_, new_n12641_,
    new_n12642_, new_n12643_, new_n12644_, new_n12645_, new_n12646_,
    new_n12647_, new_n12648_, new_n12649_, new_n12650_, new_n12651_,
    new_n12652_, new_n12653_, new_n12654_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12664_, new_n12665_, new_n12666_,
    new_n12667_, new_n12668_, new_n12669_, new_n12670_, new_n12671_,
    new_n12672_, new_n12673_, new_n12674_, new_n12675_, new_n12676_,
    new_n12677_, new_n12678_, new_n12679_, new_n12680_, new_n12681_,
    new_n12682_, new_n12683_, new_n12684_, new_n12685_, new_n12686_,
    new_n12687_, new_n12688_, new_n12689_, new_n12690_, new_n12691_,
    new_n12692_, new_n12693_, new_n12694_, new_n12695_, new_n12696_,
    new_n12697_, new_n12698_, new_n12699_, new_n12700_, new_n12701_,
    new_n12702_, new_n12703_, new_n12704_, new_n12705_, new_n12706_,
    new_n12707_, new_n12708_, new_n12709_, new_n12710_, new_n12711_,
    new_n12712_, new_n12713_, new_n12714_, new_n12715_, new_n12716_,
    new_n12717_, new_n12718_, new_n12719_, new_n12720_, new_n12721_,
    new_n12722_, new_n12723_, new_n12724_, new_n12725_, new_n12726_,
    new_n12727_, new_n12728_, new_n12729_, new_n12730_, new_n12731_,
    new_n12732_, new_n12733_, new_n12734_, new_n12735_, new_n12736_,
    new_n12737_, new_n12738_, new_n12739_, new_n12740_, new_n12741_,
    new_n12742_, new_n12743_, new_n12744_, new_n12745_, new_n12746_,
    new_n12747_, new_n12748_, new_n12749_, new_n12750_, new_n12751_,
    new_n12752_, new_n12753_, new_n12754_, new_n12755_, new_n12756_,
    new_n12757_, new_n12758_, new_n12759_, new_n12760_, new_n12761_,
    new_n12762_, new_n12763_, new_n12764_, new_n12765_, new_n12766_,
    new_n12767_, new_n12768_, new_n12769_, new_n12770_, new_n12771_,
    new_n12772_, new_n12773_, new_n12774_, new_n12775_, new_n12776_,
    new_n12777_, new_n12778_, new_n12779_, new_n12780_, new_n12781_,
    new_n12782_, new_n12783_, new_n12784_, new_n12785_, new_n12786_,
    new_n12787_, new_n12788_, new_n12789_, new_n12790_, new_n12791_,
    new_n12792_, new_n12793_, new_n12794_, new_n12795_, new_n12796_,
    new_n12797_, new_n12798_, new_n12799_, new_n12800_, new_n12801_,
    new_n12802_, new_n12803_, new_n12804_, new_n12805_, new_n12806_,
    new_n12807_, new_n12808_, new_n12809_, new_n12810_, new_n12811_,
    new_n12812_, new_n12813_, new_n12814_, new_n12815_, new_n12816_,
    new_n12817_, new_n12818_, new_n12819_, new_n12820_, new_n12821_,
    new_n12822_, new_n12823_, new_n12824_, new_n12825_, new_n12826_,
    new_n12827_, new_n12828_, new_n12829_, new_n12830_, new_n12831_,
    new_n12832_, new_n12833_, new_n12834_, new_n12835_, new_n12836_,
    new_n12837_, new_n12838_, new_n12839_, new_n12840_, new_n12841_,
    new_n12842_, new_n12843_, new_n12844_, new_n12845_, new_n12846_,
    new_n12847_, new_n12848_, new_n12849_, new_n12850_, new_n12851_,
    new_n12852_, new_n12853_, new_n12854_, new_n12855_, new_n12856_,
    new_n12857_, new_n12858_, new_n12859_, new_n12860_, new_n12861_,
    new_n12862_, new_n12863_, new_n12864_, new_n12865_, new_n12866_,
    new_n12867_, new_n12868_, new_n12869_, new_n12870_, new_n12871_,
    new_n12872_, new_n12873_, new_n12874_, new_n12875_, new_n12876_,
    new_n12877_, new_n12878_, new_n12879_, new_n12880_, new_n12881_,
    new_n12882_, new_n12883_, new_n12884_, new_n12885_, new_n12886_,
    new_n12887_, new_n12888_, new_n12889_, new_n12890_, new_n12891_,
    new_n12892_, new_n12893_, new_n12894_, new_n12895_, new_n12896_,
    new_n12897_, new_n12898_, new_n12899_, new_n12900_, new_n12901_,
    new_n12902_, new_n12903_, new_n12904_, new_n12905_, new_n12906_,
    new_n12907_, new_n12908_, new_n12909_, new_n12910_, new_n12911_,
    new_n12912_, new_n12913_, new_n12914_, new_n12915_, new_n12916_,
    new_n12917_, new_n12918_, new_n12919_, new_n12920_, new_n12921_,
    new_n12922_, new_n12923_, new_n12924_, new_n12925_, new_n12926_,
    new_n12927_, new_n12928_, new_n12929_, new_n12930_, new_n12931_,
    new_n12932_, new_n12933_, new_n12934_, new_n12935_, new_n12936_,
    new_n12937_, new_n12938_, new_n12939_, new_n12940_, new_n12941_,
    new_n12942_, new_n12943_, new_n12944_, new_n12945_, new_n12946_,
    new_n12947_, new_n12948_, new_n12949_, new_n12950_, new_n12951_,
    new_n12952_, new_n12953_, new_n12954_, new_n12955_, new_n12956_,
    new_n12957_, new_n12958_, new_n12959_, new_n12960_, new_n12961_,
    new_n12962_, new_n12963_, new_n12964_, new_n12965_, new_n12966_,
    new_n12967_, new_n12968_, new_n12969_, new_n12970_, new_n12971_,
    new_n12972_, new_n12973_, new_n12974_, new_n12975_, new_n12976_,
    new_n12977_, new_n12978_, new_n12979_, new_n12980_, new_n12981_,
    new_n12982_, new_n12983_, new_n12984_, new_n12985_, new_n12986_,
    new_n12987_, new_n12988_, new_n12989_, new_n12990_, new_n12991_,
    new_n12992_, new_n12993_, new_n12994_, new_n12995_, new_n12996_,
    new_n12997_, new_n12998_, new_n12999_, new_n13000_, new_n13001_,
    new_n13002_, new_n13003_, new_n13004_, new_n13005_, new_n13006_,
    new_n13007_, new_n13008_, new_n13009_, new_n13010_, new_n13011_,
    new_n13012_, new_n13013_, new_n13014_, new_n13015_, new_n13016_,
    new_n13017_, new_n13018_, new_n13019_, new_n13020_, new_n13021_,
    new_n13022_, new_n13023_, new_n13024_, new_n13025_, new_n13026_,
    new_n13027_, new_n13028_, new_n13029_, new_n13030_, new_n13031_,
    new_n13032_, new_n13033_, new_n13034_, new_n13035_, new_n13036_,
    new_n13037_, new_n13038_, new_n13039_, new_n13040_, new_n13041_,
    new_n13042_, new_n13043_, new_n13044_, new_n13045_, new_n13046_,
    new_n13047_, new_n13048_, new_n13049_, new_n13050_, new_n13051_,
    new_n13052_, new_n13053_, new_n13054_, new_n13055_, new_n13056_,
    new_n13057_, new_n13058_, new_n13059_, new_n13060_, new_n13061_,
    new_n13062_, new_n13063_, new_n13064_, new_n13065_, new_n13066_,
    new_n13067_, new_n13068_, new_n13069_, new_n13070_, new_n13071_,
    new_n13072_, new_n13073_, new_n13074_, new_n13075_, new_n13076_,
    new_n13077_, new_n13078_, new_n13079_, new_n13080_, new_n13081_,
    new_n13082_, new_n13083_, new_n13084_, new_n13085_, new_n13086_,
    new_n13087_, new_n13088_, new_n13089_, new_n13090_, new_n13091_,
    new_n13092_, new_n13093_, new_n13094_, new_n13095_, new_n13096_,
    new_n13097_, new_n13098_, new_n13099_, new_n13100_, new_n13101_,
    new_n13102_, new_n13103_, new_n13104_, new_n13105_, new_n13106_,
    new_n13107_, new_n13108_, new_n13109_, new_n13110_, new_n13111_,
    new_n13112_, new_n13113_, new_n13114_, new_n13115_, new_n13116_,
    new_n13117_, new_n13118_, new_n13119_, new_n13120_, new_n13121_,
    new_n13122_, new_n13123_, new_n13124_, new_n13125_, new_n13126_,
    new_n13127_, new_n13128_, new_n13129_, new_n13130_, new_n13131_,
    new_n13132_, new_n13133_, new_n13134_, new_n13135_, new_n13136_,
    new_n13137_, new_n13138_, new_n13139_, new_n13140_, new_n13141_,
    new_n13142_, new_n13143_, new_n13144_, new_n13145_, new_n13146_,
    new_n13147_, new_n13148_, new_n13149_, new_n13150_, new_n13151_,
    new_n13152_, new_n13153_, new_n13154_, new_n13155_, new_n13156_,
    new_n13157_, new_n13158_, new_n13159_, new_n13160_, new_n13161_,
    new_n13162_, new_n13163_, new_n13164_, new_n13165_, new_n13166_,
    new_n13167_, new_n13168_, new_n13169_, new_n13170_, new_n13171_,
    new_n13172_, new_n13173_, new_n13174_, new_n13175_, new_n13176_,
    new_n13177_, new_n13178_, new_n13179_, new_n13180_, new_n13181_,
    new_n13182_, new_n13183_, new_n13184_, new_n13185_, new_n13186_,
    new_n13187_, new_n13188_, new_n13189_, new_n13190_, new_n13191_,
    new_n13192_, new_n13193_, new_n13194_, new_n13195_, new_n13196_,
    new_n13197_, new_n13198_, new_n13199_, new_n13200_, new_n13201_,
    new_n13202_, new_n13203_, new_n13204_, new_n13205_, new_n13206_,
    new_n13207_, new_n13208_, new_n13209_, new_n13210_, new_n13211_,
    new_n13212_, new_n13213_, new_n13214_, new_n13215_, new_n13216_,
    new_n13217_, new_n13218_, new_n13219_, new_n13220_, new_n13221_,
    new_n13222_, new_n13223_, new_n13224_, new_n13225_, new_n13226_,
    new_n13227_, new_n13228_, new_n13229_, new_n13230_, new_n13231_,
    new_n13232_, new_n13233_, new_n13234_, new_n13235_, new_n13236_,
    new_n13237_, new_n13238_, new_n13239_, new_n13240_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13245_, new_n13246_,
    new_n13247_, new_n13248_, new_n13249_, new_n13250_, new_n13251_,
    new_n13252_, new_n13253_, new_n13254_, new_n13255_, new_n13256_,
    new_n13257_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13262_, new_n13263_, new_n13264_, new_n13265_, new_n13266_,
    new_n13267_, new_n13268_, new_n13269_, new_n13270_, new_n13271_,
    new_n13272_, new_n13273_, new_n13274_, new_n13275_, new_n13276_,
    new_n13277_, new_n13278_, new_n13279_, new_n13280_, new_n13281_,
    new_n13282_, new_n13283_, new_n13284_, new_n13285_, new_n13286_,
    new_n13287_, new_n13288_, new_n13289_, new_n13290_, new_n13291_,
    new_n13292_, new_n13293_, new_n13294_, new_n13295_, new_n13296_,
    new_n13297_, new_n13298_, new_n13299_, new_n13300_, new_n13301_,
    new_n13302_, new_n13303_, new_n13304_, new_n13305_, new_n13306_,
    new_n13307_, new_n13308_, new_n13309_, new_n13310_, new_n13311_,
    new_n13312_, new_n13313_, new_n13314_, new_n13315_, new_n13316_,
    new_n13317_, new_n13318_, new_n13319_, new_n13320_, new_n13321_,
    new_n13322_, new_n13323_, new_n13324_, new_n13325_, new_n13326_,
    new_n13327_, new_n13328_, new_n13329_, new_n13330_, new_n13331_,
    new_n13332_, new_n13333_, new_n13334_, new_n13335_, new_n13336_,
    new_n13337_, new_n13338_, new_n13339_, new_n13340_, new_n13341_,
    new_n13342_, new_n13343_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13354_, new_n13355_, new_n13356_,
    new_n13357_, new_n13358_, new_n13359_, new_n13360_, new_n13361_,
    new_n13362_, new_n13363_, new_n13364_, new_n13365_, new_n13366_,
    new_n13367_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13373_, new_n13374_, new_n13375_, new_n13376_,
    new_n13377_, new_n13378_, new_n13379_, new_n13380_, new_n13381_,
    new_n13382_, new_n13383_, new_n13384_, new_n13385_, new_n13386_,
    new_n13387_, new_n13388_, new_n13389_, new_n13390_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13395_, new_n13396_,
    new_n13397_, new_n13398_, new_n13399_, new_n13400_, new_n13401_,
    new_n13402_, new_n13403_, new_n13404_, new_n13405_, new_n13406_,
    new_n13407_, new_n13408_, new_n13409_, new_n13410_, new_n13411_,
    new_n13412_, new_n13413_, new_n13414_, new_n13415_, new_n13416_,
    new_n13417_, new_n13418_, new_n13419_, new_n13420_, new_n13421_,
    new_n13422_, new_n13423_, new_n13424_, new_n13425_, new_n13426_,
    new_n13427_, new_n13428_, new_n13429_, new_n13430_, new_n13431_,
    new_n13432_, new_n13433_, new_n13434_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13473_, new_n13474_, new_n13475_, new_n13476_,
    new_n13477_, new_n13478_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14445_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14456_,
    new_n14457_, new_n14458_, new_n14459_, new_n14460_, new_n14461_,
    new_n14462_, new_n14463_, new_n14464_, new_n14465_, new_n14466_,
    new_n14467_, new_n14468_, new_n14469_, new_n14470_, new_n14471_,
    new_n14472_, new_n14473_, new_n14474_, new_n14475_, new_n14476_,
    new_n14477_, new_n14478_, new_n14479_, new_n14480_, new_n14481_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14487_, new_n14488_, new_n14489_, new_n14490_, new_n14491_,
    new_n14492_, new_n14493_, new_n14494_, new_n14495_, new_n14496_,
    new_n14497_, new_n14498_, new_n14499_, new_n14500_, new_n14501_,
    new_n14502_, new_n14503_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14522_, new_n14523_, new_n14524_, new_n14525_, new_n14526_,
    new_n14527_, new_n14528_, new_n14529_, new_n14530_, new_n14531_,
    new_n14532_, new_n14533_, new_n14534_, new_n14535_, new_n14536_,
    new_n14537_, new_n14538_, new_n14539_, new_n14540_, new_n14541_,
    new_n14542_, new_n14543_, new_n14544_, new_n14545_, new_n14546_,
    new_n14547_, new_n14548_, new_n14549_, new_n14550_, new_n14551_,
    new_n14552_, new_n14553_, new_n14554_, new_n14555_, new_n14556_,
    new_n14557_, new_n14558_, new_n14559_, new_n14560_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14575_, new_n14576_,
    new_n14577_, new_n14578_, new_n14579_, new_n14580_, new_n14581_,
    new_n14582_, new_n14583_, new_n14584_, new_n14585_, new_n14586_,
    new_n14587_, new_n14588_, new_n14589_, new_n14590_, new_n14591_,
    new_n14592_, new_n14593_, new_n14594_, new_n14595_, new_n14596_,
    new_n14597_, new_n14598_, new_n14599_, new_n14600_, new_n14601_,
    new_n14602_, new_n14603_, new_n14604_, new_n14605_, new_n14606_,
    new_n14607_, new_n14608_, new_n14609_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14620_, new_n14621_,
    new_n14622_, new_n14623_, new_n14624_, new_n14625_, new_n14626_,
    new_n14627_, new_n14628_, new_n14629_, new_n14630_, new_n14631_,
    new_n14632_, new_n14633_, new_n14634_, new_n14635_, new_n14636_,
    new_n14637_, new_n14638_, new_n14639_, new_n14640_, new_n14641_,
    new_n14642_, new_n14643_, new_n14644_, new_n14645_, new_n14646_,
    new_n14647_, new_n14648_, new_n14649_, new_n14650_, new_n14651_,
    new_n14652_, new_n14653_, new_n14654_, new_n14655_, new_n14656_,
    new_n14657_, new_n14658_, new_n14659_, new_n14660_, new_n14661_,
    new_n14662_, new_n14663_, new_n14664_, new_n14665_, new_n14666_,
    new_n14667_, new_n14668_, new_n14669_, new_n14670_, new_n14671_,
    new_n14672_, new_n14673_, new_n14674_, new_n14675_, new_n14676_,
    new_n14677_, new_n14678_, new_n14679_, new_n14680_, new_n14681_,
    new_n14682_, new_n14683_, new_n14684_, new_n14685_, new_n14686_,
    new_n14687_, new_n14688_, new_n14689_, new_n14690_, new_n14691_,
    new_n14692_, new_n14693_, new_n14694_, new_n14695_, new_n14696_,
    new_n14697_, new_n14698_, new_n14699_, new_n14700_, new_n14701_,
    new_n14702_, new_n14703_, new_n14704_, new_n14705_, new_n14706_,
    new_n14707_, new_n14708_, new_n14709_, new_n14710_, new_n14711_,
    new_n14712_, new_n14713_, new_n14714_, new_n14715_, new_n14716_,
    new_n14717_, new_n14718_, new_n14719_, new_n14720_, new_n14721_,
    new_n14722_, new_n14723_, new_n14724_, new_n14725_, new_n14726_,
    new_n14727_, new_n14728_, new_n14729_, new_n14730_, new_n14731_,
    new_n14732_, new_n14733_, new_n14734_, new_n14735_, new_n14736_,
    new_n14737_, new_n14738_, new_n14739_, new_n14740_, new_n14741_,
    new_n14742_, new_n14743_, new_n14744_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14781_,
    new_n14782_, new_n14783_, new_n14784_, new_n14785_, new_n14786_,
    new_n14787_, new_n14788_, new_n14789_, new_n14790_, new_n14791_,
    new_n14792_, new_n14793_, new_n14794_, new_n14795_, new_n14796_,
    new_n14797_, new_n14798_, new_n14799_, new_n14800_, new_n14801_,
    new_n14802_, new_n14803_, new_n14804_, new_n14805_, new_n14806_,
    new_n14807_, new_n14808_, new_n14809_, new_n14810_, new_n14811_,
    new_n14812_, new_n14813_, new_n14814_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14958_, new_n14959_, new_n14960_, new_n14961_,
    new_n14962_, new_n14963_, new_n14964_, new_n14965_, new_n14966_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14976_,
    new_n14977_, new_n14978_, new_n14979_, new_n14980_, new_n14981_,
    new_n14982_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15113_, new_n15114_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15127_, new_n15128_, new_n15129_, new_n15130_, new_n15131_,
    new_n15132_, new_n15133_, new_n15134_, new_n15135_, new_n15136_,
    new_n15137_, new_n15138_, new_n15139_, new_n15140_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15179_, new_n15180_, new_n15181_,
    new_n15182_, new_n15183_, new_n15184_, new_n15185_, new_n15186_,
    new_n15187_, new_n15188_, new_n15189_, new_n15190_, new_n15191_,
    new_n15192_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15206_,
    new_n15207_, new_n15208_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15213_, new_n15214_, new_n15215_, new_n15216_,
    new_n15217_, new_n15218_, new_n15219_, new_n15220_, new_n15221_,
    new_n15222_, new_n15223_, new_n15224_, new_n15225_, new_n15226_,
    new_n15227_, new_n15228_, new_n15229_, new_n15230_, new_n15231_,
    new_n15232_, new_n15233_, new_n15234_, new_n15235_, new_n15236_,
    new_n15237_, new_n15238_, new_n15239_, new_n15240_, new_n15241_,
    new_n15242_, new_n15243_, new_n15244_, new_n15245_, new_n15246_,
    new_n15247_, new_n15248_, new_n15249_, new_n15250_, new_n15251_,
    new_n15252_, new_n15253_, new_n15254_, new_n15255_, new_n15256_,
    new_n15257_, new_n15258_, new_n15259_, new_n15260_, new_n15261_,
    new_n15262_, new_n15263_, new_n15264_, new_n15265_, new_n15266_,
    new_n15267_, new_n15268_, new_n15269_, new_n15270_, new_n15271_,
    new_n15272_, new_n15273_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15280_, new_n15281_,
    new_n15282_, new_n15283_, new_n15284_, new_n15285_, new_n15286_,
    new_n15287_, new_n15288_, new_n15289_, new_n15290_, new_n15291_,
    new_n15292_, new_n15293_, new_n15294_, new_n15295_, new_n15296_,
    new_n15297_, new_n15298_, new_n15299_, new_n15300_, new_n15301_,
    new_n15302_, new_n15303_, new_n15304_, new_n15305_, new_n15306_,
    new_n15307_, new_n15308_, new_n15309_, new_n15310_, new_n15311_,
    new_n15312_, new_n15313_, new_n15314_, new_n15315_, new_n15316_,
    new_n15317_, new_n15318_, new_n15319_, new_n15320_, new_n15321_,
    new_n15322_, new_n15323_, new_n15324_, new_n15325_, new_n15326_,
    new_n15327_, new_n15328_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15434_, new_n15435_, new_n15436_,
    new_n15437_, new_n15438_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15470_, new_n15471_,
    new_n15472_, new_n15473_, new_n15474_, new_n15475_, new_n15476_,
    new_n15477_, new_n15478_, new_n15479_, new_n15480_, new_n15481_,
    new_n15482_, new_n15483_, new_n15484_, new_n15485_, new_n15486_,
    new_n15487_, new_n15488_, new_n15489_, new_n15490_, new_n15491_,
    new_n15492_, new_n15493_, new_n15494_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15544_, new_n15545_, new_n15546_,
    new_n15547_, new_n15548_, new_n15549_, new_n15550_, new_n15551_,
    new_n15552_, new_n15553_, new_n15554_, new_n15555_, new_n15556_,
    new_n15557_, new_n15558_, new_n15559_, new_n15560_, new_n15561_,
    new_n15562_, new_n15563_, new_n15564_, new_n15565_, new_n15566_,
    new_n15567_, new_n15568_, new_n15569_, new_n15570_, new_n15571_,
    new_n15572_, new_n15573_, new_n15574_, new_n15575_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15580_, new_n15581_,
    new_n15582_, new_n15583_, new_n15584_, new_n15585_, new_n15586_,
    new_n15587_, new_n15588_, new_n15589_, new_n15590_, new_n15591_,
    new_n15592_, new_n15593_, new_n15594_, new_n15595_, new_n15596_,
    new_n15597_, new_n15598_, new_n15599_, new_n15600_, new_n15601_,
    new_n15602_, new_n15603_, new_n15604_, new_n15605_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15611_,
    new_n15612_, new_n15613_, new_n15614_, new_n15615_, new_n15616_,
    new_n15617_, new_n15618_, new_n15619_, new_n15620_, new_n15621_,
    new_n15622_, new_n15623_, new_n15624_, new_n15625_, new_n15626_,
    new_n15627_, new_n15628_, new_n15629_, new_n15630_, new_n15631_,
    new_n15632_, new_n15633_, new_n15634_, new_n15635_, new_n15636_,
    new_n15637_, new_n15638_, new_n15639_, new_n15640_, new_n15641_,
    new_n15642_, new_n15643_, new_n15644_, new_n15645_, new_n15646_,
    new_n15647_, new_n15648_, new_n15649_, new_n15650_, new_n15651_,
    new_n15652_, new_n15653_, new_n15654_, new_n15655_, new_n15656_,
    new_n15657_, new_n15658_, new_n15659_, new_n15660_, new_n15661_,
    new_n15662_, new_n15663_, new_n15664_, new_n15665_, new_n15666_,
    new_n15667_, new_n15668_, new_n15669_, new_n15670_, new_n15671_,
    new_n15672_, new_n15673_, new_n15674_, new_n15675_, new_n15676_,
    new_n15677_, new_n15678_, new_n15679_, new_n15680_, new_n15681_,
    new_n15682_, new_n15683_, new_n15684_, new_n15685_, new_n15686_,
    new_n15687_, new_n15688_, new_n15689_, new_n15690_, new_n15691_,
    new_n15692_, new_n15693_, new_n15694_, new_n15695_, new_n15696_,
    new_n15697_, new_n15698_, new_n15699_, new_n15700_, new_n15701_,
    new_n15702_, new_n15703_, new_n15704_, new_n15705_, new_n15706_,
    new_n15707_, new_n15708_, new_n15709_, new_n15710_, new_n15711_,
    new_n15712_, new_n15713_, new_n15714_, new_n15715_, new_n15716_,
    new_n15717_, new_n15718_, new_n15719_, new_n15720_, new_n15721_,
    new_n15722_, new_n15723_, new_n15724_, new_n15725_, new_n15726_,
    new_n15727_, new_n15728_, new_n15729_, new_n15730_, new_n15731_,
    new_n15732_, new_n15733_, new_n15734_, new_n15735_, new_n15736_,
    new_n15737_, new_n15738_, new_n15739_, new_n15740_, new_n15741_,
    new_n15742_, new_n15743_, new_n15744_, new_n15745_, new_n15746_,
    new_n15747_, new_n15748_, new_n15749_, new_n15750_, new_n15751_,
    new_n15752_, new_n15753_, new_n15754_, new_n15755_, new_n15756_,
    new_n15757_, new_n15758_, new_n15759_, new_n15760_, new_n15761_,
    new_n15762_, new_n15763_, new_n15764_, new_n15765_, new_n15766_,
    new_n15767_, new_n15768_, new_n15769_, new_n15770_, new_n15771_,
    new_n15772_, new_n15773_, new_n15774_, new_n15775_, new_n15776_,
    new_n15777_, new_n15778_, new_n15779_, new_n15780_, new_n15781_,
    new_n15782_, new_n15783_, new_n15784_, new_n15785_, new_n15786_,
    new_n15787_, new_n15788_, new_n15789_, new_n15790_, new_n15791_,
    new_n15792_, new_n15793_, new_n15794_, new_n15795_, new_n15796_,
    new_n15797_, new_n15798_, new_n15799_, new_n15800_, new_n15801_,
    new_n15802_, new_n15803_, new_n15804_, new_n15805_, new_n15806_,
    new_n15807_, new_n15808_, new_n15809_, new_n15810_, new_n15811_,
    new_n15812_, new_n15813_, new_n15814_, new_n15815_, new_n15816_,
    new_n15817_, new_n15818_, new_n15819_, new_n15820_, new_n15821_,
    new_n15822_, new_n15823_, new_n15824_, new_n15825_, new_n15826_,
    new_n15827_, new_n15828_, new_n15829_, new_n15830_, new_n15831_,
    new_n15832_, new_n15833_, new_n15834_, new_n15835_, new_n15836_,
    new_n15837_, new_n15838_, new_n15839_, new_n15840_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15850_, new_n15851_,
    new_n15852_, new_n15853_, new_n15854_, new_n15855_, new_n15856_,
    new_n15857_, new_n15858_, new_n15859_, new_n15860_, new_n15861_,
    new_n15862_, new_n15863_, new_n15864_, new_n15865_, new_n15866_,
    new_n15867_, new_n15868_, new_n15869_, new_n15870_, new_n15871_,
    new_n15872_, new_n15873_, new_n15874_, new_n15875_, new_n15876_,
    new_n15877_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15889_, new_n15890_, new_n15891_,
    new_n15892_, new_n15893_, new_n15894_, new_n15895_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15925_, new_n15926_,
    new_n15927_, new_n15928_, new_n15929_, new_n15930_, new_n15931_,
    new_n15932_, new_n15933_, new_n15934_, new_n15935_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16011_,
    new_n16012_, new_n16013_, new_n16014_, new_n16015_, new_n16016_,
    new_n16017_, new_n16018_, new_n16019_, new_n16020_, new_n16021_,
    new_n16022_, new_n16023_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16040_, new_n16041_,
    new_n16042_, new_n16043_, new_n16044_, new_n16045_, new_n16046_,
    new_n16047_, new_n16048_, new_n16049_, new_n16050_, new_n16051_,
    new_n16052_, new_n16053_, new_n16054_, new_n16055_, new_n16056_,
    new_n16057_, new_n16058_, new_n16059_, new_n16060_, new_n16061_,
    new_n16062_, new_n16063_, new_n16064_, new_n16065_, new_n16066_,
    new_n16067_, new_n16068_, new_n16069_, new_n16070_, new_n16071_,
    new_n16072_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16082_, new_n16083_, new_n16084_, new_n16085_, new_n16086_,
    new_n16087_, new_n16088_, new_n16089_, new_n16090_, new_n16091_,
    new_n16092_, new_n16093_, new_n16094_, new_n16095_, new_n16096_,
    new_n16097_, new_n16098_, new_n16099_, new_n16100_, new_n16101_,
    new_n16102_, new_n16103_, new_n16104_, new_n16105_, new_n16106_,
    new_n16107_, new_n16108_, new_n16109_, new_n16110_, new_n16111_,
    new_n16112_, new_n16113_, new_n16114_, new_n16115_, new_n16116_,
    new_n16117_, new_n16118_, new_n16119_, new_n16120_, new_n16121_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16164_, new_n16165_, new_n16166_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16295_, new_n16296_,
    new_n16297_, new_n16298_, new_n16299_, new_n16300_, new_n16301_,
    new_n16302_, new_n16303_, new_n16304_, new_n16305_, new_n16306_,
    new_n16307_, new_n16308_, new_n16309_, new_n16310_, new_n16311_,
    new_n16312_, new_n16313_, new_n16314_, new_n16315_, new_n16316_,
    new_n16317_, new_n16318_, new_n16319_, new_n16320_, new_n16321_,
    new_n16322_, new_n16323_, new_n16324_, new_n16325_, new_n16326_,
    new_n16327_, new_n16328_, new_n16329_, new_n16330_, new_n16331_,
    new_n16332_, new_n16333_, new_n16334_, new_n16335_, new_n16336_,
    new_n16337_, new_n16338_, new_n16339_, new_n16340_, new_n16341_,
    new_n16342_, new_n16343_, new_n16344_, new_n16345_, new_n16346_,
    new_n16347_, new_n16348_, new_n16349_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17283_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17328_, new_n17329_, new_n17330_, new_n17331_,
    new_n17332_, new_n17333_, new_n17334_, new_n17335_, new_n17336_,
    new_n17337_, new_n17338_, new_n17339_, new_n17340_, new_n17341_,
    new_n17342_, new_n17343_, new_n17344_, new_n17345_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17361_,
    new_n17362_, new_n17363_, new_n17364_, new_n17365_, new_n17366_,
    new_n17367_, new_n17368_, new_n17369_, new_n17370_, new_n17371_,
    new_n17372_, new_n17373_, new_n17374_, new_n17375_, new_n17376_,
    new_n17377_, new_n17378_, new_n17379_, new_n17380_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17398_, new_n17399_, new_n17400_, new_n17401_,
    new_n17402_, new_n17403_, new_n17404_, new_n17405_, new_n17406_,
    new_n17407_, new_n17408_, new_n17409_, new_n17410_, new_n17411_,
    new_n17412_, new_n17413_, new_n17414_, new_n17415_, new_n17416_,
    new_n17417_, new_n17418_, new_n17419_, new_n17420_, new_n17421_,
    new_n17422_, new_n17423_, new_n17424_, new_n17425_, new_n17426_,
    new_n17427_, new_n17428_, new_n17429_, new_n17430_, new_n17431_,
    new_n17432_, new_n17433_, new_n17434_, new_n17435_, new_n17436_,
    new_n17437_, new_n17438_, new_n17439_, new_n17440_, new_n17441_,
    new_n17442_, new_n17443_, new_n17444_, new_n17445_, new_n17446_,
    new_n17447_, new_n17448_, new_n17449_, new_n17450_, new_n17451_,
    new_n17452_, new_n17453_, new_n17454_, new_n17455_, new_n17456_,
    new_n17457_, new_n17458_, new_n17459_, new_n17460_, new_n17461_,
    new_n17462_, new_n17463_, new_n17464_, new_n17465_, new_n17466_,
    new_n17467_, new_n17468_, new_n17469_, new_n17470_, new_n17471_,
    new_n17472_, new_n17473_, new_n17474_, new_n17475_, new_n17476_,
    new_n17477_, new_n17478_, new_n17479_, new_n17480_, new_n17481_,
    new_n17482_, new_n17483_, new_n17484_, new_n17485_, new_n17486_,
    new_n17487_, new_n17488_, new_n17489_, new_n17490_, new_n17491_,
    new_n17492_, new_n17493_, new_n17494_, new_n17495_, new_n17496_,
    new_n17497_, new_n17498_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17504_, new_n17505_, new_n17506_,
    new_n17507_, new_n17508_, new_n17509_, new_n17510_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17516_,
    new_n17517_, new_n17518_, new_n17519_, new_n17520_, new_n17521_,
    new_n17522_, new_n17523_, new_n17524_, new_n17525_, new_n17526_,
    new_n17527_, new_n17528_, new_n17529_, new_n17530_, new_n17531_,
    new_n17532_, new_n17533_, new_n17534_, new_n17535_, new_n17536_,
    new_n17537_, new_n17538_, new_n17539_, new_n17540_, new_n17541_,
    new_n17542_, new_n17543_, new_n17544_, new_n17545_, new_n17546_,
    new_n17547_, new_n17548_, new_n17549_, new_n17550_, new_n17551_,
    new_n17552_, new_n17553_, new_n17554_, new_n17555_, new_n17556_,
    new_n17557_, new_n17558_, new_n17559_, new_n17560_, new_n17561_,
    new_n17562_, new_n17563_, new_n17564_, new_n17565_, new_n17566_,
    new_n17567_, new_n17568_, new_n17569_, new_n17570_, new_n17571_,
    new_n17572_, new_n17573_, new_n17574_, new_n17575_, new_n17576_,
    new_n17577_, new_n17578_, new_n17579_, new_n17580_, new_n17581_,
    new_n17582_, new_n17583_, new_n17584_, new_n17585_, new_n17586_,
    new_n17587_, new_n17588_, new_n17589_, new_n17590_, new_n17591_,
    new_n17592_, new_n17593_, new_n17594_, new_n17595_, new_n17596_,
    new_n17597_, new_n17598_, new_n17599_, new_n17600_, new_n17601_,
    new_n17602_, new_n17603_, new_n17604_, new_n17605_, new_n17606_,
    new_n17607_, new_n17608_, new_n17609_, new_n17610_, new_n17611_,
    new_n17612_, new_n17613_, new_n17614_, new_n17615_, new_n17616_,
    new_n17617_, new_n17618_, new_n17619_, new_n17620_, new_n17621_,
    new_n17622_, new_n17623_, new_n17624_, new_n17625_, new_n17626_,
    new_n17627_, new_n17628_, new_n17629_, new_n17630_, new_n17631_,
    new_n17632_, new_n17633_, new_n17634_, new_n17635_, new_n17636_,
    new_n17637_, new_n17638_, new_n17639_, new_n17640_, new_n17641_,
    new_n17642_, new_n17643_, new_n17644_, new_n17645_, new_n17646_,
    new_n17647_, new_n17648_, new_n17649_, new_n17650_, new_n17651_,
    new_n17652_, new_n17653_, new_n17654_, new_n17655_, new_n17656_,
    new_n17657_, new_n17658_, new_n17659_, new_n17660_, new_n17661_,
    new_n17662_, new_n17663_, new_n17664_, new_n17665_, new_n17666_,
    new_n17667_, new_n17668_, new_n17669_, new_n17670_, new_n17671_,
    new_n17672_, new_n17673_, new_n17674_, new_n17675_, new_n17676_,
    new_n17677_, new_n17678_, new_n17679_, new_n17680_, new_n17681_,
    new_n17682_, new_n17683_, new_n17684_, new_n17685_, new_n17686_,
    new_n17687_, new_n17688_, new_n17689_, new_n17690_, new_n17691_,
    new_n17692_, new_n17693_, new_n17694_, new_n17695_, new_n17696_,
    new_n17697_, new_n17698_, new_n17699_, new_n17700_, new_n17701_,
    new_n17702_, new_n17703_, new_n17704_, new_n17705_, new_n17706_,
    new_n17707_, new_n17708_, new_n17709_, new_n17710_, new_n17711_,
    new_n17712_, new_n17713_, new_n17714_, new_n17715_, new_n17716_,
    new_n17717_, new_n17718_, new_n17719_, new_n17720_, new_n17721_,
    new_n17722_, new_n17723_, new_n17724_, new_n17725_, new_n17726_,
    new_n17727_, new_n17728_, new_n17729_, new_n17730_, new_n17731_,
    new_n17732_, new_n17733_, new_n17734_, new_n17735_, new_n17736_,
    new_n17737_, new_n17738_, new_n17739_, new_n17740_, new_n17741_,
    new_n17742_, new_n17743_, new_n17744_, new_n17745_, new_n17746_,
    new_n17747_, new_n17748_, new_n17749_, new_n17750_, new_n17751_,
    new_n17752_, new_n17753_, new_n17754_, new_n17755_, new_n17756_,
    new_n17757_, new_n17758_, new_n17759_, new_n17760_, new_n17761_,
    new_n17762_, new_n17763_, new_n17764_, new_n17765_, new_n17766_,
    new_n17767_, new_n17768_, new_n17769_, new_n17770_, new_n17771_,
    new_n17772_, new_n17773_, new_n17774_, new_n17775_, new_n17776_,
    new_n17777_, new_n17778_, new_n17779_, new_n17780_, new_n17781_,
    new_n17782_, new_n17783_, new_n17784_, new_n17785_, new_n17786_,
    new_n17787_, new_n17788_, new_n17789_, new_n17790_, new_n17791_,
    new_n17792_, new_n17793_, new_n17794_, new_n17795_, new_n17796_,
    new_n17797_, new_n17798_, new_n17799_, new_n17800_, new_n17801_,
    new_n17802_, new_n17803_, new_n17804_, new_n17805_, new_n17806_,
    new_n17807_, new_n17808_, new_n17809_, new_n17810_, new_n17811_,
    new_n17812_, new_n17813_, new_n17814_, new_n17815_, new_n17816_,
    new_n17817_, new_n17818_, new_n17819_, new_n17820_, new_n17821_,
    new_n17822_, new_n17823_, new_n17824_, new_n17825_, new_n17826_,
    new_n17827_, new_n17828_, new_n17829_, new_n17830_, new_n17831_,
    new_n17832_, new_n17833_, new_n17834_, new_n17835_, new_n17836_,
    new_n17837_, new_n17838_, new_n17839_, new_n17840_, new_n17841_,
    new_n17842_, new_n17843_, new_n17844_, new_n17845_, new_n17846_,
    new_n17847_, new_n17848_, new_n17849_, new_n17850_, new_n17851_,
    new_n17852_, new_n17853_, new_n17854_, new_n17855_, new_n17856_,
    new_n17857_, new_n17858_, new_n17859_, new_n17860_, new_n17861_,
    new_n17862_, new_n17863_, new_n17864_, new_n17865_, new_n17866_,
    new_n17867_, new_n17868_, new_n17869_, new_n17870_, new_n17871_,
    new_n17872_, new_n17873_, new_n17874_, new_n17875_, new_n17876_,
    new_n17877_, new_n17878_, new_n17879_, new_n17880_, new_n17881_,
    new_n17882_, new_n17883_, new_n17884_, new_n17885_, new_n17886_,
    new_n17887_, new_n17888_, new_n17889_, new_n17890_, new_n17891_,
    new_n17892_, new_n17893_, new_n17894_, new_n17895_, new_n17896_,
    new_n17897_, new_n17898_, new_n17899_, new_n17900_, new_n17901_,
    new_n17902_, new_n17903_, new_n17904_, new_n17905_, new_n17906_,
    new_n17907_, new_n17908_, new_n17909_, new_n17910_, new_n17911_,
    new_n17912_, new_n17913_, new_n17914_, new_n17915_, new_n17916_,
    new_n17917_, new_n17918_, new_n17919_, new_n17920_, new_n17921_,
    new_n17922_, new_n17923_, new_n17924_, new_n17925_, new_n17926_,
    new_n17927_, new_n17928_, new_n17929_, new_n17930_, new_n17931_,
    new_n17932_, new_n17933_, new_n17934_, new_n17935_, new_n17936_,
    new_n17937_, new_n17938_, new_n17939_, new_n17940_, new_n17941_,
    new_n17942_, new_n17943_, new_n17944_, new_n17945_, new_n17946_,
    new_n17947_, new_n17948_, new_n17949_, new_n17950_, new_n17951_,
    new_n17952_, new_n17953_, new_n17954_, new_n17955_, new_n17956_,
    new_n17957_, new_n17958_, new_n17959_, new_n17960_, new_n17961_,
    new_n17962_, new_n17963_, new_n17964_, new_n17965_, new_n17966_,
    new_n17967_, new_n17968_, new_n17969_, new_n17970_, new_n17971_,
    new_n17972_, new_n17973_, new_n17974_, new_n17975_, new_n17976_,
    new_n17977_, new_n17978_, new_n17979_, new_n17980_, new_n17981_,
    new_n17982_, new_n17983_, new_n17984_, new_n17985_, new_n17986_,
    new_n17987_, new_n17988_, new_n17989_, new_n17990_, new_n17991_,
    new_n17992_, new_n17993_, new_n17994_, new_n17995_, new_n17996_,
    new_n17997_, new_n17998_, new_n17999_, new_n18000_, new_n18001_,
    new_n18002_, new_n18003_, new_n18004_, new_n18005_, new_n18006_,
    new_n18007_, new_n18008_, new_n18009_, new_n18010_, new_n18011_,
    new_n18012_, new_n18013_, new_n18014_, new_n18015_, new_n18016_,
    new_n18017_, new_n18018_, new_n18019_, new_n18020_, new_n18021_,
    new_n18022_, new_n18023_, new_n18024_, new_n18025_, new_n18026_,
    new_n18027_, new_n18028_, new_n18029_, new_n18030_, new_n18031_,
    new_n18032_, new_n18033_, new_n18034_, new_n18035_, new_n18036_,
    new_n18037_, new_n18038_, new_n18039_, new_n18040_, new_n18041_,
    new_n18042_, new_n18043_, new_n18044_, new_n18045_, new_n18046_,
    new_n18047_, new_n18048_, new_n18049_, new_n18050_, new_n18051_,
    new_n18052_, new_n18053_, new_n18054_, new_n18055_, new_n18056_,
    new_n18057_, new_n18058_, new_n18059_, new_n18060_, new_n18061_,
    new_n18062_, new_n18063_, new_n18064_, new_n18065_, new_n18066_,
    new_n18067_, new_n18068_, new_n18069_, new_n18070_, new_n18071_,
    new_n18072_, new_n18073_, new_n18074_, new_n18075_, new_n18076_,
    new_n18077_, new_n18078_, new_n18079_, new_n18080_, new_n18081_,
    new_n18082_, new_n18083_, new_n18084_, new_n18085_, new_n18086_,
    new_n18087_, new_n18088_, new_n18089_, new_n18090_, new_n18091_,
    new_n18092_, new_n18093_, new_n18094_, new_n18095_, new_n18096_,
    new_n18097_, new_n18098_, new_n18099_, new_n18100_, new_n18101_,
    new_n18102_, new_n18103_, new_n18104_, new_n18105_, new_n18106_,
    new_n18107_, new_n18108_, new_n18109_, new_n18110_, new_n18111_,
    new_n18112_, new_n18113_, new_n18114_, new_n18115_, new_n18116_,
    new_n18117_, new_n18118_, new_n18119_, new_n18120_, new_n18121_,
    new_n18122_, new_n18123_, new_n18124_, new_n18125_, new_n18126_,
    new_n18127_, new_n18128_, new_n18129_, new_n18130_, new_n18131_,
    new_n18132_, new_n18133_, new_n18134_, new_n18135_, new_n18136_,
    new_n18137_, new_n18138_, new_n18139_, new_n18140_, new_n18141_,
    new_n18142_, new_n18143_, new_n18144_, new_n18145_, new_n18146_,
    new_n18147_, new_n18148_, new_n18149_, new_n18150_, new_n18151_,
    new_n18152_, new_n18153_, new_n18154_, new_n18155_, new_n18156_,
    new_n18157_, new_n18158_, new_n18159_, new_n18160_, new_n18161_,
    new_n18162_, new_n18163_, new_n18164_, new_n18165_, new_n18166_,
    new_n18167_, new_n18168_, new_n18169_, new_n18170_, new_n18171_,
    new_n18172_, new_n18173_, new_n18174_, new_n18175_, new_n18176_,
    new_n18177_, new_n18178_, new_n18179_, new_n18180_, new_n18181_,
    new_n18182_, new_n18183_, new_n18184_, new_n18185_, new_n18186_,
    new_n18187_, new_n18188_, new_n18189_, new_n18190_, new_n18191_,
    new_n18192_, new_n18193_, new_n18194_, new_n18195_, new_n18196_,
    new_n18197_, new_n18198_, new_n18199_, new_n18200_, new_n18201_,
    new_n18202_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18210_, new_n18211_,
    new_n18212_, new_n18213_, new_n18214_, new_n18215_, new_n18216_,
    new_n18217_, new_n18218_, new_n18219_, new_n18220_, new_n18221_,
    new_n18222_, new_n18223_, new_n18224_, new_n18225_, new_n18226_,
    new_n18227_, new_n18228_, new_n18229_, new_n18230_, new_n18231_,
    new_n18232_, new_n18233_, new_n18234_, new_n18235_, new_n18236_,
    new_n18237_, new_n18238_, new_n18239_, new_n18240_, new_n18241_,
    new_n18242_, new_n18243_, new_n18244_, new_n18245_, new_n18246_,
    new_n18247_, new_n18248_, new_n18249_, new_n18250_, new_n18251_,
    new_n18252_, new_n18253_, new_n18254_, new_n18255_, new_n18256_,
    new_n18257_, new_n18258_, new_n18259_, new_n18260_, new_n18261_,
    new_n18262_, new_n18263_, new_n18264_, new_n18265_, new_n18266_,
    new_n18267_, new_n18268_, new_n18269_, new_n18270_, new_n18271_,
    new_n18272_, new_n18273_, new_n18274_, new_n18275_, new_n18276_,
    new_n18277_, new_n18278_, new_n18279_, new_n18280_, new_n18281_,
    new_n18282_, new_n18283_, new_n18284_, new_n18285_, new_n18286_,
    new_n18287_, new_n18288_, new_n18289_, new_n18290_, new_n18291_,
    new_n18292_, new_n18293_, new_n18294_, new_n18295_, new_n18296_,
    new_n18297_, new_n18298_, new_n18299_, new_n18300_, new_n18301_,
    new_n18302_, new_n18303_, new_n18304_, new_n18305_, new_n18306_,
    new_n18307_, new_n18308_, new_n18309_, new_n18310_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18315_, new_n18316_,
    new_n18317_, new_n18318_, new_n18319_, new_n18320_, new_n18321_,
    new_n18322_, new_n18323_, new_n18324_, new_n18325_, new_n18326_,
    new_n18327_, new_n18328_, new_n18329_, new_n18330_, new_n18331_,
    new_n18332_, new_n18333_, new_n18334_, new_n18335_, new_n18336_,
    new_n18337_, new_n18338_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18577_, new_n18578_, new_n18579_, new_n18580_, new_n18581_,
    new_n18582_, new_n18583_, new_n18584_, new_n18585_, new_n18586_,
    new_n18587_, new_n18588_, new_n18589_, new_n18590_, new_n18591_,
    new_n18592_, new_n18593_, new_n18594_, new_n18595_, new_n18596_,
    new_n18597_, new_n18598_, new_n18599_, new_n18600_, new_n18601_,
    new_n18602_, new_n18603_, new_n18604_, new_n18605_, new_n18606_,
    new_n18607_, new_n18608_, new_n18609_, new_n18610_, new_n18611_,
    new_n18612_, new_n18613_, new_n18614_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18620_, new_n18621_,
    new_n18622_, new_n18623_, new_n18624_, new_n18625_, new_n18626_,
    new_n18627_, new_n18628_, new_n18629_, new_n18630_, new_n18631_,
    new_n18632_, new_n18633_, new_n18634_, new_n18635_, new_n18636_,
    new_n18637_, new_n18638_, new_n18639_, new_n18640_, new_n18641_,
    new_n18642_, new_n18643_, new_n18644_, new_n18645_, new_n18646_,
    new_n18647_, new_n18648_, new_n18649_, new_n18650_, new_n18651_,
    new_n18652_, new_n18653_, new_n18654_, new_n18655_, new_n18656_,
    new_n18657_, new_n18658_, new_n18659_, new_n18660_, new_n18661_,
    new_n18662_, new_n18663_, new_n18664_, new_n18665_, new_n18666_,
    new_n18667_, new_n18668_, new_n18669_, new_n18670_, new_n18671_,
    new_n18672_, new_n18673_, new_n18674_, new_n18675_, new_n18676_,
    new_n18677_, new_n18678_, new_n18679_, new_n18680_, new_n18681_,
    new_n18682_, new_n18683_, new_n18684_, new_n18685_, new_n18686_,
    new_n18687_, new_n18688_, new_n18689_, new_n18690_, new_n18691_,
    new_n18692_, new_n18693_, new_n18694_, new_n18695_, new_n18696_,
    new_n18697_, new_n18698_, new_n18699_, new_n18700_, new_n18701_,
    new_n18702_, new_n18703_, new_n18704_, new_n18705_, new_n18706_,
    new_n18707_, new_n18708_, new_n18709_, new_n18710_, new_n18711_,
    new_n18712_, new_n18713_, new_n18714_, new_n18715_, new_n18716_,
    new_n18717_, new_n18718_, new_n18719_, new_n18720_, new_n18721_,
    new_n18722_, new_n18723_, new_n18724_, new_n18725_, new_n18726_,
    new_n18727_, new_n18728_, new_n18729_, new_n18730_, new_n18731_,
    new_n18732_, new_n18733_, new_n18734_, new_n18735_, new_n18736_,
    new_n18737_, new_n18738_, new_n18739_, new_n18740_, new_n18741_,
    new_n18742_, new_n18743_, new_n18744_, new_n18745_, new_n18746_,
    new_n18747_, new_n18748_, new_n18749_, new_n18750_, new_n18751_,
    new_n18752_, new_n18753_, new_n18754_, new_n18755_, new_n18756_,
    new_n18757_, new_n18758_, new_n18759_, new_n18760_, new_n18761_,
    new_n18762_, new_n18763_, new_n18764_, new_n18765_, new_n18766_,
    new_n18767_, new_n18768_, new_n18769_, new_n18770_, new_n18771_,
    new_n18772_, new_n18773_, new_n18774_, new_n18775_, new_n18776_,
    new_n18777_, new_n18778_, new_n18779_, new_n18780_, new_n18781_,
    new_n18782_, new_n18783_, new_n18784_, new_n18785_, new_n18786_,
    new_n18787_, new_n18788_, new_n18789_, new_n18790_, new_n18791_,
    new_n18792_, new_n18793_, new_n18794_, new_n18795_, new_n18796_,
    new_n18797_, new_n18798_, new_n18799_, new_n18800_, new_n18801_,
    new_n18802_, new_n18803_, new_n18804_, new_n18805_, new_n18806_,
    new_n18807_, new_n18808_, new_n18809_, new_n18810_, new_n18811_,
    new_n18812_, new_n18813_, new_n18814_, new_n18815_, new_n18816_,
    new_n18817_, new_n18818_, new_n18819_, new_n18820_, new_n18821_,
    new_n18822_, new_n18823_, new_n18824_, new_n18825_, new_n18826_,
    new_n18827_, new_n18828_, new_n18829_, new_n18830_, new_n18831_,
    new_n18832_, new_n18833_, new_n18834_, new_n18835_, new_n18836_,
    new_n18837_, new_n18838_, new_n18839_, new_n18840_, new_n18841_,
    new_n18842_, new_n18843_, new_n18844_, new_n18845_, new_n18846_,
    new_n18847_, new_n18848_, new_n18849_, new_n18850_, new_n18851_,
    new_n18852_, new_n18853_, new_n18854_, new_n18855_, new_n18856_,
    new_n18857_, new_n18858_, new_n18859_, new_n18860_, new_n18861_,
    new_n18862_, new_n18863_, new_n18864_, new_n18865_, new_n18866_,
    new_n18867_, new_n18868_, new_n18869_, new_n18870_, new_n18871_,
    new_n18872_, new_n18873_, new_n18874_, new_n18875_, new_n18876_,
    new_n18877_, new_n18878_, new_n18879_, new_n18880_, new_n18881_,
    new_n18882_, new_n18883_, new_n18884_, new_n18885_, new_n18886_,
    new_n18887_, new_n18888_, new_n18889_, new_n18890_, new_n18891_,
    new_n18892_, new_n18893_, new_n18894_, new_n18895_, new_n18896_,
    new_n18897_, new_n18898_, new_n18899_, new_n18900_, new_n18901_,
    new_n18902_, new_n18903_, new_n18904_, new_n18905_, new_n18906_,
    new_n18907_, new_n18908_, new_n18909_, new_n18910_, new_n18911_,
    new_n18912_, new_n18913_, new_n18914_, new_n18915_, new_n18916_,
    new_n18917_, new_n18918_, new_n18919_, new_n18920_, new_n18921_,
    new_n18922_, new_n18923_, new_n18924_, new_n18925_, new_n18926_,
    new_n18927_, new_n18928_, new_n18929_, new_n18930_, new_n18931_,
    new_n18932_, new_n18933_, new_n18934_, new_n18935_, new_n18936_,
    new_n18937_, new_n18938_, new_n18939_, new_n18940_, new_n18941_,
    new_n18942_, new_n18943_, new_n18944_, new_n18945_, new_n18946_,
    new_n18947_, new_n18948_, new_n18949_, new_n18950_, new_n18951_,
    new_n18952_, new_n18953_, new_n18954_, new_n18955_, new_n18956_,
    new_n18957_, new_n18958_, new_n18959_, new_n18960_, new_n18961_,
    new_n18962_, new_n18963_, new_n18964_, new_n18965_, new_n18966_,
    new_n18967_, new_n18968_, new_n18969_, new_n18970_, new_n18971_,
    new_n18972_, new_n18973_, new_n18974_, new_n18975_, new_n18976_,
    new_n18977_, new_n18978_, new_n18979_, new_n18980_, new_n18981_,
    new_n18982_, new_n18983_, new_n18984_, new_n18985_, new_n18986_,
    new_n18987_, new_n18988_, new_n18989_, new_n18990_, new_n18991_,
    new_n18992_, new_n18993_, new_n18994_, new_n18995_, new_n18996_,
    new_n18997_, new_n18998_, new_n18999_, new_n19000_, new_n19001_,
    new_n19002_, new_n19003_, new_n19004_, new_n19005_, new_n19006_,
    new_n19007_, new_n19008_, new_n19009_, new_n19010_, new_n19011_,
    new_n19012_, new_n19013_, new_n19014_, new_n19015_, new_n19016_,
    new_n19017_, new_n19018_, new_n19019_, new_n19020_, new_n19021_,
    new_n19022_, new_n19023_, new_n19024_, new_n19025_, new_n19026_,
    new_n19027_, new_n19028_, new_n19029_, new_n19030_, new_n19031_,
    new_n19032_, new_n19033_, new_n19034_, new_n19035_, new_n19036_,
    new_n19037_, new_n19038_, new_n19039_, new_n19040_, new_n19041_,
    new_n19042_, new_n19043_, new_n19044_, new_n19045_, new_n19046_,
    new_n19047_, new_n19048_, new_n19049_, new_n19050_, new_n19051_,
    new_n19052_, new_n19053_, new_n19054_, new_n19055_, new_n19056_,
    new_n19057_, new_n19058_, new_n19059_, new_n19060_, new_n19061_,
    new_n19062_, new_n19063_, new_n19064_, new_n19065_, new_n19066_,
    new_n19067_, new_n19068_, new_n19069_, new_n19070_, new_n19071_,
    new_n19072_, new_n19073_, new_n19074_, new_n19075_, new_n19076_,
    new_n19077_, new_n19078_, new_n19079_, new_n19080_, new_n19081_,
    new_n19082_, new_n19083_, new_n19084_, new_n19085_, new_n19086_,
    new_n19087_, new_n19088_, new_n19089_, new_n19090_, new_n19091_,
    new_n19092_, new_n19093_, new_n19094_, new_n19095_, new_n19096_,
    new_n19097_, new_n19098_, new_n19099_, new_n19100_, new_n19101_,
    new_n19102_, new_n19103_, new_n19104_, new_n19105_, new_n19106_,
    new_n19107_, new_n19108_, new_n19109_, new_n19110_, new_n19111_,
    new_n19112_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19140_, new_n19141_,
    new_n19142_, new_n19143_, new_n19144_, new_n19145_, new_n19146_,
    new_n19147_, new_n19148_, new_n19149_, new_n19150_, new_n19151_,
    new_n19152_, new_n19153_, new_n19154_, new_n19155_, new_n19156_,
    new_n19157_, new_n19158_, new_n19159_, new_n19160_, new_n19161_,
    new_n19162_, new_n19163_, new_n19164_, new_n19165_, new_n19166_,
    new_n19167_, new_n19168_, new_n19169_, new_n19170_, new_n19171_,
    new_n19172_, new_n19173_, new_n19174_, new_n19175_, new_n19176_,
    new_n19177_, new_n19178_, new_n19179_, new_n19180_, new_n19181_,
    new_n19182_, new_n19183_, new_n19184_, new_n19185_, new_n19186_,
    new_n19187_, new_n19188_, new_n19189_, new_n19190_, new_n19191_,
    new_n19192_, new_n19193_, new_n19194_, new_n19195_, new_n19196_,
    new_n19197_, new_n19198_, new_n19199_, new_n19200_, new_n19201_,
    new_n19202_, new_n19203_, new_n19204_, new_n19205_, new_n19206_,
    new_n19207_, new_n19208_, new_n19209_, new_n19210_, new_n19211_,
    new_n19212_, new_n19213_, new_n19214_, new_n19215_, new_n19216_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19227_, new_n19228_, new_n19229_, new_n19230_, new_n19231_,
    new_n19232_, new_n19233_, new_n19234_, new_n19235_, new_n19236_,
    new_n19237_, new_n19238_, new_n19239_, new_n19240_, new_n19241_,
    new_n19242_, new_n19243_, new_n19244_, new_n19245_, new_n19246_,
    new_n19247_, new_n19248_, new_n19249_, new_n19250_, new_n19251_,
    new_n19252_, new_n19253_, new_n19254_, new_n19255_, new_n19256_,
    new_n19257_, new_n19258_, new_n19259_, new_n19260_, new_n19261_,
    new_n19262_, new_n19263_, new_n19264_, new_n19265_, new_n19266_,
    new_n19267_, new_n19268_, new_n19269_, new_n19270_, new_n19271_,
    new_n19272_, new_n19273_, new_n19274_, new_n19275_, new_n19276_,
    new_n19277_, new_n19278_, new_n19279_, new_n19280_, new_n19281_,
    new_n19282_, new_n19283_, new_n19284_, new_n19285_, new_n19286_,
    new_n19287_, new_n19288_, new_n19289_, new_n19290_, new_n19291_,
    new_n19292_, new_n19293_, new_n19294_, new_n19295_, new_n19296_,
    new_n19297_, new_n19298_, new_n19299_, new_n19300_, new_n19301_,
    new_n19302_, new_n19303_, new_n19304_, new_n19305_, new_n19306_,
    new_n19307_, new_n19308_, new_n19309_, new_n19310_, new_n19311_,
    new_n19312_, new_n19313_, new_n19314_, new_n19315_, new_n19316_,
    new_n19317_, new_n19318_, new_n19319_, new_n19320_, new_n19321_,
    new_n19322_, new_n19323_, new_n19324_, new_n19325_, new_n19326_,
    new_n19327_, new_n19328_, new_n19329_, new_n19330_, new_n19331_,
    new_n19332_, new_n19333_, new_n19334_, new_n19335_, new_n19336_,
    new_n19337_, new_n19338_, new_n19339_, new_n19340_, new_n19341_,
    new_n19342_, new_n19343_, new_n19344_, new_n19345_, new_n19346_,
    new_n19347_, new_n19348_, new_n19349_, new_n19350_, new_n19351_,
    new_n19352_, new_n19353_, new_n19354_, new_n19355_, new_n19356_,
    new_n19357_, new_n19358_, new_n19359_, new_n19360_, new_n19361_,
    new_n19362_, new_n19363_, new_n19364_, new_n19365_, new_n19366_,
    new_n19367_, new_n19368_, new_n19369_, new_n19370_, new_n19371_,
    new_n19372_, new_n19373_, new_n19374_, new_n19375_, new_n19376_,
    new_n19377_, new_n19378_, new_n19379_, new_n19380_, new_n19381_,
    new_n19382_, new_n19383_, new_n19384_, new_n19385_, new_n19386_,
    new_n19387_, new_n19388_, new_n19389_, new_n19390_, new_n19391_,
    new_n19392_, new_n19393_, new_n19394_, new_n19395_, new_n19396_,
    new_n19397_, new_n19398_, new_n19399_, new_n19400_, new_n19401_,
    new_n19402_, new_n19403_, new_n19404_, new_n19405_, new_n19406_,
    new_n19407_, new_n19408_, new_n19409_, new_n19410_, new_n19411_,
    new_n19412_, new_n19413_, new_n19414_, new_n19415_, new_n19416_,
    new_n19417_, new_n19418_, new_n19419_, new_n19420_, new_n19421_,
    new_n19422_, new_n19423_, new_n19424_, new_n19425_, new_n19426_,
    new_n19427_, new_n19428_, new_n19429_, new_n19430_, new_n19431_,
    new_n19432_, new_n19433_, new_n19434_, new_n19435_, new_n19436_,
    new_n19437_, new_n19438_, new_n19439_, new_n19440_, new_n19441_,
    new_n19442_, new_n19443_, new_n19444_, new_n19445_, new_n19446_,
    new_n19447_, new_n19448_, new_n19449_, new_n19450_, new_n19451_,
    new_n19452_, new_n19453_, new_n19454_, new_n19455_, new_n19456_,
    new_n19457_, new_n19458_, new_n19459_, new_n19460_, new_n19461_,
    new_n19462_, new_n19463_, new_n19464_, new_n19465_, new_n19466_,
    new_n19467_, new_n19468_, new_n19469_, new_n19470_, new_n19471_,
    new_n19472_, new_n19473_, new_n19474_, new_n19475_, new_n19476_,
    new_n19477_, new_n19478_, new_n19479_, new_n19480_, new_n19481_,
    new_n19482_, new_n19483_, new_n19484_, new_n19485_, new_n19486_,
    new_n19487_, new_n19488_, new_n19489_, new_n19490_, new_n19491_,
    new_n19492_, new_n19493_, new_n19494_, new_n19495_, new_n19496_,
    new_n19497_, new_n19498_, new_n19499_, new_n19500_, new_n19501_,
    new_n19502_, new_n19503_, new_n19504_, new_n19505_, new_n19506_,
    new_n19507_, new_n19508_, new_n19509_, new_n19510_, new_n19511_,
    new_n19512_, new_n19513_, new_n19514_, new_n19515_, new_n19516_,
    new_n19517_, new_n19518_, new_n19519_, new_n19520_, new_n19521_,
    new_n19522_, new_n19523_, new_n19524_, new_n19525_, new_n19526_,
    new_n19527_, new_n19528_, new_n19529_, new_n19530_, new_n19531_,
    new_n19532_, new_n19533_, new_n19534_, new_n19535_, new_n19536_,
    new_n19537_, new_n19538_, new_n19539_, new_n19540_, new_n19541_,
    new_n19542_, new_n19543_, new_n19544_, new_n19545_, new_n19546_,
    new_n19547_, new_n19548_, new_n19549_, new_n19550_, new_n19551_,
    new_n19552_, new_n19553_, new_n19554_, new_n19555_, new_n19556_,
    new_n19557_, new_n19558_, new_n19559_, new_n19560_, new_n19561_,
    new_n19562_, new_n19563_, new_n19564_, new_n19565_, new_n19566_,
    new_n19567_, new_n19568_, new_n19569_, new_n19570_, new_n19571_,
    new_n19572_, new_n19573_, new_n19574_, new_n19575_, new_n19576_,
    new_n19577_, new_n19578_, new_n19579_, new_n19580_, new_n19581_,
    new_n19582_, new_n19583_, new_n19584_, new_n19585_, new_n19586_,
    new_n19587_, new_n19588_, new_n19589_, new_n19590_, new_n19591_,
    new_n19592_, new_n19593_, new_n19594_, new_n19595_, new_n19596_,
    new_n19597_, new_n19598_, new_n19599_, new_n19600_, new_n19601_,
    new_n19602_, new_n19603_, new_n19604_, new_n19605_, new_n19606_,
    new_n19607_, new_n19608_, new_n19609_, new_n19610_, new_n19611_,
    new_n19612_, new_n19613_, new_n19614_, new_n19615_, new_n19616_,
    new_n19617_, new_n19618_, new_n19619_, new_n19620_, new_n19621_,
    new_n19622_, new_n19623_, new_n19624_, new_n19625_, new_n19626_,
    new_n19627_, new_n19628_, new_n19629_, new_n19630_, new_n19631_,
    new_n19632_, new_n19633_, new_n19634_, new_n19635_, new_n19636_,
    new_n19637_, new_n19638_, new_n19639_, new_n19640_, new_n19641_,
    new_n19642_, new_n19643_, new_n19644_, new_n19645_, new_n19646_,
    new_n19647_, new_n19648_, new_n19649_, new_n19650_, new_n19651_,
    new_n19652_, new_n19653_, new_n19654_, new_n19655_, new_n19656_,
    new_n19657_, new_n19658_, new_n19659_, new_n19660_, new_n19661_,
    new_n19662_, new_n19663_, new_n19664_, new_n19665_, new_n19666_,
    new_n19667_, new_n19668_, new_n19669_, new_n19670_, new_n19671_,
    new_n19672_, new_n19673_, new_n19674_, new_n19675_, new_n19676_,
    new_n19677_, new_n19678_, new_n19679_, new_n19680_, new_n19681_,
    new_n19682_, new_n19683_, new_n19684_, new_n19685_, new_n19686_,
    new_n19687_, new_n19688_, new_n19689_, new_n19690_, new_n19691_,
    new_n19692_, new_n19693_, new_n19694_, new_n19695_, new_n19696_,
    new_n19697_, new_n19698_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20321_,
    new_n20322_, new_n20323_, new_n20324_, new_n20325_, new_n20326_,
    new_n20327_, new_n20328_, new_n20329_, new_n20330_, new_n20331_,
    new_n20332_, new_n20333_, new_n20334_, new_n20335_, new_n20336_,
    new_n20337_, new_n20338_, new_n20339_, new_n20340_, new_n20341_,
    new_n20342_, new_n20343_, new_n20344_, new_n20345_, new_n20346_,
    new_n20347_, new_n20348_, new_n20349_, new_n20350_, new_n20351_,
    new_n20352_, new_n20353_, new_n20354_, new_n20355_, new_n20356_,
    new_n20357_, new_n20358_, new_n20359_, new_n20360_, new_n20361_,
    new_n20362_, new_n20363_, new_n20364_, new_n20365_, new_n20366_,
    new_n20367_, new_n20368_, new_n20369_, new_n20370_, new_n20371_,
    new_n20372_, new_n20373_, new_n20374_, new_n20375_, new_n20376_,
    new_n20377_, new_n20378_, new_n20379_, new_n20380_, new_n20381_,
    new_n20382_, new_n20383_, new_n20384_, new_n20385_, new_n20386_,
    new_n20387_, new_n20388_, new_n20389_, new_n20390_, new_n20391_,
    new_n20392_, new_n20393_, new_n20394_, new_n20395_, new_n20396_,
    new_n20397_, new_n20398_, new_n20399_, new_n20400_, new_n20401_,
    new_n20402_, new_n20403_, new_n20404_, new_n20405_, new_n20406_,
    new_n20407_, new_n20408_, new_n20409_, new_n20410_, new_n20411_,
    new_n20412_, new_n20413_, new_n20414_, new_n20415_, new_n20416_,
    new_n20417_, new_n20418_, new_n20419_, new_n20420_, new_n20421_,
    new_n20422_, new_n20423_, new_n20424_, new_n20425_, new_n20426_,
    new_n20427_, new_n20428_, new_n20429_, new_n20430_, new_n20431_,
    new_n20432_, new_n20433_, new_n20434_, new_n20435_, new_n20436_,
    new_n20437_, new_n20438_, new_n20439_, new_n20440_, new_n20441_,
    new_n20442_, new_n20443_, new_n20444_, new_n20445_, new_n20446_,
    new_n20447_, new_n20448_, new_n20449_, new_n20450_, new_n20451_,
    new_n20452_, new_n20453_, new_n20454_, new_n20455_, new_n20456_,
    new_n20457_, new_n20458_, new_n20459_, new_n20460_, new_n20461_,
    new_n20462_, new_n20463_, new_n20464_, new_n20465_, new_n20466_,
    new_n20467_, new_n20468_, new_n20469_, new_n20470_, new_n20471_,
    new_n20472_, new_n20473_, new_n20474_, new_n20475_, new_n20476_,
    new_n20477_, new_n20478_, new_n20479_, new_n20480_, new_n20481_,
    new_n20482_, new_n20483_, new_n20484_, new_n20485_, new_n20486_,
    new_n20487_, new_n20488_, new_n20489_, new_n20490_, new_n20491_,
    new_n20492_, new_n20493_, new_n20494_, new_n20495_, new_n20496_,
    new_n20497_, new_n20498_, new_n20499_, new_n20500_, new_n20501_,
    new_n20502_, new_n20503_, new_n20504_, new_n20505_, new_n20506_,
    new_n20507_, new_n20508_, new_n20509_, new_n20510_, new_n20511_,
    new_n20512_, new_n20513_, new_n20514_, new_n20515_, new_n20516_,
    new_n20517_, new_n20518_, new_n20519_, new_n20520_, new_n20521_,
    new_n20522_, new_n20523_, new_n20524_, new_n20525_, new_n20526_,
    new_n20527_, new_n20528_, new_n20529_, new_n20530_, new_n20531_,
    new_n20532_, new_n20533_, new_n20534_, new_n20535_, new_n20536_,
    new_n20537_, new_n20538_, new_n20539_, new_n20540_, new_n20541_,
    new_n20542_, new_n20543_, new_n20544_, new_n20545_, new_n20546_,
    new_n20547_, new_n20548_, new_n20549_, new_n20550_, new_n20551_,
    new_n20552_, new_n20553_, new_n20554_, new_n20555_, new_n20556_,
    new_n20557_, new_n20558_, new_n20559_, new_n20560_, new_n20561_,
    new_n20562_, new_n20563_, new_n20564_, new_n20565_, new_n20566_,
    new_n20567_, new_n20568_, new_n20569_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20679_, new_n20680_, new_n20681_,
    new_n20682_, new_n20683_, new_n20684_, new_n20685_, new_n20686_,
    new_n20687_, new_n20688_, new_n20689_, new_n20690_, new_n20691_,
    new_n20692_, new_n20693_, new_n20694_, new_n20695_, new_n20696_,
    new_n20697_, new_n20698_, new_n20699_, new_n20700_, new_n20701_,
    new_n20702_, new_n20703_, new_n20704_, new_n20705_, new_n20706_,
    new_n20707_, new_n20708_, new_n20709_, new_n20710_, new_n20711_,
    new_n20712_, new_n20713_, new_n20714_, new_n20715_, new_n20716_,
    new_n20717_, new_n20718_, new_n20719_, new_n20720_, new_n20721_,
    new_n20722_, new_n20723_, new_n20724_, new_n20725_, new_n20726_,
    new_n20727_, new_n20728_, new_n20729_, new_n20730_, new_n20731_,
    new_n20732_, new_n20733_, new_n20734_, new_n20735_, new_n20736_,
    new_n20737_, new_n20738_, new_n20739_, new_n20740_, new_n20741_,
    new_n20742_, new_n20743_, new_n20744_, new_n20745_, new_n20746_,
    new_n20747_, new_n20748_, new_n20749_, new_n20750_, new_n20751_,
    new_n20752_, new_n20753_, new_n20754_, new_n20755_, new_n20756_,
    new_n20757_, new_n20758_, new_n20759_, new_n20760_, new_n20761_,
    new_n20762_, new_n20763_, new_n20764_, new_n20765_, new_n20766_,
    new_n20767_, new_n20768_, new_n20769_, new_n20770_, new_n20771_,
    new_n20772_, new_n20773_, new_n20774_, new_n20775_, new_n20776_,
    new_n20777_, new_n20778_, new_n20779_, new_n20780_, new_n20781_,
    new_n20782_, new_n20783_, new_n20784_, new_n20785_, new_n20786_,
    new_n20787_, new_n20788_, new_n20789_, new_n20790_, new_n20791_,
    new_n20792_, new_n20793_, new_n20794_, new_n20795_, new_n20796_,
    new_n20797_, new_n20798_, new_n20799_, new_n20800_, new_n20801_,
    new_n20802_, new_n20803_, new_n20804_, new_n20805_, new_n20806_,
    new_n20807_, new_n20808_, new_n20809_, new_n20810_, new_n20811_,
    new_n20812_, new_n20813_, new_n20814_, new_n20815_, new_n20816_,
    new_n20817_, new_n20818_, new_n20819_, new_n20820_, new_n20821_,
    new_n20822_, new_n20823_, new_n20824_, new_n20825_, new_n20826_,
    new_n20827_, new_n20828_, new_n20829_, new_n20830_, new_n20831_,
    new_n20832_, new_n20833_, new_n20834_, new_n20835_, new_n20836_,
    new_n20837_, new_n20838_, new_n20839_, new_n20840_, new_n20841_,
    new_n20842_, new_n20843_, new_n20844_, new_n20845_, new_n20846_,
    new_n20847_, new_n20848_, new_n20849_, new_n20850_, new_n20851_,
    new_n20852_, new_n20853_, new_n20854_, new_n20855_, new_n20856_,
    new_n20857_, new_n20858_, new_n20859_, new_n20860_, new_n20861_,
    new_n20862_, new_n20863_, new_n20864_, new_n20865_, new_n20866_,
    new_n20867_, new_n20868_, new_n20869_, new_n20870_, new_n20871_,
    new_n20872_, new_n20873_, new_n20874_, new_n20875_, new_n20876_,
    new_n20877_, new_n20878_, new_n20879_, new_n20880_, new_n20881_,
    new_n20882_, new_n20883_, new_n20884_, new_n20885_, new_n20886_,
    new_n20887_, new_n20888_, new_n20889_, new_n20890_, new_n20891_,
    new_n20892_, new_n20893_, new_n20894_, new_n20895_, new_n20896_,
    new_n20897_, new_n20898_, new_n20899_, new_n20900_, new_n20901_,
    new_n20902_, new_n20903_, new_n20904_, new_n20905_, new_n20906_,
    new_n20907_, new_n20908_, new_n20909_, new_n20910_, new_n20911_,
    new_n20912_, new_n20913_, new_n20914_, new_n20915_, new_n20916_,
    new_n20917_, new_n20918_, new_n20919_, new_n20920_, new_n20921_,
    new_n20922_, new_n20923_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20969_, new_n20970_, new_n20971_,
    new_n20972_, new_n20973_, new_n20974_, new_n20975_, new_n20976_,
    new_n20977_, new_n20978_, new_n20979_, new_n20980_, new_n20981_,
    new_n20982_, new_n20983_, new_n20984_, new_n20985_, new_n20986_,
    new_n20987_, new_n20988_, new_n20989_, new_n20990_, new_n20991_,
    new_n20992_, new_n20993_, new_n20994_, new_n20995_, new_n20996_,
    new_n20997_, new_n20998_, new_n20999_, new_n21000_, new_n21001_,
    new_n21002_, new_n21003_, new_n21004_, new_n21005_, new_n21006_,
    new_n21007_, new_n21008_, new_n21009_, new_n21010_, new_n21011_,
    new_n21012_, new_n21013_, new_n21014_, new_n21015_, new_n21016_,
    new_n21017_, new_n21018_, new_n21019_, new_n21020_, new_n21021_,
    new_n21022_, new_n21023_, new_n21024_, new_n21025_, new_n21026_,
    new_n21027_, new_n21028_, new_n21029_, new_n21030_, new_n21031_,
    new_n21032_, new_n21033_, new_n21034_, new_n21035_, new_n21036_,
    new_n21037_, new_n21038_, new_n21039_, new_n21040_, new_n21041_,
    new_n21042_, new_n21043_, new_n21044_, new_n21045_, new_n21046_,
    new_n21047_, new_n21048_, new_n21049_, new_n21050_, new_n21051_,
    new_n21052_, new_n21053_, new_n21054_, new_n21055_, new_n21056_,
    new_n21057_, new_n21058_, new_n21059_, new_n21060_, new_n21061_,
    new_n21062_, new_n21063_, new_n21064_, new_n21065_, new_n21066_,
    new_n21067_, new_n21068_, new_n21069_, new_n21070_, new_n21071_,
    new_n21072_, new_n21073_, new_n21074_, new_n21075_, new_n21076_,
    new_n21077_, new_n21078_, new_n21079_, new_n21080_, new_n21081_,
    new_n21082_, new_n21083_, new_n21084_, new_n21085_, new_n21086_,
    new_n21087_, new_n21088_, new_n21089_, new_n21090_, new_n21091_,
    new_n21092_, new_n21093_, new_n21094_, new_n21095_, new_n21096_,
    new_n21097_, new_n21098_, new_n21099_, new_n21100_, new_n21101_,
    new_n21102_, new_n21103_, new_n21104_, new_n21105_, new_n21106_,
    new_n21107_, new_n21108_, new_n21109_, new_n21110_, new_n21111_,
    new_n21112_, new_n21113_, new_n21114_, new_n21115_, new_n21116_,
    new_n21117_, new_n21118_, new_n21119_, new_n21120_, new_n21121_,
    new_n21122_, new_n21123_, new_n21124_, new_n21125_, new_n21126_,
    new_n21127_, new_n21128_, new_n21129_, new_n21130_, new_n21131_,
    new_n21132_, new_n21133_, new_n21134_, new_n21135_, new_n21136_,
    new_n21137_, new_n21138_, new_n21139_, new_n21140_, new_n21141_,
    new_n21142_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21178_, new_n21179_, new_n21180_, new_n21181_,
    new_n21182_, new_n21183_, new_n21184_, new_n21185_, new_n21186_,
    new_n21187_, new_n21188_, new_n21189_, new_n21190_, new_n21191_,
    new_n21192_, new_n21193_, new_n21194_, new_n21195_, new_n21196_,
    new_n21197_, new_n21198_, new_n21199_, new_n21200_, new_n21201_,
    new_n21202_, new_n21203_, new_n21204_, new_n21205_, new_n21206_,
    new_n21207_, new_n21208_, new_n21209_, new_n21210_, new_n21211_,
    new_n21212_, new_n21213_, new_n21214_, new_n21215_, new_n21216_,
    new_n21217_, new_n21218_, new_n21219_, new_n21220_, new_n21221_,
    new_n21222_, new_n21223_, new_n21224_, new_n21225_, new_n21226_,
    new_n21227_, new_n21228_, new_n21229_, new_n21230_, new_n21231_,
    new_n21232_, new_n21233_, new_n21234_, new_n21235_, new_n21236_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21385_, new_n21386_,
    new_n21387_, new_n21388_, new_n21389_, new_n21390_, new_n21391_,
    new_n21392_, new_n21393_, new_n21394_, new_n21395_, new_n21396_,
    new_n21397_, new_n21398_, new_n21399_, new_n21400_, new_n21401_,
    new_n21402_, new_n21403_, new_n21404_, new_n21405_, new_n21406_,
    new_n21407_, new_n21408_, new_n21409_, new_n21410_, new_n21411_,
    new_n21412_, new_n21413_, new_n21414_, new_n21415_, new_n21416_,
    new_n21417_, new_n21418_, new_n21419_, new_n21420_, new_n21421_,
    new_n21422_, new_n21423_, new_n21424_, new_n21425_, new_n21426_,
    new_n21427_, new_n21428_, new_n21429_, new_n21430_, new_n21431_,
    new_n21432_, new_n21433_, new_n21434_, new_n21435_, new_n21436_,
    new_n21437_, new_n21438_, new_n21439_, new_n21440_, new_n21441_,
    new_n21442_, new_n21443_, new_n21444_, new_n21445_, new_n21446_,
    new_n21447_, new_n21448_, new_n21449_, new_n21450_, new_n21451_,
    new_n21452_, new_n21453_, new_n21454_, new_n21455_, new_n21456_,
    new_n21457_, new_n21458_, new_n21459_, new_n21460_, new_n21461_,
    new_n21462_, new_n21463_, new_n21464_, new_n21465_, new_n21466_,
    new_n21467_, new_n21468_, new_n21469_, new_n21470_, new_n21471_,
    new_n21472_, new_n21473_, new_n21474_, new_n21475_, new_n21476_,
    new_n21477_, new_n21478_, new_n21479_, new_n21480_, new_n21481_,
    new_n21482_, new_n21483_, new_n21484_, new_n21485_, new_n21486_,
    new_n21487_, new_n21488_, new_n21489_, new_n21490_, new_n21491_,
    new_n21492_, new_n21493_, new_n21494_, new_n21495_, new_n21496_,
    new_n21497_, new_n21498_, new_n21499_, new_n21500_, new_n21501_,
    new_n21502_, new_n21503_, new_n21504_, new_n21505_, new_n21506_,
    new_n21507_, new_n21508_, new_n21509_, new_n21510_, new_n21511_,
    new_n21512_, new_n21513_, new_n21514_, new_n21515_, new_n21516_,
    new_n21517_, new_n21518_, new_n21519_, new_n21520_, new_n21521_,
    new_n21522_, new_n21523_, new_n21524_, new_n21525_, new_n21526_,
    new_n21527_, new_n21528_, new_n21529_, new_n21530_, new_n21531_,
    new_n21532_, new_n21533_, new_n21534_, new_n21535_, new_n21536_,
    new_n21537_, new_n21538_, new_n21539_, new_n21540_, new_n21541_,
    new_n21542_, new_n21543_, new_n21544_, new_n21545_, new_n21546_,
    new_n21547_, new_n21548_, new_n21549_, new_n21550_, new_n21551_,
    new_n21552_, new_n21553_, new_n21554_, new_n21555_, new_n21556_,
    new_n21557_, new_n21558_, new_n21559_, new_n21560_, new_n21561_,
    new_n21562_, new_n21563_, new_n21564_, new_n21565_, new_n21566_,
    new_n21567_, new_n21568_, new_n21569_, new_n21570_, new_n21571_,
    new_n21572_, new_n21573_, new_n21574_, new_n21575_, new_n21576_,
    new_n21577_, new_n21578_, new_n21579_, new_n21580_, new_n21581_,
    new_n21582_, new_n21583_, new_n21584_, new_n21585_, new_n21586_,
    new_n21587_, new_n21588_, new_n21589_, new_n21590_, new_n21591_,
    new_n21592_, new_n21593_, new_n21594_, new_n21595_, new_n21596_,
    new_n21597_, new_n21598_, new_n21599_, new_n21600_, new_n21601_,
    new_n21602_, new_n21603_, new_n21604_, new_n21605_, new_n21606_,
    new_n21607_, new_n21608_, new_n21609_, new_n21610_, new_n21611_,
    new_n21612_, new_n21613_, new_n21614_, new_n21615_, new_n21616_,
    new_n21617_, new_n21618_, new_n21619_, new_n21620_, new_n21621_,
    new_n21622_, new_n21623_, new_n21624_, new_n21625_, new_n21626_,
    new_n21627_, new_n21628_, new_n21629_, new_n21630_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21691_,
    new_n21692_, new_n21693_, new_n21694_, new_n21695_, new_n21696_,
    new_n21697_, new_n21698_, new_n21699_, new_n21700_, new_n21701_,
    new_n21702_, new_n21703_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21776_,
    new_n21777_, new_n21778_, new_n21779_, new_n21780_, new_n21781_,
    new_n21782_, new_n21783_, new_n21784_, new_n21785_, new_n21786_,
    new_n21787_, new_n21788_, new_n21789_, new_n21790_, new_n21791_,
    new_n21792_, new_n21793_, new_n21794_, new_n21795_, new_n21796_,
    new_n21797_, new_n21798_, new_n21799_, new_n21800_, new_n21801_,
    new_n21802_, new_n21803_, new_n21804_, new_n21805_, new_n21806_,
    new_n21807_, new_n21808_, new_n21809_, new_n21810_, new_n21811_,
    new_n21812_, new_n21813_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21880_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22304_, new_n22305_, new_n22306_,
    new_n22307_, new_n22308_, new_n22309_, new_n22310_, new_n22311_,
    new_n22312_, new_n22313_, new_n22314_, new_n22315_, new_n22316_,
    new_n22317_, new_n22318_, new_n22319_, new_n22320_, new_n22321_,
    new_n22322_, new_n22323_, new_n22324_, new_n22325_, new_n22326_,
    new_n22327_, new_n22328_, new_n22329_, new_n22330_, new_n22331_,
    new_n22332_, new_n22333_, new_n22334_, new_n22335_, new_n22336_,
    new_n22337_, new_n22338_, new_n22339_, new_n22340_, new_n22341_,
    new_n22342_, new_n22343_, new_n22344_, new_n22345_, new_n22346_,
    new_n22347_, new_n22348_, new_n22349_, new_n22350_, new_n22351_,
    new_n22352_, new_n22353_, new_n22354_, new_n22355_, new_n22356_,
    new_n22357_, new_n22358_, new_n22359_, new_n22360_, new_n22361_,
    new_n22362_, new_n22363_, new_n22364_, new_n22365_, new_n22366_,
    new_n22367_, new_n22368_, new_n22369_, new_n22370_, new_n22371_,
    new_n22372_, new_n22373_, new_n22374_, new_n22375_, new_n22376_,
    new_n22377_, new_n22378_, new_n22379_, new_n22380_, new_n22381_,
    new_n22382_, new_n22383_, new_n22384_, new_n22385_, new_n22386_,
    new_n22387_, new_n22388_, new_n22389_, new_n22390_, new_n22391_,
    new_n22392_, new_n22393_, new_n22394_, new_n22395_, new_n22396_,
    new_n22397_, new_n22398_, new_n22399_, new_n22400_, new_n22401_,
    new_n22402_, new_n22403_, new_n22404_, new_n22405_, new_n22406_,
    new_n22407_, new_n22408_, new_n22409_, new_n22410_, new_n22411_,
    new_n22412_, new_n22413_, new_n22414_, new_n22415_, new_n22416_,
    new_n22417_, new_n22418_, new_n22419_, new_n22420_, new_n22421_,
    new_n22422_, new_n22423_, new_n22424_, new_n22425_, new_n22426_,
    new_n22427_, new_n22428_, new_n22429_, new_n22430_, new_n22431_,
    new_n22432_, new_n22433_, new_n22434_, new_n22435_, new_n22436_,
    new_n22437_, new_n22438_, new_n22439_, new_n22440_, new_n22441_,
    new_n22442_, new_n22443_, new_n22444_, new_n22445_, new_n22446_,
    new_n22447_, new_n22448_, new_n22449_, new_n22450_, new_n22451_,
    new_n22452_, new_n22453_, new_n22454_, new_n22455_, new_n22456_,
    new_n22457_, new_n22458_, new_n22459_, new_n22460_, new_n22461_,
    new_n22462_, new_n22463_, new_n22464_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22471_,
    new_n22472_, new_n22473_, new_n22474_, new_n22475_, new_n22476_,
    new_n22477_, new_n22478_, new_n22479_, new_n22480_, new_n22481_,
    new_n22482_, new_n22483_, new_n22484_, new_n22485_, new_n22486_,
    new_n22487_, new_n22488_, new_n22489_, new_n22490_, new_n22491_,
    new_n22492_, new_n22493_, new_n22494_, new_n22495_, new_n22496_,
    new_n22497_, new_n22498_, new_n22499_, new_n22500_, new_n22501_,
    new_n22502_, new_n22503_, new_n22504_, new_n22505_, new_n22506_,
    new_n22507_, new_n22508_, new_n22509_, new_n22510_, new_n22511_,
    new_n22512_, new_n22513_, new_n22514_, new_n22515_, new_n22516_,
    new_n22517_, new_n22518_, new_n22519_, new_n22520_, new_n22521_,
    new_n22522_, new_n22523_, new_n22524_, new_n22525_, new_n22526_,
    new_n22527_, new_n22528_, new_n22529_, new_n22530_, new_n22531_,
    new_n22532_, new_n22533_, new_n22534_, new_n22535_, new_n22536_,
    new_n22537_, new_n22538_, new_n22539_, new_n22540_, new_n22541_,
    new_n22542_, new_n22543_, new_n22544_, new_n22545_, new_n22546_,
    new_n22547_, new_n22548_, new_n22549_, new_n22550_, new_n22551_,
    new_n22552_, new_n22553_, new_n22554_, new_n22555_, new_n22556_,
    new_n22557_, new_n22558_, new_n22559_, new_n22560_, new_n22561_,
    new_n22562_, new_n22563_, new_n22564_, new_n22565_, new_n22566_,
    new_n22567_, new_n22568_, new_n22569_, new_n22570_, new_n22571_,
    new_n22572_, new_n22573_, new_n22574_, new_n22575_, new_n22576_,
    new_n22577_, new_n22578_, new_n22579_, new_n22580_, new_n22581_,
    new_n22582_, new_n22583_, new_n22584_, new_n22585_, new_n22586_,
    new_n22587_, new_n22588_, new_n22589_, new_n22590_, new_n22591_,
    new_n22592_, new_n22593_, new_n22594_, new_n22595_, new_n22596_,
    new_n22597_, new_n22598_, new_n22599_, new_n22600_, new_n22601_,
    new_n22602_, new_n22603_, new_n22604_, new_n22605_, new_n22606_,
    new_n22607_, new_n22608_, new_n22609_, new_n22610_, new_n22611_,
    new_n22612_, new_n22613_, new_n22614_, new_n22615_, new_n22616_,
    new_n22617_, new_n22618_, new_n22619_, new_n22620_, new_n22621_,
    new_n22622_, new_n22623_, new_n22624_, new_n22625_, new_n22626_,
    new_n22627_, new_n22628_, new_n22629_, new_n22630_, new_n22631_,
    new_n22632_, new_n22633_, new_n22634_, new_n22635_, new_n22636_,
    new_n22637_, new_n22638_, new_n22639_, new_n22640_, new_n22641_,
    new_n22642_, new_n22643_, new_n22644_, new_n22645_, new_n22646_,
    new_n22647_, new_n22648_, new_n22649_, new_n22650_, new_n22651_,
    new_n22652_, new_n22653_, new_n22654_, new_n22655_, new_n22656_,
    new_n22657_, new_n22658_, new_n22659_, new_n22660_, new_n22661_,
    new_n22662_, new_n22663_, new_n22664_, new_n22665_, new_n22666_,
    new_n22667_, new_n22668_, new_n22669_, new_n22670_, new_n22671_,
    new_n22672_, new_n22673_, new_n22674_, new_n22675_, new_n22676_,
    new_n22677_, new_n22678_, new_n22679_, new_n22680_, new_n22681_,
    new_n22682_, new_n22683_, new_n22684_, new_n22685_, new_n22686_,
    new_n22687_, new_n22688_, new_n22689_, new_n22690_, new_n22691_,
    new_n22692_, new_n22693_, new_n22694_, new_n22695_, new_n22696_,
    new_n22697_, new_n22698_, new_n22699_, new_n22700_, new_n22701_,
    new_n22702_, new_n22703_, new_n22704_, new_n22705_, new_n22706_,
    new_n22707_, new_n22708_, new_n22709_, new_n22710_, new_n22711_,
    new_n22712_, new_n22713_, new_n22714_, new_n22715_, new_n22716_,
    new_n22717_, new_n22718_, new_n22719_, new_n22720_, new_n22721_,
    new_n22722_, new_n22723_, new_n22724_, new_n22725_, new_n22726_,
    new_n22727_, new_n22728_, new_n22729_, new_n22730_, new_n22731_,
    new_n22732_, new_n22733_, new_n22734_, new_n22735_, new_n22736_,
    new_n22737_, new_n22738_, new_n22739_, new_n22740_, new_n22741_,
    new_n22742_, new_n22743_, new_n22744_, new_n22745_, new_n22746_,
    new_n22747_, new_n22748_, new_n22749_, new_n22750_, new_n22751_,
    new_n22752_, new_n22753_, new_n22754_, new_n22755_, new_n22756_,
    new_n22757_, new_n22758_, new_n22759_, new_n22760_, new_n22761_,
    new_n22762_, new_n22763_, new_n22764_, new_n22765_, new_n22766_,
    new_n22767_, new_n22768_, new_n22769_, new_n22770_, new_n22771_,
    new_n22772_, new_n22773_, new_n22774_, new_n22775_, new_n22776_,
    new_n22777_, new_n22778_, new_n22779_, new_n22780_, new_n22781_,
    new_n22782_, new_n22783_, new_n22784_, new_n22785_, new_n22786_,
    new_n22787_, new_n22788_, new_n22789_, new_n22790_, new_n22791_,
    new_n22792_, new_n22793_, new_n22794_, new_n22795_, new_n22796_,
    new_n22797_, new_n22798_, new_n22799_, new_n22800_, new_n22801_,
    new_n22802_, new_n22803_, new_n22804_, new_n22805_, new_n22806_,
    new_n22807_, new_n22808_, new_n22809_, new_n22810_, new_n22811_,
    new_n22812_, new_n22813_, new_n22814_, new_n22815_, new_n22816_,
    new_n22817_, new_n22818_, new_n22819_, new_n22820_, new_n22821_,
    new_n22822_, new_n22823_, new_n22824_, new_n22825_, new_n22826_,
    new_n22827_, new_n22828_, new_n22829_, new_n22830_, new_n22831_,
    new_n22832_, new_n22833_, new_n22834_, new_n22835_, new_n22836_,
    new_n22837_, new_n22838_, new_n22839_, new_n22840_, new_n22841_,
    new_n22842_, new_n22843_, new_n22844_, new_n22845_, new_n22846_,
    new_n22847_, new_n22848_, new_n22849_, new_n22850_, new_n22851_,
    new_n22852_, new_n22853_, new_n22854_, new_n22855_, new_n22856_,
    new_n22857_, new_n22858_, new_n22859_, new_n22860_, new_n22861_,
    new_n22862_, new_n22863_, new_n22864_, new_n22865_, new_n22866_,
    new_n22867_, new_n22868_, new_n22869_, new_n22870_, new_n22871_,
    new_n22872_, new_n22873_, new_n22874_, new_n22875_, new_n22876_,
    new_n22877_, new_n22878_, new_n22879_, new_n22880_, new_n22881_,
    new_n22882_, new_n22883_, new_n22884_, new_n22885_, new_n22886_,
    new_n22887_, new_n22888_, new_n22889_, new_n22890_, new_n22891_,
    new_n22892_, new_n22893_, new_n22894_, new_n22895_, new_n22896_,
    new_n22897_, new_n22898_, new_n22899_, new_n22900_, new_n22901_,
    new_n22902_, new_n22903_, new_n22904_, new_n22905_, new_n22906_,
    new_n22907_, new_n22908_, new_n22909_, new_n22910_, new_n22911_,
    new_n22912_, new_n22913_, new_n22914_, new_n22915_, new_n22916_,
    new_n22917_, new_n22918_, new_n22919_, new_n22920_, new_n22921_,
    new_n22922_, new_n22923_, new_n22924_, new_n22925_, new_n22926_,
    new_n22927_, new_n22928_, new_n22929_, new_n22930_, new_n22931_,
    new_n22932_, new_n22933_, new_n22934_, new_n22935_, new_n22936_,
    new_n22937_, new_n22938_, new_n22939_, new_n22940_, new_n22941_,
    new_n22942_, new_n22943_, new_n22944_, new_n22945_, new_n22946_,
    new_n22947_, new_n22948_, new_n22949_, new_n22950_, new_n22951_,
    new_n22952_, new_n22953_, new_n22954_, new_n22955_, new_n22956_,
    new_n22957_, new_n22958_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23023_, new_n23024_, new_n23025_, new_n23026_,
    new_n23027_, new_n23028_, new_n23029_, new_n23030_, new_n23031_,
    new_n23032_, new_n23033_, new_n23034_, new_n23035_, new_n23036_,
    new_n23037_, new_n23038_, new_n23039_, new_n23040_, new_n23041_,
    new_n23042_, new_n23043_, new_n23044_, new_n23045_, new_n23046_,
    new_n23047_, new_n23048_, new_n23049_, new_n23050_, new_n23051_,
    new_n23052_, new_n23053_, new_n23054_, new_n23055_, new_n23056_,
    new_n23057_, new_n23058_, new_n23059_, new_n23060_, new_n23061_,
    new_n23062_, new_n23063_, new_n23064_, new_n23065_, new_n23066_,
    new_n23067_, new_n23068_, new_n23069_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23097_, new_n23098_, new_n23099_, new_n23100_, new_n23101_,
    new_n23102_, new_n23103_, new_n23104_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23150_, new_n23151_,
    new_n23152_, new_n23153_, new_n23154_, new_n23155_, new_n23156_,
    new_n23157_, new_n23158_, new_n23159_, new_n23160_, new_n23161_,
    new_n23162_, new_n23163_, new_n23164_, new_n23165_, new_n23166_,
    new_n23167_, new_n23168_, new_n23169_, new_n23170_, new_n23171_,
    new_n23172_, new_n23173_, new_n23174_, new_n23175_, new_n23176_,
    new_n23177_, new_n23178_, new_n23179_, new_n23180_, new_n23181_,
    new_n23182_, new_n23183_, new_n23184_, new_n23185_, new_n23186_,
    new_n23187_, new_n23188_, new_n23189_, new_n23190_, new_n23191_,
    new_n23192_, new_n23193_, new_n23194_, new_n23195_, new_n23196_,
    new_n23197_, new_n23198_, new_n23199_, new_n23200_, new_n23201_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23213_, new_n23214_, new_n23215_, new_n23216_,
    new_n23217_, new_n23218_, new_n23219_, new_n23220_, new_n23221_,
    new_n23222_, new_n23223_, new_n23224_, new_n23225_, new_n23226_,
    new_n23227_, new_n23228_, new_n23229_, new_n23230_, new_n23231_,
    new_n23232_, new_n23233_, new_n23234_, new_n23235_, new_n23236_,
    new_n23237_, new_n23238_, new_n23239_, new_n23240_, new_n23241_,
    new_n23242_, new_n23243_, new_n23244_, new_n23245_, new_n23246_,
    new_n23247_, new_n23248_, new_n23249_, new_n23250_, new_n23251_,
    new_n23252_, new_n23253_, new_n23254_, new_n23255_, new_n23256_,
    new_n23257_, new_n23258_, new_n23259_, new_n23260_, new_n23261_,
    new_n23262_, new_n23263_, new_n23264_, new_n23265_, new_n23266_,
    new_n23267_, new_n23268_, new_n23269_, new_n23270_, new_n23271_,
    new_n23272_, new_n23273_, new_n23274_, new_n23275_, new_n23276_,
    new_n23277_, new_n23278_, new_n23279_, new_n23280_, new_n23281_,
    new_n23282_, new_n23283_, new_n23284_, new_n23285_, new_n23286_,
    new_n23287_, new_n23288_, new_n23289_, new_n23290_, new_n23291_,
    new_n23292_, new_n23293_, new_n23294_, new_n23295_, new_n23296_,
    new_n23297_, new_n23298_, new_n23299_, new_n23300_, new_n23301_,
    new_n23302_, new_n23303_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23313_, new_n23314_, new_n23315_, new_n23316_,
    new_n23317_, new_n23318_, new_n23319_, new_n23320_, new_n23321_,
    new_n23322_, new_n23323_, new_n23324_, new_n23325_, new_n23326_,
    new_n23327_, new_n23328_, new_n23329_, new_n23330_, new_n23331_,
    new_n23332_, new_n23333_, new_n23334_, new_n23335_, new_n23336_,
    new_n23337_, new_n23338_, new_n23339_, new_n23340_, new_n23341_,
    new_n23342_, new_n23343_, new_n23344_, new_n23345_, new_n23346_,
    new_n23347_, new_n23348_, new_n23349_, new_n23350_, new_n23351_,
    new_n23352_, new_n23353_, new_n23354_, new_n23355_, new_n23356_,
    new_n23357_, new_n23358_, new_n23359_, new_n23360_, new_n23361_,
    new_n23362_, new_n23363_, new_n23364_, new_n23365_, new_n23366_,
    new_n23367_, new_n23368_, new_n23369_, new_n23370_, new_n23371_,
    new_n23372_, new_n23373_, new_n23374_, new_n23375_, new_n23376_,
    new_n23377_, new_n23378_, new_n23379_, new_n23380_, new_n23381_,
    new_n23382_, new_n23383_, new_n23384_, new_n23385_, new_n23386_,
    new_n23387_, new_n23388_, new_n23389_, new_n23390_, new_n23391_,
    new_n23392_, new_n23393_, new_n23394_, new_n23395_, new_n23396_,
    new_n23397_, new_n23398_, new_n23399_, new_n23400_, new_n23401_,
    new_n23402_, new_n23403_, new_n23404_, new_n23405_, new_n23406_,
    new_n23407_, new_n23408_, new_n23409_, new_n23410_, new_n23411_,
    new_n23412_, new_n23413_, new_n23414_, new_n23415_, new_n23416_,
    new_n23417_, new_n23418_, new_n23419_, new_n23420_, new_n23421_,
    new_n23422_, new_n23423_, new_n23424_, new_n23425_, new_n23426_,
    new_n23427_, new_n23428_, new_n23429_, new_n23430_, new_n23431_,
    new_n23432_, new_n23433_, new_n23434_, new_n23435_, new_n23436_,
    new_n23437_, new_n23438_, new_n23439_, new_n23440_, new_n23441_,
    new_n23442_, new_n23443_, new_n23444_, new_n23445_, new_n23446_,
    new_n23447_, new_n23448_, new_n23449_, new_n23450_, new_n23451_,
    new_n23452_, new_n23453_, new_n23454_, new_n23455_, new_n23456_,
    new_n23457_, new_n23458_, new_n23459_, new_n23460_, new_n23461_,
    new_n23462_, new_n23463_, new_n23464_, new_n23465_, new_n23466_,
    new_n23467_, new_n23468_, new_n23469_, new_n23470_, new_n23471_,
    new_n23472_, new_n23473_, new_n23474_, new_n23475_, new_n23476_,
    new_n23477_, new_n23478_, new_n23479_, new_n23480_, new_n23481_,
    new_n23482_, new_n23483_, new_n23484_, new_n23485_, new_n23486_,
    new_n23487_, new_n23488_, new_n23489_, new_n23490_, new_n23491_,
    new_n23492_, new_n23493_, new_n23494_, new_n23495_, new_n23496_,
    new_n23497_, new_n23498_, new_n23499_, new_n23500_, new_n23501_,
    new_n23502_, new_n23503_, new_n23504_, new_n23505_, new_n23506_,
    new_n23507_, new_n23508_, new_n23509_, new_n23510_, new_n23511_,
    new_n23512_, new_n23513_, new_n23514_, new_n23515_, new_n23516_,
    new_n23517_, new_n23518_, new_n23519_, new_n23520_, new_n23521_,
    new_n23522_, new_n23523_, new_n23524_, new_n23525_, new_n23526_,
    new_n23527_, new_n23528_, new_n23529_, new_n23530_, new_n23531_,
    new_n23532_, new_n23533_, new_n23534_, new_n23535_, new_n23536_,
    new_n23537_, new_n23538_, new_n23539_, new_n23540_, new_n23541_,
    new_n23542_, new_n23543_, new_n23544_, new_n23545_, new_n23546_,
    new_n23547_, new_n23548_, new_n23549_, new_n23550_, new_n23551_,
    new_n23552_, new_n23553_, new_n23554_, new_n23555_, new_n23556_,
    new_n23557_, new_n23558_, new_n23559_, new_n23560_, new_n23561_,
    new_n23562_, new_n23563_, new_n23564_, new_n23565_, new_n23566_,
    new_n23567_, new_n23568_, new_n23569_, new_n23570_, new_n23571_,
    new_n23572_, new_n23573_, new_n23574_, new_n23575_, new_n23576_,
    new_n23577_, new_n23578_, new_n23579_, new_n23580_, new_n23581_,
    new_n23582_, new_n23583_, new_n23584_, new_n23585_, new_n23586_,
    new_n23587_, new_n23588_, new_n23589_, new_n23590_, new_n23591_,
    new_n23592_, new_n23593_, new_n23594_, new_n23595_, new_n23596_,
    new_n23597_, new_n23598_, new_n23599_, new_n23600_, new_n23601_,
    new_n23602_, new_n23603_, new_n23604_, new_n23605_, new_n23606_,
    new_n23607_, new_n23608_, new_n23609_, new_n23610_, new_n23611_,
    new_n23612_, new_n23613_, new_n23614_, new_n23615_, new_n23616_,
    new_n23617_, new_n23618_, new_n23619_, new_n23620_, new_n23621_,
    new_n23622_, new_n23623_, new_n23624_, new_n23625_, new_n23626_,
    new_n23627_, new_n23628_, new_n23629_, new_n23630_, new_n23631_,
    new_n23632_, new_n23633_, new_n23634_, new_n23635_, new_n23636_,
    new_n23637_, new_n23638_, new_n23639_, new_n23640_, new_n23641_,
    new_n23642_, new_n23643_, new_n23644_, new_n23645_, new_n23646_,
    new_n23647_, new_n23648_, new_n23649_, new_n23650_, new_n23651_,
    new_n23652_, new_n23653_, new_n23654_, new_n23655_, new_n23656_,
    new_n23657_, new_n23658_, new_n23659_, new_n23660_, new_n23661_,
    new_n23662_, new_n23663_, new_n23664_, new_n23665_, new_n23666_,
    new_n23667_, new_n23668_, new_n23669_, new_n23670_, new_n23671_,
    new_n23672_, new_n23673_, new_n23674_, new_n23675_, new_n23676_,
    new_n23677_, new_n23678_, new_n23679_, new_n23680_, new_n23681_,
    new_n23682_, new_n23683_, new_n23684_, new_n23685_, new_n23686_,
    new_n23687_, new_n23688_, new_n23689_, new_n23690_, new_n23691_,
    new_n23692_, new_n23693_, new_n23694_, new_n23695_, new_n23696_,
    new_n23697_, new_n23698_, new_n23699_, new_n23700_, new_n23701_,
    new_n23702_, new_n23703_, new_n23704_, new_n23705_, new_n23706_,
    new_n23707_, new_n23708_, new_n23709_, new_n23710_, new_n23711_,
    new_n23712_, new_n23713_, new_n23714_, new_n23715_, new_n23716_,
    new_n23717_, new_n23718_, new_n23719_, new_n23720_, new_n23721_,
    new_n23722_, new_n23723_, new_n23724_, new_n23725_, new_n23726_,
    new_n23727_, new_n23728_, new_n23729_, new_n23730_, new_n23731_,
    new_n23732_, new_n23733_, new_n23734_, new_n23735_, new_n23736_,
    new_n23737_, new_n23738_, new_n23739_, new_n23740_, new_n23741_,
    new_n23742_, new_n23743_, new_n23744_, new_n23745_, new_n23746_,
    new_n23747_, new_n23748_, new_n23749_, new_n23750_, new_n23751_,
    new_n23752_, new_n23753_, new_n23754_, new_n23755_, new_n23756_,
    new_n23757_, new_n23758_, new_n23759_, new_n23760_, new_n23761_,
    new_n23762_, new_n23763_, new_n23764_, new_n23765_, new_n23766_,
    new_n23767_, new_n23768_, new_n23769_, new_n23770_, new_n23771_,
    new_n23772_, new_n23773_, new_n23774_, new_n23775_, new_n23776_,
    new_n23777_, new_n23778_, new_n23779_, new_n23780_, new_n23781_,
    new_n23782_, new_n23783_, new_n23784_, new_n23785_, new_n23786_,
    new_n23787_, new_n23788_, new_n23789_, new_n23790_, new_n23791_,
    new_n23792_, new_n23793_, new_n23794_, new_n23795_, new_n23796_,
    new_n23797_, new_n23798_, new_n23799_, new_n23800_, new_n23801_,
    new_n23802_, new_n23803_, new_n23804_, new_n23805_, new_n23806_,
    new_n23807_, new_n23808_, new_n23809_, new_n23810_, new_n23811_,
    new_n23812_, new_n23813_, new_n23814_, new_n23815_, new_n23816_,
    new_n23817_, new_n23818_, new_n23819_, new_n23820_, new_n23821_,
    new_n23822_, new_n23823_, new_n23824_, new_n23825_, new_n23826_,
    new_n23827_, new_n23828_, new_n23829_, new_n23830_, new_n23831_,
    new_n23832_, new_n23833_, new_n23834_, new_n23835_, new_n23836_,
    new_n23837_, new_n23838_, new_n23839_, new_n23840_, new_n23841_,
    new_n23842_, new_n23843_, new_n23844_, new_n23845_, new_n23846_,
    new_n23847_, new_n23848_, new_n23849_, new_n23850_, new_n23851_,
    new_n23852_, new_n23853_, new_n23854_, new_n23855_, new_n23856_,
    new_n23857_, new_n23858_, new_n23859_, new_n23860_, new_n23861_,
    new_n23862_, new_n23863_, new_n23864_, new_n23865_, new_n23866_,
    new_n23867_, new_n23868_, new_n23869_, new_n23870_, new_n23871_,
    new_n23872_, new_n23873_, new_n23874_, new_n23875_, new_n23876_,
    new_n23877_, new_n23878_, new_n23879_, new_n23880_, new_n23881_,
    new_n23882_, new_n23883_, new_n23884_, new_n23885_, new_n23886_,
    new_n23887_, new_n23888_, new_n23889_, new_n23890_, new_n23891_,
    new_n23892_, new_n23893_, new_n23894_, new_n23895_, new_n23896_,
    new_n23897_, new_n23898_, new_n23899_, new_n23900_, new_n23901_,
    new_n23902_, new_n23903_, new_n23904_, new_n23905_, new_n23906_,
    new_n23907_, new_n23908_, new_n23909_, new_n23910_, new_n23911_,
    new_n23912_, new_n23913_, new_n23914_, new_n23915_, new_n23916_,
    new_n23917_, new_n23918_, new_n23919_, new_n23920_, new_n23921_,
    new_n23922_, new_n23923_, new_n23924_, new_n23925_, new_n23926_,
    new_n23927_, new_n23928_, new_n23929_, new_n23930_, new_n23931_,
    new_n23932_, new_n23933_, new_n23934_, new_n23935_, new_n23936_,
    new_n23937_, new_n23938_, new_n23939_, new_n23940_, new_n23941_,
    new_n23942_, new_n23943_, new_n23944_, new_n23945_, new_n23946_,
    new_n23947_, new_n23948_, new_n23949_, new_n23950_, new_n23951_,
    new_n23952_, new_n23953_, new_n23954_, new_n23955_, new_n23956_,
    new_n23957_, new_n23958_, new_n23959_, new_n23960_, new_n23961_,
    new_n23962_, new_n23963_, new_n23964_, new_n23965_, new_n23966_,
    new_n23967_, new_n23968_, new_n23969_, new_n23970_, new_n23971_,
    new_n23972_, new_n23973_, new_n23974_, new_n23975_, new_n23976_,
    new_n23977_, new_n23978_, new_n23979_, new_n23980_, new_n23981_,
    new_n23982_, new_n23983_, new_n23984_, new_n23985_, new_n23986_,
    new_n23987_, new_n23988_, new_n23989_, new_n23990_, new_n23991_,
    new_n23992_, new_n23993_, new_n23994_, new_n23995_, new_n23996_,
    new_n23997_, new_n23998_, new_n23999_, new_n24000_, new_n24001_,
    new_n24002_, new_n24003_, new_n24004_, new_n24005_, new_n24006_,
    new_n24007_, new_n24008_, new_n24009_, new_n24010_, new_n24011_,
    new_n24012_, new_n24013_, new_n24014_, new_n24015_, new_n24016_,
    new_n24017_, new_n24018_, new_n24019_, new_n24020_, new_n24021_,
    new_n24022_, new_n24023_, new_n24024_, new_n24025_, new_n24026_,
    new_n24027_, new_n24028_, new_n24029_, new_n24030_, new_n24031_,
    new_n24032_, new_n24033_, new_n24034_, new_n24035_, new_n24036_,
    new_n24037_, new_n24038_, new_n24039_, new_n24040_, new_n24041_,
    new_n24042_, new_n24043_, new_n24044_, new_n24045_, new_n24046_,
    new_n24047_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24074_, new_n24075_, new_n24076_,
    new_n24077_, new_n24078_, new_n24079_, new_n24080_, new_n24081_,
    new_n24082_, new_n24083_, new_n24084_, new_n24085_, new_n24086_,
    new_n24087_, new_n24088_, new_n24089_, new_n24090_, new_n24091_,
    new_n24092_, new_n24093_, new_n24094_, new_n24095_, new_n24096_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24240_, new_n24241_,
    new_n24242_, new_n24243_, new_n24244_, new_n24245_, new_n24246_,
    new_n24247_, new_n24248_, new_n24249_, new_n24250_, new_n24251_,
    new_n24252_, new_n24253_, new_n24254_, new_n24255_, new_n24256_,
    new_n24257_, new_n24258_, new_n24259_, new_n24260_, new_n24261_,
    new_n24262_, new_n24263_, new_n24264_, new_n24265_, new_n24266_,
    new_n24267_, new_n24268_, new_n24269_, new_n24270_, new_n24271_,
    new_n24272_, new_n24273_, new_n24274_, new_n24275_, new_n24276_,
    new_n24277_, new_n24278_, new_n24279_, new_n24280_, new_n24281_,
    new_n24282_, new_n24283_, new_n24284_, new_n24285_, new_n24286_,
    new_n24287_, new_n24288_, new_n24289_, new_n24290_, new_n24291_,
    new_n24292_, new_n24293_, new_n24294_, new_n24295_, new_n24296_,
    new_n24297_, new_n24298_, new_n24299_, new_n24300_, new_n24301_,
    new_n24302_, new_n24303_, new_n24304_, new_n24305_, new_n24306_,
    new_n24307_, new_n24308_, new_n24309_, new_n24310_, new_n24311_,
    new_n24312_, new_n24313_, new_n24314_, new_n24315_, new_n24316_,
    new_n24317_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24336_,
    new_n24337_, new_n24338_, new_n24339_, new_n24340_, new_n24341_,
    new_n24342_, new_n24343_, new_n24344_, new_n24345_, new_n24346_,
    new_n24347_, new_n24348_, new_n24349_, new_n24350_, new_n24351_,
    new_n24352_, new_n24353_, new_n24354_, new_n24355_, new_n24356_,
    new_n24357_, new_n24358_, new_n24359_, new_n24360_, new_n24361_,
    new_n24362_, new_n24363_, new_n24364_, new_n24365_, new_n24366_,
    new_n24367_, new_n24368_, new_n24369_, new_n24370_, new_n24371_,
    new_n24372_, new_n24373_, new_n24374_, new_n24375_, new_n24376_,
    new_n24377_, new_n24378_, new_n24379_, new_n24380_, new_n24381_,
    new_n24382_, new_n24383_, new_n24384_, new_n24385_, new_n24386_,
    new_n24387_, new_n24388_, new_n24389_, new_n24390_, new_n24391_,
    new_n24392_, new_n24393_, new_n24394_, new_n24395_, new_n24396_,
    new_n24397_, new_n24398_, new_n24399_, new_n24400_, new_n24401_,
    new_n24402_, new_n24403_, new_n24404_, new_n24405_, new_n24406_,
    new_n24407_, new_n24408_, new_n24409_, new_n24410_, new_n24411_,
    new_n24412_, new_n24413_, new_n24414_, new_n24415_, new_n24416_,
    new_n24417_, new_n24418_, new_n24419_, new_n24420_, new_n24421_,
    new_n24422_, new_n24423_, new_n24424_, new_n24425_, new_n24426_,
    new_n24427_, new_n24428_, new_n24429_, new_n24430_, new_n24431_,
    new_n24432_, new_n24433_, new_n24434_, new_n24435_, new_n24436_,
    new_n24437_, new_n24438_, new_n24439_, new_n24440_, new_n24441_,
    new_n24442_, new_n24443_, new_n24444_, new_n24445_, new_n24446_,
    new_n24447_, new_n24448_, new_n24449_, new_n24450_, new_n24451_,
    new_n24452_, new_n24453_, new_n24454_, new_n24455_, new_n24456_,
    new_n24457_, new_n24458_, new_n24459_, new_n24460_, new_n24461_,
    new_n24462_, new_n24463_, new_n24464_, new_n24465_, new_n24466_,
    new_n24467_, new_n24468_, new_n24469_, new_n24470_, new_n24471_,
    new_n24472_, new_n24473_, new_n24474_, new_n24475_, new_n24476_,
    new_n24477_, new_n24478_, new_n24479_, new_n24480_, new_n24481_,
    new_n24482_, new_n24483_, new_n24484_, new_n24485_, new_n24486_,
    new_n24487_, new_n24488_, new_n24489_, new_n24490_, new_n24491_,
    new_n24492_, new_n24493_, new_n24494_, new_n24495_, new_n24496_,
    new_n24497_, new_n24498_, new_n24499_, new_n24500_, new_n24501_,
    new_n24502_, new_n24503_, new_n24504_, new_n24505_, new_n24506_,
    new_n24507_, new_n24508_, new_n24509_, new_n24510_, new_n24511_,
    new_n24512_, new_n24513_, new_n24514_, new_n24515_, new_n24516_,
    new_n24517_, new_n24518_, new_n24519_, new_n24520_, new_n24521_,
    new_n24522_, new_n24523_, new_n24524_, new_n24525_, new_n24526_,
    new_n24527_, new_n24528_, new_n24529_, new_n24530_, new_n24531_,
    new_n24532_, new_n24533_, new_n24534_, new_n24535_, new_n24536_,
    new_n24537_, new_n24538_, new_n24539_, new_n24540_, new_n24541_,
    new_n24542_, new_n24543_, new_n24544_, new_n24545_, new_n24546_,
    new_n24547_, new_n24548_, new_n24549_, new_n24550_, new_n24551_,
    new_n24552_, new_n24553_, new_n24554_, new_n24555_, new_n24556_,
    new_n24557_, new_n24558_, new_n24559_, new_n24560_, new_n24561_,
    new_n24562_, new_n24563_, new_n24564_, new_n24565_, new_n24566_,
    new_n24567_, new_n24568_, new_n24569_, new_n24570_, new_n24571_,
    new_n24572_, new_n24573_, new_n24574_, new_n24575_, new_n24576_,
    new_n24577_, new_n24578_, new_n24579_, new_n24580_, new_n24581_,
    new_n24582_, new_n24583_, new_n24584_, new_n24585_, new_n24586_,
    new_n24587_, new_n24588_, new_n24589_, new_n24590_, new_n24591_,
    new_n24592_, new_n24593_, new_n24594_, new_n24595_, new_n24596_,
    new_n24597_, new_n24598_, new_n24599_, new_n24600_, new_n24601_,
    new_n24602_, new_n24603_, new_n24604_, new_n24605_, new_n24606_,
    new_n24607_, new_n24608_, new_n24609_, new_n24610_, new_n24611_,
    new_n24612_, new_n24613_, new_n24614_, new_n24615_, new_n24616_,
    new_n24617_, new_n24618_, new_n24619_, new_n24620_, new_n24621_,
    new_n24622_, new_n24623_, new_n24624_, new_n24625_, new_n24626_,
    new_n24627_, new_n24628_, new_n24629_, new_n24630_, new_n24631_,
    new_n24632_, new_n24633_, new_n24634_, new_n24635_, new_n24636_,
    new_n24637_, new_n24638_, new_n24639_, new_n24640_, new_n24641_,
    new_n24642_, new_n24643_, new_n24644_, new_n24645_, new_n24646_,
    new_n24647_, new_n24648_, new_n24649_, new_n24650_, new_n24651_,
    new_n24652_, new_n24653_, new_n24654_, new_n24655_, new_n24656_,
    new_n24657_, new_n24658_, new_n24659_, new_n24660_, new_n24661_,
    new_n24662_, new_n24663_, new_n24664_, new_n24665_, new_n24666_,
    new_n24667_, new_n24668_, new_n24669_, new_n24670_, new_n24671_,
    new_n24672_, new_n24673_, new_n24674_, new_n24675_, new_n24676_,
    new_n24677_, new_n24678_, new_n24679_, new_n24680_, new_n24681_,
    new_n24682_, new_n24683_, new_n24684_, new_n24685_, new_n24686_,
    new_n24687_, new_n24688_, new_n24689_, new_n24690_, new_n24691_,
    new_n24692_, new_n24693_, new_n24694_, new_n24695_, new_n24696_,
    new_n24697_, new_n24698_, new_n24699_, new_n24700_, new_n24701_,
    new_n24702_, new_n24703_, new_n24704_, new_n24705_, new_n24706_,
    new_n24707_, new_n24708_, new_n24709_, new_n24710_, new_n24711_,
    new_n24712_, new_n24713_, new_n24714_, new_n24715_, new_n24716_,
    new_n24717_, new_n24718_, new_n24719_, new_n24720_, new_n24721_,
    new_n24722_, new_n24723_, new_n24724_, new_n24725_, new_n24726_,
    new_n24727_, new_n24728_, new_n24729_, new_n24730_, new_n24731_,
    new_n24732_, new_n24733_, new_n24734_, new_n24735_, new_n24736_,
    new_n24737_, new_n24738_, new_n24739_, new_n24740_, new_n24741_,
    new_n24742_, new_n24743_, new_n24744_, new_n24745_, new_n24746_,
    new_n24747_, new_n24748_, new_n24749_, new_n24750_, new_n24751_,
    new_n24752_, new_n24753_, new_n24754_, new_n24755_, new_n24756_,
    new_n24757_, new_n24758_, new_n24759_, new_n24760_, new_n24761_,
    new_n24762_, new_n24763_, new_n24764_, new_n24765_, new_n24766_,
    new_n24767_, new_n24768_, new_n24769_, new_n24770_, new_n24771_,
    new_n24772_, new_n24773_, new_n24774_, new_n24775_, new_n24776_,
    new_n24777_, new_n24778_, new_n24779_, new_n24780_, new_n24781_,
    new_n24782_, new_n24783_, new_n24784_, new_n24785_, new_n24786_,
    new_n24787_, new_n24788_, new_n24789_, new_n24790_, new_n24791_,
    new_n24792_, new_n24793_, new_n24794_, new_n24795_, new_n24796_,
    new_n24797_, new_n24798_, new_n24799_, new_n24800_, new_n24801_,
    new_n24802_, new_n24803_, new_n24804_, new_n24805_, new_n24806_,
    new_n24807_, new_n24808_, new_n24809_, new_n24810_, new_n24811_,
    new_n24812_, new_n24813_, new_n24814_, new_n24815_, new_n24816_,
    new_n24817_, new_n24818_, new_n24819_, new_n24820_, new_n24821_,
    new_n24822_, new_n24823_, new_n24824_, new_n24825_, new_n24826_,
    new_n24827_, new_n24828_, new_n24829_, new_n24830_, new_n24831_,
    new_n24832_, new_n24833_, new_n24834_, new_n24835_, new_n24836_,
    new_n24837_, new_n24838_, new_n24839_, new_n24840_, new_n24841_,
    new_n24842_, new_n24843_, new_n24844_, new_n24845_, new_n24846_,
    new_n24847_, new_n24848_, new_n24849_, new_n24850_, new_n24851_,
    new_n24852_, new_n24853_, new_n24854_, new_n24855_, new_n24856_,
    new_n24857_, new_n24858_, new_n24859_, new_n24860_, new_n24861_,
    new_n24862_, new_n24863_, new_n24864_, new_n24865_, new_n24866_,
    new_n24867_, new_n24868_, new_n24869_, new_n24870_, new_n24871_,
    new_n24872_, new_n24873_, new_n24874_, new_n24875_, new_n24876_,
    new_n24877_, new_n24878_, new_n24879_, new_n24880_, new_n24881_,
    new_n24882_, new_n24883_, new_n24884_, new_n24885_, new_n24886_,
    new_n24887_, new_n24888_, new_n24889_, new_n24890_, new_n24891_,
    new_n24892_, new_n24893_, new_n24894_, new_n24895_, new_n24896_,
    new_n24897_, new_n24898_, new_n24899_, new_n24900_, new_n24901_,
    new_n24902_, new_n24903_, new_n24904_, new_n24905_, new_n24906_,
    new_n24907_, new_n24908_, new_n24909_, new_n24910_, new_n24911_,
    new_n24912_, new_n24913_, new_n24914_, new_n24915_, new_n24916_,
    new_n24917_, new_n24918_, new_n24919_, new_n24920_, new_n24921_,
    new_n24922_, new_n24923_, new_n24924_, new_n24925_, new_n24926_,
    new_n24927_, new_n24928_, new_n24929_, new_n24930_, new_n24931_,
    new_n24932_, new_n24933_, new_n24934_, new_n24935_, new_n24936_,
    new_n24937_, new_n24938_, new_n24939_, new_n24940_, new_n24941_,
    new_n24942_, new_n24943_, new_n24944_, new_n24945_, new_n24946_,
    new_n24947_, new_n24948_, new_n24949_, new_n24950_, new_n24951_,
    new_n24952_, new_n24953_, new_n24954_, new_n24955_, new_n24956_,
    new_n24957_, new_n24958_, new_n24959_, new_n24960_, new_n24961_,
    new_n24962_, new_n24963_, new_n24964_, new_n24965_, new_n24966_,
    new_n24967_, new_n24968_, new_n24969_, new_n24970_, new_n24971_,
    new_n24972_, new_n24973_, new_n24974_, new_n24975_, new_n24976_,
    new_n24977_, new_n24978_, new_n24979_, new_n24980_, new_n24981_,
    new_n24982_, new_n24983_, new_n24984_, new_n24985_, new_n24986_,
    new_n24987_, new_n24988_, new_n24989_, new_n24990_, new_n24991_,
    new_n24992_, new_n24993_, new_n24994_, new_n24995_, new_n24996_,
    new_n24997_, new_n24998_, new_n24999_, new_n25000_, new_n25001_,
    new_n25002_, new_n25003_, new_n25004_, new_n25005_, new_n25006_,
    new_n25007_, new_n25008_, new_n25009_, new_n25010_, new_n25011_,
    new_n25012_, new_n25013_, new_n25014_, new_n25015_, new_n25016_,
    new_n25017_, new_n25018_, new_n25019_, new_n25020_, new_n25021_,
    new_n25022_, new_n25023_, new_n25024_, new_n25025_, new_n25026_,
    new_n25027_, new_n25028_, new_n25029_, new_n25030_, new_n25031_,
    new_n25032_, new_n25033_, new_n25034_, new_n25035_, new_n25036_,
    new_n25037_, new_n25038_, new_n25039_, new_n25040_, new_n25041_,
    new_n25042_, new_n25043_, new_n25044_, new_n25045_, new_n25046_,
    new_n25047_, new_n25048_, new_n25049_, new_n25050_, new_n25051_,
    new_n25052_, new_n25053_, new_n25054_, new_n25055_, new_n25056_,
    new_n25057_, new_n25058_, new_n25059_, new_n25060_, new_n25061_,
    new_n25062_, new_n25063_, new_n25064_, new_n25065_, new_n25066_,
    new_n25067_, new_n25068_, new_n25069_, new_n25070_, new_n25071_,
    new_n25072_, new_n25073_, new_n25074_, new_n25075_, new_n25076_,
    new_n25077_, new_n25078_, new_n25079_, new_n25080_, new_n25081_,
    new_n25082_, new_n25083_, new_n25084_, new_n25085_, new_n25086_,
    new_n25087_, new_n25088_, new_n25089_, new_n25090_, new_n25091_,
    new_n25092_, new_n25093_, new_n25094_, new_n25095_, new_n25096_,
    new_n25097_, new_n25098_, new_n25099_, new_n25100_, new_n25101_,
    new_n25102_, new_n25103_, new_n25104_, new_n25105_, new_n25106_,
    new_n25107_, new_n25108_, new_n25109_, new_n25110_, new_n25111_,
    new_n25112_, new_n25113_, new_n25114_, new_n25115_, new_n25116_,
    new_n25117_, new_n25118_, new_n25119_, new_n25120_, new_n25121_,
    new_n25122_, new_n25123_, new_n25124_, new_n25125_, new_n25126_,
    new_n25127_, new_n25128_, new_n25129_, new_n25130_, new_n25131_,
    new_n25132_, new_n25133_, new_n25134_, new_n25135_, new_n25136_,
    new_n25137_, new_n25138_, new_n25139_, new_n25140_, new_n25141_,
    new_n25142_, new_n25143_, new_n25144_, new_n25145_, new_n25146_,
    new_n25147_, new_n25148_, new_n25149_, new_n25150_, new_n25151_,
    new_n25152_, new_n25153_, new_n25154_, new_n25155_;
  assign new_n27_ = A302 & ~A301;
  assign new_n28_ = ~A300 & new_n27_;
  assign new_n29_ = A299 & ~A298;
  assign new_n30_ = new_n28_ & new_n29_;
  assign new_n31_ = A269 & ~A268;
  assign new_n32_ = A267 & A236;
  assign new_n33_ = new_n31_ & new_n32_;
  assign new_n34_ = new_n30_ & new_n33_;
  assign new_n35_ = ~A235 & ~A234;
  assign new_n36_ = ~A233 & new_n35_;
  assign new_n37_ = A232 & A166;
  assign new_n38_ = new_n36_ & new_n37_;
  assign new_n39_ = ~A167 & ~A168;
  assign new_n40_ = ~A169 & ~A170;
  assign new_n41_ = new_n39_ & new_n40_;
  assign new_n42_ = new_n38_ & new_n41_;
  assign new_n43_ = new_n34_ & new_n42_;
  assign new_n44_ = A300 & new_n27_;
  assign new_n45_ = new_n31_ & new_n44_;
  assign new_n46_ = ~A267 & ~A266;
  assign new_n47_ = A265 & A236;
  assign new_n48_ = new_n46_ & new_n47_;
  assign new_n49_ = new_n45_ & new_n48_;
  assign new_n50_ = new_n42_ & new_n49_;
  assign new_n51_ = ~A267 & A266;
  assign new_n52_ = ~A265 & A236;
  assign new_n53_ = new_n51_ & new_n52_;
  assign new_n54_ = new_n45_ & new_n53_;
  assign new_n55_ = new_n42_ & new_n54_;
  assign new_n56_ = ~new_n50_ & ~new_n55_;
  assign new_n57_ = ~new_n43_ & new_n56_;
  assign new_n58_ = A233 & new_n35_;
  assign new_n59_ = ~A232 & A166;
  assign new_n60_ = new_n58_ & new_n59_;
  assign new_n61_ = new_n41_ & new_n60_;
  assign new_n62_ = new_n54_ & new_n61_;
  assign new_n63_ = ~A299 & A298;
  assign new_n64_ = new_n28_ & new_n63_;
  assign new_n65_ = new_n33_ & new_n64_;
  assign new_n66_ = new_n42_ & new_n65_;
  assign new_n67_ = new_n49_ & new_n61_;
  assign new_n68_ = ~new_n66_ & ~new_n67_;
  assign new_n69_ = ~new_n62_ & new_n68_;
  assign new_n70_ = new_n57_ & new_n69_;
  assign new_n71_ = A232 & ~A166;
  assign new_n72_ = new_n36_ & new_n71_;
  assign new_n73_ = A167 & ~A168;
  assign new_n74_ = new_n40_ & new_n73_;
  assign new_n75_ = new_n72_ & new_n74_;
  assign new_n76_ = new_n49_ & new_n75_;
  assign new_n77_ = new_n34_ & new_n61_;
  assign new_n78_ = new_n61_ & new_n65_;
  assign new_n79_ = ~new_n77_ & ~new_n78_;
  assign new_n80_ = ~new_n76_ & new_n79_;
  assign new_n81_ = new_n65_ & new_n75_;
  assign new_n82_ = new_n54_ & new_n75_;
  assign new_n83_ = new_n34_ & new_n75_;
  assign new_n84_ = ~new_n82_ & ~new_n83_;
  assign new_n85_ = ~new_n81_ & new_n84_;
  assign new_n86_ = new_n80_ & new_n85_;
  assign new_n87_ = new_n70_ & new_n86_;
  assign new_n88_ = ~A232 & ~A166;
  assign new_n89_ = new_n58_ & new_n88_;
  assign new_n90_ = new_n74_ & new_n89_;
  assign new_n91_ = new_n34_ & new_n90_;
  assign new_n92_ = new_n49_ & new_n90_;
  assign new_n93_ = new_n54_ & new_n90_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ~new_n91_ & new_n94_;
  assign new_n96_ = A232 & A203;
  assign new_n97_ = new_n36_ & new_n96_;
  assign new_n98_ = ~A202 & ~A201;
  assign new_n99_ = ~A200 & A199;
  assign new_n100_ = new_n98_ & new_n99_;
  assign new_n101_ = new_n97_ & new_n100_;
  assign new_n102_ = new_n54_ & new_n101_;
  assign new_n103_ = new_n65_ & new_n90_;
  assign new_n104_ = new_n49_ & new_n101_;
  assign new_n105_ = ~new_n103_ & ~new_n104_;
  assign new_n106_ = ~new_n102_ & new_n105_;
  assign new_n107_ = new_n95_ & new_n106_;
  assign new_n108_ = ~A232 & A203;
  assign new_n109_ = new_n58_ & new_n108_;
  assign new_n110_ = new_n100_ & new_n109_;
  assign new_n111_ = new_n49_ & new_n110_;
  assign new_n112_ = new_n34_ & new_n101_;
  assign new_n113_ = new_n65_ & new_n101_;
  assign new_n114_ = ~new_n112_ & ~new_n113_;
  assign new_n115_ = ~new_n111_ & new_n114_;
  assign new_n116_ = new_n65_ & new_n110_;
  assign new_n117_ = new_n54_ & new_n110_;
  assign new_n118_ = new_n34_ & new_n110_;
  assign new_n119_ = ~new_n117_ & ~new_n118_;
  assign new_n120_ = ~new_n116_ & new_n119_;
  assign new_n121_ = new_n115_ & new_n120_;
  assign new_n122_ = new_n107_ & new_n121_;
  assign new_n123_ = new_n87_ & new_n122_;
  assign new_n124_ = A200 & ~A199;
  assign new_n125_ = new_n98_ & new_n124_;
  assign new_n126_ = new_n97_ & new_n125_;
  assign new_n127_ = new_n34_ & new_n126_;
  assign new_n128_ = new_n49_ & new_n126_;
  assign new_n129_ = new_n54_ & new_n126_;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_ = ~new_n127_ & new_n130_;
  assign new_n132_ = new_n109_ & new_n125_;
  assign new_n133_ = new_n54_ & new_n132_;
  assign new_n134_ = new_n65_ & new_n126_;
  assign new_n135_ = new_n49_ & new_n132_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = ~new_n133_ & new_n136_;
  assign new_n138_ = new_n131_ & new_n137_;
  assign new_n139_ = ~A266 & ~A265;
  assign new_n140_ = A236 & ~A235;
  assign new_n141_ = new_n139_ & new_n140_;
  assign new_n142_ = new_n30_ & new_n141_;
  assign new_n143_ = ~A234 & ~A233;
  assign new_n144_ = new_n37_ & new_n143_;
  assign new_n145_ = new_n41_ & new_n144_;
  assign new_n146_ = new_n142_ & new_n145_;
  assign new_n147_ = new_n34_ & new_n132_;
  assign new_n148_ = new_n65_ & new_n132_;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_ = ~new_n146_ & new_n149_;
  assign new_n151_ = A299 & A298;
  assign new_n152_ = A269 & new_n151_;
  assign new_n153_ = ~A268 & ~A267;
  assign new_n154_ = new_n152_ & new_n153_;
  assign new_n155_ = ~A266 & A265;
  assign new_n156_ = new_n140_ & new_n155_;
  assign new_n157_ = new_n154_ & new_n156_;
  assign new_n158_ = new_n145_ & new_n157_;
  assign new_n159_ = new_n64_ & new_n141_;
  assign new_n160_ = new_n145_ & new_n159_;
  assign new_n161_ = ~A299 & ~A298;
  assign new_n162_ = A269 & new_n161_;
  assign new_n163_ = new_n153_ & new_n162_;
  assign new_n164_ = new_n156_ & new_n163_;
  assign new_n165_ = new_n145_ & new_n164_;
  assign new_n166_ = ~new_n160_ & ~new_n165_;
  assign new_n167_ = ~new_n158_ & new_n166_;
  assign new_n168_ = new_n150_ & new_n167_;
  assign new_n169_ = new_n138_ & new_n168_;
  assign new_n170_ = ~A269 & A267;
  assign new_n171_ = new_n44_ & new_n170_;
  assign new_n172_ = new_n156_ & new_n171_;
  assign new_n173_ = new_n145_ & new_n172_;
  assign new_n174_ = ~A302 & ~A300;
  assign new_n175_ = A269 & new_n174_;
  assign new_n176_ = new_n153_ & new_n175_;
  assign new_n177_ = new_n156_ & new_n176_;
  assign new_n178_ = new_n145_ & new_n177_;
  assign new_n179_ = A301 & ~A300;
  assign new_n180_ = A269 & new_n179_;
  assign new_n181_ = new_n153_ & new_n180_;
  assign new_n182_ = new_n156_ & new_n181_;
  assign new_n183_ = new_n145_ & new_n182_;
  assign new_n184_ = ~new_n178_ & ~new_n183_;
  assign new_n185_ = ~new_n173_ & new_n184_;
  assign new_n186_ = A266 & ~A265;
  assign new_n187_ = new_n140_ & new_n186_;
  assign new_n188_ = new_n154_ & new_n187_;
  assign new_n189_ = new_n145_ & new_n188_;
  assign new_n190_ = A268 & A267;
  assign new_n191_ = new_n44_ & new_n190_;
  assign new_n192_ = new_n156_ & new_n191_;
  assign new_n193_ = new_n145_ & new_n192_;
  assign new_n194_ = new_n163_ & new_n187_;
  assign new_n195_ = new_n145_ & new_n194_;
  assign new_n196_ = ~new_n193_ & ~new_n195_;
  assign new_n197_ = ~new_n189_ & new_n196_;
  assign new_n198_ = new_n185_ & new_n197_;
  assign new_n199_ = new_n171_ & new_n187_;
  assign new_n200_ = new_n145_ & new_n199_;
  assign new_n201_ = new_n176_ & new_n187_;
  assign new_n202_ = new_n145_ & new_n201_;
  assign new_n203_ = new_n181_ & new_n187_;
  assign new_n204_ = new_n145_ & new_n203_;
  assign new_n205_ = ~new_n202_ & ~new_n204_;
  assign new_n206_ = ~new_n200_ & new_n205_;
  assign new_n207_ = new_n187_ & new_n191_;
  assign new_n208_ = new_n145_ & new_n207_;
  assign new_n209_ = A266 & A265;
  assign new_n210_ = new_n140_ & new_n209_;
  assign new_n211_ = new_n30_ & new_n210_;
  assign new_n212_ = new_n145_ & new_n211_;
  assign new_n213_ = ~new_n208_ & ~new_n212_;
  assign new_n214_ = new_n206_ & new_n213_;
  assign new_n215_ = new_n198_ & new_n214_;
  assign new_n216_ = new_n169_ & new_n215_;
  assign new_n217_ = new_n123_ & new_n216_;
  assign new_n218_ = ~A269 & ~A267;
  assign new_n219_ = new_n140_ & new_n218_;
  assign new_n220_ = new_n64_ & new_n219_;
  assign new_n221_ = new_n145_ & new_n220_;
  assign new_n222_ = new_n64_ & new_n210_;
  assign new_n223_ = new_n145_ & new_n222_;
  assign new_n224_ = new_n30_ & new_n219_;
  assign new_n225_ = new_n145_ & new_n224_;
  assign new_n226_ = ~new_n223_ & ~new_n225_;
  assign new_n227_ = ~new_n221_ & new_n226_;
  assign new_n228_ = ~A302 & A300;
  assign new_n229_ = A299 & new_n228_;
  assign new_n230_ = ~A298 & A269;
  assign new_n231_ = new_n229_ & new_n230_;
  assign new_n232_ = ~A268 & A267;
  assign new_n233_ = new_n140_ & new_n232_;
  assign new_n234_ = new_n231_ & new_n233_;
  assign new_n235_ = new_n145_ & new_n234_;
  assign new_n236_ = A268 & ~A267;
  assign new_n237_ = new_n140_ & new_n236_;
  assign new_n238_ = new_n30_ & new_n237_;
  assign new_n239_ = new_n145_ & new_n238_;
  assign new_n240_ = new_n64_ & new_n237_;
  assign new_n241_ = new_n145_ & new_n240_;
  assign new_n242_ = ~new_n239_ & ~new_n241_;
  assign new_n243_ = ~new_n235_ & new_n242_;
  assign new_n244_ = new_n227_ & new_n243_;
  assign new_n245_ = A301 & A300;
  assign new_n246_ = ~A299 & new_n245_;
  assign new_n247_ = A298 & A269;
  assign new_n248_ = new_n246_ & new_n247_;
  assign new_n249_ = new_n233_ & new_n248_;
  assign new_n250_ = new_n145_ & new_n249_;
  assign new_n251_ = A299 & new_n245_;
  assign new_n252_ = new_n230_ & new_n251_;
  assign new_n253_ = new_n233_ & new_n252_;
  assign new_n254_ = new_n145_ & new_n253_;
  assign new_n255_ = ~A299 & new_n228_;
  assign new_n256_ = new_n247_ & new_n255_;
  assign new_n257_ = new_n233_ & new_n256_;
  assign new_n258_ = new_n145_ & new_n257_;
  assign new_n259_ = ~new_n254_ & ~new_n258_;
  assign new_n260_ = ~new_n250_ & new_n259_;
  assign new_n261_ = A267 & ~A236;
  assign new_n262_ = new_n31_ & new_n261_;
  assign new_n263_ = new_n30_ & new_n262_;
  assign new_n264_ = A234 & ~A233;
  assign new_n265_ = new_n37_ & new_n264_;
  assign new_n266_ = new_n41_ & new_n265_;
  assign new_n267_ = new_n263_ & new_n266_;
  assign new_n268_ = A265 & ~A236;
  assign new_n269_ = new_n46_ & new_n268_;
  assign new_n270_ = new_n45_ & new_n269_;
  assign new_n271_ = new_n266_ & new_n270_;
  assign new_n272_ = ~A265 & ~A236;
  assign new_n273_ = new_n51_ & new_n272_;
  assign new_n274_ = new_n45_ & new_n273_;
  assign new_n275_ = new_n266_ & new_n274_;
  assign new_n276_ = ~new_n271_ & ~new_n275_;
  assign new_n277_ = ~new_n267_ & new_n276_;
  assign new_n278_ = new_n260_ & new_n277_;
  assign new_n279_ = new_n244_ & new_n278_;
  assign new_n280_ = ~A265 & A235;
  assign new_n281_ = new_n51_ & new_n280_;
  assign new_n282_ = new_n45_ & new_n281_;
  assign new_n283_ = new_n266_ & new_n282_;
  assign new_n284_ = new_n64_ & new_n262_;
  assign new_n285_ = new_n266_ & new_n284_;
  assign new_n286_ = A265 & A235;
  assign new_n287_ = new_n46_ & new_n286_;
  assign new_n288_ = new_n45_ & new_n287_;
  assign new_n289_ = new_n266_ & new_n288_;
  assign new_n290_ = ~new_n285_ & ~new_n289_;
  assign new_n291_ = ~new_n283_ & new_n290_;
  assign new_n292_ = ~A234 & A233;
  assign new_n293_ = new_n59_ & new_n292_;
  assign new_n294_ = new_n41_ & new_n293_;
  assign new_n295_ = new_n142_ & new_n294_;
  assign new_n296_ = A267 & A235;
  assign new_n297_ = new_n31_ & new_n296_;
  assign new_n298_ = new_n30_ & new_n297_;
  assign new_n299_ = new_n266_ & new_n298_;
  assign new_n300_ = new_n64_ & new_n297_;
  assign new_n301_ = new_n266_ & new_n300_;
  assign new_n302_ = ~new_n299_ & ~new_n301_;
  assign new_n303_ = ~new_n295_ & new_n302_;
  assign new_n304_ = new_n291_ & new_n303_;
  assign new_n305_ = new_n157_ & new_n294_;
  assign new_n306_ = new_n159_ & new_n294_;
  assign new_n307_ = new_n164_ & new_n294_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = ~new_n305_ & new_n308_;
  assign new_n310_ = new_n177_ & new_n294_;
  assign new_n311_ = new_n182_ & new_n294_;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign new_n313_ = new_n309_ & new_n312_;
  assign new_n314_ = new_n304_ & new_n313_;
  assign new_n315_ = new_n279_ & new_n314_;
  assign new_n316_ = new_n194_ & new_n294_;
  assign new_n317_ = new_n172_ & new_n294_;
  assign new_n318_ = new_n192_ & new_n294_;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = ~new_n316_ & new_n319_;
  assign new_n321_ = new_n203_ & new_n294_;
  assign new_n322_ = new_n188_ & new_n294_;
  assign new_n323_ = new_n201_ & new_n294_;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign new_n325_ = ~new_n321_ & new_n324_;
  assign new_n326_ = new_n320_ & new_n325_;
  assign new_n327_ = new_n211_ & new_n294_;
  assign new_n328_ = new_n199_ & new_n294_;
  assign new_n329_ = new_n207_ & new_n294_;
  assign new_n330_ = ~new_n328_ & ~new_n329_;
  assign new_n331_ = ~new_n327_ & new_n330_;
  assign new_n332_ = new_n220_ & new_n294_;
  assign new_n333_ = new_n222_ & new_n294_;
  assign new_n334_ = new_n224_ & new_n294_;
  assign new_n335_ = ~new_n333_ & ~new_n334_;
  assign new_n336_ = ~new_n332_ & new_n335_;
  assign new_n337_ = new_n331_ & new_n336_;
  assign new_n338_ = new_n326_ & new_n337_;
  assign new_n339_ = new_n234_ & new_n294_;
  assign new_n340_ = new_n238_ & new_n294_;
  assign new_n341_ = new_n240_ & new_n294_;
  assign new_n342_ = ~new_n340_ & ~new_n341_;
  assign new_n343_ = ~new_n339_ & new_n342_;
  assign new_n344_ = new_n249_ & new_n294_;
  assign new_n345_ = new_n253_ & new_n294_;
  assign new_n346_ = new_n257_ & new_n294_;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = ~new_n344_ & new_n347_;
  assign new_n349_ = new_n343_ & new_n348_;
  assign new_n350_ = A234 & A233;
  assign new_n351_ = new_n59_ & new_n350_;
  assign new_n352_ = new_n41_ & new_n351_;
  assign new_n353_ = new_n263_ & new_n352_;
  assign new_n354_ = new_n270_ & new_n352_;
  assign new_n355_ = new_n274_ & new_n352_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = ~new_n353_ & new_n356_;
  assign new_n358_ = new_n284_ & new_n352_;
  assign new_n359_ = new_n288_ & new_n352_;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = new_n357_ & new_n360_;
  assign new_n362_ = new_n349_ & new_n361_;
  assign new_n363_ = new_n338_ & new_n362_;
  assign new_n364_ = new_n315_ & new_n363_;
  assign new_n365_ = new_n217_ & new_n364_;
  assign new_n366_ = new_n300_ & new_n352_;
  assign new_n367_ = new_n282_ & new_n352_;
  assign new_n368_ = new_n298_ & new_n352_;
  assign new_n369_ = ~new_n367_ & ~new_n368_;
  assign new_n370_ = ~new_n366_ & new_n369_;
  assign new_n371_ = new_n71_ & new_n143_;
  assign new_n372_ = new_n74_ & new_n371_;
  assign new_n373_ = new_n164_ & new_n372_;
  assign new_n374_ = new_n142_ & new_n372_;
  assign new_n375_ = new_n159_ & new_n372_;
  assign new_n376_ = ~new_n374_ & ~new_n375_;
  assign new_n377_ = ~new_n373_ & new_n376_;
  assign new_n378_ = new_n370_ & new_n377_;
  assign new_n379_ = new_n182_ & new_n372_;
  assign new_n380_ = new_n157_ & new_n372_;
  assign new_n381_ = new_n177_ & new_n372_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = ~new_n379_ & new_n382_;
  assign new_n384_ = new_n194_ & new_n372_;
  assign new_n385_ = new_n172_ & new_n372_;
  assign new_n386_ = new_n192_ & new_n372_;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign new_n388_ = ~new_n384_ & new_n387_;
  assign new_n389_ = new_n383_ & new_n388_;
  assign new_n390_ = new_n378_ & new_n389_;
  assign new_n391_ = new_n203_ & new_n372_;
  assign new_n392_ = new_n188_ & new_n372_;
  assign new_n393_ = new_n201_ & new_n372_;
  assign new_n394_ = ~new_n392_ & ~new_n393_;
  assign new_n395_ = ~new_n391_ & new_n394_;
  assign new_n396_ = new_n211_ & new_n372_;
  assign new_n397_ = new_n199_ & new_n372_;
  assign new_n398_ = new_n207_ & new_n372_;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = ~new_n396_ & new_n399_;
  assign new_n401_ = new_n395_ & new_n400_;
  assign new_n402_ = new_n220_ & new_n372_;
  assign new_n403_ = new_n222_ & new_n372_;
  assign new_n404_ = new_n224_ & new_n372_;
  assign new_n405_ = ~new_n403_ & ~new_n404_;
  assign new_n406_ = ~new_n402_ & new_n405_;
  assign new_n407_ = new_n238_ & new_n372_;
  assign new_n408_ = new_n240_ & new_n372_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = new_n406_ & new_n409_;
  assign new_n411_ = new_n401_ & new_n410_;
  assign new_n412_ = new_n390_ & new_n411_;
  assign new_n413_ = new_n257_ & new_n372_;
  assign new_n414_ = new_n234_ & new_n372_;
  assign new_n415_ = new_n253_ & new_n372_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~new_n413_ & new_n416_;
  assign new_n418_ = new_n71_ & new_n264_;
  assign new_n419_ = new_n74_ & new_n418_;
  assign new_n420_ = new_n274_ & new_n419_;
  assign new_n421_ = new_n249_ & new_n372_;
  assign new_n422_ = new_n270_ & new_n419_;
  assign new_n423_ = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~new_n420_ & new_n423_;
  assign new_n425_ = new_n417_ & new_n424_;
  assign new_n426_ = new_n288_ & new_n419_;
  assign new_n427_ = new_n263_ & new_n419_;
  assign new_n428_ = new_n284_ & new_n419_;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = ~new_n426_ & new_n429_;
  assign new_n431_ = new_n300_ & new_n419_;
  assign new_n432_ = new_n282_ & new_n419_;
  assign new_n433_ = new_n298_ & new_n419_;
  assign new_n434_ = ~new_n432_ & ~new_n433_;
  assign new_n435_ = ~new_n431_ & new_n434_;
  assign new_n436_ = new_n430_ & new_n435_;
  assign new_n437_ = new_n425_ & new_n436_;
  assign new_n438_ = new_n88_ & new_n292_;
  assign new_n439_ = new_n74_ & new_n438_;
  assign new_n440_ = new_n164_ & new_n439_;
  assign new_n441_ = new_n142_ & new_n439_;
  assign new_n442_ = new_n159_ & new_n439_;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign new_n444_ = ~new_n440_ & new_n443_;
  assign new_n445_ = new_n182_ & new_n439_;
  assign new_n446_ = new_n157_ & new_n439_;
  assign new_n447_ = new_n177_ & new_n439_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = ~new_n445_ & new_n448_;
  assign new_n450_ = new_n444_ & new_n449_;
  assign new_n451_ = new_n194_ & new_n439_;
  assign new_n452_ = new_n172_ & new_n439_;
  assign new_n453_ = new_n192_ & new_n439_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~new_n451_ & new_n454_;
  assign new_n456_ = new_n188_ & new_n439_;
  assign new_n457_ = new_n201_ & new_n439_;
  assign new_n458_ = ~new_n456_ & ~new_n457_;
  assign new_n459_ = new_n455_ & new_n458_;
  assign new_n460_ = new_n450_ & new_n459_;
  assign new_n461_ = new_n437_ & new_n460_;
  assign new_n462_ = new_n412_ & new_n461_;
  assign new_n463_ = new_n207_ & new_n439_;
  assign new_n464_ = new_n203_ & new_n439_;
  assign new_n465_ = new_n199_ & new_n439_;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign new_n467_ = ~new_n463_ & new_n466_;
  assign new_n468_ = new_n224_ & new_n439_;
  assign new_n469_ = new_n211_ & new_n439_;
  assign new_n470_ = new_n222_ & new_n439_;
  assign new_n471_ = ~new_n469_ & ~new_n470_;
  assign new_n472_ = ~new_n468_ & new_n471_;
  assign new_n473_ = new_n467_ & new_n472_;
  assign new_n474_ = new_n240_ & new_n439_;
  assign new_n475_ = new_n220_ & new_n439_;
  assign new_n476_ = new_n238_ & new_n439_;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign new_n478_ = ~new_n474_ & new_n477_;
  assign new_n479_ = new_n257_ & new_n439_;
  assign new_n480_ = new_n234_ & new_n439_;
  assign new_n481_ = new_n253_ & new_n439_;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = ~new_n479_ & new_n482_;
  assign new_n484_ = new_n478_ & new_n483_;
  assign new_n485_ = new_n473_ & new_n484_;
  assign new_n486_ = new_n88_ & new_n350_;
  assign new_n487_ = new_n74_ & new_n486_;
  assign new_n488_ = new_n274_ & new_n487_;
  assign new_n489_ = new_n249_ & new_n439_;
  assign new_n490_ = new_n270_ & new_n487_;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = ~new_n488_ & new_n491_;
  assign new_n493_ = new_n288_ & new_n487_;
  assign new_n494_ = new_n263_ & new_n487_;
  assign new_n495_ = new_n284_ & new_n487_;
  assign new_n496_ = ~new_n494_ & ~new_n495_;
  assign new_n497_ = ~new_n493_ & new_n496_;
  assign new_n498_ = new_n492_ & new_n497_;
  assign new_n499_ = new_n300_ & new_n487_;
  assign new_n500_ = new_n282_ & new_n487_;
  assign new_n501_ = new_n298_ & new_n487_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n499_ & new_n502_;
  assign new_n504_ = ~A235 & A234;
  assign new_n505_ = A203 & ~A202;
  assign new_n506_ = new_n504_ & new_n505_;
  assign new_n507_ = A201 & A168;
  assign new_n508_ = new_n40_ & new_n507_;
  assign new_n509_ = new_n506_ & new_n508_;
  assign new_n510_ = new_n49_ & new_n509_;
  assign new_n511_ = new_n54_ & new_n509_;
  assign new_n512_ = ~new_n510_ & ~new_n511_;
  assign new_n513_ = new_n503_ & new_n512_;
  assign new_n514_ = new_n498_ & new_n513_;
  assign new_n515_ = new_n485_ & new_n514_;
  assign new_n516_ = ~A233 & A232;
  assign new_n517_ = new_n35_ & new_n516_;
  assign new_n518_ = A166 & ~A167;
  assign new_n519_ = A168 & A169;
  assign new_n520_ = new_n518_ & new_n519_;
  assign new_n521_ = new_n517_ & new_n520_;
  assign new_n522_ = new_n49_ & new_n521_;
  assign new_n523_ = new_n34_ & new_n509_;
  assign new_n524_ = new_n65_ & new_n509_;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign new_n526_ = ~new_n522_ & new_n525_;
  assign new_n527_ = new_n65_ & new_n521_;
  assign new_n528_ = new_n54_ & new_n521_;
  assign new_n529_ = new_n34_ & new_n521_;
  assign new_n530_ = ~new_n528_ & ~new_n529_;
  assign new_n531_ = ~new_n527_ & new_n530_;
  assign new_n532_ = new_n526_ & new_n531_;
  assign new_n533_ = A233 & ~A232;
  assign new_n534_ = new_n35_ & new_n533_;
  assign new_n535_ = new_n520_ & new_n534_;
  assign new_n536_ = new_n34_ & new_n535_;
  assign new_n537_ = new_n49_ & new_n535_;
  assign new_n538_ = new_n54_ & new_n535_;
  assign new_n539_ = ~new_n537_ & ~new_n538_;
  assign new_n540_ = ~new_n536_ & new_n539_;
  assign new_n541_ = ~A166 & A167;
  assign new_n542_ = new_n519_ & new_n541_;
  assign new_n543_ = new_n517_ & new_n542_;
  assign new_n544_ = new_n54_ & new_n543_;
  assign new_n545_ = new_n65_ & new_n535_;
  assign new_n546_ = new_n49_ & new_n543_;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = ~new_n544_ & new_n547_;
  assign new_n549_ = new_n540_ & new_n548_;
  assign new_n550_ = new_n532_ & new_n549_;
  assign new_n551_ = new_n534_ & new_n542_;
  assign new_n552_ = new_n49_ & new_n551_;
  assign new_n553_ = new_n34_ & new_n543_;
  assign new_n554_ = new_n65_ & new_n543_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = ~new_n552_ & new_n555_;
  assign new_n557_ = new_n65_ & new_n551_;
  assign new_n558_ = new_n54_ & new_n551_;
  assign new_n559_ = new_n34_ & new_n551_;
  assign new_n560_ = ~new_n558_ & ~new_n559_;
  assign new_n561_ = ~new_n557_ & new_n560_;
  assign new_n562_ = new_n556_ & new_n561_;
  assign new_n563_ = A168 & A170;
  assign new_n564_ = new_n518_ & new_n563_;
  assign new_n565_ = new_n517_ & new_n564_;
  assign new_n566_ = new_n34_ & new_n565_;
  assign new_n567_ = new_n49_ & new_n565_;
  assign new_n568_ = new_n54_ & new_n565_;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = ~new_n566_ & new_n569_;
  assign new_n571_ = new_n65_ & new_n565_;
  assign new_n572_ = new_n534_ & new_n564_;
  assign new_n573_ = new_n49_ & new_n572_;
  assign new_n574_ = ~new_n571_ & ~new_n573_;
  assign new_n575_ = new_n570_ & new_n574_;
  assign new_n576_ = new_n562_ & new_n575_;
  assign new_n577_ = new_n550_ & new_n576_;
  assign new_n578_ = new_n515_ & new_n577_;
  assign new_n579_ = new_n462_ & new_n578_;
  assign new_n580_ = new_n365_ & new_n579_;
  assign new_n581_ = new_n65_ & new_n572_;
  assign new_n582_ = new_n54_ & new_n572_;
  assign new_n583_ = new_n34_ & new_n572_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = ~new_n581_ & new_n584_;
  assign new_n586_ = new_n541_ & new_n563_;
  assign new_n587_ = new_n517_ & new_n586_;
  assign new_n588_ = new_n34_ & new_n587_;
  assign new_n589_ = new_n49_ & new_n587_;
  assign new_n590_ = new_n54_ & new_n587_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~new_n588_ & new_n591_;
  assign new_n593_ = new_n585_ & new_n592_;
  assign new_n594_ = new_n534_ & new_n586_;
  assign new_n595_ = new_n54_ & new_n594_;
  assign new_n596_ = new_n65_ & new_n587_;
  assign new_n597_ = new_n49_ & new_n594_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~new_n595_ & new_n598_;
  assign new_n600_ = new_n96_ & new_n143_;
  assign new_n601_ = new_n100_ & new_n600_;
  assign new_n602_ = new_n142_ & new_n601_;
  assign new_n603_ = new_n34_ & new_n594_;
  assign new_n604_ = new_n65_ & new_n594_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n602_ & new_n605_;
  assign new_n607_ = new_n599_ & new_n606_;
  assign new_n608_ = new_n593_ & new_n607_;
  assign new_n609_ = new_n157_ & new_n601_;
  assign new_n610_ = new_n159_ & new_n601_;
  assign new_n611_ = new_n164_ & new_n601_;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = ~new_n609_ & new_n612_;
  assign new_n614_ = new_n172_ & new_n601_;
  assign new_n615_ = new_n177_ & new_n601_;
  assign new_n616_ = new_n182_ & new_n601_;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = ~new_n614_ & new_n617_;
  assign new_n619_ = new_n613_ & new_n618_;
  assign new_n620_ = new_n188_ & new_n601_;
  assign new_n621_ = new_n192_ & new_n601_;
  assign new_n622_ = new_n194_ & new_n601_;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_ = ~new_n620_ & new_n623_;
  assign new_n625_ = new_n199_ & new_n601_;
  assign new_n626_ = new_n201_ & new_n601_;
  assign new_n627_ = new_n203_ & new_n601_;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = ~new_n625_ & new_n628_;
  assign new_n630_ = new_n624_ & new_n629_;
  assign new_n631_ = new_n619_ & new_n630_;
  assign new_n632_ = new_n608_ & new_n631_;
  assign new_n633_ = new_n222_ & new_n601_;
  assign new_n634_ = new_n207_ & new_n601_;
  assign new_n635_ = new_n211_ & new_n601_;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = ~new_n633_ & new_n636_;
  assign new_n638_ = new_n238_ & new_n601_;
  assign new_n639_ = new_n224_ & new_n601_;
  assign new_n640_ = new_n220_ & new_n601_;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n638_ & new_n641_;
  assign new_n643_ = new_n637_ & new_n642_;
  assign new_n644_ = new_n253_ & new_n601_;
  assign new_n645_ = new_n240_ & new_n601_;
  assign new_n646_ = new_n234_ & new_n601_;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = ~new_n644_ & new_n647_;
  assign new_n649_ = new_n96_ & new_n264_;
  assign new_n650_ = new_n100_ & new_n649_;
  assign new_n651_ = new_n270_ & new_n650_;
  assign new_n652_ = new_n257_ & new_n601_;
  assign new_n653_ = new_n249_ & new_n601_;
  assign new_n654_ = ~new_n652_ & ~new_n653_;
  assign new_n655_ = ~new_n651_ & new_n654_;
  assign new_n656_ = new_n648_ & new_n655_;
  assign new_n657_ = new_n643_ & new_n656_;
  assign new_n658_ = new_n284_ & new_n650_;
  assign new_n659_ = new_n274_ & new_n650_;
  assign new_n660_ = new_n263_ & new_n650_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = ~new_n658_ & new_n661_;
  assign new_n663_ = new_n298_ & new_n650_;
  assign new_n664_ = new_n288_ & new_n650_;
  assign new_n665_ = new_n282_ & new_n650_;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = ~new_n663_ & new_n666_;
  assign new_n668_ = new_n662_ & new_n667_;
  assign new_n669_ = new_n108_ & new_n292_;
  assign new_n670_ = new_n100_ & new_n669_;
  assign new_n671_ = new_n159_ & new_n670_;
  assign new_n672_ = new_n300_ & new_n650_;
  assign new_n673_ = new_n142_ & new_n670_;
  assign new_n674_ = ~new_n672_ & ~new_n673_;
  assign new_n675_ = ~new_n671_ & new_n674_;
  assign new_n676_ = new_n164_ & new_n670_;
  assign new_n677_ = new_n157_ & new_n670_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = new_n675_ & new_n678_;
  assign new_n680_ = new_n668_ & new_n679_;
  assign new_n681_ = new_n657_ & new_n680_;
  assign new_n682_ = new_n632_ & new_n681_;
  assign new_n683_ = new_n172_ & new_n670_;
  assign new_n684_ = new_n177_ & new_n670_;
  assign new_n685_ = new_n182_ & new_n670_;
  assign new_n686_ = ~new_n684_ & ~new_n685_;
  assign new_n687_ = ~new_n683_ & new_n686_;
  assign new_n688_ = new_n188_ & new_n670_;
  assign new_n689_ = new_n192_ & new_n670_;
  assign new_n690_ = new_n194_ & new_n670_;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = ~new_n688_ & new_n691_;
  assign new_n693_ = new_n687_ & new_n692_;
  assign new_n694_ = new_n199_ & new_n670_;
  assign new_n695_ = new_n201_ & new_n670_;
  assign new_n696_ = new_n203_ & new_n670_;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~new_n694_ & new_n697_;
  assign new_n699_ = new_n222_ & new_n670_;
  assign new_n700_ = new_n207_ & new_n670_;
  assign new_n701_ = new_n211_ & new_n670_;
  assign new_n702_ = ~new_n700_ & ~new_n701_;
  assign new_n703_ = ~new_n699_ & new_n702_;
  assign new_n704_ = new_n698_ & new_n703_;
  assign new_n705_ = new_n693_ & new_n704_;
  assign new_n706_ = new_n238_ & new_n670_;
  assign new_n707_ = new_n224_ & new_n670_;
  assign new_n708_ = new_n220_ & new_n670_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = ~new_n706_ & new_n709_;
  assign new_n711_ = new_n253_ & new_n670_;
  assign new_n712_ = new_n240_ & new_n670_;
  assign new_n713_ = new_n234_ & new_n670_;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = ~new_n711_ & new_n714_;
  assign new_n716_ = new_n710_ & new_n715_;
  assign new_n717_ = new_n108_ & new_n350_;
  assign new_n718_ = new_n100_ & new_n717_;
  assign new_n719_ = new_n270_ & new_n718_;
  assign new_n720_ = new_n257_ & new_n670_;
  assign new_n721_ = new_n249_ & new_n670_;
  assign new_n722_ = ~new_n720_ & ~new_n721_;
  assign new_n723_ = ~new_n719_ & new_n722_;
  assign new_n724_ = new_n274_ & new_n718_;
  assign new_n725_ = new_n263_ & new_n718_;
  assign new_n726_ = ~new_n724_ & ~new_n725_;
  assign new_n727_ = new_n723_ & new_n726_;
  assign new_n728_ = new_n716_ & new_n727_;
  assign new_n729_ = new_n705_ & new_n728_;
  assign new_n730_ = new_n282_ & new_n718_;
  assign new_n731_ = new_n284_ & new_n718_;
  assign new_n732_ = new_n288_ & new_n718_;
  assign new_n733_ = ~new_n731_ & ~new_n732_;
  assign new_n734_ = ~new_n730_ & new_n733_;
  assign new_n735_ = ~A203 & A201;
  assign new_n736_ = new_n99_ & new_n735_;
  assign new_n737_ = new_n517_ & new_n736_;
  assign new_n738_ = new_n49_ & new_n737_;
  assign new_n739_ = new_n298_ & new_n718_;
  assign new_n740_ = new_n300_ & new_n718_;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = ~new_n738_ & new_n741_;
  assign new_n743_ = new_n734_ & new_n742_;
  assign new_n744_ = new_n65_ & new_n737_;
  assign new_n745_ = new_n54_ & new_n737_;
  assign new_n746_ = new_n34_ & new_n737_;
  assign new_n747_ = ~new_n745_ & ~new_n746_;
  assign new_n748_ = ~new_n744_ & new_n747_;
  assign new_n749_ = new_n534_ & new_n736_;
  assign new_n750_ = new_n34_ & new_n749_;
  assign new_n751_ = new_n49_ & new_n749_;
  assign new_n752_ = new_n54_ & new_n749_;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = ~new_n750_ & new_n753_;
  assign new_n755_ = new_n748_ & new_n754_;
  assign new_n756_ = new_n743_ & new_n755_;
  assign new_n757_ = A202 & A201;
  assign new_n758_ = new_n99_ & new_n757_;
  assign new_n759_ = new_n517_ & new_n758_;
  assign new_n760_ = new_n54_ & new_n759_;
  assign new_n761_ = new_n65_ & new_n749_;
  assign new_n762_ = new_n49_ & new_n759_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = ~new_n760_ & new_n763_;
  assign new_n765_ = new_n534_ & new_n758_;
  assign new_n766_ = new_n49_ & new_n765_;
  assign new_n767_ = new_n34_ & new_n759_;
  assign new_n768_ = new_n65_ & new_n759_;
  assign new_n769_ = ~new_n767_ & ~new_n768_;
  assign new_n770_ = ~new_n766_ & new_n769_;
  assign new_n771_ = new_n764_ & new_n770_;
  assign new_n772_ = new_n65_ & new_n765_;
  assign new_n773_ = new_n54_ & new_n765_;
  assign new_n774_ = new_n34_ & new_n765_;
  assign new_n775_ = ~new_n773_ & ~new_n774_;
  assign new_n776_ = ~new_n772_ & new_n775_;
  assign new_n777_ = new_n125_ & new_n600_;
  assign new_n778_ = new_n142_ & new_n777_;
  assign new_n779_ = new_n159_ & new_n777_;
  assign new_n780_ = ~new_n778_ & ~new_n779_;
  assign new_n781_ = new_n776_ & new_n780_;
  assign new_n782_ = new_n771_ & new_n781_;
  assign new_n783_ = new_n756_ & new_n782_;
  assign new_n784_ = new_n729_ & new_n783_;
  assign new_n785_ = new_n682_ & new_n784_;
  assign new_n786_ = new_n177_ & new_n777_;
  assign new_n787_ = new_n164_ & new_n777_;
  assign new_n788_ = new_n157_ & new_n777_;
  assign new_n789_ = ~new_n787_ & ~new_n788_;
  assign new_n790_ = ~new_n786_ & new_n789_;
  assign new_n791_ = new_n192_ & new_n777_;
  assign new_n792_ = new_n182_ & new_n777_;
  assign new_n793_ = new_n172_ & new_n777_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = ~new_n791_ & new_n794_;
  assign new_n796_ = new_n790_ & new_n795_;
  assign new_n797_ = new_n201_ & new_n777_;
  assign new_n798_ = new_n194_ & new_n777_;
  assign new_n799_ = new_n188_ & new_n777_;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = ~new_n797_ & new_n800_;
  assign new_n802_ = new_n207_ & new_n777_;
  assign new_n803_ = new_n203_ & new_n777_;
  assign new_n804_ = new_n199_ & new_n777_;
  assign new_n805_ = ~new_n803_ & ~new_n804_;
  assign new_n806_ = ~new_n802_ & new_n805_;
  assign new_n807_ = new_n801_ & new_n806_;
  assign new_n808_ = new_n796_ & new_n807_;
  assign new_n809_ = new_n224_ & new_n777_;
  assign new_n810_ = new_n211_ & new_n777_;
  assign new_n811_ = new_n222_ & new_n777_;
  assign new_n812_ = ~new_n810_ & ~new_n811_;
  assign new_n813_ = ~new_n809_ & new_n812_;
  assign new_n814_ = new_n240_ & new_n777_;
  assign new_n815_ = new_n220_ & new_n777_;
  assign new_n816_ = new_n238_ & new_n777_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~new_n814_ & new_n817_;
  assign new_n819_ = new_n813_ & new_n818_;
  assign new_n820_ = new_n257_ & new_n777_;
  assign new_n821_ = new_n234_ & new_n777_;
  assign new_n822_ = new_n253_ & new_n777_;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = ~new_n820_ & new_n823_;
  assign new_n825_ = new_n249_ & new_n777_;
  assign new_n826_ = new_n125_ & new_n649_;
  assign new_n827_ = new_n270_ & new_n826_;
  assign new_n828_ = ~new_n825_ & ~new_n827_;
  assign new_n829_ = new_n824_ & new_n828_;
  assign new_n830_ = new_n819_ & new_n829_;
  assign new_n831_ = new_n808_ & new_n830_;
  assign new_n832_ = new_n284_ & new_n826_;
  assign new_n833_ = new_n274_ & new_n826_;
  assign new_n834_ = new_n263_ & new_n826_;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = ~new_n832_ & new_n835_;
  assign new_n837_ = new_n298_ & new_n826_;
  assign new_n838_ = new_n288_ & new_n826_;
  assign new_n839_ = new_n282_ & new_n826_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = ~new_n837_ & new_n840_;
  assign new_n842_ = new_n836_ & new_n841_;
  assign new_n843_ = new_n125_ & new_n669_;
  assign new_n844_ = new_n159_ & new_n843_;
  assign new_n845_ = new_n300_ & new_n826_;
  assign new_n846_ = new_n142_ & new_n843_;
  assign new_n847_ = ~new_n845_ & ~new_n846_;
  assign new_n848_ = ~new_n844_ & new_n847_;
  assign new_n849_ = new_n177_ & new_n843_;
  assign new_n850_ = new_n164_ & new_n843_;
  assign new_n851_ = new_n157_ & new_n843_;
  assign new_n852_ = ~new_n850_ & ~new_n851_;
  assign new_n853_ = ~new_n849_ & new_n852_;
  assign new_n854_ = new_n848_ & new_n853_;
  assign new_n855_ = new_n842_ & new_n854_;
  assign new_n856_ = new_n192_ & new_n843_;
  assign new_n857_ = new_n182_ & new_n843_;
  assign new_n858_ = new_n172_ & new_n843_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~new_n856_ & new_n859_;
  assign new_n861_ = new_n201_ & new_n843_;
  assign new_n862_ = new_n194_ & new_n843_;
  assign new_n863_ = new_n188_ & new_n843_;
  assign new_n864_ = ~new_n862_ & ~new_n863_;
  assign new_n865_ = ~new_n861_ & new_n864_;
  assign new_n866_ = new_n860_ & new_n865_;
  assign new_n867_ = new_n207_ & new_n843_;
  assign new_n868_ = new_n203_ & new_n843_;
  assign new_n869_ = new_n199_ & new_n843_;
  assign new_n870_ = ~new_n868_ & ~new_n869_;
  assign new_n871_ = ~new_n867_ & new_n870_;
  assign new_n872_ = new_n211_ & new_n843_;
  assign new_n873_ = new_n222_ & new_n843_;
  assign new_n874_ = ~new_n872_ & ~new_n873_;
  assign new_n875_ = new_n871_ & new_n874_;
  assign new_n876_ = new_n866_ & new_n875_;
  assign new_n877_ = new_n855_ & new_n876_;
  assign new_n878_ = new_n831_ & new_n877_;
  assign new_n879_ = new_n238_ & new_n843_;
  assign new_n880_ = new_n224_ & new_n843_;
  assign new_n881_ = new_n220_ & new_n843_;
  assign new_n882_ = ~new_n880_ & ~new_n881_;
  assign new_n883_ = ~new_n879_ & new_n882_;
  assign new_n884_ = new_n253_ & new_n843_;
  assign new_n885_ = new_n240_ & new_n843_;
  assign new_n886_ = new_n234_ & new_n843_;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = ~new_n884_ & new_n887_;
  assign new_n889_ = new_n883_ & new_n888_;
  assign new_n890_ = new_n125_ & new_n717_;
  assign new_n891_ = new_n270_ & new_n890_;
  assign new_n892_ = new_n257_ & new_n843_;
  assign new_n893_ = new_n249_ & new_n843_;
  assign new_n894_ = ~new_n892_ & ~new_n893_;
  assign new_n895_ = ~new_n891_ & new_n894_;
  assign new_n896_ = new_n284_ & new_n890_;
  assign new_n897_ = new_n274_ & new_n890_;
  assign new_n898_ = new_n263_ & new_n890_;
  assign new_n899_ = ~new_n897_ & ~new_n898_;
  assign new_n900_ = ~new_n896_ & new_n899_;
  assign new_n901_ = new_n895_ & new_n900_;
  assign new_n902_ = new_n889_ & new_n901_;
  assign new_n903_ = new_n298_ & new_n890_;
  assign new_n904_ = new_n288_ & new_n890_;
  assign new_n905_ = new_n282_ & new_n890_;
  assign new_n906_ = ~new_n904_ & ~new_n905_;
  assign new_n907_ = ~new_n903_ & new_n906_;
  assign new_n908_ = new_n124_ & new_n735_;
  assign new_n909_ = new_n517_ & new_n908_;
  assign new_n910_ = new_n54_ & new_n909_;
  assign new_n911_ = new_n300_ & new_n890_;
  assign new_n912_ = new_n49_ & new_n909_;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = ~new_n910_ & new_n913_;
  assign new_n915_ = new_n907_ & new_n914_;
  assign new_n916_ = new_n534_ & new_n908_;
  assign new_n917_ = new_n49_ & new_n916_;
  assign new_n918_ = new_n34_ & new_n909_;
  assign new_n919_ = new_n65_ & new_n909_;
  assign new_n920_ = ~new_n918_ & ~new_n919_;
  assign new_n921_ = ~new_n917_ & new_n920_;
  assign new_n922_ = new_n54_ & new_n916_;
  assign new_n923_ = new_n34_ & new_n916_;
  assign new_n924_ = ~new_n922_ & ~new_n923_;
  assign new_n925_ = new_n921_ & new_n924_;
  assign new_n926_ = new_n915_ & new_n925_;
  assign new_n927_ = new_n902_ & new_n926_;
  assign new_n928_ = new_n124_ & new_n757_;
  assign new_n929_ = new_n517_ & new_n928_;
  assign new_n930_ = new_n54_ & new_n929_;
  assign new_n931_ = new_n65_ & new_n916_;
  assign new_n932_ = new_n49_ & new_n929_;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign new_n934_ = ~new_n930_ & new_n933_;
  assign new_n935_ = new_n534_ & new_n928_;
  assign new_n936_ = new_n49_ & new_n935_;
  assign new_n937_ = new_n34_ & new_n929_;
  assign new_n938_ = new_n65_ & new_n929_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = ~new_n936_ & new_n939_;
  assign new_n941_ = new_n934_ & new_n940_;
  assign new_n942_ = new_n65_ & new_n935_;
  assign new_n943_ = new_n54_ & new_n935_;
  assign new_n944_ = new_n34_ & new_n935_;
  assign new_n945_ = ~new_n943_ & ~new_n944_;
  assign new_n946_ = ~new_n942_ & new_n945_;
  assign new_n947_ = new_n63_ & new_n228_;
  assign new_n948_ = new_n141_ & new_n947_;
  assign new_n949_ = new_n145_ & new_n948_;
  assign new_n950_ = new_n29_ & new_n228_;
  assign new_n951_ = new_n141_ & new_n950_;
  assign new_n952_ = new_n145_ & new_n951_;
  assign new_n953_ = new_n29_ & new_n245_;
  assign new_n954_ = new_n141_ & new_n953_;
  assign new_n955_ = new_n145_ & new_n954_;
  assign new_n956_ = ~new_n952_ & ~new_n955_;
  assign new_n957_ = ~new_n949_ & new_n956_;
  assign new_n958_ = new_n946_ & new_n957_;
  assign new_n959_ = new_n941_ & new_n958_;
  assign new_n960_ = new_n151_ & new_n170_;
  assign new_n961_ = new_n156_ & new_n960_;
  assign new_n962_ = new_n145_ & new_n961_;
  assign new_n963_ = new_n63_ & new_n245_;
  assign new_n964_ = new_n141_ & new_n963_;
  assign new_n965_ = new_n145_ & new_n964_;
  assign new_n966_ = new_n161_ & new_n170_;
  assign new_n967_ = new_n156_ & new_n966_;
  assign new_n968_ = new_n145_ & new_n967_;
  assign new_n969_ = ~new_n965_ & ~new_n968_;
  assign new_n970_ = ~new_n962_ & new_n969_;
  assign new_n971_ = new_n161_ & new_n190_;
  assign new_n972_ = new_n156_ & new_n971_;
  assign new_n973_ = new_n145_ & new_n972_;
  assign new_n974_ = new_n170_ & new_n174_;
  assign new_n975_ = new_n156_ & new_n974_;
  assign new_n976_ = new_n145_ & new_n975_;
  assign new_n977_ = new_n170_ & new_n179_;
  assign new_n978_ = new_n156_ & new_n977_;
  assign new_n979_ = new_n145_ & new_n978_;
  assign new_n980_ = ~new_n976_ & ~new_n979_;
  assign new_n981_ = ~new_n973_ & new_n980_;
  assign new_n982_ = new_n970_ & new_n981_;
  assign new_n983_ = new_n179_ & new_n190_;
  assign new_n984_ = new_n156_ & new_n983_;
  assign new_n985_ = new_n145_ & new_n984_;
  assign new_n986_ = new_n151_ & new_n190_;
  assign new_n987_ = new_n156_ & new_n986_;
  assign new_n988_ = new_n145_ & new_n987_;
  assign new_n989_ = new_n174_ & new_n190_;
  assign new_n990_ = new_n156_ & new_n989_;
  assign new_n991_ = new_n145_ & new_n990_;
  assign new_n992_ = ~new_n988_ & ~new_n991_;
  assign new_n993_ = ~new_n985_ & new_n992_;
  assign new_n994_ = new_n187_ & new_n966_;
  assign new_n995_ = new_n145_ & new_n994_;
  assign new_n996_ = new_n187_ & new_n960_;
  assign new_n997_ = new_n145_ & new_n996_;
  assign new_n998_ = ~new_n995_ & ~new_n997_;
  assign new_n999_ = new_n993_ & new_n998_;
  assign new_n1000_ = new_n982_ & new_n999_;
  assign new_n1001_ = new_n959_ & new_n1000_;
  assign new_n1002_ = new_n927_ & new_n1001_;
  assign new_n1003_ = new_n878_ & new_n1002_;
  assign new_n1004_ = new_n785_ & new_n1003_;
  assign new_n1005_ = new_n580_ & new_n1004_;
  assign new_n1006_ = new_n187_ & new_n971_;
  assign new_n1007_ = new_n145_ & new_n1006_;
  assign new_n1008_ = new_n187_ & new_n974_;
  assign new_n1009_ = new_n145_ & new_n1008_;
  assign new_n1010_ = new_n187_ & new_n977_;
  assign new_n1011_ = new_n145_ & new_n1010_;
  assign new_n1012_ = ~new_n1009_ & ~new_n1011_;
  assign new_n1013_ = ~new_n1007_ & new_n1012_;
  assign new_n1014_ = new_n187_ & new_n983_;
  assign new_n1015_ = new_n145_ & new_n1014_;
  assign new_n1016_ = new_n187_ & new_n986_;
  assign new_n1017_ = new_n145_ & new_n1016_;
  assign new_n1018_ = new_n187_ & new_n989_;
  assign new_n1019_ = new_n145_ & new_n1018_;
  assign new_n1020_ = ~new_n1017_ & ~new_n1019_;
  assign new_n1021_ = ~new_n1015_ & new_n1020_;
  assign new_n1022_ = new_n1013_ & new_n1021_;
  assign new_n1023_ = new_n210_ & new_n947_;
  assign new_n1024_ = new_n145_ & new_n1023_;
  assign new_n1025_ = new_n210_ & new_n950_;
  assign new_n1026_ = new_n145_ & new_n1025_;
  assign new_n1027_ = new_n210_ & new_n953_;
  assign new_n1028_ = new_n145_ & new_n1027_;
  assign new_n1029_ = ~new_n1026_ & ~new_n1028_;
  assign new_n1030_ = ~new_n1024_ & new_n1029_;
  assign new_n1031_ = new_n219_ & new_n953_;
  assign new_n1032_ = new_n145_ & new_n1031_;
  assign new_n1033_ = new_n210_ & new_n963_;
  assign new_n1034_ = new_n145_ & new_n1033_;
  assign new_n1035_ = new_n219_ & new_n950_;
  assign new_n1036_ = new_n145_ & new_n1035_;
  assign new_n1037_ = ~new_n1034_ & ~new_n1036_;
  assign new_n1038_ = ~new_n1032_ & new_n1037_;
  assign new_n1039_ = new_n1030_ & new_n1038_;
  assign new_n1040_ = new_n1022_ & new_n1039_;
  assign new_n1041_ = new_n237_ & new_n950_;
  assign new_n1042_ = new_n145_ & new_n1041_;
  assign new_n1043_ = new_n219_ & new_n947_;
  assign new_n1044_ = new_n145_ & new_n1043_;
  assign new_n1045_ = new_n219_ & new_n963_;
  assign new_n1046_ = new_n145_ & new_n1045_;
  assign new_n1047_ = ~new_n1044_ & ~new_n1046_;
  assign new_n1048_ = ~new_n1042_ & new_n1047_;
  assign new_n1049_ = new_n237_ & new_n963_;
  assign new_n1050_ = new_n145_ & new_n1049_;
  assign new_n1051_ = new_n237_ & new_n953_;
  assign new_n1052_ = new_n145_ & new_n1051_;
  assign new_n1053_ = new_n237_ & new_n947_;
  assign new_n1054_ = new_n145_ & new_n1053_;
  assign new_n1055_ = ~new_n1052_ & ~new_n1054_;
  assign new_n1056_ = ~new_n1050_ & new_n1055_;
  assign new_n1057_ = new_n1048_ & new_n1056_;
  assign new_n1058_ = new_n31_ & new_n161_;
  assign new_n1059_ = new_n269_ & new_n1058_;
  assign new_n1060_ = new_n266_ & new_n1059_;
  assign new_n1061_ = ~A300 & A299;
  assign new_n1062_ = new_n27_ & new_n1061_;
  assign new_n1063_ = ~A298 & ~A266;
  assign new_n1064_ = new_n272_ & new_n1063_;
  assign new_n1065_ = new_n1062_ & new_n1064_;
  assign new_n1066_ = new_n266_ & new_n1065_;
  assign new_n1067_ = ~A300 & ~A299;
  assign new_n1068_ = new_n27_ & new_n1067_;
  assign new_n1069_ = A298 & ~A266;
  assign new_n1070_ = new_n272_ & new_n1069_;
  assign new_n1071_ = new_n1068_ & new_n1070_;
  assign new_n1072_ = new_n266_ & new_n1071_;
  assign new_n1073_ = ~new_n1066_ & ~new_n1072_;
  assign new_n1074_ = ~new_n1060_ & new_n1073_;
  assign new_n1075_ = new_n31_ & new_n179_;
  assign new_n1076_ = new_n269_ & new_n1075_;
  assign new_n1077_ = new_n266_ & new_n1076_;
  assign new_n1078_ = new_n31_ & new_n151_;
  assign new_n1079_ = new_n269_ & new_n1078_;
  assign new_n1080_ = new_n266_ & new_n1079_;
  assign new_n1081_ = new_n31_ & new_n174_;
  assign new_n1082_ = new_n269_ & new_n1081_;
  assign new_n1083_ = new_n266_ & new_n1082_;
  assign new_n1084_ = ~new_n1080_ & ~new_n1083_;
  assign new_n1085_ = ~new_n1077_ & new_n1084_;
  assign new_n1086_ = new_n1074_ & new_n1085_;
  assign new_n1087_ = new_n1057_ & new_n1086_;
  assign new_n1088_ = new_n1040_ & new_n1087_;
  assign new_n1089_ = new_n273_ & new_n1058_;
  assign new_n1090_ = new_n266_ & new_n1089_;
  assign new_n1091_ = A300 & ~A269;
  assign new_n1092_ = new_n27_ & new_n1091_;
  assign new_n1093_ = A267 & ~A266;
  assign new_n1094_ = new_n268_ & new_n1093_;
  assign new_n1095_ = new_n1092_ & new_n1094_;
  assign new_n1096_ = new_n266_ & new_n1095_;
  assign new_n1097_ = A300 & A268;
  assign new_n1098_ = new_n27_ & new_n1097_;
  assign new_n1099_ = new_n1094_ & new_n1098_;
  assign new_n1100_ = new_n266_ & new_n1099_;
  assign new_n1101_ = ~new_n1096_ & ~new_n1100_;
  assign new_n1102_ = ~new_n1090_ & new_n1101_;
  assign new_n1103_ = new_n273_ & new_n1075_;
  assign new_n1104_ = new_n266_ & new_n1103_;
  assign new_n1105_ = new_n273_ & new_n1078_;
  assign new_n1106_ = new_n266_ & new_n1105_;
  assign new_n1107_ = new_n273_ & new_n1081_;
  assign new_n1108_ = new_n266_ & new_n1107_;
  assign new_n1109_ = ~new_n1106_ & ~new_n1108_;
  assign new_n1110_ = ~new_n1104_ & new_n1109_;
  assign new_n1111_ = new_n1102_ & new_n1110_;
  assign new_n1112_ = ~A298 & A266;
  assign new_n1113_ = new_n268_ & new_n1112_;
  assign new_n1114_ = new_n1062_ & new_n1113_;
  assign new_n1115_ = new_n266_ & new_n1114_;
  assign new_n1116_ = A267 & A266;
  assign new_n1117_ = new_n272_ & new_n1116_;
  assign new_n1118_ = new_n1092_ & new_n1117_;
  assign new_n1119_ = new_n266_ & new_n1118_;
  assign new_n1120_ = new_n1098_ & new_n1117_;
  assign new_n1121_ = new_n266_ & new_n1120_;
  assign new_n1122_ = ~new_n1119_ & ~new_n1121_;
  assign new_n1123_ = ~new_n1115_ & new_n1122_;
  assign new_n1124_ = A298 & ~A269;
  assign new_n1125_ = ~A267 & ~A236;
  assign new_n1126_ = new_n1124_ & new_n1125_;
  assign new_n1127_ = new_n1068_ & new_n1126_;
  assign new_n1128_ = new_n266_ & new_n1127_;
  assign new_n1129_ = A298 & A266;
  assign new_n1130_ = new_n268_ & new_n1129_;
  assign new_n1131_ = new_n1068_ & new_n1130_;
  assign new_n1132_ = new_n266_ & new_n1131_;
  assign new_n1133_ = ~A298 & ~A269;
  assign new_n1134_ = new_n1125_ & new_n1133_;
  assign new_n1135_ = new_n1062_ & new_n1134_;
  assign new_n1136_ = new_n266_ & new_n1135_;
  assign new_n1137_ = ~new_n1132_ & ~new_n1136_;
  assign new_n1138_ = ~new_n1128_ & new_n1137_;
  assign new_n1139_ = new_n1123_ & new_n1138_;
  assign new_n1140_ = new_n1111_ & new_n1139_;
  assign new_n1141_ = new_n262_ & new_n950_;
  assign new_n1142_ = new_n266_ & new_n1141_;
  assign new_n1143_ = ~A298 & A268;
  assign new_n1144_ = new_n1125_ & new_n1143_;
  assign new_n1145_ = new_n1062_ & new_n1144_;
  assign new_n1146_ = new_n266_ & new_n1145_;
  assign new_n1147_ = A298 & A268;
  assign new_n1148_ = new_n1125_ & new_n1147_;
  assign new_n1149_ = new_n1068_ & new_n1148_;
  assign new_n1150_ = new_n266_ & new_n1149_;
  assign new_n1151_ = ~new_n1146_ & ~new_n1150_;
  assign new_n1152_ = ~new_n1142_ & new_n1151_;
  assign new_n1153_ = new_n262_ & new_n963_;
  assign new_n1154_ = new_n266_ & new_n1153_;
  assign new_n1155_ = new_n262_ & new_n953_;
  assign new_n1156_ = new_n266_ & new_n1155_;
  assign new_n1157_ = new_n262_ & new_n947_;
  assign new_n1158_ = new_n266_ & new_n1157_;
  assign new_n1159_ = ~new_n1156_ & ~new_n1158_;
  assign new_n1160_ = ~new_n1154_ & new_n1159_;
  assign new_n1161_ = new_n1152_ & new_n1160_;
  assign new_n1162_ = new_n287_ & new_n1058_;
  assign new_n1163_ = new_n266_ & new_n1162_;
  assign new_n1164_ = new_n280_ & new_n1063_;
  assign new_n1165_ = new_n1062_ & new_n1164_;
  assign new_n1166_ = new_n266_ & new_n1165_;
  assign new_n1167_ = new_n280_ & new_n1069_;
  assign new_n1168_ = new_n1068_ & new_n1167_;
  assign new_n1169_ = new_n266_ & new_n1168_;
  assign new_n1170_ = ~new_n1166_ & ~new_n1169_;
  assign new_n1171_ = ~new_n1163_ & new_n1170_;
  assign new_n1172_ = new_n287_ & new_n1078_;
  assign new_n1173_ = new_n266_ & new_n1172_;
  assign new_n1174_ = new_n287_ & new_n1081_;
  assign new_n1175_ = new_n266_ & new_n1174_;
  assign new_n1176_ = ~new_n1173_ & ~new_n1175_;
  assign new_n1177_ = new_n1171_ & new_n1176_;
  assign new_n1178_ = new_n1161_ & new_n1177_;
  assign new_n1179_ = new_n1140_ & new_n1178_;
  assign new_n1180_ = new_n1088_ & new_n1179_;
  assign new_n1181_ = new_n286_ & new_n1093_;
  assign new_n1182_ = new_n1098_ & new_n1181_;
  assign new_n1183_ = new_n266_ & new_n1182_;
  assign new_n1184_ = new_n287_ & new_n1075_;
  assign new_n1185_ = new_n266_ & new_n1184_;
  assign new_n1186_ = new_n1092_ & new_n1181_;
  assign new_n1187_ = new_n266_ & new_n1186_;
  assign new_n1188_ = ~new_n1185_ & ~new_n1187_;
  assign new_n1189_ = ~new_n1183_ & new_n1188_;
  assign new_n1190_ = new_n281_ & new_n1081_;
  assign new_n1191_ = new_n266_ & new_n1190_;
  assign new_n1192_ = new_n281_ & new_n1058_;
  assign new_n1193_ = new_n266_ & new_n1192_;
  assign new_n1194_ = new_n281_ & new_n1078_;
  assign new_n1195_ = new_n266_ & new_n1194_;
  assign new_n1196_ = ~new_n1193_ & ~new_n1195_;
  assign new_n1197_ = ~new_n1191_ & new_n1196_;
  assign new_n1198_ = new_n1189_ & new_n1197_;
  assign new_n1199_ = new_n280_ & new_n1116_;
  assign new_n1200_ = new_n1098_ & new_n1199_;
  assign new_n1201_ = new_n266_ & new_n1200_;
  assign new_n1202_ = new_n281_ & new_n1075_;
  assign new_n1203_ = new_n266_ & new_n1202_;
  assign new_n1204_ = new_n1092_ & new_n1199_;
  assign new_n1205_ = new_n266_ & new_n1204_;
  assign new_n1206_ = ~new_n1203_ & ~new_n1205_;
  assign new_n1207_ = ~new_n1201_ & new_n1206_;
  assign new_n1208_ = ~A267 & A235;
  assign new_n1209_ = new_n1133_ & new_n1208_;
  assign new_n1210_ = new_n1062_ & new_n1209_;
  assign new_n1211_ = new_n266_ & new_n1210_;
  assign new_n1212_ = new_n286_ & new_n1112_;
  assign new_n1213_ = new_n1062_ & new_n1212_;
  assign new_n1214_ = new_n266_ & new_n1213_;
  assign new_n1215_ = new_n286_ & new_n1129_;
  assign new_n1216_ = new_n1068_ & new_n1215_;
  assign new_n1217_ = new_n266_ & new_n1216_;
  assign new_n1218_ = ~new_n1214_ & ~new_n1217_;
  assign new_n1219_ = ~new_n1211_ & new_n1218_;
  assign new_n1220_ = new_n1207_ & new_n1219_;
  assign new_n1221_ = new_n1198_ & new_n1220_;
  assign new_n1222_ = new_n1147_ & new_n1208_;
  assign new_n1223_ = new_n1068_ & new_n1222_;
  assign new_n1224_ = new_n266_ & new_n1223_;
  assign new_n1225_ = new_n1124_ & new_n1208_;
  assign new_n1226_ = new_n1068_ & new_n1225_;
  assign new_n1227_ = new_n266_ & new_n1226_;
  assign new_n1228_ = new_n1143_ & new_n1208_;
  assign new_n1229_ = new_n1062_ & new_n1228_;
  assign new_n1230_ = new_n266_ & new_n1229_;
  assign new_n1231_ = ~new_n1227_ & ~new_n1230_;
  assign new_n1232_ = ~new_n1224_ & new_n1231_;
  assign new_n1233_ = new_n297_ & new_n947_;
  assign new_n1234_ = new_n266_ & new_n1233_;
  assign new_n1235_ = new_n297_ & new_n950_;
  assign new_n1236_ = new_n266_ & new_n1235_;
  assign new_n1237_ = new_n297_ & new_n953_;
  assign new_n1238_ = new_n266_ & new_n1237_;
  assign new_n1239_ = ~new_n1236_ & ~new_n1238_;
  assign new_n1240_ = ~new_n1234_ & new_n1239_;
  assign new_n1241_ = new_n1232_ & new_n1240_;
  assign new_n1242_ = new_n294_ & new_n954_;
  assign new_n1243_ = new_n297_ & new_n963_;
  assign new_n1244_ = new_n266_ & new_n1243_;
  assign new_n1245_ = new_n294_ & new_n951_;
  assign new_n1246_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1247_ = ~new_n1242_ & new_n1246_;
  assign new_n1248_ = new_n294_ & new_n948_;
  assign new_n1249_ = new_n294_ & new_n964_;
  assign new_n1250_ = ~new_n1248_ & ~new_n1249_;
  assign new_n1251_ = new_n1247_ & new_n1250_;
  assign new_n1252_ = new_n1241_ & new_n1251_;
  assign new_n1253_ = new_n1221_ & new_n1252_;
  assign new_n1254_ = new_n294_ & new_n975_;
  assign new_n1255_ = new_n294_ & new_n967_;
  assign new_n1256_ = new_n294_ & new_n961_;
  assign new_n1257_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1258_ = ~new_n1254_ & new_n1257_;
  assign new_n1259_ = new_n294_ & new_n987_;
  assign new_n1260_ = new_n294_ & new_n978_;
  assign new_n1261_ = new_n294_ & new_n972_;
  assign new_n1262_ = ~new_n1260_ & ~new_n1261_;
  assign new_n1263_ = ~new_n1259_ & new_n1262_;
  assign new_n1264_ = new_n1258_ & new_n1263_;
  assign new_n1265_ = new_n294_ & new_n994_;
  assign new_n1266_ = new_n294_ & new_n990_;
  assign new_n1267_ = new_n294_ & new_n984_;
  assign new_n1268_ = ~new_n1266_ & ~new_n1267_;
  assign new_n1269_ = ~new_n1265_ & new_n1268_;
  assign new_n1270_ = new_n294_ & new_n1010_;
  assign new_n1271_ = new_n294_ & new_n996_;
  assign new_n1272_ = new_n294_ & new_n1008_;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = ~new_n1270_ & new_n1273_;
  assign new_n1275_ = new_n1269_ & new_n1274_;
  assign new_n1276_ = new_n1264_ & new_n1275_;
  assign new_n1277_ = new_n294_ & new_n1018_;
  assign new_n1278_ = new_n294_ & new_n1006_;
  assign new_n1279_ = new_n294_ & new_n1016_;
  assign new_n1280_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1281_ = ~new_n1277_ & new_n1280_;
  assign new_n1282_ = new_n294_ & new_n1027_;
  assign new_n1283_ = new_n294_ & new_n1014_;
  assign new_n1284_ = new_n294_ & new_n1025_;
  assign new_n1285_ = ~new_n1283_ & ~new_n1284_;
  assign new_n1286_ = ~new_n1282_ & new_n1285_;
  assign new_n1287_ = new_n1281_ & new_n1286_;
  assign new_n1288_ = new_n294_ & new_n1035_;
  assign new_n1289_ = new_n294_ & new_n1023_;
  assign new_n1290_ = new_n294_ & new_n1033_;
  assign new_n1291_ = ~new_n1289_ & ~new_n1290_;
  assign new_n1292_ = ~new_n1288_ & new_n1291_;
  assign new_n1293_ = new_n294_ & new_n1031_;
  assign new_n1294_ = new_n294_ & new_n1043_;
  assign new_n1295_ = ~new_n1293_ & ~new_n1294_;
  assign new_n1296_ = new_n1292_ & new_n1295_;
  assign new_n1297_ = new_n1287_ & new_n1296_;
  assign new_n1298_ = new_n1276_ & new_n1297_;
  assign new_n1299_ = new_n1253_ & new_n1298_;
  assign new_n1300_ = new_n1180_ & new_n1299_;
  assign new_n1301_ = new_n294_ & new_n1051_;
  assign new_n1302_ = new_n294_ & new_n1045_;
  assign new_n1303_ = new_n294_ & new_n1041_;
  assign new_n1304_ = ~new_n1302_ & ~new_n1303_;
  assign new_n1305_ = ~new_n1301_ & new_n1304_;
  assign new_n1306_ = new_n352_ & new_n1065_;
  assign new_n1307_ = new_n294_ & new_n1053_;
  assign new_n1308_ = new_n294_ & new_n1049_;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign new_n1310_ = ~new_n1306_ & new_n1309_;
  assign new_n1311_ = new_n1305_ & new_n1310_;
  assign new_n1312_ = new_n352_ & new_n1079_;
  assign new_n1313_ = new_n352_ & new_n1071_;
  assign new_n1314_ = new_n352_ & new_n1059_;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1316_ = ~new_n1312_ & new_n1315_;
  assign new_n1317_ = new_n352_ & new_n1095_;
  assign new_n1318_ = new_n352_ & new_n1082_;
  assign new_n1319_ = new_n352_ & new_n1076_;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = ~new_n1317_ & new_n1320_;
  assign new_n1322_ = new_n1316_ & new_n1321_;
  assign new_n1323_ = new_n1311_ & new_n1322_;
  assign new_n1324_ = new_n352_ & new_n1105_;
  assign new_n1325_ = new_n352_ & new_n1099_;
  assign new_n1326_ = new_n352_ & new_n1089_;
  assign new_n1327_ = ~new_n1325_ & ~new_n1326_;
  assign new_n1328_ = ~new_n1324_ & new_n1327_;
  assign new_n1329_ = new_n352_ & new_n1118_;
  assign new_n1330_ = new_n352_ & new_n1107_;
  assign new_n1331_ = new_n352_ & new_n1103_;
  assign new_n1332_ = ~new_n1330_ & ~new_n1331_;
  assign new_n1333_ = ~new_n1329_ & new_n1332_;
  assign new_n1334_ = new_n1328_ & new_n1333_;
  assign new_n1335_ = new_n352_ & new_n1131_;
  assign new_n1336_ = new_n352_ & new_n1120_;
  assign new_n1337_ = new_n352_ & new_n1114_;
  assign new_n1338_ = ~new_n1336_ & ~new_n1337_;
  assign new_n1339_ = ~new_n1335_ & new_n1338_;
  assign new_n1340_ = new_n352_ & new_n1135_;
  assign new_n1341_ = new_n352_ & new_n1127_;
  assign new_n1342_ = ~new_n1340_ & ~new_n1341_;
  assign new_n1343_ = new_n1339_ & new_n1342_;
  assign new_n1344_ = new_n1334_ & new_n1343_;
  assign new_n1345_ = new_n1323_ & new_n1344_;
  assign new_n1346_ = new_n352_ & new_n1141_;
  assign new_n1347_ = new_n352_ & new_n1145_;
  assign new_n1348_ = new_n352_ & new_n1149_;
  assign new_n1349_ = ~new_n1347_ & ~new_n1348_;
  assign new_n1350_ = ~new_n1346_ & new_n1349_;
  assign new_n1351_ = new_n352_ & new_n1153_;
  assign new_n1352_ = new_n352_ & new_n1155_;
  assign new_n1353_ = new_n352_ & new_n1157_;
  assign new_n1354_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1355_ = ~new_n1351_ & new_n1354_;
  assign new_n1356_ = new_n1350_ & new_n1355_;
  assign new_n1357_ = new_n352_ & new_n1162_;
  assign new_n1358_ = new_n352_ & new_n1165_;
  assign new_n1359_ = new_n352_ & new_n1168_;
  assign new_n1360_ = ~new_n1358_ & ~new_n1359_;
  assign new_n1361_ = ~new_n1357_ & new_n1360_;
  assign new_n1362_ = new_n352_ & new_n1184_;
  assign new_n1363_ = new_n352_ & new_n1172_;
  assign new_n1364_ = new_n352_ & new_n1174_;
  assign new_n1365_ = ~new_n1363_ & ~new_n1364_;
  assign new_n1366_ = ~new_n1362_ & new_n1365_;
  assign new_n1367_ = new_n1361_ & new_n1366_;
  assign new_n1368_ = new_n1356_ & new_n1367_;
  assign new_n1369_ = new_n352_ & new_n1192_;
  assign new_n1370_ = new_n352_ & new_n1186_;
  assign new_n1371_ = new_n352_ & new_n1182_;
  assign new_n1372_ = ~new_n1370_ & ~new_n1371_;
  assign new_n1373_ = ~new_n1369_ & new_n1372_;
  assign new_n1374_ = new_n352_ & new_n1202_;
  assign new_n1375_ = new_n352_ & new_n1194_;
  assign new_n1376_ = new_n352_ & new_n1190_;
  assign new_n1377_ = ~new_n1375_ & ~new_n1376_;
  assign new_n1378_ = ~new_n1374_ & new_n1377_;
  assign new_n1379_ = new_n1373_ & new_n1378_;
  assign new_n1380_ = new_n352_ & new_n1213_;
  assign new_n1381_ = new_n352_ & new_n1204_;
  assign new_n1382_ = new_n352_ & new_n1200_;
  assign new_n1383_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1384_ = ~new_n1380_ & new_n1383_;
  assign new_n1385_ = new_n352_ & new_n1216_;
  assign new_n1386_ = new_n352_ & new_n1210_;
  assign new_n1387_ = ~new_n1385_ & ~new_n1386_;
  assign new_n1388_ = new_n1384_ & new_n1387_;
  assign new_n1389_ = new_n1379_ & new_n1388_;
  assign new_n1390_ = new_n1368_ & new_n1389_;
  assign new_n1391_ = new_n1345_ & new_n1390_;
  assign new_n1392_ = new_n352_ & new_n1223_;
  assign new_n1393_ = new_n352_ & new_n1226_;
  assign new_n1394_ = new_n352_ & new_n1229_;
  assign new_n1395_ = ~new_n1393_ & ~new_n1394_;
  assign new_n1396_ = ~new_n1392_ & new_n1395_;
  assign new_n1397_ = new_n352_ & new_n1233_;
  assign new_n1398_ = new_n352_ & new_n1235_;
  assign new_n1399_ = new_n352_ & new_n1237_;
  assign new_n1400_ = ~new_n1398_ & ~new_n1399_;
  assign new_n1401_ = ~new_n1397_ & new_n1400_;
  assign new_n1402_ = new_n1396_ & new_n1401_;
  assign new_n1403_ = new_n372_ & new_n954_;
  assign new_n1404_ = new_n352_ & new_n1243_;
  assign new_n1405_ = new_n372_ & new_n951_;
  assign new_n1406_ = ~new_n1404_ & ~new_n1405_;
  assign new_n1407_ = ~new_n1403_ & new_n1406_;
  assign new_n1408_ = new_n372_ & new_n967_;
  assign new_n1409_ = new_n372_ & new_n948_;
  assign new_n1410_ = new_n372_ & new_n964_;
  assign new_n1411_ = ~new_n1409_ & ~new_n1410_;
  assign new_n1412_ = ~new_n1408_ & new_n1411_;
  assign new_n1413_ = new_n1407_ & new_n1412_;
  assign new_n1414_ = new_n1402_ & new_n1413_;
  assign new_n1415_ = new_n372_ & new_n978_;
  assign new_n1416_ = new_n372_ & new_n961_;
  assign new_n1417_ = new_n372_ & new_n975_;
  assign new_n1418_ = ~new_n1416_ & ~new_n1417_;
  assign new_n1419_ = ~new_n1415_ & new_n1418_;
  assign new_n1420_ = new_n372_ & new_n990_;
  assign new_n1421_ = new_n372_ & new_n972_;
  assign new_n1422_ = new_n372_ & new_n987_;
  assign new_n1423_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1424_ = ~new_n1420_ & new_n1423_;
  assign new_n1425_ = new_n1419_ & new_n1424_;
  assign new_n1426_ = new_n372_ & new_n996_;
  assign new_n1427_ = new_n372_ & new_n984_;
  assign new_n1428_ = new_n372_ & new_n994_;
  assign new_n1429_ = ~new_n1427_ & ~new_n1428_;
  assign new_n1430_ = ~new_n1426_ & new_n1429_;
  assign new_n1431_ = new_n372_ & new_n1008_;
  assign new_n1432_ = new_n372_ & new_n1010_;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = new_n1430_ & new_n1433_;
  assign new_n1435_ = new_n1425_ & new_n1434_;
  assign new_n1436_ = new_n1414_ & new_n1435_;
  assign new_n1437_ = new_n372_ & new_n1018_;
  assign new_n1438_ = new_n372_ & new_n1006_;
  assign new_n1439_ = new_n372_ & new_n1016_;
  assign new_n1440_ = ~new_n1438_ & ~new_n1439_;
  assign new_n1441_ = ~new_n1437_ & new_n1440_;
  assign new_n1442_ = new_n372_ & new_n1027_;
  assign new_n1443_ = new_n372_ & new_n1014_;
  assign new_n1444_ = new_n372_ & new_n1025_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = ~new_n1442_ & new_n1445_;
  assign new_n1447_ = new_n1441_ & new_n1446_;
  assign new_n1448_ = new_n372_ & new_n1035_;
  assign new_n1449_ = new_n372_ & new_n1023_;
  assign new_n1450_ = new_n372_ & new_n1033_;
  assign new_n1451_ = ~new_n1449_ & ~new_n1450_;
  assign new_n1452_ = ~new_n1448_ & new_n1451_;
  assign new_n1453_ = new_n372_ & new_n1045_;
  assign new_n1454_ = new_n372_ & new_n1031_;
  assign new_n1455_ = new_n372_ & new_n1043_;
  assign new_n1456_ = ~new_n1454_ & ~new_n1455_;
  assign new_n1457_ = ~new_n1453_ & new_n1456_;
  assign new_n1458_ = new_n1452_ & new_n1457_;
  assign new_n1459_ = new_n1447_ & new_n1458_;
  assign new_n1460_ = new_n372_ & new_n1053_;
  assign new_n1461_ = new_n372_ & new_n1041_;
  assign new_n1462_ = new_n372_ & new_n1051_;
  assign new_n1463_ = ~new_n1461_ & ~new_n1462_;
  assign new_n1464_ = ~new_n1460_ & new_n1463_;
  assign new_n1465_ = new_n419_ & new_n1071_;
  assign new_n1466_ = new_n372_ & new_n1049_;
  assign new_n1467_ = new_n419_ & new_n1065_;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign new_n1469_ = ~new_n1465_ & new_n1468_;
  assign new_n1470_ = new_n1464_ & new_n1469_;
  assign new_n1471_ = new_n419_ & new_n1082_;
  assign new_n1472_ = new_n419_ & new_n1059_;
  assign new_n1473_ = new_n419_ & new_n1079_;
  assign new_n1474_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1475_ = ~new_n1471_ & new_n1474_;
  assign new_n1476_ = new_n419_ & new_n1076_;
  assign new_n1477_ = new_n419_ & new_n1095_;
  assign new_n1478_ = ~new_n1476_ & ~new_n1477_;
  assign new_n1479_ = new_n1475_ & new_n1478_;
  assign new_n1480_ = new_n1470_ & new_n1479_;
  assign new_n1481_ = new_n1459_ & new_n1480_;
  assign new_n1482_ = new_n1436_ & new_n1481_;
  assign new_n1483_ = new_n1391_ & new_n1482_;
  assign new_n1484_ = new_n1300_ & new_n1483_;
  assign new_n1485_ = new_n419_ & new_n1105_;
  assign new_n1486_ = new_n419_ & new_n1099_;
  assign new_n1487_ = new_n419_ & new_n1089_;
  assign new_n1488_ = ~new_n1486_ & ~new_n1487_;
  assign new_n1489_ = ~new_n1485_ & new_n1488_;
  assign new_n1490_ = new_n419_ & new_n1118_;
  assign new_n1491_ = new_n419_ & new_n1107_;
  assign new_n1492_ = new_n419_ & new_n1103_;
  assign new_n1493_ = ~new_n1491_ & ~new_n1492_;
  assign new_n1494_ = ~new_n1490_ & new_n1493_;
  assign new_n1495_ = new_n1489_ & new_n1494_;
  assign new_n1496_ = new_n419_ & new_n1131_;
  assign new_n1497_ = new_n419_ & new_n1120_;
  assign new_n1498_ = new_n419_ & new_n1114_;
  assign new_n1499_ = ~new_n1497_ & ~new_n1498_;
  assign new_n1500_ = ~new_n1496_ & new_n1499_;
  assign new_n1501_ = new_n419_ & new_n1145_;
  assign new_n1502_ = new_n419_ & new_n1135_;
  assign new_n1503_ = new_n419_ & new_n1127_;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = ~new_n1501_ & new_n1504_;
  assign new_n1506_ = new_n1500_ & new_n1505_;
  assign new_n1507_ = new_n1495_ & new_n1506_;
  assign new_n1508_ = new_n419_ & new_n1155_;
  assign new_n1509_ = new_n419_ & new_n1149_;
  assign new_n1510_ = new_n419_ & new_n1141_;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = ~new_n1508_ & new_n1511_;
  assign new_n1513_ = new_n419_ & new_n1165_;
  assign new_n1514_ = new_n419_ & new_n1157_;
  assign new_n1515_ = new_n419_ & new_n1153_;
  assign new_n1516_ = ~new_n1514_ & ~new_n1515_;
  assign new_n1517_ = ~new_n1513_ & new_n1516_;
  assign new_n1518_ = new_n1512_ & new_n1517_;
  assign new_n1519_ = new_n419_ & new_n1172_;
  assign new_n1520_ = new_n419_ & new_n1168_;
  assign new_n1521_ = new_n419_ & new_n1162_;
  assign new_n1522_ = ~new_n1520_ & ~new_n1521_;
  assign new_n1523_ = ~new_n1519_ & new_n1522_;
  assign new_n1524_ = new_n419_ & new_n1174_;
  assign new_n1525_ = new_n419_ & new_n1184_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = new_n1523_ & new_n1526_;
  assign new_n1528_ = new_n1518_ & new_n1527_;
  assign new_n1529_ = new_n1507_ & new_n1528_;
  assign new_n1530_ = new_n419_ & new_n1192_;
  assign new_n1531_ = new_n419_ & new_n1186_;
  assign new_n1532_ = new_n419_ & new_n1182_;
  assign new_n1533_ = ~new_n1531_ & ~new_n1532_;
  assign new_n1534_ = ~new_n1530_ & new_n1533_;
  assign new_n1535_ = new_n419_ & new_n1202_;
  assign new_n1536_ = new_n419_ & new_n1194_;
  assign new_n1537_ = new_n419_ & new_n1190_;
  assign new_n1538_ = ~new_n1536_ & ~new_n1537_;
  assign new_n1539_ = ~new_n1535_ & new_n1538_;
  assign new_n1540_ = new_n1534_ & new_n1539_;
  assign new_n1541_ = new_n419_ & new_n1213_;
  assign new_n1542_ = new_n419_ & new_n1204_;
  assign new_n1543_ = new_n419_ & new_n1200_;
  assign new_n1544_ = ~new_n1542_ & ~new_n1543_;
  assign new_n1545_ = ~new_n1541_ & new_n1544_;
  assign new_n1546_ = new_n419_ & new_n1226_;
  assign new_n1547_ = new_n419_ & new_n1216_;
  assign new_n1548_ = new_n419_ & new_n1210_;
  assign new_n1549_ = ~new_n1547_ & ~new_n1548_;
  assign new_n1550_ = ~new_n1546_ & new_n1549_;
  assign new_n1551_ = new_n1545_ & new_n1550_;
  assign new_n1552_ = new_n1540_ & new_n1551_;
  assign new_n1553_ = new_n419_ & new_n1235_;
  assign new_n1554_ = new_n419_ & new_n1229_;
  assign new_n1555_ = new_n419_ & new_n1223_;
  assign new_n1556_ = ~new_n1554_ & ~new_n1555_;
  assign new_n1557_ = ~new_n1553_ & new_n1556_;
  assign new_n1558_ = new_n419_ & new_n1243_;
  assign new_n1559_ = new_n419_ & new_n1237_;
  assign new_n1560_ = new_n419_ & new_n1233_;
  assign new_n1561_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1562_ = ~new_n1558_ & new_n1561_;
  assign new_n1563_ = new_n1557_ & new_n1562_;
  assign new_n1564_ = new_n439_ & new_n948_;
  assign new_n1565_ = new_n439_ & new_n951_;
  assign new_n1566_ = new_n439_ & new_n954_;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = ~new_n1564_ & new_n1567_;
  assign new_n1569_ = new_n439_ & new_n964_;
  assign new_n1570_ = new_n439_ & new_n967_;
  assign new_n1571_ = ~new_n1569_ & ~new_n1570_;
  assign new_n1572_ = new_n1568_ & new_n1571_;
  assign new_n1573_ = new_n1563_ & new_n1572_;
  assign new_n1574_ = new_n1552_ & new_n1573_;
  assign new_n1575_ = new_n1529_ & new_n1574_;
  assign new_n1576_ = new_n439_ & new_n978_;
  assign new_n1577_ = new_n439_ & new_n961_;
  assign new_n1578_ = new_n439_ & new_n975_;
  assign new_n1579_ = ~new_n1577_ & ~new_n1578_;
  assign new_n1580_ = ~new_n1576_ & new_n1579_;
  assign new_n1581_ = new_n439_ & new_n990_;
  assign new_n1582_ = new_n439_ & new_n972_;
  assign new_n1583_ = new_n439_ & new_n987_;
  assign new_n1584_ = ~new_n1582_ & ~new_n1583_;
  assign new_n1585_ = ~new_n1581_ & new_n1584_;
  assign new_n1586_ = new_n1580_ & new_n1585_;
  assign new_n1587_ = new_n439_ & new_n996_;
  assign new_n1588_ = new_n439_ & new_n984_;
  assign new_n1589_ = new_n439_ & new_n994_;
  assign new_n1590_ = ~new_n1588_ & ~new_n1589_;
  assign new_n1591_ = ~new_n1587_ & new_n1590_;
  assign new_n1592_ = new_n439_ & new_n1006_;
  assign new_n1593_ = new_n439_ & new_n1008_;
  assign new_n1594_ = new_n439_ & new_n1010_;
  assign new_n1595_ = ~new_n1593_ & ~new_n1594_;
  assign new_n1596_ = ~new_n1592_ & new_n1595_;
  assign new_n1597_ = new_n1591_ & new_n1596_;
  assign new_n1598_ = new_n1586_ & new_n1597_;
  assign new_n1599_ = new_n439_ & new_n1014_;
  assign new_n1600_ = new_n439_ & new_n1016_;
  assign new_n1601_ = new_n439_ & new_n1018_;
  assign new_n1602_ = ~new_n1600_ & ~new_n1601_;
  assign new_n1603_ = ~new_n1599_ & new_n1602_;
  assign new_n1604_ = new_n439_ & new_n1023_;
  assign new_n1605_ = new_n439_ & new_n1025_;
  assign new_n1606_ = new_n439_ & new_n1027_;
  assign new_n1607_ = ~new_n1605_ & ~new_n1606_;
  assign new_n1608_ = ~new_n1604_ & new_n1607_;
  assign new_n1609_ = new_n1603_ & new_n1608_;
  assign new_n1610_ = new_n439_ & new_n1031_;
  assign new_n1611_ = new_n439_ & new_n1033_;
  assign new_n1612_ = new_n439_ & new_n1035_;
  assign new_n1613_ = ~new_n1611_ & ~new_n1612_;
  assign new_n1614_ = ~new_n1610_ & new_n1613_;
  assign new_n1615_ = new_n439_ & new_n1043_;
  assign new_n1616_ = new_n439_ & new_n1045_;
  assign new_n1617_ = ~new_n1615_ & ~new_n1616_;
  assign new_n1618_ = new_n1614_ & new_n1617_;
  assign new_n1619_ = new_n1609_ & new_n1618_;
  assign new_n1620_ = new_n1598_ & new_n1619_;
  assign new_n1621_ = new_n439_ & new_n1053_;
  assign new_n1622_ = new_n439_ & new_n1041_;
  assign new_n1623_ = new_n439_ & new_n1051_;
  assign new_n1624_ = ~new_n1622_ & ~new_n1623_;
  assign new_n1625_ = ~new_n1621_ & new_n1624_;
  assign new_n1626_ = new_n487_ & new_n1071_;
  assign new_n1627_ = new_n439_ & new_n1049_;
  assign new_n1628_ = new_n487_ & new_n1065_;
  assign new_n1629_ = ~new_n1627_ & ~new_n1628_;
  assign new_n1630_ = ~new_n1626_ & new_n1629_;
  assign new_n1631_ = new_n1625_ & new_n1630_;
  assign new_n1632_ = new_n487_ & new_n1082_;
  assign new_n1633_ = new_n487_ & new_n1059_;
  assign new_n1634_ = new_n487_ & new_n1079_;
  assign new_n1635_ = ~new_n1633_ & ~new_n1634_;
  assign new_n1636_ = ~new_n1632_ & new_n1635_;
  assign new_n1637_ = new_n487_ & new_n1099_;
  assign new_n1638_ = new_n487_ & new_n1076_;
  assign new_n1639_ = new_n487_ & new_n1095_;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1641_ = ~new_n1637_ & new_n1640_;
  assign new_n1642_ = new_n1636_ & new_n1641_;
  assign new_n1643_ = new_n1631_ & new_n1642_;
  assign new_n1644_ = new_n487_ & new_n1107_;
  assign new_n1645_ = new_n487_ & new_n1089_;
  assign new_n1646_ = new_n487_ & new_n1105_;
  assign new_n1647_ = ~new_n1645_ & ~new_n1646_;
  assign new_n1648_ = ~new_n1644_ & new_n1647_;
  assign new_n1649_ = new_n487_ & new_n1120_;
  assign new_n1650_ = new_n487_ & new_n1103_;
  assign new_n1651_ = new_n487_ & new_n1118_;
  assign new_n1652_ = ~new_n1650_ & ~new_n1651_;
  assign new_n1653_ = ~new_n1649_ & new_n1652_;
  assign new_n1654_ = new_n1648_ & new_n1653_;
  assign new_n1655_ = new_n487_ & new_n1135_;
  assign new_n1656_ = new_n487_ & new_n1114_;
  assign new_n1657_ = new_n487_ & new_n1131_;
  assign new_n1658_ = ~new_n1656_ & ~new_n1657_;
  assign new_n1659_ = ~new_n1655_ & new_n1658_;
  assign new_n1660_ = new_n487_ & new_n1127_;
  assign new_n1661_ = new_n487_ & new_n1145_;
  assign new_n1662_ = ~new_n1660_ & ~new_n1661_;
  assign new_n1663_ = new_n1659_ & new_n1662_;
  assign new_n1664_ = new_n1654_ & new_n1663_;
  assign new_n1665_ = new_n1643_ & new_n1664_;
  assign new_n1666_ = new_n1620_ & new_n1665_;
  assign new_n1667_ = new_n1575_ & new_n1666_;
  assign new_n1668_ = new_n487_ & new_n1155_;
  assign new_n1669_ = new_n487_ & new_n1149_;
  assign new_n1670_ = new_n487_ & new_n1141_;
  assign new_n1671_ = ~new_n1669_ & ~new_n1670_;
  assign new_n1672_ = ~new_n1668_ & new_n1671_;
  assign new_n1673_ = new_n487_ & new_n1165_;
  assign new_n1674_ = new_n487_ & new_n1157_;
  assign new_n1675_ = new_n487_ & new_n1153_;
  assign new_n1676_ = ~new_n1674_ & ~new_n1675_;
  assign new_n1677_ = ~new_n1673_ & new_n1676_;
  assign new_n1678_ = new_n1672_ & new_n1677_;
  assign new_n1679_ = new_n487_ & new_n1172_;
  assign new_n1680_ = new_n487_ & new_n1168_;
  assign new_n1681_ = new_n487_ & new_n1162_;
  assign new_n1682_ = ~new_n1680_ & ~new_n1681_;
  assign new_n1683_ = ~new_n1679_ & new_n1682_;
  assign new_n1684_ = new_n487_ & new_n1186_;
  assign new_n1685_ = new_n487_ & new_n1174_;
  assign new_n1686_ = new_n487_ & new_n1184_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = ~new_n1684_ & new_n1687_;
  assign new_n1689_ = new_n1683_ & new_n1688_;
  assign new_n1690_ = new_n1678_ & new_n1689_;
  assign new_n1691_ = new_n487_ & new_n1194_;
  assign new_n1692_ = new_n487_ & new_n1182_;
  assign new_n1693_ = new_n487_ & new_n1192_;
  assign new_n1694_ = ~new_n1692_ & ~new_n1693_;
  assign new_n1695_ = ~new_n1691_ & new_n1694_;
  assign new_n1696_ = new_n487_ & new_n1204_;
  assign new_n1697_ = new_n487_ & new_n1190_;
  assign new_n1698_ = new_n487_ & new_n1202_;
  assign new_n1699_ = ~new_n1697_ & ~new_n1698_;
  assign new_n1700_ = ~new_n1696_ & new_n1699_;
  assign new_n1701_ = new_n1695_ & new_n1700_;
  assign new_n1702_ = new_n487_ & new_n1216_;
  assign new_n1703_ = new_n487_ & new_n1200_;
  assign new_n1704_ = new_n487_ & new_n1213_;
  assign new_n1705_ = ~new_n1703_ & ~new_n1704_;
  assign new_n1706_ = ~new_n1702_ & new_n1705_;
  assign new_n1707_ = new_n487_ & new_n1210_;
  assign new_n1708_ = new_n487_ & new_n1226_;
  assign new_n1709_ = ~new_n1707_ & ~new_n1708_;
  assign new_n1710_ = new_n1706_ & new_n1709_;
  assign new_n1711_ = new_n1701_ & new_n1710_;
  assign new_n1712_ = new_n1690_ & new_n1711_;
  assign new_n1713_ = new_n487_ & new_n1235_;
  assign new_n1714_ = new_n487_ & new_n1229_;
  assign new_n1715_ = new_n487_ & new_n1223_;
  assign new_n1716_ = ~new_n1714_ & ~new_n1715_;
  assign new_n1717_ = ~new_n1713_ & new_n1716_;
  assign new_n1718_ = new_n487_ & new_n1243_;
  assign new_n1719_ = new_n487_ & new_n1237_;
  assign new_n1720_ = new_n487_ & new_n1233_;
  assign new_n1721_ = ~new_n1719_ & ~new_n1720_;
  assign new_n1722_ = ~new_n1718_ & new_n1721_;
  assign new_n1723_ = new_n1717_ & new_n1722_;
  assign new_n1724_ = new_n230_ & new_n232_;
  assign new_n1725_ = new_n1062_ & new_n1724_;
  assign new_n1726_ = A234 & ~A200;
  assign new_n1727_ = new_n140_ & new_n1726_;
  assign new_n1728_ = ~A199 & A168;
  assign new_n1729_ = new_n40_ & new_n1728_;
  assign new_n1730_ = new_n1727_ & new_n1729_;
  assign new_n1731_ = new_n1725_ & new_n1730_;
  assign new_n1732_ = A300 & A269;
  assign new_n1733_ = new_n27_ & new_n1732_;
  assign new_n1734_ = new_n153_ & new_n155_;
  assign new_n1735_ = new_n1733_ & new_n1734_;
  assign new_n1736_ = new_n1730_ & new_n1735_;
  assign new_n1737_ = new_n153_ & new_n186_;
  assign new_n1738_ = new_n1733_ & new_n1737_;
  assign new_n1739_ = new_n1730_ & new_n1738_;
  assign new_n1740_ = ~new_n1736_ & ~new_n1739_;
  assign new_n1741_ = ~new_n1731_ & new_n1740_;
  assign new_n1742_ = A234 & A200;
  assign new_n1743_ = new_n140_ & new_n1742_;
  assign new_n1744_ = A199 & A168;
  assign new_n1745_ = new_n40_ & new_n1744_;
  assign new_n1746_ = new_n1743_ & new_n1745_;
  assign new_n1747_ = new_n1738_ & new_n1746_;
  assign new_n1748_ = new_n232_ & new_n247_;
  assign new_n1749_ = new_n1068_ & new_n1748_;
  assign new_n1750_ = new_n1730_ & new_n1749_;
  assign new_n1751_ = new_n1735_ & new_n1746_;
  assign new_n1752_ = ~new_n1750_ & ~new_n1751_;
  assign new_n1753_ = ~new_n1747_ & new_n1752_;
  assign new_n1754_ = new_n1741_ & new_n1753_;
  assign new_n1755_ = new_n1723_ & new_n1754_;
  assign new_n1756_ = A234 & ~A203;
  assign new_n1757_ = new_n140_ & new_n1756_;
  assign new_n1758_ = ~A201 & A168;
  assign new_n1759_ = new_n40_ & new_n1758_;
  assign new_n1760_ = new_n1757_ & new_n1759_;
  assign new_n1761_ = new_n1735_ & new_n1760_;
  assign new_n1762_ = new_n1725_ & new_n1746_;
  assign new_n1763_ = new_n1746_ & new_n1749_;
  assign new_n1764_ = ~new_n1762_ & ~new_n1763_;
  assign new_n1765_ = ~new_n1761_ & new_n1764_;
  assign new_n1766_ = new_n1749_ & new_n1760_;
  assign new_n1767_ = new_n1738_ & new_n1760_;
  assign new_n1768_ = new_n1725_ & new_n1760_;
  assign new_n1769_ = ~new_n1767_ & ~new_n1768_;
  assign new_n1770_ = ~new_n1766_ & new_n1769_;
  assign new_n1771_ = new_n1765_ & new_n1770_;
  assign new_n1772_ = A234 & A202;
  assign new_n1773_ = new_n140_ & new_n1772_;
  assign new_n1774_ = new_n1759_ & new_n1773_;
  assign new_n1775_ = new_n1725_ & new_n1774_;
  assign new_n1776_ = new_n1735_ & new_n1774_;
  assign new_n1777_ = new_n1738_ & new_n1774_;
  assign new_n1778_ = ~new_n1776_ & ~new_n1777_;
  assign new_n1779_ = ~new_n1775_ & new_n1778_;
  assign new_n1780_ = new_n1749_ & new_n1774_;
  assign new_n1781_ = ~A233 & ~A232;
  assign new_n1782_ = new_n505_ & new_n1781_;
  assign new_n1783_ = new_n508_ & new_n1782_;
  assign new_n1784_ = new_n1735_ & new_n1783_;
  assign new_n1785_ = ~new_n1780_ & ~new_n1784_;
  assign new_n1786_ = new_n1779_ & new_n1785_;
  assign new_n1787_ = new_n1771_ & new_n1786_;
  assign new_n1788_ = new_n1755_ & new_n1787_;
  assign new_n1789_ = new_n1712_ & new_n1788_;
  assign new_n1790_ = new_n1749_ & new_n1783_;
  assign new_n1791_ = new_n1738_ & new_n1783_;
  assign new_n1792_ = new_n1725_ & new_n1783_;
  assign new_n1793_ = ~new_n1791_ & ~new_n1792_;
  assign new_n1794_ = ~new_n1790_ & new_n1793_;
  assign new_n1795_ = A233 & A232;
  assign new_n1796_ = new_n505_ & new_n1795_;
  assign new_n1797_ = new_n508_ & new_n1796_;
  assign new_n1798_ = new_n1725_ & new_n1797_;
  assign new_n1799_ = new_n1735_ & new_n1797_;
  assign new_n1800_ = new_n1738_ & new_n1797_;
  assign new_n1801_ = ~new_n1799_ & ~new_n1800_;
  assign new_n1802_ = ~new_n1798_ & new_n1801_;
  assign new_n1803_ = new_n1794_ & new_n1802_;
  assign new_n1804_ = ~A236 & ~A234;
  assign new_n1805_ = new_n505_ & new_n1804_;
  assign new_n1806_ = new_n508_ & new_n1805_;
  assign new_n1807_ = new_n1738_ & new_n1806_;
  assign new_n1808_ = new_n1749_ & new_n1797_;
  assign new_n1809_ = new_n1735_ & new_n1806_;
  assign new_n1810_ = ~new_n1808_ & ~new_n1809_;
  assign new_n1811_ = ~new_n1807_ & new_n1810_;
  assign new_n1812_ = A235 & ~A234;
  assign new_n1813_ = new_n505_ & new_n1812_;
  assign new_n1814_ = new_n508_ & new_n1813_;
  assign new_n1815_ = new_n1735_ & new_n1814_;
  assign new_n1816_ = new_n1725_ & new_n1806_;
  assign new_n1817_ = new_n1749_ & new_n1806_;
  assign new_n1818_ = ~new_n1816_ & ~new_n1817_;
  assign new_n1819_ = ~new_n1815_ & new_n1818_;
  assign new_n1820_ = new_n1811_ & new_n1819_;
  assign new_n1821_ = new_n1803_ & new_n1820_;
  assign new_n1822_ = new_n1749_ & new_n1814_;
  assign new_n1823_ = new_n1738_ & new_n1814_;
  assign new_n1824_ = new_n1725_ & new_n1814_;
  assign new_n1825_ = ~new_n1823_ & ~new_n1824_;
  assign new_n1826_ = ~new_n1822_ & new_n1825_;
  assign new_n1827_ = new_n48_ & new_n1058_;
  assign new_n1828_ = new_n509_ & new_n1827_;
  assign new_n1829_ = new_n52_ & new_n1063_;
  assign new_n1830_ = new_n1062_ & new_n1829_;
  assign new_n1831_ = new_n509_ & new_n1830_;
  assign new_n1832_ = new_n52_ & new_n1069_;
  assign new_n1833_ = new_n1068_ & new_n1832_;
  assign new_n1834_ = new_n509_ & new_n1833_;
  assign new_n1835_ = ~new_n1831_ & ~new_n1834_;
  assign new_n1836_ = ~new_n1828_ & new_n1835_;
  assign new_n1837_ = new_n1826_ & new_n1836_;
  assign new_n1838_ = new_n48_ & new_n1075_;
  assign new_n1839_ = new_n509_ & new_n1838_;
  assign new_n1840_ = new_n48_ & new_n1078_;
  assign new_n1841_ = new_n509_ & new_n1840_;
  assign new_n1842_ = new_n48_ & new_n1081_;
  assign new_n1843_ = new_n509_ & new_n1842_;
  assign new_n1844_ = ~new_n1841_ & ~new_n1843_;
  assign new_n1845_ = ~new_n1839_ & new_n1844_;
  assign new_n1846_ = new_n47_ & new_n1093_;
  assign new_n1847_ = new_n1092_ & new_n1846_;
  assign new_n1848_ = new_n509_ & new_n1847_;
  assign new_n1849_ = new_n1098_ & new_n1846_;
  assign new_n1850_ = new_n509_ & new_n1849_;
  assign new_n1851_ = ~new_n1848_ & ~new_n1850_;
  assign new_n1852_ = new_n1845_ & new_n1851_;
  assign new_n1853_ = new_n1837_ & new_n1852_;
  assign new_n1854_ = new_n1821_ & new_n1853_;
  assign new_n1855_ = new_n53_ & new_n1081_;
  assign new_n1856_ = new_n509_ & new_n1855_;
  assign new_n1857_ = new_n53_ & new_n1058_;
  assign new_n1858_ = new_n509_ & new_n1857_;
  assign new_n1859_ = new_n53_ & new_n1078_;
  assign new_n1860_ = new_n509_ & new_n1859_;
  assign new_n1861_ = ~new_n1858_ & ~new_n1860_;
  assign new_n1862_ = ~new_n1856_ & new_n1861_;
  assign new_n1863_ = new_n52_ & new_n1116_;
  assign new_n1864_ = new_n1098_ & new_n1863_;
  assign new_n1865_ = new_n509_ & new_n1864_;
  assign new_n1866_ = new_n53_ & new_n1075_;
  assign new_n1867_ = new_n509_ & new_n1866_;
  assign new_n1868_ = new_n1092_ & new_n1863_;
  assign new_n1869_ = new_n509_ & new_n1868_;
  assign new_n1870_ = ~new_n1867_ & ~new_n1869_;
  assign new_n1871_ = ~new_n1865_ & new_n1870_;
  assign new_n1872_ = new_n1862_ & new_n1871_;
  assign new_n1873_ = ~A267 & A236;
  assign new_n1874_ = new_n1133_ & new_n1873_;
  assign new_n1875_ = new_n1062_ & new_n1874_;
  assign new_n1876_ = new_n509_ & new_n1875_;
  assign new_n1877_ = new_n47_ & new_n1112_;
  assign new_n1878_ = new_n1062_ & new_n1877_;
  assign new_n1879_ = new_n509_ & new_n1878_;
  assign new_n1880_ = new_n47_ & new_n1129_;
  assign new_n1881_ = new_n1068_ & new_n1880_;
  assign new_n1882_ = new_n509_ & new_n1881_;
  assign new_n1883_ = ~new_n1879_ & ~new_n1882_;
  assign new_n1884_ = ~new_n1876_ & new_n1883_;
  assign new_n1885_ = new_n1147_ & new_n1873_;
  assign new_n1886_ = new_n1068_ & new_n1885_;
  assign new_n1887_ = new_n509_ & new_n1886_;
  assign new_n1888_ = new_n1124_ & new_n1873_;
  assign new_n1889_ = new_n1068_ & new_n1888_;
  assign new_n1890_ = new_n509_ & new_n1889_;
  assign new_n1891_ = new_n1143_ & new_n1873_;
  assign new_n1892_ = new_n1062_ & new_n1891_;
  assign new_n1893_ = new_n509_ & new_n1892_;
  assign new_n1894_ = ~new_n1890_ & ~new_n1893_;
  assign new_n1895_ = ~new_n1887_ & new_n1894_;
  assign new_n1896_ = new_n1884_ & new_n1895_;
  assign new_n1897_ = new_n1872_ & new_n1896_;
  assign new_n1898_ = new_n33_ & new_n947_;
  assign new_n1899_ = new_n509_ & new_n1898_;
  assign new_n1900_ = new_n33_ & new_n950_;
  assign new_n1901_ = new_n509_ & new_n1900_;
  assign new_n1902_ = new_n33_ & new_n953_;
  assign new_n1903_ = new_n509_ & new_n1902_;
  assign new_n1904_ = ~new_n1901_ & ~new_n1903_;
  assign new_n1905_ = ~new_n1899_ & new_n1904_;
  assign new_n1906_ = A234 & A203;
  assign new_n1907_ = new_n140_ & new_n1906_;
  assign new_n1908_ = ~A202 & A201;
  assign new_n1909_ = ~A168 & A169;
  assign new_n1910_ = new_n1908_ & new_n1909_;
  assign new_n1911_ = new_n1907_ & new_n1910_;
  assign new_n1912_ = new_n1738_ & new_n1911_;
  assign new_n1913_ = new_n33_ & new_n963_;
  assign new_n1914_ = new_n509_ & new_n1913_;
  assign new_n1915_ = new_n1735_ & new_n1911_;
  assign new_n1916_ = ~new_n1914_ & ~new_n1915_;
  assign new_n1917_ = ~new_n1912_ & new_n1916_;
  assign new_n1918_ = new_n1905_ & new_n1917_;
  assign new_n1919_ = new_n521_ & new_n1830_;
  assign new_n1920_ = new_n1725_ & new_n1911_;
  assign new_n1921_ = new_n1749_ & new_n1911_;
  assign new_n1922_ = ~new_n1920_ & ~new_n1921_;
  assign new_n1923_ = ~new_n1919_ & new_n1922_;
  assign new_n1924_ = new_n521_ & new_n1833_;
  assign new_n1925_ = new_n521_ & new_n1827_;
  assign new_n1926_ = ~new_n1924_ & ~new_n1925_;
  assign new_n1927_ = new_n1923_ & new_n1926_;
  assign new_n1928_ = new_n1918_ & new_n1927_;
  assign new_n1929_ = new_n1897_ & new_n1928_;
  assign new_n1930_ = new_n1854_ & new_n1929_;
  assign new_n1931_ = new_n1789_ & new_n1930_;
  assign new_n1932_ = new_n1667_ & new_n1931_;
  assign new_n1933_ = new_n1484_ & new_n1932_;
  assign new_n1934_ = new_n1005_ & new_n1933_;
  assign new_n1935_ = new_n521_ & new_n1838_;
  assign new_n1936_ = new_n521_ & new_n1840_;
  assign new_n1937_ = new_n521_ & new_n1842_;
  assign new_n1938_ = ~new_n1936_ & ~new_n1937_;
  assign new_n1939_ = ~new_n1935_ & new_n1938_;
  assign new_n1940_ = new_n521_ & new_n1857_;
  assign new_n1941_ = new_n521_ & new_n1847_;
  assign new_n1942_ = new_n521_ & new_n1849_;
  assign new_n1943_ = ~new_n1941_ & ~new_n1942_;
  assign new_n1944_ = ~new_n1940_ & new_n1943_;
  assign new_n1945_ = new_n1939_ & new_n1944_;
  assign new_n1946_ = new_n521_ & new_n1866_;
  assign new_n1947_ = new_n521_ & new_n1859_;
  assign new_n1948_ = new_n521_ & new_n1855_;
  assign new_n1949_ = ~new_n1947_ & ~new_n1948_;
  assign new_n1950_ = ~new_n1946_ & new_n1949_;
  assign new_n1951_ = new_n521_ & new_n1878_;
  assign new_n1952_ = new_n521_ & new_n1868_;
  assign new_n1953_ = new_n521_ & new_n1864_;
  assign new_n1954_ = ~new_n1952_ & ~new_n1953_;
  assign new_n1955_ = ~new_n1951_ & new_n1954_;
  assign new_n1956_ = new_n1950_ & new_n1955_;
  assign new_n1957_ = new_n1945_ & new_n1956_;
  assign new_n1958_ = new_n521_ & new_n1889_;
  assign new_n1959_ = new_n521_ & new_n1881_;
  assign new_n1960_ = new_n521_ & new_n1875_;
  assign new_n1961_ = ~new_n1959_ & ~new_n1960_;
  assign new_n1962_ = ~new_n1958_ & new_n1961_;
  assign new_n1963_ = new_n521_ & new_n1900_;
  assign new_n1964_ = new_n521_ & new_n1892_;
  assign new_n1965_ = new_n521_ & new_n1886_;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_;
  assign new_n1967_ = ~new_n1963_ & new_n1966_;
  assign new_n1968_ = new_n1962_ & new_n1967_;
  assign new_n1969_ = new_n521_ & new_n1913_;
  assign new_n1970_ = new_n521_ & new_n1902_;
  assign new_n1971_ = new_n521_ & new_n1898_;
  assign new_n1972_ = ~new_n1970_ & ~new_n1971_;
  assign new_n1973_ = ~new_n1969_ & new_n1972_;
  assign new_n1974_ = ~A236 & A234;
  assign new_n1975_ = new_n516_ & new_n1974_;
  assign new_n1976_ = new_n520_ & new_n1975_;
  assign new_n1977_ = new_n1725_ & new_n1976_;
  assign new_n1978_ = new_n1735_ & new_n1976_;
  assign new_n1979_ = new_n1738_ & new_n1976_;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = ~new_n1977_ & new_n1980_;
  assign new_n1982_ = new_n1973_ & new_n1981_;
  assign new_n1983_ = new_n1968_ & new_n1982_;
  assign new_n1984_ = new_n1957_ & new_n1983_;
  assign new_n1985_ = A235 & A234;
  assign new_n1986_ = new_n516_ & new_n1985_;
  assign new_n1987_ = new_n520_ & new_n1986_;
  assign new_n1988_ = new_n1738_ & new_n1987_;
  assign new_n1989_ = new_n1749_ & new_n1976_;
  assign new_n1990_ = new_n1735_ & new_n1987_;
  assign new_n1991_ = ~new_n1989_ & ~new_n1990_;
  assign new_n1992_ = ~new_n1988_ & new_n1991_;
  assign new_n1993_ = new_n535_ & new_n1830_;
  assign new_n1994_ = new_n1725_ & new_n1987_;
  assign new_n1995_ = new_n1749_ & new_n1987_;
  assign new_n1996_ = ~new_n1994_ & ~new_n1995_;
  assign new_n1997_ = ~new_n1993_ & new_n1996_;
  assign new_n1998_ = new_n1992_ & new_n1997_;
  assign new_n1999_ = new_n535_ & new_n1840_;
  assign new_n2000_ = new_n535_ & new_n1833_;
  assign new_n2001_ = new_n535_ & new_n1827_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = ~new_n1999_ & new_n2002_;
  assign new_n2004_ = new_n535_ & new_n1847_;
  assign new_n2005_ = new_n535_ & new_n1842_;
  assign new_n2006_ = new_n535_ & new_n1838_;
  assign new_n2007_ = ~new_n2005_ & ~new_n2006_;
  assign new_n2008_ = ~new_n2004_ & new_n2007_;
  assign new_n2009_ = new_n2003_ & new_n2008_;
  assign new_n2010_ = new_n1998_ & new_n2009_;
  assign new_n2011_ = new_n535_ & new_n1859_;
  assign new_n2012_ = new_n535_ & new_n1849_;
  assign new_n2013_ = new_n535_ & new_n1857_;
  assign new_n2014_ = ~new_n2012_ & ~new_n2013_;
  assign new_n2015_ = ~new_n2011_ & new_n2014_;
  assign new_n2016_ = new_n535_ & new_n1868_;
  assign new_n2017_ = new_n535_ & new_n1855_;
  assign new_n2018_ = new_n535_ & new_n1866_;
  assign new_n2019_ = ~new_n2017_ & ~new_n2018_;
  assign new_n2020_ = ~new_n2016_ & new_n2019_;
  assign new_n2021_ = new_n2015_ & new_n2020_;
  assign new_n2022_ = new_n535_ & new_n1881_;
  assign new_n2023_ = new_n535_ & new_n1864_;
  assign new_n2024_ = new_n535_ & new_n1878_;
  assign new_n2025_ = ~new_n2023_ & ~new_n2024_;
  assign new_n2026_ = ~new_n2022_ & new_n2025_;
  assign new_n2027_ = new_n535_ & new_n1875_;
  assign new_n2028_ = new_n535_ & new_n1889_;
  assign new_n2029_ = ~new_n2027_ & ~new_n2028_;
  assign new_n2030_ = new_n2026_ & new_n2029_;
  assign new_n2031_ = new_n2021_ & new_n2030_;
  assign new_n2032_ = new_n2010_ & new_n2031_;
  assign new_n2033_ = new_n1984_ & new_n2032_;
  assign new_n2034_ = new_n535_ & new_n1900_;
  assign new_n2035_ = new_n535_ & new_n1892_;
  assign new_n2036_ = new_n535_ & new_n1886_;
  assign new_n2037_ = ~new_n2035_ & ~new_n2036_;
  assign new_n2038_ = ~new_n2034_ & new_n2037_;
  assign new_n2039_ = new_n535_ & new_n1913_;
  assign new_n2040_ = new_n535_ & new_n1902_;
  assign new_n2041_ = new_n535_ & new_n1898_;
  assign new_n2042_ = ~new_n2040_ & ~new_n2041_;
  assign new_n2043_ = ~new_n2039_ & new_n2042_;
  assign new_n2044_ = new_n2038_ & new_n2043_;
  assign new_n2045_ = new_n533_ & new_n1974_;
  assign new_n2046_ = new_n520_ & new_n2045_;
  assign new_n2047_ = new_n1725_ & new_n2046_;
  assign new_n2048_ = new_n1735_ & new_n2046_;
  assign new_n2049_ = new_n1738_ & new_n2046_;
  assign new_n2050_ = ~new_n2048_ & ~new_n2049_;
  assign new_n2051_ = ~new_n2047_ & new_n2050_;
  assign new_n2052_ = new_n533_ & new_n1985_;
  assign new_n2053_ = new_n520_ & new_n2052_;
  assign new_n2054_ = new_n1738_ & new_n2053_;
  assign new_n2055_ = new_n1749_ & new_n2046_;
  assign new_n2056_ = new_n1735_ & new_n2053_;
  assign new_n2057_ = ~new_n2055_ & ~new_n2056_;
  assign new_n2058_ = ~new_n2054_ & new_n2057_;
  assign new_n2059_ = new_n2051_ & new_n2058_;
  assign new_n2060_ = new_n2044_ & new_n2059_;
  assign new_n2061_ = new_n543_ & new_n1830_;
  assign new_n2062_ = new_n1725_ & new_n2053_;
  assign new_n2063_ = new_n1749_ & new_n2053_;
  assign new_n2064_ = ~new_n2062_ & ~new_n2063_;
  assign new_n2065_ = ~new_n2061_ & new_n2064_;
  assign new_n2066_ = new_n543_ & new_n1840_;
  assign new_n2067_ = new_n543_ & new_n1833_;
  assign new_n2068_ = new_n543_ & new_n1827_;
  assign new_n2069_ = ~new_n2067_ & ~new_n2068_;
  assign new_n2070_ = ~new_n2066_ & new_n2069_;
  assign new_n2071_ = new_n2065_ & new_n2070_;
  assign new_n2072_ = new_n543_ & new_n1847_;
  assign new_n2073_ = new_n543_ & new_n1842_;
  assign new_n2074_ = new_n543_ & new_n1838_;
  assign new_n2075_ = ~new_n2073_ & ~new_n2074_;
  assign new_n2076_ = ~new_n2072_ & new_n2075_;
  assign new_n2077_ = new_n543_ & new_n1849_;
  assign new_n2078_ = new_n543_ & new_n1857_;
  assign new_n2079_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2080_ = new_n2076_ & new_n2079_;
  assign new_n2081_ = new_n2071_ & new_n2080_;
  assign new_n2082_ = new_n2060_ & new_n2081_;
  assign new_n2083_ = new_n543_ & new_n1866_;
  assign new_n2084_ = new_n543_ & new_n1859_;
  assign new_n2085_ = new_n543_ & new_n1855_;
  assign new_n2086_ = ~new_n2084_ & ~new_n2085_;
  assign new_n2087_ = ~new_n2083_ & new_n2086_;
  assign new_n2088_ = new_n543_ & new_n1878_;
  assign new_n2089_ = new_n543_ & new_n1868_;
  assign new_n2090_ = new_n543_ & new_n1864_;
  assign new_n2091_ = ~new_n2089_ & ~new_n2090_;
  assign new_n2092_ = ~new_n2088_ & new_n2091_;
  assign new_n2093_ = new_n2087_ & new_n2092_;
  assign new_n2094_ = new_n543_ & new_n1889_;
  assign new_n2095_ = new_n543_ & new_n1881_;
  assign new_n2096_ = new_n543_ & new_n1875_;
  assign new_n2097_ = ~new_n2095_ & ~new_n2096_;
  assign new_n2098_ = ~new_n2094_ & new_n2097_;
  assign new_n2099_ = new_n543_ & new_n1900_;
  assign new_n2100_ = new_n543_ & new_n1892_;
  assign new_n2101_ = new_n543_ & new_n1886_;
  assign new_n2102_ = ~new_n2100_ & ~new_n2101_;
  assign new_n2103_ = ~new_n2099_ & new_n2102_;
  assign new_n2104_ = new_n2098_ & new_n2103_;
  assign new_n2105_ = new_n2093_ & new_n2104_;
  assign new_n2106_ = new_n543_ & new_n1913_;
  assign new_n2107_ = new_n543_ & new_n1902_;
  assign new_n2108_ = new_n543_ & new_n1898_;
  assign new_n2109_ = ~new_n2107_ & ~new_n2108_;
  assign new_n2110_ = ~new_n2106_ & new_n2109_;
  assign new_n2111_ = new_n542_ & new_n1975_;
  assign new_n2112_ = new_n1725_ & new_n2111_;
  assign new_n2113_ = new_n1735_ & new_n2111_;
  assign new_n2114_ = new_n1738_ & new_n2111_;
  assign new_n2115_ = ~new_n2113_ & ~new_n2114_;
  assign new_n2116_ = ~new_n2112_ & new_n2115_;
  assign new_n2117_ = new_n2110_ & new_n2116_;
  assign new_n2118_ = new_n542_ & new_n1986_;
  assign new_n2119_ = new_n1738_ & new_n2118_;
  assign new_n2120_ = new_n1749_ & new_n2111_;
  assign new_n2121_ = new_n1735_ & new_n2118_;
  assign new_n2122_ = ~new_n2120_ & ~new_n2121_;
  assign new_n2123_ = ~new_n2119_ & new_n2122_;
  assign new_n2124_ = new_n1725_ & new_n2118_;
  assign new_n2125_ = new_n1749_ & new_n2118_;
  assign new_n2126_ = ~new_n2124_ & ~new_n2125_;
  assign new_n2127_ = new_n2123_ & new_n2126_;
  assign new_n2128_ = new_n2117_ & new_n2127_;
  assign new_n2129_ = new_n2105_ & new_n2128_;
  assign new_n2130_ = new_n2082_ & new_n2129_;
  assign new_n2131_ = new_n2033_ & new_n2130_;
  assign new_n2132_ = new_n551_ & new_n1827_;
  assign new_n2133_ = new_n551_ & new_n1830_;
  assign new_n2134_ = new_n551_ & new_n1833_;
  assign new_n2135_ = ~new_n2133_ & ~new_n2134_;
  assign new_n2136_ = ~new_n2132_ & new_n2135_;
  assign new_n2137_ = new_n551_ & new_n1838_;
  assign new_n2138_ = new_n551_ & new_n1840_;
  assign new_n2139_ = new_n551_ & new_n1842_;
  assign new_n2140_ = ~new_n2138_ & ~new_n2139_;
  assign new_n2141_ = ~new_n2137_ & new_n2140_;
  assign new_n2142_ = new_n2136_ & new_n2141_;
  assign new_n2143_ = new_n551_ & new_n1857_;
  assign new_n2144_ = new_n551_ & new_n1847_;
  assign new_n2145_ = new_n551_ & new_n1849_;
  assign new_n2146_ = ~new_n2144_ & ~new_n2145_;
  assign new_n2147_ = ~new_n2143_ & new_n2146_;
  assign new_n2148_ = new_n551_ & new_n1866_;
  assign new_n2149_ = new_n551_ & new_n1859_;
  assign new_n2150_ = new_n551_ & new_n1855_;
  assign new_n2151_ = ~new_n2149_ & ~new_n2150_;
  assign new_n2152_ = ~new_n2148_ & new_n2151_;
  assign new_n2153_ = new_n2147_ & new_n2152_;
  assign new_n2154_ = new_n2142_ & new_n2153_;
  assign new_n2155_ = new_n551_ & new_n1878_;
  assign new_n2156_ = new_n551_ & new_n1868_;
  assign new_n2157_ = new_n551_ & new_n1864_;
  assign new_n2158_ = ~new_n2156_ & ~new_n2157_;
  assign new_n2159_ = ~new_n2155_ & new_n2158_;
  assign new_n2160_ = new_n551_ & new_n1889_;
  assign new_n2161_ = new_n551_ & new_n1881_;
  assign new_n2162_ = new_n551_ & new_n1875_;
  assign new_n2163_ = ~new_n2161_ & ~new_n2162_;
  assign new_n2164_ = ~new_n2160_ & new_n2163_;
  assign new_n2165_ = new_n2159_ & new_n2164_;
  assign new_n2166_ = new_n551_ & new_n1900_;
  assign new_n2167_ = new_n551_ & new_n1892_;
  assign new_n2168_ = new_n551_ & new_n1886_;
  assign new_n2169_ = ~new_n2167_ & ~new_n2168_;
  assign new_n2170_ = ~new_n2166_ & new_n2169_;
  assign new_n2171_ = new_n551_ & new_n1902_;
  assign new_n2172_ = new_n551_ & new_n1898_;
  assign new_n2173_ = ~new_n2171_ & ~new_n2172_;
  assign new_n2174_ = new_n2170_ & new_n2173_;
  assign new_n2175_ = new_n2165_ & new_n2174_;
  assign new_n2176_ = new_n2154_ & new_n2175_;
  assign new_n2177_ = new_n542_ & new_n2045_;
  assign new_n2178_ = new_n1738_ & new_n2177_;
  assign new_n2179_ = new_n551_ & new_n1913_;
  assign new_n2180_ = new_n1735_ & new_n2177_;
  assign new_n2181_ = ~new_n2179_ & ~new_n2180_;
  assign new_n2182_ = ~new_n2178_ & new_n2181_;
  assign new_n2183_ = new_n542_ & new_n2052_;
  assign new_n2184_ = new_n1735_ & new_n2183_;
  assign new_n2185_ = new_n1725_ & new_n2177_;
  assign new_n2186_ = new_n1749_ & new_n2177_;
  assign new_n2187_ = ~new_n2185_ & ~new_n2186_;
  assign new_n2188_ = ~new_n2184_ & new_n2187_;
  assign new_n2189_ = new_n2182_ & new_n2188_;
  assign new_n2190_ = new_n1749_ & new_n2183_;
  assign new_n2191_ = new_n1738_ & new_n2183_;
  assign new_n2192_ = new_n1725_ & new_n2183_;
  assign new_n2193_ = ~new_n2191_ & ~new_n2192_;
  assign new_n2194_ = ~new_n2190_ & new_n2193_;
  assign new_n2195_ = ~A168 & A170;
  assign new_n2196_ = new_n1908_ & new_n2195_;
  assign new_n2197_ = new_n1907_ & new_n2196_;
  assign new_n2198_ = new_n1725_ & new_n2197_;
  assign new_n2199_ = new_n1735_ & new_n2197_;
  assign new_n2200_ = new_n1738_ & new_n2197_;
  assign new_n2201_ = ~new_n2199_ & ~new_n2200_;
  assign new_n2202_ = ~new_n2198_ & new_n2201_;
  assign new_n2203_ = new_n2194_ & new_n2202_;
  assign new_n2204_ = new_n2189_ & new_n2203_;
  assign new_n2205_ = new_n565_ & new_n1833_;
  assign new_n2206_ = new_n1749_ & new_n2197_;
  assign new_n2207_ = new_n565_ & new_n1830_;
  assign new_n2208_ = ~new_n2206_ & ~new_n2207_;
  assign new_n2209_ = ~new_n2205_ & new_n2208_;
  assign new_n2210_ = new_n565_ & new_n1842_;
  assign new_n2211_ = new_n565_ & new_n1827_;
  assign new_n2212_ = new_n565_ & new_n1840_;
  assign new_n2213_ = ~new_n2211_ & ~new_n2212_;
  assign new_n2214_ = ~new_n2210_ & new_n2213_;
  assign new_n2215_ = new_n2209_ & new_n2214_;
  assign new_n2216_ = new_n565_ & new_n1849_;
  assign new_n2217_ = new_n565_ & new_n1838_;
  assign new_n2218_ = new_n565_ & new_n1847_;
  assign new_n2219_ = ~new_n2217_ & ~new_n2218_;
  assign new_n2220_ = ~new_n2216_ & new_n2219_;
  assign new_n2221_ = new_n565_ & new_n1857_;
  assign new_n2222_ = new_n565_ & new_n1859_;
  assign new_n2223_ = ~new_n2221_ & ~new_n2222_;
  assign new_n2224_ = new_n2220_ & new_n2223_;
  assign new_n2225_ = new_n2215_ & new_n2224_;
  assign new_n2226_ = new_n2204_ & new_n2225_;
  assign new_n2227_ = new_n2176_ & new_n2226_;
  assign new_n2228_ = new_n565_ & new_n1868_;
  assign new_n2229_ = new_n565_ & new_n1855_;
  assign new_n2230_ = new_n565_ & new_n1866_;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = ~new_n2228_ & new_n2231_;
  assign new_n2233_ = new_n565_ & new_n1881_;
  assign new_n2234_ = new_n565_ & new_n1864_;
  assign new_n2235_ = new_n565_ & new_n1878_;
  assign new_n2236_ = ~new_n2234_ & ~new_n2235_;
  assign new_n2237_ = ~new_n2233_ & new_n2236_;
  assign new_n2238_ = new_n2232_ & new_n2237_;
  assign new_n2239_ = new_n565_ & new_n1892_;
  assign new_n2240_ = new_n565_ & new_n1875_;
  assign new_n2241_ = new_n565_ & new_n1889_;
  assign new_n2242_ = ~new_n2240_ & ~new_n2241_;
  assign new_n2243_ = ~new_n2239_ & new_n2242_;
  assign new_n2244_ = new_n565_ & new_n1902_;
  assign new_n2245_ = new_n565_ & new_n1886_;
  assign new_n2246_ = new_n565_ & new_n1900_;
  assign new_n2247_ = ~new_n2245_ & ~new_n2246_;
  assign new_n2248_ = ~new_n2244_ & new_n2247_;
  assign new_n2249_ = new_n2243_ & new_n2248_;
  assign new_n2250_ = new_n2238_ & new_n2249_;
  assign new_n2251_ = new_n564_ & new_n1975_;
  assign new_n2252_ = new_n1735_ & new_n2251_;
  assign new_n2253_ = new_n565_ & new_n1898_;
  assign new_n2254_ = new_n565_ & new_n1913_;
  assign new_n2255_ = ~new_n2253_ & ~new_n2254_;
  assign new_n2256_ = ~new_n2252_ & new_n2255_;
  assign new_n2257_ = new_n1749_ & new_n2251_;
  assign new_n2258_ = new_n1738_ & new_n2251_;
  assign new_n2259_ = new_n1725_ & new_n2251_;
  assign new_n2260_ = ~new_n2258_ & ~new_n2259_;
  assign new_n2261_ = ~new_n2257_ & new_n2260_;
  assign new_n2262_ = new_n2256_ & new_n2261_;
  assign new_n2263_ = new_n564_ & new_n1986_;
  assign new_n2264_ = new_n1725_ & new_n2263_;
  assign new_n2265_ = new_n1735_ & new_n2263_;
  assign new_n2266_ = new_n1738_ & new_n2263_;
  assign new_n2267_ = ~new_n2265_ & ~new_n2266_;
  assign new_n2268_ = ~new_n2264_ & new_n2267_;
  assign new_n2269_ = new_n1749_ & new_n2263_;
  assign new_n2270_ = new_n572_ & new_n1830_;
  assign new_n2271_ = ~new_n2269_ & ~new_n2270_;
  assign new_n2272_ = new_n2268_ & new_n2271_;
  assign new_n2273_ = new_n2262_ & new_n2272_;
  assign new_n2274_ = new_n2250_ & new_n2273_;
  assign new_n2275_ = new_n572_ & new_n1840_;
  assign new_n2276_ = new_n572_ & new_n1833_;
  assign new_n2277_ = new_n572_ & new_n1827_;
  assign new_n2278_ = ~new_n2276_ & ~new_n2277_;
  assign new_n2279_ = ~new_n2275_ & new_n2278_;
  assign new_n2280_ = new_n572_ & new_n1847_;
  assign new_n2281_ = new_n572_ & new_n1842_;
  assign new_n2282_ = new_n572_ & new_n1838_;
  assign new_n2283_ = ~new_n2281_ & ~new_n2282_;
  assign new_n2284_ = ~new_n2280_ & new_n2283_;
  assign new_n2285_ = new_n2279_ & new_n2284_;
  assign new_n2286_ = new_n572_ & new_n1859_;
  assign new_n2287_ = new_n572_ & new_n1849_;
  assign new_n2288_ = new_n572_ & new_n1857_;
  assign new_n2289_ = ~new_n2287_ & ~new_n2288_;
  assign new_n2290_ = ~new_n2286_ & new_n2289_;
  assign new_n2291_ = new_n572_ & new_n1868_;
  assign new_n2292_ = new_n572_ & new_n1855_;
  assign new_n2293_ = new_n572_ & new_n1866_;
  assign new_n2294_ = ~new_n2292_ & ~new_n2293_;
  assign new_n2295_ = ~new_n2291_ & new_n2294_;
  assign new_n2296_ = new_n2290_ & new_n2295_;
  assign new_n2297_ = new_n2285_ & new_n2296_;
  assign new_n2298_ = new_n572_ & new_n1881_;
  assign new_n2299_ = new_n572_ & new_n1864_;
  assign new_n2300_ = new_n572_ & new_n1878_;
  assign new_n2301_ = ~new_n2299_ & ~new_n2300_;
  assign new_n2302_ = ~new_n2298_ & new_n2301_;
  assign new_n2303_ = new_n572_ & new_n1892_;
  assign new_n2304_ = new_n572_ & new_n1875_;
  assign new_n2305_ = new_n572_ & new_n1889_;
  assign new_n2306_ = ~new_n2304_ & ~new_n2305_;
  assign new_n2307_ = ~new_n2303_ & new_n2306_;
  assign new_n2308_ = new_n2302_ & new_n2307_;
  assign new_n2309_ = new_n572_ & new_n1902_;
  assign new_n2310_ = new_n572_ & new_n1886_;
  assign new_n2311_ = new_n572_ & new_n1900_;
  assign new_n2312_ = ~new_n2310_ & ~new_n2311_;
  assign new_n2313_ = ~new_n2309_ & new_n2312_;
  assign new_n2314_ = new_n572_ & new_n1898_;
  assign new_n2315_ = new_n572_ & new_n1913_;
  assign new_n2316_ = ~new_n2314_ & ~new_n2315_;
  assign new_n2317_ = new_n2313_ & new_n2316_;
  assign new_n2318_ = new_n2308_ & new_n2317_;
  assign new_n2319_ = new_n2297_ & new_n2318_;
  assign new_n2320_ = new_n2274_ & new_n2319_;
  assign new_n2321_ = new_n2227_ & new_n2320_;
  assign new_n2322_ = new_n2131_ & new_n2321_;
  assign new_n2323_ = new_n564_ & new_n2045_;
  assign new_n2324_ = new_n1725_ & new_n2323_;
  assign new_n2325_ = new_n1735_ & new_n2323_;
  assign new_n2326_ = new_n1738_ & new_n2323_;
  assign new_n2327_ = ~new_n2325_ & ~new_n2326_;
  assign new_n2328_ = ~new_n2324_ & new_n2327_;
  assign new_n2329_ = new_n564_ & new_n2052_;
  assign new_n2330_ = new_n1738_ & new_n2329_;
  assign new_n2331_ = new_n1749_ & new_n2323_;
  assign new_n2332_ = new_n1735_ & new_n2329_;
  assign new_n2333_ = ~new_n2331_ & ~new_n2332_;
  assign new_n2334_ = ~new_n2330_ & new_n2333_;
  assign new_n2335_ = new_n2328_ & new_n2334_;
  assign new_n2336_ = new_n587_ & new_n1830_;
  assign new_n2337_ = new_n1725_ & new_n2329_;
  assign new_n2338_ = new_n1749_ & new_n2329_;
  assign new_n2339_ = ~new_n2337_ & ~new_n2338_;
  assign new_n2340_ = ~new_n2336_ & new_n2339_;
  assign new_n2341_ = new_n587_ & new_n1840_;
  assign new_n2342_ = new_n587_ & new_n1833_;
  assign new_n2343_ = new_n587_ & new_n1827_;
  assign new_n2344_ = ~new_n2342_ & ~new_n2343_;
  assign new_n2345_ = ~new_n2341_ & new_n2344_;
  assign new_n2346_ = new_n2340_ & new_n2345_;
  assign new_n2347_ = new_n2335_ & new_n2346_;
  assign new_n2348_ = new_n587_ & new_n1847_;
  assign new_n2349_ = new_n587_ & new_n1842_;
  assign new_n2350_ = new_n587_ & new_n1838_;
  assign new_n2351_ = ~new_n2349_ & ~new_n2350_;
  assign new_n2352_ = ~new_n2348_ & new_n2351_;
  assign new_n2353_ = new_n587_ & new_n1859_;
  assign new_n2354_ = new_n587_ & new_n1849_;
  assign new_n2355_ = new_n587_ & new_n1857_;
  assign new_n2356_ = ~new_n2354_ & ~new_n2355_;
  assign new_n2357_ = ~new_n2353_ & new_n2356_;
  assign new_n2358_ = new_n2352_ & new_n2357_;
  assign new_n2359_ = new_n587_ & new_n1868_;
  assign new_n2360_ = new_n587_ & new_n1855_;
  assign new_n2361_ = new_n587_ & new_n1866_;
  assign new_n2362_ = ~new_n2360_ & ~new_n2361_;
  assign new_n2363_ = ~new_n2359_ & new_n2362_;
  assign new_n2364_ = new_n587_ & new_n1881_;
  assign new_n2365_ = new_n587_ & new_n1864_;
  assign new_n2366_ = new_n587_ & new_n1878_;
  assign new_n2367_ = ~new_n2365_ & ~new_n2366_;
  assign new_n2368_ = ~new_n2364_ & new_n2367_;
  assign new_n2369_ = new_n2363_ & new_n2368_;
  assign new_n2370_ = new_n2358_ & new_n2369_;
  assign new_n2371_ = new_n2347_ & new_n2370_;
  assign new_n2372_ = new_n587_ & new_n1892_;
  assign new_n2373_ = new_n587_ & new_n1875_;
  assign new_n2374_ = new_n587_ & new_n1889_;
  assign new_n2375_ = ~new_n2373_ & ~new_n2374_;
  assign new_n2376_ = ~new_n2372_ & new_n2375_;
  assign new_n2377_ = new_n587_ & new_n1902_;
  assign new_n2378_ = new_n587_ & new_n1886_;
  assign new_n2379_ = new_n587_ & new_n1900_;
  assign new_n2380_ = ~new_n2378_ & ~new_n2379_;
  assign new_n2381_ = ~new_n2377_ & new_n2380_;
  assign new_n2382_ = new_n2376_ & new_n2381_;
  assign new_n2383_ = new_n586_ & new_n1975_;
  assign new_n2384_ = new_n1735_ & new_n2383_;
  assign new_n2385_ = new_n587_ & new_n1898_;
  assign new_n2386_ = new_n587_ & new_n1913_;
  assign new_n2387_ = ~new_n2385_ & ~new_n2386_;
  assign new_n2388_ = ~new_n2384_ & new_n2387_;
  assign new_n2389_ = new_n1749_ & new_n2383_;
  assign new_n2390_ = new_n1738_ & new_n2383_;
  assign new_n2391_ = new_n1725_ & new_n2383_;
  assign new_n2392_ = ~new_n2390_ & ~new_n2391_;
  assign new_n2393_ = ~new_n2389_ & new_n2392_;
  assign new_n2394_ = new_n2388_ & new_n2393_;
  assign new_n2395_ = new_n2382_ & new_n2394_;
  assign new_n2396_ = new_n586_ & new_n1986_;
  assign new_n2397_ = new_n1725_ & new_n2396_;
  assign new_n2398_ = new_n1735_ & new_n2396_;
  assign new_n2399_ = new_n1738_ & new_n2396_;
  assign new_n2400_ = ~new_n2398_ & ~new_n2399_;
  assign new_n2401_ = ~new_n2397_ & new_n2400_;
  assign new_n2402_ = new_n594_ & new_n1833_;
  assign new_n2403_ = new_n1749_ & new_n2396_;
  assign new_n2404_ = new_n594_ & new_n1830_;
  assign new_n2405_ = ~new_n2403_ & ~new_n2404_;
  assign new_n2406_ = ~new_n2402_ & new_n2405_;
  assign new_n2407_ = new_n2401_ & new_n2406_;
  assign new_n2408_ = new_n594_ & new_n1842_;
  assign new_n2409_ = new_n594_ & new_n1827_;
  assign new_n2410_ = new_n594_ & new_n1840_;
  assign new_n2411_ = ~new_n2409_ & ~new_n2410_;
  assign new_n2412_ = ~new_n2408_ & new_n2411_;
  assign new_n2413_ = new_n594_ & new_n1838_;
  assign new_n2414_ = new_n594_ & new_n1847_;
  assign new_n2415_ = ~new_n2413_ & ~new_n2414_;
  assign new_n2416_ = new_n2412_ & new_n2415_;
  assign new_n2417_ = new_n2407_ & new_n2416_;
  assign new_n2418_ = new_n2395_ & new_n2417_;
  assign new_n2419_ = new_n2371_ & new_n2418_;
  assign new_n2420_ = new_n594_ & new_n1859_;
  assign new_n2421_ = new_n594_ & new_n1849_;
  assign new_n2422_ = new_n594_ & new_n1857_;
  assign new_n2423_ = ~new_n2421_ & ~new_n2422_;
  assign new_n2424_ = ~new_n2420_ & new_n2423_;
  assign new_n2425_ = new_n594_ & new_n1868_;
  assign new_n2426_ = new_n594_ & new_n1855_;
  assign new_n2427_ = new_n594_ & new_n1866_;
  assign new_n2428_ = ~new_n2426_ & ~new_n2427_;
  assign new_n2429_ = ~new_n2425_ & new_n2428_;
  assign new_n2430_ = new_n2424_ & new_n2429_;
  assign new_n2431_ = new_n594_ & new_n1881_;
  assign new_n2432_ = new_n594_ & new_n1864_;
  assign new_n2433_ = new_n594_ & new_n1878_;
  assign new_n2434_ = ~new_n2432_ & ~new_n2433_;
  assign new_n2435_ = ~new_n2431_ & new_n2434_;
  assign new_n2436_ = new_n594_ & new_n1892_;
  assign new_n2437_ = new_n594_ & new_n1875_;
  assign new_n2438_ = new_n594_ & new_n1889_;
  assign new_n2439_ = ~new_n2437_ & ~new_n2438_;
  assign new_n2440_ = ~new_n2436_ & new_n2439_;
  assign new_n2441_ = new_n2435_ & new_n2440_;
  assign new_n2442_ = new_n2430_ & new_n2441_;
  assign new_n2443_ = new_n594_ & new_n1902_;
  assign new_n2444_ = new_n594_ & new_n1886_;
  assign new_n2445_ = new_n594_ & new_n1900_;
  assign new_n2446_ = ~new_n2444_ & ~new_n2445_;
  assign new_n2447_ = ~new_n2443_ & new_n2446_;
  assign new_n2448_ = new_n586_ & new_n2045_;
  assign new_n2449_ = new_n1735_ & new_n2448_;
  assign new_n2450_ = new_n594_ & new_n1898_;
  assign new_n2451_ = new_n594_ & new_n1913_;
  assign new_n2452_ = ~new_n2450_ & ~new_n2451_;
  assign new_n2453_ = ~new_n2449_ & new_n2452_;
  assign new_n2454_ = new_n2447_ & new_n2453_;
  assign new_n2455_ = new_n1749_ & new_n2448_;
  assign new_n2456_ = new_n1738_ & new_n2448_;
  assign new_n2457_ = new_n1725_ & new_n2448_;
  assign new_n2458_ = ~new_n2456_ & ~new_n2457_;
  assign new_n2459_ = ~new_n2455_ & new_n2458_;
  assign new_n2460_ = new_n586_ & new_n2052_;
  assign new_n2461_ = new_n1735_ & new_n2460_;
  assign new_n2462_ = new_n1738_ & new_n2460_;
  assign new_n2463_ = ~new_n2461_ & ~new_n2462_;
  assign new_n2464_ = new_n2459_ & new_n2463_;
  assign new_n2465_ = new_n2454_ & new_n2464_;
  assign new_n2466_ = new_n2442_ & new_n2465_;
  assign new_n2467_ = ~A166 & ~A167;
  assign new_n2468_ = new_n1908_ & new_n2467_;
  assign new_n2469_ = new_n1907_ & new_n2468_;
  assign new_n2470_ = new_n1735_ & new_n2469_;
  assign new_n2471_ = new_n1725_ & new_n2460_;
  assign new_n2472_ = new_n1749_ & new_n2460_;
  assign new_n2473_ = ~new_n2471_ & ~new_n2472_;
  assign new_n2474_ = ~new_n2470_ & new_n2473_;
  assign new_n2475_ = new_n1749_ & new_n2469_;
  assign new_n2476_ = new_n1738_ & new_n2469_;
  assign new_n2477_ = new_n1725_ & new_n2469_;
  assign new_n2478_ = ~new_n2476_ & ~new_n2477_;
  assign new_n2479_ = ~new_n2475_ & new_n2478_;
  assign new_n2480_ = new_n2474_ & new_n2479_;
  assign new_n2481_ = A166 & A167;
  assign new_n2482_ = new_n1908_ & new_n2481_;
  assign new_n2483_ = new_n1907_ & new_n2482_;
  assign new_n2484_ = new_n1725_ & new_n2483_;
  assign new_n2485_ = new_n1735_ & new_n2483_;
  assign new_n2486_ = new_n1738_ & new_n2483_;
  assign new_n2487_ = ~new_n2485_ & ~new_n2486_;
  assign new_n2488_ = ~new_n2484_ & new_n2487_;
  assign new_n2489_ = new_n601_ & new_n954_;
  assign new_n2490_ = new_n1749_ & new_n2483_;
  assign new_n2491_ = new_n601_ & new_n951_;
  assign new_n2492_ = ~new_n2490_ & ~new_n2491_;
  assign new_n2493_ = ~new_n2489_ & new_n2492_;
  assign new_n2494_ = new_n2488_ & new_n2493_;
  assign new_n2495_ = new_n2480_ & new_n2494_;
  assign new_n2496_ = new_n601_ & new_n967_;
  assign new_n2497_ = new_n601_ & new_n948_;
  assign new_n2498_ = new_n601_ & new_n964_;
  assign new_n2499_ = ~new_n2497_ & ~new_n2498_;
  assign new_n2500_ = ~new_n2496_ & new_n2499_;
  assign new_n2501_ = new_n601_ & new_n978_;
  assign new_n2502_ = new_n601_ & new_n961_;
  assign new_n2503_ = new_n601_ & new_n975_;
  assign new_n2504_ = ~new_n2502_ & ~new_n2503_;
  assign new_n2505_ = ~new_n2501_ & new_n2504_;
  assign new_n2506_ = new_n2500_ & new_n2505_;
  assign new_n2507_ = new_n601_ & new_n990_;
  assign new_n2508_ = new_n601_ & new_n972_;
  assign new_n2509_ = new_n601_ & new_n987_;
  assign new_n2510_ = ~new_n2508_ & ~new_n2509_;
  assign new_n2511_ = ~new_n2507_ & new_n2510_;
  assign new_n2512_ = new_n601_ & new_n984_;
  assign new_n2513_ = new_n601_ & new_n994_;
  assign new_n2514_ = ~new_n2512_ & ~new_n2513_;
  assign new_n2515_ = new_n2511_ & new_n2514_;
  assign new_n2516_ = new_n2506_ & new_n2515_;
  assign new_n2517_ = new_n2495_ & new_n2516_;
  assign new_n2518_ = new_n2466_ & new_n2517_;
  assign new_n2519_ = new_n2419_ & new_n2518_;
  assign new_n2520_ = new_n601_ & new_n1010_;
  assign new_n2521_ = new_n601_ & new_n996_;
  assign new_n2522_ = new_n601_ & new_n1008_;
  assign new_n2523_ = ~new_n2521_ & ~new_n2522_;
  assign new_n2524_ = ~new_n2520_ & new_n2523_;
  assign new_n2525_ = new_n601_ & new_n1018_;
  assign new_n2526_ = new_n601_ & new_n1006_;
  assign new_n2527_ = new_n601_ & new_n1016_;
  assign new_n2528_ = ~new_n2526_ & ~new_n2527_;
  assign new_n2529_ = ~new_n2525_ & new_n2528_;
  assign new_n2530_ = new_n2524_ & new_n2529_;
  assign new_n2531_ = new_n601_ & new_n1027_;
  assign new_n2532_ = new_n601_ & new_n1014_;
  assign new_n2533_ = new_n601_ & new_n1025_;
  assign new_n2534_ = ~new_n2532_ & ~new_n2533_;
  assign new_n2535_ = ~new_n2531_ & new_n2534_;
  assign new_n2536_ = new_n601_ & new_n1035_;
  assign new_n2537_ = new_n601_ & new_n1023_;
  assign new_n2538_ = new_n601_ & new_n1033_;
  assign new_n2539_ = ~new_n2537_ & ~new_n2538_;
  assign new_n2540_ = ~new_n2536_ & new_n2539_;
  assign new_n2541_ = new_n2535_ & new_n2540_;
  assign new_n2542_ = new_n2530_ & new_n2541_;
  assign new_n2543_ = new_n601_ & new_n1045_;
  assign new_n2544_ = new_n601_ & new_n1031_;
  assign new_n2545_ = new_n601_ & new_n1043_;
  assign new_n2546_ = ~new_n2544_ & ~new_n2545_;
  assign new_n2547_ = ~new_n2543_ & new_n2546_;
  assign new_n2548_ = new_n601_ & new_n1053_;
  assign new_n2549_ = new_n601_ & new_n1041_;
  assign new_n2550_ = new_n601_ & new_n1051_;
  assign new_n2551_ = ~new_n2549_ & ~new_n2550_;
  assign new_n2552_ = ~new_n2548_ & new_n2551_;
  assign new_n2553_ = new_n2547_ & new_n2552_;
  assign new_n2554_ = new_n650_ & new_n1071_;
  assign new_n2555_ = new_n601_ & new_n1049_;
  assign new_n2556_ = new_n650_ & new_n1065_;
  assign new_n2557_ = ~new_n2555_ & ~new_n2556_;
  assign new_n2558_ = ~new_n2554_ & new_n2557_;
  assign new_n2559_ = new_n650_ & new_n1059_;
  assign new_n2560_ = new_n650_ & new_n1079_;
  assign new_n2561_ = ~new_n2559_ & ~new_n2560_;
  assign new_n2562_ = new_n2558_ & new_n2561_;
  assign new_n2563_ = new_n2553_ & new_n2562_;
  assign new_n2564_ = new_n2542_ & new_n2563_;
  assign new_n2565_ = new_n650_ & new_n1095_;
  assign new_n2566_ = new_n650_ & new_n1082_;
  assign new_n2567_ = new_n650_ & new_n1076_;
  assign new_n2568_ = ~new_n2566_ & ~new_n2567_;
  assign new_n2569_ = ~new_n2565_ & new_n2568_;
  assign new_n2570_ = new_n650_ & new_n1105_;
  assign new_n2571_ = new_n650_ & new_n1099_;
  assign new_n2572_ = new_n650_ & new_n1089_;
  assign new_n2573_ = ~new_n2571_ & ~new_n2572_;
  assign new_n2574_ = ~new_n2570_ & new_n2573_;
  assign new_n2575_ = new_n2569_ & new_n2574_;
  assign new_n2576_ = new_n650_ & new_n1118_;
  assign new_n2577_ = new_n650_ & new_n1107_;
  assign new_n2578_ = new_n650_ & new_n1103_;
  assign new_n2579_ = ~new_n2577_ & ~new_n2578_;
  assign new_n2580_ = ~new_n2576_ & new_n2579_;
  assign new_n2581_ = new_n650_ & new_n1131_;
  assign new_n2582_ = new_n650_ & new_n1120_;
  assign new_n2583_ = new_n650_ & new_n1114_;
  assign new_n2584_ = ~new_n2582_ & ~new_n2583_;
  assign new_n2585_ = ~new_n2581_ & new_n2584_;
  assign new_n2586_ = new_n2580_ & new_n2585_;
  assign new_n2587_ = new_n2575_ & new_n2586_;
  assign new_n2588_ = new_n650_ & new_n1145_;
  assign new_n2589_ = new_n650_ & new_n1135_;
  assign new_n2590_ = new_n650_ & new_n1127_;
  assign new_n2591_ = ~new_n2589_ & ~new_n2590_;
  assign new_n2592_ = ~new_n2588_ & new_n2591_;
  assign new_n2593_ = new_n650_ & new_n1155_;
  assign new_n2594_ = new_n650_ & new_n1149_;
  assign new_n2595_ = new_n650_ & new_n1141_;
  assign new_n2596_ = ~new_n2594_ & ~new_n2595_;
  assign new_n2597_ = ~new_n2593_ & new_n2596_;
  assign new_n2598_ = new_n2592_ & new_n2597_;
  assign new_n2599_ = new_n650_ & new_n1165_;
  assign new_n2600_ = new_n650_ & new_n1157_;
  assign new_n2601_ = new_n650_ & new_n1153_;
  assign new_n2602_ = ~new_n2600_ & ~new_n2601_;
  assign new_n2603_ = ~new_n2599_ & new_n2602_;
  assign new_n2604_ = new_n650_ & new_n1168_;
  assign new_n2605_ = new_n650_ & new_n1162_;
  assign new_n2606_ = ~new_n2604_ & ~new_n2605_;
  assign new_n2607_ = new_n2603_ & new_n2606_;
  assign new_n2608_ = new_n2598_ & new_n2607_;
  assign new_n2609_ = new_n2587_ & new_n2608_;
  assign new_n2610_ = new_n2564_ & new_n2609_;
  assign new_n2611_ = new_n650_ & new_n1184_;
  assign new_n2612_ = new_n650_ & new_n1172_;
  assign new_n2613_ = new_n650_ & new_n1174_;
  assign new_n2614_ = ~new_n2612_ & ~new_n2613_;
  assign new_n2615_ = ~new_n2611_ & new_n2614_;
  assign new_n2616_ = new_n650_ & new_n1192_;
  assign new_n2617_ = new_n650_ & new_n1186_;
  assign new_n2618_ = new_n650_ & new_n1182_;
  assign new_n2619_ = ~new_n2617_ & ~new_n2618_;
  assign new_n2620_ = ~new_n2616_ & new_n2619_;
  assign new_n2621_ = new_n2615_ & new_n2620_;
  assign new_n2622_ = new_n650_ & new_n1202_;
  assign new_n2623_ = new_n650_ & new_n1194_;
  assign new_n2624_ = new_n650_ & new_n1190_;
  assign new_n2625_ = ~new_n2623_ & ~new_n2624_;
  assign new_n2626_ = ~new_n2622_ & new_n2625_;
  assign new_n2627_ = new_n650_ & new_n1213_;
  assign new_n2628_ = new_n650_ & new_n1204_;
  assign new_n2629_ = new_n650_ & new_n1200_;
  assign new_n2630_ = ~new_n2628_ & ~new_n2629_;
  assign new_n2631_ = ~new_n2627_ & new_n2630_;
  assign new_n2632_ = new_n2626_ & new_n2631_;
  assign new_n2633_ = new_n2621_ & new_n2632_;
  assign new_n2634_ = new_n650_ & new_n1226_;
  assign new_n2635_ = new_n650_ & new_n1216_;
  assign new_n2636_ = new_n650_ & new_n1210_;
  assign new_n2637_ = ~new_n2635_ & ~new_n2636_;
  assign new_n2638_ = ~new_n2634_ & new_n2637_;
  assign new_n2639_ = new_n650_ & new_n1235_;
  assign new_n2640_ = new_n650_ & new_n1229_;
  assign new_n2641_ = new_n650_ & new_n1223_;
  assign new_n2642_ = ~new_n2640_ & ~new_n2641_;
  assign new_n2643_ = ~new_n2639_ & new_n2642_;
  assign new_n2644_ = new_n2638_ & new_n2643_;
  assign new_n2645_ = new_n650_ & new_n1243_;
  assign new_n2646_ = new_n650_ & new_n1237_;
  assign new_n2647_ = new_n650_ & new_n1233_;
  assign new_n2648_ = ~new_n2646_ & ~new_n2647_;
  assign new_n2649_ = ~new_n2645_ & new_n2648_;
  assign new_n2650_ = new_n670_ & new_n951_;
  assign new_n2651_ = new_n670_ & new_n954_;
  assign new_n2652_ = ~new_n2650_ & ~new_n2651_;
  assign new_n2653_ = new_n2649_ & new_n2652_;
  assign new_n2654_ = new_n2644_ & new_n2653_;
  assign new_n2655_ = new_n2633_ & new_n2654_;
  assign new_n2656_ = new_n670_ & new_n967_;
  assign new_n2657_ = new_n670_ & new_n948_;
  assign new_n2658_ = new_n670_ & new_n964_;
  assign new_n2659_ = ~new_n2657_ & ~new_n2658_;
  assign new_n2660_ = ~new_n2656_ & new_n2659_;
  assign new_n2661_ = new_n670_ & new_n978_;
  assign new_n2662_ = new_n670_ & new_n961_;
  assign new_n2663_ = new_n670_ & new_n975_;
  assign new_n2664_ = ~new_n2662_ & ~new_n2663_;
  assign new_n2665_ = ~new_n2661_ & new_n2664_;
  assign new_n2666_ = new_n2660_ & new_n2665_;
  assign new_n2667_ = new_n670_ & new_n990_;
  assign new_n2668_ = new_n670_ & new_n972_;
  assign new_n2669_ = new_n670_ & new_n987_;
  assign new_n2670_ = ~new_n2668_ & ~new_n2669_;
  assign new_n2671_ = ~new_n2667_ & new_n2670_;
  assign new_n2672_ = new_n670_ & new_n996_;
  assign new_n2673_ = new_n670_ & new_n984_;
  assign new_n2674_ = new_n670_ & new_n994_;
  assign new_n2675_ = ~new_n2673_ & ~new_n2674_;
  assign new_n2676_ = ~new_n2672_ & new_n2675_;
  assign new_n2677_ = new_n2671_ & new_n2676_;
  assign new_n2678_ = new_n2666_ & new_n2677_;
  assign new_n2679_ = new_n670_ & new_n1006_;
  assign new_n2680_ = new_n670_ & new_n1008_;
  assign new_n2681_ = new_n670_ & new_n1010_;
  assign new_n2682_ = ~new_n2680_ & ~new_n2681_;
  assign new_n2683_ = ~new_n2679_ & new_n2682_;
  assign new_n2684_ = new_n670_ & new_n1014_;
  assign new_n2685_ = new_n670_ & new_n1016_;
  assign new_n2686_ = new_n670_ & new_n1018_;
  assign new_n2687_ = ~new_n2685_ & ~new_n2686_;
  assign new_n2688_ = ~new_n2684_ & new_n2687_;
  assign new_n2689_ = new_n2683_ & new_n2688_;
  assign new_n2690_ = new_n670_ & new_n1023_;
  assign new_n2691_ = new_n670_ & new_n1025_;
  assign new_n2692_ = new_n670_ & new_n1027_;
  assign new_n2693_ = ~new_n2691_ & ~new_n2692_;
  assign new_n2694_ = ~new_n2690_ & new_n2693_;
  assign new_n2695_ = new_n670_ & new_n1033_;
  assign new_n2696_ = new_n670_ & new_n1035_;
  assign new_n2697_ = ~new_n2695_ & ~new_n2696_;
  assign new_n2698_ = new_n2694_ & new_n2697_;
  assign new_n2699_ = new_n2689_ & new_n2698_;
  assign new_n2700_ = new_n2678_ & new_n2699_;
  assign new_n2701_ = new_n2655_ & new_n2700_;
  assign new_n2702_ = new_n2610_ & new_n2701_;
  assign new_n2703_ = new_n2519_ & new_n2702_;
  assign new_n2704_ = new_n2322_ & new_n2703_;
  assign new_n2705_ = new_n670_ & new_n1045_;
  assign new_n2706_ = new_n670_ & new_n1031_;
  assign new_n2707_ = new_n670_ & new_n1043_;
  assign new_n2708_ = ~new_n2706_ & ~new_n2707_;
  assign new_n2709_ = ~new_n2705_ & new_n2708_;
  assign new_n2710_ = new_n670_ & new_n1053_;
  assign new_n2711_ = new_n670_ & new_n1041_;
  assign new_n2712_ = new_n670_ & new_n1051_;
  assign new_n2713_ = ~new_n2711_ & ~new_n2712_;
  assign new_n2714_ = ~new_n2710_ & new_n2713_;
  assign new_n2715_ = new_n2709_ & new_n2714_;
  assign new_n2716_ = new_n718_ & new_n1071_;
  assign new_n2717_ = new_n670_ & new_n1049_;
  assign new_n2718_ = new_n718_ & new_n1065_;
  assign new_n2719_ = ~new_n2717_ & ~new_n2718_;
  assign new_n2720_ = ~new_n2716_ & new_n2719_;
  assign new_n2721_ = new_n718_ & new_n1082_;
  assign new_n2722_ = new_n718_ & new_n1059_;
  assign new_n2723_ = new_n718_ & new_n1079_;
  assign new_n2724_ = ~new_n2722_ & ~new_n2723_;
  assign new_n2725_ = ~new_n2721_ & new_n2724_;
  assign new_n2726_ = new_n2720_ & new_n2725_;
  assign new_n2727_ = new_n2715_ & new_n2726_;
  assign new_n2728_ = new_n718_ & new_n1099_;
  assign new_n2729_ = new_n718_ & new_n1076_;
  assign new_n2730_ = new_n718_ & new_n1095_;
  assign new_n2731_ = ~new_n2729_ & ~new_n2730_;
  assign new_n2732_ = ~new_n2728_ & new_n2731_;
  assign new_n2733_ = new_n718_ & new_n1107_;
  assign new_n2734_ = new_n718_ & new_n1089_;
  assign new_n2735_ = new_n718_ & new_n1105_;
  assign new_n2736_ = ~new_n2734_ & ~new_n2735_;
  assign new_n2737_ = ~new_n2733_ & new_n2736_;
  assign new_n2738_ = new_n2732_ & new_n2737_;
  assign new_n2739_ = new_n718_ & new_n1120_;
  assign new_n2740_ = new_n718_ & new_n1103_;
  assign new_n2741_ = new_n718_ & new_n1118_;
  assign new_n2742_ = ~new_n2740_ & ~new_n2741_;
  assign new_n2743_ = ~new_n2739_ & new_n2742_;
  assign new_n2744_ = new_n718_ & new_n1135_;
  assign new_n2745_ = new_n718_ & new_n1114_;
  assign new_n2746_ = new_n718_ & new_n1131_;
  assign new_n2747_ = ~new_n2745_ & ~new_n2746_;
  assign new_n2748_ = ~new_n2744_ & new_n2747_;
  assign new_n2749_ = new_n2743_ & new_n2748_;
  assign new_n2750_ = new_n2738_ & new_n2749_;
  assign new_n2751_ = new_n2727_ & new_n2750_;
  assign new_n2752_ = new_n718_ & new_n1149_;
  assign new_n2753_ = new_n718_ & new_n1127_;
  assign new_n2754_ = new_n718_ & new_n1145_;
  assign new_n2755_ = ~new_n2753_ & ~new_n2754_;
  assign new_n2756_ = ~new_n2752_ & new_n2755_;
  assign new_n2757_ = new_n718_ & new_n1157_;
  assign new_n2758_ = new_n718_ & new_n1141_;
  assign new_n2759_ = new_n718_ & new_n1155_;
  assign new_n2760_ = ~new_n2758_ & ~new_n2759_;
  assign new_n2761_ = ~new_n2757_ & new_n2760_;
  assign new_n2762_ = new_n2756_ & new_n2761_;
  assign new_n2763_ = new_n718_ & new_n1168_;
  assign new_n2764_ = new_n718_ & new_n1153_;
  assign new_n2765_ = new_n718_ & new_n1165_;
  assign new_n2766_ = ~new_n2764_ & ~new_n2765_;
  assign new_n2767_ = ~new_n2763_ & new_n2766_;
  assign new_n2768_ = new_n718_ & new_n1174_;
  assign new_n2769_ = new_n718_ & new_n1162_;
  assign new_n2770_ = new_n718_ & new_n1172_;
  assign new_n2771_ = ~new_n2769_ & ~new_n2770_;
  assign new_n2772_ = ~new_n2768_ & new_n2771_;
  assign new_n2773_ = new_n2767_ & new_n2772_;
  assign new_n2774_ = new_n2762_ & new_n2773_;
  assign new_n2775_ = new_n718_ & new_n1182_;
  assign new_n2776_ = new_n718_ & new_n1184_;
  assign new_n2777_ = new_n718_ & new_n1186_;
  assign new_n2778_ = ~new_n2776_ & ~new_n2777_;
  assign new_n2779_ = ~new_n2775_ & new_n2778_;
  assign new_n2780_ = new_n718_ & new_n1190_;
  assign new_n2781_ = new_n718_ & new_n1192_;
  assign new_n2782_ = new_n718_ & new_n1194_;
  assign new_n2783_ = ~new_n2781_ & ~new_n2782_;
  assign new_n2784_ = ~new_n2780_ & new_n2783_;
  assign new_n2785_ = new_n2779_ & new_n2784_;
  assign new_n2786_ = new_n718_ & new_n1200_;
  assign new_n2787_ = new_n718_ & new_n1202_;
  assign new_n2788_ = new_n718_ & new_n1204_;
  assign new_n2789_ = ~new_n2787_ & ~new_n2788_;
  assign new_n2790_ = ~new_n2786_ & new_n2789_;
  assign new_n2791_ = new_n718_ & new_n1213_;
  assign new_n2792_ = new_n718_ & new_n1216_;
  assign new_n2793_ = ~new_n2791_ & ~new_n2792_;
  assign new_n2794_ = new_n2790_ & new_n2793_;
  assign new_n2795_ = new_n2785_ & new_n2794_;
  assign new_n2796_ = new_n2774_ & new_n2795_;
  assign new_n2797_ = new_n2751_ & new_n2796_;
  assign new_n2798_ = new_n718_ & new_n1229_;
  assign new_n2799_ = new_n718_ & new_n1210_;
  assign new_n2800_ = new_n718_ & new_n1226_;
  assign new_n2801_ = ~new_n2799_ & ~new_n2800_;
  assign new_n2802_ = ~new_n2798_ & new_n2801_;
  assign new_n2803_ = new_n718_ & new_n1237_;
  assign new_n2804_ = new_n718_ & new_n1223_;
  assign new_n2805_ = new_n718_ & new_n1235_;
  assign new_n2806_ = ~new_n2804_ & ~new_n2805_;
  assign new_n2807_ = ~new_n2803_ & new_n2806_;
  assign new_n2808_ = new_n2802_ & new_n2807_;
  assign new_n2809_ = new_n737_ & new_n1830_;
  assign new_n2810_ = new_n718_ & new_n1233_;
  assign new_n2811_ = new_n718_ & new_n1243_;
  assign new_n2812_ = ~new_n2810_ & ~new_n2811_;
  assign new_n2813_ = ~new_n2809_ & new_n2812_;
  assign new_n2814_ = new_n737_ & new_n1840_;
  assign new_n2815_ = new_n737_ & new_n1833_;
  assign new_n2816_ = new_n737_ & new_n1827_;
  assign new_n2817_ = ~new_n2815_ & ~new_n2816_;
  assign new_n2818_ = ~new_n2814_ & new_n2817_;
  assign new_n2819_ = new_n2813_ & new_n2818_;
  assign new_n2820_ = new_n2808_ & new_n2819_;
  assign new_n2821_ = new_n737_ & new_n1847_;
  assign new_n2822_ = new_n737_ & new_n1842_;
  assign new_n2823_ = new_n737_ & new_n1838_;
  assign new_n2824_ = ~new_n2822_ & ~new_n2823_;
  assign new_n2825_ = ~new_n2821_ & new_n2824_;
  assign new_n2826_ = new_n737_ & new_n1859_;
  assign new_n2827_ = new_n737_ & new_n1849_;
  assign new_n2828_ = new_n737_ & new_n1857_;
  assign new_n2829_ = ~new_n2827_ & ~new_n2828_;
  assign new_n2830_ = ~new_n2826_ & new_n2829_;
  assign new_n2831_ = new_n2825_ & new_n2830_;
  assign new_n2832_ = new_n737_ & new_n1868_;
  assign new_n2833_ = new_n737_ & new_n1855_;
  assign new_n2834_ = new_n737_ & new_n1866_;
  assign new_n2835_ = ~new_n2833_ & ~new_n2834_;
  assign new_n2836_ = ~new_n2832_ & new_n2835_;
  assign new_n2837_ = new_n737_ & new_n1864_;
  assign new_n2838_ = new_n737_ & new_n1878_;
  assign new_n2839_ = ~new_n2837_ & ~new_n2838_;
  assign new_n2840_ = new_n2836_ & new_n2839_;
  assign new_n2841_ = new_n2831_ & new_n2840_;
  assign new_n2842_ = new_n2820_ & new_n2841_;
  assign new_n2843_ = new_n737_ & new_n1889_;
  assign new_n2844_ = new_n737_ & new_n1881_;
  assign new_n2845_ = new_n737_ & new_n1875_;
  assign new_n2846_ = ~new_n2844_ & ~new_n2845_;
  assign new_n2847_ = ~new_n2843_ & new_n2846_;
  assign new_n2848_ = new_n737_ & new_n1900_;
  assign new_n2849_ = new_n737_ & new_n1892_;
  assign new_n2850_ = new_n737_ & new_n1886_;
  assign new_n2851_ = ~new_n2849_ & ~new_n2850_;
  assign new_n2852_ = ~new_n2848_ & new_n2851_;
  assign new_n2853_ = new_n2847_ & new_n2852_;
  assign new_n2854_ = new_n737_ & new_n1913_;
  assign new_n2855_ = new_n737_ & new_n1902_;
  assign new_n2856_ = new_n737_ & new_n1898_;
  assign new_n2857_ = ~new_n2855_ & ~new_n2856_;
  assign new_n2858_ = ~new_n2854_ & new_n2857_;
  assign new_n2859_ = new_n736_ & new_n1975_;
  assign new_n2860_ = new_n1725_ & new_n2859_;
  assign new_n2861_ = new_n1735_ & new_n2859_;
  assign new_n2862_ = new_n1738_ & new_n2859_;
  assign new_n2863_ = ~new_n2861_ & ~new_n2862_;
  assign new_n2864_ = ~new_n2860_ & new_n2863_;
  assign new_n2865_ = new_n2858_ & new_n2864_;
  assign new_n2866_ = new_n2853_ & new_n2865_;
  assign new_n2867_ = new_n736_ & new_n1986_;
  assign new_n2868_ = new_n1738_ & new_n2867_;
  assign new_n2869_ = new_n1749_ & new_n2859_;
  assign new_n2870_ = new_n1735_ & new_n2867_;
  assign new_n2871_ = ~new_n2869_ & ~new_n2870_;
  assign new_n2872_ = ~new_n2868_ & new_n2871_;
  assign new_n2873_ = new_n749_ & new_n1830_;
  assign new_n2874_ = new_n1725_ & new_n2867_;
  assign new_n2875_ = new_n1749_ & new_n2867_;
  assign new_n2876_ = ~new_n2874_ & ~new_n2875_;
  assign new_n2877_ = ~new_n2873_ & new_n2876_;
  assign new_n2878_ = new_n2872_ & new_n2877_;
  assign new_n2879_ = new_n749_ & new_n1840_;
  assign new_n2880_ = new_n749_ & new_n1833_;
  assign new_n2881_ = new_n749_ & new_n1827_;
  assign new_n2882_ = ~new_n2880_ & ~new_n2881_;
  assign new_n2883_ = ~new_n2879_ & new_n2882_;
  assign new_n2884_ = new_n749_ & new_n1842_;
  assign new_n2885_ = new_n749_ & new_n1838_;
  assign new_n2886_ = ~new_n2884_ & ~new_n2885_;
  assign new_n2887_ = new_n2883_ & new_n2886_;
  assign new_n2888_ = new_n2878_ & new_n2887_;
  assign new_n2889_ = new_n2866_ & new_n2888_;
  assign new_n2890_ = new_n2842_ & new_n2889_;
  assign new_n2891_ = new_n2797_ & new_n2890_;
  assign new_n2892_ = new_n749_ & new_n1857_;
  assign new_n2893_ = new_n749_ & new_n1847_;
  assign new_n2894_ = new_n749_ & new_n1849_;
  assign new_n2895_ = ~new_n2893_ & ~new_n2894_;
  assign new_n2896_ = ~new_n2892_ & new_n2895_;
  assign new_n2897_ = new_n749_ & new_n1866_;
  assign new_n2898_ = new_n749_ & new_n1859_;
  assign new_n2899_ = new_n749_ & new_n1855_;
  assign new_n2900_ = ~new_n2898_ & ~new_n2899_;
  assign new_n2901_ = ~new_n2897_ & new_n2900_;
  assign new_n2902_ = new_n2896_ & new_n2901_;
  assign new_n2903_ = new_n749_ & new_n1878_;
  assign new_n2904_ = new_n749_ & new_n1868_;
  assign new_n2905_ = new_n749_ & new_n1864_;
  assign new_n2906_ = ~new_n2904_ & ~new_n2905_;
  assign new_n2907_ = ~new_n2903_ & new_n2906_;
  assign new_n2908_ = new_n749_ & new_n1889_;
  assign new_n2909_ = new_n749_ & new_n1881_;
  assign new_n2910_ = new_n749_ & new_n1875_;
  assign new_n2911_ = ~new_n2909_ & ~new_n2910_;
  assign new_n2912_ = ~new_n2908_ & new_n2911_;
  assign new_n2913_ = new_n2907_ & new_n2912_;
  assign new_n2914_ = new_n2902_ & new_n2913_;
  assign new_n2915_ = new_n749_ & new_n1900_;
  assign new_n2916_ = new_n749_ & new_n1892_;
  assign new_n2917_ = new_n749_ & new_n1886_;
  assign new_n2918_ = ~new_n2916_ & ~new_n2917_;
  assign new_n2919_ = ~new_n2915_ & new_n2918_;
  assign new_n2920_ = new_n749_ & new_n1913_;
  assign new_n2921_ = new_n749_ & new_n1902_;
  assign new_n2922_ = new_n749_ & new_n1898_;
  assign new_n2923_ = ~new_n2921_ & ~new_n2922_;
  assign new_n2924_ = ~new_n2920_ & new_n2923_;
  assign new_n2925_ = new_n2919_ & new_n2924_;
  assign new_n2926_ = new_n736_ & new_n2045_;
  assign new_n2927_ = new_n1725_ & new_n2926_;
  assign new_n2928_ = new_n1735_ & new_n2926_;
  assign new_n2929_ = new_n1738_ & new_n2926_;
  assign new_n2930_ = ~new_n2928_ & ~new_n2929_;
  assign new_n2931_ = ~new_n2927_ & new_n2930_;
  assign new_n2932_ = new_n1749_ & new_n2926_;
  assign new_n2933_ = new_n736_ & new_n2052_;
  assign new_n2934_ = new_n1735_ & new_n2933_;
  assign new_n2935_ = ~new_n2932_ & ~new_n2934_;
  assign new_n2936_ = new_n2931_ & new_n2935_;
  assign new_n2937_ = new_n2925_ & new_n2936_;
  assign new_n2938_ = new_n2914_ & new_n2937_;
  assign new_n2939_ = new_n1749_ & new_n2933_;
  assign new_n2940_ = new_n1738_ & new_n2933_;
  assign new_n2941_ = new_n1725_ & new_n2933_;
  assign new_n2942_ = ~new_n2940_ & ~new_n2941_;
  assign new_n2943_ = ~new_n2939_ & new_n2942_;
  assign new_n2944_ = new_n759_ & new_n1827_;
  assign new_n2945_ = new_n759_ & new_n1830_;
  assign new_n2946_ = new_n759_ & new_n1833_;
  assign new_n2947_ = ~new_n2945_ & ~new_n2946_;
  assign new_n2948_ = ~new_n2944_ & new_n2947_;
  assign new_n2949_ = new_n2943_ & new_n2948_;
  assign new_n2950_ = new_n759_ & new_n1838_;
  assign new_n2951_ = new_n759_ & new_n1840_;
  assign new_n2952_ = new_n759_ & new_n1842_;
  assign new_n2953_ = ~new_n2951_ & ~new_n2952_;
  assign new_n2954_ = ~new_n2950_ & new_n2953_;
  assign new_n2955_ = new_n759_ & new_n1857_;
  assign new_n2956_ = new_n759_ & new_n1847_;
  assign new_n2957_ = new_n759_ & new_n1849_;
  assign new_n2958_ = ~new_n2956_ & ~new_n2957_;
  assign new_n2959_ = ~new_n2955_ & new_n2958_;
  assign new_n2960_ = new_n2954_ & new_n2959_;
  assign new_n2961_ = new_n2949_ & new_n2960_;
  assign new_n2962_ = new_n759_ & new_n1866_;
  assign new_n2963_ = new_n759_ & new_n1859_;
  assign new_n2964_ = new_n759_ & new_n1855_;
  assign new_n2965_ = ~new_n2963_ & ~new_n2964_;
  assign new_n2966_ = ~new_n2962_ & new_n2965_;
  assign new_n2967_ = new_n759_ & new_n1878_;
  assign new_n2968_ = new_n759_ & new_n1868_;
  assign new_n2969_ = new_n759_ & new_n1864_;
  assign new_n2970_ = ~new_n2968_ & ~new_n2969_;
  assign new_n2971_ = ~new_n2967_ & new_n2970_;
  assign new_n2972_ = new_n2966_ & new_n2971_;
  assign new_n2973_ = new_n759_ & new_n1889_;
  assign new_n2974_ = new_n759_ & new_n1881_;
  assign new_n2975_ = new_n759_ & new_n1875_;
  assign new_n2976_ = ~new_n2974_ & ~new_n2975_;
  assign new_n2977_ = ~new_n2973_ & new_n2976_;
  assign new_n2978_ = new_n759_ & new_n1892_;
  assign new_n2979_ = new_n759_ & new_n1886_;
  assign new_n2980_ = ~new_n2978_ & ~new_n2979_;
  assign new_n2981_ = new_n2977_ & new_n2980_;
  assign new_n2982_ = new_n2972_ & new_n2981_;
  assign new_n2983_ = new_n2961_ & new_n2982_;
  assign new_n2984_ = new_n2938_ & new_n2983_;
  assign new_n2985_ = new_n759_ & new_n1898_;
  assign new_n2986_ = new_n759_ & new_n1900_;
  assign new_n2987_ = new_n759_ & new_n1902_;
  assign new_n2988_ = ~new_n2986_ & ~new_n2987_;
  assign new_n2989_ = ~new_n2985_ & new_n2988_;
  assign new_n2990_ = new_n758_ & new_n1975_;
  assign new_n2991_ = new_n1738_ & new_n2990_;
  assign new_n2992_ = new_n759_ & new_n1913_;
  assign new_n2993_ = new_n1735_ & new_n2990_;
  assign new_n2994_ = ~new_n2992_ & ~new_n2993_;
  assign new_n2995_ = ~new_n2991_ & new_n2994_;
  assign new_n2996_ = new_n2989_ & new_n2995_;
  assign new_n2997_ = new_n758_ & new_n1986_;
  assign new_n2998_ = new_n1735_ & new_n2997_;
  assign new_n2999_ = new_n1725_ & new_n2990_;
  assign new_n3000_ = new_n1749_ & new_n2990_;
  assign new_n3001_ = ~new_n2999_ & ~new_n3000_;
  assign new_n3002_ = ~new_n2998_ & new_n3001_;
  assign new_n3003_ = new_n1749_ & new_n2997_;
  assign new_n3004_ = new_n1738_ & new_n2997_;
  assign new_n3005_ = new_n1725_ & new_n2997_;
  assign new_n3006_ = ~new_n3004_ & ~new_n3005_;
  assign new_n3007_ = ~new_n3003_ & new_n3006_;
  assign new_n3008_ = new_n3002_ & new_n3007_;
  assign new_n3009_ = new_n2996_ & new_n3008_;
  assign new_n3010_ = new_n765_ & new_n1827_;
  assign new_n3011_ = new_n765_ & new_n1830_;
  assign new_n3012_ = new_n765_ & new_n1833_;
  assign new_n3013_ = ~new_n3011_ & ~new_n3012_;
  assign new_n3014_ = ~new_n3010_ & new_n3013_;
  assign new_n3015_ = new_n765_ & new_n1838_;
  assign new_n3016_ = new_n765_ & new_n1840_;
  assign new_n3017_ = new_n765_ & new_n1842_;
  assign new_n3018_ = ~new_n3016_ & ~new_n3017_;
  assign new_n3019_ = ~new_n3015_ & new_n3018_;
  assign new_n3020_ = new_n3014_ & new_n3019_;
  assign new_n3021_ = new_n765_ & new_n1857_;
  assign new_n3022_ = new_n765_ & new_n1847_;
  assign new_n3023_ = new_n765_ & new_n1849_;
  assign new_n3024_ = ~new_n3022_ & ~new_n3023_;
  assign new_n3025_ = ~new_n3021_ & new_n3024_;
  assign new_n3026_ = new_n765_ & new_n1859_;
  assign new_n3027_ = new_n765_ & new_n1855_;
  assign new_n3028_ = ~new_n3026_ & ~new_n3027_;
  assign new_n3029_ = new_n3025_ & new_n3028_;
  assign new_n3030_ = new_n3020_ & new_n3029_;
  assign new_n3031_ = new_n3009_ & new_n3030_;
  assign new_n3032_ = new_n765_ & new_n1864_;
  assign new_n3033_ = new_n765_ & new_n1866_;
  assign new_n3034_ = new_n765_ & new_n1868_;
  assign new_n3035_ = ~new_n3033_ & ~new_n3034_;
  assign new_n3036_ = ~new_n3032_ & new_n3035_;
  assign new_n3037_ = new_n765_ & new_n1875_;
  assign new_n3038_ = new_n765_ & new_n1878_;
  assign new_n3039_ = new_n765_ & new_n1881_;
  assign new_n3040_ = ~new_n3038_ & ~new_n3039_;
  assign new_n3041_ = ~new_n3037_ & new_n3040_;
  assign new_n3042_ = new_n3036_ & new_n3041_;
  assign new_n3043_ = new_n765_ & new_n1886_;
  assign new_n3044_ = new_n765_ & new_n1889_;
  assign new_n3045_ = new_n765_ & new_n1892_;
  assign new_n3046_ = ~new_n3044_ & ~new_n3045_;
  assign new_n3047_ = ~new_n3043_ & new_n3046_;
  assign new_n3048_ = new_n765_ & new_n1898_;
  assign new_n3049_ = new_n765_ & new_n1900_;
  assign new_n3050_ = new_n765_ & new_n1902_;
  assign new_n3051_ = ~new_n3049_ & ~new_n3050_;
  assign new_n3052_ = ~new_n3048_ & new_n3051_;
  assign new_n3053_ = new_n3047_ & new_n3052_;
  assign new_n3054_ = new_n3042_ & new_n3053_;
  assign new_n3055_ = new_n758_ & new_n2045_;
  assign new_n3056_ = new_n1738_ & new_n3055_;
  assign new_n3057_ = new_n765_ & new_n1913_;
  assign new_n3058_ = new_n1735_ & new_n3055_;
  assign new_n3059_ = ~new_n3057_ & ~new_n3058_;
  assign new_n3060_ = ~new_n3056_ & new_n3059_;
  assign new_n3061_ = new_n758_ & new_n2052_;
  assign new_n3062_ = new_n1735_ & new_n3061_;
  assign new_n3063_ = new_n1725_ & new_n3055_;
  assign new_n3064_ = new_n1749_ & new_n3055_;
  assign new_n3065_ = ~new_n3063_ & ~new_n3064_;
  assign new_n3066_ = ~new_n3062_ & new_n3065_;
  assign new_n3067_ = new_n3060_ & new_n3066_;
  assign new_n3068_ = new_n1749_ & new_n3061_;
  assign new_n3069_ = new_n1738_ & new_n3061_;
  assign new_n3070_ = new_n1725_ & new_n3061_;
  assign new_n3071_ = ~new_n3069_ & ~new_n3070_;
  assign new_n3072_ = ~new_n3068_ & new_n3071_;
  assign new_n3073_ = new_n777_ & new_n951_;
  assign new_n3074_ = new_n777_ & new_n954_;
  assign new_n3075_ = ~new_n3073_ & ~new_n3074_;
  assign new_n3076_ = new_n3072_ & new_n3075_;
  assign new_n3077_ = new_n3067_ & new_n3076_;
  assign new_n3078_ = new_n3054_ & new_n3077_;
  assign new_n3079_ = new_n3031_ & new_n3078_;
  assign new_n3080_ = new_n2984_ & new_n3079_;
  assign new_n3081_ = new_n2891_ & new_n3080_;
  assign new_n3082_ = new_n777_ & new_n967_;
  assign new_n3083_ = new_n777_ & new_n948_;
  assign new_n3084_ = new_n777_ & new_n964_;
  assign new_n3085_ = ~new_n3083_ & ~new_n3084_;
  assign new_n3086_ = ~new_n3082_ & new_n3085_;
  assign new_n3087_ = new_n777_ & new_n978_;
  assign new_n3088_ = new_n777_ & new_n961_;
  assign new_n3089_ = new_n777_ & new_n975_;
  assign new_n3090_ = ~new_n3088_ & ~new_n3089_;
  assign new_n3091_ = ~new_n3087_ & new_n3090_;
  assign new_n3092_ = new_n3086_ & new_n3091_;
  assign new_n3093_ = new_n777_ & new_n990_;
  assign new_n3094_ = new_n777_ & new_n972_;
  assign new_n3095_ = new_n777_ & new_n987_;
  assign new_n3096_ = ~new_n3094_ & ~new_n3095_;
  assign new_n3097_ = ~new_n3093_ & new_n3096_;
  assign new_n3098_ = new_n777_ & new_n996_;
  assign new_n3099_ = new_n777_ & new_n984_;
  assign new_n3100_ = new_n777_ & new_n994_;
  assign new_n3101_ = ~new_n3099_ & ~new_n3100_;
  assign new_n3102_ = ~new_n3098_ & new_n3101_;
  assign new_n3103_ = new_n3097_ & new_n3102_;
  assign new_n3104_ = new_n3092_ & new_n3103_;
  assign new_n3105_ = new_n777_ & new_n1006_;
  assign new_n3106_ = new_n777_ & new_n1008_;
  assign new_n3107_ = new_n777_ & new_n1010_;
  assign new_n3108_ = ~new_n3106_ & ~new_n3107_;
  assign new_n3109_ = ~new_n3105_ & new_n3108_;
  assign new_n3110_ = new_n777_ & new_n1014_;
  assign new_n3111_ = new_n777_ & new_n1016_;
  assign new_n3112_ = new_n777_ & new_n1018_;
  assign new_n3113_ = ~new_n3111_ & ~new_n3112_;
  assign new_n3114_ = ~new_n3110_ & new_n3113_;
  assign new_n3115_ = new_n3109_ & new_n3114_;
  assign new_n3116_ = new_n777_ & new_n1023_;
  assign new_n3117_ = new_n777_ & new_n1025_;
  assign new_n3118_ = new_n777_ & new_n1027_;
  assign new_n3119_ = ~new_n3117_ & ~new_n3118_;
  assign new_n3120_ = ~new_n3116_ & new_n3119_;
  assign new_n3121_ = new_n777_ & new_n1033_;
  assign new_n3122_ = new_n777_ & new_n1035_;
  assign new_n3123_ = ~new_n3121_ & ~new_n3122_;
  assign new_n3124_ = new_n3120_ & new_n3123_;
  assign new_n3125_ = new_n3115_ & new_n3124_;
  assign new_n3126_ = new_n3104_ & new_n3125_;
  assign new_n3127_ = new_n777_ & new_n1045_;
  assign new_n3128_ = new_n777_ & new_n1031_;
  assign new_n3129_ = new_n777_ & new_n1043_;
  assign new_n3130_ = ~new_n3128_ & ~new_n3129_;
  assign new_n3131_ = ~new_n3127_ & new_n3130_;
  assign new_n3132_ = new_n777_ & new_n1053_;
  assign new_n3133_ = new_n777_ & new_n1041_;
  assign new_n3134_ = new_n777_ & new_n1051_;
  assign new_n3135_ = ~new_n3133_ & ~new_n3134_;
  assign new_n3136_ = ~new_n3132_ & new_n3135_;
  assign new_n3137_ = new_n3131_ & new_n3136_;
  assign new_n3138_ = new_n826_ & new_n1071_;
  assign new_n3139_ = new_n777_ & new_n1049_;
  assign new_n3140_ = new_n826_ & new_n1065_;
  assign new_n3141_ = ~new_n3139_ & ~new_n3140_;
  assign new_n3142_ = ~new_n3138_ & new_n3141_;
  assign new_n3143_ = new_n826_ & new_n1082_;
  assign new_n3144_ = new_n826_ & new_n1059_;
  assign new_n3145_ = new_n826_ & new_n1079_;
  assign new_n3146_ = ~new_n3144_ & ~new_n3145_;
  assign new_n3147_ = ~new_n3143_ & new_n3146_;
  assign new_n3148_ = new_n3142_ & new_n3147_;
  assign new_n3149_ = new_n3137_ & new_n3148_;
  assign new_n3150_ = new_n826_ & new_n1099_;
  assign new_n3151_ = new_n826_ & new_n1076_;
  assign new_n3152_ = new_n826_ & new_n1095_;
  assign new_n3153_ = ~new_n3151_ & ~new_n3152_;
  assign new_n3154_ = ~new_n3150_ & new_n3153_;
  assign new_n3155_ = new_n826_ & new_n1107_;
  assign new_n3156_ = new_n826_ & new_n1089_;
  assign new_n3157_ = new_n826_ & new_n1105_;
  assign new_n3158_ = ~new_n3156_ & ~new_n3157_;
  assign new_n3159_ = ~new_n3155_ & new_n3158_;
  assign new_n3160_ = new_n3154_ & new_n3159_;
  assign new_n3161_ = new_n826_ & new_n1120_;
  assign new_n3162_ = new_n826_ & new_n1103_;
  assign new_n3163_ = new_n826_ & new_n1118_;
  assign new_n3164_ = ~new_n3162_ & ~new_n3163_;
  assign new_n3165_ = ~new_n3161_ & new_n3164_;
  assign new_n3166_ = new_n826_ & new_n1114_;
  assign new_n3167_ = new_n826_ & new_n1131_;
  assign new_n3168_ = ~new_n3166_ & ~new_n3167_;
  assign new_n3169_ = new_n3165_ & new_n3168_;
  assign new_n3170_ = new_n3160_ & new_n3169_;
  assign new_n3171_ = new_n3149_ & new_n3170_;
  assign new_n3172_ = new_n3126_ & new_n3171_;
  assign new_n3173_ = new_n826_ & new_n1145_;
  assign new_n3174_ = new_n826_ & new_n1135_;
  assign new_n3175_ = new_n826_ & new_n1127_;
  assign new_n3176_ = ~new_n3174_ & ~new_n3175_;
  assign new_n3177_ = ~new_n3173_ & new_n3176_;
  assign new_n3178_ = new_n826_ & new_n1155_;
  assign new_n3179_ = new_n826_ & new_n1149_;
  assign new_n3180_ = new_n826_ & new_n1141_;
  assign new_n3181_ = ~new_n3179_ & ~new_n3180_;
  assign new_n3182_ = ~new_n3178_ & new_n3181_;
  assign new_n3183_ = new_n3177_ & new_n3182_;
  assign new_n3184_ = new_n826_ & new_n1165_;
  assign new_n3185_ = new_n826_ & new_n1157_;
  assign new_n3186_ = new_n826_ & new_n1153_;
  assign new_n3187_ = ~new_n3185_ & ~new_n3186_;
  assign new_n3188_ = ~new_n3184_ & new_n3187_;
  assign new_n3189_ = new_n826_ & new_n1172_;
  assign new_n3190_ = new_n826_ & new_n1168_;
  assign new_n3191_ = new_n826_ & new_n1162_;
  assign new_n3192_ = ~new_n3190_ & ~new_n3191_;
  assign new_n3193_ = ~new_n3189_ & new_n3192_;
  assign new_n3194_ = new_n3188_ & new_n3193_;
  assign new_n3195_ = new_n3183_ & new_n3194_;
  assign new_n3196_ = new_n826_ & new_n1186_;
  assign new_n3197_ = new_n826_ & new_n1174_;
  assign new_n3198_ = new_n826_ & new_n1184_;
  assign new_n3199_ = ~new_n3197_ & ~new_n3198_;
  assign new_n3200_ = ~new_n3196_ & new_n3199_;
  assign new_n3201_ = new_n826_ & new_n1194_;
  assign new_n3202_ = new_n826_ & new_n1182_;
  assign new_n3203_ = new_n826_ & new_n1192_;
  assign new_n3204_ = ~new_n3202_ & ~new_n3203_;
  assign new_n3205_ = ~new_n3201_ & new_n3204_;
  assign new_n3206_ = new_n3200_ & new_n3205_;
  assign new_n3207_ = new_n826_ & new_n1204_;
  assign new_n3208_ = new_n826_ & new_n1190_;
  assign new_n3209_ = new_n826_ & new_n1202_;
  assign new_n3210_ = ~new_n3208_ & ~new_n3209_;
  assign new_n3211_ = ~new_n3207_ & new_n3210_;
  assign new_n3212_ = new_n826_ & new_n1200_;
  assign new_n3213_ = new_n826_ & new_n1213_;
  assign new_n3214_ = ~new_n3212_ & ~new_n3213_;
  assign new_n3215_ = new_n3211_ & new_n3214_;
  assign new_n3216_ = new_n3206_ & new_n3215_;
  assign new_n3217_ = new_n3195_ & new_n3216_;
  assign new_n3218_ = new_n826_ & new_n1226_;
  assign new_n3219_ = new_n826_ & new_n1216_;
  assign new_n3220_ = new_n826_ & new_n1210_;
  assign new_n3221_ = ~new_n3219_ & ~new_n3220_;
  assign new_n3222_ = ~new_n3218_ & new_n3221_;
  assign new_n3223_ = new_n826_ & new_n1235_;
  assign new_n3224_ = new_n826_ & new_n1229_;
  assign new_n3225_ = new_n826_ & new_n1223_;
  assign new_n3226_ = ~new_n3224_ & ~new_n3225_;
  assign new_n3227_ = ~new_n3223_ & new_n3226_;
  assign new_n3228_ = new_n3222_ & new_n3227_;
  assign new_n3229_ = new_n826_ & new_n1243_;
  assign new_n3230_ = new_n826_ & new_n1237_;
  assign new_n3231_ = new_n826_ & new_n1233_;
  assign new_n3232_ = ~new_n3230_ & ~new_n3231_;
  assign new_n3233_ = ~new_n3229_ & new_n3232_;
  assign new_n3234_ = new_n843_ & new_n948_;
  assign new_n3235_ = new_n843_ & new_n951_;
  assign new_n3236_ = new_n843_ & new_n954_;
  assign new_n3237_ = ~new_n3235_ & ~new_n3236_;
  assign new_n3238_ = ~new_n3234_ & new_n3237_;
  assign new_n3239_ = new_n3233_ & new_n3238_;
  assign new_n3240_ = new_n3228_ & new_n3239_;
  assign new_n3241_ = new_n843_ & new_n961_;
  assign new_n3242_ = new_n843_ & new_n964_;
  assign new_n3243_ = new_n843_ & new_n967_;
  assign new_n3244_ = ~new_n3242_ & ~new_n3243_;
  assign new_n3245_ = ~new_n3241_ & new_n3244_;
  assign new_n3246_ = new_n843_ & new_n972_;
  assign new_n3247_ = new_n843_ & new_n975_;
  assign new_n3248_ = new_n843_ & new_n978_;
  assign new_n3249_ = ~new_n3247_ & ~new_n3248_;
  assign new_n3250_ = ~new_n3246_ & new_n3249_;
  assign new_n3251_ = new_n3245_ & new_n3250_;
  assign new_n3252_ = new_n843_ & new_n984_;
  assign new_n3253_ = new_n843_ & new_n987_;
  assign new_n3254_ = new_n843_ & new_n990_;
  assign new_n3255_ = ~new_n3253_ & ~new_n3254_;
  assign new_n3256_ = ~new_n3252_ & new_n3255_;
  assign new_n3257_ = new_n843_ & new_n994_;
  assign new_n3258_ = new_n843_ & new_n996_;
  assign new_n3259_ = ~new_n3257_ & ~new_n3258_;
  assign new_n3260_ = new_n3256_ & new_n3259_;
  assign new_n3261_ = new_n3251_ & new_n3260_;
  assign new_n3262_ = new_n3240_ & new_n3261_;
  assign new_n3263_ = new_n3217_ & new_n3262_;
  assign new_n3264_ = new_n3172_ & new_n3263_;
  assign new_n3265_ = new_n843_ & new_n1006_;
  assign new_n3266_ = new_n843_ & new_n1008_;
  assign new_n3267_ = new_n843_ & new_n1010_;
  assign new_n3268_ = ~new_n3266_ & ~new_n3267_;
  assign new_n3269_ = ~new_n3265_ & new_n3268_;
  assign new_n3270_ = new_n843_ & new_n1014_;
  assign new_n3271_ = new_n843_ & new_n1016_;
  assign new_n3272_ = new_n843_ & new_n1018_;
  assign new_n3273_ = ~new_n3271_ & ~new_n3272_;
  assign new_n3274_ = ~new_n3270_ & new_n3273_;
  assign new_n3275_ = new_n3269_ & new_n3274_;
  assign new_n3276_ = new_n843_ & new_n1023_;
  assign new_n3277_ = new_n843_ & new_n1025_;
  assign new_n3278_ = new_n843_ & new_n1027_;
  assign new_n3279_ = ~new_n3277_ & ~new_n3278_;
  assign new_n3280_ = ~new_n3276_ & new_n3279_;
  assign new_n3281_ = new_n843_ & new_n1031_;
  assign new_n3282_ = new_n843_ & new_n1033_;
  assign new_n3283_ = new_n843_ & new_n1035_;
  assign new_n3284_ = ~new_n3282_ & ~new_n3283_;
  assign new_n3285_ = ~new_n3281_ & new_n3284_;
  assign new_n3286_ = new_n3280_ & new_n3285_;
  assign new_n3287_ = new_n3275_ & new_n3286_;
  assign new_n3288_ = new_n843_ & new_n1041_;
  assign new_n3289_ = new_n843_ & new_n1043_;
  assign new_n3290_ = new_n843_ & new_n1045_;
  assign new_n3291_ = ~new_n3289_ & ~new_n3290_;
  assign new_n3292_ = ~new_n3288_ & new_n3291_;
  assign new_n3293_ = new_n843_ & new_n1049_;
  assign new_n3294_ = new_n843_ & new_n1051_;
  assign new_n3295_ = new_n843_ & new_n1053_;
  assign new_n3296_ = ~new_n3294_ & ~new_n3295_;
  assign new_n3297_ = ~new_n3293_ & new_n3296_;
  assign new_n3298_ = new_n3292_ & new_n3297_;
  assign new_n3299_ = new_n890_ & new_n1059_;
  assign new_n3300_ = new_n890_ & new_n1065_;
  assign new_n3301_ = new_n890_ & new_n1071_;
  assign new_n3302_ = ~new_n3300_ & ~new_n3301_;
  assign new_n3303_ = ~new_n3299_ & new_n3302_;
  assign new_n3304_ = new_n890_ & new_n1079_;
  assign new_n3305_ = new_n890_ & new_n1082_;
  assign new_n3306_ = ~new_n3304_ & ~new_n3305_;
  assign new_n3307_ = new_n3303_ & new_n3306_;
  assign new_n3308_ = new_n3298_ & new_n3307_;
  assign new_n3309_ = new_n3287_ & new_n3308_;
  assign new_n3310_ = new_n890_ & new_n1099_;
  assign new_n3311_ = new_n890_ & new_n1076_;
  assign new_n3312_ = new_n890_ & new_n1095_;
  assign new_n3313_ = ~new_n3311_ & ~new_n3312_;
  assign new_n3314_ = ~new_n3310_ & new_n3313_;
  assign new_n3315_ = new_n890_ & new_n1107_;
  assign new_n3316_ = new_n890_ & new_n1089_;
  assign new_n3317_ = new_n890_ & new_n1105_;
  assign new_n3318_ = ~new_n3316_ & ~new_n3317_;
  assign new_n3319_ = ~new_n3315_ & new_n3318_;
  assign new_n3320_ = new_n3314_ & new_n3319_;
  assign new_n3321_ = new_n890_ & new_n1120_;
  assign new_n3322_ = new_n890_ & new_n1103_;
  assign new_n3323_ = new_n890_ & new_n1118_;
  assign new_n3324_ = ~new_n3322_ & ~new_n3323_;
  assign new_n3325_ = ~new_n3321_ & new_n3324_;
  assign new_n3326_ = new_n890_ & new_n1135_;
  assign new_n3327_ = new_n890_ & new_n1114_;
  assign new_n3328_ = new_n890_ & new_n1131_;
  assign new_n3329_ = ~new_n3327_ & ~new_n3328_;
  assign new_n3330_ = ~new_n3326_ & new_n3329_;
  assign new_n3331_ = new_n3325_ & new_n3330_;
  assign new_n3332_ = new_n3320_ & new_n3331_;
  assign new_n3333_ = new_n890_ & new_n1149_;
  assign new_n3334_ = new_n890_ & new_n1127_;
  assign new_n3335_ = new_n890_ & new_n1145_;
  assign new_n3336_ = ~new_n3334_ & ~new_n3335_;
  assign new_n3337_ = ~new_n3333_ & new_n3336_;
  assign new_n3338_ = new_n890_ & new_n1157_;
  assign new_n3339_ = new_n890_ & new_n1141_;
  assign new_n3340_ = new_n890_ & new_n1155_;
  assign new_n3341_ = ~new_n3339_ & ~new_n3340_;
  assign new_n3342_ = ~new_n3338_ & new_n3341_;
  assign new_n3343_ = new_n3337_ & new_n3342_;
  assign new_n3344_ = new_n890_ & new_n1168_;
  assign new_n3345_ = new_n890_ & new_n1153_;
  assign new_n3346_ = new_n890_ & new_n1165_;
  assign new_n3347_ = ~new_n3345_ & ~new_n3346_;
  assign new_n3348_ = ~new_n3344_ & new_n3347_;
  assign new_n3349_ = new_n890_ & new_n1162_;
  assign new_n3350_ = new_n890_ & new_n1172_;
  assign new_n3351_ = ~new_n3349_ & ~new_n3350_;
  assign new_n3352_ = new_n3348_ & new_n3351_;
  assign new_n3353_ = new_n3343_ & new_n3352_;
  assign new_n3354_ = new_n3332_ & new_n3353_;
  assign new_n3355_ = new_n3309_ & new_n3354_;
  assign new_n3356_ = new_n890_ & new_n1186_;
  assign new_n3357_ = new_n890_ & new_n1174_;
  assign new_n3358_ = new_n890_ & new_n1184_;
  assign new_n3359_ = ~new_n3357_ & ~new_n3358_;
  assign new_n3360_ = ~new_n3356_ & new_n3359_;
  assign new_n3361_ = new_n890_ & new_n1194_;
  assign new_n3362_ = new_n890_ & new_n1182_;
  assign new_n3363_ = new_n890_ & new_n1192_;
  assign new_n3364_ = ~new_n3362_ & ~new_n3363_;
  assign new_n3365_ = ~new_n3361_ & new_n3364_;
  assign new_n3366_ = new_n3360_ & new_n3365_;
  assign new_n3367_ = new_n890_ & new_n1204_;
  assign new_n3368_ = new_n890_ & new_n1190_;
  assign new_n3369_ = new_n890_ & new_n1202_;
  assign new_n3370_ = ~new_n3368_ & ~new_n3369_;
  assign new_n3371_ = ~new_n3367_ & new_n3370_;
  assign new_n3372_ = new_n890_ & new_n1216_;
  assign new_n3373_ = new_n890_ & new_n1200_;
  assign new_n3374_ = new_n890_ & new_n1213_;
  assign new_n3375_ = ~new_n3373_ & ~new_n3374_;
  assign new_n3376_ = ~new_n3372_ & new_n3375_;
  assign new_n3377_ = new_n3371_ & new_n3376_;
  assign new_n3378_ = new_n3366_ & new_n3377_;
  assign new_n3379_ = new_n890_ & new_n1229_;
  assign new_n3380_ = new_n890_ & new_n1210_;
  assign new_n3381_ = new_n890_ & new_n1226_;
  assign new_n3382_ = ~new_n3380_ & ~new_n3381_;
  assign new_n3383_ = ~new_n3379_ & new_n3382_;
  assign new_n3384_ = new_n890_ & new_n1237_;
  assign new_n3385_ = new_n890_ & new_n1223_;
  assign new_n3386_ = new_n890_ & new_n1235_;
  assign new_n3387_ = ~new_n3385_ & ~new_n3386_;
  assign new_n3388_ = ~new_n3384_ & new_n3387_;
  assign new_n3389_ = new_n3383_ & new_n3388_;
  assign new_n3390_ = new_n909_ & new_n1830_;
  assign new_n3391_ = new_n890_ & new_n1233_;
  assign new_n3392_ = new_n890_ & new_n1243_;
  assign new_n3393_ = ~new_n3391_ & ~new_n3392_;
  assign new_n3394_ = ~new_n3390_ & new_n3393_;
  assign new_n3395_ = new_n909_ & new_n1833_;
  assign new_n3396_ = new_n909_ & new_n1827_;
  assign new_n3397_ = ~new_n3395_ & ~new_n3396_;
  assign new_n3398_ = new_n3394_ & new_n3397_;
  assign new_n3399_ = new_n3389_ & new_n3398_;
  assign new_n3400_ = new_n3378_ & new_n3399_;
  assign new_n3401_ = new_n909_ & new_n1838_;
  assign new_n3402_ = new_n909_ & new_n1840_;
  assign new_n3403_ = new_n909_ & new_n1842_;
  assign new_n3404_ = ~new_n3402_ & ~new_n3403_;
  assign new_n3405_ = ~new_n3401_ & new_n3404_;
  assign new_n3406_ = new_n909_ & new_n1857_;
  assign new_n3407_ = new_n909_ & new_n1847_;
  assign new_n3408_ = new_n909_ & new_n1849_;
  assign new_n3409_ = ~new_n3407_ & ~new_n3408_;
  assign new_n3410_ = ~new_n3406_ & new_n3409_;
  assign new_n3411_ = new_n3405_ & new_n3410_;
  assign new_n3412_ = new_n909_ & new_n1866_;
  assign new_n3413_ = new_n909_ & new_n1859_;
  assign new_n3414_ = new_n909_ & new_n1855_;
  assign new_n3415_ = ~new_n3413_ & ~new_n3414_;
  assign new_n3416_ = ~new_n3412_ & new_n3415_;
  assign new_n3417_ = new_n909_ & new_n1878_;
  assign new_n3418_ = new_n909_ & new_n1868_;
  assign new_n3419_ = new_n909_ & new_n1864_;
  assign new_n3420_ = ~new_n3418_ & ~new_n3419_;
  assign new_n3421_ = ~new_n3417_ & new_n3420_;
  assign new_n3422_ = new_n3416_ & new_n3421_;
  assign new_n3423_ = new_n3411_ & new_n3422_;
  assign new_n3424_ = new_n909_ & new_n1889_;
  assign new_n3425_ = new_n909_ & new_n1881_;
  assign new_n3426_ = new_n909_ & new_n1875_;
  assign new_n3427_ = ~new_n3425_ & ~new_n3426_;
  assign new_n3428_ = ~new_n3424_ & new_n3427_;
  assign new_n3429_ = new_n909_ & new_n1900_;
  assign new_n3430_ = new_n909_ & new_n1892_;
  assign new_n3431_ = new_n909_ & new_n1886_;
  assign new_n3432_ = ~new_n3430_ & ~new_n3431_;
  assign new_n3433_ = ~new_n3429_ & new_n3432_;
  assign new_n3434_ = new_n3428_ & new_n3433_;
  assign new_n3435_ = new_n909_ & new_n1913_;
  assign new_n3436_ = new_n909_ & new_n1902_;
  assign new_n3437_ = new_n909_ & new_n1898_;
  assign new_n3438_ = ~new_n3436_ & ~new_n3437_;
  assign new_n3439_ = ~new_n3435_ & new_n3438_;
  assign new_n3440_ = new_n908_ & new_n1975_;
  assign new_n3441_ = new_n1735_ & new_n3440_;
  assign new_n3442_ = new_n1738_ & new_n3440_;
  assign new_n3443_ = ~new_n3441_ & ~new_n3442_;
  assign new_n3444_ = new_n3439_ & new_n3443_;
  assign new_n3445_ = new_n3434_ & new_n3444_;
  assign new_n3446_ = new_n3423_ & new_n3445_;
  assign new_n3447_ = new_n3400_ & new_n3446_;
  assign new_n3448_ = new_n3355_ & new_n3447_;
  assign new_n3449_ = new_n3264_ & new_n3448_;
  assign new_n3450_ = new_n3081_ & new_n3449_;
  assign new_n3451_ = new_n2704_ & new_n3450_;
  assign new_n3452_ = new_n1934_ & new_n3451_;
  assign new_n3453_ = new_n908_ & new_n1986_;
  assign new_n3454_ = new_n1735_ & new_n3453_;
  assign new_n3455_ = new_n1725_ & new_n3440_;
  assign new_n3456_ = new_n1749_ & new_n3440_;
  assign new_n3457_ = ~new_n3455_ & ~new_n3456_;
  assign new_n3458_ = ~new_n3454_ & new_n3457_;
  assign new_n3459_ = new_n1749_ & new_n3453_;
  assign new_n3460_ = new_n1738_ & new_n3453_;
  assign new_n3461_ = new_n1725_ & new_n3453_;
  assign new_n3462_ = ~new_n3460_ & ~new_n3461_;
  assign new_n3463_ = ~new_n3459_ & new_n3462_;
  assign new_n3464_ = new_n3458_ & new_n3463_;
  assign new_n3465_ = new_n916_ & new_n1827_;
  assign new_n3466_ = new_n916_ & new_n1830_;
  assign new_n3467_ = new_n916_ & new_n1833_;
  assign new_n3468_ = ~new_n3466_ & ~new_n3467_;
  assign new_n3469_ = ~new_n3465_ & new_n3468_;
  assign new_n3470_ = new_n916_ & new_n1838_;
  assign new_n3471_ = new_n916_ & new_n1840_;
  assign new_n3472_ = new_n916_ & new_n1842_;
  assign new_n3473_ = ~new_n3471_ & ~new_n3472_;
  assign new_n3474_ = ~new_n3470_ & new_n3473_;
  assign new_n3475_ = new_n3469_ & new_n3474_;
  assign new_n3476_ = new_n3464_ & new_n3475_;
  assign new_n3477_ = new_n916_ & new_n1857_;
  assign new_n3478_ = new_n916_ & new_n1847_;
  assign new_n3479_ = new_n916_ & new_n1849_;
  assign new_n3480_ = ~new_n3478_ & ~new_n3479_;
  assign new_n3481_ = ~new_n3477_ & new_n3480_;
  assign new_n3482_ = new_n916_ & new_n1866_;
  assign new_n3483_ = new_n916_ & new_n1859_;
  assign new_n3484_ = new_n916_ & new_n1855_;
  assign new_n3485_ = ~new_n3483_ & ~new_n3484_;
  assign new_n3486_ = ~new_n3482_ & new_n3485_;
  assign new_n3487_ = new_n3481_ & new_n3486_;
  assign new_n3488_ = new_n916_ & new_n1878_;
  assign new_n3489_ = new_n916_ & new_n1868_;
  assign new_n3490_ = new_n916_ & new_n1864_;
  assign new_n3491_ = ~new_n3489_ & ~new_n3490_;
  assign new_n3492_ = ~new_n3488_ & new_n3491_;
  assign new_n3493_ = new_n916_ & new_n1889_;
  assign new_n3494_ = new_n916_ & new_n1881_;
  assign new_n3495_ = new_n916_ & new_n1875_;
  assign new_n3496_ = ~new_n3494_ & ~new_n3495_;
  assign new_n3497_ = ~new_n3493_ & new_n3496_;
  assign new_n3498_ = new_n3492_ & new_n3497_;
  assign new_n3499_ = new_n3487_ & new_n3498_;
  assign new_n3500_ = new_n3476_ & new_n3499_;
  assign new_n3501_ = new_n916_ & new_n1900_;
  assign new_n3502_ = new_n916_ & new_n1892_;
  assign new_n3503_ = new_n916_ & new_n1886_;
  assign new_n3504_ = ~new_n3502_ & ~new_n3503_;
  assign new_n3505_ = ~new_n3501_ & new_n3504_;
  assign new_n3506_ = new_n916_ & new_n1913_;
  assign new_n3507_ = new_n916_ & new_n1902_;
  assign new_n3508_ = new_n916_ & new_n1898_;
  assign new_n3509_ = ~new_n3507_ & ~new_n3508_;
  assign new_n3510_ = ~new_n3506_ & new_n3509_;
  assign new_n3511_ = new_n3505_ & new_n3510_;
  assign new_n3512_ = new_n908_ & new_n2045_;
  assign new_n3513_ = new_n1725_ & new_n3512_;
  assign new_n3514_ = new_n1735_ & new_n3512_;
  assign new_n3515_ = new_n1738_ & new_n3512_;
  assign new_n3516_ = ~new_n3514_ & ~new_n3515_;
  assign new_n3517_ = ~new_n3513_ & new_n3516_;
  assign new_n3518_ = new_n908_ & new_n2052_;
  assign new_n3519_ = new_n1738_ & new_n3518_;
  assign new_n3520_ = new_n1749_ & new_n3512_;
  assign new_n3521_ = new_n1735_ & new_n3518_;
  assign new_n3522_ = ~new_n3520_ & ~new_n3521_;
  assign new_n3523_ = ~new_n3519_ & new_n3522_;
  assign new_n3524_ = new_n3517_ & new_n3523_;
  assign new_n3525_ = new_n3511_ & new_n3524_;
  assign new_n3526_ = new_n929_ & new_n1830_;
  assign new_n3527_ = new_n1725_ & new_n3518_;
  assign new_n3528_ = new_n1749_ & new_n3518_;
  assign new_n3529_ = ~new_n3527_ & ~new_n3528_;
  assign new_n3530_ = ~new_n3526_ & new_n3529_;
  assign new_n3531_ = new_n929_ & new_n1840_;
  assign new_n3532_ = new_n929_ & new_n1833_;
  assign new_n3533_ = new_n929_ & new_n1827_;
  assign new_n3534_ = ~new_n3532_ & ~new_n3533_;
  assign new_n3535_ = ~new_n3531_ & new_n3534_;
  assign new_n3536_ = new_n3530_ & new_n3535_;
  assign new_n3537_ = new_n929_ & new_n1847_;
  assign new_n3538_ = new_n929_ & new_n1842_;
  assign new_n3539_ = new_n929_ & new_n1838_;
  assign new_n3540_ = ~new_n3538_ & ~new_n3539_;
  assign new_n3541_ = ~new_n3537_ & new_n3540_;
  assign new_n3542_ = new_n929_ & new_n1849_;
  assign new_n3543_ = new_n929_ & new_n1857_;
  assign new_n3544_ = ~new_n3542_ & ~new_n3543_;
  assign new_n3545_ = new_n3541_ & new_n3544_;
  assign new_n3546_ = new_n3536_ & new_n3545_;
  assign new_n3547_ = new_n3525_ & new_n3546_;
  assign new_n3548_ = new_n3500_ & new_n3547_;
  assign new_n3549_ = new_n929_ & new_n1866_;
  assign new_n3550_ = new_n929_ & new_n1859_;
  assign new_n3551_ = new_n929_ & new_n1855_;
  assign new_n3552_ = ~new_n3550_ & ~new_n3551_;
  assign new_n3553_ = ~new_n3549_ & new_n3552_;
  assign new_n3554_ = new_n929_ & new_n1878_;
  assign new_n3555_ = new_n929_ & new_n1868_;
  assign new_n3556_ = new_n929_ & new_n1864_;
  assign new_n3557_ = ~new_n3555_ & ~new_n3556_;
  assign new_n3558_ = ~new_n3554_ & new_n3557_;
  assign new_n3559_ = new_n3553_ & new_n3558_;
  assign new_n3560_ = new_n929_ & new_n1889_;
  assign new_n3561_ = new_n929_ & new_n1881_;
  assign new_n3562_ = new_n929_ & new_n1875_;
  assign new_n3563_ = ~new_n3561_ & ~new_n3562_;
  assign new_n3564_ = ~new_n3560_ & new_n3563_;
  assign new_n3565_ = new_n929_ & new_n1900_;
  assign new_n3566_ = new_n929_ & new_n1892_;
  assign new_n3567_ = new_n929_ & new_n1886_;
  assign new_n3568_ = ~new_n3566_ & ~new_n3567_;
  assign new_n3569_ = ~new_n3565_ & new_n3568_;
  assign new_n3570_ = new_n3564_ & new_n3569_;
  assign new_n3571_ = new_n3559_ & new_n3570_;
  assign new_n3572_ = new_n929_ & new_n1913_;
  assign new_n3573_ = new_n929_ & new_n1902_;
  assign new_n3574_ = new_n929_ & new_n1898_;
  assign new_n3575_ = ~new_n3573_ & ~new_n3574_;
  assign new_n3576_ = ~new_n3572_ & new_n3575_;
  assign new_n3577_ = new_n928_ & new_n1975_;
  assign new_n3578_ = new_n1725_ & new_n3577_;
  assign new_n3579_ = new_n1735_ & new_n3577_;
  assign new_n3580_ = new_n1738_ & new_n3577_;
  assign new_n3581_ = ~new_n3579_ & ~new_n3580_;
  assign new_n3582_ = ~new_n3578_ & new_n3581_;
  assign new_n3583_ = new_n3576_ & new_n3582_;
  assign new_n3584_ = new_n928_ & new_n1986_;
  assign new_n3585_ = new_n1738_ & new_n3584_;
  assign new_n3586_ = new_n1749_ & new_n3577_;
  assign new_n3587_ = new_n1735_ & new_n3584_;
  assign new_n3588_ = ~new_n3586_ & ~new_n3587_;
  assign new_n3589_ = ~new_n3585_ & new_n3588_;
  assign new_n3590_ = new_n1725_ & new_n3584_;
  assign new_n3591_ = new_n1749_ & new_n3584_;
  assign new_n3592_ = ~new_n3590_ & ~new_n3591_;
  assign new_n3593_ = new_n3589_ & new_n3592_;
  assign new_n3594_ = new_n3583_ & new_n3593_;
  assign new_n3595_ = new_n3571_ & new_n3594_;
  assign new_n3596_ = new_n935_ & new_n1827_;
  assign new_n3597_ = new_n935_ & new_n1830_;
  assign new_n3598_ = new_n935_ & new_n1833_;
  assign new_n3599_ = ~new_n3597_ & ~new_n3598_;
  assign new_n3600_ = ~new_n3596_ & new_n3599_;
  assign new_n3601_ = new_n935_ & new_n1838_;
  assign new_n3602_ = new_n935_ & new_n1840_;
  assign new_n3603_ = new_n935_ & new_n1842_;
  assign new_n3604_ = ~new_n3602_ & ~new_n3603_;
  assign new_n3605_ = ~new_n3601_ & new_n3604_;
  assign new_n3606_ = new_n3600_ & new_n3605_;
  assign new_n3607_ = new_n935_ & new_n1857_;
  assign new_n3608_ = new_n935_ & new_n1847_;
  assign new_n3609_ = new_n935_ & new_n1849_;
  assign new_n3610_ = ~new_n3608_ & ~new_n3609_;
  assign new_n3611_ = ~new_n3607_ & new_n3610_;
  assign new_n3612_ = new_n935_ & new_n1866_;
  assign new_n3613_ = new_n935_ & new_n1859_;
  assign new_n3614_ = new_n935_ & new_n1855_;
  assign new_n3615_ = ~new_n3613_ & ~new_n3614_;
  assign new_n3616_ = ~new_n3612_ & new_n3615_;
  assign new_n3617_ = new_n3611_ & new_n3616_;
  assign new_n3618_ = new_n3606_ & new_n3617_;
  assign new_n3619_ = new_n935_ & new_n1878_;
  assign new_n3620_ = new_n935_ & new_n1868_;
  assign new_n3621_ = new_n935_ & new_n1864_;
  assign new_n3622_ = ~new_n3620_ & ~new_n3621_;
  assign new_n3623_ = ~new_n3619_ & new_n3622_;
  assign new_n3624_ = new_n935_ & new_n1889_;
  assign new_n3625_ = new_n935_ & new_n1881_;
  assign new_n3626_ = new_n935_ & new_n1875_;
  assign new_n3627_ = ~new_n3625_ & ~new_n3626_;
  assign new_n3628_ = ~new_n3624_ & new_n3627_;
  assign new_n3629_ = new_n3623_ & new_n3628_;
  assign new_n3630_ = new_n935_ & new_n1900_;
  assign new_n3631_ = new_n935_ & new_n1892_;
  assign new_n3632_ = new_n935_ & new_n1886_;
  assign new_n3633_ = ~new_n3631_ & ~new_n3632_;
  assign new_n3634_ = ~new_n3630_ & new_n3633_;
  assign new_n3635_ = new_n935_ & new_n1902_;
  assign new_n3636_ = new_n935_ & new_n1898_;
  assign new_n3637_ = ~new_n3635_ & ~new_n3636_;
  assign new_n3638_ = new_n3634_ & new_n3637_;
  assign new_n3639_ = new_n3629_ & new_n3638_;
  assign new_n3640_ = new_n3618_ & new_n3639_;
  assign new_n3641_ = new_n3595_ & new_n3640_;
  assign new_n3642_ = new_n3548_ & new_n3641_;
  assign new_n3643_ = new_n928_ & new_n2045_;
  assign new_n3644_ = new_n1738_ & new_n3643_;
  assign new_n3645_ = new_n935_ & new_n1913_;
  assign new_n3646_ = new_n1735_ & new_n3643_;
  assign new_n3647_ = ~new_n3645_ & ~new_n3646_;
  assign new_n3648_ = ~new_n3644_ & new_n3647_;
  assign new_n3649_ = new_n928_ & new_n2052_;
  assign new_n3650_ = new_n1735_ & new_n3649_;
  assign new_n3651_ = new_n1725_ & new_n3643_;
  assign new_n3652_ = new_n1749_ & new_n3643_;
  assign new_n3653_ = ~new_n3651_ & ~new_n3652_;
  assign new_n3654_ = ~new_n3650_ & new_n3653_;
  assign new_n3655_ = new_n3648_ & new_n3654_;
  assign new_n3656_ = new_n1749_ & new_n3649_;
  assign new_n3657_ = new_n1738_ & new_n3649_;
  assign new_n3658_ = new_n1725_ & new_n3649_;
  assign new_n3659_ = ~new_n3657_ & ~new_n3658_;
  assign new_n3660_ = ~new_n3656_ & new_n3659_;
  assign new_n3661_ = new_n139_ & new_n1974_;
  assign new_n3662_ = new_n947_ & new_n3661_;
  assign new_n3663_ = new_n516_ & new_n518_;
  assign new_n3664_ = ~A168 & ~A169;
  assign new_n3665_ = ~A170 & new_n3664_;
  assign new_n3666_ = new_n3663_ & new_n3665_;
  assign new_n3667_ = new_n3662_ & new_n3666_;
  assign new_n3668_ = new_n950_ & new_n3661_;
  assign new_n3669_ = new_n3666_ & new_n3668_;
  assign new_n3670_ = new_n953_ & new_n3661_;
  assign new_n3671_ = new_n3666_ & new_n3670_;
  assign new_n3672_ = ~new_n3669_ & ~new_n3671_;
  assign new_n3673_ = ~new_n3667_ & new_n3672_;
  assign new_n3674_ = new_n3660_ & new_n3673_;
  assign new_n3675_ = new_n3655_ & new_n3674_;
  assign new_n3676_ = new_n155_ & new_n1974_;
  assign new_n3677_ = new_n960_ & new_n3676_;
  assign new_n3678_ = new_n3666_ & new_n3677_;
  assign new_n3679_ = new_n963_ & new_n3661_;
  assign new_n3680_ = new_n3666_ & new_n3679_;
  assign new_n3681_ = new_n966_ & new_n3676_;
  assign new_n3682_ = new_n3666_ & new_n3681_;
  assign new_n3683_ = ~new_n3680_ & ~new_n3682_;
  assign new_n3684_ = ~new_n3678_ & new_n3683_;
  assign new_n3685_ = new_n971_ & new_n3676_;
  assign new_n3686_ = new_n3666_ & new_n3685_;
  assign new_n3687_ = new_n974_ & new_n3676_;
  assign new_n3688_ = new_n3666_ & new_n3687_;
  assign new_n3689_ = new_n977_ & new_n3676_;
  assign new_n3690_ = new_n3666_ & new_n3689_;
  assign new_n3691_ = ~new_n3688_ & ~new_n3690_;
  assign new_n3692_ = ~new_n3686_ & new_n3691_;
  assign new_n3693_ = new_n3684_ & new_n3692_;
  assign new_n3694_ = new_n983_ & new_n3676_;
  assign new_n3695_ = new_n3666_ & new_n3694_;
  assign new_n3696_ = new_n986_ & new_n3676_;
  assign new_n3697_ = new_n3666_ & new_n3696_;
  assign new_n3698_ = new_n989_ & new_n3676_;
  assign new_n3699_ = new_n3666_ & new_n3698_;
  assign new_n3700_ = ~new_n3697_ & ~new_n3699_;
  assign new_n3701_ = ~new_n3695_ & new_n3700_;
  assign new_n3702_ = new_n186_ & new_n1974_;
  assign new_n3703_ = new_n966_ & new_n3702_;
  assign new_n3704_ = new_n3666_ & new_n3703_;
  assign new_n3705_ = new_n960_ & new_n3702_;
  assign new_n3706_ = new_n3666_ & new_n3705_;
  assign new_n3707_ = ~new_n3704_ & ~new_n3706_;
  assign new_n3708_ = new_n3701_ & new_n3707_;
  assign new_n3709_ = new_n3693_ & new_n3708_;
  assign new_n3710_ = new_n3675_ & new_n3709_;
  assign new_n3711_ = new_n971_ & new_n3702_;
  assign new_n3712_ = new_n3666_ & new_n3711_;
  assign new_n3713_ = new_n974_ & new_n3702_;
  assign new_n3714_ = new_n3666_ & new_n3713_;
  assign new_n3715_ = new_n977_ & new_n3702_;
  assign new_n3716_ = new_n3666_ & new_n3715_;
  assign new_n3717_ = ~new_n3714_ & ~new_n3716_;
  assign new_n3718_ = ~new_n3712_ & new_n3717_;
  assign new_n3719_ = new_n983_ & new_n3702_;
  assign new_n3720_ = new_n3666_ & new_n3719_;
  assign new_n3721_ = new_n986_ & new_n3702_;
  assign new_n3722_ = new_n3666_ & new_n3721_;
  assign new_n3723_ = new_n989_ & new_n3702_;
  assign new_n3724_ = new_n3666_ & new_n3723_;
  assign new_n3725_ = ~new_n3722_ & ~new_n3724_;
  assign new_n3726_ = ~new_n3720_ & new_n3725_;
  assign new_n3727_ = new_n3718_ & new_n3726_;
  assign new_n3728_ = new_n209_ & new_n1974_;
  assign new_n3729_ = new_n947_ & new_n3728_;
  assign new_n3730_ = new_n3666_ & new_n3729_;
  assign new_n3731_ = new_n950_ & new_n3728_;
  assign new_n3732_ = new_n3666_ & new_n3731_;
  assign new_n3733_ = new_n953_ & new_n3728_;
  assign new_n3734_ = new_n3666_ & new_n3733_;
  assign new_n3735_ = ~new_n3732_ & ~new_n3734_;
  assign new_n3736_ = ~new_n3730_ & new_n3735_;
  assign new_n3737_ = new_n218_ & new_n1974_;
  assign new_n3738_ = new_n953_ & new_n3737_;
  assign new_n3739_ = new_n3666_ & new_n3738_;
  assign new_n3740_ = new_n963_ & new_n3728_;
  assign new_n3741_ = new_n3666_ & new_n3740_;
  assign new_n3742_ = new_n950_ & new_n3737_;
  assign new_n3743_ = new_n3666_ & new_n3742_;
  assign new_n3744_ = ~new_n3741_ & ~new_n3743_;
  assign new_n3745_ = ~new_n3739_ & new_n3744_;
  assign new_n3746_ = new_n3736_ & new_n3745_;
  assign new_n3747_ = new_n3727_ & new_n3746_;
  assign new_n3748_ = new_n236_ & new_n1974_;
  assign new_n3749_ = new_n950_ & new_n3748_;
  assign new_n3750_ = new_n3666_ & new_n3749_;
  assign new_n3751_ = new_n947_ & new_n3737_;
  assign new_n3752_ = new_n3666_ & new_n3751_;
  assign new_n3753_ = new_n963_ & new_n3737_;
  assign new_n3754_ = new_n3666_ & new_n3753_;
  assign new_n3755_ = ~new_n3752_ & ~new_n3754_;
  assign new_n3756_ = ~new_n3750_ & new_n3755_;
  assign new_n3757_ = new_n963_ & new_n3748_;
  assign new_n3758_ = new_n3666_ & new_n3757_;
  assign new_n3759_ = new_n953_ & new_n3748_;
  assign new_n3760_ = new_n3666_ & new_n3759_;
  assign new_n3761_ = new_n947_ & new_n3748_;
  assign new_n3762_ = new_n3666_ & new_n3761_;
  assign new_n3763_ = ~new_n3760_ & ~new_n3762_;
  assign new_n3764_ = ~new_n3758_ & new_n3763_;
  assign new_n3765_ = new_n3756_ & new_n3764_;
  assign new_n3766_ = new_n139_ & new_n1985_;
  assign new_n3767_ = new_n947_ & new_n3766_;
  assign new_n3768_ = new_n3666_ & new_n3767_;
  assign new_n3769_ = new_n950_ & new_n3766_;
  assign new_n3770_ = new_n3666_ & new_n3769_;
  assign new_n3771_ = new_n953_ & new_n3766_;
  assign new_n3772_ = new_n3666_ & new_n3771_;
  assign new_n3773_ = ~new_n3770_ & ~new_n3772_;
  assign new_n3774_ = ~new_n3768_ & new_n3773_;
  assign new_n3775_ = new_n963_ & new_n3766_;
  assign new_n3776_ = new_n3666_ & new_n3775_;
  assign new_n3777_ = new_n155_ & new_n1985_;
  assign new_n3778_ = new_n966_ & new_n3777_;
  assign new_n3779_ = new_n3666_ & new_n3778_;
  assign new_n3780_ = ~new_n3776_ & ~new_n3779_;
  assign new_n3781_ = new_n3774_ & new_n3780_;
  assign new_n3782_ = new_n3765_ & new_n3781_;
  assign new_n3783_ = new_n3747_ & new_n3782_;
  assign new_n3784_ = new_n3710_ & new_n3783_;
  assign new_n3785_ = new_n977_ & new_n3777_;
  assign new_n3786_ = new_n3666_ & new_n3785_;
  assign new_n3787_ = new_n960_ & new_n3777_;
  assign new_n3788_ = new_n3666_ & new_n3787_;
  assign new_n3789_ = new_n974_ & new_n3777_;
  assign new_n3790_ = new_n3666_ & new_n3789_;
  assign new_n3791_ = ~new_n3788_ & ~new_n3790_;
  assign new_n3792_ = ~new_n3786_ & new_n3791_;
  assign new_n3793_ = new_n989_ & new_n3777_;
  assign new_n3794_ = new_n3666_ & new_n3793_;
  assign new_n3795_ = new_n971_ & new_n3777_;
  assign new_n3796_ = new_n3666_ & new_n3795_;
  assign new_n3797_ = new_n986_ & new_n3777_;
  assign new_n3798_ = new_n3666_ & new_n3797_;
  assign new_n3799_ = ~new_n3796_ & ~new_n3798_;
  assign new_n3800_ = ~new_n3794_ & new_n3799_;
  assign new_n3801_ = new_n3792_ & new_n3800_;
  assign new_n3802_ = new_n186_ & new_n1985_;
  assign new_n3803_ = new_n960_ & new_n3802_;
  assign new_n3804_ = new_n3666_ & new_n3803_;
  assign new_n3805_ = new_n983_ & new_n3777_;
  assign new_n3806_ = new_n3666_ & new_n3805_;
  assign new_n3807_ = new_n966_ & new_n3802_;
  assign new_n3808_ = new_n3666_ & new_n3807_;
  assign new_n3809_ = ~new_n3806_ & ~new_n3808_;
  assign new_n3810_ = ~new_n3804_ & new_n3809_;
  assign new_n3811_ = new_n971_ & new_n3802_;
  assign new_n3812_ = new_n3666_ & new_n3811_;
  assign new_n3813_ = new_n974_ & new_n3802_;
  assign new_n3814_ = new_n3666_ & new_n3813_;
  assign new_n3815_ = new_n977_ & new_n3802_;
  assign new_n3816_ = new_n3666_ & new_n3815_;
  assign new_n3817_ = ~new_n3814_ & ~new_n3816_;
  assign new_n3818_ = ~new_n3812_ & new_n3817_;
  assign new_n3819_ = new_n3810_ & new_n3818_;
  assign new_n3820_ = new_n3801_ & new_n3819_;
  assign new_n3821_ = new_n983_ & new_n3802_;
  assign new_n3822_ = new_n3666_ & new_n3821_;
  assign new_n3823_ = new_n986_ & new_n3802_;
  assign new_n3824_ = new_n3666_ & new_n3823_;
  assign new_n3825_ = new_n989_ & new_n3802_;
  assign new_n3826_ = new_n3666_ & new_n3825_;
  assign new_n3827_ = ~new_n3824_ & ~new_n3826_;
  assign new_n3828_ = ~new_n3822_ & new_n3827_;
  assign new_n3829_ = new_n209_ & new_n1985_;
  assign new_n3830_ = new_n947_ & new_n3829_;
  assign new_n3831_ = new_n3666_ & new_n3830_;
  assign new_n3832_ = new_n950_ & new_n3829_;
  assign new_n3833_ = new_n3666_ & new_n3832_;
  assign new_n3834_ = new_n953_ & new_n3829_;
  assign new_n3835_ = new_n3666_ & new_n3834_;
  assign new_n3836_ = ~new_n3833_ & ~new_n3835_;
  assign new_n3837_ = ~new_n3831_ & new_n3836_;
  assign new_n3838_ = new_n3828_ & new_n3837_;
  assign new_n3839_ = new_n218_ & new_n1985_;
  assign new_n3840_ = new_n953_ & new_n3839_;
  assign new_n3841_ = new_n3666_ & new_n3840_;
  assign new_n3842_ = new_n963_ & new_n3829_;
  assign new_n3843_ = new_n3666_ & new_n3842_;
  assign new_n3844_ = new_n950_ & new_n3839_;
  assign new_n3845_ = new_n3666_ & new_n3844_;
  assign new_n3846_ = ~new_n3843_ & ~new_n3845_;
  assign new_n3847_ = ~new_n3841_ & new_n3846_;
  assign new_n3848_ = new_n947_ & new_n3839_;
  assign new_n3849_ = new_n3666_ & new_n3848_;
  assign new_n3850_ = new_n963_ & new_n3839_;
  assign new_n3851_ = new_n3666_ & new_n3850_;
  assign new_n3852_ = ~new_n3849_ & ~new_n3851_;
  assign new_n3853_ = new_n3847_ & new_n3852_;
  assign new_n3854_ = new_n3838_ & new_n3853_;
  assign new_n3855_ = new_n3820_ & new_n3854_;
  assign new_n3856_ = new_n236_ & new_n1985_;
  assign new_n3857_ = new_n947_ & new_n3856_;
  assign new_n3858_ = new_n3666_ & new_n3857_;
  assign new_n3859_ = new_n950_ & new_n3856_;
  assign new_n3860_ = new_n3666_ & new_n3859_;
  assign new_n3861_ = new_n953_ & new_n3856_;
  assign new_n3862_ = new_n3666_ & new_n3861_;
  assign new_n3863_ = ~new_n3860_ & ~new_n3862_;
  assign new_n3864_ = ~new_n3858_ & new_n3863_;
  assign new_n3865_ = new_n518_ & new_n533_;
  assign new_n3866_ = new_n3665_ & new_n3865_;
  assign new_n3867_ = new_n3670_ & new_n3866_;
  assign new_n3868_ = new_n963_ & new_n3856_;
  assign new_n3869_ = new_n3666_ & new_n3868_;
  assign new_n3870_ = new_n3668_ & new_n3866_;
  assign new_n3871_ = ~new_n3869_ & ~new_n3870_;
  assign new_n3872_ = ~new_n3867_ & new_n3871_;
  assign new_n3873_ = new_n3864_ & new_n3872_;
  assign new_n3874_ = new_n3681_ & new_n3866_;
  assign new_n3875_ = new_n3662_ & new_n3866_;
  assign new_n3876_ = new_n3679_ & new_n3866_;
  assign new_n3877_ = ~new_n3875_ & ~new_n3876_;
  assign new_n3878_ = ~new_n3874_ & new_n3877_;
  assign new_n3879_ = new_n3689_ & new_n3866_;
  assign new_n3880_ = new_n3677_ & new_n3866_;
  assign new_n3881_ = new_n3687_ & new_n3866_;
  assign new_n3882_ = ~new_n3880_ & ~new_n3881_;
  assign new_n3883_ = ~new_n3879_ & new_n3882_;
  assign new_n3884_ = new_n3878_ & new_n3883_;
  assign new_n3885_ = new_n3873_ & new_n3884_;
  assign new_n3886_ = new_n3698_ & new_n3866_;
  assign new_n3887_ = new_n3685_ & new_n3866_;
  assign new_n3888_ = new_n3696_ & new_n3866_;
  assign new_n3889_ = ~new_n3887_ & ~new_n3888_;
  assign new_n3890_ = ~new_n3886_ & new_n3889_;
  assign new_n3891_ = new_n3705_ & new_n3866_;
  assign new_n3892_ = new_n3694_ & new_n3866_;
  assign new_n3893_ = new_n3703_ & new_n3866_;
  assign new_n3894_ = ~new_n3892_ & ~new_n3893_;
  assign new_n3895_ = ~new_n3891_ & new_n3894_;
  assign new_n3896_ = new_n3890_ & new_n3895_;
  assign new_n3897_ = new_n3711_ & new_n3866_;
  assign new_n3898_ = new_n3713_ & new_n3866_;
  assign new_n3899_ = new_n3715_ & new_n3866_;
  assign new_n3900_ = ~new_n3898_ & ~new_n3899_;
  assign new_n3901_ = ~new_n3897_ & new_n3900_;
  assign new_n3902_ = new_n3721_ & new_n3866_;
  assign new_n3903_ = new_n3723_ & new_n3866_;
  assign new_n3904_ = ~new_n3902_ & ~new_n3903_;
  assign new_n3905_ = new_n3901_ & new_n3904_;
  assign new_n3906_ = new_n3896_ & new_n3905_;
  assign new_n3907_ = new_n3885_ & new_n3906_;
  assign new_n3908_ = new_n3855_ & new_n3907_;
  assign new_n3909_ = new_n3784_ & new_n3908_;
  assign new_n3910_ = new_n3642_ & new_n3909_;
  assign new_n3911_ = new_n3733_ & new_n3866_;
  assign new_n3912_ = new_n3719_ & new_n3866_;
  assign new_n3913_ = new_n3731_ & new_n3866_;
  assign new_n3914_ = ~new_n3912_ & ~new_n3913_;
  assign new_n3915_ = ~new_n3911_ & new_n3914_;
  assign new_n3916_ = new_n3742_ & new_n3866_;
  assign new_n3917_ = new_n3729_ & new_n3866_;
  assign new_n3918_ = new_n3740_ & new_n3866_;
  assign new_n3919_ = ~new_n3917_ & ~new_n3918_;
  assign new_n3920_ = ~new_n3916_ & new_n3919_;
  assign new_n3921_ = new_n3915_ & new_n3920_;
  assign new_n3922_ = new_n3753_ & new_n3866_;
  assign new_n3923_ = new_n3738_ & new_n3866_;
  assign new_n3924_ = new_n3751_ & new_n3866_;
  assign new_n3925_ = ~new_n3923_ & ~new_n3924_;
  assign new_n3926_ = ~new_n3922_ & new_n3925_;
  assign new_n3927_ = new_n3761_ & new_n3866_;
  assign new_n3928_ = new_n3749_ & new_n3866_;
  assign new_n3929_ = new_n3759_ & new_n3866_;
  assign new_n3930_ = ~new_n3928_ & ~new_n3929_;
  assign new_n3931_ = ~new_n3927_ & new_n3930_;
  assign new_n3932_ = new_n3926_ & new_n3931_;
  assign new_n3933_ = new_n3921_ & new_n3932_;
  assign new_n3934_ = new_n3771_ & new_n3866_;
  assign new_n3935_ = new_n3757_ & new_n3866_;
  assign new_n3936_ = new_n3769_ & new_n3866_;
  assign new_n3937_ = ~new_n3935_ & ~new_n3936_;
  assign new_n3938_ = ~new_n3934_ & new_n3937_;
  assign new_n3939_ = new_n3778_ & new_n3866_;
  assign new_n3940_ = new_n3767_ & new_n3866_;
  assign new_n3941_ = new_n3775_ & new_n3866_;
  assign new_n3942_ = ~new_n3940_ & ~new_n3941_;
  assign new_n3943_ = ~new_n3939_ & new_n3942_;
  assign new_n3944_ = new_n3938_ & new_n3943_;
  assign new_n3945_ = new_n3785_ & new_n3866_;
  assign new_n3946_ = new_n3787_ & new_n3866_;
  assign new_n3947_ = new_n3789_ & new_n3866_;
  assign new_n3948_ = ~new_n3946_ & ~new_n3947_;
  assign new_n3949_ = ~new_n3945_ & new_n3948_;
  assign new_n3950_ = new_n3793_ & new_n3866_;
  assign new_n3951_ = new_n3795_ & new_n3866_;
  assign new_n3952_ = new_n3797_ & new_n3866_;
  assign new_n3953_ = ~new_n3951_ & ~new_n3952_;
  assign new_n3954_ = ~new_n3950_ & new_n3953_;
  assign new_n3955_ = new_n3949_ & new_n3954_;
  assign new_n3956_ = new_n3944_ & new_n3955_;
  assign new_n3957_ = new_n3933_ & new_n3956_;
  assign new_n3958_ = new_n3803_ & new_n3866_;
  assign new_n3959_ = new_n3805_ & new_n3866_;
  assign new_n3960_ = new_n3807_ & new_n3866_;
  assign new_n3961_ = ~new_n3959_ & ~new_n3960_;
  assign new_n3962_ = ~new_n3958_ & new_n3961_;
  assign new_n3963_ = new_n3811_ & new_n3866_;
  assign new_n3964_ = new_n3813_ & new_n3866_;
  assign new_n3965_ = new_n3815_ & new_n3866_;
  assign new_n3966_ = ~new_n3964_ & ~new_n3965_;
  assign new_n3967_ = ~new_n3963_ & new_n3966_;
  assign new_n3968_ = new_n3962_ & new_n3967_;
  assign new_n3969_ = new_n3821_ & new_n3866_;
  assign new_n3970_ = new_n3823_ & new_n3866_;
  assign new_n3971_ = new_n3825_ & new_n3866_;
  assign new_n3972_ = ~new_n3970_ & ~new_n3971_;
  assign new_n3973_ = ~new_n3969_ & new_n3972_;
  assign new_n3974_ = new_n3830_ & new_n3866_;
  assign new_n3975_ = new_n3832_ & new_n3866_;
  assign new_n3976_ = new_n3834_ & new_n3866_;
  assign new_n3977_ = ~new_n3975_ & ~new_n3976_;
  assign new_n3978_ = ~new_n3974_ & new_n3977_;
  assign new_n3979_ = new_n3973_ & new_n3978_;
  assign new_n3980_ = new_n3968_ & new_n3979_;
  assign new_n3981_ = new_n3840_ & new_n3866_;
  assign new_n3982_ = new_n3842_ & new_n3866_;
  assign new_n3983_ = new_n3844_ & new_n3866_;
  assign new_n3984_ = ~new_n3982_ & ~new_n3983_;
  assign new_n3985_ = ~new_n3981_ & new_n3984_;
  assign new_n3986_ = new_n3859_ & new_n3866_;
  assign new_n3987_ = new_n3848_ & new_n3866_;
  assign new_n3988_ = new_n3850_ & new_n3866_;
  assign new_n3989_ = ~new_n3987_ & ~new_n3988_;
  assign new_n3990_ = ~new_n3986_ & new_n3989_;
  assign new_n3991_ = new_n3985_ & new_n3990_;
  assign new_n3992_ = new_n3866_ & new_n3868_;
  assign new_n3993_ = new_n3861_ & new_n3866_;
  assign new_n3994_ = new_n3857_ & new_n3866_;
  assign new_n3995_ = ~new_n3993_ & ~new_n3994_;
  assign new_n3996_ = ~new_n3992_ & new_n3995_;
  assign new_n3997_ = new_n516_ & new_n541_;
  assign new_n3998_ = new_n3665_ & new_n3997_;
  assign new_n3999_ = new_n3668_ & new_n3998_;
  assign new_n4000_ = new_n3670_ & new_n3998_;
  assign new_n4001_ = ~new_n3999_ & ~new_n4000_;
  assign new_n4002_ = new_n3996_ & new_n4001_;
  assign new_n4003_ = new_n3991_ & new_n4002_;
  assign new_n4004_ = new_n3980_ & new_n4003_;
  assign new_n4005_ = new_n3957_ & new_n4004_;
  assign new_n4006_ = new_n3681_ & new_n3998_;
  assign new_n4007_ = new_n3662_ & new_n3998_;
  assign new_n4008_ = new_n3679_ & new_n3998_;
  assign new_n4009_ = ~new_n4007_ & ~new_n4008_;
  assign new_n4010_ = ~new_n4006_ & new_n4009_;
  assign new_n4011_ = new_n3689_ & new_n3998_;
  assign new_n4012_ = new_n3677_ & new_n3998_;
  assign new_n4013_ = new_n3687_ & new_n3998_;
  assign new_n4014_ = ~new_n4012_ & ~new_n4013_;
  assign new_n4015_ = ~new_n4011_ & new_n4014_;
  assign new_n4016_ = new_n4010_ & new_n4015_;
  assign new_n4017_ = new_n3698_ & new_n3998_;
  assign new_n4018_ = new_n3685_ & new_n3998_;
  assign new_n4019_ = new_n3696_ & new_n3998_;
  assign new_n4020_ = ~new_n4018_ & ~new_n4019_;
  assign new_n4021_ = ~new_n4017_ & new_n4020_;
  assign new_n4022_ = new_n3705_ & new_n3998_;
  assign new_n4023_ = new_n3694_ & new_n3998_;
  assign new_n4024_ = new_n3703_ & new_n3998_;
  assign new_n4025_ = ~new_n4023_ & ~new_n4024_;
  assign new_n4026_ = ~new_n4022_ & new_n4025_;
  assign new_n4027_ = new_n4021_ & new_n4026_;
  assign new_n4028_ = new_n4016_ & new_n4027_;
  assign new_n4029_ = new_n3711_ & new_n3998_;
  assign new_n4030_ = new_n3713_ & new_n3998_;
  assign new_n4031_ = new_n3715_ & new_n3998_;
  assign new_n4032_ = ~new_n4030_ & ~new_n4031_;
  assign new_n4033_ = ~new_n4029_ & new_n4032_;
  assign new_n4034_ = new_n3719_ & new_n3998_;
  assign new_n4035_ = new_n3721_ & new_n3998_;
  assign new_n4036_ = new_n3723_ & new_n3998_;
  assign new_n4037_ = ~new_n4035_ & ~new_n4036_;
  assign new_n4038_ = ~new_n4034_ & new_n4037_;
  assign new_n4039_ = new_n4033_ & new_n4038_;
  assign new_n4040_ = new_n3729_ & new_n3998_;
  assign new_n4041_ = new_n3731_ & new_n3998_;
  assign new_n4042_ = new_n3733_ & new_n3998_;
  assign new_n4043_ = ~new_n4041_ & ~new_n4042_;
  assign new_n4044_ = ~new_n4040_ & new_n4043_;
  assign new_n4045_ = new_n3740_ & new_n3998_;
  assign new_n4046_ = new_n3742_ & new_n3998_;
  assign new_n4047_ = ~new_n4045_ & ~new_n4046_;
  assign new_n4048_ = new_n4044_ & new_n4047_;
  assign new_n4049_ = new_n4039_ & new_n4048_;
  assign new_n4050_ = new_n4028_ & new_n4049_;
  assign new_n4051_ = new_n3753_ & new_n3998_;
  assign new_n4052_ = new_n3738_ & new_n3998_;
  assign new_n4053_ = new_n3751_ & new_n3998_;
  assign new_n4054_ = ~new_n4052_ & ~new_n4053_;
  assign new_n4055_ = ~new_n4051_ & new_n4054_;
  assign new_n4056_ = new_n3761_ & new_n3998_;
  assign new_n4057_ = new_n3749_ & new_n3998_;
  assign new_n4058_ = new_n3759_ & new_n3998_;
  assign new_n4059_ = ~new_n4057_ & ~new_n4058_;
  assign new_n4060_ = ~new_n4056_ & new_n4059_;
  assign new_n4061_ = new_n4055_ & new_n4060_;
  assign new_n4062_ = new_n3771_ & new_n3998_;
  assign new_n4063_ = new_n3757_ & new_n3998_;
  assign new_n4064_ = new_n3769_ & new_n3998_;
  assign new_n4065_ = ~new_n4063_ & ~new_n4064_;
  assign new_n4066_ = ~new_n4062_ & new_n4065_;
  assign new_n4067_ = new_n3778_ & new_n3998_;
  assign new_n4068_ = new_n3767_ & new_n3998_;
  assign new_n4069_ = new_n3775_ & new_n3998_;
  assign new_n4070_ = ~new_n4068_ & ~new_n4069_;
  assign new_n4071_ = ~new_n4067_ & new_n4070_;
  assign new_n4072_ = new_n4066_ & new_n4071_;
  assign new_n4073_ = new_n4061_ & new_n4072_;
  assign new_n4074_ = new_n3785_ & new_n3998_;
  assign new_n4075_ = new_n3787_ & new_n3998_;
  assign new_n4076_ = new_n3789_ & new_n3998_;
  assign new_n4077_ = ~new_n4075_ & ~new_n4076_;
  assign new_n4078_ = ~new_n4074_ & new_n4077_;
  assign new_n4079_ = new_n3793_ & new_n3998_;
  assign new_n4080_ = new_n3795_ & new_n3998_;
  assign new_n4081_ = new_n3797_ & new_n3998_;
  assign new_n4082_ = ~new_n4080_ & ~new_n4081_;
  assign new_n4083_ = ~new_n4079_ & new_n4082_;
  assign new_n4084_ = new_n4078_ & new_n4083_;
  assign new_n4085_ = new_n3803_ & new_n3998_;
  assign new_n4086_ = new_n3805_ & new_n3998_;
  assign new_n4087_ = new_n3807_ & new_n3998_;
  assign new_n4088_ = ~new_n4086_ & ~new_n4087_;
  assign new_n4089_ = ~new_n4085_ & new_n4088_;
  assign new_n4090_ = new_n3813_ & new_n3998_;
  assign new_n4091_ = new_n3815_ & new_n3998_;
  assign new_n4092_ = ~new_n4090_ & ~new_n4091_;
  assign new_n4093_ = new_n4089_ & new_n4092_;
  assign new_n4094_ = new_n4084_ & new_n4093_;
  assign new_n4095_ = new_n4073_ & new_n4094_;
  assign new_n4096_ = new_n4050_ & new_n4095_;
  assign new_n4097_ = new_n4005_ & new_n4096_;
  assign new_n4098_ = new_n3825_ & new_n3998_;
  assign new_n4099_ = new_n3811_ & new_n3998_;
  assign new_n4100_ = new_n3823_ & new_n3998_;
  assign new_n4101_ = ~new_n4099_ & ~new_n4100_;
  assign new_n4102_ = ~new_n4098_ & new_n4101_;
  assign new_n4103_ = new_n3834_ & new_n3998_;
  assign new_n4104_ = new_n3821_ & new_n3998_;
  assign new_n4105_ = new_n3832_ & new_n3998_;
  assign new_n4106_ = ~new_n4104_ & ~new_n4105_;
  assign new_n4107_ = ~new_n4103_ & new_n4106_;
  assign new_n4108_ = new_n4102_ & new_n4107_;
  assign new_n4109_ = new_n3844_ & new_n3998_;
  assign new_n4110_ = new_n3830_ & new_n3998_;
  assign new_n4111_ = new_n3842_ & new_n3998_;
  assign new_n4112_ = ~new_n4110_ & ~new_n4111_;
  assign new_n4113_ = ~new_n4109_ & new_n4112_;
  assign new_n4114_ = new_n3850_ & new_n3998_;
  assign new_n4115_ = new_n3840_ & new_n3998_;
  assign new_n4116_ = new_n3848_ & new_n3998_;
  assign new_n4117_ = ~new_n4115_ & ~new_n4116_;
  assign new_n4118_ = ~new_n4114_ & new_n4117_;
  assign new_n4119_ = new_n4113_ & new_n4118_;
  assign new_n4120_ = new_n4108_ & new_n4119_;
  assign new_n4121_ = new_n3857_ & new_n3998_;
  assign new_n4122_ = new_n3859_ & new_n3998_;
  assign new_n4123_ = new_n3861_ & new_n3998_;
  assign new_n4124_ = ~new_n4122_ & ~new_n4123_;
  assign new_n4125_ = ~new_n4121_ & new_n4124_;
  assign new_n4126_ = new_n533_ & new_n541_;
  assign new_n4127_ = new_n3665_ & new_n4126_;
  assign new_n4128_ = new_n3670_ & new_n4127_;
  assign new_n4129_ = new_n3868_ & new_n3998_;
  assign new_n4130_ = new_n3668_ & new_n4127_;
  assign new_n4131_ = ~new_n4129_ & ~new_n4130_;
  assign new_n4132_ = ~new_n4128_ & new_n4131_;
  assign new_n4133_ = new_n4125_ & new_n4132_;
  assign new_n4134_ = new_n3681_ & new_n4127_;
  assign new_n4135_ = new_n3662_ & new_n4127_;
  assign new_n4136_ = new_n3679_ & new_n4127_;
  assign new_n4137_ = ~new_n4135_ & ~new_n4136_;
  assign new_n4138_ = ~new_n4134_ & new_n4137_;
  assign new_n4139_ = new_n3677_ & new_n4127_;
  assign new_n4140_ = new_n3687_ & new_n4127_;
  assign new_n4141_ = ~new_n4139_ & ~new_n4140_;
  assign new_n4142_ = new_n4138_ & new_n4141_;
  assign new_n4143_ = new_n4133_ & new_n4142_;
  assign new_n4144_ = new_n4120_ & new_n4143_;
  assign new_n4145_ = new_n3696_ & new_n4127_;
  assign new_n4146_ = new_n3689_ & new_n4127_;
  assign new_n4147_ = new_n3685_ & new_n4127_;
  assign new_n4148_ = ~new_n4146_ & ~new_n4147_;
  assign new_n4149_ = ~new_n4145_ & new_n4148_;
  assign new_n4150_ = new_n3703_ & new_n4127_;
  assign new_n4151_ = new_n3698_ & new_n4127_;
  assign new_n4152_ = new_n3694_ & new_n4127_;
  assign new_n4153_ = ~new_n4151_ & ~new_n4152_;
  assign new_n4154_ = ~new_n4150_ & new_n4153_;
  assign new_n4155_ = new_n4149_ & new_n4154_;
  assign new_n4156_ = new_n3715_ & new_n4127_;
  assign new_n4157_ = new_n3705_ & new_n4127_;
  assign new_n4158_ = new_n3713_ & new_n4127_;
  assign new_n4159_ = ~new_n4157_ & ~new_n4158_;
  assign new_n4160_ = ~new_n4156_ & new_n4159_;
  assign new_n4161_ = new_n3723_ & new_n4127_;
  assign new_n4162_ = new_n3711_ & new_n4127_;
  assign new_n4163_ = new_n3721_ & new_n4127_;
  assign new_n4164_ = ~new_n4162_ & ~new_n4163_;
  assign new_n4165_ = ~new_n4161_ & new_n4164_;
  assign new_n4166_ = new_n4160_ & new_n4165_;
  assign new_n4167_ = new_n4155_ & new_n4166_;
  assign new_n4168_ = new_n3733_ & new_n4127_;
  assign new_n4169_ = new_n3719_ & new_n4127_;
  assign new_n4170_ = new_n3731_ & new_n4127_;
  assign new_n4171_ = ~new_n4169_ & ~new_n4170_;
  assign new_n4172_ = ~new_n4168_ & new_n4171_;
  assign new_n4173_ = new_n3742_ & new_n4127_;
  assign new_n4174_ = new_n3729_ & new_n4127_;
  assign new_n4175_ = new_n3740_ & new_n4127_;
  assign new_n4176_ = ~new_n4174_ & ~new_n4175_;
  assign new_n4177_ = ~new_n4173_ & new_n4176_;
  assign new_n4178_ = new_n4172_ & new_n4177_;
  assign new_n4179_ = new_n3753_ & new_n4127_;
  assign new_n4180_ = new_n3738_ & new_n4127_;
  assign new_n4181_ = new_n3751_ & new_n4127_;
  assign new_n4182_ = ~new_n4180_ & ~new_n4181_;
  assign new_n4183_ = ~new_n4179_ & new_n4182_;
  assign new_n4184_ = new_n3749_ & new_n4127_;
  assign new_n4185_ = new_n3759_ & new_n4127_;
  assign new_n4186_ = ~new_n4184_ & ~new_n4185_;
  assign new_n4187_ = new_n4183_ & new_n4186_;
  assign new_n4188_ = new_n4178_ & new_n4187_;
  assign new_n4189_ = new_n4167_ & new_n4188_;
  assign new_n4190_ = new_n4144_ & new_n4189_;
  assign new_n4191_ = new_n3769_ & new_n4127_;
  assign new_n4192_ = new_n3761_ & new_n4127_;
  assign new_n4193_ = new_n3757_ & new_n4127_;
  assign new_n4194_ = ~new_n4192_ & ~new_n4193_;
  assign new_n4195_ = ~new_n4191_ & new_n4194_;
  assign new_n4196_ = new_n3775_ & new_n4127_;
  assign new_n4197_ = new_n3771_ & new_n4127_;
  assign new_n4198_ = new_n3767_ & new_n4127_;
  assign new_n4199_ = ~new_n4197_ & ~new_n4198_;
  assign new_n4200_ = ~new_n4196_ & new_n4199_;
  assign new_n4201_ = new_n4195_ & new_n4200_;
  assign new_n4202_ = new_n3789_ & new_n4127_;
  assign new_n4203_ = new_n3778_ & new_n4127_;
  assign new_n4204_ = new_n3787_ & new_n4127_;
  assign new_n4205_ = ~new_n4203_ & ~new_n4204_;
  assign new_n4206_ = ~new_n4202_ & new_n4205_;
  assign new_n4207_ = new_n3797_ & new_n4127_;
  assign new_n4208_ = new_n3785_ & new_n4127_;
  assign new_n4209_ = new_n3795_ & new_n4127_;
  assign new_n4210_ = ~new_n4208_ & ~new_n4209_;
  assign new_n4211_ = ~new_n4207_ & new_n4210_;
  assign new_n4212_ = new_n4206_ & new_n4211_;
  assign new_n4213_ = new_n4201_ & new_n4212_;
  assign new_n4214_ = new_n3807_ & new_n4127_;
  assign new_n4215_ = new_n3793_ & new_n4127_;
  assign new_n4216_ = new_n3805_ & new_n4127_;
  assign new_n4217_ = ~new_n4215_ & ~new_n4216_;
  assign new_n4218_ = ~new_n4214_ & new_n4217_;
  assign new_n4219_ = new_n3815_ & new_n4127_;
  assign new_n4220_ = new_n3803_ & new_n4127_;
  assign new_n4221_ = new_n3813_ & new_n4127_;
  assign new_n4222_ = ~new_n4220_ & ~new_n4221_;
  assign new_n4223_ = ~new_n4219_ & new_n4222_;
  assign new_n4224_ = new_n4218_ & new_n4223_;
  assign new_n4225_ = new_n3825_ & new_n4127_;
  assign new_n4226_ = new_n3811_ & new_n4127_;
  assign new_n4227_ = new_n3823_ & new_n4127_;
  assign new_n4228_ = ~new_n4226_ & ~new_n4227_;
  assign new_n4229_ = ~new_n4225_ & new_n4228_;
  assign new_n4230_ = new_n3821_ & new_n4127_;
  assign new_n4231_ = new_n3832_ & new_n4127_;
  assign new_n4232_ = ~new_n4230_ & ~new_n4231_;
  assign new_n4233_ = new_n4229_ & new_n4232_;
  assign new_n4234_ = new_n4224_ & new_n4233_;
  assign new_n4235_ = new_n4213_ & new_n4234_;
  assign new_n4236_ = new_n3842_ & new_n4127_;
  assign new_n4237_ = new_n3834_ & new_n4127_;
  assign new_n4238_ = new_n3830_ & new_n4127_;
  assign new_n4239_ = ~new_n4237_ & ~new_n4238_;
  assign new_n4240_ = ~new_n4236_ & new_n4239_;
  assign new_n4241_ = new_n3848_ & new_n4127_;
  assign new_n4242_ = new_n3844_ & new_n4127_;
  assign new_n4243_ = new_n3840_ & new_n4127_;
  assign new_n4244_ = ~new_n4242_ & ~new_n4243_;
  assign new_n4245_ = ~new_n4241_ & new_n4244_;
  assign new_n4246_ = new_n4240_ & new_n4245_;
  assign new_n4247_ = new_n3861_ & new_n4127_;
  assign new_n4248_ = new_n3850_ & new_n4127_;
  assign new_n4249_ = new_n3859_ & new_n4127_;
  assign new_n4250_ = ~new_n4248_ & ~new_n4249_;
  assign new_n4251_ = ~new_n4247_ & new_n4250_;
  assign new_n4252_ = ~A200 & ~A199;
  assign new_n4253_ = new_n1781_ & new_n4252_;
  assign new_n4254_ = A168 & ~A169;
  assign new_n4255_ = ~A170 & new_n4254_;
  assign new_n4256_ = new_n4253_ & new_n4255_;
  assign new_n4257_ = new_n1735_ & new_n4256_;
  assign new_n4258_ = new_n3857_ & new_n4127_;
  assign new_n4259_ = new_n3868_ & new_n4127_;
  assign new_n4260_ = ~new_n4258_ & ~new_n4259_;
  assign new_n4261_ = ~new_n4257_ & new_n4260_;
  assign new_n4262_ = new_n4251_ & new_n4261_;
  assign new_n4263_ = new_n4246_ & new_n4262_;
  assign new_n4264_ = new_n1749_ & new_n4256_;
  assign new_n4265_ = new_n1738_ & new_n4256_;
  assign new_n4266_ = new_n1725_ & new_n4256_;
  assign new_n4267_ = ~new_n4265_ & ~new_n4266_;
  assign new_n4268_ = ~new_n4264_ & new_n4267_;
  assign new_n4269_ = new_n1795_ & new_n4252_;
  assign new_n4270_ = new_n4255_ & new_n4269_;
  assign new_n4271_ = new_n1725_ & new_n4270_;
  assign new_n4272_ = new_n1735_ & new_n4270_;
  assign new_n4273_ = new_n1738_ & new_n4270_;
  assign new_n4274_ = ~new_n4272_ & ~new_n4273_;
  assign new_n4275_ = ~new_n4271_ & new_n4274_;
  assign new_n4276_ = new_n4268_ & new_n4275_;
  assign new_n4277_ = new_n1804_ & new_n4252_;
  assign new_n4278_ = new_n4255_ & new_n4277_;
  assign new_n4279_ = new_n1738_ & new_n4278_;
  assign new_n4280_ = new_n1749_ & new_n4270_;
  assign new_n4281_ = new_n1735_ & new_n4278_;
  assign new_n4282_ = ~new_n4280_ & ~new_n4281_;
  assign new_n4283_ = ~new_n4279_ & new_n4282_;
  assign new_n4284_ = new_n1725_ & new_n4278_;
  assign new_n4285_ = new_n1749_ & new_n4278_;
  assign new_n4286_ = ~new_n4284_ & ~new_n4285_;
  assign new_n4287_ = new_n4283_ & new_n4286_;
  assign new_n4288_ = new_n4276_ & new_n4287_;
  assign new_n4289_ = new_n4263_ & new_n4288_;
  assign new_n4290_ = new_n4235_ & new_n4289_;
  assign new_n4291_ = new_n4190_ & new_n4290_;
  assign new_n4292_ = new_n4097_ & new_n4291_;
  assign new_n4293_ = new_n3910_ & new_n4292_;
  assign new_n4294_ = new_n1812_ & new_n4252_;
  assign new_n4295_ = new_n4255_ & new_n4294_;
  assign new_n4296_ = new_n1725_ & new_n4295_;
  assign new_n4297_ = new_n1735_ & new_n4295_;
  assign new_n4298_ = new_n1738_ & new_n4295_;
  assign new_n4299_ = ~new_n4297_ & ~new_n4298_;
  assign new_n4300_ = ~new_n4296_ & new_n4299_;
  assign new_n4301_ = new_n504_ & new_n4252_;
  assign new_n4302_ = new_n4255_ & new_n4301_;
  assign new_n4303_ = new_n1833_ & new_n4302_;
  assign new_n4304_ = new_n1749_ & new_n4295_;
  assign new_n4305_ = new_n1830_ & new_n4302_;
  assign new_n4306_ = ~new_n4304_ & ~new_n4305_;
  assign new_n4307_ = ~new_n4303_ & new_n4306_;
  assign new_n4308_ = new_n4300_ & new_n4307_;
  assign new_n4309_ = new_n1842_ & new_n4302_;
  assign new_n4310_ = new_n1827_ & new_n4302_;
  assign new_n4311_ = new_n1840_ & new_n4302_;
  assign new_n4312_ = ~new_n4310_ & ~new_n4311_;
  assign new_n4313_ = ~new_n4309_ & new_n4312_;
  assign new_n4314_ = new_n1849_ & new_n4302_;
  assign new_n4315_ = new_n1838_ & new_n4302_;
  assign new_n4316_ = new_n1847_ & new_n4302_;
  assign new_n4317_ = ~new_n4315_ & ~new_n4316_;
  assign new_n4318_ = ~new_n4314_ & new_n4317_;
  assign new_n4319_ = new_n4313_ & new_n4318_;
  assign new_n4320_ = new_n4308_ & new_n4319_;
  assign new_n4321_ = new_n1855_ & new_n4302_;
  assign new_n4322_ = new_n1857_ & new_n4302_;
  assign new_n4323_ = new_n1859_ & new_n4302_;
  assign new_n4324_ = ~new_n4322_ & ~new_n4323_;
  assign new_n4325_ = ~new_n4321_ & new_n4324_;
  assign new_n4326_ = new_n1864_ & new_n4302_;
  assign new_n4327_ = new_n1866_ & new_n4302_;
  assign new_n4328_ = new_n1868_ & new_n4302_;
  assign new_n4329_ = ~new_n4327_ & ~new_n4328_;
  assign new_n4330_ = ~new_n4326_ & new_n4329_;
  assign new_n4331_ = new_n4325_ & new_n4330_;
  assign new_n4332_ = new_n1875_ & new_n4302_;
  assign new_n4333_ = new_n1878_ & new_n4302_;
  assign new_n4334_ = new_n1881_ & new_n4302_;
  assign new_n4335_ = ~new_n4333_ & ~new_n4334_;
  assign new_n4336_ = ~new_n4332_ & new_n4335_;
  assign new_n4337_ = new_n1886_ & new_n4302_;
  assign new_n4338_ = new_n1889_ & new_n4302_;
  assign new_n4339_ = new_n1892_ & new_n4302_;
  assign new_n4340_ = ~new_n4338_ & ~new_n4339_;
  assign new_n4341_ = ~new_n4337_ & new_n4340_;
  assign new_n4342_ = new_n4336_ & new_n4341_;
  assign new_n4343_ = new_n4331_ & new_n4342_;
  assign new_n4344_ = new_n4320_ & new_n4343_;
  assign new_n4345_ = new_n1898_ & new_n4302_;
  assign new_n4346_ = new_n1900_ & new_n4302_;
  assign new_n4347_ = new_n1902_ & new_n4302_;
  assign new_n4348_ = ~new_n4346_ & ~new_n4347_;
  assign new_n4349_ = ~new_n4345_ & new_n4348_;
  assign new_n4350_ = A200 & A199;
  assign new_n4351_ = new_n1781_ & new_n4350_;
  assign new_n4352_ = new_n4255_ & new_n4351_;
  assign new_n4353_ = new_n1738_ & new_n4352_;
  assign new_n4354_ = new_n1913_ & new_n4302_;
  assign new_n4355_ = new_n1735_ & new_n4352_;
  assign new_n4356_ = ~new_n4354_ & ~new_n4355_;
  assign new_n4357_ = ~new_n4353_ & new_n4356_;
  assign new_n4358_ = new_n4349_ & new_n4357_;
  assign new_n4359_ = new_n1795_ & new_n4350_;
  assign new_n4360_ = new_n4255_ & new_n4359_;
  assign new_n4361_ = new_n1735_ & new_n4360_;
  assign new_n4362_ = new_n1725_ & new_n4352_;
  assign new_n4363_ = new_n1749_ & new_n4352_;
  assign new_n4364_ = ~new_n4362_ & ~new_n4363_;
  assign new_n4365_ = ~new_n4361_ & new_n4364_;
  assign new_n4366_ = new_n1749_ & new_n4360_;
  assign new_n4367_ = new_n1738_ & new_n4360_;
  assign new_n4368_ = new_n1725_ & new_n4360_;
  assign new_n4369_ = ~new_n4367_ & ~new_n4368_;
  assign new_n4370_ = ~new_n4366_ & new_n4369_;
  assign new_n4371_ = new_n4365_ & new_n4370_;
  assign new_n4372_ = new_n4358_ & new_n4371_;
  assign new_n4373_ = new_n1804_ & new_n4350_;
  assign new_n4374_ = new_n4255_ & new_n4373_;
  assign new_n4375_ = new_n1725_ & new_n4374_;
  assign new_n4376_ = new_n1735_ & new_n4374_;
  assign new_n4377_ = new_n1738_ & new_n4374_;
  assign new_n4378_ = ~new_n4376_ & ~new_n4377_;
  assign new_n4379_ = ~new_n4375_ & new_n4378_;
  assign new_n4380_ = new_n1812_ & new_n4350_;
  assign new_n4381_ = new_n4255_ & new_n4380_;
  assign new_n4382_ = new_n1738_ & new_n4381_;
  assign new_n4383_ = new_n1749_ & new_n4374_;
  assign new_n4384_ = new_n1735_ & new_n4381_;
  assign new_n4385_ = ~new_n4383_ & ~new_n4384_;
  assign new_n4386_ = ~new_n4382_ & new_n4385_;
  assign new_n4387_ = new_n4379_ & new_n4386_;
  assign new_n4388_ = new_n504_ & new_n4350_;
  assign new_n4389_ = new_n4255_ & new_n4388_;
  assign new_n4390_ = new_n1830_ & new_n4389_;
  assign new_n4391_ = new_n1725_ & new_n4381_;
  assign new_n4392_ = new_n1749_ & new_n4381_;
  assign new_n4393_ = ~new_n4391_ & ~new_n4392_;
  assign new_n4394_ = ~new_n4390_ & new_n4393_;
  assign new_n4395_ = new_n1833_ & new_n4389_;
  assign new_n4396_ = new_n1827_ & new_n4389_;
  assign new_n4397_ = ~new_n4395_ & ~new_n4396_;
  assign new_n4398_ = new_n4394_ & new_n4397_;
  assign new_n4399_ = new_n4387_ & new_n4398_;
  assign new_n4400_ = new_n4372_ & new_n4399_;
  assign new_n4401_ = new_n4344_ & new_n4400_;
  assign new_n4402_ = new_n1838_ & new_n4389_;
  assign new_n4403_ = new_n1840_ & new_n4389_;
  assign new_n4404_ = new_n1842_ & new_n4389_;
  assign new_n4405_ = ~new_n4403_ & ~new_n4404_;
  assign new_n4406_ = ~new_n4402_ & new_n4405_;
  assign new_n4407_ = new_n1857_ & new_n4389_;
  assign new_n4408_ = new_n1847_ & new_n4389_;
  assign new_n4409_ = new_n1849_ & new_n4389_;
  assign new_n4410_ = ~new_n4408_ & ~new_n4409_;
  assign new_n4411_ = ~new_n4407_ & new_n4410_;
  assign new_n4412_ = new_n4406_ & new_n4411_;
  assign new_n4413_ = new_n1866_ & new_n4389_;
  assign new_n4414_ = new_n1859_ & new_n4389_;
  assign new_n4415_ = new_n1855_ & new_n4389_;
  assign new_n4416_ = ~new_n4414_ & ~new_n4415_;
  assign new_n4417_ = ~new_n4413_ & new_n4416_;
  assign new_n4418_ = new_n1878_ & new_n4389_;
  assign new_n4419_ = new_n1868_ & new_n4389_;
  assign new_n4420_ = new_n1864_ & new_n4389_;
  assign new_n4421_ = ~new_n4419_ & ~new_n4420_;
  assign new_n4422_ = ~new_n4418_ & new_n4421_;
  assign new_n4423_ = new_n4417_ & new_n4422_;
  assign new_n4424_ = new_n4412_ & new_n4423_;
  assign new_n4425_ = new_n1889_ & new_n4389_;
  assign new_n4426_ = new_n1881_ & new_n4389_;
  assign new_n4427_ = new_n1875_ & new_n4389_;
  assign new_n4428_ = ~new_n4426_ & ~new_n4427_;
  assign new_n4429_ = ~new_n4425_ & new_n4428_;
  assign new_n4430_ = new_n1900_ & new_n4389_;
  assign new_n4431_ = new_n1892_ & new_n4389_;
  assign new_n4432_ = new_n1886_ & new_n4389_;
  assign new_n4433_ = ~new_n4431_ & ~new_n4432_;
  assign new_n4434_ = ~new_n4430_ & new_n4433_;
  assign new_n4435_ = new_n4429_ & new_n4434_;
  assign new_n4436_ = new_n1913_ & new_n4389_;
  assign new_n4437_ = new_n1902_ & new_n4389_;
  assign new_n4438_ = new_n1898_ & new_n4389_;
  assign new_n4439_ = ~new_n4437_ & ~new_n4438_;
  assign new_n4440_ = ~new_n4436_ & new_n4439_;
  assign new_n4441_ = ~A203 & ~A201;
  assign new_n4442_ = new_n1781_ & new_n4441_;
  assign new_n4443_ = new_n4255_ & new_n4442_;
  assign new_n4444_ = new_n1735_ & new_n4443_;
  assign new_n4445_ = new_n1738_ & new_n4443_;
  assign new_n4446_ = ~new_n4444_ & ~new_n4445_;
  assign new_n4447_ = new_n4440_ & new_n4446_;
  assign new_n4448_ = new_n4435_ & new_n4447_;
  assign new_n4449_ = new_n4424_ & new_n4448_;
  assign new_n4450_ = new_n1795_ & new_n4441_;
  assign new_n4451_ = new_n4255_ & new_n4450_;
  assign new_n4452_ = new_n1735_ & new_n4451_;
  assign new_n4453_ = new_n1725_ & new_n4443_;
  assign new_n4454_ = new_n1749_ & new_n4443_;
  assign new_n4455_ = ~new_n4453_ & ~new_n4454_;
  assign new_n4456_ = ~new_n4452_ & new_n4455_;
  assign new_n4457_ = new_n1749_ & new_n4451_;
  assign new_n4458_ = new_n1738_ & new_n4451_;
  assign new_n4459_ = new_n1725_ & new_n4451_;
  assign new_n4460_ = ~new_n4458_ & ~new_n4459_;
  assign new_n4461_ = ~new_n4457_ & new_n4460_;
  assign new_n4462_ = new_n4456_ & new_n4461_;
  assign new_n4463_ = new_n1804_ & new_n4441_;
  assign new_n4464_ = new_n4255_ & new_n4463_;
  assign new_n4465_ = new_n1725_ & new_n4464_;
  assign new_n4466_ = new_n1735_ & new_n4464_;
  assign new_n4467_ = new_n1738_ & new_n4464_;
  assign new_n4468_ = ~new_n4466_ & ~new_n4467_;
  assign new_n4469_ = ~new_n4465_ & new_n4468_;
  assign new_n4470_ = new_n1812_ & new_n4441_;
  assign new_n4471_ = new_n4255_ & new_n4470_;
  assign new_n4472_ = new_n1738_ & new_n4471_;
  assign new_n4473_ = new_n1749_ & new_n4464_;
  assign new_n4474_ = new_n1735_ & new_n4471_;
  assign new_n4475_ = ~new_n4473_ & ~new_n4474_;
  assign new_n4476_ = ~new_n4472_ & new_n4475_;
  assign new_n4477_ = new_n4469_ & new_n4476_;
  assign new_n4478_ = new_n4462_ & new_n4477_;
  assign new_n4479_ = new_n504_ & new_n4441_;
  assign new_n4480_ = new_n4255_ & new_n4479_;
  assign new_n4481_ = new_n1830_ & new_n4480_;
  assign new_n4482_ = new_n1725_ & new_n4471_;
  assign new_n4483_ = new_n1749_ & new_n4471_;
  assign new_n4484_ = ~new_n4482_ & ~new_n4483_;
  assign new_n4485_ = ~new_n4481_ & new_n4484_;
  assign new_n4486_ = new_n1840_ & new_n4480_;
  assign new_n4487_ = new_n1833_ & new_n4480_;
  assign new_n4488_ = new_n1827_ & new_n4480_;
  assign new_n4489_ = ~new_n4487_ & ~new_n4488_;
  assign new_n4490_ = ~new_n4486_ & new_n4489_;
  assign new_n4491_ = new_n4485_ & new_n4490_;
  assign new_n4492_ = new_n1847_ & new_n4480_;
  assign new_n4493_ = new_n1842_ & new_n4480_;
  assign new_n4494_ = new_n1838_ & new_n4480_;
  assign new_n4495_ = ~new_n4493_ & ~new_n4494_;
  assign new_n4496_ = ~new_n4492_ & new_n4495_;
  assign new_n4497_ = new_n1849_ & new_n4480_;
  assign new_n4498_ = new_n1857_ & new_n4480_;
  assign new_n4499_ = ~new_n4497_ & ~new_n4498_;
  assign new_n4500_ = new_n4496_ & new_n4499_;
  assign new_n4501_ = new_n4491_ & new_n4500_;
  assign new_n4502_ = new_n4478_ & new_n4501_;
  assign new_n4503_ = new_n4449_ & new_n4502_;
  assign new_n4504_ = new_n4401_ & new_n4503_;
  assign new_n4505_ = new_n1866_ & new_n4480_;
  assign new_n4506_ = new_n1859_ & new_n4480_;
  assign new_n4507_ = new_n1855_ & new_n4480_;
  assign new_n4508_ = ~new_n4506_ & ~new_n4507_;
  assign new_n4509_ = ~new_n4505_ & new_n4508_;
  assign new_n4510_ = new_n1878_ & new_n4480_;
  assign new_n4511_ = new_n1868_ & new_n4480_;
  assign new_n4512_ = new_n1864_ & new_n4480_;
  assign new_n4513_ = ~new_n4511_ & ~new_n4512_;
  assign new_n4514_ = ~new_n4510_ & new_n4513_;
  assign new_n4515_ = new_n4509_ & new_n4514_;
  assign new_n4516_ = new_n1889_ & new_n4480_;
  assign new_n4517_ = new_n1881_ & new_n4480_;
  assign new_n4518_ = new_n1875_ & new_n4480_;
  assign new_n4519_ = ~new_n4517_ & ~new_n4518_;
  assign new_n4520_ = ~new_n4516_ & new_n4519_;
  assign new_n4521_ = new_n1900_ & new_n4480_;
  assign new_n4522_ = new_n1892_ & new_n4480_;
  assign new_n4523_ = new_n1886_ & new_n4480_;
  assign new_n4524_ = ~new_n4522_ & ~new_n4523_;
  assign new_n4525_ = ~new_n4521_ & new_n4524_;
  assign new_n4526_ = new_n4520_ & new_n4525_;
  assign new_n4527_ = new_n4515_ & new_n4526_;
  assign new_n4528_ = new_n1913_ & new_n4480_;
  assign new_n4529_ = new_n1902_ & new_n4480_;
  assign new_n4530_ = new_n1898_ & new_n4480_;
  assign new_n4531_ = ~new_n4529_ & ~new_n4530_;
  assign new_n4532_ = ~new_n4528_ & new_n4531_;
  assign new_n4533_ = A202 & ~A201;
  assign new_n4534_ = new_n1781_ & new_n4533_;
  assign new_n4535_ = new_n4255_ & new_n4534_;
  assign new_n4536_ = new_n1725_ & new_n4535_;
  assign new_n4537_ = new_n1735_ & new_n4535_;
  assign new_n4538_ = new_n1738_ & new_n4535_;
  assign new_n4539_ = ~new_n4537_ & ~new_n4538_;
  assign new_n4540_ = ~new_n4536_ & new_n4539_;
  assign new_n4541_ = new_n4532_ & new_n4540_;
  assign new_n4542_ = new_n1795_ & new_n4533_;
  assign new_n4543_ = new_n4255_ & new_n4542_;
  assign new_n4544_ = new_n1738_ & new_n4543_;
  assign new_n4545_ = new_n1749_ & new_n4535_;
  assign new_n4546_ = new_n1735_ & new_n4543_;
  assign new_n4547_ = ~new_n4545_ & ~new_n4546_;
  assign new_n4548_ = ~new_n4544_ & new_n4547_;
  assign new_n4549_ = new_n1725_ & new_n4543_;
  assign new_n4550_ = new_n1749_ & new_n4543_;
  assign new_n4551_ = ~new_n4549_ & ~new_n4550_;
  assign new_n4552_ = new_n4548_ & new_n4551_;
  assign new_n4553_ = new_n4541_ & new_n4552_;
  assign new_n4554_ = new_n4527_ & new_n4553_;
  assign new_n4555_ = new_n1804_ & new_n4533_;
  assign new_n4556_ = new_n4255_ & new_n4555_;
  assign new_n4557_ = new_n1725_ & new_n4556_;
  assign new_n4558_ = new_n1735_ & new_n4556_;
  assign new_n4559_ = new_n1738_ & new_n4556_;
  assign new_n4560_ = ~new_n4558_ & ~new_n4559_;
  assign new_n4561_ = ~new_n4557_ & new_n4560_;
  assign new_n4562_ = new_n1812_ & new_n4533_;
  assign new_n4563_ = new_n4255_ & new_n4562_;
  assign new_n4564_ = new_n1738_ & new_n4563_;
  assign new_n4565_ = new_n1749_ & new_n4556_;
  assign new_n4566_ = new_n1735_ & new_n4563_;
  assign new_n4567_ = ~new_n4565_ & ~new_n4566_;
  assign new_n4568_ = ~new_n4564_ & new_n4567_;
  assign new_n4569_ = new_n4561_ & new_n4568_;
  assign new_n4570_ = new_n504_ & new_n4533_;
  assign new_n4571_ = new_n4255_ & new_n4570_;
  assign new_n4572_ = new_n1830_ & new_n4571_;
  assign new_n4573_ = new_n1725_ & new_n4563_;
  assign new_n4574_ = new_n1749_ & new_n4563_;
  assign new_n4575_ = ~new_n4573_ & ~new_n4574_;
  assign new_n4576_ = ~new_n4572_ & new_n4575_;
  assign new_n4577_ = new_n1840_ & new_n4571_;
  assign new_n4578_ = new_n1833_ & new_n4571_;
  assign new_n4579_ = new_n1827_ & new_n4571_;
  assign new_n4580_ = ~new_n4578_ & ~new_n4579_;
  assign new_n4581_ = ~new_n4577_ & new_n4580_;
  assign new_n4582_ = new_n4576_ & new_n4581_;
  assign new_n4583_ = new_n4569_ & new_n4582_;
  assign new_n4584_ = new_n1847_ & new_n4571_;
  assign new_n4585_ = new_n1842_ & new_n4571_;
  assign new_n4586_ = new_n1838_ & new_n4571_;
  assign new_n4587_ = ~new_n4585_ & ~new_n4586_;
  assign new_n4588_ = ~new_n4584_ & new_n4587_;
  assign new_n4589_ = new_n1859_ & new_n4571_;
  assign new_n4590_ = new_n1849_ & new_n4571_;
  assign new_n4591_ = new_n1857_ & new_n4571_;
  assign new_n4592_ = ~new_n4590_ & ~new_n4591_;
  assign new_n4593_ = ~new_n4589_ & new_n4592_;
  assign new_n4594_ = new_n4588_ & new_n4593_;
  assign new_n4595_ = new_n1868_ & new_n4571_;
  assign new_n4596_ = new_n1855_ & new_n4571_;
  assign new_n4597_ = new_n1866_ & new_n4571_;
  assign new_n4598_ = ~new_n4596_ & ~new_n4597_;
  assign new_n4599_ = ~new_n4595_ & new_n4598_;
  assign new_n4600_ = new_n1864_ & new_n4571_;
  assign new_n4601_ = new_n1878_ & new_n4571_;
  assign new_n4602_ = ~new_n4600_ & ~new_n4601_;
  assign new_n4603_ = new_n4599_ & new_n4602_;
  assign new_n4604_ = new_n4594_ & new_n4603_;
  assign new_n4605_ = new_n4583_ & new_n4604_;
  assign new_n4606_ = new_n4554_ & new_n4605_;
  assign new_n4607_ = new_n1889_ & new_n4571_;
  assign new_n4608_ = new_n1881_ & new_n4571_;
  assign new_n4609_ = new_n1875_ & new_n4571_;
  assign new_n4610_ = ~new_n4608_ & ~new_n4609_;
  assign new_n4611_ = ~new_n4607_ & new_n4610_;
  assign new_n4612_ = new_n1900_ & new_n4571_;
  assign new_n4613_ = new_n1892_ & new_n4571_;
  assign new_n4614_ = new_n1886_ & new_n4571_;
  assign new_n4615_ = ~new_n4613_ & ~new_n4614_;
  assign new_n4616_ = ~new_n4612_ & new_n4615_;
  assign new_n4617_ = new_n4611_ & new_n4616_;
  assign new_n4618_ = new_n1913_ & new_n4571_;
  assign new_n4619_ = new_n1902_ & new_n4571_;
  assign new_n4620_ = new_n1898_ & new_n4571_;
  assign new_n4621_ = ~new_n4619_ & ~new_n4620_;
  assign new_n4622_ = ~new_n4618_ & new_n4621_;
  assign new_n4623_ = A265 & ~A233;
  assign new_n4624_ = new_n46_ & new_n4623_;
  assign new_n4625_ = new_n1058_ & new_n4624_;
  assign new_n4626_ = new_n108_ & new_n1908_;
  assign new_n4627_ = new_n4255_ & new_n4626_;
  assign new_n4628_ = new_n4625_ & new_n4627_;
  assign new_n4629_ = ~A265 & ~A233;
  assign new_n4630_ = new_n1063_ & new_n4629_;
  assign new_n4631_ = new_n1062_ & new_n4630_;
  assign new_n4632_ = new_n4627_ & new_n4631_;
  assign new_n4633_ = new_n1069_ & new_n4629_;
  assign new_n4634_ = new_n1068_ & new_n4633_;
  assign new_n4635_ = new_n4627_ & new_n4634_;
  assign new_n4636_ = ~new_n4632_ & ~new_n4635_;
  assign new_n4637_ = ~new_n4628_ & new_n4636_;
  assign new_n4638_ = new_n4622_ & new_n4637_;
  assign new_n4639_ = new_n4617_ & new_n4638_;
  assign new_n4640_ = new_n1075_ & new_n4624_;
  assign new_n4641_ = new_n4627_ & new_n4640_;
  assign new_n4642_ = new_n1078_ & new_n4624_;
  assign new_n4643_ = new_n4627_ & new_n4642_;
  assign new_n4644_ = new_n1081_ & new_n4624_;
  assign new_n4645_ = new_n4627_ & new_n4644_;
  assign new_n4646_ = ~new_n4643_ & ~new_n4645_;
  assign new_n4647_ = ~new_n4641_ & new_n4646_;
  assign new_n4648_ = new_n51_ & new_n4629_;
  assign new_n4649_ = new_n1058_ & new_n4648_;
  assign new_n4650_ = new_n4627_ & new_n4649_;
  assign new_n4651_ = new_n1093_ & new_n4623_;
  assign new_n4652_ = new_n1092_ & new_n4651_;
  assign new_n4653_ = new_n4627_ & new_n4652_;
  assign new_n4654_ = new_n1098_ & new_n4651_;
  assign new_n4655_ = new_n4627_ & new_n4654_;
  assign new_n4656_ = ~new_n4653_ & ~new_n4655_;
  assign new_n4657_ = ~new_n4650_ & new_n4656_;
  assign new_n4658_ = new_n4647_ & new_n4657_;
  assign new_n4659_ = new_n1075_ & new_n4648_;
  assign new_n4660_ = new_n4627_ & new_n4659_;
  assign new_n4661_ = new_n1078_ & new_n4648_;
  assign new_n4662_ = new_n4627_ & new_n4661_;
  assign new_n4663_ = new_n1081_ & new_n4648_;
  assign new_n4664_ = new_n4627_ & new_n4663_;
  assign new_n4665_ = ~new_n4662_ & ~new_n4664_;
  assign new_n4666_ = ~new_n4660_ & new_n4665_;
  assign new_n4667_ = new_n1116_ & new_n4629_;
  assign new_n4668_ = new_n1092_ & new_n4667_;
  assign new_n4669_ = new_n4627_ & new_n4668_;
  assign new_n4670_ = new_n1098_ & new_n4667_;
  assign new_n4671_ = new_n4627_ & new_n4670_;
  assign new_n4672_ = ~new_n4669_ & ~new_n4671_;
  assign new_n4673_ = new_n4666_ & new_n4672_;
  assign new_n4674_ = new_n4658_ & new_n4673_;
  assign new_n4675_ = new_n4639_ & new_n4674_;
  assign new_n4676_ = ~A267 & ~A233;
  assign new_n4677_ = new_n1133_ & new_n4676_;
  assign new_n4678_ = new_n1062_ & new_n4677_;
  assign new_n4679_ = new_n4627_ & new_n4678_;
  assign new_n4680_ = new_n1112_ & new_n4623_;
  assign new_n4681_ = new_n1062_ & new_n4680_;
  assign new_n4682_ = new_n4627_ & new_n4681_;
  assign new_n4683_ = new_n1129_ & new_n4623_;
  assign new_n4684_ = new_n1068_ & new_n4683_;
  assign new_n4685_ = new_n4627_ & new_n4684_;
  assign new_n4686_ = ~new_n4682_ & ~new_n4685_;
  assign new_n4687_ = ~new_n4679_ & new_n4686_;
  assign new_n4688_ = new_n1147_ & new_n4676_;
  assign new_n4689_ = new_n1068_ & new_n4688_;
  assign new_n4690_ = new_n4627_ & new_n4689_;
  assign new_n4691_ = new_n1124_ & new_n4676_;
  assign new_n4692_ = new_n1068_ & new_n4691_;
  assign new_n4693_ = new_n4627_ & new_n4692_;
  assign new_n4694_ = new_n1143_ & new_n4676_;
  assign new_n4695_ = new_n1062_ & new_n4694_;
  assign new_n4696_ = new_n4627_ & new_n4695_;
  assign new_n4697_ = ~new_n4693_ & ~new_n4696_;
  assign new_n4698_ = ~new_n4690_ & new_n4697_;
  assign new_n4699_ = new_n4687_ & new_n4698_;
  assign new_n4700_ = A267 & ~A233;
  assign new_n4701_ = new_n31_ & new_n4700_;
  assign new_n4702_ = new_n947_ & new_n4701_;
  assign new_n4703_ = new_n4627_ & new_n4702_;
  assign new_n4704_ = new_n950_ & new_n4701_;
  assign new_n4705_ = new_n4627_ & new_n4704_;
  assign new_n4706_ = new_n953_ & new_n4701_;
  assign new_n4707_ = new_n4627_ & new_n4706_;
  assign new_n4708_ = ~new_n4705_ & ~new_n4707_;
  assign new_n4709_ = ~new_n4703_ & new_n4708_;
  assign new_n4710_ = ~A265 & A233;
  assign new_n4711_ = new_n1069_ & new_n4710_;
  assign new_n4712_ = new_n1068_ & new_n4711_;
  assign new_n4713_ = new_n96_ & new_n1908_;
  assign new_n4714_ = new_n4255_ & new_n4713_;
  assign new_n4715_ = new_n4712_ & new_n4714_;
  assign new_n4716_ = new_n963_ & new_n4701_;
  assign new_n4717_ = new_n4627_ & new_n4716_;
  assign new_n4718_ = new_n1063_ & new_n4710_;
  assign new_n4719_ = new_n1062_ & new_n4718_;
  assign new_n4720_ = new_n4714_ & new_n4719_;
  assign new_n4721_ = ~new_n4717_ & ~new_n4720_;
  assign new_n4722_ = ~new_n4715_ & new_n4721_;
  assign new_n4723_ = new_n4709_ & new_n4722_;
  assign new_n4724_ = new_n4699_ & new_n4723_;
  assign new_n4725_ = A265 & A233;
  assign new_n4726_ = new_n46_ & new_n4725_;
  assign new_n4727_ = new_n1081_ & new_n4726_;
  assign new_n4728_ = new_n4714_ & new_n4727_;
  assign new_n4729_ = new_n1058_ & new_n4726_;
  assign new_n4730_ = new_n4714_ & new_n4729_;
  assign new_n4731_ = new_n1078_ & new_n4726_;
  assign new_n4732_ = new_n4714_ & new_n4731_;
  assign new_n4733_ = ~new_n4730_ & ~new_n4732_;
  assign new_n4734_ = ~new_n4728_ & new_n4733_;
  assign new_n4735_ = new_n1093_ & new_n4725_;
  assign new_n4736_ = new_n1098_ & new_n4735_;
  assign new_n4737_ = new_n4714_ & new_n4736_;
  assign new_n4738_ = new_n1075_ & new_n4726_;
  assign new_n4739_ = new_n4714_ & new_n4738_;
  assign new_n4740_ = new_n1092_ & new_n4735_;
  assign new_n4741_ = new_n4714_ & new_n4740_;
  assign new_n4742_ = ~new_n4739_ & ~new_n4741_;
  assign new_n4743_ = ~new_n4737_ & new_n4742_;
  assign new_n4744_ = new_n4734_ & new_n4743_;
  assign new_n4745_ = new_n51_ & new_n4710_;
  assign new_n4746_ = new_n1081_ & new_n4745_;
  assign new_n4747_ = new_n4714_ & new_n4746_;
  assign new_n4748_ = new_n1058_ & new_n4745_;
  assign new_n4749_ = new_n4714_ & new_n4748_;
  assign new_n4750_ = new_n1078_ & new_n4745_;
  assign new_n4751_ = new_n4714_ & new_n4750_;
  assign new_n4752_ = ~new_n4749_ & ~new_n4751_;
  assign new_n4753_ = ~new_n4747_ & new_n4752_;
  assign new_n4754_ = new_n1075_ & new_n4745_;
  assign new_n4755_ = new_n4714_ & new_n4754_;
  assign new_n4756_ = new_n1116_ & new_n4710_;
  assign new_n4757_ = new_n1092_ & new_n4756_;
  assign new_n4758_ = new_n4714_ & new_n4757_;
  assign new_n4759_ = ~new_n4755_ & ~new_n4758_;
  assign new_n4760_ = new_n4753_ & new_n4759_;
  assign new_n4761_ = new_n4744_ & new_n4760_;
  assign new_n4762_ = new_n4724_ & new_n4761_;
  assign new_n4763_ = new_n4675_ & new_n4762_;
  assign new_n4764_ = new_n4606_ & new_n4763_;
  assign new_n4765_ = new_n4504_ & new_n4764_;
  assign new_n4766_ = new_n1129_ & new_n4725_;
  assign new_n4767_ = new_n1068_ & new_n4766_;
  assign new_n4768_ = new_n4714_ & new_n4767_;
  assign new_n4769_ = new_n1098_ & new_n4756_;
  assign new_n4770_ = new_n4714_ & new_n4769_;
  assign new_n4771_ = new_n1112_ & new_n4725_;
  assign new_n4772_ = new_n1062_ & new_n4771_;
  assign new_n4773_ = new_n4714_ & new_n4772_;
  assign new_n4774_ = ~new_n4770_ & ~new_n4773_;
  assign new_n4775_ = ~new_n4768_ & new_n4774_;
  assign new_n4776_ = ~A267 & A233;
  assign new_n4777_ = new_n1143_ & new_n4776_;
  assign new_n4778_ = new_n1062_ & new_n4777_;
  assign new_n4779_ = new_n4714_ & new_n4778_;
  assign new_n4780_ = new_n1133_ & new_n4776_;
  assign new_n4781_ = new_n1062_ & new_n4780_;
  assign new_n4782_ = new_n4714_ & new_n4781_;
  assign new_n4783_ = new_n1124_ & new_n4776_;
  assign new_n4784_ = new_n1068_ & new_n4783_;
  assign new_n4785_ = new_n4714_ & new_n4784_;
  assign new_n4786_ = ~new_n4782_ & ~new_n4785_;
  assign new_n4787_ = ~new_n4779_ & new_n4786_;
  assign new_n4788_ = new_n4775_ & new_n4787_;
  assign new_n4789_ = A267 & A233;
  assign new_n4790_ = new_n31_ & new_n4789_;
  assign new_n4791_ = new_n953_ & new_n4790_;
  assign new_n4792_ = new_n4714_ & new_n4791_;
  assign new_n4793_ = new_n1147_ & new_n4776_;
  assign new_n4794_ = new_n1068_ & new_n4793_;
  assign new_n4795_ = new_n4714_ & new_n4794_;
  assign new_n4796_ = new_n950_ & new_n4790_;
  assign new_n4797_ = new_n4714_ & new_n4796_;
  assign new_n4798_ = ~new_n4795_ & ~new_n4797_;
  assign new_n4799_ = ~new_n4792_ & new_n4798_;
  assign new_n4800_ = ~A234 & A203;
  assign new_n4801_ = new_n1908_ & new_n4800_;
  assign new_n4802_ = new_n4255_ & new_n4801_;
  assign new_n4803_ = new_n1065_ & new_n4802_;
  assign new_n4804_ = new_n947_ & new_n4790_;
  assign new_n4805_ = new_n4714_ & new_n4804_;
  assign new_n4806_ = new_n963_ & new_n4790_;
  assign new_n4807_ = new_n4714_ & new_n4806_;
  assign new_n4808_ = ~new_n4805_ & ~new_n4807_;
  assign new_n4809_ = ~new_n4803_ & new_n4808_;
  assign new_n4810_ = new_n4799_ & new_n4809_;
  assign new_n4811_ = new_n4788_ & new_n4810_;
  assign new_n4812_ = new_n1079_ & new_n4802_;
  assign new_n4813_ = new_n1071_ & new_n4802_;
  assign new_n4814_ = new_n1059_ & new_n4802_;
  assign new_n4815_ = ~new_n4813_ & ~new_n4814_;
  assign new_n4816_ = ~new_n4812_ & new_n4815_;
  assign new_n4817_ = new_n1095_ & new_n4802_;
  assign new_n4818_ = new_n1082_ & new_n4802_;
  assign new_n4819_ = new_n1076_ & new_n4802_;
  assign new_n4820_ = ~new_n4818_ & ~new_n4819_;
  assign new_n4821_ = ~new_n4817_ & new_n4820_;
  assign new_n4822_ = new_n4816_ & new_n4821_;
  assign new_n4823_ = new_n1105_ & new_n4802_;
  assign new_n4824_ = new_n1099_ & new_n4802_;
  assign new_n4825_ = new_n1089_ & new_n4802_;
  assign new_n4826_ = ~new_n4824_ & ~new_n4825_;
  assign new_n4827_ = ~new_n4823_ & new_n4826_;
  assign new_n4828_ = new_n1107_ & new_n4802_;
  assign new_n4829_ = new_n1103_ & new_n4802_;
  assign new_n4830_ = ~new_n4828_ & ~new_n4829_;
  assign new_n4831_ = new_n4827_ & new_n4830_;
  assign new_n4832_ = new_n4822_ & new_n4831_;
  assign new_n4833_ = new_n4811_ & new_n4832_;
  assign new_n4834_ = new_n1114_ & new_n4802_;
  assign new_n4835_ = new_n1118_ & new_n4802_;
  assign new_n4836_ = new_n1120_ & new_n4802_;
  assign new_n4837_ = ~new_n4835_ & ~new_n4836_;
  assign new_n4838_ = ~new_n4834_ & new_n4837_;
  assign new_n4839_ = new_n1127_ & new_n4802_;
  assign new_n4840_ = new_n1131_ & new_n4802_;
  assign new_n4841_ = new_n1135_ & new_n4802_;
  assign new_n4842_ = ~new_n4840_ & ~new_n4841_;
  assign new_n4843_ = ~new_n4839_ & new_n4842_;
  assign new_n4844_ = new_n4838_ & new_n4843_;
  assign new_n4845_ = new_n1141_ & new_n4802_;
  assign new_n4846_ = new_n1145_ & new_n4802_;
  assign new_n4847_ = new_n1149_ & new_n4802_;
  assign new_n4848_ = ~new_n4846_ & ~new_n4847_;
  assign new_n4849_ = ~new_n4845_ & new_n4848_;
  assign new_n4850_ = new_n1153_ & new_n4802_;
  assign new_n4851_ = new_n1155_ & new_n4802_;
  assign new_n4852_ = new_n1157_ & new_n4802_;
  assign new_n4853_ = ~new_n4851_ & ~new_n4852_;
  assign new_n4854_ = ~new_n4850_ & new_n4853_;
  assign new_n4855_ = new_n4849_ & new_n4854_;
  assign new_n4856_ = new_n4844_ & new_n4855_;
  assign new_n4857_ = new_n1162_ & new_n4802_;
  assign new_n4858_ = new_n1165_ & new_n4802_;
  assign new_n4859_ = new_n1168_ & new_n4802_;
  assign new_n4860_ = ~new_n4858_ & ~new_n4859_;
  assign new_n4861_ = ~new_n4857_ & new_n4860_;
  assign new_n4862_ = new_n1184_ & new_n4802_;
  assign new_n4863_ = new_n1172_ & new_n4802_;
  assign new_n4864_ = new_n1174_ & new_n4802_;
  assign new_n4865_ = ~new_n4863_ & ~new_n4864_;
  assign new_n4866_ = ~new_n4862_ & new_n4865_;
  assign new_n4867_ = new_n4861_ & new_n4866_;
  assign new_n4868_ = new_n1192_ & new_n4802_;
  assign new_n4869_ = new_n1186_ & new_n4802_;
  assign new_n4870_ = new_n1182_ & new_n4802_;
  assign new_n4871_ = ~new_n4869_ & ~new_n4870_;
  assign new_n4872_ = ~new_n4868_ & new_n4871_;
  assign new_n4873_ = new_n1194_ & new_n4802_;
  assign new_n4874_ = new_n1190_ & new_n4802_;
  assign new_n4875_ = ~new_n4873_ & ~new_n4874_;
  assign new_n4876_ = new_n4872_ & new_n4875_;
  assign new_n4877_ = new_n4867_ & new_n4876_;
  assign new_n4878_ = new_n4856_ & new_n4877_;
  assign new_n4879_ = new_n4833_ & new_n4878_;
  assign new_n4880_ = new_n1200_ & new_n4802_;
  assign new_n4881_ = new_n1202_ & new_n4802_;
  assign new_n4882_ = new_n1204_ & new_n4802_;
  assign new_n4883_ = ~new_n4881_ & ~new_n4882_;
  assign new_n4884_ = ~new_n4880_ & new_n4883_;
  assign new_n4885_ = new_n1210_ & new_n4802_;
  assign new_n4886_ = new_n1213_ & new_n4802_;
  assign new_n4887_ = new_n1216_ & new_n4802_;
  assign new_n4888_ = ~new_n4886_ & ~new_n4887_;
  assign new_n4889_ = ~new_n4885_ & new_n4888_;
  assign new_n4890_ = new_n4884_ & new_n4889_;
  assign new_n4891_ = new_n1223_ & new_n4802_;
  assign new_n4892_ = new_n1226_ & new_n4802_;
  assign new_n4893_ = new_n1229_ & new_n4802_;
  assign new_n4894_ = ~new_n4892_ & ~new_n4893_;
  assign new_n4895_ = ~new_n4891_ & new_n4894_;
  assign new_n4896_ = new_n1233_ & new_n4802_;
  assign new_n4897_ = new_n1235_ & new_n4802_;
  assign new_n4898_ = new_n1237_ & new_n4802_;
  assign new_n4899_ = ~new_n4897_ & ~new_n4898_;
  assign new_n4900_ = ~new_n4896_ & new_n4899_;
  assign new_n4901_ = new_n4895_ & new_n4900_;
  assign new_n4902_ = new_n4890_ & new_n4901_;
  assign new_n4903_ = new_n1906_ & new_n1908_;
  assign new_n4904_ = new_n4255_ & new_n4903_;
  assign new_n4905_ = new_n954_ & new_n4904_;
  assign new_n4906_ = new_n1243_ & new_n4802_;
  assign new_n4907_ = new_n951_ & new_n4904_;
  assign new_n4908_ = ~new_n4906_ & ~new_n4907_;
  assign new_n4909_ = ~new_n4905_ & new_n4908_;
  assign new_n4910_ = new_n967_ & new_n4904_;
  assign new_n4911_ = new_n948_ & new_n4904_;
  assign new_n4912_ = new_n964_ & new_n4904_;
  assign new_n4913_ = ~new_n4911_ & ~new_n4912_;
  assign new_n4914_ = ~new_n4910_ & new_n4913_;
  assign new_n4915_ = new_n4909_ & new_n4914_;
  assign new_n4916_ = new_n978_ & new_n4904_;
  assign new_n4917_ = new_n961_ & new_n4904_;
  assign new_n4918_ = new_n975_ & new_n4904_;
  assign new_n4919_ = ~new_n4917_ & ~new_n4918_;
  assign new_n4920_ = ~new_n4916_ & new_n4919_;
  assign new_n4921_ = new_n972_ & new_n4904_;
  assign new_n4922_ = new_n987_ & new_n4904_;
  assign new_n4923_ = ~new_n4921_ & ~new_n4922_;
  assign new_n4924_ = new_n4920_ & new_n4923_;
  assign new_n4925_ = new_n4915_ & new_n4924_;
  assign new_n4926_ = new_n4902_ & new_n4925_;
  assign new_n4927_ = new_n994_ & new_n4904_;
  assign new_n4928_ = new_n990_ & new_n4904_;
  assign new_n4929_ = new_n984_ & new_n4904_;
  assign new_n4930_ = ~new_n4928_ & ~new_n4929_;
  assign new_n4931_ = ~new_n4927_ & new_n4930_;
  assign new_n4932_ = new_n1010_ & new_n4904_;
  assign new_n4933_ = new_n996_ & new_n4904_;
  assign new_n4934_ = new_n1008_ & new_n4904_;
  assign new_n4935_ = ~new_n4933_ & ~new_n4934_;
  assign new_n4936_ = ~new_n4932_ & new_n4935_;
  assign new_n4937_ = new_n4931_ & new_n4936_;
  assign new_n4938_ = new_n1018_ & new_n4904_;
  assign new_n4939_ = new_n1006_ & new_n4904_;
  assign new_n4940_ = new_n1016_ & new_n4904_;
  assign new_n4941_ = ~new_n4939_ & ~new_n4940_;
  assign new_n4942_ = ~new_n4938_ & new_n4941_;
  assign new_n4943_ = new_n1027_ & new_n4904_;
  assign new_n4944_ = new_n1014_ & new_n4904_;
  assign new_n4945_ = new_n1025_ & new_n4904_;
  assign new_n4946_ = ~new_n4944_ & ~new_n4945_;
  assign new_n4947_ = ~new_n4943_ & new_n4946_;
  assign new_n4948_ = new_n4942_ & new_n4947_;
  assign new_n4949_ = new_n4937_ & new_n4948_;
  assign new_n4950_ = new_n1035_ & new_n4904_;
  assign new_n4951_ = new_n1023_ & new_n4904_;
  assign new_n4952_ = new_n1033_ & new_n4904_;
  assign new_n4953_ = ~new_n4951_ & ~new_n4952_;
  assign new_n4954_ = ~new_n4950_ & new_n4953_;
  assign new_n4955_ = new_n1045_ & new_n4904_;
  assign new_n4956_ = new_n1031_ & new_n4904_;
  assign new_n4957_ = new_n1043_ & new_n4904_;
  assign new_n4958_ = ~new_n4956_ & ~new_n4957_;
  assign new_n4959_ = ~new_n4955_ & new_n4958_;
  assign new_n4960_ = new_n4954_ & new_n4959_;
  assign new_n4961_ = new_n1053_ & new_n4904_;
  assign new_n4962_ = new_n1041_ & new_n4904_;
  assign new_n4963_ = new_n1051_ & new_n4904_;
  assign new_n4964_ = ~new_n4962_ & ~new_n4963_;
  assign new_n4965_ = ~new_n4961_ & new_n4964_;
  assign new_n4966_ = new_n1049_ & new_n4904_;
  assign new_n4967_ = ~A199 & ~A168;
  assign new_n4968_ = A169 & new_n4967_;
  assign new_n4969_ = new_n1727_ & new_n4968_;
  assign new_n4970_ = new_n1735_ & new_n4969_;
  assign new_n4971_ = ~new_n4966_ & ~new_n4970_;
  assign new_n4972_ = new_n4965_ & new_n4971_;
  assign new_n4973_ = new_n4960_ & new_n4972_;
  assign new_n4974_ = new_n4949_ & new_n4973_;
  assign new_n4975_ = new_n4926_ & new_n4974_;
  assign new_n4976_ = new_n4879_ & new_n4975_;
  assign new_n4977_ = new_n1749_ & new_n4969_;
  assign new_n4978_ = new_n1738_ & new_n4969_;
  assign new_n4979_ = new_n1725_ & new_n4969_;
  assign new_n4980_ = ~new_n4978_ & ~new_n4979_;
  assign new_n4981_ = ~new_n4977_ & new_n4980_;
  assign new_n4982_ = A199 & ~A168;
  assign new_n4983_ = A169 & new_n4982_;
  assign new_n4984_ = new_n1743_ & new_n4983_;
  assign new_n4985_ = new_n1725_ & new_n4984_;
  assign new_n4986_ = new_n1735_ & new_n4984_;
  assign new_n4987_ = new_n1738_ & new_n4984_;
  assign new_n4988_ = ~new_n4986_ & ~new_n4987_;
  assign new_n4989_ = ~new_n4985_ & new_n4988_;
  assign new_n4990_ = new_n4981_ & new_n4989_;
  assign new_n4991_ = ~A201 & ~A168;
  assign new_n4992_ = A169 & new_n4991_;
  assign new_n4993_ = new_n1757_ & new_n4992_;
  assign new_n4994_ = new_n1738_ & new_n4993_;
  assign new_n4995_ = new_n1749_ & new_n4984_;
  assign new_n4996_ = new_n1735_ & new_n4993_;
  assign new_n4997_ = ~new_n4995_ & ~new_n4996_;
  assign new_n4998_ = ~new_n4994_ & new_n4997_;
  assign new_n4999_ = new_n1773_ & new_n4992_;
  assign new_n5000_ = new_n1735_ & new_n4999_;
  assign new_n5001_ = new_n1725_ & new_n4993_;
  assign new_n5002_ = new_n1749_ & new_n4993_;
  assign new_n5003_ = ~new_n5001_ & ~new_n5002_;
  assign new_n5004_ = ~new_n5000_ & new_n5003_;
  assign new_n5005_ = new_n4998_ & new_n5004_;
  assign new_n5006_ = new_n4990_ & new_n5005_;
  assign new_n5007_ = new_n1749_ & new_n4999_;
  assign new_n5008_ = new_n1738_ & new_n4999_;
  assign new_n5009_ = new_n1725_ & new_n4999_;
  assign new_n5010_ = ~new_n5008_ & ~new_n5009_;
  assign new_n5011_ = ~new_n5007_ & new_n5010_;
  assign new_n5012_ = A201 & ~A168;
  assign new_n5013_ = A169 & new_n5012_;
  assign new_n5014_ = new_n1782_ & new_n5013_;
  assign new_n5015_ = new_n1725_ & new_n5014_;
  assign new_n5016_ = new_n1735_ & new_n5014_;
  assign new_n5017_ = new_n1738_ & new_n5014_;
  assign new_n5018_ = ~new_n5016_ & ~new_n5017_;
  assign new_n5019_ = ~new_n5015_ & new_n5018_;
  assign new_n5020_ = new_n5011_ & new_n5019_;
  assign new_n5021_ = new_n1796_ & new_n5013_;
  assign new_n5022_ = new_n1738_ & new_n5021_;
  assign new_n5023_ = new_n1749_ & new_n5014_;
  assign new_n5024_ = new_n1735_ & new_n5021_;
  assign new_n5025_ = ~new_n5023_ & ~new_n5024_;
  assign new_n5026_ = ~new_n5022_ & new_n5025_;
  assign new_n5027_ = new_n1725_ & new_n5021_;
  assign new_n5028_ = new_n1749_ & new_n5021_;
  assign new_n5029_ = ~new_n5027_ & ~new_n5028_;
  assign new_n5030_ = new_n5026_ & new_n5029_;
  assign new_n5031_ = new_n5020_ & new_n5030_;
  assign new_n5032_ = new_n5006_ & new_n5031_;
  assign new_n5033_ = new_n1805_ & new_n5013_;
  assign new_n5034_ = new_n1725_ & new_n5033_;
  assign new_n5035_ = new_n1735_ & new_n5033_;
  assign new_n5036_ = new_n1738_ & new_n5033_;
  assign new_n5037_ = ~new_n5035_ & ~new_n5036_;
  assign new_n5038_ = ~new_n5034_ & new_n5037_;
  assign new_n5039_ = new_n1813_ & new_n5013_;
  assign new_n5040_ = new_n1738_ & new_n5039_;
  assign new_n5041_ = new_n1749_ & new_n5033_;
  assign new_n5042_ = new_n1735_ & new_n5039_;
  assign new_n5043_ = ~new_n5041_ & ~new_n5042_;
  assign new_n5044_ = ~new_n5040_ & new_n5043_;
  assign new_n5045_ = new_n5038_ & new_n5044_;
  assign new_n5046_ = new_n506_ & new_n5013_;
  assign new_n5047_ = new_n1830_ & new_n5046_;
  assign new_n5048_ = new_n1725_ & new_n5039_;
  assign new_n5049_ = new_n1749_ & new_n5039_;
  assign new_n5050_ = ~new_n5048_ & ~new_n5049_;
  assign new_n5051_ = ~new_n5047_ & new_n5050_;
  assign new_n5052_ = new_n1840_ & new_n5046_;
  assign new_n5053_ = new_n1833_ & new_n5046_;
  assign new_n5054_ = new_n1827_ & new_n5046_;
  assign new_n5055_ = ~new_n5053_ & ~new_n5054_;
  assign new_n5056_ = ~new_n5052_ & new_n5055_;
  assign new_n5057_ = new_n5051_ & new_n5056_;
  assign new_n5058_ = new_n5045_ & new_n5057_;
  assign new_n5059_ = new_n1847_ & new_n5046_;
  assign new_n5060_ = new_n1842_ & new_n5046_;
  assign new_n5061_ = new_n1838_ & new_n5046_;
  assign new_n5062_ = ~new_n5060_ & ~new_n5061_;
  assign new_n5063_ = ~new_n5059_ & new_n5062_;
  assign new_n5064_ = new_n1859_ & new_n5046_;
  assign new_n5065_ = new_n1849_ & new_n5046_;
  assign new_n5066_ = new_n1857_ & new_n5046_;
  assign new_n5067_ = ~new_n5065_ & ~new_n5066_;
  assign new_n5068_ = ~new_n5064_ & new_n5067_;
  assign new_n5069_ = new_n5063_ & new_n5068_;
  assign new_n5070_ = new_n1868_ & new_n5046_;
  assign new_n5071_ = new_n1855_ & new_n5046_;
  assign new_n5072_ = new_n1866_ & new_n5046_;
  assign new_n5073_ = ~new_n5071_ & ~new_n5072_;
  assign new_n5074_ = ~new_n5070_ & new_n5073_;
  assign new_n5075_ = new_n1864_ & new_n5046_;
  assign new_n5076_ = new_n1878_ & new_n5046_;
  assign new_n5077_ = ~new_n5075_ & ~new_n5076_;
  assign new_n5078_ = new_n5074_ & new_n5077_;
  assign new_n5079_ = new_n5069_ & new_n5078_;
  assign new_n5080_ = new_n5058_ & new_n5079_;
  assign new_n5081_ = new_n5032_ & new_n5080_;
  assign new_n5082_ = new_n1889_ & new_n5046_;
  assign new_n5083_ = new_n1881_ & new_n5046_;
  assign new_n5084_ = new_n1875_ & new_n5046_;
  assign new_n5085_ = ~new_n5083_ & ~new_n5084_;
  assign new_n5086_ = ~new_n5082_ & new_n5085_;
  assign new_n5087_ = new_n1900_ & new_n5046_;
  assign new_n5088_ = new_n1892_ & new_n5046_;
  assign new_n5089_ = new_n1886_ & new_n5046_;
  assign new_n5090_ = ~new_n5088_ & ~new_n5089_;
  assign new_n5091_ = ~new_n5087_ & new_n5090_;
  assign new_n5092_ = new_n5086_ & new_n5091_;
  assign new_n5093_ = new_n1913_ & new_n5046_;
  assign new_n5094_ = new_n1902_ & new_n5046_;
  assign new_n5095_ = new_n1898_ & new_n5046_;
  assign new_n5096_ = ~new_n5094_ & ~new_n5095_;
  assign new_n5097_ = ~new_n5093_ & new_n5096_;
  assign new_n5098_ = ~A167 & A168;
  assign new_n5099_ = A169 & new_n5098_;
  assign new_n5100_ = new_n144_ & new_n5099_;
  assign new_n5101_ = new_n948_ & new_n5100_;
  assign new_n5102_ = new_n951_ & new_n5100_;
  assign new_n5103_ = new_n954_ & new_n5100_;
  assign new_n5104_ = ~new_n5102_ & ~new_n5103_;
  assign new_n5105_ = ~new_n5101_ & new_n5104_;
  assign new_n5106_ = new_n5097_ & new_n5105_;
  assign new_n5107_ = new_n5092_ & new_n5106_;
  assign new_n5108_ = new_n961_ & new_n5100_;
  assign new_n5109_ = new_n964_ & new_n5100_;
  assign new_n5110_ = new_n967_ & new_n5100_;
  assign new_n5111_ = ~new_n5109_ & ~new_n5110_;
  assign new_n5112_ = ~new_n5108_ & new_n5111_;
  assign new_n5113_ = new_n972_ & new_n5100_;
  assign new_n5114_ = new_n975_ & new_n5100_;
  assign new_n5115_ = new_n978_ & new_n5100_;
  assign new_n5116_ = ~new_n5114_ & ~new_n5115_;
  assign new_n5117_ = ~new_n5113_ & new_n5116_;
  assign new_n5118_ = new_n5112_ & new_n5117_;
  assign new_n5119_ = new_n984_ & new_n5100_;
  assign new_n5120_ = new_n987_ & new_n5100_;
  assign new_n5121_ = new_n990_ & new_n5100_;
  assign new_n5122_ = ~new_n5120_ & ~new_n5121_;
  assign new_n5123_ = ~new_n5119_ & new_n5122_;
  assign new_n5124_ = new_n994_ & new_n5100_;
  assign new_n5125_ = new_n996_ & new_n5100_;
  assign new_n5126_ = ~new_n5124_ & ~new_n5125_;
  assign new_n5127_ = new_n5123_ & new_n5126_;
  assign new_n5128_ = new_n5118_ & new_n5127_;
  assign new_n5129_ = new_n5107_ & new_n5128_;
  assign new_n5130_ = new_n1006_ & new_n5100_;
  assign new_n5131_ = new_n1008_ & new_n5100_;
  assign new_n5132_ = new_n1010_ & new_n5100_;
  assign new_n5133_ = ~new_n5131_ & ~new_n5132_;
  assign new_n5134_ = ~new_n5130_ & new_n5133_;
  assign new_n5135_ = new_n1014_ & new_n5100_;
  assign new_n5136_ = new_n1016_ & new_n5100_;
  assign new_n5137_ = new_n1018_ & new_n5100_;
  assign new_n5138_ = ~new_n5136_ & ~new_n5137_;
  assign new_n5139_ = ~new_n5135_ & new_n5138_;
  assign new_n5140_ = new_n5134_ & new_n5139_;
  assign new_n5141_ = new_n1023_ & new_n5100_;
  assign new_n5142_ = new_n1025_ & new_n5100_;
  assign new_n5143_ = new_n1027_ & new_n5100_;
  assign new_n5144_ = ~new_n5142_ & ~new_n5143_;
  assign new_n5145_ = ~new_n5141_ & new_n5144_;
  assign new_n5146_ = new_n1031_ & new_n5100_;
  assign new_n5147_ = new_n1033_ & new_n5100_;
  assign new_n5148_ = new_n1035_ & new_n5100_;
  assign new_n5149_ = ~new_n5147_ & ~new_n5148_;
  assign new_n5150_ = ~new_n5146_ & new_n5149_;
  assign new_n5151_ = new_n5145_ & new_n5150_;
  assign new_n5152_ = new_n5140_ & new_n5151_;
  assign new_n5153_ = new_n1041_ & new_n5100_;
  assign new_n5154_ = new_n1043_ & new_n5100_;
  assign new_n5155_ = new_n1045_ & new_n5100_;
  assign new_n5156_ = ~new_n5154_ & ~new_n5155_;
  assign new_n5157_ = ~new_n5153_ & new_n5156_;
  assign new_n5158_ = new_n1049_ & new_n5100_;
  assign new_n5159_ = new_n1051_ & new_n5100_;
  assign new_n5160_ = new_n1053_ & new_n5100_;
  assign new_n5161_ = ~new_n5159_ & ~new_n5160_;
  assign new_n5162_ = ~new_n5158_ & new_n5161_;
  assign new_n5163_ = new_n5157_ & new_n5162_;
  assign new_n5164_ = new_n265_ & new_n5099_;
  assign new_n5165_ = new_n1059_ & new_n5164_;
  assign new_n5166_ = new_n1065_ & new_n5164_;
  assign new_n5167_ = new_n1071_ & new_n5164_;
  assign new_n5168_ = ~new_n5166_ & ~new_n5167_;
  assign new_n5169_ = ~new_n5165_ & new_n5168_;
  assign new_n5170_ = new_n1079_ & new_n5164_;
  assign new_n5171_ = new_n1082_ & new_n5164_;
  assign new_n5172_ = ~new_n5170_ & ~new_n5171_;
  assign new_n5173_ = new_n5169_ & new_n5172_;
  assign new_n5174_ = new_n5163_ & new_n5173_;
  assign new_n5175_ = new_n5152_ & new_n5174_;
  assign new_n5176_ = new_n5129_ & new_n5175_;
  assign new_n5177_ = new_n5081_ & new_n5176_;
  assign new_n5178_ = new_n4976_ & new_n5177_;
  assign new_n5179_ = new_n4765_ & new_n5178_;
  assign new_n5180_ = new_n4293_ & new_n5179_;
  assign new_n5181_ = new_n1099_ & new_n5164_;
  assign new_n5182_ = new_n1076_ & new_n5164_;
  assign new_n5183_ = new_n1095_ & new_n5164_;
  assign new_n5184_ = ~new_n5182_ & ~new_n5183_;
  assign new_n5185_ = ~new_n5181_ & new_n5184_;
  assign new_n5186_ = new_n1107_ & new_n5164_;
  assign new_n5187_ = new_n1089_ & new_n5164_;
  assign new_n5188_ = new_n1105_ & new_n5164_;
  assign new_n5189_ = ~new_n5187_ & ~new_n5188_;
  assign new_n5190_ = ~new_n5186_ & new_n5189_;
  assign new_n5191_ = new_n5185_ & new_n5190_;
  assign new_n5192_ = new_n1120_ & new_n5164_;
  assign new_n5193_ = new_n1103_ & new_n5164_;
  assign new_n5194_ = new_n1118_ & new_n5164_;
  assign new_n5195_ = ~new_n5193_ & ~new_n5194_;
  assign new_n5196_ = ~new_n5192_ & new_n5195_;
  assign new_n5197_ = new_n1135_ & new_n5164_;
  assign new_n5198_ = new_n1114_ & new_n5164_;
  assign new_n5199_ = new_n1131_ & new_n5164_;
  assign new_n5200_ = ~new_n5198_ & ~new_n5199_;
  assign new_n5201_ = ~new_n5197_ & new_n5200_;
  assign new_n5202_ = new_n5196_ & new_n5201_;
  assign new_n5203_ = new_n5191_ & new_n5202_;
  assign new_n5204_ = new_n1149_ & new_n5164_;
  assign new_n5205_ = new_n1127_ & new_n5164_;
  assign new_n5206_ = new_n1145_ & new_n5164_;
  assign new_n5207_ = ~new_n5205_ & ~new_n5206_;
  assign new_n5208_ = ~new_n5204_ & new_n5207_;
  assign new_n5209_ = new_n1157_ & new_n5164_;
  assign new_n5210_ = new_n1141_ & new_n5164_;
  assign new_n5211_ = new_n1155_ & new_n5164_;
  assign new_n5212_ = ~new_n5210_ & ~new_n5211_;
  assign new_n5213_ = ~new_n5209_ & new_n5212_;
  assign new_n5214_ = new_n5208_ & new_n5213_;
  assign new_n5215_ = new_n1168_ & new_n5164_;
  assign new_n5216_ = new_n1153_ & new_n5164_;
  assign new_n5217_ = new_n1165_ & new_n5164_;
  assign new_n5218_ = ~new_n5216_ & ~new_n5217_;
  assign new_n5219_ = ~new_n5215_ & new_n5218_;
  assign new_n5220_ = new_n1174_ & new_n5164_;
  assign new_n5221_ = new_n1162_ & new_n5164_;
  assign new_n5222_ = new_n1172_ & new_n5164_;
  assign new_n5223_ = ~new_n5221_ & ~new_n5222_;
  assign new_n5224_ = ~new_n5220_ & new_n5223_;
  assign new_n5225_ = new_n5219_ & new_n5224_;
  assign new_n5226_ = new_n5214_ & new_n5225_;
  assign new_n5227_ = new_n5203_ & new_n5226_;
  assign new_n5228_ = new_n1182_ & new_n5164_;
  assign new_n5229_ = new_n1184_ & new_n5164_;
  assign new_n5230_ = new_n1186_ & new_n5164_;
  assign new_n5231_ = ~new_n5229_ & ~new_n5230_;
  assign new_n5232_ = ~new_n5228_ & new_n5231_;
  assign new_n5233_ = new_n1190_ & new_n5164_;
  assign new_n5234_ = new_n1192_ & new_n5164_;
  assign new_n5235_ = new_n1194_ & new_n5164_;
  assign new_n5236_ = ~new_n5234_ & ~new_n5235_;
  assign new_n5237_ = ~new_n5233_ & new_n5236_;
  assign new_n5238_ = new_n5232_ & new_n5237_;
  assign new_n5239_ = new_n1200_ & new_n5164_;
  assign new_n5240_ = new_n1202_ & new_n5164_;
  assign new_n5241_ = new_n1204_ & new_n5164_;
  assign new_n5242_ = ~new_n5240_ & ~new_n5241_;
  assign new_n5243_ = ~new_n5239_ & new_n5242_;
  assign new_n5244_ = new_n1210_ & new_n5164_;
  assign new_n5245_ = new_n1213_ & new_n5164_;
  assign new_n5246_ = new_n1216_ & new_n5164_;
  assign new_n5247_ = ~new_n5245_ & ~new_n5246_;
  assign new_n5248_ = ~new_n5244_ & new_n5247_;
  assign new_n5249_ = new_n5243_ & new_n5248_;
  assign new_n5250_ = new_n5238_ & new_n5249_;
  assign new_n5251_ = new_n1223_ & new_n5164_;
  assign new_n5252_ = new_n1226_ & new_n5164_;
  assign new_n5253_ = new_n1229_ & new_n5164_;
  assign new_n5254_ = ~new_n5252_ & ~new_n5253_;
  assign new_n5255_ = ~new_n5251_ & new_n5254_;
  assign new_n5256_ = new_n1233_ & new_n5164_;
  assign new_n5257_ = new_n1235_ & new_n5164_;
  assign new_n5258_ = new_n1237_ & new_n5164_;
  assign new_n5259_ = ~new_n5257_ & ~new_n5258_;
  assign new_n5260_ = ~new_n5256_ & new_n5259_;
  assign new_n5261_ = new_n5255_ & new_n5260_;
  assign new_n5262_ = new_n293_ & new_n5099_;
  assign new_n5263_ = new_n954_ & new_n5262_;
  assign new_n5264_ = new_n1243_ & new_n5164_;
  assign new_n5265_ = new_n951_ & new_n5262_;
  assign new_n5266_ = ~new_n5264_ & ~new_n5265_;
  assign new_n5267_ = ~new_n5263_ & new_n5266_;
  assign new_n5268_ = new_n948_ & new_n5262_;
  assign new_n5269_ = new_n964_ & new_n5262_;
  assign new_n5270_ = ~new_n5268_ & ~new_n5269_;
  assign new_n5271_ = new_n5267_ & new_n5270_;
  assign new_n5272_ = new_n5261_ & new_n5271_;
  assign new_n5273_ = new_n5250_ & new_n5272_;
  assign new_n5274_ = new_n5227_ & new_n5273_;
  assign new_n5275_ = new_n975_ & new_n5262_;
  assign new_n5276_ = new_n967_ & new_n5262_;
  assign new_n5277_ = new_n961_ & new_n5262_;
  assign new_n5278_ = ~new_n5276_ & ~new_n5277_;
  assign new_n5279_ = ~new_n5275_ & new_n5278_;
  assign new_n5280_ = new_n987_ & new_n5262_;
  assign new_n5281_ = new_n978_ & new_n5262_;
  assign new_n5282_ = new_n972_ & new_n5262_;
  assign new_n5283_ = ~new_n5281_ & ~new_n5282_;
  assign new_n5284_ = ~new_n5280_ & new_n5283_;
  assign new_n5285_ = new_n5279_ & new_n5284_;
  assign new_n5286_ = new_n994_ & new_n5262_;
  assign new_n5287_ = new_n990_ & new_n5262_;
  assign new_n5288_ = new_n984_ & new_n5262_;
  assign new_n5289_ = ~new_n5287_ & ~new_n5288_;
  assign new_n5290_ = ~new_n5286_ & new_n5289_;
  assign new_n5291_ = new_n1010_ & new_n5262_;
  assign new_n5292_ = new_n996_ & new_n5262_;
  assign new_n5293_ = new_n1008_ & new_n5262_;
  assign new_n5294_ = ~new_n5292_ & ~new_n5293_;
  assign new_n5295_ = ~new_n5291_ & new_n5294_;
  assign new_n5296_ = new_n5290_ & new_n5295_;
  assign new_n5297_ = new_n5285_ & new_n5296_;
  assign new_n5298_ = new_n1018_ & new_n5262_;
  assign new_n5299_ = new_n1006_ & new_n5262_;
  assign new_n5300_ = new_n1016_ & new_n5262_;
  assign new_n5301_ = ~new_n5299_ & ~new_n5300_;
  assign new_n5302_ = ~new_n5298_ & new_n5301_;
  assign new_n5303_ = new_n1027_ & new_n5262_;
  assign new_n5304_ = new_n1014_ & new_n5262_;
  assign new_n5305_ = new_n1025_ & new_n5262_;
  assign new_n5306_ = ~new_n5304_ & ~new_n5305_;
  assign new_n5307_ = ~new_n5303_ & new_n5306_;
  assign new_n5308_ = new_n5302_ & new_n5307_;
  assign new_n5309_ = new_n1035_ & new_n5262_;
  assign new_n5310_ = new_n1023_ & new_n5262_;
  assign new_n5311_ = new_n1033_ & new_n5262_;
  assign new_n5312_ = ~new_n5310_ & ~new_n5311_;
  assign new_n5313_ = ~new_n5309_ & new_n5312_;
  assign new_n5314_ = new_n1031_ & new_n5262_;
  assign new_n5315_ = new_n1043_ & new_n5262_;
  assign new_n5316_ = ~new_n5314_ & ~new_n5315_;
  assign new_n5317_ = new_n5313_ & new_n5316_;
  assign new_n5318_ = new_n5308_ & new_n5317_;
  assign new_n5319_ = new_n5297_ & new_n5318_;
  assign new_n5320_ = new_n1051_ & new_n5262_;
  assign new_n5321_ = new_n1045_ & new_n5262_;
  assign new_n5322_ = new_n1041_ & new_n5262_;
  assign new_n5323_ = ~new_n5321_ & ~new_n5322_;
  assign new_n5324_ = ~new_n5320_ & new_n5323_;
  assign new_n5325_ = new_n351_ & new_n5099_;
  assign new_n5326_ = new_n1065_ & new_n5325_;
  assign new_n5327_ = new_n1053_ & new_n5262_;
  assign new_n5328_ = new_n1049_ & new_n5262_;
  assign new_n5329_ = ~new_n5327_ & ~new_n5328_;
  assign new_n5330_ = ~new_n5326_ & new_n5329_;
  assign new_n5331_ = new_n5324_ & new_n5330_;
  assign new_n5332_ = new_n1079_ & new_n5325_;
  assign new_n5333_ = new_n1071_ & new_n5325_;
  assign new_n5334_ = new_n1059_ & new_n5325_;
  assign new_n5335_ = ~new_n5333_ & ~new_n5334_;
  assign new_n5336_ = ~new_n5332_ & new_n5335_;
  assign new_n5337_ = new_n1095_ & new_n5325_;
  assign new_n5338_ = new_n1082_ & new_n5325_;
  assign new_n5339_ = new_n1076_ & new_n5325_;
  assign new_n5340_ = ~new_n5338_ & ~new_n5339_;
  assign new_n5341_ = ~new_n5337_ & new_n5340_;
  assign new_n5342_ = new_n5336_ & new_n5341_;
  assign new_n5343_ = new_n5331_ & new_n5342_;
  assign new_n5344_ = new_n1105_ & new_n5325_;
  assign new_n5345_ = new_n1099_ & new_n5325_;
  assign new_n5346_ = new_n1089_ & new_n5325_;
  assign new_n5347_ = ~new_n5345_ & ~new_n5346_;
  assign new_n5348_ = ~new_n5344_ & new_n5347_;
  assign new_n5349_ = new_n1118_ & new_n5325_;
  assign new_n5350_ = new_n1107_ & new_n5325_;
  assign new_n5351_ = new_n1103_ & new_n5325_;
  assign new_n5352_ = ~new_n5350_ & ~new_n5351_;
  assign new_n5353_ = ~new_n5349_ & new_n5352_;
  assign new_n5354_ = new_n5348_ & new_n5353_;
  assign new_n5355_ = new_n1131_ & new_n5325_;
  assign new_n5356_ = new_n1120_ & new_n5325_;
  assign new_n5357_ = new_n1114_ & new_n5325_;
  assign new_n5358_ = ~new_n5356_ & ~new_n5357_;
  assign new_n5359_ = ~new_n5355_ & new_n5358_;
  assign new_n5360_ = new_n1135_ & new_n5325_;
  assign new_n5361_ = new_n1127_ & new_n5325_;
  assign new_n5362_ = ~new_n5360_ & ~new_n5361_;
  assign new_n5363_ = new_n5359_ & new_n5362_;
  assign new_n5364_ = new_n5354_ & new_n5363_;
  assign new_n5365_ = new_n5343_ & new_n5364_;
  assign new_n5366_ = new_n5319_ & new_n5365_;
  assign new_n5367_ = new_n5274_ & new_n5366_;
  assign new_n5368_ = new_n1141_ & new_n5325_;
  assign new_n5369_ = new_n1145_ & new_n5325_;
  assign new_n5370_ = new_n1149_ & new_n5325_;
  assign new_n5371_ = ~new_n5369_ & ~new_n5370_;
  assign new_n5372_ = ~new_n5368_ & new_n5371_;
  assign new_n5373_ = new_n1153_ & new_n5325_;
  assign new_n5374_ = new_n1155_ & new_n5325_;
  assign new_n5375_ = new_n1157_ & new_n5325_;
  assign new_n5376_ = ~new_n5374_ & ~new_n5375_;
  assign new_n5377_ = ~new_n5373_ & new_n5376_;
  assign new_n5378_ = new_n5372_ & new_n5377_;
  assign new_n5379_ = new_n1162_ & new_n5325_;
  assign new_n5380_ = new_n1165_ & new_n5325_;
  assign new_n5381_ = new_n1168_ & new_n5325_;
  assign new_n5382_ = ~new_n5380_ & ~new_n5381_;
  assign new_n5383_ = ~new_n5379_ & new_n5382_;
  assign new_n5384_ = new_n1184_ & new_n5325_;
  assign new_n5385_ = new_n1172_ & new_n5325_;
  assign new_n5386_ = new_n1174_ & new_n5325_;
  assign new_n5387_ = ~new_n5385_ & ~new_n5386_;
  assign new_n5388_ = ~new_n5384_ & new_n5387_;
  assign new_n5389_ = new_n5383_ & new_n5388_;
  assign new_n5390_ = new_n5378_ & new_n5389_;
  assign new_n5391_ = new_n1192_ & new_n5325_;
  assign new_n5392_ = new_n1186_ & new_n5325_;
  assign new_n5393_ = new_n1182_ & new_n5325_;
  assign new_n5394_ = ~new_n5392_ & ~new_n5393_;
  assign new_n5395_ = ~new_n5391_ & new_n5394_;
  assign new_n5396_ = new_n1202_ & new_n5325_;
  assign new_n5397_ = new_n1194_ & new_n5325_;
  assign new_n5398_ = new_n1190_ & new_n5325_;
  assign new_n5399_ = ~new_n5397_ & ~new_n5398_;
  assign new_n5400_ = ~new_n5396_ & new_n5399_;
  assign new_n5401_ = new_n5395_ & new_n5400_;
  assign new_n5402_ = new_n1213_ & new_n5325_;
  assign new_n5403_ = new_n1204_ & new_n5325_;
  assign new_n5404_ = new_n1200_ & new_n5325_;
  assign new_n5405_ = ~new_n5403_ & ~new_n5404_;
  assign new_n5406_ = ~new_n5402_ & new_n5405_;
  assign new_n5407_ = new_n1216_ & new_n5325_;
  assign new_n5408_ = new_n1210_ & new_n5325_;
  assign new_n5409_ = ~new_n5407_ & ~new_n5408_;
  assign new_n5410_ = new_n5406_ & new_n5409_;
  assign new_n5411_ = new_n5401_ & new_n5410_;
  assign new_n5412_ = new_n5390_ & new_n5411_;
  assign new_n5413_ = new_n1223_ & new_n5325_;
  assign new_n5414_ = new_n1226_ & new_n5325_;
  assign new_n5415_ = new_n1229_ & new_n5325_;
  assign new_n5416_ = ~new_n5414_ & ~new_n5415_;
  assign new_n5417_ = ~new_n5413_ & new_n5416_;
  assign new_n5418_ = new_n1233_ & new_n5325_;
  assign new_n5419_ = new_n1235_ & new_n5325_;
  assign new_n5420_ = new_n1237_ & new_n5325_;
  assign new_n5421_ = ~new_n5419_ & ~new_n5420_;
  assign new_n5422_ = ~new_n5418_ & new_n5421_;
  assign new_n5423_ = new_n5417_ & new_n5422_;
  assign new_n5424_ = A167 & A168;
  assign new_n5425_ = A169 & new_n5424_;
  assign new_n5426_ = new_n371_ & new_n5425_;
  assign new_n5427_ = new_n954_ & new_n5426_;
  assign new_n5428_ = new_n1243_ & new_n5325_;
  assign new_n5429_ = new_n951_ & new_n5426_;
  assign new_n5430_ = ~new_n5428_ & ~new_n5429_;
  assign new_n5431_ = ~new_n5427_ & new_n5430_;
  assign new_n5432_ = new_n967_ & new_n5426_;
  assign new_n5433_ = new_n948_ & new_n5426_;
  assign new_n5434_ = new_n964_ & new_n5426_;
  assign new_n5435_ = ~new_n5433_ & ~new_n5434_;
  assign new_n5436_ = ~new_n5432_ & new_n5435_;
  assign new_n5437_ = new_n5431_ & new_n5436_;
  assign new_n5438_ = new_n5423_ & new_n5437_;
  assign new_n5439_ = new_n978_ & new_n5426_;
  assign new_n5440_ = new_n961_ & new_n5426_;
  assign new_n5441_ = new_n975_ & new_n5426_;
  assign new_n5442_ = ~new_n5440_ & ~new_n5441_;
  assign new_n5443_ = ~new_n5439_ & new_n5442_;
  assign new_n5444_ = new_n990_ & new_n5426_;
  assign new_n5445_ = new_n972_ & new_n5426_;
  assign new_n5446_ = new_n987_ & new_n5426_;
  assign new_n5447_ = ~new_n5445_ & ~new_n5446_;
  assign new_n5448_ = ~new_n5444_ & new_n5447_;
  assign new_n5449_ = new_n5443_ & new_n5448_;
  assign new_n5450_ = new_n996_ & new_n5426_;
  assign new_n5451_ = new_n984_ & new_n5426_;
  assign new_n5452_ = new_n994_ & new_n5426_;
  assign new_n5453_ = ~new_n5451_ & ~new_n5452_;
  assign new_n5454_ = ~new_n5450_ & new_n5453_;
  assign new_n5455_ = new_n1008_ & new_n5426_;
  assign new_n5456_ = new_n1010_ & new_n5426_;
  assign new_n5457_ = ~new_n5455_ & ~new_n5456_;
  assign new_n5458_ = new_n5454_ & new_n5457_;
  assign new_n5459_ = new_n5449_ & new_n5458_;
  assign new_n5460_ = new_n5438_ & new_n5459_;
  assign new_n5461_ = new_n5412_ & new_n5460_;
  assign new_n5462_ = new_n1018_ & new_n5426_;
  assign new_n5463_ = new_n1006_ & new_n5426_;
  assign new_n5464_ = new_n1016_ & new_n5426_;
  assign new_n5465_ = ~new_n5463_ & ~new_n5464_;
  assign new_n5466_ = ~new_n5462_ & new_n5465_;
  assign new_n5467_ = new_n1027_ & new_n5426_;
  assign new_n5468_ = new_n1014_ & new_n5426_;
  assign new_n5469_ = new_n1025_ & new_n5426_;
  assign new_n5470_ = ~new_n5468_ & ~new_n5469_;
  assign new_n5471_ = ~new_n5467_ & new_n5470_;
  assign new_n5472_ = new_n5466_ & new_n5471_;
  assign new_n5473_ = new_n1035_ & new_n5426_;
  assign new_n5474_ = new_n1023_ & new_n5426_;
  assign new_n5475_ = new_n1033_ & new_n5426_;
  assign new_n5476_ = ~new_n5474_ & ~new_n5475_;
  assign new_n5477_ = ~new_n5473_ & new_n5476_;
  assign new_n5478_ = new_n1045_ & new_n5426_;
  assign new_n5479_ = new_n1031_ & new_n5426_;
  assign new_n5480_ = new_n1043_ & new_n5426_;
  assign new_n5481_ = ~new_n5479_ & ~new_n5480_;
  assign new_n5482_ = ~new_n5478_ & new_n5481_;
  assign new_n5483_ = new_n5477_ & new_n5482_;
  assign new_n5484_ = new_n5472_ & new_n5483_;
  assign new_n5485_ = new_n1053_ & new_n5426_;
  assign new_n5486_ = new_n1041_ & new_n5426_;
  assign new_n5487_ = new_n1051_ & new_n5426_;
  assign new_n5488_ = ~new_n5486_ & ~new_n5487_;
  assign new_n5489_ = ~new_n5485_ & new_n5488_;
  assign new_n5490_ = new_n418_ & new_n5425_;
  assign new_n5491_ = new_n1071_ & new_n5490_;
  assign new_n5492_ = new_n1049_ & new_n5426_;
  assign new_n5493_ = new_n1065_ & new_n5490_;
  assign new_n5494_ = ~new_n5492_ & ~new_n5493_;
  assign new_n5495_ = ~new_n5491_ & new_n5494_;
  assign new_n5496_ = new_n5489_ & new_n5495_;
  assign new_n5497_ = new_n1082_ & new_n5490_;
  assign new_n5498_ = new_n1059_ & new_n5490_;
  assign new_n5499_ = new_n1079_ & new_n5490_;
  assign new_n5500_ = ~new_n5498_ & ~new_n5499_;
  assign new_n5501_ = ~new_n5497_ & new_n5500_;
  assign new_n5502_ = new_n1076_ & new_n5490_;
  assign new_n5503_ = new_n1095_ & new_n5490_;
  assign new_n5504_ = ~new_n5502_ & ~new_n5503_;
  assign new_n5505_ = new_n5501_ & new_n5504_;
  assign new_n5506_ = new_n5496_ & new_n5505_;
  assign new_n5507_ = new_n5484_ & new_n5506_;
  assign new_n5508_ = new_n1105_ & new_n5490_;
  assign new_n5509_ = new_n1099_ & new_n5490_;
  assign new_n5510_ = new_n1089_ & new_n5490_;
  assign new_n5511_ = ~new_n5509_ & ~new_n5510_;
  assign new_n5512_ = ~new_n5508_ & new_n5511_;
  assign new_n5513_ = new_n1118_ & new_n5490_;
  assign new_n5514_ = new_n1107_ & new_n5490_;
  assign new_n5515_ = new_n1103_ & new_n5490_;
  assign new_n5516_ = ~new_n5514_ & ~new_n5515_;
  assign new_n5517_ = ~new_n5513_ & new_n5516_;
  assign new_n5518_ = new_n5512_ & new_n5517_;
  assign new_n5519_ = new_n1131_ & new_n5490_;
  assign new_n5520_ = new_n1120_ & new_n5490_;
  assign new_n5521_ = new_n1114_ & new_n5490_;
  assign new_n5522_ = ~new_n5520_ & ~new_n5521_;
  assign new_n5523_ = ~new_n5519_ & new_n5522_;
  assign new_n5524_ = new_n1145_ & new_n5490_;
  assign new_n5525_ = new_n1135_ & new_n5490_;
  assign new_n5526_ = new_n1127_ & new_n5490_;
  assign new_n5527_ = ~new_n5525_ & ~new_n5526_;
  assign new_n5528_ = ~new_n5524_ & new_n5527_;
  assign new_n5529_ = new_n5523_ & new_n5528_;
  assign new_n5530_ = new_n5518_ & new_n5529_;
  assign new_n5531_ = new_n1155_ & new_n5490_;
  assign new_n5532_ = new_n1149_ & new_n5490_;
  assign new_n5533_ = new_n1141_ & new_n5490_;
  assign new_n5534_ = ~new_n5532_ & ~new_n5533_;
  assign new_n5535_ = ~new_n5531_ & new_n5534_;
  assign new_n5536_ = new_n1165_ & new_n5490_;
  assign new_n5537_ = new_n1157_ & new_n5490_;
  assign new_n5538_ = new_n1153_ & new_n5490_;
  assign new_n5539_ = ~new_n5537_ & ~new_n5538_;
  assign new_n5540_ = ~new_n5536_ & new_n5539_;
  assign new_n5541_ = new_n5535_ & new_n5540_;
  assign new_n5542_ = new_n1172_ & new_n5490_;
  assign new_n5543_ = new_n1168_ & new_n5490_;
  assign new_n5544_ = new_n1162_ & new_n5490_;
  assign new_n5545_ = ~new_n5543_ & ~new_n5544_;
  assign new_n5546_ = ~new_n5542_ & new_n5545_;
  assign new_n5547_ = new_n1174_ & new_n5490_;
  assign new_n5548_ = new_n1184_ & new_n5490_;
  assign new_n5549_ = ~new_n5547_ & ~new_n5548_;
  assign new_n5550_ = new_n5546_ & new_n5549_;
  assign new_n5551_ = new_n5541_ & new_n5550_;
  assign new_n5552_ = new_n5530_ & new_n5551_;
  assign new_n5553_ = new_n5507_ & new_n5552_;
  assign new_n5554_ = new_n5461_ & new_n5553_;
  assign new_n5555_ = new_n5367_ & new_n5554_;
  assign new_n5556_ = new_n1192_ & new_n5490_;
  assign new_n5557_ = new_n1186_ & new_n5490_;
  assign new_n5558_ = new_n1182_ & new_n5490_;
  assign new_n5559_ = ~new_n5557_ & ~new_n5558_;
  assign new_n5560_ = ~new_n5556_ & new_n5559_;
  assign new_n5561_ = new_n1202_ & new_n5490_;
  assign new_n5562_ = new_n1194_ & new_n5490_;
  assign new_n5563_ = new_n1190_ & new_n5490_;
  assign new_n5564_ = ~new_n5562_ & ~new_n5563_;
  assign new_n5565_ = ~new_n5561_ & new_n5564_;
  assign new_n5566_ = new_n5560_ & new_n5565_;
  assign new_n5567_ = new_n1213_ & new_n5490_;
  assign new_n5568_ = new_n1204_ & new_n5490_;
  assign new_n5569_ = new_n1200_ & new_n5490_;
  assign new_n5570_ = ~new_n5568_ & ~new_n5569_;
  assign new_n5571_ = ~new_n5567_ & new_n5570_;
  assign new_n5572_ = new_n1226_ & new_n5490_;
  assign new_n5573_ = new_n1216_ & new_n5490_;
  assign new_n5574_ = new_n1210_ & new_n5490_;
  assign new_n5575_ = ~new_n5573_ & ~new_n5574_;
  assign new_n5576_ = ~new_n5572_ & new_n5575_;
  assign new_n5577_ = new_n5571_ & new_n5576_;
  assign new_n5578_ = new_n5566_ & new_n5577_;
  assign new_n5579_ = new_n1235_ & new_n5490_;
  assign new_n5580_ = new_n1229_ & new_n5490_;
  assign new_n5581_ = new_n1223_ & new_n5490_;
  assign new_n5582_ = ~new_n5580_ & ~new_n5581_;
  assign new_n5583_ = ~new_n5579_ & new_n5582_;
  assign new_n5584_ = new_n1243_ & new_n5490_;
  assign new_n5585_ = new_n1237_ & new_n5490_;
  assign new_n5586_ = new_n1233_ & new_n5490_;
  assign new_n5587_ = ~new_n5585_ & ~new_n5586_;
  assign new_n5588_ = ~new_n5584_ & new_n5587_;
  assign new_n5589_ = new_n5583_ & new_n5588_;
  assign new_n5590_ = new_n438_ & new_n5425_;
  assign new_n5591_ = new_n948_ & new_n5590_;
  assign new_n5592_ = new_n951_ & new_n5590_;
  assign new_n5593_ = new_n954_ & new_n5590_;
  assign new_n5594_ = ~new_n5592_ & ~new_n5593_;
  assign new_n5595_ = ~new_n5591_ & new_n5594_;
  assign new_n5596_ = new_n964_ & new_n5590_;
  assign new_n5597_ = new_n967_ & new_n5590_;
  assign new_n5598_ = ~new_n5596_ & ~new_n5597_;
  assign new_n5599_ = new_n5595_ & new_n5598_;
  assign new_n5600_ = new_n5589_ & new_n5599_;
  assign new_n5601_ = new_n5578_ & new_n5600_;
  assign new_n5602_ = new_n978_ & new_n5590_;
  assign new_n5603_ = new_n961_ & new_n5590_;
  assign new_n5604_ = new_n975_ & new_n5590_;
  assign new_n5605_ = ~new_n5603_ & ~new_n5604_;
  assign new_n5606_ = ~new_n5602_ & new_n5605_;
  assign new_n5607_ = new_n990_ & new_n5590_;
  assign new_n5608_ = new_n972_ & new_n5590_;
  assign new_n5609_ = new_n987_ & new_n5590_;
  assign new_n5610_ = ~new_n5608_ & ~new_n5609_;
  assign new_n5611_ = ~new_n5607_ & new_n5610_;
  assign new_n5612_ = new_n5606_ & new_n5611_;
  assign new_n5613_ = new_n996_ & new_n5590_;
  assign new_n5614_ = new_n984_ & new_n5590_;
  assign new_n5615_ = new_n994_ & new_n5590_;
  assign new_n5616_ = ~new_n5614_ & ~new_n5615_;
  assign new_n5617_ = ~new_n5613_ & new_n5616_;
  assign new_n5618_ = new_n1006_ & new_n5590_;
  assign new_n5619_ = new_n1008_ & new_n5590_;
  assign new_n5620_ = new_n1010_ & new_n5590_;
  assign new_n5621_ = ~new_n5619_ & ~new_n5620_;
  assign new_n5622_ = ~new_n5618_ & new_n5621_;
  assign new_n5623_ = new_n5617_ & new_n5622_;
  assign new_n5624_ = new_n5612_ & new_n5623_;
  assign new_n5625_ = new_n1014_ & new_n5590_;
  assign new_n5626_ = new_n1016_ & new_n5590_;
  assign new_n5627_ = new_n1018_ & new_n5590_;
  assign new_n5628_ = ~new_n5626_ & ~new_n5627_;
  assign new_n5629_ = ~new_n5625_ & new_n5628_;
  assign new_n5630_ = new_n1023_ & new_n5590_;
  assign new_n5631_ = new_n1025_ & new_n5590_;
  assign new_n5632_ = new_n1027_ & new_n5590_;
  assign new_n5633_ = ~new_n5631_ & ~new_n5632_;
  assign new_n5634_ = ~new_n5630_ & new_n5633_;
  assign new_n5635_ = new_n5629_ & new_n5634_;
  assign new_n5636_ = new_n1031_ & new_n5590_;
  assign new_n5637_ = new_n1033_ & new_n5590_;
  assign new_n5638_ = new_n1035_ & new_n5590_;
  assign new_n5639_ = ~new_n5637_ & ~new_n5638_;
  assign new_n5640_ = ~new_n5636_ & new_n5639_;
  assign new_n5641_ = new_n1043_ & new_n5590_;
  assign new_n5642_ = new_n1045_ & new_n5590_;
  assign new_n5643_ = ~new_n5641_ & ~new_n5642_;
  assign new_n5644_ = new_n5640_ & new_n5643_;
  assign new_n5645_ = new_n5635_ & new_n5644_;
  assign new_n5646_ = new_n5624_ & new_n5645_;
  assign new_n5647_ = new_n5601_ & new_n5646_;
  assign new_n5648_ = new_n1053_ & new_n5590_;
  assign new_n5649_ = new_n1041_ & new_n5590_;
  assign new_n5650_ = new_n1051_ & new_n5590_;
  assign new_n5651_ = ~new_n5649_ & ~new_n5650_;
  assign new_n5652_ = ~new_n5648_ & new_n5651_;
  assign new_n5653_ = new_n486_ & new_n5425_;
  assign new_n5654_ = new_n1071_ & new_n5653_;
  assign new_n5655_ = new_n1049_ & new_n5590_;
  assign new_n5656_ = new_n1065_ & new_n5653_;
  assign new_n5657_ = ~new_n5655_ & ~new_n5656_;
  assign new_n5658_ = ~new_n5654_ & new_n5657_;
  assign new_n5659_ = new_n5652_ & new_n5658_;
  assign new_n5660_ = new_n1082_ & new_n5653_;
  assign new_n5661_ = new_n1059_ & new_n5653_;
  assign new_n5662_ = new_n1079_ & new_n5653_;
  assign new_n5663_ = ~new_n5661_ & ~new_n5662_;
  assign new_n5664_ = ~new_n5660_ & new_n5663_;
  assign new_n5665_ = new_n1099_ & new_n5653_;
  assign new_n5666_ = new_n1076_ & new_n5653_;
  assign new_n5667_ = new_n1095_ & new_n5653_;
  assign new_n5668_ = ~new_n5666_ & ~new_n5667_;
  assign new_n5669_ = ~new_n5665_ & new_n5668_;
  assign new_n5670_ = new_n5664_ & new_n5669_;
  assign new_n5671_ = new_n5659_ & new_n5670_;
  assign new_n5672_ = new_n1107_ & new_n5653_;
  assign new_n5673_ = new_n1089_ & new_n5653_;
  assign new_n5674_ = new_n1105_ & new_n5653_;
  assign new_n5675_ = ~new_n5673_ & ~new_n5674_;
  assign new_n5676_ = ~new_n5672_ & new_n5675_;
  assign new_n5677_ = new_n1120_ & new_n5653_;
  assign new_n5678_ = new_n1103_ & new_n5653_;
  assign new_n5679_ = new_n1118_ & new_n5653_;
  assign new_n5680_ = ~new_n5678_ & ~new_n5679_;
  assign new_n5681_ = ~new_n5677_ & new_n5680_;
  assign new_n5682_ = new_n5676_ & new_n5681_;
  assign new_n5683_ = new_n1135_ & new_n5653_;
  assign new_n5684_ = new_n1114_ & new_n5653_;
  assign new_n5685_ = new_n1131_ & new_n5653_;
  assign new_n5686_ = ~new_n5684_ & ~new_n5685_;
  assign new_n5687_ = ~new_n5683_ & new_n5686_;
  assign new_n5688_ = new_n1127_ & new_n5653_;
  assign new_n5689_ = new_n1145_ & new_n5653_;
  assign new_n5690_ = ~new_n5688_ & ~new_n5689_;
  assign new_n5691_ = new_n5687_ & new_n5690_;
  assign new_n5692_ = new_n5682_ & new_n5691_;
  assign new_n5693_ = new_n5671_ & new_n5692_;
  assign new_n5694_ = new_n1155_ & new_n5653_;
  assign new_n5695_ = new_n1149_ & new_n5653_;
  assign new_n5696_ = new_n1141_ & new_n5653_;
  assign new_n5697_ = ~new_n5695_ & ~new_n5696_;
  assign new_n5698_ = ~new_n5694_ & new_n5697_;
  assign new_n5699_ = new_n1165_ & new_n5653_;
  assign new_n5700_ = new_n1157_ & new_n5653_;
  assign new_n5701_ = new_n1153_ & new_n5653_;
  assign new_n5702_ = ~new_n5700_ & ~new_n5701_;
  assign new_n5703_ = ~new_n5699_ & new_n5702_;
  assign new_n5704_ = new_n5698_ & new_n5703_;
  assign new_n5705_ = new_n1172_ & new_n5653_;
  assign new_n5706_ = new_n1168_ & new_n5653_;
  assign new_n5707_ = new_n1162_ & new_n5653_;
  assign new_n5708_ = ~new_n5706_ & ~new_n5707_;
  assign new_n5709_ = ~new_n5705_ & new_n5708_;
  assign new_n5710_ = new_n1186_ & new_n5653_;
  assign new_n5711_ = new_n1174_ & new_n5653_;
  assign new_n5712_ = new_n1184_ & new_n5653_;
  assign new_n5713_ = ~new_n5711_ & ~new_n5712_;
  assign new_n5714_ = ~new_n5710_ & new_n5713_;
  assign new_n5715_ = new_n5709_ & new_n5714_;
  assign new_n5716_ = new_n5704_ & new_n5715_;
  assign new_n5717_ = new_n1194_ & new_n5653_;
  assign new_n5718_ = new_n1182_ & new_n5653_;
  assign new_n5719_ = new_n1192_ & new_n5653_;
  assign new_n5720_ = ~new_n5718_ & ~new_n5719_;
  assign new_n5721_ = ~new_n5717_ & new_n5720_;
  assign new_n5722_ = new_n1204_ & new_n5653_;
  assign new_n5723_ = new_n1190_ & new_n5653_;
  assign new_n5724_ = new_n1202_ & new_n5653_;
  assign new_n5725_ = ~new_n5723_ & ~new_n5724_;
  assign new_n5726_ = ~new_n5722_ & new_n5725_;
  assign new_n5727_ = new_n5721_ & new_n5726_;
  assign new_n5728_ = new_n1216_ & new_n5653_;
  assign new_n5729_ = new_n1200_ & new_n5653_;
  assign new_n5730_ = new_n1213_ & new_n5653_;
  assign new_n5731_ = ~new_n5729_ & ~new_n5730_;
  assign new_n5732_ = ~new_n5728_ & new_n5731_;
  assign new_n5733_ = new_n1210_ & new_n5653_;
  assign new_n5734_ = new_n1226_ & new_n5653_;
  assign new_n5735_ = ~new_n5733_ & ~new_n5734_;
  assign new_n5736_ = new_n5732_ & new_n5735_;
  assign new_n5737_ = new_n5727_ & new_n5736_;
  assign new_n5738_ = new_n5716_ & new_n5737_;
  assign new_n5739_ = new_n5693_ & new_n5738_;
  assign new_n5740_ = new_n5647_ & new_n5739_;
  assign new_n5741_ = new_n1235_ & new_n5653_;
  assign new_n5742_ = new_n1229_ & new_n5653_;
  assign new_n5743_ = new_n1223_ & new_n5653_;
  assign new_n5744_ = ~new_n5742_ & ~new_n5743_;
  assign new_n5745_ = ~new_n5741_ & new_n5744_;
  assign new_n5746_ = new_n1243_ & new_n5653_;
  assign new_n5747_ = new_n1237_ & new_n5653_;
  assign new_n5748_ = new_n1233_ & new_n5653_;
  assign new_n5749_ = ~new_n5747_ & ~new_n5748_;
  assign new_n5750_ = ~new_n5746_ & new_n5749_;
  assign new_n5751_ = new_n5745_ & new_n5750_;
  assign new_n5752_ = A170 & new_n4967_;
  assign new_n5753_ = new_n1727_ & new_n5752_;
  assign new_n5754_ = new_n1725_ & new_n5753_;
  assign new_n5755_ = new_n1735_ & new_n5753_;
  assign new_n5756_ = new_n1738_ & new_n5753_;
  assign new_n5757_ = ~new_n5755_ & ~new_n5756_;
  assign new_n5758_ = ~new_n5754_ & new_n5757_;
  assign new_n5759_ = A170 & new_n4982_;
  assign new_n5760_ = new_n1743_ & new_n5759_;
  assign new_n5761_ = new_n1738_ & new_n5760_;
  assign new_n5762_ = new_n1749_ & new_n5753_;
  assign new_n5763_ = new_n1735_ & new_n5760_;
  assign new_n5764_ = ~new_n5762_ & ~new_n5763_;
  assign new_n5765_ = ~new_n5761_ & new_n5764_;
  assign new_n5766_ = new_n5758_ & new_n5765_;
  assign new_n5767_ = new_n5751_ & new_n5766_;
  assign new_n5768_ = A170 & new_n4991_;
  assign new_n5769_ = new_n1757_ & new_n5768_;
  assign new_n5770_ = new_n1735_ & new_n5769_;
  assign new_n5771_ = new_n1725_ & new_n5760_;
  assign new_n5772_ = new_n1749_ & new_n5760_;
  assign new_n5773_ = ~new_n5771_ & ~new_n5772_;
  assign new_n5774_ = ~new_n5770_ & new_n5773_;
  assign new_n5775_ = new_n1749_ & new_n5769_;
  assign new_n5776_ = new_n1738_ & new_n5769_;
  assign new_n5777_ = new_n1725_ & new_n5769_;
  assign new_n5778_ = ~new_n5776_ & ~new_n5777_;
  assign new_n5779_ = ~new_n5775_ & new_n5778_;
  assign new_n5780_ = new_n5774_ & new_n5779_;
  assign new_n5781_ = new_n1773_ & new_n5768_;
  assign new_n5782_ = new_n1725_ & new_n5781_;
  assign new_n5783_ = new_n1735_ & new_n5781_;
  assign new_n5784_ = new_n1738_ & new_n5781_;
  assign new_n5785_ = ~new_n5783_ & ~new_n5784_;
  assign new_n5786_ = ~new_n5782_ & new_n5785_;
  assign new_n5787_ = new_n1749_ & new_n5781_;
  assign new_n5788_ = A170 & new_n5012_;
  assign new_n5789_ = new_n1782_ & new_n5788_;
  assign new_n5790_ = new_n1735_ & new_n5789_;
  assign new_n5791_ = ~new_n5787_ & ~new_n5790_;
  assign new_n5792_ = new_n5786_ & new_n5791_;
  assign new_n5793_ = new_n5780_ & new_n5792_;
  assign new_n5794_ = new_n5767_ & new_n5793_;
  assign new_n5795_ = new_n1749_ & new_n5789_;
  assign new_n5796_ = new_n1738_ & new_n5789_;
  assign new_n5797_ = new_n1725_ & new_n5789_;
  assign new_n5798_ = ~new_n5796_ & ~new_n5797_;
  assign new_n5799_ = ~new_n5795_ & new_n5798_;
  assign new_n5800_ = new_n1796_ & new_n5788_;
  assign new_n5801_ = new_n1725_ & new_n5800_;
  assign new_n5802_ = new_n1735_ & new_n5800_;
  assign new_n5803_ = new_n1738_ & new_n5800_;
  assign new_n5804_ = ~new_n5802_ & ~new_n5803_;
  assign new_n5805_ = ~new_n5801_ & new_n5804_;
  assign new_n5806_ = new_n5799_ & new_n5805_;
  assign new_n5807_ = new_n1805_ & new_n5788_;
  assign new_n5808_ = new_n1738_ & new_n5807_;
  assign new_n5809_ = new_n1749_ & new_n5800_;
  assign new_n5810_ = new_n1735_ & new_n5807_;
  assign new_n5811_ = ~new_n5809_ & ~new_n5810_;
  assign new_n5812_ = ~new_n5808_ & new_n5811_;
  assign new_n5813_ = new_n1813_ & new_n5788_;
  assign new_n5814_ = new_n1735_ & new_n5813_;
  assign new_n5815_ = new_n1725_ & new_n5807_;
  assign new_n5816_ = new_n1749_ & new_n5807_;
  assign new_n5817_ = ~new_n5815_ & ~new_n5816_;
  assign new_n5818_ = ~new_n5814_ & new_n5817_;
  assign new_n5819_ = new_n5812_ & new_n5818_;
  assign new_n5820_ = new_n5806_ & new_n5819_;
  assign new_n5821_ = new_n1749_ & new_n5813_;
  assign new_n5822_ = new_n1738_ & new_n5813_;
  assign new_n5823_ = new_n1725_ & new_n5813_;
  assign new_n5824_ = ~new_n5822_ & ~new_n5823_;
  assign new_n5825_ = ~new_n5821_ & new_n5824_;
  assign new_n5826_ = new_n506_ & new_n5788_;
  assign new_n5827_ = new_n1827_ & new_n5826_;
  assign new_n5828_ = new_n1830_ & new_n5826_;
  assign new_n5829_ = new_n1833_ & new_n5826_;
  assign new_n5830_ = ~new_n5828_ & ~new_n5829_;
  assign new_n5831_ = ~new_n5827_ & new_n5830_;
  assign new_n5832_ = new_n5825_ & new_n5831_;
  assign new_n5833_ = new_n1838_ & new_n5826_;
  assign new_n5834_ = new_n1840_ & new_n5826_;
  assign new_n5835_ = new_n1842_ & new_n5826_;
  assign new_n5836_ = ~new_n5834_ & ~new_n5835_;
  assign new_n5837_ = ~new_n5833_ & new_n5836_;
  assign new_n5838_ = new_n1847_ & new_n5826_;
  assign new_n5839_ = new_n1849_ & new_n5826_;
  assign new_n5840_ = ~new_n5838_ & ~new_n5839_;
  assign new_n5841_ = new_n5837_ & new_n5840_;
  assign new_n5842_ = new_n5832_ & new_n5841_;
  assign new_n5843_ = new_n5820_ & new_n5842_;
  assign new_n5844_ = new_n5794_ & new_n5843_;
  assign new_n5845_ = new_n1855_ & new_n5826_;
  assign new_n5846_ = new_n1857_ & new_n5826_;
  assign new_n5847_ = new_n1859_ & new_n5826_;
  assign new_n5848_ = ~new_n5846_ & ~new_n5847_;
  assign new_n5849_ = ~new_n5845_ & new_n5848_;
  assign new_n5850_ = new_n1864_ & new_n5826_;
  assign new_n5851_ = new_n1866_ & new_n5826_;
  assign new_n5852_ = new_n1868_ & new_n5826_;
  assign new_n5853_ = ~new_n5851_ & ~new_n5852_;
  assign new_n5854_ = ~new_n5850_ & new_n5853_;
  assign new_n5855_ = new_n5849_ & new_n5854_;
  assign new_n5856_ = new_n1875_ & new_n5826_;
  assign new_n5857_ = new_n1878_ & new_n5826_;
  assign new_n5858_ = new_n1881_ & new_n5826_;
  assign new_n5859_ = ~new_n5857_ & ~new_n5858_;
  assign new_n5860_ = ~new_n5856_ & new_n5859_;
  assign new_n5861_ = new_n1886_ & new_n5826_;
  assign new_n5862_ = new_n1889_ & new_n5826_;
  assign new_n5863_ = new_n1892_ & new_n5826_;
  assign new_n5864_ = ~new_n5862_ & ~new_n5863_;
  assign new_n5865_ = ~new_n5861_ & new_n5864_;
  assign new_n5866_ = new_n5860_ & new_n5865_;
  assign new_n5867_ = new_n5855_ & new_n5866_;
  assign new_n5868_ = new_n1898_ & new_n5826_;
  assign new_n5869_ = new_n1900_ & new_n5826_;
  assign new_n5870_ = new_n1902_ & new_n5826_;
  assign new_n5871_ = ~new_n5869_ & ~new_n5870_;
  assign new_n5872_ = ~new_n5868_ & new_n5871_;
  assign new_n5873_ = A170 & new_n5098_;
  assign new_n5874_ = new_n144_ & new_n5873_;
  assign new_n5875_ = new_n954_ & new_n5874_;
  assign new_n5876_ = new_n1913_ & new_n5826_;
  assign new_n5877_ = new_n951_ & new_n5874_;
  assign new_n5878_ = ~new_n5876_ & ~new_n5877_;
  assign new_n5879_ = ~new_n5875_ & new_n5878_;
  assign new_n5880_ = new_n5872_ & new_n5879_;
  assign new_n5881_ = new_n967_ & new_n5874_;
  assign new_n5882_ = new_n948_ & new_n5874_;
  assign new_n5883_ = new_n964_ & new_n5874_;
  assign new_n5884_ = ~new_n5882_ & ~new_n5883_;
  assign new_n5885_ = ~new_n5881_ & new_n5884_;
  assign new_n5886_ = new_n961_ & new_n5874_;
  assign new_n5887_ = new_n975_ & new_n5874_;
  assign new_n5888_ = ~new_n5886_ & ~new_n5887_;
  assign new_n5889_ = new_n5885_ & new_n5888_;
  assign new_n5890_ = new_n5880_ & new_n5889_;
  assign new_n5891_ = new_n5867_ & new_n5890_;
  assign new_n5892_ = new_n987_ & new_n5874_;
  assign new_n5893_ = new_n978_ & new_n5874_;
  assign new_n5894_ = new_n972_ & new_n5874_;
  assign new_n5895_ = ~new_n5893_ & ~new_n5894_;
  assign new_n5896_ = ~new_n5892_ & new_n5895_;
  assign new_n5897_ = new_n994_ & new_n5874_;
  assign new_n5898_ = new_n990_ & new_n5874_;
  assign new_n5899_ = new_n984_ & new_n5874_;
  assign new_n5900_ = ~new_n5898_ & ~new_n5899_;
  assign new_n5901_ = ~new_n5897_ & new_n5900_;
  assign new_n5902_ = new_n5896_ & new_n5901_;
  assign new_n5903_ = new_n1010_ & new_n5874_;
  assign new_n5904_ = new_n996_ & new_n5874_;
  assign new_n5905_ = new_n1008_ & new_n5874_;
  assign new_n5906_ = ~new_n5904_ & ~new_n5905_;
  assign new_n5907_ = ~new_n5903_ & new_n5906_;
  assign new_n5908_ = new_n1018_ & new_n5874_;
  assign new_n5909_ = new_n1006_ & new_n5874_;
  assign new_n5910_ = new_n1016_ & new_n5874_;
  assign new_n5911_ = ~new_n5909_ & ~new_n5910_;
  assign new_n5912_ = ~new_n5908_ & new_n5911_;
  assign new_n5913_ = new_n5907_ & new_n5912_;
  assign new_n5914_ = new_n5902_ & new_n5913_;
  assign new_n5915_ = new_n1027_ & new_n5874_;
  assign new_n5916_ = new_n1014_ & new_n5874_;
  assign new_n5917_ = new_n1025_ & new_n5874_;
  assign new_n5918_ = ~new_n5916_ & ~new_n5917_;
  assign new_n5919_ = ~new_n5915_ & new_n5918_;
  assign new_n5920_ = new_n1035_ & new_n5874_;
  assign new_n5921_ = new_n1023_ & new_n5874_;
  assign new_n5922_ = new_n1033_ & new_n5874_;
  assign new_n5923_ = ~new_n5921_ & ~new_n5922_;
  assign new_n5924_ = ~new_n5920_ & new_n5923_;
  assign new_n5925_ = new_n5919_ & new_n5924_;
  assign new_n5926_ = new_n1045_ & new_n5874_;
  assign new_n5927_ = new_n1031_ & new_n5874_;
  assign new_n5928_ = new_n1043_ & new_n5874_;
  assign new_n5929_ = ~new_n5927_ & ~new_n5928_;
  assign new_n5930_ = ~new_n5926_ & new_n5929_;
  assign new_n5931_ = new_n1041_ & new_n5874_;
  assign new_n5932_ = new_n1051_ & new_n5874_;
  assign new_n5933_ = ~new_n5931_ & ~new_n5932_;
  assign new_n5934_ = new_n5930_ & new_n5933_;
  assign new_n5935_ = new_n5925_ & new_n5934_;
  assign new_n5936_ = new_n5914_ & new_n5935_;
  assign new_n5937_ = new_n5891_ & new_n5936_;
  assign new_n5938_ = new_n5844_ & new_n5937_;
  assign new_n5939_ = new_n5740_ & new_n5938_;
  assign new_n5940_ = new_n5555_ & new_n5939_;
  assign new_n5941_ = new_n265_ & new_n5873_;
  assign new_n5942_ = new_n1065_ & new_n5941_;
  assign new_n5943_ = new_n1053_ & new_n5874_;
  assign new_n5944_ = new_n1049_ & new_n5874_;
  assign new_n5945_ = ~new_n5943_ & ~new_n5944_;
  assign new_n5946_ = ~new_n5942_ & new_n5945_;
  assign new_n5947_ = new_n1079_ & new_n5941_;
  assign new_n5948_ = new_n1071_ & new_n5941_;
  assign new_n5949_ = new_n1059_ & new_n5941_;
  assign new_n5950_ = ~new_n5948_ & ~new_n5949_;
  assign new_n5951_ = ~new_n5947_ & new_n5950_;
  assign new_n5952_ = new_n5946_ & new_n5951_;
  assign new_n5953_ = new_n1095_ & new_n5941_;
  assign new_n5954_ = new_n1082_ & new_n5941_;
  assign new_n5955_ = new_n1076_ & new_n5941_;
  assign new_n5956_ = ~new_n5954_ & ~new_n5955_;
  assign new_n5957_ = ~new_n5953_ & new_n5956_;
  assign new_n5958_ = new_n1105_ & new_n5941_;
  assign new_n5959_ = new_n1099_ & new_n5941_;
  assign new_n5960_ = new_n1089_ & new_n5941_;
  assign new_n5961_ = ~new_n5959_ & ~new_n5960_;
  assign new_n5962_ = ~new_n5958_ & new_n5961_;
  assign new_n5963_ = new_n5957_ & new_n5962_;
  assign new_n5964_ = new_n5952_ & new_n5963_;
  assign new_n5965_ = new_n1118_ & new_n5941_;
  assign new_n5966_ = new_n1107_ & new_n5941_;
  assign new_n5967_ = new_n1103_ & new_n5941_;
  assign new_n5968_ = ~new_n5966_ & ~new_n5967_;
  assign new_n5969_ = ~new_n5965_ & new_n5968_;
  assign new_n5970_ = new_n1131_ & new_n5941_;
  assign new_n5971_ = new_n1120_ & new_n5941_;
  assign new_n5972_ = new_n1114_ & new_n5941_;
  assign new_n5973_ = ~new_n5971_ & ~new_n5972_;
  assign new_n5974_ = ~new_n5970_ & new_n5973_;
  assign new_n5975_ = new_n5969_ & new_n5974_;
  assign new_n5976_ = new_n1145_ & new_n5941_;
  assign new_n5977_ = new_n1135_ & new_n5941_;
  assign new_n5978_ = new_n1127_ & new_n5941_;
  assign new_n5979_ = ~new_n5977_ & ~new_n5978_;
  assign new_n5980_ = ~new_n5976_ & new_n5979_;
  assign new_n5981_ = new_n1155_ & new_n5941_;
  assign new_n5982_ = new_n1149_ & new_n5941_;
  assign new_n5983_ = new_n1141_ & new_n5941_;
  assign new_n5984_ = ~new_n5982_ & ~new_n5983_;
  assign new_n5985_ = ~new_n5981_ & new_n5984_;
  assign new_n5986_ = new_n5980_ & new_n5985_;
  assign new_n5987_ = new_n5975_ & new_n5986_;
  assign new_n5988_ = new_n5964_ & new_n5987_;
  assign new_n5989_ = new_n1165_ & new_n5941_;
  assign new_n5990_ = new_n1157_ & new_n5941_;
  assign new_n5991_ = new_n1153_ & new_n5941_;
  assign new_n5992_ = ~new_n5990_ & ~new_n5991_;
  assign new_n5993_ = ~new_n5989_ & new_n5992_;
  assign new_n5994_ = new_n1172_ & new_n5941_;
  assign new_n5995_ = new_n1168_ & new_n5941_;
  assign new_n5996_ = new_n1162_ & new_n5941_;
  assign new_n5997_ = ~new_n5995_ & ~new_n5996_;
  assign new_n5998_ = ~new_n5994_ & new_n5997_;
  assign new_n5999_ = new_n5993_ & new_n5998_;
  assign new_n6000_ = new_n1186_ & new_n5941_;
  assign new_n6001_ = new_n1174_ & new_n5941_;
  assign new_n6002_ = new_n1184_ & new_n5941_;
  assign new_n6003_ = ~new_n6001_ & ~new_n6002_;
  assign new_n6004_ = ~new_n6000_ & new_n6003_;
  assign new_n6005_ = new_n1194_ & new_n5941_;
  assign new_n6006_ = new_n1182_ & new_n5941_;
  assign new_n6007_ = new_n1192_ & new_n5941_;
  assign new_n6008_ = ~new_n6006_ & ~new_n6007_;
  assign new_n6009_ = ~new_n6005_ & new_n6008_;
  assign new_n6010_ = new_n6004_ & new_n6009_;
  assign new_n6011_ = new_n5999_ & new_n6010_;
  assign new_n6012_ = new_n1204_ & new_n5941_;
  assign new_n6013_ = new_n1190_ & new_n5941_;
  assign new_n6014_ = new_n1202_ & new_n5941_;
  assign new_n6015_ = ~new_n6013_ & ~new_n6014_;
  assign new_n6016_ = ~new_n6012_ & new_n6015_;
  assign new_n6017_ = new_n1216_ & new_n5941_;
  assign new_n6018_ = new_n1200_ & new_n5941_;
  assign new_n6019_ = new_n1213_ & new_n5941_;
  assign new_n6020_ = ~new_n6018_ & ~new_n6019_;
  assign new_n6021_ = ~new_n6017_ & new_n6020_;
  assign new_n6022_ = new_n6016_ & new_n6021_;
  assign new_n6023_ = new_n1229_ & new_n5941_;
  assign new_n6024_ = new_n1210_ & new_n5941_;
  assign new_n6025_ = new_n1226_ & new_n5941_;
  assign new_n6026_ = ~new_n6024_ & ~new_n6025_;
  assign new_n6027_ = ~new_n6023_ & new_n6026_;
  assign new_n6028_ = new_n1223_ & new_n5941_;
  assign new_n6029_ = new_n1235_ & new_n5941_;
  assign new_n6030_ = ~new_n6028_ & ~new_n6029_;
  assign new_n6031_ = new_n6027_ & new_n6030_;
  assign new_n6032_ = new_n6022_ & new_n6031_;
  assign new_n6033_ = new_n6011_ & new_n6032_;
  assign new_n6034_ = new_n5988_ & new_n6033_;
  assign new_n6035_ = new_n1243_ & new_n5941_;
  assign new_n6036_ = new_n1237_ & new_n5941_;
  assign new_n6037_ = new_n1233_ & new_n5941_;
  assign new_n6038_ = ~new_n6036_ & ~new_n6037_;
  assign new_n6039_ = ~new_n6035_ & new_n6038_;
  assign new_n6040_ = new_n293_ & new_n5873_;
  assign new_n6041_ = new_n948_ & new_n6040_;
  assign new_n6042_ = new_n951_ & new_n6040_;
  assign new_n6043_ = new_n954_ & new_n6040_;
  assign new_n6044_ = ~new_n6042_ & ~new_n6043_;
  assign new_n6045_ = ~new_n6041_ & new_n6044_;
  assign new_n6046_ = new_n6039_ & new_n6045_;
  assign new_n6047_ = new_n961_ & new_n6040_;
  assign new_n6048_ = new_n964_ & new_n6040_;
  assign new_n6049_ = new_n967_ & new_n6040_;
  assign new_n6050_ = ~new_n6048_ & ~new_n6049_;
  assign new_n6051_ = ~new_n6047_ & new_n6050_;
  assign new_n6052_ = new_n972_ & new_n6040_;
  assign new_n6053_ = new_n975_ & new_n6040_;
  assign new_n6054_ = new_n978_ & new_n6040_;
  assign new_n6055_ = ~new_n6053_ & ~new_n6054_;
  assign new_n6056_ = ~new_n6052_ & new_n6055_;
  assign new_n6057_ = new_n6051_ & new_n6056_;
  assign new_n6058_ = new_n6046_ & new_n6057_;
  assign new_n6059_ = new_n984_ & new_n6040_;
  assign new_n6060_ = new_n987_ & new_n6040_;
  assign new_n6061_ = new_n990_ & new_n6040_;
  assign new_n6062_ = ~new_n6060_ & ~new_n6061_;
  assign new_n6063_ = ~new_n6059_ & new_n6062_;
  assign new_n6064_ = new_n1008_ & new_n6040_;
  assign new_n6065_ = new_n994_ & new_n6040_;
  assign new_n6066_ = new_n996_ & new_n6040_;
  assign new_n6067_ = ~new_n6065_ & ~new_n6066_;
  assign new_n6068_ = ~new_n6064_ & new_n6067_;
  assign new_n6069_ = new_n6063_ & new_n6068_;
  assign new_n6070_ = new_n1016_ & new_n6040_;
  assign new_n6071_ = new_n1010_ & new_n6040_;
  assign new_n6072_ = new_n1006_ & new_n6040_;
  assign new_n6073_ = ~new_n6071_ & ~new_n6072_;
  assign new_n6074_ = ~new_n6070_ & new_n6073_;
  assign new_n6075_ = new_n1018_ & new_n6040_;
  assign new_n6076_ = new_n1014_ & new_n6040_;
  assign new_n6077_ = ~new_n6075_ & ~new_n6076_;
  assign new_n6078_ = new_n6074_ & new_n6077_;
  assign new_n6079_ = new_n6069_ & new_n6078_;
  assign new_n6080_ = new_n6058_ & new_n6079_;
  assign new_n6081_ = new_n1023_ & new_n6040_;
  assign new_n6082_ = new_n1025_ & new_n6040_;
  assign new_n6083_ = new_n1027_ & new_n6040_;
  assign new_n6084_ = ~new_n6082_ & ~new_n6083_;
  assign new_n6085_ = ~new_n6081_ & new_n6084_;
  assign new_n6086_ = new_n1031_ & new_n6040_;
  assign new_n6087_ = new_n1033_ & new_n6040_;
  assign new_n6088_ = new_n1035_ & new_n6040_;
  assign new_n6089_ = ~new_n6087_ & ~new_n6088_;
  assign new_n6090_ = ~new_n6086_ & new_n6089_;
  assign new_n6091_ = new_n6085_ & new_n6090_;
  assign new_n6092_ = new_n1041_ & new_n6040_;
  assign new_n6093_ = new_n1043_ & new_n6040_;
  assign new_n6094_ = new_n1045_ & new_n6040_;
  assign new_n6095_ = ~new_n6093_ & ~new_n6094_;
  assign new_n6096_ = ~new_n6092_ & new_n6095_;
  assign new_n6097_ = new_n1049_ & new_n6040_;
  assign new_n6098_ = new_n1051_ & new_n6040_;
  assign new_n6099_ = new_n1053_ & new_n6040_;
  assign new_n6100_ = ~new_n6098_ & ~new_n6099_;
  assign new_n6101_ = ~new_n6097_ & new_n6100_;
  assign new_n6102_ = new_n6096_ & new_n6101_;
  assign new_n6103_ = new_n6091_ & new_n6102_;
  assign new_n6104_ = new_n351_ & new_n5873_;
  assign new_n6105_ = new_n1059_ & new_n6104_;
  assign new_n6106_ = new_n1065_ & new_n6104_;
  assign new_n6107_ = new_n1071_ & new_n6104_;
  assign new_n6108_ = ~new_n6106_ & ~new_n6107_;
  assign new_n6109_ = ~new_n6105_ & new_n6108_;
  assign new_n6110_ = new_n1076_ & new_n6104_;
  assign new_n6111_ = new_n1079_ & new_n6104_;
  assign new_n6112_ = new_n1082_ & new_n6104_;
  assign new_n6113_ = ~new_n6111_ & ~new_n6112_;
  assign new_n6114_ = ~new_n6110_ & new_n6113_;
  assign new_n6115_ = new_n6109_ & new_n6114_;
  assign new_n6116_ = new_n1089_ & new_n6104_;
  assign new_n6117_ = new_n1095_ & new_n6104_;
  assign new_n6118_ = new_n1099_ & new_n6104_;
  assign new_n6119_ = ~new_n6117_ & ~new_n6118_;
  assign new_n6120_ = ~new_n6116_ & new_n6119_;
  assign new_n6121_ = new_n1105_ & new_n6104_;
  assign new_n6122_ = new_n1107_ & new_n6104_;
  assign new_n6123_ = ~new_n6121_ & ~new_n6122_;
  assign new_n6124_ = new_n6120_ & new_n6123_;
  assign new_n6125_ = new_n6115_ & new_n6124_;
  assign new_n6126_ = new_n6103_ & new_n6125_;
  assign new_n6127_ = new_n6080_ & new_n6126_;
  assign new_n6128_ = new_n6034_ & new_n6127_;
  assign new_n6129_ = new_n1120_ & new_n6104_;
  assign new_n6130_ = new_n1103_ & new_n6104_;
  assign new_n6131_ = new_n1118_ & new_n6104_;
  assign new_n6132_ = ~new_n6130_ & ~new_n6131_;
  assign new_n6133_ = ~new_n6129_ & new_n6132_;
  assign new_n6134_ = new_n1135_ & new_n6104_;
  assign new_n6135_ = new_n1114_ & new_n6104_;
  assign new_n6136_ = new_n1131_ & new_n6104_;
  assign new_n6137_ = ~new_n6135_ & ~new_n6136_;
  assign new_n6138_ = ~new_n6134_ & new_n6137_;
  assign new_n6139_ = new_n6133_ & new_n6138_;
  assign new_n6140_ = new_n1149_ & new_n6104_;
  assign new_n6141_ = new_n1127_ & new_n6104_;
  assign new_n6142_ = new_n1145_ & new_n6104_;
  assign new_n6143_ = ~new_n6141_ & ~new_n6142_;
  assign new_n6144_ = ~new_n6140_ & new_n6143_;
  assign new_n6145_ = new_n1157_ & new_n6104_;
  assign new_n6146_ = new_n1141_ & new_n6104_;
  assign new_n6147_ = new_n1155_ & new_n6104_;
  assign new_n6148_ = ~new_n6146_ & ~new_n6147_;
  assign new_n6149_ = ~new_n6145_ & new_n6148_;
  assign new_n6150_ = new_n6144_ & new_n6149_;
  assign new_n6151_ = new_n6139_ & new_n6150_;
  assign new_n6152_ = new_n1168_ & new_n6104_;
  assign new_n6153_ = new_n1153_ & new_n6104_;
  assign new_n6154_ = new_n1165_ & new_n6104_;
  assign new_n6155_ = ~new_n6153_ & ~new_n6154_;
  assign new_n6156_ = ~new_n6152_ & new_n6155_;
  assign new_n6157_ = new_n1174_ & new_n6104_;
  assign new_n6158_ = new_n1162_ & new_n6104_;
  assign new_n6159_ = new_n1172_ & new_n6104_;
  assign new_n6160_ = ~new_n6158_ & ~new_n6159_;
  assign new_n6161_ = ~new_n6157_ & new_n6160_;
  assign new_n6162_ = new_n6156_ & new_n6161_;
  assign new_n6163_ = new_n1182_ & new_n6104_;
  assign new_n6164_ = new_n1184_ & new_n6104_;
  assign new_n6165_ = new_n1186_ & new_n6104_;
  assign new_n6166_ = ~new_n6164_ & ~new_n6165_;
  assign new_n6167_ = ~new_n6163_ & new_n6166_;
  assign new_n6168_ = new_n1192_ & new_n6104_;
  assign new_n6169_ = new_n1194_ & new_n6104_;
  assign new_n6170_ = ~new_n6168_ & ~new_n6169_;
  assign new_n6171_ = new_n6167_ & new_n6170_;
  assign new_n6172_ = new_n6162_ & new_n6171_;
  assign new_n6173_ = new_n6151_ & new_n6172_;
  assign new_n6174_ = new_n1204_ & new_n6104_;
  assign new_n6175_ = new_n1190_ & new_n6104_;
  assign new_n6176_ = new_n1202_ & new_n6104_;
  assign new_n6177_ = ~new_n6175_ & ~new_n6176_;
  assign new_n6178_ = ~new_n6174_ & new_n6177_;
  assign new_n6179_ = new_n1216_ & new_n6104_;
  assign new_n6180_ = new_n1200_ & new_n6104_;
  assign new_n6181_ = new_n1213_ & new_n6104_;
  assign new_n6182_ = ~new_n6180_ & ~new_n6181_;
  assign new_n6183_ = ~new_n6179_ & new_n6182_;
  assign new_n6184_ = new_n6178_ & new_n6183_;
  assign new_n6185_ = new_n1229_ & new_n6104_;
  assign new_n6186_ = new_n1210_ & new_n6104_;
  assign new_n6187_ = new_n1226_ & new_n6104_;
  assign new_n6188_ = ~new_n6186_ & ~new_n6187_;
  assign new_n6189_ = ~new_n6185_ & new_n6188_;
  assign new_n6190_ = new_n1237_ & new_n6104_;
  assign new_n6191_ = new_n1223_ & new_n6104_;
  assign new_n6192_ = new_n1235_ & new_n6104_;
  assign new_n6193_ = ~new_n6191_ & ~new_n6192_;
  assign new_n6194_ = ~new_n6190_ & new_n6193_;
  assign new_n6195_ = new_n6189_ & new_n6194_;
  assign new_n6196_ = new_n6184_ & new_n6195_;
  assign new_n6197_ = A170 & new_n5424_;
  assign new_n6198_ = new_n371_ & new_n6197_;
  assign new_n6199_ = new_n951_ & new_n6198_;
  assign new_n6200_ = new_n1233_ & new_n6104_;
  assign new_n6201_ = new_n1243_ & new_n6104_;
  assign new_n6202_ = ~new_n6200_ & ~new_n6201_;
  assign new_n6203_ = ~new_n6199_ & new_n6202_;
  assign new_n6204_ = new_n964_ & new_n6198_;
  assign new_n6205_ = new_n954_ & new_n6198_;
  assign new_n6206_ = new_n948_ & new_n6198_;
  assign new_n6207_ = ~new_n6205_ & ~new_n6206_;
  assign new_n6208_ = ~new_n6204_ & new_n6207_;
  assign new_n6209_ = new_n6203_ & new_n6208_;
  assign new_n6210_ = new_n975_ & new_n6198_;
  assign new_n6211_ = new_n967_ & new_n6198_;
  assign new_n6212_ = new_n961_ & new_n6198_;
  assign new_n6213_ = ~new_n6211_ & ~new_n6212_;
  assign new_n6214_ = ~new_n6210_ & new_n6213_;
  assign new_n6215_ = new_n978_ & new_n6198_;
  assign new_n6216_ = new_n972_ & new_n6198_;
  assign new_n6217_ = ~new_n6215_ & ~new_n6216_;
  assign new_n6218_ = new_n6214_ & new_n6217_;
  assign new_n6219_ = new_n6209_ & new_n6218_;
  assign new_n6220_ = new_n6196_ & new_n6219_;
  assign new_n6221_ = new_n6173_ & new_n6220_;
  assign new_n6222_ = new_n984_ & new_n6198_;
  assign new_n6223_ = new_n987_ & new_n6198_;
  assign new_n6224_ = new_n990_ & new_n6198_;
  assign new_n6225_ = ~new_n6223_ & ~new_n6224_;
  assign new_n6226_ = ~new_n6222_ & new_n6225_;
  assign new_n6227_ = new_n1008_ & new_n6198_;
  assign new_n6228_ = new_n994_ & new_n6198_;
  assign new_n6229_ = new_n996_ & new_n6198_;
  assign new_n6230_ = ~new_n6228_ & ~new_n6229_;
  assign new_n6231_ = ~new_n6227_ & new_n6230_;
  assign new_n6232_ = new_n6226_ & new_n6231_;
  assign new_n6233_ = new_n1016_ & new_n6198_;
  assign new_n6234_ = new_n1010_ & new_n6198_;
  assign new_n6235_ = new_n1006_ & new_n6198_;
  assign new_n6236_ = ~new_n6234_ & ~new_n6235_;
  assign new_n6237_ = ~new_n6233_ & new_n6236_;
  assign new_n6238_ = new_n1025_ & new_n6198_;
  assign new_n6239_ = new_n1018_ & new_n6198_;
  assign new_n6240_ = new_n1014_ & new_n6198_;
  assign new_n6241_ = ~new_n6239_ & ~new_n6240_;
  assign new_n6242_ = ~new_n6238_ & new_n6241_;
  assign new_n6243_ = new_n6237_ & new_n6242_;
  assign new_n6244_ = new_n6232_ & new_n6243_;
  assign new_n6245_ = new_n1033_ & new_n6198_;
  assign new_n6246_ = new_n1027_ & new_n6198_;
  assign new_n6247_ = new_n1023_ & new_n6198_;
  assign new_n6248_ = ~new_n6246_ & ~new_n6247_;
  assign new_n6249_ = ~new_n6245_ & new_n6248_;
  assign new_n6250_ = new_n1043_ & new_n6198_;
  assign new_n6251_ = new_n1035_ & new_n6198_;
  assign new_n6252_ = new_n1031_ & new_n6198_;
  assign new_n6253_ = ~new_n6251_ & ~new_n6252_;
  assign new_n6254_ = ~new_n6250_ & new_n6253_;
  assign new_n6255_ = new_n6249_ & new_n6254_;
  assign new_n6256_ = new_n1051_ & new_n6198_;
  assign new_n6257_ = new_n1045_ & new_n6198_;
  assign new_n6258_ = new_n1041_ & new_n6198_;
  assign new_n6259_ = ~new_n6257_ & ~new_n6258_;
  assign new_n6260_ = ~new_n6256_ & new_n6259_;
  assign new_n6261_ = new_n1053_ & new_n6198_;
  assign new_n6262_ = new_n1049_ & new_n6198_;
  assign new_n6263_ = ~new_n6261_ & ~new_n6262_;
  assign new_n6264_ = new_n6260_ & new_n6263_;
  assign new_n6265_ = new_n6255_ & new_n6264_;
  assign new_n6266_ = new_n6244_ & new_n6265_;
  assign new_n6267_ = new_n418_ & new_n6197_;
  assign new_n6268_ = new_n1059_ & new_n6267_;
  assign new_n6269_ = new_n1065_ & new_n6267_;
  assign new_n6270_ = new_n1071_ & new_n6267_;
  assign new_n6271_ = ~new_n6269_ & ~new_n6270_;
  assign new_n6272_ = ~new_n6268_ & new_n6271_;
  assign new_n6273_ = new_n1076_ & new_n6267_;
  assign new_n6274_ = new_n1079_ & new_n6267_;
  assign new_n6275_ = new_n1082_ & new_n6267_;
  assign new_n6276_ = ~new_n6274_ & ~new_n6275_;
  assign new_n6277_ = ~new_n6273_ & new_n6276_;
  assign new_n6278_ = new_n6272_ & new_n6277_;
  assign new_n6279_ = new_n1089_ & new_n6267_;
  assign new_n6280_ = new_n1095_ & new_n6267_;
  assign new_n6281_ = new_n1099_ & new_n6267_;
  assign new_n6282_ = ~new_n6280_ & ~new_n6281_;
  assign new_n6283_ = ~new_n6279_ & new_n6282_;
  assign new_n6284_ = new_n1103_ & new_n6267_;
  assign new_n6285_ = new_n1105_ & new_n6267_;
  assign new_n6286_ = new_n1107_ & new_n6267_;
  assign new_n6287_ = ~new_n6285_ & ~new_n6286_;
  assign new_n6288_ = ~new_n6284_ & new_n6287_;
  assign new_n6289_ = new_n6283_ & new_n6288_;
  assign new_n6290_ = new_n6278_ & new_n6289_;
  assign new_n6291_ = new_n1114_ & new_n6267_;
  assign new_n6292_ = new_n1118_ & new_n6267_;
  assign new_n6293_ = new_n1120_ & new_n6267_;
  assign new_n6294_ = ~new_n6292_ & ~new_n6293_;
  assign new_n6295_ = ~new_n6291_ & new_n6294_;
  assign new_n6296_ = new_n1127_ & new_n6267_;
  assign new_n6297_ = new_n1131_ & new_n6267_;
  assign new_n6298_ = new_n1135_ & new_n6267_;
  assign new_n6299_ = ~new_n6297_ & ~new_n6298_;
  assign new_n6300_ = ~new_n6296_ & new_n6299_;
  assign new_n6301_ = new_n6295_ & new_n6300_;
  assign new_n6302_ = new_n1141_ & new_n6267_;
  assign new_n6303_ = new_n1145_ & new_n6267_;
  assign new_n6304_ = new_n1149_ & new_n6267_;
  assign new_n6305_ = ~new_n6303_ & ~new_n6304_;
  assign new_n6306_ = ~new_n6302_ & new_n6305_;
  assign new_n6307_ = new_n1155_ & new_n6267_;
  assign new_n6308_ = new_n1157_ & new_n6267_;
  assign new_n6309_ = ~new_n6307_ & ~new_n6308_;
  assign new_n6310_ = new_n6306_ & new_n6309_;
  assign new_n6311_ = new_n6301_ & new_n6310_;
  assign new_n6312_ = new_n6290_ & new_n6311_;
  assign new_n6313_ = new_n6266_ & new_n6312_;
  assign new_n6314_ = new_n6221_ & new_n6313_;
  assign new_n6315_ = new_n6128_ & new_n6314_;
  assign new_n6316_ = new_n1168_ & new_n6267_;
  assign new_n6317_ = new_n1153_ & new_n6267_;
  assign new_n6318_ = new_n1165_ & new_n6267_;
  assign new_n6319_ = ~new_n6317_ & ~new_n6318_;
  assign new_n6320_ = ~new_n6316_ & new_n6319_;
  assign new_n6321_ = new_n1174_ & new_n6267_;
  assign new_n6322_ = new_n1162_ & new_n6267_;
  assign new_n6323_ = new_n1172_ & new_n6267_;
  assign new_n6324_ = ~new_n6322_ & ~new_n6323_;
  assign new_n6325_ = ~new_n6321_ & new_n6324_;
  assign new_n6326_ = new_n6320_ & new_n6325_;
  assign new_n6327_ = new_n1182_ & new_n6267_;
  assign new_n6328_ = new_n1184_ & new_n6267_;
  assign new_n6329_ = new_n1186_ & new_n6267_;
  assign new_n6330_ = ~new_n6328_ & ~new_n6329_;
  assign new_n6331_ = ~new_n6327_ & new_n6330_;
  assign new_n6332_ = new_n1190_ & new_n6267_;
  assign new_n6333_ = new_n1192_ & new_n6267_;
  assign new_n6334_ = new_n1194_ & new_n6267_;
  assign new_n6335_ = ~new_n6333_ & ~new_n6334_;
  assign new_n6336_ = ~new_n6332_ & new_n6335_;
  assign new_n6337_ = new_n6331_ & new_n6336_;
  assign new_n6338_ = new_n6326_ & new_n6337_;
  assign new_n6339_ = new_n1200_ & new_n6267_;
  assign new_n6340_ = new_n1202_ & new_n6267_;
  assign new_n6341_ = new_n1204_ & new_n6267_;
  assign new_n6342_ = ~new_n6340_ & ~new_n6341_;
  assign new_n6343_ = ~new_n6339_ & new_n6342_;
  assign new_n6344_ = new_n1210_ & new_n6267_;
  assign new_n6345_ = new_n1213_ & new_n6267_;
  assign new_n6346_ = new_n1216_ & new_n6267_;
  assign new_n6347_ = ~new_n6345_ & ~new_n6346_;
  assign new_n6348_ = ~new_n6344_ & new_n6347_;
  assign new_n6349_ = new_n6343_ & new_n6348_;
  assign new_n6350_ = new_n1223_ & new_n6267_;
  assign new_n6351_ = new_n1226_ & new_n6267_;
  assign new_n6352_ = new_n1229_ & new_n6267_;
  assign new_n6353_ = ~new_n6351_ & ~new_n6352_;
  assign new_n6354_ = ~new_n6350_ & new_n6353_;
  assign new_n6355_ = new_n1235_ & new_n6267_;
  assign new_n6356_ = new_n1237_ & new_n6267_;
  assign new_n6357_ = ~new_n6355_ & ~new_n6356_;
  assign new_n6358_ = new_n6354_ & new_n6357_;
  assign new_n6359_ = new_n6349_ & new_n6358_;
  assign new_n6360_ = new_n6338_ & new_n6359_;
  assign new_n6361_ = new_n438_ & new_n6197_;
  assign new_n6362_ = new_n951_ & new_n6361_;
  assign new_n6363_ = new_n1233_ & new_n6267_;
  assign new_n6364_ = new_n1243_ & new_n6267_;
  assign new_n6365_ = ~new_n6363_ & ~new_n6364_;
  assign new_n6366_ = ~new_n6362_ & new_n6365_;
  assign new_n6367_ = new_n964_ & new_n6361_;
  assign new_n6368_ = new_n954_ & new_n6361_;
  assign new_n6369_ = new_n948_ & new_n6361_;
  assign new_n6370_ = ~new_n6368_ & ~new_n6369_;
  assign new_n6371_ = ~new_n6367_ & new_n6370_;
  assign new_n6372_ = new_n6366_ & new_n6371_;
  assign new_n6373_ = new_n975_ & new_n6361_;
  assign new_n6374_ = new_n967_ & new_n6361_;
  assign new_n6375_ = new_n961_ & new_n6361_;
  assign new_n6376_ = ~new_n6374_ & ~new_n6375_;
  assign new_n6377_ = ~new_n6373_ & new_n6376_;
  assign new_n6378_ = new_n987_ & new_n6361_;
  assign new_n6379_ = new_n978_ & new_n6361_;
  assign new_n6380_ = new_n972_ & new_n6361_;
  assign new_n6381_ = ~new_n6379_ & ~new_n6380_;
  assign new_n6382_ = ~new_n6378_ & new_n6381_;
  assign new_n6383_ = new_n6377_ & new_n6382_;
  assign new_n6384_ = new_n6372_ & new_n6383_;
  assign new_n6385_ = new_n994_ & new_n6361_;
  assign new_n6386_ = new_n990_ & new_n6361_;
  assign new_n6387_ = new_n984_ & new_n6361_;
  assign new_n6388_ = ~new_n6386_ & ~new_n6387_;
  assign new_n6389_ = ~new_n6385_ & new_n6388_;
  assign new_n6390_ = new_n1010_ & new_n6361_;
  assign new_n6391_ = new_n996_ & new_n6361_;
  assign new_n6392_ = new_n1008_ & new_n6361_;
  assign new_n6393_ = ~new_n6391_ & ~new_n6392_;
  assign new_n6394_ = ~new_n6390_ & new_n6393_;
  assign new_n6395_ = new_n6389_ & new_n6394_;
  assign new_n6396_ = new_n1018_ & new_n6361_;
  assign new_n6397_ = new_n1006_ & new_n6361_;
  assign new_n6398_ = new_n1016_ & new_n6361_;
  assign new_n6399_ = ~new_n6397_ & ~new_n6398_;
  assign new_n6400_ = ~new_n6396_ & new_n6399_;
  assign new_n6401_ = new_n1014_ & new_n6361_;
  assign new_n6402_ = new_n1025_ & new_n6361_;
  assign new_n6403_ = ~new_n6401_ & ~new_n6402_;
  assign new_n6404_ = new_n6400_ & new_n6403_;
  assign new_n6405_ = new_n6395_ & new_n6404_;
  assign new_n6406_ = new_n6384_ & new_n6405_;
  assign new_n6407_ = new_n6360_ & new_n6406_;
  assign new_n6408_ = new_n1033_ & new_n6361_;
  assign new_n6409_ = new_n1027_ & new_n6361_;
  assign new_n6410_ = new_n1023_ & new_n6361_;
  assign new_n6411_ = ~new_n6409_ & ~new_n6410_;
  assign new_n6412_ = ~new_n6408_ & new_n6411_;
  assign new_n6413_ = new_n1043_ & new_n6361_;
  assign new_n6414_ = new_n1035_ & new_n6361_;
  assign new_n6415_ = new_n1031_ & new_n6361_;
  assign new_n6416_ = ~new_n6414_ & ~new_n6415_;
  assign new_n6417_ = ~new_n6413_ & new_n6416_;
  assign new_n6418_ = new_n6412_ & new_n6417_;
  assign new_n6419_ = new_n1051_ & new_n6361_;
  assign new_n6420_ = new_n1045_ & new_n6361_;
  assign new_n6421_ = new_n1041_ & new_n6361_;
  assign new_n6422_ = ~new_n6420_ & ~new_n6421_;
  assign new_n6423_ = ~new_n6419_ & new_n6422_;
  assign new_n6424_ = new_n486_ & new_n6197_;
  assign new_n6425_ = new_n1065_ & new_n6424_;
  assign new_n6426_ = new_n1053_ & new_n6361_;
  assign new_n6427_ = new_n1049_ & new_n6361_;
  assign new_n6428_ = ~new_n6426_ & ~new_n6427_;
  assign new_n6429_ = ~new_n6425_ & new_n6428_;
  assign new_n6430_ = new_n6423_ & new_n6429_;
  assign new_n6431_ = new_n6418_ & new_n6430_;
  assign new_n6432_ = new_n1079_ & new_n6424_;
  assign new_n6433_ = new_n1071_ & new_n6424_;
  assign new_n6434_ = new_n1059_ & new_n6424_;
  assign new_n6435_ = ~new_n6433_ & ~new_n6434_;
  assign new_n6436_ = ~new_n6432_ & new_n6435_;
  assign new_n6437_ = new_n1095_ & new_n6424_;
  assign new_n6438_ = new_n1082_ & new_n6424_;
  assign new_n6439_ = new_n1076_ & new_n6424_;
  assign new_n6440_ = ~new_n6438_ & ~new_n6439_;
  assign new_n6441_ = ~new_n6437_ & new_n6440_;
  assign new_n6442_ = new_n6436_ & new_n6441_;
  assign new_n6443_ = new_n1105_ & new_n6424_;
  assign new_n6444_ = new_n1099_ & new_n6424_;
  assign new_n6445_ = new_n1089_ & new_n6424_;
  assign new_n6446_ = ~new_n6444_ & ~new_n6445_;
  assign new_n6447_ = ~new_n6443_ & new_n6446_;
  assign new_n6448_ = new_n1107_ & new_n6424_;
  assign new_n6449_ = new_n1103_ & new_n6424_;
  assign new_n6450_ = ~new_n6448_ & ~new_n6449_;
  assign new_n6451_ = new_n6447_ & new_n6450_;
  assign new_n6452_ = new_n6442_ & new_n6451_;
  assign new_n6453_ = new_n6431_ & new_n6452_;
  assign new_n6454_ = new_n1114_ & new_n6424_;
  assign new_n6455_ = new_n1118_ & new_n6424_;
  assign new_n6456_ = new_n1120_ & new_n6424_;
  assign new_n6457_ = ~new_n6455_ & ~new_n6456_;
  assign new_n6458_ = ~new_n6454_ & new_n6457_;
  assign new_n6459_ = new_n1127_ & new_n6424_;
  assign new_n6460_ = new_n1131_ & new_n6424_;
  assign new_n6461_ = new_n1135_ & new_n6424_;
  assign new_n6462_ = ~new_n6460_ & ~new_n6461_;
  assign new_n6463_ = ~new_n6459_ & new_n6462_;
  assign new_n6464_ = new_n6458_ & new_n6463_;
  assign new_n6465_ = new_n1141_ & new_n6424_;
  assign new_n6466_ = new_n1145_ & new_n6424_;
  assign new_n6467_ = new_n1149_ & new_n6424_;
  assign new_n6468_ = ~new_n6466_ & ~new_n6467_;
  assign new_n6469_ = ~new_n6465_ & new_n6468_;
  assign new_n6470_ = new_n1153_ & new_n6424_;
  assign new_n6471_ = new_n1155_ & new_n6424_;
  assign new_n6472_ = new_n1157_ & new_n6424_;
  assign new_n6473_ = ~new_n6471_ & ~new_n6472_;
  assign new_n6474_ = ~new_n6470_ & new_n6473_;
  assign new_n6475_ = new_n6469_ & new_n6474_;
  assign new_n6476_ = new_n6464_ & new_n6475_;
  assign new_n6477_ = new_n1162_ & new_n6424_;
  assign new_n6478_ = new_n1165_ & new_n6424_;
  assign new_n6479_ = new_n1168_ & new_n6424_;
  assign new_n6480_ = ~new_n6478_ & ~new_n6479_;
  assign new_n6481_ = ~new_n6477_ & new_n6480_;
  assign new_n6482_ = new_n1184_ & new_n6424_;
  assign new_n6483_ = new_n1172_ & new_n6424_;
  assign new_n6484_ = new_n1174_ & new_n6424_;
  assign new_n6485_ = ~new_n6483_ & ~new_n6484_;
  assign new_n6486_ = ~new_n6482_ & new_n6485_;
  assign new_n6487_ = new_n6481_ & new_n6486_;
  assign new_n6488_ = new_n1192_ & new_n6424_;
  assign new_n6489_ = new_n1186_ & new_n6424_;
  assign new_n6490_ = new_n1182_ & new_n6424_;
  assign new_n6491_ = ~new_n6489_ & ~new_n6490_;
  assign new_n6492_ = ~new_n6488_ & new_n6491_;
  assign new_n6493_ = new_n1194_ & new_n6424_;
  assign new_n6494_ = new_n1190_ & new_n6424_;
  assign new_n6495_ = ~new_n6493_ & ~new_n6494_;
  assign new_n6496_ = new_n6492_ & new_n6495_;
  assign new_n6497_ = new_n6487_ & new_n6496_;
  assign new_n6498_ = new_n6476_ & new_n6497_;
  assign new_n6499_ = new_n6453_ & new_n6498_;
  assign new_n6500_ = new_n6407_ & new_n6499_;
  assign new_n6501_ = new_n1200_ & new_n6424_;
  assign new_n6502_ = new_n1202_ & new_n6424_;
  assign new_n6503_ = new_n1204_ & new_n6424_;
  assign new_n6504_ = ~new_n6502_ & ~new_n6503_;
  assign new_n6505_ = ~new_n6501_ & new_n6504_;
  assign new_n6506_ = new_n1210_ & new_n6424_;
  assign new_n6507_ = new_n1213_ & new_n6424_;
  assign new_n6508_ = new_n1216_ & new_n6424_;
  assign new_n6509_ = ~new_n6507_ & ~new_n6508_;
  assign new_n6510_ = ~new_n6506_ & new_n6509_;
  assign new_n6511_ = new_n6505_ & new_n6510_;
  assign new_n6512_ = new_n1223_ & new_n6424_;
  assign new_n6513_ = new_n1226_ & new_n6424_;
  assign new_n6514_ = new_n1229_ & new_n6424_;
  assign new_n6515_ = ~new_n6513_ & ~new_n6514_;
  assign new_n6516_ = ~new_n6512_ & new_n6515_;
  assign new_n6517_ = new_n1233_ & new_n6424_;
  assign new_n6518_ = new_n1235_ & new_n6424_;
  assign new_n6519_ = new_n1237_ & new_n6424_;
  assign new_n6520_ = ~new_n6518_ & ~new_n6519_;
  assign new_n6521_ = ~new_n6517_ & new_n6520_;
  assign new_n6522_ = new_n6516_ & new_n6521_;
  assign new_n6523_ = new_n6511_ & new_n6522_;
  assign new_n6524_ = ~A199 & ~A166;
  assign new_n6525_ = ~A167 & new_n6524_;
  assign new_n6526_ = new_n1727_ & new_n6525_;
  assign new_n6527_ = new_n1738_ & new_n6526_;
  assign new_n6528_ = new_n1243_ & new_n6424_;
  assign new_n6529_ = new_n1735_ & new_n6526_;
  assign new_n6530_ = ~new_n6528_ & ~new_n6529_;
  assign new_n6531_ = ~new_n6527_ & new_n6530_;
  assign new_n6532_ = A199 & ~A166;
  assign new_n6533_ = ~A167 & new_n6532_;
  assign new_n6534_ = new_n1743_ & new_n6533_;
  assign new_n6535_ = new_n1735_ & new_n6534_;
  assign new_n6536_ = new_n1725_ & new_n6526_;
  assign new_n6537_ = new_n1749_ & new_n6526_;
  assign new_n6538_ = ~new_n6536_ & ~new_n6537_;
  assign new_n6539_ = ~new_n6535_ & new_n6538_;
  assign new_n6540_ = new_n6531_ & new_n6539_;
  assign new_n6541_ = new_n1749_ & new_n6534_;
  assign new_n6542_ = new_n1738_ & new_n6534_;
  assign new_n6543_ = new_n1725_ & new_n6534_;
  assign new_n6544_ = ~new_n6542_ & ~new_n6543_;
  assign new_n6545_ = ~new_n6541_ & new_n6544_;
  assign new_n6546_ = ~A201 & ~A166;
  assign new_n6547_ = ~A167 & new_n6546_;
  assign new_n6548_ = new_n1757_ & new_n6547_;
  assign new_n6549_ = new_n1735_ & new_n6548_;
  assign new_n6550_ = new_n1738_ & new_n6548_;
  assign new_n6551_ = ~new_n6549_ & ~new_n6550_;
  assign new_n6552_ = new_n6545_ & new_n6551_;
  assign new_n6553_ = new_n6540_ & new_n6552_;
  assign new_n6554_ = new_n6523_ & new_n6553_;
  assign new_n6555_ = new_n1773_ & new_n6547_;
  assign new_n6556_ = new_n1735_ & new_n6555_;
  assign new_n6557_ = new_n1725_ & new_n6548_;
  assign new_n6558_ = new_n1749_ & new_n6548_;
  assign new_n6559_ = ~new_n6557_ & ~new_n6558_;
  assign new_n6560_ = ~new_n6556_ & new_n6559_;
  assign new_n6561_ = new_n1749_ & new_n6555_;
  assign new_n6562_ = new_n1738_ & new_n6555_;
  assign new_n6563_ = new_n1725_ & new_n6555_;
  assign new_n6564_ = ~new_n6562_ & ~new_n6563_;
  assign new_n6565_ = ~new_n6561_ & new_n6564_;
  assign new_n6566_ = new_n6560_ & new_n6565_;
  assign new_n6567_ = A201 & ~A166;
  assign new_n6568_ = ~A167 & new_n6567_;
  assign new_n6569_ = new_n1782_ & new_n6568_;
  assign new_n6570_ = new_n1725_ & new_n6569_;
  assign new_n6571_ = new_n1735_ & new_n6569_;
  assign new_n6572_ = new_n1738_ & new_n6569_;
  assign new_n6573_ = ~new_n6571_ & ~new_n6572_;
  assign new_n6574_ = ~new_n6570_ & new_n6573_;
  assign new_n6575_ = new_n1796_ & new_n6568_;
  assign new_n6576_ = new_n1738_ & new_n6575_;
  assign new_n6577_ = new_n1749_ & new_n6569_;
  assign new_n6578_ = new_n1735_ & new_n6575_;
  assign new_n6579_ = ~new_n6577_ & ~new_n6578_;
  assign new_n6580_ = ~new_n6576_ & new_n6579_;
  assign new_n6581_ = new_n6574_ & new_n6580_;
  assign new_n6582_ = new_n6566_ & new_n6581_;
  assign new_n6583_ = new_n1805_ & new_n6568_;
  assign new_n6584_ = new_n1735_ & new_n6583_;
  assign new_n6585_ = new_n1725_ & new_n6575_;
  assign new_n6586_ = new_n1749_ & new_n6575_;
  assign new_n6587_ = ~new_n6585_ & ~new_n6586_;
  assign new_n6588_ = ~new_n6584_ & new_n6587_;
  assign new_n6589_ = new_n1749_ & new_n6583_;
  assign new_n6590_ = new_n1738_ & new_n6583_;
  assign new_n6591_ = new_n1725_ & new_n6583_;
  assign new_n6592_ = ~new_n6590_ & ~new_n6591_;
  assign new_n6593_ = ~new_n6589_ & new_n6592_;
  assign new_n6594_ = new_n6588_ & new_n6593_;
  assign new_n6595_ = new_n1813_ & new_n6568_;
  assign new_n6596_ = new_n1725_ & new_n6595_;
  assign new_n6597_ = new_n1735_ & new_n6595_;
  assign new_n6598_ = new_n1738_ & new_n6595_;
  assign new_n6599_ = ~new_n6597_ & ~new_n6598_;
  assign new_n6600_ = ~new_n6596_ & new_n6599_;
  assign new_n6601_ = new_n1749_ & new_n6595_;
  assign new_n6602_ = new_n506_ & new_n6568_;
  assign new_n6603_ = new_n1830_ & new_n6602_;
  assign new_n6604_ = ~new_n6601_ & ~new_n6603_;
  assign new_n6605_ = new_n6600_ & new_n6604_;
  assign new_n6606_ = new_n6594_ & new_n6605_;
  assign new_n6607_ = new_n6582_ & new_n6606_;
  assign new_n6608_ = new_n6554_ & new_n6607_;
  assign new_n6609_ = new_n1840_ & new_n6602_;
  assign new_n6610_ = new_n1833_ & new_n6602_;
  assign new_n6611_ = new_n1827_ & new_n6602_;
  assign new_n6612_ = ~new_n6610_ & ~new_n6611_;
  assign new_n6613_ = ~new_n6609_ & new_n6612_;
  assign new_n6614_ = new_n1847_ & new_n6602_;
  assign new_n6615_ = new_n1842_ & new_n6602_;
  assign new_n6616_ = new_n1838_ & new_n6602_;
  assign new_n6617_ = ~new_n6615_ & ~new_n6616_;
  assign new_n6618_ = ~new_n6614_ & new_n6617_;
  assign new_n6619_ = new_n6613_ & new_n6618_;
  assign new_n6620_ = new_n1859_ & new_n6602_;
  assign new_n6621_ = new_n1849_ & new_n6602_;
  assign new_n6622_ = new_n1857_ & new_n6602_;
  assign new_n6623_ = ~new_n6621_ & ~new_n6622_;
  assign new_n6624_ = ~new_n6620_ & new_n6623_;
  assign new_n6625_ = new_n1868_ & new_n6602_;
  assign new_n6626_ = new_n1855_ & new_n6602_;
  assign new_n6627_ = new_n1866_ & new_n6602_;
  assign new_n6628_ = ~new_n6626_ & ~new_n6627_;
  assign new_n6629_ = ~new_n6625_ & new_n6628_;
  assign new_n6630_ = new_n6624_ & new_n6629_;
  assign new_n6631_ = new_n6619_ & new_n6630_;
  assign new_n6632_ = new_n1881_ & new_n6602_;
  assign new_n6633_ = new_n1864_ & new_n6602_;
  assign new_n6634_ = new_n1878_ & new_n6602_;
  assign new_n6635_ = ~new_n6633_ & ~new_n6634_;
  assign new_n6636_ = ~new_n6632_ & new_n6635_;
  assign new_n6637_ = new_n1892_ & new_n6602_;
  assign new_n6638_ = new_n1875_ & new_n6602_;
  assign new_n6639_ = new_n1889_ & new_n6602_;
  assign new_n6640_ = ~new_n6638_ & ~new_n6639_;
  assign new_n6641_ = ~new_n6637_ & new_n6640_;
  assign new_n6642_ = new_n6636_ & new_n6641_;
  assign new_n6643_ = new_n1902_ & new_n6602_;
  assign new_n6644_ = new_n1886_ & new_n6602_;
  assign new_n6645_ = new_n1900_ & new_n6602_;
  assign new_n6646_ = ~new_n6644_ & ~new_n6645_;
  assign new_n6647_ = ~new_n6643_ & new_n6646_;
  assign new_n6648_ = new_n1898_ & new_n6602_;
  assign new_n6649_ = new_n1913_ & new_n6602_;
  assign new_n6650_ = ~new_n6648_ & ~new_n6649_;
  assign new_n6651_ = new_n6647_ & new_n6650_;
  assign new_n6652_ = new_n6642_ & new_n6651_;
  assign new_n6653_ = new_n6631_ & new_n6652_;
  assign new_n6654_ = ~A199 & A166;
  assign new_n6655_ = A167 & new_n6654_;
  assign new_n6656_ = new_n1727_ & new_n6655_;
  assign new_n6657_ = new_n1725_ & new_n6656_;
  assign new_n6658_ = new_n1735_ & new_n6656_;
  assign new_n6659_ = new_n1738_ & new_n6656_;
  assign new_n6660_ = ~new_n6658_ & ~new_n6659_;
  assign new_n6661_ = ~new_n6657_ & new_n6660_;
  assign new_n6662_ = A199 & A166;
  assign new_n6663_ = A167 & new_n6662_;
  assign new_n6664_ = new_n1743_ & new_n6663_;
  assign new_n6665_ = new_n1738_ & new_n6664_;
  assign new_n6666_ = new_n1749_ & new_n6656_;
  assign new_n6667_ = new_n1735_ & new_n6664_;
  assign new_n6668_ = ~new_n6666_ & ~new_n6667_;
  assign new_n6669_ = ~new_n6665_ & new_n6668_;
  assign new_n6670_ = new_n6661_ & new_n6669_;
  assign new_n6671_ = ~A201 & A166;
  assign new_n6672_ = A167 & new_n6671_;
  assign new_n6673_ = new_n1757_ & new_n6672_;
  assign new_n6674_ = new_n1735_ & new_n6673_;
  assign new_n6675_ = new_n1725_ & new_n6664_;
  assign new_n6676_ = new_n1749_ & new_n6664_;
  assign new_n6677_ = ~new_n6675_ & ~new_n6676_;
  assign new_n6678_ = ~new_n6674_ & new_n6677_;
  assign new_n6679_ = new_n1749_ & new_n6673_;
  assign new_n6680_ = new_n1738_ & new_n6673_;
  assign new_n6681_ = new_n1725_ & new_n6673_;
  assign new_n6682_ = ~new_n6680_ & ~new_n6681_;
  assign new_n6683_ = ~new_n6679_ & new_n6682_;
  assign new_n6684_ = new_n6678_ & new_n6683_;
  assign new_n6685_ = new_n6670_ & new_n6684_;
  assign new_n6686_ = new_n1773_ & new_n6672_;
  assign new_n6687_ = new_n1725_ & new_n6686_;
  assign new_n6688_ = new_n1735_ & new_n6686_;
  assign new_n6689_ = new_n1738_ & new_n6686_;
  assign new_n6690_ = ~new_n6688_ & ~new_n6689_;
  assign new_n6691_ = ~new_n6687_ & new_n6690_;
  assign new_n6692_ = A201 & A166;
  assign new_n6693_ = A167 & new_n6692_;
  assign new_n6694_ = new_n1782_ & new_n6693_;
  assign new_n6695_ = new_n1738_ & new_n6694_;
  assign new_n6696_ = new_n1749_ & new_n6686_;
  assign new_n6697_ = new_n1735_ & new_n6694_;
  assign new_n6698_ = ~new_n6696_ & ~new_n6697_;
  assign new_n6699_ = ~new_n6695_ & new_n6698_;
  assign new_n6700_ = new_n6691_ & new_n6699_;
  assign new_n6701_ = new_n1796_ & new_n6693_;
  assign new_n6702_ = new_n1735_ & new_n6701_;
  assign new_n6703_ = new_n1725_ & new_n6694_;
  assign new_n6704_ = new_n1749_ & new_n6694_;
  assign new_n6705_ = ~new_n6703_ & ~new_n6704_;
  assign new_n6706_ = ~new_n6702_ & new_n6705_;
  assign new_n6707_ = new_n1738_ & new_n6701_;
  assign new_n6708_ = new_n1725_ & new_n6701_;
  assign new_n6709_ = ~new_n6707_ & ~new_n6708_;
  assign new_n6710_ = new_n6706_ & new_n6709_;
  assign new_n6711_ = new_n6700_ & new_n6710_;
  assign new_n6712_ = new_n6685_ & new_n6711_;
  assign new_n6713_ = new_n6653_ & new_n6712_;
  assign new_n6714_ = new_n6608_ & new_n6713_;
  assign new_n6715_ = new_n6500_ & new_n6714_;
  assign new_n6716_ = new_n6315_ & new_n6715_;
  assign new_n6717_ = new_n5940_ & new_n6716_;
  assign new_n6718_ = new_n5180_ & new_n6717_;
  assign new_n6719_ = new_n3452_ & new_n6718_;
  assign new_n6720_ = new_n1805_ & new_n6693_;
  assign new_n6721_ = new_n1738_ & new_n6720_;
  assign new_n6722_ = new_n1749_ & new_n6701_;
  assign new_n6723_ = new_n1735_ & new_n6720_;
  assign new_n6724_ = ~new_n6722_ & ~new_n6723_;
  assign new_n6725_ = ~new_n6721_ & new_n6724_;
  assign new_n6726_ = new_n1813_ & new_n6693_;
  assign new_n6727_ = new_n1735_ & new_n6726_;
  assign new_n6728_ = new_n1725_ & new_n6720_;
  assign new_n6729_ = new_n1749_ & new_n6720_;
  assign new_n6730_ = ~new_n6728_ & ~new_n6729_;
  assign new_n6731_ = ~new_n6727_ & new_n6730_;
  assign new_n6732_ = new_n6725_ & new_n6731_;
  assign new_n6733_ = new_n1749_ & new_n6726_;
  assign new_n6734_ = new_n1738_ & new_n6726_;
  assign new_n6735_ = new_n1725_ & new_n6726_;
  assign new_n6736_ = ~new_n6734_ & ~new_n6735_;
  assign new_n6737_ = ~new_n6733_ & new_n6736_;
  assign new_n6738_ = new_n506_ & new_n6693_;
  assign new_n6739_ = new_n1827_ & new_n6738_;
  assign new_n6740_ = new_n1830_ & new_n6738_;
  assign new_n6741_ = new_n1833_ & new_n6738_;
  assign new_n6742_ = ~new_n6740_ & ~new_n6741_;
  assign new_n6743_ = ~new_n6739_ & new_n6742_;
  assign new_n6744_ = new_n6737_ & new_n6743_;
  assign new_n6745_ = new_n6732_ & new_n6744_;
  assign new_n6746_ = new_n1838_ & new_n6738_;
  assign new_n6747_ = new_n1840_ & new_n6738_;
  assign new_n6748_ = new_n1842_ & new_n6738_;
  assign new_n6749_ = ~new_n6747_ & ~new_n6748_;
  assign new_n6750_ = ~new_n6746_ & new_n6749_;
  assign new_n6751_ = new_n1857_ & new_n6738_;
  assign new_n6752_ = new_n1847_ & new_n6738_;
  assign new_n6753_ = new_n1849_ & new_n6738_;
  assign new_n6754_ = ~new_n6752_ & ~new_n6753_;
  assign new_n6755_ = ~new_n6751_ & new_n6754_;
  assign new_n6756_ = new_n6750_ & new_n6755_;
  assign new_n6757_ = new_n1866_ & new_n6738_;
  assign new_n6758_ = new_n1859_ & new_n6738_;
  assign new_n6759_ = new_n1855_ & new_n6738_;
  assign new_n6760_ = ~new_n6758_ & ~new_n6759_;
  assign new_n6761_ = ~new_n6757_ & new_n6760_;
  assign new_n6762_ = new_n1878_ & new_n6738_;
  assign new_n6763_ = new_n1868_ & new_n6738_;
  assign new_n6764_ = new_n1864_ & new_n6738_;
  assign new_n6765_ = ~new_n6763_ & ~new_n6764_;
  assign new_n6766_ = ~new_n6762_ & new_n6765_;
  assign new_n6767_ = new_n6761_ & new_n6766_;
  assign new_n6768_ = new_n6756_ & new_n6767_;
  assign new_n6769_ = new_n6745_ & new_n6768_;
  assign new_n6770_ = new_n1889_ & new_n6738_;
  assign new_n6771_ = new_n1881_ & new_n6738_;
  assign new_n6772_ = new_n1875_ & new_n6738_;
  assign new_n6773_ = ~new_n6771_ & ~new_n6772_;
  assign new_n6774_ = ~new_n6770_ & new_n6773_;
  assign new_n6775_ = new_n1900_ & new_n6738_;
  assign new_n6776_ = new_n1892_ & new_n6738_;
  assign new_n6777_ = new_n1886_ & new_n6738_;
  assign new_n6778_ = ~new_n6776_ & ~new_n6777_;
  assign new_n6779_ = ~new_n6775_ & new_n6778_;
  assign new_n6780_ = new_n6774_ & new_n6779_;
  assign new_n6781_ = new_n1913_ & new_n6738_;
  assign new_n6782_ = new_n1902_ & new_n6738_;
  assign new_n6783_ = new_n1898_ & new_n6738_;
  assign new_n6784_ = ~new_n6782_ & ~new_n6783_;
  assign new_n6785_ = ~new_n6781_ & new_n6784_;
  assign new_n6786_ = new_n505_ & new_n516_;
  assign new_n6787_ = ~A201 & ~A200;
  assign new_n6788_ = A199 & new_n6787_;
  assign new_n6789_ = new_n6786_ & new_n6788_;
  assign new_n6790_ = new_n3662_ & new_n6789_;
  assign new_n6791_ = new_n3668_ & new_n6789_;
  assign new_n6792_ = new_n3670_ & new_n6789_;
  assign new_n6793_ = ~new_n6791_ & ~new_n6792_;
  assign new_n6794_ = ~new_n6790_ & new_n6793_;
  assign new_n6795_ = new_n6785_ & new_n6794_;
  assign new_n6796_ = new_n6780_ & new_n6795_;
  assign new_n6797_ = new_n3677_ & new_n6789_;
  assign new_n6798_ = new_n3679_ & new_n6789_;
  assign new_n6799_ = new_n3681_ & new_n6789_;
  assign new_n6800_ = ~new_n6798_ & ~new_n6799_;
  assign new_n6801_ = ~new_n6797_ & new_n6800_;
  assign new_n6802_ = new_n3685_ & new_n6789_;
  assign new_n6803_ = new_n3687_ & new_n6789_;
  assign new_n6804_ = new_n3689_ & new_n6789_;
  assign new_n6805_ = ~new_n6803_ & ~new_n6804_;
  assign new_n6806_ = ~new_n6802_ & new_n6805_;
  assign new_n6807_ = new_n6801_ & new_n6806_;
  assign new_n6808_ = new_n3694_ & new_n6789_;
  assign new_n6809_ = new_n3696_ & new_n6789_;
  assign new_n6810_ = new_n3698_ & new_n6789_;
  assign new_n6811_ = ~new_n6809_ & ~new_n6810_;
  assign new_n6812_ = ~new_n6808_ & new_n6811_;
  assign new_n6813_ = new_n3703_ & new_n6789_;
  assign new_n6814_ = new_n3705_ & new_n6789_;
  assign new_n6815_ = ~new_n6813_ & ~new_n6814_;
  assign new_n6816_ = new_n6812_ & new_n6815_;
  assign new_n6817_ = new_n6807_ & new_n6816_;
  assign new_n6818_ = new_n6796_ & new_n6817_;
  assign new_n6819_ = new_n6769_ & new_n6818_;
  assign new_n6820_ = new_n3711_ & new_n6789_;
  assign new_n6821_ = new_n3713_ & new_n6789_;
  assign new_n6822_ = new_n3715_ & new_n6789_;
  assign new_n6823_ = ~new_n6821_ & ~new_n6822_;
  assign new_n6824_ = ~new_n6820_ & new_n6823_;
  assign new_n6825_ = new_n3719_ & new_n6789_;
  assign new_n6826_ = new_n3721_ & new_n6789_;
  assign new_n6827_ = new_n3723_ & new_n6789_;
  assign new_n6828_ = ~new_n6826_ & ~new_n6827_;
  assign new_n6829_ = ~new_n6825_ & new_n6828_;
  assign new_n6830_ = new_n6824_ & new_n6829_;
  assign new_n6831_ = new_n3729_ & new_n6789_;
  assign new_n6832_ = new_n3731_ & new_n6789_;
  assign new_n6833_ = new_n3733_ & new_n6789_;
  assign new_n6834_ = ~new_n6832_ & ~new_n6833_;
  assign new_n6835_ = ~new_n6831_ & new_n6834_;
  assign new_n6836_ = new_n3738_ & new_n6789_;
  assign new_n6837_ = new_n3740_ & new_n6789_;
  assign new_n6838_ = new_n3742_ & new_n6789_;
  assign new_n6839_ = ~new_n6837_ & ~new_n6838_;
  assign new_n6840_ = ~new_n6836_ & new_n6839_;
  assign new_n6841_ = new_n6835_ & new_n6840_;
  assign new_n6842_ = new_n6830_ & new_n6841_;
  assign new_n6843_ = new_n3749_ & new_n6789_;
  assign new_n6844_ = new_n3751_ & new_n6789_;
  assign new_n6845_ = new_n3753_ & new_n6789_;
  assign new_n6846_ = ~new_n6844_ & ~new_n6845_;
  assign new_n6847_ = ~new_n6843_ & new_n6846_;
  assign new_n6848_ = new_n3757_ & new_n6789_;
  assign new_n6849_ = new_n3759_ & new_n6789_;
  assign new_n6850_ = new_n3761_ & new_n6789_;
  assign new_n6851_ = ~new_n6849_ & ~new_n6850_;
  assign new_n6852_ = ~new_n6848_ & new_n6851_;
  assign new_n6853_ = new_n6847_ & new_n6852_;
  assign new_n6854_ = new_n3767_ & new_n6789_;
  assign new_n6855_ = new_n3769_ & new_n6789_;
  assign new_n6856_ = new_n3771_ & new_n6789_;
  assign new_n6857_ = ~new_n6855_ & ~new_n6856_;
  assign new_n6858_ = ~new_n6854_ & new_n6857_;
  assign new_n6859_ = new_n3775_ & new_n6789_;
  assign new_n6860_ = new_n3778_ & new_n6789_;
  assign new_n6861_ = ~new_n6859_ & ~new_n6860_;
  assign new_n6862_ = new_n6858_ & new_n6861_;
  assign new_n6863_ = new_n6853_ & new_n6862_;
  assign new_n6864_ = new_n6842_ & new_n6863_;
  assign new_n6865_ = new_n3785_ & new_n6789_;
  assign new_n6866_ = new_n3787_ & new_n6789_;
  assign new_n6867_ = new_n3789_ & new_n6789_;
  assign new_n6868_ = ~new_n6866_ & ~new_n6867_;
  assign new_n6869_ = ~new_n6865_ & new_n6868_;
  assign new_n6870_ = new_n3793_ & new_n6789_;
  assign new_n6871_ = new_n3795_ & new_n6789_;
  assign new_n6872_ = new_n3797_ & new_n6789_;
  assign new_n6873_ = ~new_n6871_ & ~new_n6872_;
  assign new_n6874_ = ~new_n6870_ & new_n6873_;
  assign new_n6875_ = new_n6869_ & new_n6874_;
  assign new_n6876_ = new_n3803_ & new_n6789_;
  assign new_n6877_ = new_n3805_ & new_n6789_;
  assign new_n6878_ = new_n3807_ & new_n6789_;
  assign new_n6879_ = ~new_n6877_ & ~new_n6878_;
  assign new_n6880_ = ~new_n6876_ & new_n6879_;
  assign new_n6881_ = new_n3811_ & new_n6789_;
  assign new_n6882_ = new_n3813_ & new_n6789_;
  assign new_n6883_ = new_n3815_ & new_n6789_;
  assign new_n6884_ = ~new_n6882_ & ~new_n6883_;
  assign new_n6885_ = ~new_n6881_ & new_n6884_;
  assign new_n6886_ = new_n6880_ & new_n6885_;
  assign new_n6887_ = new_n6875_ & new_n6886_;
  assign new_n6888_ = new_n3821_ & new_n6789_;
  assign new_n6889_ = new_n3823_ & new_n6789_;
  assign new_n6890_ = new_n3825_ & new_n6789_;
  assign new_n6891_ = ~new_n6889_ & ~new_n6890_;
  assign new_n6892_ = ~new_n6888_ & new_n6891_;
  assign new_n6893_ = new_n3830_ & new_n6789_;
  assign new_n6894_ = new_n3832_ & new_n6789_;
  assign new_n6895_ = new_n3834_ & new_n6789_;
  assign new_n6896_ = ~new_n6894_ & ~new_n6895_;
  assign new_n6897_ = ~new_n6893_ & new_n6896_;
  assign new_n6898_ = new_n6892_ & new_n6897_;
  assign new_n6899_ = new_n3840_ & new_n6789_;
  assign new_n6900_ = new_n3842_ & new_n6789_;
  assign new_n6901_ = new_n3844_ & new_n6789_;
  assign new_n6902_ = ~new_n6900_ & ~new_n6901_;
  assign new_n6903_ = ~new_n6899_ & new_n6902_;
  assign new_n6904_ = new_n3848_ & new_n6789_;
  assign new_n6905_ = new_n3850_ & new_n6789_;
  assign new_n6906_ = ~new_n6904_ & ~new_n6905_;
  assign new_n6907_ = new_n6903_ & new_n6906_;
  assign new_n6908_ = new_n6898_ & new_n6907_;
  assign new_n6909_ = new_n6887_ & new_n6908_;
  assign new_n6910_ = new_n6864_ & new_n6909_;
  assign new_n6911_ = new_n6819_ & new_n6910_;
  assign new_n6912_ = new_n3857_ & new_n6789_;
  assign new_n6913_ = new_n3859_ & new_n6789_;
  assign new_n6914_ = new_n3861_ & new_n6789_;
  assign new_n6915_ = ~new_n6913_ & ~new_n6914_;
  assign new_n6916_ = ~new_n6912_ & new_n6915_;
  assign new_n6917_ = new_n505_ & new_n533_;
  assign new_n6918_ = new_n6788_ & new_n6917_;
  assign new_n6919_ = new_n3670_ & new_n6918_;
  assign new_n6920_ = new_n3868_ & new_n6789_;
  assign new_n6921_ = new_n3668_ & new_n6918_;
  assign new_n6922_ = ~new_n6920_ & ~new_n6921_;
  assign new_n6923_ = ~new_n6919_ & new_n6922_;
  assign new_n6924_ = new_n6916_ & new_n6923_;
  assign new_n6925_ = new_n3681_ & new_n6918_;
  assign new_n6926_ = new_n3662_ & new_n6918_;
  assign new_n6927_ = new_n3679_ & new_n6918_;
  assign new_n6928_ = ~new_n6926_ & ~new_n6927_;
  assign new_n6929_ = ~new_n6925_ & new_n6928_;
  assign new_n6930_ = new_n3689_ & new_n6918_;
  assign new_n6931_ = new_n3677_ & new_n6918_;
  assign new_n6932_ = new_n3687_ & new_n6918_;
  assign new_n6933_ = ~new_n6931_ & ~new_n6932_;
  assign new_n6934_ = ~new_n6930_ & new_n6933_;
  assign new_n6935_ = new_n6929_ & new_n6934_;
  assign new_n6936_ = new_n6924_ & new_n6935_;
  assign new_n6937_ = new_n3698_ & new_n6918_;
  assign new_n6938_ = new_n3685_ & new_n6918_;
  assign new_n6939_ = new_n3696_ & new_n6918_;
  assign new_n6940_ = ~new_n6938_ & ~new_n6939_;
  assign new_n6941_ = ~new_n6937_ & new_n6940_;
  assign new_n6942_ = new_n3705_ & new_n6918_;
  assign new_n6943_ = new_n3694_ & new_n6918_;
  assign new_n6944_ = new_n3703_ & new_n6918_;
  assign new_n6945_ = ~new_n6943_ & ~new_n6944_;
  assign new_n6946_ = ~new_n6942_ & new_n6945_;
  assign new_n6947_ = new_n6941_ & new_n6946_;
  assign new_n6948_ = new_n3711_ & new_n6918_;
  assign new_n6949_ = new_n3713_ & new_n6918_;
  assign new_n6950_ = new_n3715_ & new_n6918_;
  assign new_n6951_ = ~new_n6949_ & ~new_n6950_;
  assign new_n6952_ = ~new_n6948_ & new_n6951_;
  assign new_n6953_ = new_n3721_ & new_n6918_;
  assign new_n6954_ = new_n3723_ & new_n6918_;
  assign new_n6955_ = ~new_n6953_ & ~new_n6954_;
  assign new_n6956_ = new_n6952_ & new_n6955_;
  assign new_n6957_ = new_n6947_ & new_n6956_;
  assign new_n6958_ = new_n6936_ & new_n6957_;
  assign new_n6959_ = new_n3733_ & new_n6918_;
  assign new_n6960_ = new_n3719_ & new_n6918_;
  assign new_n6961_ = new_n3731_ & new_n6918_;
  assign new_n6962_ = ~new_n6960_ & ~new_n6961_;
  assign new_n6963_ = ~new_n6959_ & new_n6962_;
  assign new_n6964_ = new_n3742_ & new_n6918_;
  assign new_n6965_ = new_n3729_ & new_n6918_;
  assign new_n6966_ = new_n3740_ & new_n6918_;
  assign new_n6967_ = ~new_n6965_ & ~new_n6966_;
  assign new_n6968_ = ~new_n6964_ & new_n6967_;
  assign new_n6969_ = new_n6963_ & new_n6968_;
  assign new_n6970_ = new_n3753_ & new_n6918_;
  assign new_n6971_ = new_n3738_ & new_n6918_;
  assign new_n6972_ = new_n3751_ & new_n6918_;
  assign new_n6973_ = ~new_n6971_ & ~new_n6972_;
  assign new_n6974_ = ~new_n6970_ & new_n6973_;
  assign new_n6975_ = new_n3761_ & new_n6918_;
  assign new_n6976_ = new_n3749_ & new_n6918_;
  assign new_n6977_ = new_n3759_ & new_n6918_;
  assign new_n6978_ = ~new_n6976_ & ~new_n6977_;
  assign new_n6979_ = ~new_n6975_ & new_n6978_;
  assign new_n6980_ = new_n6974_ & new_n6979_;
  assign new_n6981_ = new_n6969_ & new_n6980_;
  assign new_n6982_ = new_n3771_ & new_n6918_;
  assign new_n6983_ = new_n3757_ & new_n6918_;
  assign new_n6984_ = new_n3769_ & new_n6918_;
  assign new_n6985_ = ~new_n6983_ & ~new_n6984_;
  assign new_n6986_ = ~new_n6982_ & new_n6985_;
  assign new_n6987_ = new_n3778_ & new_n6918_;
  assign new_n6988_ = new_n3767_ & new_n6918_;
  assign new_n6989_ = new_n3775_ & new_n6918_;
  assign new_n6990_ = ~new_n6988_ & ~new_n6989_;
  assign new_n6991_ = ~new_n6987_ & new_n6990_;
  assign new_n6992_ = new_n6986_ & new_n6991_;
  assign new_n6993_ = new_n3785_ & new_n6918_;
  assign new_n6994_ = new_n3787_ & new_n6918_;
  assign new_n6995_ = new_n3789_ & new_n6918_;
  assign new_n6996_ = ~new_n6994_ & ~new_n6995_;
  assign new_n6997_ = ~new_n6993_ & new_n6996_;
  assign new_n6998_ = new_n3795_ & new_n6918_;
  assign new_n6999_ = new_n3797_ & new_n6918_;
  assign new_n7000_ = ~new_n6998_ & ~new_n6999_;
  assign new_n7001_ = new_n6997_ & new_n7000_;
  assign new_n7002_ = new_n6992_ & new_n7001_;
  assign new_n7003_ = new_n6981_ & new_n7002_;
  assign new_n7004_ = new_n6958_ & new_n7003_;
  assign new_n7005_ = new_n3807_ & new_n6918_;
  assign new_n7006_ = new_n3793_ & new_n6918_;
  assign new_n7007_ = new_n3805_ & new_n6918_;
  assign new_n7008_ = ~new_n7006_ & ~new_n7007_;
  assign new_n7009_ = ~new_n7005_ & new_n7008_;
  assign new_n7010_ = new_n3815_ & new_n6918_;
  assign new_n7011_ = new_n3803_ & new_n6918_;
  assign new_n7012_ = new_n3813_ & new_n6918_;
  assign new_n7013_ = ~new_n7011_ & ~new_n7012_;
  assign new_n7014_ = ~new_n7010_ & new_n7013_;
  assign new_n7015_ = new_n7009_ & new_n7014_;
  assign new_n7016_ = new_n3825_ & new_n6918_;
  assign new_n7017_ = new_n3811_ & new_n6918_;
  assign new_n7018_ = new_n3823_ & new_n6918_;
  assign new_n7019_ = ~new_n7017_ & ~new_n7018_;
  assign new_n7020_ = ~new_n7016_ & new_n7019_;
  assign new_n7021_ = new_n3834_ & new_n6918_;
  assign new_n7022_ = new_n3821_ & new_n6918_;
  assign new_n7023_ = new_n3832_ & new_n6918_;
  assign new_n7024_ = ~new_n7022_ & ~new_n7023_;
  assign new_n7025_ = ~new_n7021_ & new_n7024_;
  assign new_n7026_ = new_n7020_ & new_n7025_;
  assign new_n7027_ = new_n7015_ & new_n7026_;
  assign new_n7028_ = new_n3844_ & new_n6918_;
  assign new_n7029_ = new_n3830_ & new_n6918_;
  assign new_n7030_ = new_n3842_ & new_n6918_;
  assign new_n7031_ = ~new_n7029_ & ~new_n7030_;
  assign new_n7032_ = ~new_n7028_ & new_n7031_;
  assign new_n7033_ = new_n3850_ & new_n6918_;
  assign new_n7034_ = new_n3840_ & new_n6918_;
  assign new_n7035_ = new_n3848_ & new_n6918_;
  assign new_n7036_ = ~new_n7034_ & ~new_n7035_;
  assign new_n7037_ = ~new_n7033_ & new_n7036_;
  assign new_n7038_ = new_n7032_ & new_n7037_;
  assign new_n7039_ = new_n3857_ & new_n6918_;
  assign new_n7040_ = new_n3859_ & new_n6918_;
  assign new_n7041_ = new_n3861_ & new_n6918_;
  assign new_n7042_ = ~new_n7040_ & ~new_n7041_;
  assign new_n7043_ = ~new_n7039_ & new_n7042_;
  assign new_n7044_ = new_n3868_ & new_n6918_;
  assign new_n7045_ = A232 & ~A203;
  assign new_n7046_ = new_n143_ & new_n7045_;
  assign new_n7047_ = A201 & ~A200;
  assign new_n7048_ = A199 & new_n7047_;
  assign new_n7049_ = new_n7046_ & new_n7048_;
  assign new_n7050_ = new_n951_ & new_n7049_;
  assign new_n7051_ = ~new_n7044_ & ~new_n7050_;
  assign new_n7052_ = new_n7043_ & new_n7051_;
  assign new_n7053_ = new_n7038_ & new_n7052_;
  assign new_n7054_ = new_n7027_ & new_n7053_;
  assign new_n7055_ = new_n964_ & new_n7049_;
  assign new_n7056_ = new_n954_ & new_n7049_;
  assign new_n7057_ = new_n948_ & new_n7049_;
  assign new_n7058_ = ~new_n7056_ & ~new_n7057_;
  assign new_n7059_ = ~new_n7055_ & new_n7058_;
  assign new_n7060_ = new_n975_ & new_n7049_;
  assign new_n7061_ = new_n967_ & new_n7049_;
  assign new_n7062_ = new_n961_ & new_n7049_;
  assign new_n7063_ = ~new_n7061_ & ~new_n7062_;
  assign new_n7064_ = ~new_n7060_ & new_n7063_;
  assign new_n7065_ = new_n7059_ & new_n7064_;
  assign new_n7066_ = new_n987_ & new_n7049_;
  assign new_n7067_ = new_n978_ & new_n7049_;
  assign new_n7068_ = new_n972_ & new_n7049_;
  assign new_n7069_ = ~new_n7067_ & ~new_n7068_;
  assign new_n7070_ = ~new_n7066_ & new_n7069_;
  assign new_n7071_ = new_n994_ & new_n7049_;
  assign new_n7072_ = new_n990_ & new_n7049_;
  assign new_n7073_ = new_n984_ & new_n7049_;
  assign new_n7074_ = ~new_n7072_ & ~new_n7073_;
  assign new_n7075_ = ~new_n7071_ & new_n7074_;
  assign new_n7076_ = new_n7070_ & new_n7075_;
  assign new_n7077_ = new_n7065_ & new_n7076_;
  assign new_n7078_ = new_n1010_ & new_n7049_;
  assign new_n7079_ = new_n996_ & new_n7049_;
  assign new_n7080_ = new_n1008_ & new_n7049_;
  assign new_n7081_ = ~new_n7079_ & ~new_n7080_;
  assign new_n7082_ = ~new_n7078_ & new_n7081_;
  assign new_n7083_ = new_n1018_ & new_n7049_;
  assign new_n7084_ = new_n1006_ & new_n7049_;
  assign new_n7085_ = new_n1016_ & new_n7049_;
  assign new_n7086_ = ~new_n7084_ & ~new_n7085_;
  assign new_n7087_ = ~new_n7083_ & new_n7086_;
  assign new_n7088_ = new_n7082_ & new_n7087_;
  assign new_n7089_ = new_n1027_ & new_n7049_;
  assign new_n7090_ = new_n1014_ & new_n7049_;
  assign new_n7091_ = new_n1025_ & new_n7049_;
  assign new_n7092_ = ~new_n7090_ & ~new_n7091_;
  assign new_n7093_ = ~new_n7089_ & new_n7092_;
  assign new_n7094_ = new_n1023_ & new_n7049_;
  assign new_n7095_ = new_n1033_ & new_n7049_;
  assign new_n7096_ = ~new_n7094_ & ~new_n7095_;
  assign new_n7097_ = new_n7093_ & new_n7096_;
  assign new_n7098_ = new_n7088_ & new_n7097_;
  assign new_n7099_ = new_n7077_ & new_n7098_;
  assign new_n7100_ = new_n7054_ & new_n7099_;
  assign new_n7101_ = new_n7004_ & new_n7100_;
  assign new_n7102_ = new_n6911_ & new_n7101_;
  assign new_n7103_ = new_n1043_ & new_n7049_;
  assign new_n7104_ = new_n1035_ & new_n7049_;
  assign new_n7105_ = new_n1031_ & new_n7049_;
  assign new_n7106_ = ~new_n7104_ & ~new_n7105_;
  assign new_n7107_ = ~new_n7103_ & new_n7106_;
  assign new_n7108_ = new_n1051_ & new_n7049_;
  assign new_n7109_ = new_n1045_ & new_n7049_;
  assign new_n7110_ = new_n1041_ & new_n7049_;
  assign new_n7111_ = ~new_n7109_ & ~new_n7110_;
  assign new_n7112_ = ~new_n7108_ & new_n7111_;
  assign new_n7113_ = new_n7107_ & new_n7112_;
  assign new_n7114_ = new_n264_ & new_n7045_;
  assign new_n7115_ = new_n7048_ & new_n7114_;
  assign new_n7116_ = new_n1065_ & new_n7115_;
  assign new_n7117_ = new_n1053_ & new_n7049_;
  assign new_n7118_ = new_n1049_ & new_n7049_;
  assign new_n7119_ = ~new_n7117_ & ~new_n7118_;
  assign new_n7120_ = ~new_n7116_ & new_n7119_;
  assign new_n7121_ = new_n1079_ & new_n7115_;
  assign new_n7122_ = new_n1071_ & new_n7115_;
  assign new_n7123_ = new_n1059_ & new_n7115_;
  assign new_n7124_ = ~new_n7122_ & ~new_n7123_;
  assign new_n7125_ = ~new_n7121_ & new_n7124_;
  assign new_n7126_ = new_n7120_ & new_n7125_;
  assign new_n7127_ = new_n7113_ & new_n7126_;
  assign new_n7128_ = new_n1095_ & new_n7115_;
  assign new_n7129_ = new_n1082_ & new_n7115_;
  assign new_n7130_ = new_n1076_ & new_n7115_;
  assign new_n7131_ = ~new_n7129_ & ~new_n7130_;
  assign new_n7132_ = ~new_n7128_ & new_n7131_;
  assign new_n7133_ = new_n1105_ & new_n7115_;
  assign new_n7134_ = new_n1099_ & new_n7115_;
  assign new_n7135_ = new_n1089_ & new_n7115_;
  assign new_n7136_ = ~new_n7134_ & ~new_n7135_;
  assign new_n7137_ = ~new_n7133_ & new_n7136_;
  assign new_n7138_ = new_n7132_ & new_n7137_;
  assign new_n7139_ = new_n1118_ & new_n7115_;
  assign new_n7140_ = new_n1107_ & new_n7115_;
  assign new_n7141_ = new_n1103_ & new_n7115_;
  assign new_n7142_ = ~new_n7140_ & ~new_n7141_;
  assign new_n7143_ = ~new_n7139_ & new_n7142_;
  assign new_n7144_ = new_n1131_ & new_n7115_;
  assign new_n7145_ = new_n1120_ & new_n7115_;
  assign new_n7146_ = new_n1114_ & new_n7115_;
  assign new_n7147_ = ~new_n7145_ & ~new_n7146_;
  assign new_n7148_ = ~new_n7144_ & new_n7147_;
  assign new_n7149_ = new_n7143_ & new_n7148_;
  assign new_n7150_ = new_n7138_ & new_n7149_;
  assign new_n7151_ = new_n7127_ & new_n7150_;
  assign new_n7152_ = new_n1145_ & new_n7115_;
  assign new_n7153_ = new_n1135_ & new_n7115_;
  assign new_n7154_ = new_n1127_ & new_n7115_;
  assign new_n7155_ = ~new_n7153_ & ~new_n7154_;
  assign new_n7156_ = ~new_n7152_ & new_n7155_;
  assign new_n7157_ = new_n1155_ & new_n7115_;
  assign new_n7158_ = new_n1149_ & new_n7115_;
  assign new_n7159_ = new_n1141_ & new_n7115_;
  assign new_n7160_ = ~new_n7158_ & ~new_n7159_;
  assign new_n7161_ = ~new_n7157_ & new_n7160_;
  assign new_n7162_ = new_n7156_ & new_n7161_;
  assign new_n7163_ = new_n1165_ & new_n7115_;
  assign new_n7164_ = new_n1157_ & new_n7115_;
  assign new_n7165_ = new_n1153_ & new_n7115_;
  assign new_n7166_ = ~new_n7164_ & ~new_n7165_;
  assign new_n7167_ = ~new_n7163_ & new_n7166_;
  assign new_n7168_ = new_n1172_ & new_n7115_;
  assign new_n7169_ = new_n1168_ & new_n7115_;
  assign new_n7170_ = new_n1162_ & new_n7115_;
  assign new_n7171_ = ~new_n7169_ & ~new_n7170_;
  assign new_n7172_ = ~new_n7168_ & new_n7171_;
  assign new_n7173_ = new_n7167_ & new_n7172_;
  assign new_n7174_ = new_n7162_ & new_n7173_;
  assign new_n7175_ = new_n1186_ & new_n7115_;
  assign new_n7176_ = new_n1174_ & new_n7115_;
  assign new_n7177_ = new_n1184_ & new_n7115_;
  assign new_n7178_ = ~new_n7176_ & ~new_n7177_;
  assign new_n7179_ = ~new_n7175_ & new_n7178_;
  assign new_n7180_ = new_n1194_ & new_n7115_;
  assign new_n7181_ = new_n1182_ & new_n7115_;
  assign new_n7182_ = new_n1192_ & new_n7115_;
  assign new_n7183_ = ~new_n7181_ & ~new_n7182_;
  assign new_n7184_ = ~new_n7180_ & new_n7183_;
  assign new_n7185_ = new_n7179_ & new_n7184_;
  assign new_n7186_ = new_n1204_ & new_n7115_;
  assign new_n7187_ = new_n1190_ & new_n7115_;
  assign new_n7188_ = new_n1202_ & new_n7115_;
  assign new_n7189_ = ~new_n7187_ & ~new_n7188_;
  assign new_n7190_ = ~new_n7186_ & new_n7189_;
  assign new_n7191_ = new_n1200_ & new_n7115_;
  assign new_n7192_ = new_n1213_ & new_n7115_;
  assign new_n7193_ = ~new_n7191_ & ~new_n7192_;
  assign new_n7194_ = new_n7190_ & new_n7193_;
  assign new_n7195_ = new_n7185_ & new_n7194_;
  assign new_n7196_ = new_n7174_ & new_n7195_;
  assign new_n7197_ = new_n7151_ & new_n7196_;
  assign new_n7198_ = new_n1226_ & new_n7115_;
  assign new_n7199_ = new_n1216_ & new_n7115_;
  assign new_n7200_ = new_n1210_ & new_n7115_;
  assign new_n7201_ = ~new_n7199_ & ~new_n7200_;
  assign new_n7202_ = ~new_n7198_ & new_n7201_;
  assign new_n7203_ = new_n1235_ & new_n7115_;
  assign new_n7204_ = new_n1229_ & new_n7115_;
  assign new_n7205_ = new_n1223_ & new_n7115_;
  assign new_n7206_ = ~new_n7204_ & ~new_n7205_;
  assign new_n7207_ = ~new_n7203_ & new_n7206_;
  assign new_n7208_ = new_n7202_ & new_n7207_;
  assign new_n7209_ = new_n1243_ & new_n7115_;
  assign new_n7210_ = new_n1237_ & new_n7115_;
  assign new_n7211_ = new_n1233_ & new_n7115_;
  assign new_n7212_ = ~new_n7210_ & ~new_n7211_;
  assign new_n7213_ = ~new_n7209_ & new_n7212_;
  assign new_n7214_ = ~A232 & ~A203;
  assign new_n7215_ = new_n292_ & new_n7214_;
  assign new_n7216_ = new_n7048_ & new_n7215_;
  assign new_n7217_ = new_n948_ & new_n7216_;
  assign new_n7218_ = new_n951_ & new_n7216_;
  assign new_n7219_ = new_n954_ & new_n7216_;
  assign new_n7220_ = ~new_n7218_ & ~new_n7219_;
  assign new_n7221_ = ~new_n7217_ & new_n7220_;
  assign new_n7222_ = new_n7213_ & new_n7221_;
  assign new_n7223_ = new_n7208_ & new_n7222_;
  assign new_n7224_ = new_n961_ & new_n7216_;
  assign new_n7225_ = new_n964_ & new_n7216_;
  assign new_n7226_ = new_n967_ & new_n7216_;
  assign new_n7227_ = ~new_n7225_ & ~new_n7226_;
  assign new_n7228_ = ~new_n7224_ & new_n7227_;
  assign new_n7229_ = new_n972_ & new_n7216_;
  assign new_n7230_ = new_n975_ & new_n7216_;
  assign new_n7231_ = new_n978_ & new_n7216_;
  assign new_n7232_ = ~new_n7230_ & ~new_n7231_;
  assign new_n7233_ = ~new_n7229_ & new_n7232_;
  assign new_n7234_ = new_n7228_ & new_n7233_;
  assign new_n7235_ = new_n984_ & new_n7216_;
  assign new_n7236_ = new_n987_ & new_n7216_;
  assign new_n7237_ = new_n990_ & new_n7216_;
  assign new_n7238_ = ~new_n7236_ & ~new_n7237_;
  assign new_n7239_ = ~new_n7235_ & new_n7238_;
  assign new_n7240_ = new_n994_ & new_n7216_;
  assign new_n7241_ = new_n996_ & new_n7216_;
  assign new_n7242_ = ~new_n7240_ & ~new_n7241_;
  assign new_n7243_ = new_n7239_ & new_n7242_;
  assign new_n7244_ = new_n7234_ & new_n7243_;
  assign new_n7245_ = new_n7223_ & new_n7244_;
  assign new_n7246_ = new_n1006_ & new_n7216_;
  assign new_n7247_ = new_n1008_ & new_n7216_;
  assign new_n7248_ = new_n1010_ & new_n7216_;
  assign new_n7249_ = ~new_n7247_ & ~new_n7248_;
  assign new_n7250_ = ~new_n7246_ & new_n7249_;
  assign new_n7251_ = new_n1014_ & new_n7216_;
  assign new_n7252_ = new_n1016_ & new_n7216_;
  assign new_n7253_ = new_n1018_ & new_n7216_;
  assign new_n7254_ = ~new_n7252_ & ~new_n7253_;
  assign new_n7255_ = ~new_n7251_ & new_n7254_;
  assign new_n7256_ = new_n7250_ & new_n7255_;
  assign new_n7257_ = new_n1023_ & new_n7216_;
  assign new_n7258_ = new_n1025_ & new_n7216_;
  assign new_n7259_ = new_n1027_ & new_n7216_;
  assign new_n7260_ = ~new_n7258_ & ~new_n7259_;
  assign new_n7261_ = ~new_n7257_ & new_n7260_;
  assign new_n7262_ = new_n1031_ & new_n7216_;
  assign new_n7263_ = new_n1033_ & new_n7216_;
  assign new_n7264_ = new_n1035_ & new_n7216_;
  assign new_n7265_ = ~new_n7263_ & ~new_n7264_;
  assign new_n7266_ = ~new_n7262_ & new_n7265_;
  assign new_n7267_ = new_n7261_ & new_n7266_;
  assign new_n7268_ = new_n7256_ & new_n7267_;
  assign new_n7269_ = new_n1041_ & new_n7216_;
  assign new_n7270_ = new_n1043_ & new_n7216_;
  assign new_n7271_ = new_n1045_ & new_n7216_;
  assign new_n7272_ = ~new_n7270_ & ~new_n7271_;
  assign new_n7273_ = ~new_n7269_ & new_n7272_;
  assign new_n7274_ = new_n1049_ & new_n7216_;
  assign new_n7275_ = new_n1051_ & new_n7216_;
  assign new_n7276_ = new_n1053_ & new_n7216_;
  assign new_n7277_ = ~new_n7275_ & ~new_n7276_;
  assign new_n7278_ = ~new_n7274_ & new_n7277_;
  assign new_n7279_ = new_n7273_ & new_n7278_;
  assign new_n7280_ = new_n350_ & new_n7214_;
  assign new_n7281_ = new_n7048_ & new_n7280_;
  assign new_n7282_ = new_n1059_ & new_n7281_;
  assign new_n7283_ = new_n1065_ & new_n7281_;
  assign new_n7284_ = new_n1071_ & new_n7281_;
  assign new_n7285_ = ~new_n7283_ & ~new_n7284_;
  assign new_n7286_ = ~new_n7282_ & new_n7285_;
  assign new_n7287_ = new_n1079_ & new_n7281_;
  assign new_n7288_ = new_n1082_ & new_n7281_;
  assign new_n7289_ = ~new_n7287_ & ~new_n7288_;
  assign new_n7290_ = new_n7286_ & new_n7289_;
  assign new_n7291_ = new_n7279_ & new_n7290_;
  assign new_n7292_ = new_n7268_ & new_n7291_;
  assign new_n7293_ = new_n7245_ & new_n7292_;
  assign new_n7294_ = new_n7197_ & new_n7293_;
  assign new_n7295_ = new_n1099_ & new_n7281_;
  assign new_n7296_ = new_n1076_ & new_n7281_;
  assign new_n7297_ = new_n1095_ & new_n7281_;
  assign new_n7298_ = ~new_n7296_ & ~new_n7297_;
  assign new_n7299_ = ~new_n7295_ & new_n7298_;
  assign new_n7300_ = new_n1107_ & new_n7281_;
  assign new_n7301_ = new_n1089_ & new_n7281_;
  assign new_n7302_ = new_n1105_ & new_n7281_;
  assign new_n7303_ = ~new_n7301_ & ~new_n7302_;
  assign new_n7304_ = ~new_n7300_ & new_n7303_;
  assign new_n7305_ = new_n7299_ & new_n7304_;
  assign new_n7306_ = new_n1120_ & new_n7281_;
  assign new_n7307_ = new_n1103_ & new_n7281_;
  assign new_n7308_ = new_n1118_ & new_n7281_;
  assign new_n7309_ = ~new_n7307_ & ~new_n7308_;
  assign new_n7310_ = ~new_n7306_ & new_n7309_;
  assign new_n7311_ = new_n1135_ & new_n7281_;
  assign new_n7312_ = new_n1114_ & new_n7281_;
  assign new_n7313_ = new_n1131_ & new_n7281_;
  assign new_n7314_ = ~new_n7312_ & ~new_n7313_;
  assign new_n7315_ = ~new_n7311_ & new_n7314_;
  assign new_n7316_ = new_n7310_ & new_n7315_;
  assign new_n7317_ = new_n7305_ & new_n7316_;
  assign new_n7318_ = new_n1149_ & new_n7281_;
  assign new_n7319_ = new_n1127_ & new_n7281_;
  assign new_n7320_ = new_n1145_ & new_n7281_;
  assign new_n7321_ = ~new_n7319_ & ~new_n7320_;
  assign new_n7322_ = ~new_n7318_ & new_n7321_;
  assign new_n7323_ = new_n1157_ & new_n7281_;
  assign new_n7324_ = new_n1141_ & new_n7281_;
  assign new_n7325_ = new_n1155_ & new_n7281_;
  assign new_n7326_ = ~new_n7324_ & ~new_n7325_;
  assign new_n7327_ = ~new_n7323_ & new_n7326_;
  assign new_n7328_ = new_n7322_ & new_n7327_;
  assign new_n7329_ = new_n1168_ & new_n7281_;
  assign new_n7330_ = new_n1153_ & new_n7281_;
  assign new_n7331_ = new_n1165_ & new_n7281_;
  assign new_n7332_ = ~new_n7330_ & ~new_n7331_;
  assign new_n7333_ = ~new_n7329_ & new_n7332_;
  assign new_n7334_ = new_n1162_ & new_n7281_;
  assign new_n7335_ = new_n1172_ & new_n7281_;
  assign new_n7336_ = ~new_n7334_ & ~new_n7335_;
  assign new_n7337_ = new_n7333_ & new_n7336_;
  assign new_n7338_ = new_n7328_ & new_n7337_;
  assign new_n7339_ = new_n7317_ & new_n7338_;
  assign new_n7340_ = new_n1186_ & new_n7281_;
  assign new_n7341_ = new_n1174_ & new_n7281_;
  assign new_n7342_ = new_n1184_ & new_n7281_;
  assign new_n7343_ = ~new_n7341_ & ~new_n7342_;
  assign new_n7344_ = ~new_n7340_ & new_n7343_;
  assign new_n7345_ = new_n1194_ & new_n7281_;
  assign new_n7346_ = new_n1182_ & new_n7281_;
  assign new_n7347_ = new_n1192_ & new_n7281_;
  assign new_n7348_ = ~new_n7346_ & ~new_n7347_;
  assign new_n7349_ = ~new_n7345_ & new_n7348_;
  assign new_n7350_ = new_n7344_ & new_n7349_;
  assign new_n7351_ = new_n1204_ & new_n7281_;
  assign new_n7352_ = new_n1190_ & new_n7281_;
  assign new_n7353_ = new_n1202_ & new_n7281_;
  assign new_n7354_ = ~new_n7352_ & ~new_n7353_;
  assign new_n7355_ = ~new_n7351_ & new_n7354_;
  assign new_n7356_ = new_n1216_ & new_n7281_;
  assign new_n7357_ = new_n1200_ & new_n7281_;
  assign new_n7358_ = new_n1213_ & new_n7281_;
  assign new_n7359_ = ~new_n7357_ & ~new_n7358_;
  assign new_n7360_ = ~new_n7356_ & new_n7359_;
  assign new_n7361_ = new_n7355_ & new_n7360_;
  assign new_n7362_ = new_n7350_ & new_n7361_;
  assign new_n7363_ = new_n1229_ & new_n7281_;
  assign new_n7364_ = new_n1210_ & new_n7281_;
  assign new_n7365_ = new_n1226_ & new_n7281_;
  assign new_n7366_ = ~new_n7364_ & ~new_n7365_;
  assign new_n7367_ = ~new_n7363_ & new_n7366_;
  assign new_n7368_ = new_n1237_ & new_n7281_;
  assign new_n7369_ = new_n1223_ & new_n7281_;
  assign new_n7370_ = new_n1235_ & new_n7281_;
  assign new_n7371_ = ~new_n7369_ & ~new_n7370_;
  assign new_n7372_ = ~new_n7368_ & new_n7371_;
  assign new_n7373_ = new_n7367_ & new_n7372_;
  assign new_n7374_ = A232 & A202;
  assign new_n7375_ = new_n143_ & new_n7374_;
  assign new_n7376_ = new_n7048_ & new_n7375_;
  assign new_n7377_ = new_n951_ & new_n7376_;
  assign new_n7378_ = new_n1233_ & new_n7281_;
  assign new_n7379_ = new_n1243_ & new_n7281_;
  assign new_n7380_ = ~new_n7378_ & ~new_n7379_;
  assign new_n7381_ = ~new_n7377_ & new_n7380_;
  assign new_n7382_ = new_n954_ & new_n7376_;
  assign new_n7383_ = new_n948_ & new_n7376_;
  assign new_n7384_ = ~new_n7382_ & ~new_n7383_;
  assign new_n7385_ = new_n7381_ & new_n7384_;
  assign new_n7386_ = new_n7373_ & new_n7385_;
  assign new_n7387_ = new_n7362_ & new_n7386_;
  assign new_n7388_ = new_n7339_ & new_n7387_;
  assign new_n7389_ = new_n961_ & new_n7376_;
  assign new_n7390_ = new_n964_ & new_n7376_;
  assign new_n7391_ = new_n967_ & new_n7376_;
  assign new_n7392_ = ~new_n7390_ & ~new_n7391_;
  assign new_n7393_ = ~new_n7389_ & new_n7392_;
  assign new_n7394_ = new_n972_ & new_n7376_;
  assign new_n7395_ = new_n975_ & new_n7376_;
  assign new_n7396_ = new_n978_ & new_n7376_;
  assign new_n7397_ = ~new_n7395_ & ~new_n7396_;
  assign new_n7398_ = ~new_n7394_ & new_n7397_;
  assign new_n7399_ = new_n7393_ & new_n7398_;
  assign new_n7400_ = new_n984_ & new_n7376_;
  assign new_n7401_ = new_n987_ & new_n7376_;
  assign new_n7402_ = new_n990_ & new_n7376_;
  assign new_n7403_ = ~new_n7401_ & ~new_n7402_;
  assign new_n7404_ = ~new_n7400_ & new_n7403_;
  assign new_n7405_ = new_n1008_ & new_n7376_;
  assign new_n7406_ = new_n994_ & new_n7376_;
  assign new_n7407_ = new_n996_ & new_n7376_;
  assign new_n7408_ = ~new_n7406_ & ~new_n7407_;
  assign new_n7409_ = ~new_n7405_ & new_n7408_;
  assign new_n7410_ = new_n7404_ & new_n7409_;
  assign new_n7411_ = new_n7399_ & new_n7410_;
  assign new_n7412_ = new_n1016_ & new_n7376_;
  assign new_n7413_ = new_n1010_ & new_n7376_;
  assign new_n7414_ = new_n1006_ & new_n7376_;
  assign new_n7415_ = ~new_n7413_ & ~new_n7414_;
  assign new_n7416_ = ~new_n7412_ & new_n7415_;
  assign new_n7417_ = new_n1025_ & new_n7376_;
  assign new_n7418_ = new_n1018_ & new_n7376_;
  assign new_n7419_ = new_n1014_ & new_n7376_;
  assign new_n7420_ = ~new_n7418_ & ~new_n7419_;
  assign new_n7421_ = ~new_n7417_ & new_n7420_;
  assign new_n7422_ = new_n7416_ & new_n7421_;
  assign new_n7423_ = new_n1033_ & new_n7376_;
  assign new_n7424_ = new_n1027_ & new_n7376_;
  assign new_n7425_ = new_n1023_ & new_n7376_;
  assign new_n7426_ = ~new_n7424_ & ~new_n7425_;
  assign new_n7427_ = ~new_n7423_ & new_n7426_;
  assign new_n7428_ = new_n1035_ & new_n7376_;
  assign new_n7429_ = new_n1031_ & new_n7376_;
  assign new_n7430_ = ~new_n7428_ & ~new_n7429_;
  assign new_n7431_ = new_n7427_ & new_n7430_;
  assign new_n7432_ = new_n7422_ & new_n7431_;
  assign new_n7433_ = new_n7411_ & new_n7432_;
  assign new_n7434_ = new_n1041_ & new_n7376_;
  assign new_n7435_ = new_n1043_ & new_n7376_;
  assign new_n7436_ = new_n1045_ & new_n7376_;
  assign new_n7437_ = ~new_n7435_ & ~new_n7436_;
  assign new_n7438_ = ~new_n7434_ & new_n7437_;
  assign new_n7439_ = new_n1049_ & new_n7376_;
  assign new_n7440_ = new_n1051_ & new_n7376_;
  assign new_n7441_ = new_n1053_ & new_n7376_;
  assign new_n7442_ = ~new_n7440_ & ~new_n7441_;
  assign new_n7443_ = ~new_n7439_ & new_n7442_;
  assign new_n7444_ = new_n7438_ & new_n7443_;
  assign new_n7445_ = new_n264_ & new_n7374_;
  assign new_n7446_ = new_n7048_ & new_n7445_;
  assign new_n7447_ = new_n1059_ & new_n7446_;
  assign new_n7448_ = new_n1065_ & new_n7446_;
  assign new_n7449_ = new_n1071_ & new_n7446_;
  assign new_n7450_ = ~new_n7448_ & ~new_n7449_;
  assign new_n7451_ = ~new_n7447_ & new_n7450_;
  assign new_n7452_ = new_n1076_ & new_n7446_;
  assign new_n7453_ = new_n1079_ & new_n7446_;
  assign new_n7454_ = new_n1082_ & new_n7446_;
  assign new_n7455_ = ~new_n7453_ & ~new_n7454_;
  assign new_n7456_ = ~new_n7452_ & new_n7455_;
  assign new_n7457_ = new_n7451_ & new_n7456_;
  assign new_n7458_ = new_n7444_ & new_n7457_;
  assign new_n7459_ = new_n1089_ & new_n7446_;
  assign new_n7460_ = new_n1095_ & new_n7446_;
  assign new_n7461_ = new_n1099_ & new_n7446_;
  assign new_n7462_ = ~new_n7460_ & ~new_n7461_;
  assign new_n7463_ = ~new_n7459_ & new_n7462_;
  assign new_n7464_ = new_n1103_ & new_n7446_;
  assign new_n7465_ = new_n1105_ & new_n7446_;
  assign new_n7466_ = new_n1107_ & new_n7446_;
  assign new_n7467_ = ~new_n7465_ & ~new_n7466_;
  assign new_n7468_ = ~new_n7464_ & new_n7467_;
  assign new_n7469_ = new_n7463_ & new_n7468_;
  assign new_n7470_ = new_n1114_ & new_n7446_;
  assign new_n7471_ = new_n1118_ & new_n7446_;
  assign new_n7472_ = new_n1120_ & new_n7446_;
  assign new_n7473_ = ~new_n7471_ & ~new_n7472_;
  assign new_n7474_ = ~new_n7470_ & new_n7473_;
  assign new_n7475_ = new_n1131_ & new_n7446_;
  assign new_n7476_ = new_n1135_ & new_n7446_;
  assign new_n7477_ = ~new_n7475_ & ~new_n7476_;
  assign new_n7478_ = new_n7474_ & new_n7477_;
  assign new_n7479_ = new_n7469_ & new_n7478_;
  assign new_n7480_ = new_n7458_ & new_n7479_;
  assign new_n7481_ = new_n7433_ & new_n7480_;
  assign new_n7482_ = new_n7388_ & new_n7481_;
  assign new_n7483_ = new_n7294_ & new_n7482_;
  assign new_n7484_ = new_n7102_ & new_n7483_;
  assign new_n7485_ = new_n1149_ & new_n7446_;
  assign new_n7486_ = new_n1127_ & new_n7446_;
  assign new_n7487_ = new_n1145_ & new_n7446_;
  assign new_n7488_ = ~new_n7486_ & ~new_n7487_;
  assign new_n7489_ = ~new_n7485_ & new_n7488_;
  assign new_n7490_ = new_n1157_ & new_n7446_;
  assign new_n7491_ = new_n1141_ & new_n7446_;
  assign new_n7492_ = new_n1155_ & new_n7446_;
  assign new_n7493_ = ~new_n7491_ & ~new_n7492_;
  assign new_n7494_ = ~new_n7490_ & new_n7493_;
  assign new_n7495_ = new_n7489_ & new_n7494_;
  assign new_n7496_ = new_n1168_ & new_n7446_;
  assign new_n7497_ = new_n1153_ & new_n7446_;
  assign new_n7498_ = new_n1165_ & new_n7446_;
  assign new_n7499_ = ~new_n7497_ & ~new_n7498_;
  assign new_n7500_ = ~new_n7496_ & new_n7499_;
  assign new_n7501_ = new_n1174_ & new_n7446_;
  assign new_n7502_ = new_n1162_ & new_n7446_;
  assign new_n7503_ = new_n1172_ & new_n7446_;
  assign new_n7504_ = ~new_n7502_ & ~new_n7503_;
  assign new_n7505_ = ~new_n7501_ & new_n7504_;
  assign new_n7506_ = new_n7500_ & new_n7505_;
  assign new_n7507_ = new_n7495_ & new_n7506_;
  assign new_n7508_ = new_n1182_ & new_n7446_;
  assign new_n7509_ = new_n1184_ & new_n7446_;
  assign new_n7510_ = new_n1186_ & new_n7446_;
  assign new_n7511_ = ~new_n7509_ & ~new_n7510_;
  assign new_n7512_ = ~new_n7508_ & new_n7511_;
  assign new_n7513_ = new_n1190_ & new_n7446_;
  assign new_n7514_ = new_n1192_ & new_n7446_;
  assign new_n7515_ = new_n1194_ & new_n7446_;
  assign new_n7516_ = ~new_n7514_ & ~new_n7515_;
  assign new_n7517_ = ~new_n7513_ & new_n7516_;
  assign new_n7518_ = new_n7512_ & new_n7517_;
  assign new_n7519_ = new_n1200_ & new_n7446_;
  assign new_n7520_ = new_n1202_ & new_n7446_;
  assign new_n7521_ = new_n1204_ & new_n7446_;
  assign new_n7522_ = ~new_n7520_ & ~new_n7521_;
  assign new_n7523_ = ~new_n7519_ & new_n7522_;
  assign new_n7524_ = new_n1210_ & new_n7446_;
  assign new_n7525_ = new_n1213_ & new_n7446_;
  assign new_n7526_ = new_n1216_ & new_n7446_;
  assign new_n7527_ = ~new_n7525_ & ~new_n7526_;
  assign new_n7528_ = ~new_n7524_ & new_n7527_;
  assign new_n7529_ = new_n7523_ & new_n7528_;
  assign new_n7530_ = new_n7518_ & new_n7529_;
  assign new_n7531_ = new_n7507_ & new_n7530_;
  assign new_n7532_ = new_n1223_ & new_n7446_;
  assign new_n7533_ = new_n1226_ & new_n7446_;
  assign new_n7534_ = new_n1229_ & new_n7446_;
  assign new_n7535_ = ~new_n7533_ & ~new_n7534_;
  assign new_n7536_ = ~new_n7532_ & new_n7535_;
  assign new_n7537_ = new_n1233_ & new_n7446_;
  assign new_n7538_ = new_n1235_ & new_n7446_;
  assign new_n7539_ = new_n1237_ & new_n7446_;
  assign new_n7540_ = ~new_n7538_ & ~new_n7539_;
  assign new_n7541_ = ~new_n7537_ & new_n7540_;
  assign new_n7542_ = new_n7536_ & new_n7541_;
  assign new_n7543_ = ~A232 & A202;
  assign new_n7544_ = new_n292_ & new_n7543_;
  assign new_n7545_ = new_n7048_ & new_n7544_;
  assign new_n7546_ = new_n954_ & new_n7545_;
  assign new_n7547_ = new_n1243_ & new_n7446_;
  assign new_n7548_ = new_n951_ & new_n7545_;
  assign new_n7549_ = ~new_n7547_ & ~new_n7548_;
  assign new_n7550_ = ~new_n7546_ & new_n7549_;
  assign new_n7551_ = new_n967_ & new_n7545_;
  assign new_n7552_ = new_n948_ & new_n7545_;
  assign new_n7553_ = new_n964_ & new_n7545_;
  assign new_n7554_ = ~new_n7552_ & ~new_n7553_;
  assign new_n7555_ = ~new_n7551_ & new_n7554_;
  assign new_n7556_ = new_n7550_ & new_n7555_;
  assign new_n7557_ = new_n7542_ & new_n7556_;
  assign new_n7558_ = new_n978_ & new_n7545_;
  assign new_n7559_ = new_n961_ & new_n7545_;
  assign new_n7560_ = new_n975_ & new_n7545_;
  assign new_n7561_ = ~new_n7559_ & ~new_n7560_;
  assign new_n7562_ = ~new_n7558_ & new_n7561_;
  assign new_n7563_ = new_n990_ & new_n7545_;
  assign new_n7564_ = new_n972_ & new_n7545_;
  assign new_n7565_ = new_n987_ & new_n7545_;
  assign new_n7566_ = ~new_n7564_ & ~new_n7565_;
  assign new_n7567_ = ~new_n7563_ & new_n7566_;
  assign new_n7568_ = new_n7562_ & new_n7567_;
  assign new_n7569_ = new_n996_ & new_n7545_;
  assign new_n7570_ = new_n984_ & new_n7545_;
  assign new_n7571_ = new_n994_ & new_n7545_;
  assign new_n7572_ = ~new_n7570_ & ~new_n7571_;
  assign new_n7573_ = ~new_n7569_ & new_n7572_;
  assign new_n7574_ = new_n1008_ & new_n7545_;
  assign new_n7575_ = new_n1010_ & new_n7545_;
  assign new_n7576_ = ~new_n7574_ & ~new_n7575_;
  assign new_n7577_ = new_n7573_ & new_n7576_;
  assign new_n7578_ = new_n7568_ & new_n7577_;
  assign new_n7579_ = new_n7557_ & new_n7578_;
  assign new_n7580_ = new_n7531_ & new_n7579_;
  assign new_n7581_ = new_n1018_ & new_n7545_;
  assign new_n7582_ = new_n1006_ & new_n7545_;
  assign new_n7583_ = new_n1016_ & new_n7545_;
  assign new_n7584_ = ~new_n7582_ & ~new_n7583_;
  assign new_n7585_ = ~new_n7581_ & new_n7584_;
  assign new_n7586_ = new_n1027_ & new_n7545_;
  assign new_n7587_ = new_n1014_ & new_n7545_;
  assign new_n7588_ = new_n1025_ & new_n7545_;
  assign new_n7589_ = ~new_n7587_ & ~new_n7588_;
  assign new_n7590_ = ~new_n7586_ & new_n7589_;
  assign new_n7591_ = new_n7585_ & new_n7590_;
  assign new_n7592_ = new_n1035_ & new_n7545_;
  assign new_n7593_ = new_n1023_ & new_n7545_;
  assign new_n7594_ = new_n1033_ & new_n7545_;
  assign new_n7595_ = ~new_n7593_ & ~new_n7594_;
  assign new_n7596_ = ~new_n7592_ & new_n7595_;
  assign new_n7597_ = new_n1045_ & new_n7545_;
  assign new_n7598_ = new_n1031_ & new_n7545_;
  assign new_n7599_ = new_n1043_ & new_n7545_;
  assign new_n7600_ = ~new_n7598_ & ~new_n7599_;
  assign new_n7601_ = ~new_n7597_ & new_n7600_;
  assign new_n7602_ = new_n7596_ & new_n7601_;
  assign new_n7603_ = new_n7591_ & new_n7602_;
  assign new_n7604_ = new_n1053_ & new_n7545_;
  assign new_n7605_ = new_n1041_ & new_n7545_;
  assign new_n7606_ = new_n1051_ & new_n7545_;
  assign new_n7607_ = ~new_n7605_ & ~new_n7606_;
  assign new_n7608_ = ~new_n7604_ & new_n7607_;
  assign new_n7609_ = new_n350_ & new_n7543_;
  assign new_n7610_ = new_n7048_ & new_n7609_;
  assign new_n7611_ = new_n1071_ & new_n7610_;
  assign new_n7612_ = new_n1049_ & new_n7545_;
  assign new_n7613_ = new_n1065_ & new_n7610_;
  assign new_n7614_ = ~new_n7612_ & ~new_n7613_;
  assign new_n7615_ = ~new_n7611_ & new_n7614_;
  assign new_n7616_ = new_n7608_ & new_n7615_;
  assign new_n7617_ = new_n1082_ & new_n7610_;
  assign new_n7618_ = new_n1059_ & new_n7610_;
  assign new_n7619_ = new_n1079_ & new_n7610_;
  assign new_n7620_ = ~new_n7618_ & ~new_n7619_;
  assign new_n7621_ = ~new_n7617_ & new_n7620_;
  assign new_n7622_ = new_n1076_ & new_n7610_;
  assign new_n7623_ = new_n1095_ & new_n7610_;
  assign new_n7624_ = ~new_n7622_ & ~new_n7623_;
  assign new_n7625_ = new_n7621_ & new_n7624_;
  assign new_n7626_ = new_n7616_ & new_n7625_;
  assign new_n7627_ = new_n7603_ & new_n7626_;
  assign new_n7628_ = new_n1105_ & new_n7610_;
  assign new_n7629_ = new_n1099_ & new_n7610_;
  assign new_n7630_ = new_n1089_ & new_n7610_;
  assign new_n7631_ = ~new_n7629_ & ~new_n7630_;
  assign new_n7632_ = ~new_n7628_ & new_n7631_;
  assign new_n7633_ = new_n1118_ & new_n7610_;
  assign new_n7634_ = new_n1107_ & new_n7610_;
  assign new_n7635_ = new_n1103_ & new_n7610_;
  assign new_n7636_ = ~new_n7634_ & ~new_n7635_;
  assign new_n7637_ = ~new_n7633_ & new_n7636_;
  assign new_n7638_ = new_n7632_ & new_n7637_;
  assign new_n7639_ = new_n1131_ & new_n7610_;
  assign new_n7640_ = new_n1120_ & new_n7610_;
  assign new_n7641_ = new_n1114_ & new_n7610_;
  assign new_n7642_ = ~new_n7640_ & ~new_n7641_;
  assign new_n7643_ = ~new_n7639_ & new_n7642_;
  assign new_n7644_ = new_n1145_ & new_n7610_;
  assign new_n7645_ = new_n1135_ & new_n7610_;
  assign new_n7646_ = new_n1127_ & new_n7610_;
  assign new_n7647_ = ~new_n7645_ & ~new_n7646_;
  assign new_n7648_ = ~new_n7644_ & new_n7647_;
  assign new_n7649_ = new_n7643_ & new_n7648_;
  assign new_n7650_ = new_n7638_ & new_n7649_;
  assign new_n7651_ = new_n1155_ & new_n7610_;
  assign new_n7652_ = new_n1149_ & new_n7610_;
  assign new_n7653_ = new_n1141_ & new_n7610_;
  assign new_n7654_ = ~new_n7652_ & ~new_n7653_;
  assign new_n7655_ = ~new_n7651_ & new_n7654_;
  assign new_n7656_ = new_n1165_ & new_n7610_;
  assign new_n7657_ = new_n1157_ & new_n7610_;
  assign new_n7658_ = new_n1153_ & new_n7610_;
  assign new_n7659_ = ~new_n7657_ & ~new_n7658_;
  assign new_n7660_ = ~new_n7656_ & new_n7659_;
  assign new_n7661_ = new_n7655_ & new_n7660_;
  assign new_n7662_ = new_n1172_ & new_n7610_;
  assign new_n7663_ = new_n1168_ & new_n7610_;
  assign new_n7664_ = new_n1162_ & new_n7610_;
  assign new_n7665_ = ~new_n7663_ & ~new_n7664_;
  assign new_n7666_ = ~new_n7662_ & new_n7665_;
  assign new_n7667_ = new_n1174_ & new_n7610_;
  assign new_n7668_ = new_n1184_ & new_n7610_;
  assign new_n7669_ = ~new_n7667_ & ~new_n7668_;
  assign new_n7670_ = new_n7666_ & new_n7669_;
  assign new_n7671_ = new_n7661_ & new_n7670_;
  assign new_n7672_ = new_n7650_ & new_n7671_;
  assign new_n7673_ = new_n7627_ & new_n7672_;
  assign new_n7674_ = new_n7580_ & new_n7673_;
  assign new_n7675_ = new_n1192_ & new_n7610_;
  assign new_n7676_ = new_n1186_ & new_n7610_;
  assign new_n7677_ = new_n1182_ & new_n7610_;
  assign new_n7678_ = ~new_n7676_ & ~new_n7677_;
  assign new_n7679_ = ~new_n7675_ & new_n7678_;
  assign new_n7680_ = new_n1202_ & new_n7610_;
  assign new_n7681_ = new_n1194_ & new_n7610_;
  assign new_n7682_ = new_n1190_ & new_n7610_;
  assign new_n7683_ = ~new_n7681_ & ~new_n7682_;
  assign new_n7684_ = ~new_n7680_ & new_n7683_;
  assign new_n7685_ = new_n7679_ & new_n7684_;
  assign new_n7686_ = new_n1213_ & new_n7610_;
  assign new_n7687_ = new_n1204_ & new_n7610_;
  assign new_n7688_ = new_n1200_ & new_n7610_;
  assign new_n7689_ = ~new_n7687_ & ~new_n7688_;
  assign new_n7690_ = ~new_n7686_ & new_n7689_;
  assign new_n7691_ = new_n1226_ & new_n7610_;
  assign new_n7692_ = new_n1216_ & new_n7610_;
  assign new_n7693_ = new_n1210_ & new_n7610_;
  assign new_n7694_ = ~new_n7692_ & ~new_n7693_;
  assign new_n7695_ = ~new_n7691_ & new_n7694_;
  assign new_n7696_ = new_n7690_ & new_n7695_;
  assign new_n7697_ = new_n7685_ & new_n7696_;
  assign new_n7698_ = new_n1235_ & new_n7610_;
  assign new_n7699_ = new_n1229_ & new_n7610_;
  assign new_n7700_ = new_n1223_ & new_n7610_;
  assign new_n7701_ = ~new_n7699_ & ~new_n7700_;
  assign new_n7702_ = ~new_n7698_ & new_n7701_;
  assign new_n7703_ = new_n1243_ & new_n7610_;
  assign new_n7704_ = new_n1237_ & new_n7610_;
  assign new_n7705_ = new_n1233_ & new_n7610_;
  assign new_n7706_ = ~new_n7704_ & ~new_n7705_;
  assign new_n7707_ = ~new_n7703_ & new_n7706_;
  assign new_n7708_ = new_n7702_ & new_n7707_;
  assign new_n7709_ = ~A201 & A200;
  assign new_n7710_ = ~A199 & new_n7709_;
  assign new_n7711_ = new_n6786_ & new_n7710_;
  assign new_n7712_ = new_n3662_ & new_n7711_;
  assign new_n7713_ = new_n3668_ & new_n7711_;
  assign new_n7714_ = new_n3670_ & new_n7711_;
  assign new_n7715_ = ~new_n7713_ & ~new_n7714_;
  assign new_n7716_ = ~new_n7712_ & new_n7715_;
  assign new_n7717_ = new_n3679_ & new_n7711_;
  assign new_n7718_ = new_n3681_ & new_n7711_;
  assign new_n7719_ = ~new_n7717_ & ~new_n7718_;
  assign new_n7720_ = new_n7716_ & new_n7719_;
  assign new_n7721_ = new_n7708_ & new_n7720_;
  assign new_n7722_ = new_n7697_ & new_n7721_;
  assign new_n7723_ = new_n3689_ & new_n7711_;
  assign new_n7724_ = new_n3677_ & new_n7711_;
  assign new_n7725_ = new_n3687_ & new_n7711_;
  assign new_n7726_ = ~new_n7724_ & ~new_n7725_;
  assign new_n7727_ = ~new_n7723_ & new_n7726_;
  assign new_n7728_ = new_n3698_ & new_n7711_;
  assign new_n7729_ = new_n3685_ & new_n7711_;
  assign new_n7730_ = new_n3696_ & new_n7711_;
  assign new_n7731_ = ~new_n7729_ & ~new_n7730_;
  assign new_n7732_ = ~new_n7728_ & new_n7731_;
  assign new_n7733_ = new_n7727_ & new_n7732_;
  assign new_n7734_ = new_n3705_ & new_n7711_;
  assign new_n7735_ = new_n3694_ & new_n7711_;
  assign new_n7736_ = new_n3703_ & new_n7711_;
  assign new_n7737_ = ~new_n7735_ & ~new_n7736_;
  assign new_n7738_ = ~new_n7734_ & new_n7737_;
  assign new_n7739_ = new_n3711_ & new_n7711_;
  assign new_n7740_ = new_n3713_ & new_n7711_;
  assign new_n7741_ = new_n3715_ & new_n7711_;
  assign new_n7742_ = ~new_n7740_ & ~new_n7741_;
  assign new_n7743_ = ~new_n7739_ & new_n7742_;
  assign new_n7744_ = new_n7738_ & new_n7743_;
  assign new_n7745_ = new_n7733_ & new_n7744_;
  assign new_n7746_ = new_n3719_ & new_n7711_;
  assign new_n7747_ = new_n3721_ & new_n7711_;
  assign new_n7748_ = new_n3723_ & new_n7711_;
  assign new_n7749_ = ~new_n7747_ & ~new_n7748_;
  assign new_n7750_ = ~new_n7746_ & new_n7749_;
  assign new_n7751_ = new_n3729_ & new_n7711_;
  assign new_n7752_ = new_n3731_ & new_n7711_;
  assign new_n7753_ = new_n3733_ & new_n7711_;
  assign new_n7754_ = ~new_n7752_ & ~new_n7753_;
  assign new_n7755_ = ~new_n7751_ & new_n7754_;
  assign new_n7756_ = new_n7750_ & new_n7755_;
  assign new_n7757_ = new_n3738_ & new_n7711_;
  assign new_n7758_ = new_n3740_ & new_n7711_;
  assign new_n7759_ = new_n3742_ & new_n7711_;
  assign new_n7760_ = ~new_n7758_ & ~new_n7759_;
  assign new_n7761_ = ~new_n7757_ & new_n7760_;
  assign new_n7762_ = new_n3751_ & new_n7711_;
  assign new_n7763_ = new_n3753_ & new_n7711_;
  assign new_n7764_ = ~new_n7762_ & ~new_n7763_;
  assign new_n7765_ = new_n7761_ & new_n7764_;
  assign new_n7766_ = new_n7756_ & new_n7765_;
  assign new_n7767_ = new_n7745_ & new_n7766_;
  assign new_n7768_ = new_n7722_ & new_n7767_;
  assign new_n7769_ = new_n3761_ & new_n7711_;
  assign new_n7770_ = new_n3749_ & new_n7711_;
  assign new_n7771_ = new_n3759_ & new_n7711_;
  assign new_n7772_ = ~new_n7770_ & ~new_n7771_;
  assign new_n7773_ = ~new_n7769_ & new_n7772_;
  assign new_n7774_ = new_n3771_ & new_n7711_;
  assign new_n7775_ = new_n3757_ & new_n7711_;
  assign new_n7776_ = new_n3769_ & new_n7711_;
  assign new_n7777_ = ~new_n7775_ & ~new_n7776_;
  assign new_n7778_ = ~new_n7774_ & new_n7777_;
  assign new_n7779_ = new_n7773_ & new_n7778_;
  assign new_n7780_ = new_n3778_ & new_n7711_;
  assign new_n7781_ = new_n3767_ & new_n7711_;
  assign new_n7782_ = new_n3775_ & new_n7711_;
  assign new_n7783_ = ~new_n7781_ & ~new_n7782_;
  assign new_n7784_ = ~new_n7780_ & new_n7783_;
  assign new_n7785_ = new_n3785_ & new_n7711_;
  assign new_n7786_ = new_n3787_ & new_n7711_;
  assign new_n7787_ = new_n3789_ & new_n7711_;
  assign new_n7788_ = ~new_n7786_ & ~new_n7787_;
  assign new_n7789_ = ~new_n7785_ & new_n7788_;
  assign new_n7790_ = new_n7784_ & new_n7789_;
  assign new_n7791_ = new_n7779_ & new_n7790_;
  assign new_n7792_ = new_n3793_ & new_n7711_;
  assign new_n7793_ = new_n3795_ & new_n7711_;
  assign new_n7794_ = new_n3797_ & new_n7711_;
  assign new_n7795_ = ~new_n7793_ & ~new_n7794_;
  assign new_n7796_ = ~new_n7792_ & new_n7795_;
  assign new_n7797_ = new_n3803_ & new_n7711_;
  assign new_n7798_ = new_n3805_ & new_n7711_;
  assign new_n7799_ = new_n3807_ & new_n7711_;
  assign new_n7800_ = ~new_n7798_ & ~new_n7799_;
  assign new_n7801_ = ~new_n7797_ & new_n7800_;
  assign new_n7802_ = new_n7796_ & new_n7801_;
  assign new_n7803_ = new_n3811_ & new_n7711_;
  assign new_n7804_ = new_n3813_ & new_n7711_;
  assign new_n7805_ = new_n3815_ & new_n7711_;
  assign new_n7806_ = ~new_n7804_ & ~new_n7805_;
  assign new_n7807_ = ~new_n7803_ & new_n7806_;
  assign new_n7808_ = new_n3823_ & new_n7711_;
  assign new_n7809_ = new_n3825_ & new_n7711_;
  assign new_n7810_ = ~new_n7808_ & ~new_n7809_;
  assign new_n7811_ = new_n7807_ & new_n7810_;
  assign new_n7812_ = new_n7802_ & new_n7811_;
  assign new_n7813_ = new_n7791_ & new_n7812_;
  assign new_n7814_ = new_n3834_ & new_n7711_;
  assign new_n7815_ = new_n3821_ & new_n7711_;
  assign new_n7816_ = new_n3832_ & new_n7711_;
  assign new_n7817_ = ~new_n7815_ & ~new_n7816_;
  assign new_n7818_ = ~new_n7814_ & new_n7817_;
  assign new_n7819_ = new_n3844_ & new_n7711_;
  assign new_n7820_ = new_n3830_ & new_n7711_;
  assign new_n7821_ = new_n3842_ & new_n7711_;
  assign new_n7822_ = ~new_n7820_ & ~new_n7821_;
  assign new_n7823_ = ~new_n7819_ & new_n7822_;
  assign new_n7824_ = new_n7818_ & new_n7823_;
  assign new_n7825_ = new_n3850_ & new_n7711_;
  assign new_n7826_ = new_n3840_ & new_n7711_;
  assign new_n7827_ = new_n3848_ & new_n7711_;
  assign new_n7828_ = ~new_n7826_ & ~new_n7827_;
  assign new_n7829_ = ~new_n7825_ & new_n7828_;
  assign new_n7830_ = new_n3857_ & new_n7711_;
  assign new_n7831_ = new_n3859_ & new_n7711_;
  assign new_n7832_ = new_n3861_ & new_n7711_;
  assign new_n7833_ = ~new_n7831_ & ~new_n7832_;
  assign new_n7834_ = ~new_n7830_ & new_n7833_;
  assign new_n7835_ = new_n7829_ & new_n7834_;
  assign new_n7836_ = new_n7824_ & new_n7835_;
  assign new_n7837_ = new_n6917_ & new_n7710_;
  assign new_n7838_ = new_n3670_ & new_n7837_;
  assign new_n7839_ = new_n3868_ & new_n7711_;
  assign new_n7840_ = new_n3668_ & new_n7837_;
  assign new_n7841_ = ~new_n7839_ & ~new_n7840_;
  assign new_n7842_ = ~new_n7838_ & new_n7841_;
  assign new_n7843_ = new_n3681_ & new_n7837_;
  assign new_n7844_ = new_n3662_ & new_n7837_;
  assign new_n7845_ = new_n3679_ & new_n7837_;
  assign new_n7846_ = ~new_n7844_ & ~new_n7845_;
  assign new_n7847_ = ~new_n7843_ & new_n7846_;
  assign new_n7848_ = new_n7842_ & new_n7847_;
  assign new_n7849_ = new_n3689_ & new_n7837_;
  assign new_n7850_ = new_n3677_ & new_n7837_;
  assign new_n7851_ = new_n3687_ & new_n7837_;
  assign new_n7852_ = ~new_n7850_ & ~new_n7851_;
  assign new_n7853_ = ~new_n7849_ & new_n7852_;
  assign new_n7854_ = new_n3685_ & new_n7837_;
  assign new_n7855_ = new_n3696_ & new_n7837_;
  assign new_n7856_ = ~new_n7854_ & ~new_n7855_;
  assign new_n7857_ = new_n7853_ & new_n7856_;
  assign new_n7858_ = new_n7848_ & new_n7857_;
  assign new_n7859_ = new_n7836_ & new_n7858_;
  assign new_n7860_ = new_n7813_ & new_n7859_;
  assign new_n7861_ = new_n7768_ & new_n7860_;
  assign new_n7862_ = new_n7674_ & new_n7861_;
  assign new_n7863_ = new_n3703_ & new_n7837_;
  assign new_n7864_ = new_n3698_ & new_n7837_;
  assign new_n7865_ = new_n3694_ & new_n7837_;
  assign new_n7866_ = ~new_n7864_ & ~new_n7865_;
  assign new_n7867_ = ~new_n7863_ & new_n7866_;
  assign new_n7868_ = new_n3715_ & new_n7837_;
  assign new_n7869_ = new_n3705_ & new_n7837_;
  assign new_n7870_ = new_n3713_ & new_n7837_;
  assign new_n7871_ = ~new_n7869_ & ~new_n7870_;
  assign new_n7872_ = ~new_n7868_ & new_n7871_;
  assign new_n7873_ = new_n7867_ & new_n7872_;
  assign new_n7874_ = new_n3723_ & new_n7837_;
  assign new_n7875_ = new_n3711_ & new_n7837_;
  assign new_n7876_ = new_n3721_ & new_n7837_;
  assign new_n7877_ = ~new_n7875_ & ~new_n7876_;
  assign new_n7878_ = ~new_n7874_ & new_n7877_;
  assign new_n7879_ = new_n3733_ & new_n7837_;
  assign new_n7880_ = new_n3719_ & new_n7837_;
  assign new_n7881_ = new_n3731_ & new_n7837_;
  assign new_n7882_ = ~new_n7880_ & ~new_n7881_;
  assign new_n7883_ = ~new_n7879_ & new_n7882_;
  assign new_n7884_ = new_n7878_ & new_n7883_;
  assign new_n7885_ = new_n7873_ & new_n7884_;
  assign new_n7886_ = new_n3742_ & new_n7837_;
  assign new_n7887_ = new_n3729_ & new_n7837_;
  assign new_n7888_ = new_n3740_ & new_n7837_;
  assign new_n7889_ = ~new_n7887_ & ~new_n7888_;
  assign new_n7890_ = ~new_n7886_ & new_n7889_;
  assign new_n7891_ = new_n3753_ & new_n7837_;
  assign new_n7892_ = new_n3738_ & new_n7837_;
  assign new_n7893_ = new_n3751_ & new_n7837_;
  assign new_n7894_ = ~new_n7892_ & ~new_n7893_;
  assign new_n7895_ = ~new_n7891_ & new_n7894_;
  assign new_n7896_ = new_n7890_ & new_n7895_;
  assign new_n7897_ = new_n3761_ & new_n7837_;
  assign new_n7898_ = new_n3749_ & new_n7837_;
  assign new_n7899_ = new_n3759_ & new_n7837_;
  assign new_n7900_ = ~new_n7898_ & ~new_n7899_;
  assign new_n7901_ = ~new_n7897_ & new_n7900_;
  assign new_n7902_ = new_n3757_ & new_n7837_;
  assign new_n7903_ = new_n3769_ & new_n7837_;
  assign new_n7904_ = ~new_n7902_ & ~new_n7903_;
  assign new_n7905_ = new_n7901_ & new_n7904_;
  assign new_n7906_ = new_n7896_ & new_n7905_;
  assign new_n7907_ = new_n7885_ & new_n7906_;
  assign new_n7908_ = new_n3775_ & new_n7837_;
  assign new_n7909_ = new_n3771_ & new_n7837_;
  assign new_n7910_ = new_n3767_ & new_n7837_;
  assign new_n7911_ = ~new_n7909_ & ~new_n7910_;
  assign new_n7912_ = ~new_n7908_ & new_n7911_;
  assign new_n7913_ = new_n3789_ & new_n7837_;
  assign new_n7914_ = new_n3778_ & new_n7837_;
  assign new_n7915_ = new_n3787_ & new_n7837_;
  assign new_n7916_ = ~new_n7914_ & ~new_n7915_;
  assign new_n7917_ = ~new_n7913_ & new_n7916_;
  assign new_n7918_ = new_n7912_ & new_n7917_;
  assign new_n7919_ = new_n3797_ & new_n7837_;
  assign new_n7920_ = new_n3785_ & new_n7837_;
  assign new_n7921_ = new_n3795_ & new_n7837_;
  assign new_n7922_ = ~new_n7920_ & ~new_n7921_;
  assign new_n7923_ = ~new_n7919_ & new_n7922_;
  assign new_n7924_ = new_n3807_ & new_n7837_;
  assign new_n7925_ = new_n3793_ & new_n7837_;
  assign new_n7926_ = new_n3805_ & new_n7837_;
  assign new_n7927_ = ~new_n7925_ & ~new_n7926_;
  assign new_n7928_ = ~new_n7924_ & new_n7927_;
  assign new_n7929_ = new_n7923_ & new_n7928_;
  assign new_n7930_ = new_n7918_ & new_n7929_;
  assign new_n7931_ = new_n3815_ & new_n7837_;
  assign new_n7932_ = new_n3803_ & new_n7837_;
  assign new_n7933_ = new_n3813_ & new_n7837_;
  assign new_n7934_ = ~new_n7932_ & ~new_n7933_;
  assign new_n7935_ = ~new_n7931_ & new_n7934_;
  assign new_n7936_ = new_n3825_ & new_n7837_;
  assign new_n7937_ = new_n3811_ & new_n7837_;
  assign new_n7938_ = new_n3823_ & new_n7837_;
  assign new_n7939_ = ~new_n7937_ & ~new_n7938_;
  assign new_n7940_ = ~new_n7936_ & new_n7939_;
  assign new_n7941_ = new_n7935_ & new_n7940_;
  assign new_n7942_ = new_n3834_ & new_n7837_;
  assign new_n7943_ = new_n3821_ & new_n7837_;
  assign new_n7944_ = new_n3832_ & new_n7837_;
  assign new_n7945_ = ~new_n7943_ & ~new_n7944_;
  assign new_n7946_ = ~new_n7942_ & new_n7945_;
  assign new_n7947_ = new_n3830_ & new_n7837_;
  assign new_n7948_ = new_n3842_ & new_n7837_;
  assign new_n7949_ = ~new_n7947_ & ~new_n7948_;
  assign new_n7950_ = new_n7946_ & new_n7949_;
  assign new_n7951_ = new_n7941_ & new_n7950_;
  assign new_n7952_ = new_n7930_ & new_n7951_;
  assign new_n7953_ = new_n7907_ & new_n7952_;
  assign new_n7954_ = new_n3848_ & new_n7837_;
  assign new_n7955_ = new_n3844_ & new_n7837_;
  assign new_n7956_ = new_n3840_ & new_n7837_;
  assign new_n7957_ = ~new_n7955_ & ~new_n7956_;
  assign new_n7958_ = ~new_n7954_ & new_n7957_;
  assign new_n7959_ = new_n3861_ & new_n7837_;
  assign new_n7960_ = new_n3850_ & new_n7837_;
  assign new_n7961_ = new_n3859_ & new_n7837_;
  assign new_n7962_ = ~new_n7960_ & ~new_n7961_;
  assign new_n7963_ = ~new_n7959_ & new_n7962_;
  assign new_n7964_ = new_n7958_ & new_n7963_;
  assign new_n7965_ = A201 & A200;
  assign new_n7966_ = ~A199 & new_n7965_;
  assign new_n7967_ = new_n7046_ & new_n7966_;
  assign new_n7968_ = new_n951_ & new_n7967_;
  assign new_n7969_ = new_n3857_ & new_n7837_;
  assign new_n7970_ = new_n3868_ & new_n7837_;
  assign new_n7971_ = ~new_n7969_ & ~new_n7970_;
  assign new_n7972_ = ~new_n7968_ & new_n7971_;
  assign new_n7973_ = new_n964_ & new_n7967_;
  assign new_n7974_ = new_n954_ & new_n7967_;
  assign new_n7975_ = new_n948_ & new_n7967_;
  assign new_n7976_ = ~new_n7974_ & ~new_n7975_;
  assign new_n7977_ = ~new_n7973_ & new_n7976_;
  assign new_n7978_ = new_n7972_ & new_n7977_;
  assign new_n7979_ = new_n7964_ & new_n7978_;
  assign new_n7980_ = new_n975_ & new_n7967_;
  assign new_n7981_ = new_n967_ & new_n7967_;
  assign new_n7982_ = new_n961_ & new_n7967_;
  assign new_n7983_ = ~new_n7981_ & ~new_n7982_;
  assign new_n7984_ = ~new_n7980_ & new_n7983_;
  assign new_n7985_ = new_n987_ & new_n7967_;
  assign new_n7986_ = new_n978_ & new_n7967_;
  assign new_n7987_ = new_n972_ & new_n7967_;
  assign new_n7988_ = ~new_n7986_ & ~new_n7987_;
  assign new_n7989_ = ~new_n7985_ & new_n7988_;
  assign new_n7990_ = new_n7984_ & new_n7989_;
  assign new_n7991_ = new_n994_ & new_n7967_;
  assign new_n7992_ = new_n990_ & new_n7967_;
  assign new_n7993_ = new_n984_ & new_n7967_;
  assign new_n7994_ = ~new_n7992_ & ~new_n7993_;
  assign new_n7995_ = ~new_n7991_ & new_n7994_;
  assign new_n7996_ = new_n996_ & new_n7967_;
  assign new_n7997_ = new_n1008_ & new_n7967_;
  assign new_n7998_ = ~new_n7996_ & ~new_n7997_;
  assign new_n7999_ = new_n7995_ & new_n7998_;
  assign new_n8000_ = new_n7990_ & new_n7999_;
  assign new_n8001_ = new_n7979_ & new_n8000_;
  assign new_n8002_ = new_n1016_ & new_n7967_;
  assign new_n8003_ = new_n1010_ & new_n7967_;
  assign new_n8004_ = new_n1006_ & new_n7967_;
  assign new_n8005_ = ~new_n8003_ & ~new_n8004_;
  assign new_n8006_ = ~new_n8002_ & new_n8005_;
  assign new_n8007_ = new_n1025_ & new_n7967_;
  assign new_n8008_ = new_n1018_ & new_n7967_;
  assign new_n8009_ = new_n1014_ & new_n7967_;
  assign new_n8010_ = ~new_n8008_ & ~new_n8009_;
  assign new_n8011_ = ~new_n8007_ & new_n8010_;
  assign new_n8012_ = new_n8006_ & new_n8011_;
  assign new_n8013_ = new_n1033_ & new_n7967_;
  assign new_n8014_ = new_n1027_ & new_n7967_;
  assign new_n8015_ = new_n1023_ & new_n7967_;
  assign new_n8016_ = ~new_n8014_ & ~new_n8015_;
  assign new_n8017_ = ~new_n8013_ & new_n8016_;
  assign new_n8018_ = new_n1043_ & new_n7967_;
  assign new_n8019_ = new_n1035_ & new_n7967_;
  assign new_n8020_ = new_n1031_ & new_n7967_;
  assign new_n8021_ = ~new_n8019_ & ~new_n8020_;
  assign new_n8022_ = ~new_n8018_ & new_n8021_;
  assign new_n8023_ = new_n8017_ & new_n8022_;
  assign new_n8024_ = new_n8012_ & new_n8023_;
  assign new_n8025_ = new_n1051_ & new_n7967_;
  assign new_n8026_ = new_n1045_ & new_n7967_;
  assign new_n8027_ = new_n1041_ & new_n7967_;
  assign new_n8028_ = ~new_n8026_ & ~new_n8027_;
  assign new_n8029_ = ~new_n8025_ & new_n8028_;
  assign new_n8030_ = new_n7114_ & new_n7966_;
  assign new_n8031_ = new_n1065_ & new_n8030_;
  assign new_n8032_ = new_n1053_ & new_n7967_;
  assign new_n8033_ = new_n1049_ & new_n7967_;
  assign new_n8034_ = ~new_n8032_ & ~new_n8033_;
  assign new_n8035_ = ~new_n8031_ & new_n8034_;
  assign new_n8036_ = new_n8029_ & new_n8035_;
  assign new_n8037_ = new_n1079_ & new_n8030_;
  assign new_n8038_ = new_n1071_ & new_n8030_;
  assign new_n8039_ = new_n1059_ & new_n8030_;
  assign new_n8040_ = ~new_n8038_ & ~new_n8039_;
  assign new_n8041_ = ~new_n8037_ & new_n8040_;
  assign new_n8042_ = new_n1082_ & new_n8030_;
  assign new_n8043_ = new_n1076_ & new_n8030_;
  assign new_n8044_ = ~new_n8042_ & ~new_n8043_;
  assign new_n8045_ = new_n8041_ & new_n8044_;
  assign new_n8046_ = new_n8036_ & new_n8045_;
  assign new_n8047_ = new_n8024_ & new_n8046_;
  assign new_n8048_ = new_n8001_ & new_n8047_;
  assign new_n8049_ = new_n7953_ & new_n8048_;
  assign new_n8050_ = new_n1089_ & new_n8030_;
  assign new_n8051_ = new_n1095_ & new_n8030_;
  assign new_n8052_ = new_n1099_ & new_n8030_;
  assign new_n8053_ = ~new_n8051_ & ~new_n8052_;
  assign new_n8054_ = ~new_n8050_ & new_n8053_;
  assign new_n8055_ = new_n1103_ & new_n8030_;
  assign new_n8056_ = new_n1105_ & new_n8030_;
  assign new_n8057_ = new_n1107_ & new_n8030_;
  assign new_n8058_ = ~new_n8056_ & ~new_n8057_;
  assign new_n8059_ = ~new_n8055_ & new_n8058_;
  assign new_n8060_ = new_n8054_ & new_n8059_;
  assign new_n8061_ = new_n1114_ & new_n8030_;
  assign new_n8062_ = new_n1118_ & new_n8030_;
  assign new_n8063_ = new_n1120_ & new_n8030_;
  assign new_n8064_ = ~new_n8062_ & ~new_n8063_;
  assign new_n8065_ = ~new_n8061_ & new_n8064_;
  assign new_n8066_ = new_n1127_ & new_n8030_;
  assign new_n8067_ = new_n1131_ & new_n8030_;
  assign new_n8068_ = new_n1135_ & new_n8030_;
  assign new_n8069_ = ~new_n8067_ & ~new_n8068_;
  assign new_n8070_ = ~new_n8066_ & new_n8069_;
  assign new_n8071_ = new_n8065_ & new_n8070_;
  assign new_n8072_ = new_n8060_ & new_n8071_;
  assign new_n8073_ = new_n1141_ & new_n8030_;
  assign new_n8074_ = new_n1145_ & new_n8030_;
  assign new_n8075_ = new_n1149_ & new_n8030_;
  assign new_n8076_ = ~new_n8074_ & ~new_n8075_;
  assign new_n8077_ = ~new_n8073_ & new_n8076_;
  assign new_n8078_ = new_n1153_ & new_n8030_;
  assign new_n8079_ = new_n1155_ & new_n8030_;
  assign new_n8080_ = new_n1157_ & new_n8030_;
  assign new_n8081_ = ~new_n8079_ & ~new_n8080_;
  assign new_n8082_ = ~new_n8078_ & new_n8081_;
  assign new_n8083_ = new_n8077_ & new_n8082_;
  assign new_n8084_ = new_n1162_ & new_n8030_;
  assign new_n8085_ = new_n1165_ & new_n8030_;
  assign new_n8086_ = new_n1168_ & new_n8030_;
  assign new_n8087_ = ~new_n8085_ & ~new_n8086_;
  assign new_n8088_ = ~new_n8084_ & new_n8087_;
  assign new_n8089_ = new_n1172_ & new_n8030_;
  assign new_n8090_ = new_n1174_ & new_n8030_;
  assign new_n8091_ = ~new_n8089_ & ~new_n8090_;
  assign new_n8092_ = new_n8088_ & new_n8091_;
  assign new_n8093_ = new_n8083_ & new_n8092_;
  assign new_n8094_ = new_n8072_ & new_n8093_;
  assign new_n8095_ = new_n1182_ & new_n8030_;
  assign new_n8096_ = new_n1184_ & new_n8030_;
  assign new_n8097_ = new_n1186_ & new_n8030_;
  assign new_n8098_ = ~new_n8096_ & ~new_n8097_;
  assign new_n8099_ = ~new_n8095_ & new_n8098_;
  assign new_n8100_ = new_n1190_ & new_n8030_;
  assign new_n8101_ = new_n1192_ & new_n8030_;
  assign new_n8102_ = new_n1194_ & new_n8030_;
  assign new_n8103_ = ~new_n8101_ & ~new_n8102_;
  assign new_n8104_ = ~new_n8100_ & new_n8103_;
  assign new_n8105_ = new_n8099_ & new_n8104_;
  assign new_n8106_ = new_n1200_ & new_n8030_;
  assign new_n8107_ = new_n1202_ & new_n8030_;
  assign new_n8108_ = new_n1204_ & new_n8030_;
  assign new_n8109_ = ~new_n8107_ & ~new_n8108_;
  assign new_n8110_ = ~new_n8106_ & new_n8109_;
  assign new_n8111_ = new_n1210_ & new_n8030_;
  assign new_n8112_ = new_n1213_ & new_n8030_;
  assign new_n8113_ = new_n1216_ & new_n8030_;
  assign new_n8114_ = ~new_n8112_ & ~new_n8113_;
  assign new_n8115_ = ~new_n8111_ & new_n8114_;
  assign new_n8116_ = new_n8110_ & new_n8115_;
  assign new_n8117_ = new_n8105_ & new_n8116_;
  assign new_n8118_ = new_n1223_ & new_n8030_;
  assign new_n8119_ = new_n1226_ & new_n8030_;
  assign new_n8120_ = new_n1229_ & new_n8030_;
  assign new_n8121_ = ~new_n8119_ & ~new_n8120_;
  assign new_n8122_ = ~new_n8118_ & new_n8121_;
  assign new_n8123_ = new_n1233_ & new_n8030_;
  assign new_n8124_ = new_n1235_ & new_n8030_;
  assign new_n8125_ = new_n1237_ & new_n8030_;
  assign new_n8126_ = ~new_n8124_ & ~new_n8125_;
  assign new_n8127_ = ~new_n8123_ & new_n8126_;
  assign new_n8128_ = new_n8122_ & new_n8127_;
  assign new_n8129_ = new_n7215_ & new_n7966_;
  assign new_n8130_ = new_n954_ & new_n8129_;
  assign new_n8131_ = new_n1243_ & new_n8030_;
  assign new_n8132_ = new_n951_ & new_n8129_;
  assign new_n8133_ = ~new_n8131_ & ~new_n8132_;
  assign new_n8134_ = ~new_n8130_ & new_n8133_;
  assign new_n8135_ = new_n948_ & new_n8129_;
  assign new_n8136_ = new_n964_ & new_n8129_;
  assign new_n8137_ = ~new_n8135_ & ~new_n8136_;
  assign new_n8138_ = new_n8134_ & new_n8137_;
  assign new_n8139_ = new_n8128_ & new_n8138_;
  assign new_n8140_ = new_n8117_ & new_n8139_;
  assign new_n8141_ = new_n8094_ & new_n8140_;
  assign new_n8142_ = new_n975_ & new_n8129_;
  assign new_n8143_ = new_n967_ & new_n8129_;
  assign new_n8144_ = new_n961_ & new_n8129_;
  assign new_n8145_ = ~new_n8143_ & ~new_n8144_;
  assign new_n8146_ = ~new_n8142_ & new_n8145_;
  assign new_n8147_ = new_n987_ & new_n8129_;
  assign new_n8148_ = new_n978_ & new_n8129_;
  assign new_n8149_ = new_n972_ & new_n8129_;
  assign new_n8150_ = ~new_n8148_ & ~new_n8149_;
  assign new_n8151_ = ~new_n8147_ & new_n8150_;
  assign new_n8152_ = new_n8146_ & new_n8151_;
  assign new_n8153_ = new_n994_ & new_n8129_;
  assign new_n8154_ = new_n990_ & new_n8129_;
  assign new_n8155_ = new_n984_ & new_n8129_;
  assign new_n8156_ = ~new_n8154_ & ~new_n8155_;
  assign new_n8157_ = ~new_n8153_ & new_n8156_;
  assign new_n8158_ = new_n1010_ & new_n8129_;
  assign new_n8159_ = new_n996_ & new_n8129_;
  assign new_n8160_ = new_n1008_ & new_n8129_;
  assign new_n8161_ = ~new_n8159_ & ~new_n8160_;
  assign new_n8162_ = ~new_n8158_ & new_n8161_;
  assign new_n8163_ = new_n8157_ & new_n8162_;
  assign new_n8164_ = new_n8152_ & new_n8163_;
  assign new_n8165_ = new_n1018_ & new_n8129_;
  assign new_n8166_ = new_n1006_ & new_n8129_;
  assign new_n8167_ = new_n1016_ & new_n8129_;
  assign new_n8168_ = ~new_n8166_ & ~new_n8167_;
  assign new_n8169_ = ~new_n8165_ & new_n8168_;
  assign new_n8170_ = new_n1027_ & new_n8129_;
  assign new_n8171_ = new_n1014_ & new_n8129_;
  assign new_n8172_ = new_n1025_ & new_n8129_;
  assign new_n8173_ = ~new_n8171_ & ~new_n8172_;
  assign new_n8174_ = ~new_n8170_ & new_n8173_;
  assign new_n8175_ = new_n8169_ & new_n8174_;
  assign new_n8176_ = new_n1035_ & new_n8129_;
  assign new_n8177_ = new_n1023_ & new_n8129_;
  assign new_n8178_ = new_n1033_ & new_n8129_;
  assign new_n8179_ = ~new_n8177_ & ~new_n8178_;
  assign new_n8180_ = ~new_n8176_ & new_n8179_;
  assign new_n8181_ = new_n1031_ & new_n8129_;
  assign new_n8182_ = new_n1043_ & new_n8129_;
  assign new_n8183_ = ~new_n8181_ & ~new_n8182_;
  assign new_n8184_ = new_n8180_ & new_n8183_;
  assign new_n8185_ = new_n8175_ & new_n8184_;
  assign new_n8186_ = new_n8164_ & new_n8185_;
  assign new_n8187_ = new_n1051_ & new_n8129_;
  assign new_n8188_ = new_n1045_ & new_n8129_;
  assign new_n8189_ = new_n1041_ & new_n8129_;
  assign new_n8190_ = ~new_n8188_ & ~new_n8189_;
  assign new_n8191_ = ~new_n8187_ & new_n8190_;
  assign new_n8192_ = new_n7280_ & new_n7966_;
  assign new_n8193_ = new_n1065_ & new_n8192_;
  assign new_n8194_ = new_n1053_ & new_n8129_;
  assign new_n8195_ = new_n1049_ & new_n8129_;
  assign new_n8196_ = ~new_n8194_ & ~new_n8195_;
  assign new_n8197_ = ~new_n8193_ & new_n8196_;
  assign new_n8198_ = new_n8191_ & new_n8197_;
  assign new_n8199_ = new_n1079_ & new_n8192_;
  assign new_n8200_ = new_n1071_ & new_n8192_;
  assign new_n8201_ = new_n1059_ & new_n8192_;
  assign new_n8202_ = ~new_n8200_ & ~new_n8201_;
  assign new_n8203_ = ~new_n8199_ & new_n8202_;
  assign new_n8204_ = new_n1095_ & new_n8192_;
  assign new_n8205_ = new_n1082_ & new_n8192_;
  assign new_n8206_ = new_n1076_ & new_n8192_;
  assign new_n8207_ = ~new_n8205_ & ~new_n8206_;
  assign new_n8208_ = ~new_n8204_ & new_n8207_;
  assign new_n8209_ = new_n8203_ & new_n8208_;
  assign new_n8210_ = new_n8198_ & new_n8209_;
  assign new_n8211_ = new_n1105_ & new_n8192_;
  assign new_n8212_ = new_n1099_ & new_n8192_;
  assign new_n8213_ = new_n1089_ & new_n8192_;
  assign new_n8214_ = ~new_n8212_ & ~new_n8213_;
  assign new_n8215_ = ~new_n8211_ & new_n8214_;
  assign new_n8216_ = new_n1118_ & new_n8192_;
  assign new_n8217_ = new_n1107_ & new_n8192_;
  assign new_n8218_ = new_n1103_ & new_n8192_;
  assign new_n8219_ = ~new_n8217_ & ~new_n8218_;
  assign new_n8220_ = ~new_n8216_ & new_n8219_;
  assign new_n8221_ = new_n8215_ & new_n8220_;
  assign new_n8222_ = new_n1131_ & new_n8192_;
  assign new_n8223_ = new_n1120_ & new_n8192_;
  assign new_n8224_ = new_n1114_ & new_n8192_;
  assign new_n8225_ = ~new_n8223_ & ~new_n8224_;
  assign new_n8226_ = ~new_n8222_ & new_n8225_;
  assign new_n8227_ = new_n1135_ & new_n8192_;
  assign new_n8228_ = new_n1127_ & new_n8192_;
  assign new_n8229_ = ~new_n8227_ & ~new_n8228_;
  assign new_n8230_ = new_n8226_ & new_n8229_;
  assign new_n8231_ = new_n8221_ & new_n8230_;
  assign new_n8232_ = new_n8210_ & new_n8231_;
  assign new_n8233_ = new_n8186_ & new_n8232_;
  assign new_n8234_ = new_n8141_ & new_n8233_;
  assign new_n8235_ = new_n8049_ & new_n8234_;
  assign new_n8236_ = new_n7862_ & new_n8235_;
  assign new_n8237_ = new_n7484_ & new_n8236_;
  assign new_n8238_ = new_n1141_ & new_n8192_;
  assign new_n8239_ = new_n1145_ & new_n8192_;
  assign new_n8240_ = new_n1149_ & new_n8192_;
  assign new_n8241_ = ~new_n8239_ & ~new_n8240_;
  assign new_n8242_ = ~new_n8238_ & new_n8241_;
  assign new_n8243_ = new_n1153_ & new_n8192_;
  assign new_n8244_ = new_n1155_ & new_n8192_;
  assign new_n8245_ = new_n1157_ & new_n8192_;
  assign new_n8246_ = ~new_n8244_ & ~new_n8245_;
  assign new_n8247_ = ~new_n8243_ & new_n8246_;
  assign new_n8248_ = new_n8242_ & new_n8247_;
  assign new_n8249_ = new_n1162_ & new_n8192_;
  assign new_n8250_ = new_n1165_ & new_n8192_;
  assign new_n8251_ = new_n1168_ & new_n8192_;
  assign new_n8252_ = ~new_n8250_ & ~new_n8251_;
  assign new_n8253_ = ~new_n8249_ & new_n8252_;
  assign new_n8254_ = new_n1184_ & new_n8192_;
  assign new_n8255_ = new_n1172_ & new_n8192_;
  assign new_n8256_ = new_n1174_ & new_n8192_;
  assign new_n8257_ = ~new_n8255_ & ~new_n8256_;
  assign new_n8258_ = ~new_n8254_ & new_n8257_;
  assign new_n8259_ = new_n8253_ & new_n8258_;
  assign new_n8260_ = new_n8248_ & new_n8259_;
  assign new_n8261_ = new_n1192_ & new_n8192_;
  assign new_n8262_ = new_n1186_ & new_n8192_;
  assign new_n8263_ = new_n1182_ & new_n8192_;
  assign new_n8264_ = ~new_n8262_ & ~new_n8263_;
  assign new_n8265_ = ~new_n8261_ & new_n8264_;
  assign new_n8266_ = new_n1202_ & new_n8192_;
  assign new_n8267_ = new_n1194_ & new_n8192_;
  assign new_n8268_ = new_n1190_ & new_n8192_;
  assign new_n8269_ = ~new_n8267_ & ~new_n8268_;
  assign new_n8270_ = ~new_n8266_ & new_n8269_;
  assign new_n8271_ = new_n8265_ & new_n8270_;
  assign new_n8272_ = new_n1213_ & new_n8192_;
  assign new_n8273_ = new_n1204_ & new_n8192_;
  assign new_n8274_ = new_n1200_ & new_n8192_;
  assign new_n8275_ = ~new_n8273_ & ~new_n8274_;
  assign new_n8276_ = ~new_n8272_ & new_n8275_;
  assign new_n8277_ = new_n1226_ & new_n8192_;
  assign new_n8278_ = new_n1216_ & new_n8192_;
  assign new_n8279_ = new_n1210_ & new_n8192_;
  assign new_n8280_ = ~new_n8278_ & ~new_n8279_;
  assign new_n8281_ = ~new_n8277_ & new_n8280_;
  assign new_n8282_ = new_n8276_ & new_n8281_;
  assign new_n8283_ = new_n8271_ & new_n8282_;
  assign new_n8284_ = new_n8260_ & new_n8283_;
  assign new_n8285_ = new_n1235_ & new_n8192_;
  assign new_n8286_ = new_n1229_ & new_n8192_;
  assign new_n8287_ = new_n1223_ & new_n8192_;
  assign new_n8288_ = ~new_n8286_ & ~new_n8287_;
  assign new_n8289_ = ~new_n8285_ & new_n8288_;
  assign new_n8290_ = new_n1243_ & new_n8192_;
  assign new_n8291_ = new_n1237_ & new_n8192_;
  assign new_n8292_ = new_n1233_ & new_n8192_;
  assign new_n8293_ = ~new_n8291_ & ~new_n8292_;
  assign new_n8294_ = ~new_n8290_ & new_n8293_;
  assign new_n8295_ = new_n8289_ & new_n8294_;
  assign new_n8296_ = new_n7375_ & new_n7966_;
  assign new_n8297_ = new_n948_ & new_n8296_;
  assign new_n8298_ = new_n951_ & new_n8296_;
  assign new_n8299_ = new_n954_ & new_n8296_;
  assign new_n8300_ = ~new_n8298_ & ~new_n8299_;
  assign new_n8301_ = ~new_n8297_ & new_n8300_;
  assign new_n8302_ = new_n961_ & new_n8296_;
  assign new_n8303_ = new_n964_ & new_n8296_;
  assign new_n8304_ = new_n967_ & new_n8296_;
  assign new_n8305_ = ~new_n8303_ & ~new_n8304_;
  assign new_n8306_ = ~new_n8302_ & new_n8305_;
  assign new_n8307_ = new_n8301_ & new_n8306_;
  assign new_n8308_ = new_n8295_ & new_n8307_;
  assign new_n8309_ = new_n972_ & new_n8296_;
  assign new_n8310_ = new_n975_ & new_n8296_;
  assign new_n8311_ = new_n978_ & new_n8296_;
  assign new_n8312_ = ~new_n8310_ & ~new_n8311_;
  assign new_n8313_ = ~new_n8309_ & new_n8312_;
  assign new_n8314_ = new_n984_ & new_n8296_;
  assign new_n8315_ = new_n987_ & new_n8296_;
  assign new_n8316_ = new_n990_ & new_n8296_;
  assign new_n8317_ = ~new_n8315_ & ~new_n8316_;
  assign new_n8318_ = ~new_n8314_ & new_n8317_;
  assign new_n8319_ = new_n8313_ & new_n8318_;
  assign new_n8320_ = new_n1008_ & new_n8296_;
  assign new_n8321_ = new_n994_ & new_n8296_;
  assign new_n8322_ = new_n996_ & new_n8296_;
  assign new_n8323_ = ~new_n8321_ & ~new_n8322_;
  assign new_n8324_ = ~new_n8320_ & new_n8323_;
  assign new_n8325_ = new_n1010_ & new_n8296_;
  assign new_n8326_ = new_n1006_ & new_n8296_;
  assign new_n8327_ = ~new_n8325_ & ~new_n8326_;
  assign new_n8328_ = new_n8324_ & new_n8327_;
  assign new_n8329_ = new_n8319_ & new_n8328_;
  assign new_n8330_ = new_n8308_ & new_n8329_;
  assign new_n8331_ = new_n8284_ & new_n8330_;
  assign new_n8332_ = new_n1014_ & new_n8296_;
  assign new_n8333_ = new_n1016_ & new_n8296_;
  assign new_n8334_ = new_n1018_ & new_n8296_;
  assign new_n8335_ = ~new_n8333_ & ~new_n8334_;
  assign new_n8336_ = ~new_n8332_ & new_n8335_;
  assign new_n8337_ = new_n1023_ & new_n8296_;
  assign new_n8338_ = new_n1025_ & new_n8296_;
  assign new_n8339_ = new_n1027_ & new_n8296_;
  assign new_n8340_ = ~new_n8338_ & ~new_n8339_;
  assign new_n8341_ = ~new_n8337_ & new_n8340_;
  assign new_n8342_ = new_n8336_ & new_n8341_;
  assign new_n8343_ = new_n1031_ & new_n8296_;
  assign new_n8344_ = new_n1033_ & new_n8296_;
  assign new_n8345_ = new_n1035_ & new_n8296_;
  assign new_n8346_ = ~new_n8344_ & ~new_n8345_;
  assign new_n8347_ = ~new_n8343_ & new_n8346_;
  assign new_n8348_ = new_n1041_ & new_n8296_;
  assign new_n8349_ = new_n1043_ & new_n8296_;
  assign new_n8350_ = new_n1045_ & new_n8296_;
  assign new_n8351_ = ~new_n8349_ & ~new_n8350_;
  assign new_n8352_ = ~new_n8348_ & new_n8351_;
  assign new_n8353_ = new_n8347_ & new_n8352_;
  assign new_n8354_ = new_n8342_ & new_n8353_;
  assign new_n8355_ = new_n1049_ & new_n8296_;
  assign new_n8356_ = new_n1051_ & new_n8296_;
  assign new_n8357_ = new_n1053_ & new_n8296_;
  assign new_n8358_ = ~new_n8356_ & ~new_n8357_;
  assign new_n8359_ = ~new_n8355_ & new_n8358_;
  assign new_n8360_ = new_n7445_ & new_n7966_;
  assign new_n8361_ = new_n1059_ & new_n8360_;
  assign new_n8362_ = new_n1065_ & new_n8360_;
  assign new_n8363_ = new_n1071_ & new_n8360_;
  assign new_n8364_ = ~new_n8362_ & ~new_n8363_;
  assign new_n8365_ = ~new_n8361_ & new_n8364_;
  assign new_n8366_ = new_n8359_ & new_n8365_;
  assign new_n8367_ = new_n1076_ & new_n8360_;
  assign new_n8368_ = new_n1079_ & new_n8360_;
  assign new_n8369_ = new_n1082_ & new_n8360_;
  assign new_n8370_ = ~new_n8368_ & ~new_n8369_;
  assign new_n8371_ = ~new_n8367_ & new_n8370_;
  assign new_n8372_ = new_n1095_ & new_n8360_;
  assign new_n8373_ = new_n1099_ & new_n8360_;
  assign new_n8374_ = ~new_n8372_ & ~new_n8373_;
  assign new_n8375_ = new_n8371_ & new_n8374_;
  assign new_n8376_ = new_n8366_ & new_n8375_;
  assign new_n8377_ = new_n8354_ & new_n8376_;
  assign new_n8378_ = new_n1107_ & new_n8360_;
  assign new_n8379_ = new_n1089_ & new_n8360_;
  assign new_n8380_ = new_n1105_ & new_n8360_;
  assign new_n8381_ = ~new_n8379_ & ~new_n8380_;
  assign new_n8382_ = ~new_n8378_ & new_n8381_;
  assign new_n8383_ = new_n1120_ & new_n8360_;
  assign new_n8384_ = new_n1103_ & new_n8360_;
  assign new_n8385_ = new_n1118_ & new_n8360_;
  assign new_n8386_ = ~new_n8384_ & ~new_n8385_;
  assign new_n8387_ = ~new_n8383_ & new_n8386_;
  assign new_n8388_ = new_n8382_ & new_n8387_;
  assign new_n8389_ = new_n1135_ & new_n8360_;
  assign new_n8390_ = new_n1114_ & new_n8360_;
  assign new_n8391_ = new_n1131_ & new_n8360_;
  assign new_n8392_ = ~new_n8390_ & ~new_n8391_;
  assign new_n8393_ = ~new_n8389_ & new_n8392_;
  assign new_n8394_ = new_n1149_ & new_n8360_;
  assign new_n8395_ = new_n1127_ & new_n8360_;
  assign new_n8396_ = new_n1145_ & new_n8360_;
  assign new_n8397_ = ~new_n8395_ & ~new_n8396_;
  assign new_n8398_ = ~new_n8394_ & new_n8397_;
  assign new_n8399_ = new_n8393_ & new_n8398_;
  assign new_n8400_ = new_n8388_ & new_n8399_;
  assign new_n8401_ = new_n1157_ & new_n8360_;
  assign new_n8402_ = new_n1141_ & new_n8360_;
  assign new_n8403_ = new_n1155_ & new_n8360_;
  assign new_n8404_ = ~new_n8402_ & ~new_n8403_;
  assign new_n8405_ = ~new_n8401_ & new_n8404_;
  assign new_n8406_ = new_n1168_ & new_n8360_;
  assign new_n8407_ = new_n1153_ & new_n8360_;
  assign new_n8408_ = new_n1165_ & new_n8360_;
  assign new_n8409_ = ~new_n8407_ & ~new_n8408_;
  assign new_n8410_ = ~new_n8406_ & new_n8409_;
  assign new_n8411_ = new_n8405_ & new_n8410_;
  assign new_n8412_ = new_n1174_ & new_n8360_;
  assign new_n8413_ = new_n1162_ & new_n8360_;
  assign new_n8414_ = new_n1172_ & new_n8360_;
  assign new_n8415_ = ~new_n8413_ & ~new_n8414_;
  assign new_n8416_ = ~new_n8412_ & new_n8415_;
  assign new_n8417_ = new_n1184_ & new_n8360_;
  assign new_n8418_ = new_n1186_ & new_n8360_;
  assign new_n8419_ = ~new_n8417_ & ~new_n8418_;
  assign new_n8420_ = new_n8416_ & new_n8419_;
  assign new_n8421_ = new_n8411_ & new_n8420_;
  assign new_n8422_ = new_n8400_ & new_n8421_;
  assign new_n8423_ = new_n8377_ & new_n8422_;
  assign new_n8424_ = new_n8331_ & new_n8423_;
  assign new_n8425_ = new_n1194_ & new_n8360_;
  assign new_n8426_ = new_n1182_ & new_n8360_;
  assign new_n8427_ = new_n1192_ & new_n8360_;
  assign new_n8428_ = ~new_n8426_ & ~new_n8427_;
  assign new_n8429_ = ~new_n8425_ & new_n8428_;
  assign new_n8430_ = new_n1204_ & new_n8360_;
  assign new_n8431_ = new_n1190_ & new_n8360_;
  assign new_n8432_ = new_n1202_ & new_n8360_;
  assign new_n8433_ = ~new_n8431_ & ~new_n8432_;
  assign new_n8434_ = ~new_n8430_ & new_n8433_;
  assign new_n8435_ = new_n8429_ & new_n8434_;
  assign new_n8436_ = new_n1216_ & new_n8360_;
  assign new_n8437_ = new_n1200_ & new_n8360_;
  assign new_n8438_ = new_n1213_ & new_n8360_;
  assign new_n8439_ = ~new_n8437_ & ~new_n8438_;
  assign new_n8440_ = ~new_n8436_ & new_n8439_;
  assign new_n8441_ = new_n1229_ & new_n8360_;
  assign new_n8442_ = new_n1210_ & new_n8360_;
  assign new_n8443_ = new_n1226_ & new_n8360_;
  assign new_n8444_ = ~new_n8442_ & ~new_n8443_;
  assign new_n8445_ = ~new_n8441_ & new_n8444_;
  assign new_n8446_ = new_n8440_ & new_n8445_;
  assign new_n8447_ = new_n8435_ & new_n8446_;
  assign new_n8448_ = new_n1237_ & new_n8360_;
  assign new_n8449_ = new_n1223_ & new_n8360_;
  assign new_n8450_ = new_n1235_ & new_n8360_;
  assign new_n8451_ = ~new_n8449_ & ~new_n8450_;
  assign new_n8452_ = ~new_n8448_ & new_n8451_;
  assign new_n8453_ = new_n7544_ & new_n7966_;
  assign new_n8454_ = new_n951_ & new_n8453_;
  assign new_n8455_ = new_n1233_ & new_n8360_;
  assign new_n8456_ = new_n1243_ & new_n8360_;
  assign new_n8457_ = ~new_n8455_ & ~new_n8456_;
  assign new_n8458_ = ~new_n8454_ & new_n8457_;
  assign new_n8459_ = new_n8452_ & new_n8458_;
  assign new_n8460_ = new_n964_ & new_n8453_;
  assign new_n8461_ = new_n954_ & new_n8453_;
  assign new_n8462_ = new_n948_ & new_n8453_;
  assign new_n8463_ = ~new_n8461_ & ~new_n8462_;
  assign new_n8464_ = ~new_n8460_ & new_n8463_;
  assign new_n8465_ = new_n967_ & new_n8453_;
  assign new_n8466_ = new_n961_ & new_n8453_;
  assign new_n8467_ = ~new_n8465_ & ~new_n8466_;
  assign new_n8468_ = new_n8464_ & new_n8467_;
  assign new_n8469_ = new_n8459_ & new_n8468_;
  assign new_n8470_ = new_n8447_ & new_n8469_;
  assign new_n8471_ = new_n972_ & new_n8453_;
  assign new_n8472_ = new_n975_ & new_n8453_;
  assign new_n8473_ = new_n978_ & new_n8453_;
  assign new_n8474_ = ~new_n8472_ & ~new_n8473_;
  assign new_n8475_ = ~new_n8471_ & new_n8474_;
  assign new_n8476_ = new_n984_ & new_n8453_;
  assign new_n8477_ = new_n987_ & new_n8453_;
  assign new_n8478_ = new_n990_ & new_n8453_;
  assign new_n8479_ = ~new_n8477_ & ~new_n8478_;
  assign new_n8480_ = ~new_n8476_ & new_n8479_;
  assign new_n8481_ = new_n8475_ & new_n8480_;
  assign new_n8482_ = new_n1008_ & new_n8453_;
  assign new_n8483_ = new_n994_ & new_n8453_;
  assign new_n8484_ = new_n996_ & new_n8453_;
  assign new_n8485_ = ~new_n8483_ & ~new_n8484_;
  assign new_n8486_ = ~new_n8482_ & new_n8485_;
  assign new_n8487_ = new_n1016_ & new_n8453_;
  assign new_n8488_ = new_n1010_ & new_n8453_;
  assign new_n8489_ = new_n1006_ & new_n8453_;
  assign new_n8490_ = ~new_n8488_ & ~new_n8489_;
  assign new_n8491_ = ~new_n8487_ & new_n8490_;
  assign new_n8492_ = new_n8486_ & new_n8491_;
  assign new_n8493_ = new_n8481_ & new_n8492_;
  assign new_n8494_ = new_n1025_ & new_n8453_;
  assign new_n8495_ = new_n1018_ & new_n8453_;
  assign new_n8496_ = new_n1014_ & new_n8453_;
  assign new_n8497_ = ~new_n8495_ & ~new_n8496_;
  assign new_n8498_ = ~new_n8494_ & new_n8497_;
  assign new_n8499_ = new_n1033_ & new_n8453_;
  assign new_n8500_ = new_n1027_ & new_n8453_;
  assign new_n8501_ = new_n1023_ & new_n8453_;
  assign new_n8502_ = ~new_n8500_ & ~new_n8501_;
  assign new_n8503_ = ~new_n8499_ & new_n8502_;
  assign new_n8504_ = new_n8498_ & new_n8503_;
  assign new_n8505_ = new_n1043_ & new_n8453_;
  assign new_n8506_ = new_n1035_ & new_n8453_;
  assign new_n8507_ = new_n1031_ & new_n8453_;
  assign new_n8508_ = ~new_n8506_ & ~new_n8507_;
  assign new_n8509_ = ~new_n8505_ & new_n8508_;
  assign new_n8510_ = new_n1045_ & new_n8453_;
  assign new_n8511_ = new_n1041_ & new_n8453_;
  assign new_n8512_ = ~new_n8510_ & ~new_n8511_;
  assign new_n8513_ = new_n8509_ & new_n8512_;
  assign new_n8514_ = new_n8504_ & new_n8513_;
  assign new_n8515_ = new_n8493_ & new_n8514_;
  assign new_n8516_ = new_n8470_ & new_n8515_;
  assign new_n8517_ = new_n1049_ & new_n8453_;
  assign new_n8518_ = new_n1051_ & new_n8453_;
  assign new_n8519_ = new_n1053_ & new_n8453_;
  assign new_n8520_ = ~new_n8518_ & ~new_n8519_;
  assign new_n8521_ = ~new_n8517_ & new_n8520_;
  assign new_n8522_ = new_n7609_ & new_n7966_;
  assign new_n8523_ = new_n1059_ & new_n8522_;
  assign new_n8524_ = new_n1065_ & new_n8522_;
  assign new_n8525_ = new_n1071_ & new_n8522_;
  assign new_n8526_ = ~new_n8524_ & ~new_n8525_;
  assign new_n8527_ = ~new_n8523_ & new_n8526_;
  assign new_n8528_ = new_n8521_ & new_n8527_;
  assign new_n8529_ = new_n1076_ & new_n8522_;
  assign new_n8530_ = new_n1079_ & new_n8522_;
  assign new_n8531_ = new_n1082_ & new_n8522_;
  assign new_n8532_ = ~new_n8530_ & ~new_n8531_;
  assign new_n8533_ = ~new_n8529_ & new_n8532_;
  assign new_n8534_ = new_n1089_ & new_n8522_;
  assign new_n8535_ = new_n1095_ & new_n8522_;
  assign new_n8536_ = new_n1099_ & new_n8522_;
  assign new_n8537_ = ~new_n8535_ & ~new_n8536_;
  assign new_n8538_ = ~new_n8534_ & new_n8537_;
  assign new_n8539_ = new_n8533_ & new_n8538_;
  assign new_n8540_ = new_n8528_ & new_n8539_;
  assign new_n8541_ = new_n1103_ & new_n8522_;
  assign new_n8542_ = new_n1105_ & new_n8522_;
  assign new_n8543_ = new_n1107_ & new_n8522_;
  assign new_n8544_ = ~new_n8542_ & ~new_n8543_;
  assign new_n8545_ = ~new_n8541_ & new_n8544_;
  assign new_n8546_ = new_n1114_ & new_n8522_;
  assign new_n8547_ = new_n1118_ & new_n8522_;
  assign new_n8548_ = new_n1120_ & new_n8522_;
  assign new_n8549_ = ~new_n8547_ & ~new_n8548_;
  assign new_n8550_ = ~new_n8546_ & new_n8549_;
  assign new_n8551_ = new_n8545_ & new_n8550_;
  assign new_n8552_ = new_n1127_ & new_n8522_;
  assign new_n8553_ = new_n1131_ & new_n8522_;
  assign new_n8554_ = new_n1135_ & new_n8522_;
  assign new_n8555_ = ~new_n8553_ & ~new_n8554_;
  assign new_n8556_ = ~new_n8552_ & new_n8555_;
  assign new_n8557_ = new_n1145_ & new_n8522_;
  assign new_n8558_ = new_n1149_ & new_n8522_;
  assign new_n8559_ = ~new_n8557_ & ~new_n8558_;
  assign new_n8560_ = new_n8556_ & new_n8559_;
  assign new_n8561_ = new_n8551_ & new_n8560_;
  assign new_n8562_ = new_n8540_ & new_n8561_;
  assign new_n8563_ = new_n1157_ & new_n8522_;
  assign new_n8564_ = new_n1141_ & new_n8522_;
  assign new_n8565_ = new_n1155_ & new_n8522_;
  assign new_n8566_ = ~new_n8564_ & ~new_n8565_;
  assign new_n8567_ = ~new_n8563_ & new_n8566_;
  assign new_n8568_ = new_n1168_ & new_n8522_;
  assign new_n8569_ = new_n1153_ & new_n8522_;
  assign new_n8570_ = new_n1165_ & new_n8522_;
  assign new_n8571_ = ~new_n8569_ & ~new_n8570_;
  assign new_n8572_ = ~new_n8568_ & new_n8571_;
  assign new_n8573_ = new_n8567_ & new_n8572_;
  assign new_n8574_ = new_n1174_ & new_n8522_;
  assign new_n8575_ = new_n1162_ & new_n8522_;
  assign new_n8576_ = new_n1172_ & new_n8522_;
  assign new_n8577_ = ~new_n8575_ & ~new_n8576_;
  assign new_n8578_ = ~new_n8574_ & new_n8577_;
  assign new_n8579_ = new_n1182_ & new_n8522_;
  assign new_n8580_ = new_n1184_ & new_n8522_;
  assign new_n8581_ = new_n1186_ & new_n8522_;
  assign new_n8582_ = ~new_n8580_ & ~new_n8581_;
  assign new_n8583_ = ~new_n8579_ & new_n8582_;
  assign new_n8584_ = new_n8578_ & new_n8583_;
  assign new_n8585_ = new_n8573_ & new_n8584_;
  assign new_n8586_ = new_n1190_ & new_n8522_;
  assign new_n8587_ = new_n1192_ & new_n8522_;
  assign new_n8588_ = new_n1194_ & new_n8522_;
  assign new_n8589_ = ~new_n8587_ & ~new_n8588_;
  assign new_n8590_ = ~new_n8586_ & new_n8589_;
  assign new_n8591_ = new_n1200_ & new_n8522_;
  assign new_n8592_ = new_n1202_ & new_n8522_;
  assign new_n8593_ = new_n1204_ & new_n8522_;
  assign new_n8594_ = ~new_n8592_ & ~new_n8593_;
  assign new_n8595_ = ~new_n8591_ & new_n8594_;
  assign new_n8596_ = new_n8590_ & new_n8595_;
  assign new_n8597_ = new_n1210_ & new_n8522_;
  assign new_n8598_ = new_n1213_ & new_n8522_;
  assign new_n8599_ = new_n1216_ & new_n8522_;
  assign new_n8600_ = ~new_n8598_ & ~new_n8599_;
  assign new_n8601_ = ~new_n8597_ & new_n8600_;
  assign new_n8602_ = new_n1226_ & new_n8522_;
  assign new_n8603_ = new_n1229_ & new_n8522_;
  assign new_n8604_ = ~new_n8602_ & ~new_n8603_;
  assign new_n8605_ = new_n8601_ & new_n8604_;
  assign new_n8606_ = new_n8596_ & new_n8605_;
  assign new_n8607_ = new_n8585_ & new_n8606_;
  assign new_n8608_ = new_n8562_ & new_n8607_;
  assign new_n8609_ = new_n8516_ & new_n8608_;
  assign new_n8610_ = new_n8424_ & new_n8609_;
  assign new_n8611_ = new_n1237_ & new_n8522_;
  assign new_n8612_ = new_n1223_ & new_n8522_;
  assign new_n8613_ = new_n1235_ & new_n8522_;
  assign new_n8614_ = ~new_n8612_ & ~new_n8613_;
  assign new_n8615_ = ~new_n8611_ & new_n8614_;
  assign new_n8616_ = ~A265 & new_n1063_;
  assign new_n8617_ = new_n1062_ & new_n8616_;
  assign new_n8618_ = new_n4256_ & new_n8617_;
  assign new_n8619_ = new_n1233_ & new_n8522_;
  assign new_n8620_ = new_n1243_ & new_n8522_;
  assign new_n8621_ = ~new_n8619_ & ~new_n8620_;
  assign new_n8622_ = ~new_n8618_ & new_n8621_;
  assign new_n8623_ = new_n8615_ & new_n8622_;
  assign new_n8624_ = A265 & new_n46_;
  assign new_n8625_ = new_n1078_ & new_n8624_;
  assign new_n8626_ = new_n4256_ & new_n8625_;
  assign new_n8627_ = ~A265 & new_n1069_;
  assign new_n8628_ = new_n1068_ & new_n8627_;
  assign new_n8629_ = new_n4256_ & new_n8628_;
  assign new_n8630_ = new_n1058_ & new_n8624_;
  assign new_n8631_ = new_n4256_ & new_n8630_;
  assign new_n8632_ = ~new_n8629_ & ~new_n8631_;
  assign new_n8633_ = ~new_n8626_ & new_n8632_;
  assign new_n8634_ = A265 & new_n1093_;
  assign new_n8635_ = new_n1092_ & new_n8634_;
  assign new_n8636_ = new_n4256_ & new_n8635_;
  assign new_n8637_ = new_n1081_ & new_n8624_;
  assign new_n8638_ = new_n4256_ & new_n8637_;
  assign new_n8639_ = new_n1075_ & new_n8624_;
  assign new_n8640_ = new_n4256_ & new_n8639_;
  assign new_n8641_ = ~new_n8638_ & ~new_n8640_;
  assign new_n8642_ = ~new_n8636_ & new_n8641_;
  assign new_n8643_ = new_n8633_ & new_n8642_;
  assign new_n8644_ = new_n8623_ & new_n8643_;
  assign new_n8645_ = ~A265 & new_n51_;
  assign new_n8646_ = new_n1078_ & new_n8645_;
  assign new_n8647_ = new_n4256_ & new_n8646_;
  assign new_n8648_ = new_n1098_ & new_n8634_;
  assign new_n8649_ = new_n4256_ & new_n8648_;
  assign new_n8650_ = new_n1058_ & new_n8645_;
  assign new_n8651_ = new_n4256_ & new_n8650_;
  assign new_n8652_ = ~new_n8649_ & ~new_n8651_;
  assign new_n8653_ = ~new_n8647_ & new_n8652_;
  assign new_n8654_ = ~A265 & new_n1116_;
  assign new_n8655_ = new_n1092_ & new_n8654_;
  assign new_n8656_ = new_n4256_ & new_n8655_;
  assign new_n8657_ = new_n1081_ & new_n8645_;
  assign new_n8658_ = new_n4256_ & new_n8657_;
  assign new_n8659_ = new_n1075_ & new_n8645_;
  assign new_n8660_ = new_n4256_ & new_n8659_;
  assign new_n8661_ = ~new_n8658_ & ~new_n8660_;
  assign new_n8662_ = ~new_n8656_ & new_n8661_;
  assign new_n8663_ = new_n8653_ & new_n8662_;
  assign new_n8664_ = A265 & new_n1129_;
  assign new_n8665_ = new_n1068_ & new_n8664_;
  assign new_n8666_ = new_n4256_ & new_n8665_;
  assign new_n8667_ = new_n1098_ & new_n8654_;
  assign new_n8668_ = new_n4256_ & new_n8667_;
  assign new_n8669_ = A265 & new_n1112_;
  assign new_n8670_ = new_n1062_ & new_n8669_;
  assign new_n8671_ = new_n4256_ & new_n8670_;
  assign new_n8672_ = ~new_n8668_ & ~new_n8671_;
  assign new_n8673_ = ~new_n8666_ & new_n8672_;
  assign new_n8674_ = ~A267 & new_n1143_;
  assign new_n8675_ = new_n1062_ & new_n8674_;
  assign new_n8676_ = new_n4256_ & new_n8675_;
  assign new_n8677_ = ~A267 & new_n1133_;
  assign new_n8678_ = new_n1062_ & new_n8677_;
  assign new_n8679_ = new_n4256_ & new_n8678_;
  assign new_n8680_ = ~A267 & new_n1124_;
  assign new_n8681_ = new_n1068_ & new_n8680_;
  assign new_n8682_ = new_n4256_ & new_n8681_;
  assign new_n8683_ = ~new_n8679_ & ~new_n8682_;
  assign new_n8684_ = ~new_n8676_ & new_n8683_;
  assign new_n8685_ = new_n8673_ & new_n8684_;
  assign new_n8686_ = new_n8663_ & new_n8685_;
  assign new_n8687_ = new_n8644_ & new_n8686_;
  assign new_n8688_ = A267 & new_n31_;
  assign new_n8689_ = new_n953_ & new_n8688_;
  assign new_n8690_ = new_n4256_ & new_n8689_;
  assign new_n8691_ = ~A267 & new_n1147_;
  assign new_n8692_ = new_n1068_ & new_n8691_;
  assign new_n8693_ = new_n4256_ & new_n8692_;
  assign new_n8694_ = new_n950_ & new_n8688_;
  assign new_n8695_ = new_n4256_ & new_n8694_;
  assign new_n8696_ = ~new_n8693_ & ~new_n8695_;
  assign new_n8697_ = ~new_n8690_ & new_n8696_;
  assign new_n8698_ = new_n4270_ & new_n8617_;
  assign new_n8699_ = new_n947_ & new_n8688_;
  assign new_n8700_ = new_n4256_ & new_n8699_;
  assign new_n8701_ = new_n963_ & new_n8688_;
  assign new_n8702_ = new_n4256_ & new_n8701_;
  assign new_n8703_ = ~new_n8700_ & ~new_n8702_;
  assign new_n8704_ = ~new_n8698_ & new_n8703_;
  assign new_n8705_ = new_n8697_ & new_n8704_;
  assign new_n8706_ = new_n4270_ & new_n8625_;
  assign new_n8707_ = new_n4270_ & new_n8628_;
  assign new_n8708_ = new_n4270_ & new_n8630_;
  assign new_n8709_ = ~new_n8707_ & ~new_n8708_;
  assign new_n8710_ = ~new_n8706_ & new_n8709_;
  assign new_n8711_ = new_n4270_ & new_n8635_;
  assign new_n8712_ = new_n4270_ & new_n8637_;
  assign new_n8713_ = new_n4270_ & new_n8639_;
  assign new_n8714_ = ~new_n8712_ & ~new_n8713_;
  assign new_n8715_ = ~new_n8711_ & new_n8714_;
  assign new_n8716_ = new_n8710_ & new_n8715_;
  assign new_n8717_ = new_n8705_ & new_n8716_;
  assign new_n8718_ = new_n4270_ & new_n8646_;
  assign new_n8719_ = new_n4270_ & new_n8648_;
  assign new_n8720_ = new_n4270_ & new_n8650_;
  assign new_n8721_ = ~new_n8719_ & ~new_n8720_;
  assign new_n8722_ = ~new_n8718_ & new_n8721_;
  assign new_n8723_ = new_n4270_ & new_n8655_;
  assign new_n8724_ = new_n4270_ & new_n8657_;
  assign new_n8725_ = new_n4270_ & new_n8659_;
  assign new_n8726_ = ~new_n8724_ & ~new_n8725_;
  assign new_n8727_ = ~new_n8723_ & new_n8726_;
  assign new_n8728_ = new_n8722_ & new_n8727_;
  assign new_n8729_ = new_n4270_ & new_n8665_;
  assign new_n8730_ = new_n4270_ & new_n8667_;
  assign new_n8731_ = new_n4270_ & new_n8670_;
  assign new_n8732_ = ~new_n8730_ & ~new_n8731_;
  assign new_n8733_ = ~new_n8729_ & new_n8732_;
  assign new_n8734_ = new_n4270_ & new_n8678_;
  assign new_n8735_ = new_n4270_ & new_n8681_;
  assign new_n8736_ = ~new_n8734_ & ~new_n8735_;
  assign new_n8737_ = new_n8733_ & new_n8736_;
  assign new_n8738_ = new_n8728_ & new_n8737_;
  assign new_n8739_ = new_n8717_ & new_n8738_;
  assign new_n8740_ = new_n8687_ & new_n8739_;
  assign new_n8741_ = new_n4270_ & new_n8694_;
  assign new_n8742_ = new_n4270_ & new_n8675_;
  assign new_n8743_ = new_n4270_ & new_n8692_;
  assign new_n8744_ = ~new_n8742_ & ~new_n8743_;
  assign new_n8745_ = ~new_n8741_ & new_n8744_;
  assign new_n8746_ = new_n4270_ & new_n8701_;
  assign new_n8747_ = new_n4270_ & new_n8689_;
  assign new_n8748_ = new_n4270_ & new_n8699_;
  assign new_n8749_ = ~new_n8747_ & ~new_n8748_;
  assign new_n8750_ = ~new_n8746_ & new_n8749_;
  assign new_n8751_ = new_n8745_ & new_n8750_;
  assign new_n8752_ = new_n4278_ & new_n8630_;
  assign new_n8753_ = new_n4278_ & new_n8617_;
  assign new_n8754_ = new_n4278_ & new_n8628_;
  assign new_n8755_ = ~new_n8753_ & ~new_n8754_;
  assign new_n8756_ = ~new_n8752_ & new_n8755_;
  assign new_n8757_ = new_n4278_ & new_n8639_;
  assign new_n8758_ = new_n4278_ & new_n8625_;
  assign new_n8759_ = new_n4278_ & new_n8637_;
  assign new_n8760_ = ~new_n8758_ & ~new_n8759_;
  assign new_n8761_ = ~new_n8757_ & new_n8760_;
  assign new_n8762_ = new_n8756_ & new_n8761_;
  assign new_n8763_ = new_n8751_ & new_n8762_;
  assign new_n8764_ = new_n4278_ & new_n8650_;
  assign new_n8765_ = new_n4278_ & new_n8635_;
  assign new_n8766_ = new_n4278_ & new_n8648_;
  assign new_n8767_ = ~new_n8765_ & ~new_n8766_;
  assign new_n8768_ = ~new_n8764_ & new_n8767_;
  assign new_n8769_ = new_n4278_ & new_n8659_;
  assign new_n8770_ = new_n4278_ & new_n8646_;
  assign new_n8771_ = new_n4278_ & new_n8657_;
  assign new_n8772_ = ~new_n8770_ & ~new_n8771_;
  assign new_n8773_ = ~new_n8769_ & new_n8772_;
  assign new_n8774_ = new_n8768_ & new_n8773_;
  assign new_n8775_ = new_n4278_ & new_n8670_;
  assign new_n8776_ = new_n4278_ & new_n8655_;
  assign new_n8777_ = new_n4278_ & new_n8667_;
  assign new_n8778_ = ~new_n8776_ & ~new_n8777_;
  assign new_n8779_ = ~new_n8775_ & new_n8778_;
  assign new_n8780_ = new_n4278_ & new_n8665_;
  assign new_n8781_ = new_n4278_ & new_n8678_;
  assign new_n8782_ = ~new_n8780_ & ~new_n8781_;
  assign new_n8783_ = new_n8779_ & new_n8782_;
  assign new_n8784_ = new_n8774_ & new_n8783_;
  assign new_n8785_ = new_n8763_ & new_n8784_;
  assign new_n8786_ = new_n4278_ & new_n8692_;
  assign new_n8787_ = new_n4278_ & new_n8681_;
  assign new_n8788_ = new_n4278_ & new_n8675_;
  assign new_n8789_ = ~new_n8787_ & ~new_n8788_;
  assign new_n8790_ = ~new_n8786_ & new_n8789_;
  assign new_n8791_ = new_n4278_ & new_n8699_;
  assign new_n8792_ = new_n4278_ & new_n8694_;
  assign new_n8793_ = new_n4278_ & new_n8689_;
  assign new_n8794_ = ~new_n8792_ & ~new_n8793_;
  assign new_n8795_ = ~new_n8791_ & new_n8794_;
  assign new_n8796_ = new_n8790_ & new_n8795_;
  assign new_n8797_ = new_n4295_ & new_n8628_;
  assign new_n8798_ = new_n4278_ & new_n8701_;
  assign new_n8799_ = new_n4295_ & new_n8617_;
  assign new_n8800_ = ~new_n8798_ & ~new_n8799_;
  assign new_n8801_ = ~new_n8797_ & new_n8800_;
  assign new_n8802_ = new_n4295_ & new_n8637_;
  assign new_n8803_ = new_n4295_ & new_n8630_;
  assign new_n8804_ = new_n4295_ & new_n8625_;
  assign new_n8805_ = ~new_n8803_ & ~new_n8804_;
  assign new_n8806_ = ~new_n8802_ & new_n8805_;
  assign new_n8807_ = new_n8801_ & new_n8806_;
  assign new_n8808_ = new_n8796_ & new_n8807_;
  assign new_n8809_ = new_n4295_ & new_n8648_;
  assign new_n8810_ = new_n4295_ & new_n8639_;
  assign new_n8811_ = new_n4295_ & new_n8635_;
  assign new_n8812_ = ~new_n8810_ & ~new_n8811_;
  assign new_n8813_ = ~new_n8809_ & new_n8812_;
  assign new_n8814_ = new_n4295_ & new_n8657_;
  assign new_n8815_ = new_n4295_ & new_n8650_;
  assign new_n8816_ = new_n4295_ & new_n8646_;
  assign new_n8817_ = ~new_n8815_ & ~new_n8816_;
  assign new_n8818_ = ~new_n8814_ & new_n8817_;
  assign new_n8819_ = new_n8813_ & new_n8818_;
  assign new_n8820_ = new_n4295_ & new_n8667_;
  assign new_n8821_ = new_n4295_ & new_n8659_;
  assign new_n8822_ = new_n4295_ & new_n8655_;
  assign new_n8823_ = ~new_n8821_ & ~new_n8822_;
  assign new_n8824_ = ~new_n8820_ & new_n8823_;
  assign new_n8825_ = new_n4295_ & new_n8670_;
  assign new_n8826_ = new_n4295_ & new_n8665_;
  assign new_n8827_ = ~new_n8825_ & ~new_n8826_;
  assign new_n8828_ = new_n8824_ & new_n8827_;
  assign new_n8829_ = new_n8819_ & new_n8828_;
  assign new_n8830_ = new_n8808_ & new_n8829_;
  assign new_n8831_ = new_n8785_ & new_n8830_;
  assign new_n8832_ = new_n8740_ & new_n8831_;
  assign new_n8833_ = new_n4295_ & new_n8675_;
  assign new_n8834_ = new_n4295_ & new_n8678_;
  assign new_n8835_ = new_n4295_ & new_n8681_;
  assign new_n8836_ = ~new_n8834_ & ~new_n8835_;
  assign new_n8837_ = ~new_n8833_ & new_n8836_;
  assign new_n8838_ = new_n4295_ & new_n8689_;
  assign new_n8839_ = new_n4295_ & new_n8692_;
  assign new_n8840_ = new_n4295_ & new_n8694_;
  assign new_n8841_ = ~new_n8839_ & ~new_n8840_;
  assign new_n8842_ = ~new_n8838_ & new_n8841_;
  assign new_n8843_ = new_n8837_ & new_n8842_;
  assign new_n8844_ = A236 & new_n139_;
  assign new_n8845_ = new_n950_ & new_n8844_;
  assign new_n8846_ = new_n4302_ & new_n8845_;
  assign new_n8847_ = new_n4295_ & new_n8699_;
  assign new_n8848_ = new_n4295_ & new_n8701_;
  assign new_n8849_ = ~new_n8847_ & ~new_n8848_;
  assign new_n8850_ = ~new_n8846_ & new_n8849_;
  assign new_n8851_ = new_n963_ & new_n8844_;
  assign new_n8852_ = new_n4302_ & new_n8851_;
  assign new_n8853_ = new_n953_ & new_n8844_;
  assign new_n8854_ = new_n4302_ & new_n8853_;
  assign new_n8855_ = new_n947_ & new_n8844_;
  assign new_n8856_ = new_n4302_ & new_n8855_;
  assign new_n8857_ = ~new_n8854_ & ~new_n8856_;
  assign new_n8858_ = ~new_n8852_ & new_n8857_;
  assign new_n8859_ = new_n8850_ & new_n8858_;
  assign new_n8860_ = new_n8843_ & new_n8859_;
  assign new_n8861_ = A236 & new_n155_;
  assign new_n8862_ = new_n974_ & new_n8861_;
  assign new_n8863_ = new_n4302_ & new_n8862_;
  assign new_n8864_ = new_n966_ & new_n8861_;
  assign new_n8865_ = new_n4302_ & new_n8864_;
  assign new_n8866_ = new_n960_ & new_n8861_;
  assign new_n8867_ = new_n4302_ & new_n8866_;
  assign new_n8868_ = ~new_n8865_ & ~new_n8867_;
  assign new_n8869_ = ~new_n8863_ & new_n8868_;
  assign new_n8870_ = new_n986_ & new_n8861_;
  assign new_n8871_ = new_n4302_ & new_n8870_;
  assign new_n8872_ = new_n977_ & new_n8861_;
  assign new_n8873_ = new_n4302_ & new_n8872_;
  assign new_n8874_ = new_n971_ & new_n8861_;
  assign new_n8875_ = new_n4302_ & new_n8874_;
  assign new_n8876_ = ~new_n8873_ & ~new_n8875_;
  assign new_n8877_ = ~new_n8871_ & new_n8876_;
  assign new_n8878_ = new_n8869_ & new_n8877_;
  assign new_n8879_ = A236 & new_n186_;
  assign new_n8880_ = new_n966_ & new_n8879_;
  assign new_n8881_ = new_n4302_ & new_n8880_;
  assign new_n8882_ = new_n989_ & new_n8861_;
  assign new_n8883_ = new_n4302_ & new_n8882_;
  assign new_n8884_ = new_n983_ & new_n8861_;
  assign new_n8885_ = new_n4302_ & new_n8884_;
  assign new_n8886_ = ~new_n8883_ & ~new_n8885_;
  assign new_n8887_ = ~new_n8881_ & new_n8886_;
  assign new_n8888_ = new_n960_ & new_n8879_;
  assign new_n8889_ = new_n4302_ & new_n8888_;
  assign new_n8890_ = new_n974_ & new_n8879_;
  assign new_n8891_ = new_n4302_ & new_n8890_;
  assign new_n8892_ = ~new_n8889_ & ~new_n8891_;
  assign new_n8893_ = new_n8887_ & new_n8892_;
  assign new_n8894_ = new_n8878_ & new_n8893_;
  assign new_n8895_ = new_n8860_ & new_n8894_;
  assign new_n8896_ = new_n986_ & new_n8879_;
  assign new_n8897_ = new_n4302_ & new_n8896_;
  assign new_n8898_ = new_n977_ & new_n8879_;
  assign new_n8899_ = new_n4302_ & new_n8898_;
  assign new_n8900_ = new_n971_ & new_n8879_;
  assign new_n8901_ = new_n4302_ & new_n8900_;
  assign new_n8902_ = ~new_n8899_ & ~new_n8901_;
  assign new_n8903_ = ~new_n8897_ & new_n8902_;
  assign new_n8904_ = A236 & new_n209_;
  assign new_n8905_ = new_n950_ & new_n8904_;
  assign new_n8906_ = new_n4302_ & new_n8905_;
  assign new_n8907_ = new_n989_ & new_n8879_;
  assign new_n8908_ = new_n4302_ & new_n8907_;
  assign new_n8909_ = new_n983_ & new_n8879_;
  assign new_n8910_ = new_n4302_ & new_n8909_;
  assign new_n8911_ = ~new_n8908_ & ~new_n8910_;
  assign new_n8912_ = ~new_n8906_ & new_n8911_;
  assign new_n8913_ = new_n8903_ & new_n8912_;
  assign new_n8914_ = new_n963_ & new_n8904_;
  assign new_n8915_ = new_n4302_ & new_n8914_;
  assign new_n8916_ = new_n953_ & new_n8904_;
  assign new_n8917_ = new_n4302_ & new_n8916_;
  assign new_n8918_ = new_n947_ & new_n8904_;
  assign new_n8919_ = new_n4302_ & new_n8918_;
  assign new_n8920_ = ~new_n8917_ & ~new_n8919_;
  assign new_n8921_ = ~new_n8915_ & new_n8920_;
  assign new_n8922_ = A236 & new_n218_;
  assign new_n8923_ = new_n947_ & new_n8922_;
  assign new_n8924_ = new_n4302_ & new_n8923_;
  assign new_n8925_ = new_n950_ & new_n8922_;
  assign new_n8926_ = new_n4302_ & new_n8925_;
  assign new_n8927_ = new_n953_ & new_n8922_;
  assign new_n8928_ = new_n4302_ & new_n8927_;
  assign new_n8929_ = ~new_n8926_ & ~new_n8928_;
  assign new_n8930_ = ~new_n8924_ & new_n8929_;
  assign new_n8931_ = new_n8921_ & new_n8930_;
  assign new_n8932_ = new_n8913_ & new_n8931_;
  assign new_n8933_ = A236 & new_n236_;
  assign new_n8934_ = new_n953_ & new_n8933_;
  assign new_n8935_ = new_n4302_ & new_n8934_;
  assign new_n8936_ = new_n963_ & new_n8922_;
  assign new_n8937_ = new_n4302_ & new_n8936_;
  assign new_n8938_ = new_n950_ & new_n8933_;
  assign new_n8939_ = new_n4302_ & new_n8938_;
  assign new_n8940_ = ~new_n8937_ & ~new_n8939_;
  assign new_n8941_ = ~new_n8935_ & new_n8940_;
  assign new_n8942_ = new_n4352_ & new_n8617_;
  assign new_n8943_ = new_n947_ & new_n8933_;
  assign new_n8944_ = new_n4302_ & new_n8943_;
  assign new_n8945_ = new_n963_ & new_n8933_;
  assign new_n8946_ = new_n4302_ & new_n8945_;
  assign new_n8947_ = ~new_n8944_ & ~new_n8946_;
  assign new_n8948_ = ~new_n8942_ & new_n8947_;
  assign new_n8949_ = new_n8941_ & new_n8948_;
  assign new_n8950_ = new_n4352_ & new_n8625_;
  assign new_n8951_ = new_n4352_ & new_n8628_;
  assign new_n8952_ = new_n4352_ & new_n8630_;
  assign new_n8953_ = ~new_n8951_ & ~new_n8952_;
  assign new_n8954_ = ~new_n8950_ & new_n8953_;
  assign new_n8955_ = new_n4352_ & new_n8637_;
  assign new_n8956_ = new_n4352_ & new_n8639_;
  assign new_n8957_ = ~new_n8955_ & ~new_n8956_;
  assign new_n8958_ = new_n8954_ & new_n8957_;
  assign new_n8959_ = new_n8949_ & new_n8958_;
  assign new_n8960_ = new_n8932_ & new_n8959_;
  assign new_n8961_ = new_n8895_ & new_n8960_;
  assign new_n8962_ = new_n4352_ & new_n8650_;
  assign new_n8963_ = new_n4352_ & new_n8635_;
  assign new_n8964_ = new_n4352_ & new_n8648_;
  assign new_n8965_ = ~new_n8963_ & ~new_n8964_;
  assign new_n8966_ = ~new_n8962_ & new_n8965_;
  assign new_n8967_ = new_n4352_ & new_n8659_;
  assign new_n8968_ = new_n4352_ & new_n8646_;
  assign new_n8969_ = new_n4352_ & new_n8657_;
  assign new_n8970_ = ~new_n8968_ & ~new_n8969_;
  assign new_n8971_ = ~new_n8967_ & new_n8970_;
  assign new_n8972_ = new_n8966_ & new_n8971_;
  assign new_n8973_ = new_n4352_ & new_n8670_;
  assign new_n8974_ = new_n4352_ & new_n8655_;
  assign new_n8975_ = new_n4352_ & new_n8667_;
  assign new_n8976_ = ~new_n8974_ & ~new_n8975_;
  assign new_n8977_ = ~new_n8973_ & new_n8976_;
  assign new_n8978_ = new_n4352_ & new_n8681_;
  assign new_n8979_ = new_n4352_ & new_n8665_;
  assign new_n8980_ = new_n4352_ & new_n8678_;
  assign new_n8981_ = ~new_n8979_ & ~new_n8980_;
  assign new_n8982_ = ~new_n8978_ & new_n8981_;
  assign new_n8983_ = new_n8977_ & new_n8982_;
  assign new_n8984_ = new_n8972_ & new_n8983_;
  assign new_n8985_ = new_n4352_ & new_n8694_;
  assign new_n8986_ = new_n4352_ & new_n8675_;
  assign new_n8987_ = new_n4352_ & new_n8692_;
  assign new_n8988_ = ~new_n8986_ & ~new_n8987_;
  assign new_n8989_ = ~new_n8985_ & new_n8988_;
  assign new_n8990_ = new_n4352_ & new_n8701_;
  assign new_n8991_ = new_n4352_ & new_n8689_;
  assign new_n8992_ = new_n4352_ & new_n8699_;
  assign new_n8993_ = ~new_n8991_ & ~new_n8992_;
  assign new_n8994_ = ~new_n8990_ & new_n8993_;
  assign new_n8995_ = new_n8989_ & new_n8994_;
  assign new_n8996_ = new_n4360_ & new_n8630_;
  assign new_n8997_ = new_n4360_ & new_n8617_;
  assign new_n8998_ = new_n4360_ & new_n8628_;
  assign new_n8999_ = ~new_n8997_ & ~new_n8998_;
  assign new_n9000_ = ~new_n8996_ & new_n8999_;
  assign new_n9001_ = new_n4360_ & new_n8625_;
  assign new_n9002_ = new_n4360_ & new_n8637_;
  assign new_n9003_ = ~new_n9001_ & ~new_n9002_;
  assign new_n9004_ = new_n9000_ & new_n9003_;
  assign new_n9005_ = new_n8995_ & new_n9004_;
  assign new_n9006_ = new_n8984_ & new_n9005_;
  assign new_n9007_ = new_n4360_ & new_n8648_;
  assign new_n9008_ = new_n4360_ & new_n8639_;
  assign new_n9009_ = new_n4360_ & new_n8635_;
  assign new_n9010_ = ~new_n9008_ & ~new_n9009_;
  assign new_n9011_ = ~new_n9007_ & new_n9010_;
  assign new_n9012_ = new_n4360_ & new_n8657_;
  assign new_n9013_ = new_n4360_ & new_n8650_;
  assign new_n9014_ = new_n4360_ & new_n8646_;
  assign new_n9015_ = ~new_n9013_ & ~new_n9014_;
  assign new_n9016_ = ~new_n9012_ & new_n9015_;
  assign new_n9017_ = new_n9011_ & new_n9016_;
  assign new_n9018_ = new_n4360_ & new_n8667_;
  assign new_n9019_ = new_n4360_ & new_n8659_;
  assign new_n9020_ = new_n4360_ & new_n8655_;
  assign new_n9021_ = ~new_n9019_ & ~new_n9020_;
  assign new_n9022_ = ~new_n9018_ & new_n9021_;
  assign new_n9023_ = new_n4360_ & new_n8678_;
  assign new_n9024_ = new_n4360_ & new_n8670_;
  assign new_n9025_ = new_n4360_ & new_n8665_;
  assign new_n9026_ = ~new_n9024_ & ~new_n9025_;
  assign new_n9027_ = ~new_n9023_ & new_n9026_;
  assign new_n9028_ = new_n9022_ & new_n9027_;
  assign new_n9029_ = new_n9017_ & new_n9028_;
  assign new_n9030_ = new_n4360_ & new_n8692_;
  assign new_n9031_ = new_n4360_ & new_n8681_;
  assign new_n9032_ = new_n4360_ & new_n8675_;
  assign new_n9033_ = ~new_n9031_ & ~new_n9032_;
  assign new_n9034_ = ~new_n9030_ & new_n9033_;
  assign new_n9035_ = new_n4360_ & new_n8699_;
  assign new_n9036_ = new_n4360_ & new_n8694_;
  assign new_n9037_ = new_n4360_ & new_n8689_;
  assign new_n9038_ = ~new_n9036_ & ~new_n9037_;
  assign new_n9039_ = ~new_n9035_ & new_n9038_;
  assign new_n9040_ = new_n9034_ & new_n9039_;
  assign new_n9041_ = new_n4374_ & new_n8628_;
  assign new_n9042_ = new_n4360_ & new_n8701_;
  assign new_n9043_ = new_n4374_ & new_n8617_;
  assign new_n9044_ = ~new_n9042_ & ~new_n9043_;
  assign new_n9045_ = ~new_n9041_ & new_n9044_;
  assign new_n9046_ = new_n4374_ & new_n8630_;
  assign new_n9047_ = new_n4374_ & new_n8625_;
  assign new_n9048_ = ~new_n9046_ & ~new_n9047_;
  assign new_n9049_ = new_n9045_ & new_n9048_;
  assign new_n9050_ = new_n9040_ & new_n9049_;
  assign new_n9051_ = new_n9029_ & new_n9050_;
  assign new_n9052_ = new_n9006_ & new_n9051_;
  assign new_n9053_ = new_n8961_ & new_n9052_;
  assign new_n9054_ = new_n8832_ & new_n9053_;
  assign new_n9055_ = new_n8610_ & new_n9054_;
  assign new_n9056_ = new_n4374_ & new_n8635_;
  assign new_n9057_ = new_n4374_ & new_n8637_;
  assign new_n9058_ = new_n4374_ & new_n8639_;
  assign new_n9059_ = ~new_n9057_ & ~new_n9058_;
  assign new_n9060_ = ~new_n9056_ & new_n9059_;
  assign new_n9061_ = new_n4374_ & new_n8646_;
  assign new_n9062_ = new_n4374_ & new_n8648_;
  assign new_n9063_ = new_n4374_ & new_n8650_;
  assign new_n9064_ = ~new_n9062_ & ~new_n9063_;
  assign new_n9065_ = ~new_n9061_ & new_n9064_;
  assign new_n9066_ = new_n9060_ & new_n9065_;
  assign new_n9067_ = new_n4374_ & new_n8655_;
  assign new_n9068_ = new_n4374_ & new_n8657_;
  assign new_n9069_ = new_n4374_ & new_n8659_;
  assign new_n9070_ = ~new_n9068_ & ~new_n9069_;
  assign new_n9071_ = ~new_n9067_ & new_n9070_;
  assign new_n9072_ = new_n4374_ & new_n8665_;
  assign new_n9073_ = new_n4374_ & new_n8667_;
  assign new_n9074_ = new_n4374_ & new_n8670_;
  assign new_n9075_ = ~new_n9073_ & ~new_n9074_;
  assign new_n9076_ = ~new_n9072_ & new_n9075_;
  assign new_n9077_ = new_n9071_ & new_n9076_;
  assign new_n9078_ = new_n9066_ & new_n9077_;
  assign new_n9079_ = new_n4374_ & new_n8675_;
  assign new_n9080_ = new_n4374_ & new_n8678_;
  assign new_n9081_ = new_n4374_ & new_n8681_;
  assign new_n9082_ = ~new_n9080_ & ~new_n9081_;
  assign new_n9083_ = ~new_n9079_ & new_n9082_;
  assign new_n9084_ = new_n4374_ & new_n8689_;
  assign new_n9085_ = new_n4374_ & new_n8692_;
  assign new_n9086_ = new_n4374_ & new_n8694_;
  assign new_n9087_ = ~new_n9085_ & ~new_n9086_;
  assign new_n9088_ = ~new_n9084_ & new_n9087_;
  assign new_n9089_ = new_n9083_ & new_n9088_;
  assign new_n9090_ = new_n4381_ & new_n8617_;
  assign new_n9091_ = new_n4374_ & new_n8699_;
  assign new_n9092_ = new_n4374_ & new_n8701_;
  assign new_n9093_ = ~new_n9091_ & ~new_n9092_;
  assign new_n9094_ = ~new_n9090_ & new_n9093_;
  assign new_n9095_ = new_n4381_ & new_n8625_;
  assign new_n9096_ = new_n4381_ & new_n8628_;
  assign new_n9097_ = new_n4381_ & new_n8630_;
  assign new_n9098_ = ~new_n9096_ & ~new_n9097_;
  assign new_n9099_ = ~new_n9095_ & new_n9098_;
  assign new_n9100_ = new_n9094_ & new_n9099_;
  assign new_n9101_ = new_n9089_ & new_n9100_;
  assign new_n9102_ = new_n9078_ & new_n9101_;
  assign new_n9103_ = new_n4381_ & new_n8635_;
  assign new_n9104_ = new_n4381_ & new_n8637_;
  assign new_n9105_ = new_n4381_ & new_n8639_;
  assign new_n9106_ = ~new_n9104_ & ~new_n9105_;
  assign new_n9107_ = ~new_n9103_ & new_n9106_;
  assign new_n9108_ = new_n4381_ & new_n8646_;
  assign new_n9109_ = new_n4381_ & new_n8648_;
  assign new_n9110_ = new_n4381_ & new_n8650_;
  assign new_n9111_ = ~new_n9109_ & ~new_n9110_;
  assign new_n9112_ = ~new_n9108_ & new_n9111_;
  assign new_n9113_ = new_n9107_ & new_n9112_;
  assign new_n9114_ = new_n4381_ & new_n8655_;
  assign new_n9115_ = new_n4381_ & new_n8657_;
  assign new_n9116_ = new_n4381_ & new_n8659_;
  assign new_n9117_ = ~new_n9115_ & ~new_n9116_;
  assign new_n9118_ = ~new_n9114_ & new_n9117_;
  assign new_n9119_ = new_n4381_ & new_n8665_;
  assign new_n9120_ = new_n4381_ & new_n8667_;
  assign new_n9121_ = new_n4381_ & new_n8670_;
  assign new_n9122_ = ~new_n9120_ & ~new_n9121_;
  assign new_n9123_ = ~new_n9119_ & new_n9122_;
  assign new_n9124_ = new_n9118_ & new_n9123_;
  assign new_n9125_ = new_n9113_ & new_n9124_;
  assign new_n9126_ = new_n4381_ & new_n8675_;
  assign new_n9127_ = new_n4381_ & new_n8678_;
  assign new_n9128_ = new_n4381_ & new_n8681_;
  assign new_n9129_ = ~new_n9127_ & ~new_n9128_;
  assign new_n9130_ = ~new_n9126_ & new_n9129_;
  assign new_n9131_ = new_n4381_ & new_n8689_;
  assign new_n9132_ = new_n4381_ & new_n8692_;
  assign new_n9133_ = new_n4381_ & new_n8694_;
  assign new_n9134_ = ~new_n9132_ & ~new_n9133_;
  assign new_n9135_ = ~new_n9131_ & new_n9134_;
  assign new_n9136_ = new_n9130_ & new_n9135_;
  assign new_n9137_ = new_n4389_ & new_n8845_;
  assign new_n9138_ = new_n4381_ & new_n8699_;
  assign new_n9139_ = new_n4381_ & new_n8701_;
  assign new_n9140_ = ~new_n9138_ & ~new_n9139_;
  assign new_n9141_ = ~new_n9137_ & new_n9140_;
  assign new_n9142_ = new_n4389_ & new_n8853_;
  assign new_n9143_ = new_n4389_ & new_n8855_;
  assign new_n9144_ = ~new_n9142_ & ~new_n9143_;
  assign new_n9145_ = new_n9141_ & new_n9144_;
  assign new_n9146_ = new_n9136_ & new_n9145_;
  assign new_n9147_ = new_n9125_ & new_n9146_;
  assign new_n9148_ = new_n9102_ & new_n9147_;
  assign new_n9149_ = new_n4389_ & new_n8866_;
  assign new_n9150_ = new_n4389_ & new_n8851_;
  assign new_n9151_ = new_n4389_ & new_n8864_;
  assign new_n9152_ = ~new_n9150_ & ~new_n9151_;
  assign new_n9153_ = ~new_n9149_ & new_n9152_;
  assign new_n9154_ = new_n4389_ & new_n8874_;
  assign new_n9155_ = new_n4389_ & new_n8862_;
  assign new_n9156_ = new_n4389_ & new_n8872_;
  assign new_n9157_ = ~new_n9155_ & ~new_n9156_;
  assign new_n9158_ = ~new_n9154_ & new_n9157_;
  assign new_n9159_ = new_n9153_ & new_n9158_;
  assign new_n9160_ = new_n4389_ & new_n8884_;
  assign new_n9161_ = new_n4389_ & new_n8870_;
  assign new_n9162_ = new_n4389_ & new_n8882_;
  assign new_n9163_ = ~new_n9161_ & ~new_n9162_;
  assign new_n9164_ = ~new_n9160_ & new_n9163_;
  assign new_n9165_ = new_n4389_ & new_n8890_;
  assign new_n9166_ = new_n4389_ & new_n8880_;
  assign new_n9167_ = new_n4389_ & new_n8888_;
  assign new_n9168_ = ~new_n9166_ & ~new_n9167_;
  assign new_n9169_ = ~new_n9165_ & new_n9168_;
  assign new_n9170_ = new_n9164_ & new_n9169_;
  assign new_n9171_ = new_n9159_ & new_n9170_;
  assign new_n9172_ = new_n4389_ & new_n8896_;
  assign new_n9173_ = new_n4389_ & new_n8898_;
  assign new_n9174_ = new_n4389_ & new_n8900_;
  assign new_n9175_ = ~new_n9173_ & ~new_n9174_;
  assign new_n9176_ = ~new_n9172_ & new_n9175_;
  assign new_n9177_ = new_n4389_ & new_n8905_;
  assign new_n9178_ = new_n4389_ & new_n8907_;
  assign new_n9179_ = new_n4389_ & new_n8909_;
  assign new_n9180_ = ~new_n9178_ & ~new_n9179_;
  assign new_n9181_ = ~new_n9177_ & new_n9180_;
  assign new_n9182_ = new_n9176_ & new_n9181_;
  assign new_n9183_ = new_n4389_ & new_n8914_;
  assign new_n9184_ = new_n4389_ & new_n8916_;
  assign new_n9185_ = new_n4389_ & new_n8918_;
  assign new_n9186_ = ~new_n9184_ & ~new_n9185_;
  assign new_n9187_ = ~new_n9183_ & new_n9186_;
  assign new_n9188_ = new_n4389_ & new_n8925_;
  assign new_n9189_ = new_n4389_ & new_n8927_;
  assign new_n9190_ = ~new_n9188_ & ~new_n9189_;
  assign new_n9191_ = new_n9187_ & new_n9190_;
  assign new_n9192_ = new_n9182_ & new_n9191_;
  assign new_n9193_ = new_n9171_ & new_n9192_;
  assign new_n9194_ = new_n4389_ & new_n8938_;
  assign new_n9195_ = new_n4389_ & new_n8923_;
  assign new_n9196_ = new_n4389_ & new_n8936_;
  assign new_n9197_ = ~new_n9195_ & ~new_n9196_;
  assign new_n9198_ = ~new_n9194_ & new_n9197_;
  assign new_n9199_ = new_n4389_ & new_n8945_;
  assign new_n9200_ = new_n4389_ & new_n8934_;
  assign new_n9201_ = new_n4389_ & new_n8943_;
  assign new_n9202_ = ~new_n9200_ & ~new_n9201_;
  assign new_n9203_ = ~new_n9199_ & new_n9202_;
  assign new_n9204_ = new_n9198_ & new_n9203_;
  assign new_n9205_ = new_n4443_ & new_n8630_;
  assign new_n9206_ = new_n4443_ & new_n8617_;
  assign new_n9207_ = new_n4443_ & new_n8628_;
  assign new_n9208_ = ~new_n9206_ & ~new_n9207_;
  assign new_n9209_ = ~new_n9205_ & new_n9208_;
  assign new_n9210_ = new_n4443_ & new_n8639_;
  assign new_n9211_ = new_n4443_ & new_n8625_;
  assign new_n9212_ = new_n4443_ & new_n8637_;
  assign new_n9213_ = ~new_n9211_ & ~new_n9212_;
  assign new_n9214_ = ~new_n9210_ & new_n9213_;
  assign new_n9215_ = new_n9209_ & new_n9214_;
  assign new_n9216_ = new_n9204_ & new_n9215_;
  assign new_n9217_ = new_n4443_ & new_n8650_;
  assign new_n9218_ = new_n4443_ & new_n8635_;
  assign new_n9219_ = new_n4443_ & new_n8648_;
  assign new_n9220_ = ~new_n9218_ & ~new_n9219_;
  assign new_n9221_ = ~new_n9217_ & new_n9220_;
  assign new_n9222_ = new_n4443_ & new_n8659_;
  assign new_n9223_ = new_n4443_ & new_n8646_;
  assign new_n9224_ = new_n4443_ & new_n8657_;
  assign new_n9225_ = ~new_n9223_ & ~new_n9224_;
  assign new_n9226_ = ~new_n9222_ & new_n9225_;
  assign new_n9227_ = new_n9221_ & new_n9226_;
  assign new_n9228_ = new_n4443_ & new_n8670_;
  assign new_n9229_ = new_n4443_ & new_n8655_;
  assign new_n9230_ = new_n4443_ & new_n8667_;
  assign new_n9231_ = ~new_n9229_ & ~new_n9230_;
  assign new_n9232_ = ~new_n9228_ & new_n9231_;
  assign new_n9233_ = new_n4443_ & new_n8665_;
  assign new_n9234_ = new_n4443_ & new_n8678_;
  assign new_n9235_ = ~new_n9233_ & ~new_n9234_;
  assign new_n9236_ = new_n9232_ & new_n9235_;
  assign new_n9237_ = new_n9227_ & new_n9236_;
  assign new_n9238_ = new_n9216_ & new_n9237_;
  assign new_n9239_ = new_n9193_ & new_n9238_;
  assign new_n9240_ = new_n9148_ & new_n9239_;
  assign new_n9241_ = new_n4443_ & new_n8692_;
  assign new_n9242_ = new_n4443_ & new_n8681_;
  assign new_n9243_ = new_n4443_ & new_n8675_;
  assign new_n9244_ = ~new_n9242_ & ~new_n9243_;
  assign new_n9245_ = ~new_n9241_ & new_n9244_;
  assign new_n9246_ = new_n4443_ & new_n8699_;
  assign new_n9247_ = new_n4443_ & new_n8694_;
  assign new_n9248_ = new_n4443_ & new_n8689_;
  assign new_n9249_ = ~new_n9247_ & ~new_n9248_;
  assign new_n9250_ = ~new_n9246_ & new_n9249_;
  assign new_n9251_ = new_n9245_ & new_n9250_;
  assign new_n9252_ = new_n4451_ & new_n8628_;
  assign new_n9253_ = new_n4443_ & new_n8701_;
  assign new_n9254_ = new_n4451_ & new_n8617_;
  assign new_n9255_ = ~new_n9253_ & ~new_n9254_;
  assign new_n9256_ = ~new_n9252_ & new_n9255_;
  assign new_n9257_ = new_n4451_ & new_n8637_;
  assign new_n9258_ = new_n4451_ & new_n8630_;
  assign new_n9259_ = new_n4451_ & new_n8625_;
  assign new_n9260_ = ~new_n9258_ & ~new_n9259_;
  assign new_n9261_ = ~new_n9257_ & new_n9260_;
  assign new_n9262_ = new_n9256_ & new_n9261_;
  assign new_n9263_ = new_n9251_ & new_n9262_;
  assign new_n9264_ = new_n4451_ & new_n8648_;
  assign new_n9265_ = new_n4451_ & new_n8639_;
  assign new_n9266_ = new_n4451_ & new_n8635_;
  assign new_n9267_ = ~new_n9265_ & ~new_n9266_;
  assign new_n9268_ = ~new_n9264_ & new_n9267_;
  assign new_n9269_ = new_n4451_ & new_n8657_;
  assign new_n9270_ = new_n4451_ & new_n8650_;
  assign new_n9271_ = new_n4451_ & new_n8646_;
  assign new_n9272_ = ~new_n9270_ & ~new_n9271_;
  assign new_n9273_ = ~new_n9269_ & new_n9272_;
  assign new_n9274_ = new_n9268_ & new_n9273_;
  assign new_n9275_ = new_n4451_ & new_n8667_;
  assign new_n9276_ = new_n4451_ & new_n8659_;
  assign new_n9277_ = new_n4451_ & new_n8655_;
  assign new_n9278_ = ~new_n9276_ & ~new_n9277_;
  assign new_n9279_ = ~new_n9275_ & new_n9278_;
  assign new_n9280_ = new_n4451_ & new_n8670_;
  assign new_n9281_ = new_n4451_ & new_n8665_;
  assign new_n9282_ = ~new_n9280_ & ~new_n9281_;
  assign new_n9283_ = new_n9279_ & new_n9282_;
  assign new_n9284_ = new_n9274_ & new_n9283_;
  assign new_n9285_ = new_n9263_ & new_n9284_;
  assign new_n9286_ = new_n4451_ & new_n8675_;
  assign new_n9287_ = new_n4451_ & new_n8678_;
  assign new_n9288_ = new_n4451_ & new_n8681_;
  assign new_n9289_ = ~new_n9287_ & ~new_n9288_;
  assign new_n9290_ = ~new_n9286_ & new_n9289_;
  assign new_n9291_ = new_n4451_ & new_n8689_;
  assign new_n9292_ = new_n4451_ & new_n8692_;
  assign new_n9293_ = new_n4451_ & new_n8694_;
  assign new_n9294_ = ~new_n9292_ & ~new_n9293_;
  assign new_n9295_ = ~new_n9291_ & new_n9294_;
  assign new_n9296_ = new_n9290_ & new_n9295_;
  assign new_n9297_ = new_n4464_ & new_n8617_;
  assign new_n9298_ = new_n4451_ & new_n8699_;
  assign new_n9299_ = new_n4451_ & new_n8701_;
  assign new_n9300_ = ~new_n9298_ & ~new_n9299_;
  assign new_n9301_ = ~new_n9297_ & new_n9300_;
  assign new_n9302_ = new_n4464_ & new_n8625_;
  assign new_n9303_ = new_n4464_ & new_n8628_;
  assign new_n9304_ = new_n4464_ & new_n8630_;
  assign new_n9305_ = ~new_n9303_ & ~new_n9304_;
  assign new_n9306_ = ~new_n9302_ & new_n9305_;
  assign new_n9307_ = new_n9301_ & new_n9306_;
  assign new_n9308_ = new_n9296_ & new_n9307_;
  assign new_n9309_ = new_n4464_ & new_n8635_;
  assign new_n9310_ = new_n4464_ & new_n8637_;
  assign new_n9311_ = new_n4464_ & new_n8639_;
  assign new_n9312_ = ~new_n9310_ & ~new_n9311_;
  assign new_n9313_ = ~new_n9309_ & new_n9312_;
  assign new_n9314_ = new_n4464_ & new_n8646_;
  assign new_n9315_ = new_n4464_ & new_n8648_;
  assign new_n9316_ = new_n4464_ & new_n8650_;
  assign new_n9317_ = ~new_n9315_ & ~new_n9316_;
  assign new_n9318_ = ~new_n9314_ & new_n9317_;
  assign new_n9319_ = new_n9313_ & new_n9318_;
  assign new_n9320_ = new_n4464_ & new_n8655_;
  assign new_n9321_ = new_n4464_ & new_n8657_;
  assign new_n9322_ = new_n4464_ & new_n8659_;
  assign new_n9323_ = ~new_n9321_ & ~new_n9322_;
  assign new_n9324_ = ~new_n9320_ & new_n9323_;
  assign new_n9325_ = new_n4464_ & new_n8667_;
  assign new_n9326_ = new_n4464_ & new_n8670_;
  assign new_n9327_ = ~new_n9325_ & ~new_n9326_;
  assign new_n9328_ = new_n9324_ & new_n9327_;
  assign new_n9329_ = new_n9319_ & new_n9328_;
  assign new_n9330_ = new_n9308_ & new_n9329_;
  assign new_n9331_ = new_n9285_ & new_n9330_;
  assign new_n9332_ = new_n4464_ & new_n8681_;
  assign new_n9333_ = new_n4464_ & new_n8665_;
  assign new_n9334_ = new_n4464_ & new_n8678_;
  assign new_n9335_ = ~new_n9333_ & ~new_n9334_;
  assign new_n9336_ = ~new_n9332_ & new_n9335_;
  assign new_n9337_ = new_n4464_ & new_n8694_;
  assign new_n9338_ = new_n4464_ & new_n8675_;
  assign new_n9339_ = new_n4464_ & new_n8692_;
  assign new_n9340_ = ~new_n9338_ & ~new_n9339_;
  assign new_n9341_ = ~new_n9337_ & new_n9340_;
  assign new_n9342_ = new_n9336_ & new_n9341_;
  assign new_n9343_ = new_n4464_ & new_n8701_;
  assign new_n9344_ = new_n4464_ & new_n8689_;
  assign new_n9345_ = new_n4464_ & new_n8699_;
  assign new_n9346_ = ~new_n9344_ & ~new_n9345_;
  assign new_n9347_ = ~new_n9343_ & new_n9346_;
  assign new_n9348_ = new_n4471_ & new_n8630_;
  assign new_n9349_ = new_n4471_ & new_n8617_;
  assign new_n9350_ = new_n4471_ & new_n8628_;
  assign new_n9351_ = ~new_n9349_ & ~new_n9350_;
  assign new_n9352_ = ~new_n9348_ & new_n9351_;
  assign new_n9353_ = new_n9347_ & new_n9352_;
  assign new_n9354_ = new_n9342_ & new_n9353_;
  assign new_n9355_ = new_n4471_ & new_n8639_;
  assign new_n9356_ = new_n4471_ & new_n8625_;
  assign new_n9357_ = new_n4471_ & new_n8637_;
  assign new_n9358_ = ~new_n9356_ & ~new_n9357_;
  assign new_n9359_ = ~new_n9355_ & new_n9358_;
  assign new_n9360_ = new_n4471_ & new_n8650_;
  assign new_n9361_ = new_n4471_ & new_n8635_;
  assign new_n9362_ = new_n4471_ & new_n8648_;
  assign new_n9363_ = ~new_n9361_ & ~new_n9362_;
  assign new_n9364_ = ~new_n9360_ & new_n9363_;
  assign new_n9365_ = new_n9359_ & new_n9364_;
  assign new_n9366_ = new_n4471_ & new_n8659_;
  assign new_n9367_ = new_n4471_ & new_n8646_;
  assign new_n9368_ = new_n4471_ & new_n8657_;
  assign new_n9369_ = ~new_n9367_ & ~new_n9368_;
  assign new_n9370_ = ~new_n9366_ & new_n9369_;
  assign new_n9371_ = new_n4471_ & new_n8655_;
  assign new_n9372_ = new_n4471_ & new_n8667_;
  assign new_n9373_ = ~new_n9371_ & ~new_n9372_;
  assign new_n9374_ = new_n9370_ & new_n9373_;
  assign new_n9375_ = new_n9365_ & new_n9374_;
  assign new_n9376_ = new_n9354_ & new_n9375_;
  assign new_n9377_ = new_n4471_ & new_n8678_;
  assign new_n9378_ = new_n4471_ & new_n8670_;
  assign new_n9379_ = new_n4471_ & new_n8665_;
  assign new_n9380_ = ~new_n9378_ & ~new_n9379_;
  assign new_n9381_ = ~new_n9377_ & new_n9380_;
  assign new_n9382_ = new_n4471_ & new_n8692_;
  assign new_n9383_ = new_n4471_ & new_n8681_;
  assign new_n9384_ = new_n4471_ & new_n8675_;
  assign new_n9385_ = ~new_n9383_ & ~new_n9384_;
  assign new_n9386_ = ~new_n9382_ & new_n9385_;
  assign new_n9387_ = new_n9381_ & new_n9386_;
  assign new_n9388_ = new_n4471_ & new_n8699_;
  assign new_n9389_ = new_n4471_ & new_n8694_;
  assign new_n9390_ = new_n4471_ & new_n8689_;
  assign new_n9391_ = ~new_n9389_ & ~new_n9390_;
  assign new_n9392_ = ~new_n9388_ & new_n9391_;
  assign new_n9393_ = new_n4480_ & new_n8853_;
  assign new_n9394_ = new_n4471_ & new_n8701_;
  assign new_n9395_ = new_n4480_ & new_n8845_;
  assign new_n9396_ = ~new_n9394_ & ~new_n9395_;
  assign new_n9397_ = ~new_n9393_ & new_n9396_;
  assign new_n9398_ = new_n9392_ & new_n9397_;
  assign new_n9399_ = new_n9387_ & new_n9398_;
  assign new_n9400_ = new_n4480_ & new_n8864_;
  assign new_n9401_ = new_n4480_ & new_n8855_;
  assign new_n9402_ = new_n4480_ & new_n8851_;
  assign new_n9403_ = ~new_n9401_ & ~new_n9402_;
  assign new_n9404_ = ~new_n9400_ & new_n9403_;
  assign new_n9405_ = new_n4480_ & new_n8872_;
  assign new_n9406_ = new_n4480_ & new_n8866_;
  assign new_n9407_ = new_n4480_ & new_n8862_;
  assign new_n9408_ = ~new_n9406_ & ~new_n9407_;
  assign new_n9409_ = ~new_n9405_ & new_n9408_;
  assign new_n9410_ = new_n9404_ & new_n9409_;
  assign new_n9411_ = new_n4480_ & new_n8882_;
  assign new_n9412_ = new_n4480_ & new_n8874_;
  assign new_n9413_ = new_n4480_ & new_n8870_;
  assign new_n9414_ = ~new_n9412_ & ~new_n9413_;
  assign new_n9415_ = ~new_n9411_ & new_n9414_;
  assign new_n9416_ = new_n4480_ & new_n8884_;
  assign new_n9417_ = new_n4480_ & new_n8880_;
  assign new_n9418_ = ~new_n9416_ & ~new_n9417_;
  assign new_n9419_ = new_n9415_ & new_n9418_;
  assign new_n9420_ = new_n9410_ & new_n9419_;
  assign new_n9421_ = new_n9399_ & new_n9420_;
  assign new_n9422_ = new_n9376_ & new_n9421_;
  assign new_n9423_ = new_n9331_ & new_n9422_;
  assign new_n9424_ = new_n9240_ & new_n9423_;
  assign new_n9425_ = new_n4480_ & new_n8898_;
  assign new_n9426_ = new_n4480_ & new_n8888_;
  assign new_n9427_ = new_n4480_ & new_n8890_;
  assign new_n9428_ = ~new_n9426_ & ~new_n9427_;
  assign new_n9429_ = ~new_n9425_ & new_n9428_;
  assign new_n9430_ = new_n4480_ & new_n8907_;
  assign new_n9431_ = new_n4480_ & new_n8900_;
  assign new_n9432_ = new_n4480_ & new_n8896_;
  assign new_n9433_ = ~new_n9431_ & ~new_n9432_;
  assign new_n9434_ = ~new_n9430_ & new_n9433_;
  assign new_n9435_ = new_n9429_ & new_n9434_;
  assign new_n9436_ = new_n4480_ & new_n8916_;
  assign new_n9437_ = new_n4480_ & new_n8909_;
  assign new_n9438_ = new_n4480_ & new_n8905_;
  assign new_n9439_ = ~new_n9437_ & ~new_n9438_;
  assign new_n9440_ = ~new_n9436_ & new_n9439_;
  assign new_n9441_ = new_n4480_ & new_n8925_;
  assign new_n9442_ = new_n4480_ & new_n8918_;
  assign new_n9443_ = new_n4480_ & new_n8914_;
  assign new_n9444_ = ~new_n9442_ & ~new_n9443_;
  assign new_n9445_ = ~new_n9441_ & new_n9444_;
  assign new_n9446_ = new_n9440_ & new_n9445_;
  assign new_n9447_ = new_n9435_ & new_n9446_;
  assign new_n9448_ = new_n4480_ & new_n8936_;
  assign new_n9449_ = new_n4480_ & new_n8927_;
  assign new_n9450_ = new_n4480_ & new_n8923_;
  assign new_n9451_ = ~new_n9449_ & ~new_n9450_;
  assign new_n9452_ = ~new_n9448_ & new_n9451_;
  assign new_n9453_ = new_n4480_ & new_n8943_;
  assign new_n9454_ = new_n4480_ & new_n8938_;
  assign new_n9455_ = new_n4480_ & new_n8934_;
  assign new_n9456_ = ~new_n9454_ & ~new_n9455_;
  assign new_n9457_ = ~new_n9453_ & new_n9456_;
  assign new_n9458_ = new_n9452_ & new_n9457_;
  assign new_n9459_ = new_n4535_ & new_n8628_;
  assign new_n9460_ = new_n4480_ & new_n8945_;
  assign new_n9461_ = new_n4535_ & new_n8617_;
  assign new_n9462_ = ~new_n9460_ & ~new_n9461_;
  assign new_n9463_ = ~new_n9459_ & new_n9462_;
  assign new_n9464_ = new_n4535_ & new_n8630_;
  assign new_n9465_ = new_n4535_ & new_n8625_;
  assign new_n9466_ = ~new_n9464_ & ~new_n9465_;
  assign new_n9467_ = new_n9463_ & new_n9466_;
  assign new_n9468_ = new_n9458_ & new_n9467_;
  assign new_n9469_ = new_n9447_ & new_n9468_;
  assign new_n9470_ = new_n4535_ & new_n8635_;
  assign new_n9471_ = new_n4535_ & new_n8637_;
  assign new_n9472_ = new_n4535_ & new_n8639_;
  assign new_n9473_ = ~new_n9471_ & ~new_n9472_;
  assign new_n9474_ = ~new_n9470_ & new_n9473_;
  assign new_n9475_ = new_n4535_ & new_n8646_;
  assign new_n9476_ = new_n4535_ & new_n8648_;
  assign new_n9477_ = new_n4535_ & new_n8650_;
  assign new_n9478_ = ~new_n9476_ & ~new_n9477_;
  assign new_n9479_ = ~new_n9475_ & new_n9478_;
  assign new_n9480_ = new_n9474_ & new_n9479_;
  assign new_n9481_ = new_n4535_ & new_n8655_;
  assign new_n9482_ = new_n4535_ & new_n8657_;
  assign new_n9483_ = new_n4535_ & new_n8659_;
  assign new_n9484_ = ~new_n9482_ & ~new_n9483_;
  assign new_n9485_ = ~new_n9481_ & new_n9484_;
  assign new_n9486_ = new_n4535_ & new_n8665_;
  assign new_n9487_ = new_n4535_ & new_n8667_;
  assign new_n9488_ = new_n4535_ & new_n8670_;
  assign new_n9489_ = ~new_n9487_ & ~new_n9488_;
  assign new_n9490_ = ~new_n9486_ & new_n9489_;
  assign new_n9491_ = new_n9485_ & new_n9490_;
  assign new_n9492_ = new_n9480_ & new_n9491_;
  assign new_n9493_ = new_n4535_ & new_n8675_;
  assign new_n9494_ = new_n4535_ & new_n8678_;
  assign new_n9495_ = new_n4535_ & new_n8681_;
  assign new_n9496_ = ~new_n9494_ & ~new_n9495_;
  assign new_n9497_ = ~new_n9493_ & new_n9496_;
  assign new_n9498_ = new_n4535_ & new_n8689_;
  assign new_n9499_ = new_n4535_ & new_n8692_;
  assign new_n9500_ = new_n4535_ & new_n8694_;
  assign new_n9501_ = ~new_n9499_ & ~new_n9500_;
  assign new_n9502_ = ~new_n9498_ & new_n9501_;
  assign new_n9503_ = new_n9497_ & new_n9502_;
  assign new_n9504_ = new_n4543_ & new_n8617_;
  assign new_n9505_ = new_n4535_ & new_n8699_;
  assign new_n9506_ = new_n4535_ & new_n8701_;
  assign new_n9507_ = ~new_n9505_ & ~new_n9506_;
  assign new_n9508_ = ~new_n9504_ & new_n9507_;
  assign new_n9509_ = new_n4543_ & new_n8628_;
  assign new_n9510_ = new_n4543_ & new_n8630_;
  assign new_n9511_ = ~new_n9509_ & ~new_n9510_;
  assign new_n9512_ = new_n9508_ & new_n9511_;
  assign new_n9513_ = new_n9503_ & new_n9512_;
  assign new_n9514_ = new_n9492_ & new_n9513_;
  assign new_n9515_ = new_n9469_ & new_n9514_;
  assign new_n9516_ = new_n4543_ & new_n8639_;
  assign new_n9517_ = new_n4543_ & new_n8625_;
  assign new_n9518_ = new_n4543_ & new_n8637_;
  assign new_n9519_ = ~new_n9517_ & ~new_n9518_;
  assign new_n9520_ = ~new_n9516_ & new_n9519_;
  assign new_n9521_ = new_n4543_ & new_n8650_;
  assign new_n9522_ = new_n4543_ & new_n8635_;
  assign new_n9523_ = new_n4543_ & new_n8648_;
  assign new_n9524_ = ~new_n9522_ & ~new_n9523_;
  assign new_n9525_ = ~new_n9521_ & new_n9524_;
  assign new_n9526_ = new_n9520_ & new_n9525_;
  assign new_n9527_ = new_n4543_ & new_n8659_;
  assign new_n9528_ = new_n4543_ & new_n8646_;
  assign new_n9529_ = new_n4543_ & new_n8657_;
  assign new_n9530_ = ~new_n9528_ & ~new_n9529_;
  assign new_n9531_ = ~new_n9527_ & new_n9530_;
  assign new_n9532_ = new_n4543_ & new_n8670_;
  assign new_n9533_ = new_n4543_ & new_n8655_;
  assign new_n9534_ = new_n4543_ & new_n8667_;
  assign new_n9535_ = ~new_n9533_ & ~new_n9534_;
  assign new_n9536_ = ~new_n9532_ & new_n9535_;
  assign new_n9537_ = new_n9531_ & new_n9536_;
  assign new_n9538_ = new_n9526_ & new_n9537_;
  assign new_n9539_ = new_n4543_ & new_n8681_;
  assign new_n9540_ = new_n4543_ & new_n8665_;
  assign new_n9541_ = new_n4543_ & new_n8678_;
  assign new_n9542_ = ~new_n9540_ & ~new_n9541_;
  assign new_n9543_ = ~new_n9539_ & new_n9542_;
  assign new_n9544_ = new_n4543_ & new_n8694_;
  assign new_n9545_ = new_n4543_ & new_n8675_;
  assign new_n9546_ = new_n4543_ & new_n8692_;
  assign new_n9547_ = ~new_n9545_ & ~new_n9546_;
  assign new_n9548_ = ~new_n9544_ & new_n9547_;
  assign new_n9549_ = new_n9543_ & new_n9548_;
  assign new_n9550_ = new_n4543_ & new_n8701_;
  assign new_n9551_ = new_n4543_ & new_n8689_;
  assign new_n9552_ = new_n4543_ & new_n8699_;
  assign new_n9553_ = ~new_n9551_ & ~new_n9552_;
  assign new_n9554_ = ~new_n9550_ & new_n9553_;
  assign new_n9555_ = new_n4556_ & new_n8617_;
  assign new_n9556_ = new_n4556_ & new_n8628_;
  assign new_n9557_ = ~new_n9555_ & ~new_n9556_;
  assign new_n9558_ = new_n9554_ & new_n9557_;
  assign new_n9559_ = new_n9549_ & new_n9558_;
  assign new_n9560_ = new_n9538_ & new_n9559_;
  assign new_n9561_ = new_n4556_ & new_n8637_;
  assign new_n9562_ = new_n4556_ & new_n8630_;
  assign new_n9563_ = new_n4556_ & new_n8625_;
  assign new_n9564_ = ~new_n9562_ & ~new_n9563_;
  assign new_n9565_ = ~new_n9561_ & new_n9564_;
  assign new_n9566_ = new_n4556_ & new_n8648_;
  assign new_n9567_ = new_n4556_ & new_n8639_;
  assign new_n9568_ = new_n4556_ & new_n8635_;
  assign new_n9569_ = ~new_n9567_ & ~new_n9568_;
  assign new_n9570_ = ~new_n9566_ & new_n9569_;
  assign new_n9571_ = new_n9565_ & new_n9570_;
  assign new_n9572_ = new_n4556_ & new_n8657_;
  assign new_n9573_ = new_n4556_ & new_n8650_;
  assign new_n9574_ = new_n4556_ & new_n8646_;
  assign new_n9575_ = ~new_n9573_ & ~new_n9574_;
  assign new_n9576_ = ~new_n9572_ & new_n9575_;
  assign new_n9577_ = new_n4556_ & new_n8667_;
  assign new_n9578_ = new_n4556_ & new_n8659_;
  assign new_n9579_ = new_n4556_ & new_n8655_;
  assign new_n9580_ = ~new_n9578_ & ~new_n9579_;
  assign new_n9581_ = ~new_n9577_ & new_n9580_;
  assign new_n9582_ = new_n9576_ & new_n9581_;
  assign new_n9583_ = new_n9571_ & new_n9582_;
  assign new_n9584_ = new_n4556_ & new_n8678_;
  assign new_n9585_ = new_n4556_ & new_n8670_;
  assign new_n9586_ = new_n4556_ & new_n8665_;
  assign new_n9587_ = ~new_n9585_ & ~new_n9586_;
  assign new_n9588_ = ~new_n9584_ & new_n9587_;
  assign new_n9589_ = new_n4556_ & new_n8692_;
  assign new_n9590_ = new_n4556_ & new_n8681_;
  assign new_n9591_ = new_n4556_ & new_n8675_;
  assign new_n9592_ = ~new_n9590_ & ~new_n9591_;
  assign new_n9593_ = ~new_n9589_ & new_n9592_;
  assign new_n9594_ = new_n9588_ & new_n9593_;
  assign new_n9595_ = new_n4556_ & new_n8699_;
  assign new_n9596_ = new_n4556_ & new_n8694_;
  assign new_n9597_ = new_n4556_ & new_n8689_;
  assign new_n9598_ = ~new_n9596_ & ~new_n9597_;
  assign new_n9599_ = ~new_n9595_ & new_n9598_;
  assign new_n9600_ = new_n4556_ & new_n8701_;
  assign new_n9601_ = new_n4563_ & new_n8617_;
  assign new_n9602_ = ~new_n9600_ & ~new_n9601_;
  assign new_n9603_ = new_n9599_ & new_n9602_;
  assign new_n9604_ = new_n9594_ & new_n9603_;
  assign new_n9605_ = new_n9583_ & new_n9604_;
  assign new_n9606_ = new_n9560_ & new_n9605_;
  assign new_n9607_ = new_n9515_ & new_n9606_;
  assign new_n9608_ = new_n4563_ & new_n8625_;
  assign new_n9609_ = new_n4563_ & new_n8628_;
  assign new_n9610_ = new_n4563_ & new_n8630_;
  assign new_n9611_ = ~new_n9609_ & ~new_n9610_;
  assign new_n9612_ = ~new_n9608_ & new_n9611_;
  assign new_n9613_ = new_n4563_ & new_n8635_;
  assign new_n9614_ = new_n4563_ & new_n8637_;
  assign new_n9615_ = new_n4563_ & new_n8639_;
  assign new_n9616_ = ~new_n9614_ & ~new_n9615_;
  assign new_n9617_ = ~new_n9613_ & new_n9616_;
  assign new_n9618_ = new_n9612_ & new_n9617_;
  assign new_n9619_ = new_n4563_ & new_n8646_;
  assign new_n9620_ = new_n4563_ & new_n8648_;
  assign new_n9621_ = new_n4563_ & new_n8650_;
  assign new_n9622_ = ~new_n9620_ & ~new_n9621_;
  assign new_n9623_ = ~new_n9619_ & new_n9622_;
  assign new_n9624_ = new_n4563_ & new_n8655_;
  assign new_n9625_ = new_n4563_ & new_n8657_;
  assign new_n9626_ = new_n4563_ & new_n8659_;
  assign new_n9627_ = ~new_n9625_ & ~new_n9626_;
  assign new_n9628_ = ~new_n9624_ & new_n9627_;
  assign new_n9629_ = new_n9623_ & new_n9628_;
  assign new_n9630_ = new_n9618_ & new_n9629_;
  assign new_n9631_ = new_n4563_ & new_n8665_;
  assign new_n9632_ = new_n4563_ & new_n8667_;
  assign new_n9633_ = new_n4563_ & new_n8670_;
  assign new_n9634_ = ~new_n9632_ & ~new_n9633_;
  assign new_n9635_ = ~new_n9631_ & new_n9634_;
  assign new_n9636_ = new_n4563_ & new_n8675_;
  assign new_n9637_ = new_n4563_ & new_n8678_;
  assign new_n9638_ = new_n4563_ & new_n8681_;
  assign new_n9639_ = ~new_n9637_ & ~new_n9638_;
  assign new_n9640_ = ~new_n9636_ & new_n9639_;
  assign new_n9641_ = new_n9635_ & new_n9640_;
  assign new_n9642_ = new_n4563_ & new_n8689_;
  assign new_n9643_ = new_n4563_ & new_n8692_;
  assign new_n9644_ = new_n4563_ & new_n8694_;
  assign new_n9645_ = ~new_n9643_ & ~new_n9644_;
  assign new_n9646_ = ~new_n9642_ & new_n9645_;
  assign new_n9647_ = new_n4563_ & new_n8699_;
  assign new_n9648_ = new_n4563_ & new_n8701_;
  assign new_n9649_ = ~new_n9647_ & ~new_n9648_;
  assign new_n9650_ = new_n9646_ & new_n9649_;
  assign new_n9651_ = new_n9641_ & new_n9650_;
  assign new_n9652_ = new_n9630_ & new_n9651_;
  assign new_n9653_ = new_n4571_ & new_n8855_;
  assign new_n9654_ = new_n4571_ & new_n8845_;
  assign new_n9655_ = new_n4571_ & new_n8853_;
  assign new_n9656_ = ~new_n9654_ & ~new_n9655_;
  assign new_n9657_ = ~new_n9653_ & new_n9656_;
  assign new_n9658_ = new_n4571_ & new_n8866_;
  assign new_n9659_ = new_n4571_ & new_n8851_;
  assign new_n9660_ = new_n4571_ & new_n8864_;
  assign new_n9661_ = ~new_n9659_ & ~new_n9660_;
  assign new_n9662_ = ~new_n9658_ & new_n9661_;
  assign new_n9663_ = new_n9657_ & new_n9662_;
  assign new_n9664_ = new_n4571_ & new_n8874_;
  assign new_n9665_ = new_n4571_ & new_n8862_;
  assign new_n9666_ = new_n4571_ & new_n8872_;
  assign new_n9667_ = ~new_n9665_ & ~new_n9666_;
  assign new_n9668_ = ~new_n9664_ & new_n9667_;
  assign new_n9669_ = new_n4571_ & new_n8884_;
  assign new_n9670_ = new_n4571_ & new_n8870_;
  assign new_n9671_ = new_n4571_ & new_n8882_;
  assign new_n9672_ = ~new_n9670_ & ~new_n9671_;
  assign new_n9673_ = ~new_n9669_ & new_n9672_;
  assign new_n9674_ = new_n9668_ & new_n9673_;
  assign new_n9675_ = new_n9663_ & new_n9674_;
  assign new_n9676_ = new_n4571_ & new_n8890_;
  assign new_n9677_ = new_n4571_ & new_n8880_;
  assign new_n9678_ = new_n4571_ & new_n8888_;
  assign new_n9679_ = ~new_n9677_ & ~new_n9678_;
  assign new_n9680_ = ~new_n9676_ & new_n9679_;
  assign new_n9681_ = new_n4571_ & new_n8896_;
  assign new_n9682_ = new_n4571_ & new_n8898_;
  assign new_n9683_ = new_n4571_ & new_n8900_;
  assign new_n9684_ = ~new_n9682_ & ~new_n9683_;
  assign new_n9685_ = ~new_n9681_ & new_n9684_;
  assign new_n9686_ = new_n9680_ & new_n9685_;
  assign new_n9687_ = new_n4571_ & new_n8905_;
  assign new_n9688_ = new_n4571_ & new_n8907_;
  assign new_n9689_ = new_n4571_ & new_n8909_;
  assign new_n9690_ = ~new_n9688_ & ~new_n9689_;
  assign new_n9691_ = ~new_n9687_ & new_n9690_;
  assign new_n9692_ = new_n4571_ & new_n8916_;
  assign new_n9693_ = new_n4571_ & new_n8918_;
  assign new_n9694_ = ~new_n9692_ & ~new_n9693_;
  assign new_n9695_ = new_n9691_ & new_n9694_;
  assign new_n9696_ = new_n9686_ & new_n9695_;
  assign new_n9697_ = new_n9675_ & new_n9696_;
  assign new_n9698_ = new_n9652_ & new_n9697_;
  assign new_n9699_ = new_n4571_ & new_n8927_;
  assign new_n9700_ = new_n4571_ & new_n8914_;
  assign new_n9701_ = new_n4571_ & new_n8925_;
  assign new_n9702_ = ~new_n9700_ & ~new_n9701_;
  assign new_n9703_ = ~new_n9699_ & new_n9702_;
  assign new_n9704_ = new_n4571_ & new_n8938_;
  assign new_n9705_ = new_n4571_ & new_n8923_;
  assign new_n9706_ = new_n4571_ & new_n8936_;
  assign new_n9707_ = ~new_n9705_ & ~new_n9706_;
  assign new_n9708_ = ~new_n9704_ & new_n9707_;
  assign new_n9709_ = new_n9703_ & new_n9708_;
  assign new_n9710_ = new_n4571_ & new_n8945_;
  assign new_n9711_ = new_n4571_ & new_n8934_;
  assign new_n9712_ = new_n4571_ & new_n8943_;
  assign new_n9713_ = ~new_n9711_ & ~new_n9712_;
  assign new_n9714_ = ~new_n9710_ & new_n9713_;
  assign new_n9715_ = ~A233 & new_n139_;
  assign new_n9716_ = new_n947_ & new_n9715_;
  assign new_n9717_ = new_n4627_ & new_n9716_;
  assign new_n9718_ = new_n950_ & new_n9715_;
  assign new_n9719_ = new_n4627_ & new_n9718_;
  assign new_n9720_ = new_n953_ & new_n9715_;
  assign new_n9721_ = new_n4627_ & new_n9720_;
  assign new_n9722_ = ~new_n9719_ & ~new_n9721_;
  assign new_n9723_ = ~new_n9717_ & new_n9722_;
  assign new_n9724_ = new_n9714_ & new_n9723_;
  assign new_n9725_ = new_n9709_ & new_n9724_;
  assign new_n9726_ = ~A233 & new_n155_;
  assign new_n9727_ = new_n960_ & new_n9726_;
  assign new_n9728_ = new_n4627_ & new_n9727_;
  assign new_n9729_ = new_n963_ & new_n9715_;
  assign new_n9730_ = new_n4627_ & new_n9729_;
  assign new_n9731_ = new_n966_ & new_n9726_;
  assign new_n9732_ = new_n4627_ & new_n9731_;
  assign new_n9733_ = ~new_n9730_ & ~new_n9732_;
  assign new_n9734_ = ~new_n9728_ & new_n9733_;
  assign new_n9735_ = new_n971_ & new_n9726_;
  assign new_n9736_ = new_n4627_ & new_n9735_;
  assign new_n9737_ = new_n974_ & new_n9726_;
  assign new_n9738_ = new_n4627_ & new_n9737_;
  assign new_n9739_ = new_n977_ & new_n9726_;
  assign new_n9740_ = new_n4627_ & new_n9739_;
  assign new_n9741_ = ~new_n9738_ & ~new_n9740_;
  assign new_n9742_ = ~new_n9736_ & new_n9741_;
  assign new_n9743_ = new_n9734_ & new_n9742_;
  assign new_n9744_ = new_n983_ & new_n9726_;
  assign new_n9745_ = new_n4627_ & new_n9744_;
  assign new_n9746_ = new_n986_ & new_n9726_;
  assign new_n9747_ = new_n4627_ & new_n9746_;
  assign new_n9748_ = new_n989_ & new_n9726_;
  assign new_n9749_ = new_n4627_ & new_n9748_;
  assign new_n9750_ = ~new_n9747_ & ~new_n9749_;
  assign new_n9751_ = ~new_n9745_ & new_n9750_;
  assign new_n9752_ = ~A233 & new_n186_;
  assign new_n9753_ = new_n966_ & new_n9752_;
  assign new_n9754_ = new_n4627_ & new_n9753_;
  assign new_n9755_ = new_n960_ & new_n9752_;
  assign new_n9756_ = new_n4627_ & new_n9755_;
  assign new_n9757_ = ~new_n9754_ & ~new_n9756_;
  assign new_n9758_ = new_n9751_ & new_n9757_;
  assign new_n9759_ = new_n9743_ & new_n9758_;
  assign new_n9760_ = new_n9725_ & new_n9759_;
  assign new_n9761_ = new_n971_ & new_n9752_;
  assign new_n9762_ = new_n4627_ & new_n9761_;
  assign new_n9763_ = new_n974_ & new_n9752_;
  assign new_n9764_ = new_n4627_ & new_n9763_;
  assign new_n9765_ = new_n977_ & new_n9752_;
  assign new_n9766_ = new_n4627_ & new_n9765_;
  assign new_n9767_ = ~new_n9764_ & ~new_n9766_;
  assign new_n9768_ = ~new_n9762_ & new_n9767_;
  assign new_n9769_ = new_n983_ & new_n9752_;
  assign new_n9770_ = new_n4627_ & new_n9769_;
  assign new_n9771_ = new_n986_ & new_n9752_;
  assign new_n9772_ = new_n4627_ & new_n9771_;
  assign new_n9773_ = new_n989_ & new_n9752_;
  assign new_n9774_ = new_n4627_ & new_n9773_;
  assign new_n9775_ = ~new_n9772_ & ~new_n9774_;
  assign new_n9776_ = ~new_n9770_ & new_n9775_;
  assign new_n9777_ = new_n9768_ & new_n9776_;
  assign new_n9778_ = ~A233 & new_n209_;
  assign new_n9779_ = new_n947_ & new_n9778_;
  assign new_n9780_ = new_n4627_ & new_n9779_;
  assign new_n9781_ = new_n950_ & new_n9778_;
  assign new_n9782_ = new_n4627_ & new_n9781_;
  assign new_n9783_ = new_n953_ & new_n9778_;
  assign new_n9784_ = new_n4627_ & new_n9783_;
  assign new_n9785_ = ~new_n9782_ & ~new_n9784_;
  assign new_n9786_ = ~new_n9780_ & new_n9785_;
  assign new_n9787_ = ~A233 & new_n218_;
  assign new_n9788_ = new_n953_ & new_n9787_;
  assign new_n9789_ = new_n4627_ & new_n9788_;
  assign new_n9790_ = new_n963_ & new_n9778_;
  assign new_n9791_ = new_n4627_ & new_n9790_;
  assign new_n9792_ = new_n950_ & new_n9787_;
  assign new_n9793_ = new_n4627_ & new_n9792_;
  assign new_n9794_ = ~new_n9791_ & ~new_n9793_;
  assign new_n9795_ = ~new_n9789_ & new_n9794_;
  assign new_n9796_ = new_n9786_ & new_n9795_;
  assign new_n9797_ = new_n9777_ & new_n9796_;
  assign new_n9798_ = ~A233 & new_n236_;
  assign new_n9799_ = new_n950_ & new_n9798_;
  assign new_n9800_ = new_n4627_ & new_n9799_;
  assign new_n9801_ = new_n947_ & new_n9787_;
  assign new_n9802_ = new_n4627_ & new_n9801_;
  assign new_n9803_ = new_n963_ & new_n9787_;
  assign new_n9804_ = new_n4627_ & new_n9803_;
  assign new_n9805_ = ~new_n9802_ & ~new_n9804_;
  assign new_n9806_ = ~new_n9800_ & new_n9805_;
  assign new_n9807_ = new_n963_ & new_n9798_;
  assign new_n9808_ = new_n4627_ & new_n9807_;
  assign new_n9809_ = new_n953_ & new_n9798_;
  assign new_n9810_ = new_n4627_ & new_n9809_;
  assign new_n9811_ = new_n947_ & new_n9798_;
  assign new_n9812_ = new_n4627_ & new_n9811_;
  assign new_n9813_ = ~new_n9810_ & ~new_n9812_;
  assign new_n9814_ = ~new_n9808_ & new_n9813_;
  assign new_n9815_ = new_n9806_ & new_n9814_;
  assign new_n9816_ = A233 & new_n139_;
  assign new_n9817_ = new_n947_ & new_n9816_;
  assign new_n9818_ = new_n4714_ & new_n9817_;
  assign new_n9819_ = new_n950_ & new_n9816_;
  assign new_n9820_ = new_n4714_ & new_n9819_;
  assign new_n9821_ = new_n953_ & new_n9816_;
  assign new_n9822_ = new_n4714_ & new_n9821_;
  assign new_n9823_ = ~new_n9820_ & ~new_n9822_;
  assign new_n9824_ = ~new_n9818_ & new_n9823_;
  assign new_n9825_ = new_n963_ & new_n9816_;
  assign new_n9826_ = new_n4714_ & new_n9825_;
  assign new_n9827_ = A233 & new_n155_;
  assign new_n9828_ = new_n966_ & new_n9827_;
  assign new_n9829_ = new_n4714_ & new_n9828_;
  assign new_n9830_ = ~new_n9826_ & ~new_n9829_;
  assign new_n9831_ = new_n9824_ & new_n9830_;
  assign new_n9832_ = new_n9815_ & new_n9831_;
  assign new_n9833_ = new_n9797_ & new_n9832_;
  assign new_n9834_ = new_n9760_ & new_n9833_;
  assign new_n9835_ = new_n9698_ & new_n9834_;
  assign new_n9836_ = new_n9607_ & new_n9835_;
  assign new_n9837_ = new_n9424_ & new_n9836_;
  assign new_n9838_ = new_n9055_ & new_n9837_;
  assign new_n9839_ = new_n8237_ & new_n9838_;
  assign new_n9840_ = new_n977_ & new_n9827_;
  assign new_n9841_ = new_n4714_ & new_n9840_;
  assign new_n9842_ = new_n960_ & new_n9827_;
  assign new_n9843_ = new_n4714_ & new_n9842_;
  assign new_n9844_ = new_n974_ & new_n9827_;
  assign new_n9845_ = new_n4714_ & new_n9844_;
  assign new_n9846_ = ~new_n9843_ & ~new_n9845_;
  assign new_n9847_ = ~new_n9841_ & new_n9846_;
  assign new_n9848_ = new_n989_ & new_n9827_;
  assign new_n9849_ = new_n4714_ & new_n9848_;
  assign new_n9850_ = new_n971_ & new_n9827_;
  assign new_n9851_ = new_n4714_ & new_n9850_;
  assign new_n9852_ = new_n986_ & new_n9827_;
  assign new_n9853_ = new_n4714_ & new_n9852_;
  assign new_n9854_ = ~new_n9851_ & ~new_n9853_;
  assign new_n9855_ = ~new_n9849_ & new_n9854_;
  assign new_n9856_ = new_n9847_ & new_n9855_;
  assign new_n9857_ = A233 & new_n186_;
  assign new_n9858_ = new_n960_ & new_n9857_;
  assign new_n9859_ = new_n4714_ & new_n9858_;
  assign new_n9860_ = new_n983_ & new_n9827_;
  assign new_n9861_ = new_n4714_ & new_n9860_;
  assign new_n9862_ = new_n966_ & new_n9857_;
  assign new_n9863_ = new_n4714_ & new_n9862_;
  assign new_n9864_ = ~new_n9861_ & ~new_n9863_;
  assign new_n9865_ = ~new_n9859_ & new_n9864_;
  assign new_n9866_ = new_n971_ & new_n9857_;
  assign new_n9867_ = new_n4714_ & new_n9866_;
  assign new_n9868_ = new_n974_ & new_n9857_;
  assign new_n9869_ = new_n4714_ & new_n9868_;
  assign new_n9870_ = new_n977_ & new_n9857_;
  assign new_n9871_ = new_n4714_ & new_n9870_;
  assign new_n9872_ = ~new_n9869_ & ~new_n9871_;
  assign new_n9873_ = ~new_n9867_ & new_n9872_;
  assign new_n9874_ = new_n9865_ & new_n9873_;
  assign new_n9875_ = new_n9856_ & new_n9874_;
  assign new_n9876_ = new_n983_ & new_n9857_;
  assign new_n9877_ = new_n4714_ & new_n9876_;
  assign new_n9878_ = new_n986_ & new_n9857_;
  assign new_n9879_ = new_n4714_ & new_n9878_;
  assign new_n9880_ = new_n989_ & new_n9857_;
  assign new_n9881_ = new_n4714_ & new_n9880_;
  assign new_n9882_ = ~new_n9879_ & ~new_n9881_;
  assign new_n9883_ = ~new_n9877_ & new_n9882_;
  assign new_n9884_ = A233 & new_n209_;
  assign new_n9885_ = new_n947_ & new_n9884_;
  assign new_n9886_ = new_n4714_ & new_n9885_;
  assign new_n9887_ = new_n950_ & new_n9884_;
  assign new_n9888_ = new_n4714_ & new_n9887_;
  assign new_n9889_ = new_n953_ & new_n9884_;
  assign new_n9890_ = new_n4714_ & new_n9889_;
  assign new_n9891_ = ~new_n9888_ & ~new_n9890_;
  assign new_n9892_ = ~new_n9886_ & new_n9891_;
  assign new_n9893_ = new_n9883_ & new_n9892_;
  assign new_n9894_ = A233 & new_n218_;
  assign new_n9895_ = new_n953_ & new_n9894_;
  assign new_n9896_ = new_n4714_ & new_n9895_;
  assign new_n9897_ = new_n963_ & new_n9884_;
  assign new_n9898_ = new_n4714_ & new_n9897_;
  assign new_n9899_ = new_n950_ & new_n9894_;
  assign new_n9900_ = new_n4714_ & new_n9899_;
  assign new_n9901_ = ~new_n9898_ & ~new_n9900_;
  assign new_n9902_ = ~new_n9896_ & new_n9901_;
  assign new_n9903_ = A233 & new_n236_;
  assign new_n9904_ = new_n950_ & new_n9903_;
  assign new_n9905_ = new_n4714_ & new_n9904_;
  assign new_n9906_ = new_n947_ & new_n9894_;
  assign new_n9907_ = new_n4714_ & new_n9906_;
  assign new_n9908_ = new_n963_ & new_n9894_;
  assign new_n9909_ = new_n4714_ & new_n9908_;
  assign new_n9910_ = ~new_n9907_ & ~new_n9909_;
  assign new_n9911_ = ~new_n9905_ & new_n9910_;
  assign new_n9912_ = new_n9902_ & new_n9911_;
  assign new_n9913_ = new_n9893_ & new_n9912_;
  assign new_n9914_ = new_n9875_ & new_n9913_;
  assign new_n9915_ = new_n963_ & new_n9903_;
  assign new_n9916_ = new_n4714_ & new_n9915_;
  assign new_n9917_ = new_n953_ & new_n9903_;
  assign new_n9918_ = new_n4714_ & new_n9917_;
  assign new_n9919_ = new_n947_ & new_n9903_;
  assign new_n9920_ = new_n4714_ & new_n9919_;
  assign new_n9921_ = ~new_n9918_ & ~new_n9920_;
  assign new_n9922_ = ~new_n9916_ & new_n9921_;
  assign new_n9923_ = ~A236 & new_n139_;
  assign new_n9924_ = new_n947_ & new_n9923_;
  assign new_n9925_ = new_n4802_ & new_n9924_;
  assign new_n9926_ = new_n950_ & new_n9923_;
  assign new_n9927_ = new_n4802_ & new_n9926_;
  assign new_n9928_ = new_n953_ & new_n9923_;
  assign new_n9929_ = new_n4802_ & new_n9928_;
  assign new_n9930_ = ~new_n9927_ & ~new_n9929_;
  assign new_n9931_ = ~new_n9925_ & new_n9930_;
  assign new_n9932_ = new_n9922_ & new_n9931_;
  assign new_n9933_ = ~A236 & new_n155_;
  assign new_n9934_ = new_n960_ & new_n9933_;
  assign new_n9935_ = new_n4802_ & new_n9934_;
  assign new_n9936_ = new_n963_ & new_n9923_;
  assign new_n9937_ = new_n4802_ & new_n9936_;
  assign new_n9938_ = new_n966_ & new_n9933_;
  assign new_n9939_ = new_n4802_ & new_n9938_;
  assign new_n9940_ = ~new_n9937_ & ~new_n9939_;
  assign new_n9941_ = ~new_n9935_ & new_n9940_;
  assign new_n9942_ = new_n971_ & new_n9933_;
  assign new_n9943_ = new_n4802_ & new_n9942_;
  assign new_n9944_ = new_n974_ & new_n9933_;
  assign new_n9945_ = new_n4802_ & new_n9944_;
  assign new_n9946_ = new_n977_ & new_n9933_;
  assign new_n9947_ = new_n4802_ & new_n9946_;
  assign new_n9948_ = ~new_n9945_ & ~new_n9947_;
  assign new_n9949_ = ~new_n9943_ & new_n9948_;
  assign new_n9950_ = new_n9941_ & new_n9949_;
  assign new_n9951_ = new_n9932_ & new_n9950_;
  assign new_n9952_ = new_n983_ & new_n9933_;
  assign new_n9953_ = new_n4802_ & new_n9952_;
  assign new_n9954_ = new_n986_ & new_n9933_;
  assign new_n9955_ = new_n4802_ & new_n9954_;
  assign new_n9956_ = new_n989_ & new_n9933_;
  assign new_n9957_ = new_n4802_ & new_n9956_;
  assign new_n9958_ = ~new_n9955_ & ~new_n9957_;
  assign new_n9959_ = ~new_n9953_ & new_n9958_;
  assign new_n9960_ = ~A236 & new_n186_;
  assign new_n9961_ = new_n974_ & new_n9960_;
  assign new_n9962_ = new_n4802_ & new_n9961_;
  assign new_n9963_ = new_n966_ & new_n9960_;
  assign new_n9964_ = new_n4802_ & new_n9963_;
  assign new_n9965_ = new_n960_ & new_n9960_;
  assign new_n9966_ = new_n4802_ & new_n9965_;
  assign new_n9967_ = ~new_n9964_ & ~new_n9966_;
  assign new_n9968_ = ~new_n9962_ & new_n9967_;
  assign new_n9969_ = new_n9959_ & new_n9968_;
  assign new_n9970_ = new_n986_ & new_n9960_;
  assign new_n9971_ = new_n4802_ & new_n9970_;
  assign new_n9972_ = new_n977_ & new_n9960_;
  assign new_n9973_ = new_n4802_ & new_n9972_;
  assign new_n9974_ = new_n971_ & new_n9960_;
  assign new_n9975_ = new_n4802_ & new_n9974_;
  assign new_n9976_ = ~new_n9973_ & ~new_n9975_;
  assign new_n9977_ = ~new_n9971_ & new_n9976_;
  assign new_n9978_ = new_n989_ & new_n9960_;
  assign new_n9979_ = new_n4802_ & new_n9978_;
  assign new_n9980_ = new_n983_ & new_n9960_;
  assign new_n9981_ = new_n4802_ & new_n9980_;
  assign new_n9982_ = ~new_n9979_ & ~new_n9981_;
  assign new_n9983_ = new_n9977_ & new_n9982_;
  assign new_n9984_ = new_n9969_ & new_n9983_;
  assign new_n9985_ = new_n9951_ & new_n9984_;
  assign new_n9986_ = new_n9914_ & new_n9985_;
  assign new_n9987_ = ~A236 & new_n209_;
  assign new_n9988_ = new_n947_ & new_n9987_;
  assign new_n9989_ = new_n4802_ & new_n9988_;
  assign new_n9990_ = new_n950_ & new_n9987_;
  assign new_n9991_ = new_n4802_ & new_n9990_;
  assign new_n9992_ = new_n953_ & new_n9987_;
  assign new_n9993_ = new_n4802_ & new_n9992_;
  assign new_n9994_ = ~new_n9991_ & ~new_n9993_;
  assign new_n9995_ = ~new_n9989_ & new_n9994_;
  assign new_n9996_ = ~A236 & new_n218_;
  assign new_n9997_ = new_n953_ & new_n9996_;
  assign new_n9998_ = new_n4802_ & new_n9997_;
  assign new_n9999_ = new_n963_ & new_n9987_;
  assign new_n10000_ = new_n4802_ & new_n9999_;
  assign new_n10001_ = new_n950_ & new_n9996_;
  assign new_n10002_ = new_n4802_ & new_n10001_;
  assign new_n10003_ = ~new_n10000_ & ~new_n10002_;
  assign new_n10004_ = ~new_n9998_ & new_n10003_;
  assign new_n10005_ = new_n9995_ & new_n10004_;
  assign new_n10006_ = ~A236 & new_n236_;
  assign new_n10007_ = new_n950_ & new_n10006_;
  assign new_n10008_ = new_n4802_ & new_n10007_;
  assign new_n10009_ = new_n947_ & new_n9996_;
  assign new_n10010_ = new_n4802_ & new_n10009_;
  assign new_n10011_ = new_n963_ & new_n9996_;
  assign new_n10012_ = new_n4802_ & new_n10011_;
  assign new_n10013_ = ~new_n10010_ & ~new_n10012_;
  assign new_n10014_ = ~new_n10008_ & new_n10013_;
  assign new_n10015_ = new_n963_ & new_n10006_;
  assign new_n10016_ = new_n4802_ & new_n10015_;
  assign new_n10017_ = new_n953_ & new_n10006_;
  assign new_n10018_ = new_n4802_ & new_n10017_;
  assign new_n10019_ = new_n947_ & new_n10006_;
  assign new_n10020_ = new_n4802_ & new_n10019_;
  assign new_n10021_ = ~new_n10018_ & ~new_n10020_;
  assign new_n10022_ = ~new_n10016_ & new_n10021_;
  assign new_n10023_ = new_n10014_ & new_n10022_;
  assign new_n10024_ = new_n10005_ & new_n10023_;
  assign new_n10025_ = A235 & new_n139_;
  assign new_n10026_ = new_n947_ & new_n10025_;
  assign new_n10027_ = new_n4802_ & new_n10026_;
  assign new_n10028_ = new_n950_ & new_n10025_;
  assign new_n10029_ = new_n4802_ & new_n10028_;
  assign new_n10030_ = new_n953_ & new_n10025_;
  assign new_n10031_ = new_n4802_ & new_n10030_;
  assign new_n10032_ = ~new_n10029_ & ~new_n10031_;
  assign new_n10033_ = ~new_n10027_ & new_n10032_;
  assign new_n10034_ = A235 & new_n155_;
  assign new_n10035_ = new_n960_ & new_n10034_;
  assign new_n10036_ = new_n4802_ & new_n10035_;
  assign new_n10037_ = new_n963_ & new_n10025_;
  assign new_n10038_ = new_n4802_ & new_n10037_;
  assign new_n10039_ = new_n966_ & new_n10034_;
  assign new_n10040_ = new_n4802_ & new_n10039_;
  assign new_n10041_ = ~new_n10038_ & ~new_n10040_;
  assign new_n10042_ = ~new_n10036_ & new_n10041_;
  assign new_n10043_ = new_n10033_ & new_n10042_;
  assign new_n10044_ = new_n971_ & new_n10034_;
  assign new_n10045_ = new_n4802_ & new_n10044_;
  assign new_n10046_ = new_n974_ & new_n10034_;
  assign new_n10047_ = new_n4802_ & new_n10046_;
  assign new_n10048_ = new_n977_ & new_n10034_;
  assign new_n10049_ = new_n4802_ & new_n10048_;
  assign new_n10050_ = ~new_n10047_ & ~new_n10049_;
  assign new_n10051_ = ~new_n10045_ & new_n10050_;
  assign new_n10052_ = new_n986_ & new_n10034_;
  assign new_n10053_ = new_n4802_ & new_n10052_;
  assign new_n10054_ = new_n989_ & new_n10034_;
  assign new_n10055_ = new_n4802_ & new_n10054_;
  assign new_n10056_ = ~new_n10053_ & ~new_n10055_;
  assign new_n10057_ = new_n10051_ & new_n10056_;
  assign new_n10058_ = new_n10043_ & new_n10057_;
  assign new_n10059_ = new_n10024_ & new_n10058_;
  assign new_n10060_ = A235 & new_n186_;
  assign new_n10061_ = new_n960_ & new_n10060_;
  assign new_n10062_ = new_n4802_ & new_n10061_;
  assign new_n10063_ = new_n983_ & new_n10034_;
  assign new_n10064_ = new_n4802_ & new_n10063_;
  assign new_n10065_ = new_n966_ & new_n10060_;
  assign new_n10066_ = new_n4802_ & new_n10065_;
  assign new_n10067_ = ~new_n10064_ & ~new_n10066_;
  assign new_n10068_ = ~new_n10062_ & new_n10067_;
  assign new_n10069_ = new_n971_ & new_n10060_;
  assign new_n10070_ = new_n4802_ & new_n10069_;
  assign new_n10071_ = new_n974_ & new_n10060_;
  assign new_n10072_ = new_n4802_ & new_n10071_;
  assign new_n10073_ = new_n977_ & new_n10060_;
  assign new_n10074_ = new_n4802_ & new_n10073_;
  assign new_n10075_ = ~new_n10072_ & ~new_n10074_;
  assign new_n10076_ = ~new_n10070_ & new_n10075_;
  assign new_n10077_ = new_n10068_ & new_n10076_;
  assign new_n10078_ = new_n983_ & new_n10060_;
  assign new_n10079_ = new_n4802_ & new_n10078_;
  assign new_n10080_ = new_n986_ & new_n10060_;
  assign new_n10081_ = new_n4802_ & new_n10080_;
  assign new_n10082_ = new_n989_ & new_n10060_;
  assign new_n10083_ = new_n4802_ & new_n10082_;
  assign new_n10084_ = ~new_n10081_ & ~new_n10083_;
  assign new_n10085_ = ~new_n10079_ & new_n10084_;
  assign new_n10086_ = A235 & new_n209_;
  assign new_n10087_ = new_n947_ & new_n10086_;
  assign new_n10088_ = new_n4802_ & new_n10087_;
  assign new_n10089_ = new_n950_ & new_n10086_;
  assign new_n10090_ = new_n4802_ & new_n10089_;
  assign new_n10091_ = new_n953_ & new_n10086_;
  assign new_n10092_ = new_n4802_ & new_n10091_;
  assign new_n10093_ = ~new_n10090_ & ~new_n10092_;
  assign new_n10094_ = ~new_n10088_ & new_n10093_;
  assign new_n10095_ = new_n10085_ & new_n10094_;
  assign new_n10096_ = new_n10077_ & new_n10095_;
  assign new_n10097_ = A235 & new_n218_;
  assign new_n10098_ = new_n953_ & new_n10097_;
  assign new_n10099_ = new_n4802_ & new_n10098_;
  assign new_n10100_ = new_n963_ & new_n10086_;
  assign new_n10101_ = new_n4802_ & new_n10100_;
  assign new_n10102_ = new_n950_ & new_n10097_;
  assign new_n10103_ = new_n4802_ & new_n10102_;
  assign new_n10104_ = ~new_n10101_ & ~new_n10103_;
  assign new_n10105_ = ~new_n10099_ & new_n10104_;
  assign new_n10106_ = A235 & new_n236_;
  assign new_n10107_ = new_n950_ & new_n10106_;
  assign new_n10108_ = new_n4802_ & new_n10107_;
  assign new_n10109_ = new_n947_ & new_n10097_;
  assign new_n10110_ = new_n4802_ & new_n10109_;
  assign new_n10111_ = new_n963_ & new_n10097_;
  assign new_n10112_ = new_n4802_ & new_n10111_;
  assign new_n10113_ = ~new_n10110_ & ~new_n10112_;
  assign new_n10114_ = ~new_n10108_ & new_n10113_;
  assign new_n10115_ = new_n10105_ & new_n10114_;
  assign new_n10116_ = new_n963_ & new_n10106_;
  assign new_n10117_ = new_n4802_ & new_n10116_;
  assign new_n10118_ = new_n953_ & new_n10106_;
  assign new_n10119_ = new_n4802_ & new_n10118_;
  assign new_n10120_ = new_n947_ & new_n10106_;
  assign new_n10121_ = new_n4802_ & new_n10120_;
  assign new_n10122_ = ~new_n10119_ & ~new_n10121_;
  assign new_n10123_ = ~new_n10117_ & new_n10122_;
  assign new_n10124_ = ~A266 & new_n153_;
  assign new_n10125_ = new_n1733_ & new_n10124_;
  assign new_n10126_ = ~A232 & ~A200;
  assign new_n10127_ = new_n4623_ & new_n10126_;
  assign new_n10128_ = new_n4968_ & new_n10127_;
  assign new_n10129_ = new_n10125_ & new_n10128_;
  assign new_n10130_ = A266 & new_n153_;
  assign new_n10131_ = new_n1733_ & new_n10130_;
  assign new_n10132_ = new_n4629_ & new_n10126_;
  assign new_n10133_ = new_n4968_ & new_n10132_;
  assign new_n10134_ = new_n10131_ & new_n10133_;
  assign new_n10135_ = ~new_n10129_ & ~new_n10134_;
  assign new_n10136_ = new_n10123_ & new_n10135_;
  assign new_n10137_ = new_n10115_ & new_n10136_;
  assign new_n10138_ = new_n10096_ & new_n10137_;
  assign new_n10139_ = new_n10059_ & new_n10138_;
  assign new_n10140_ = new_n9986_ & new_n10139_;
  assign new_n10141_ = A232 & ~A200;
  assign new_n10142_ = new_n4725_ & new_n10141_;
  assign new_n10143_ = new_n4968_ & new_n10142_;
  assign new_n10144_ = new_n10125_ & new_n10143_;
  assign new_n10145_ = ~A268 & new_n230_;
  assign new_n10146_ = new_n1062_ & new_n10145_;
  assign new_n10147_ = new_n4700_ & new_n10126_;
  assign new_n10148_ = new_n4968_ & new_n10147_;
  assign new_n10149_ = new_n10146_ & new_n10148_;
  assign new_n10150_ = ~A268 & new_n247_;
  assign new_n10151_ = new_n1068_ & new_n10150_;
  assign new_n10152_ = new_n10148_ & new_n10151_;
  assign new_n10153_ = ~new_n10149_ & ~new_n10152_;
  assign new_n10154_ = ~new_n10144_ & new_n10153_;
  assign new_n10155_ = new_n4789_ & new_n10141_;
  assign new_n10156_ = new_n4968_ & new_n10155_;
  assign new_n10157_ = new_n10151_ & new_n10156_;
  assign new_n10158_ = new_n4710_ & new_n10141_;
  assign new_n10159_ = new_n4968_ & new_n10158_;
  assign new_n10160_ = new_n10131_ & new_n10159_;
  assign new_n10161_ = new_n10146_ & new_n10156_;
  assign new_n10162_ = ~new_n10160_ & ~new_n10161_;
  assign new_n10163_ = ~new_n10157_ & new_n10162_;
  assign new_n10164_ = new_n10154_ & new_n10163_;
  assign new_n10165_ = ~A234 & ~A200;
  assign new_n10166_ = new_n261_ & new_n10165_;
  assign new_n10167_ = new_n4968_ & new_n10166_;
  assign new_n10168_ = new_n10146_ & new_n10167_;
  assign new_n10169_ = new_n268_ & new_n10165_;
  assign new_n10170_ = new_n4968_ & new_n10169_;
  assign new_n10171_ = new_n10125_ & new_n10170_;
  assign new_n10172_ = new_n272_ & new_n10165_;
  assign new_n10173_ = new_n4968_ & new_n10172_;
  assign new_n10174_ = new_n10131_ & new_n10173_;
  assign new_n10175_ = ~new_n10171_ & ~new_n10174_;
  assign new_n10176_ = ~new_n10168_ & new_n10175_;
  assign new_n10177_ = new_n280_ & new_n10165_;
  assign new_n10178_ = new_n4968_ & new_n10177_;
  assign new_n10179_ = new_n10131_ & new_n10178_;
  assign new_n10180_ = new_n10151_ & new_n10167_;
  assign new_n10181_ = new_n286_ & new_n10165_;
  assign new_n10182_ = new_n4968_ & new_n10181_;
  assign new_n10183_ = new_n10125_ & new_n10182_;
  assign new_n10184_ = ~new_n10180_ & ~new_n10183_;
  assign new_n10185_ = ~new_n10179_ & new_n10184_;
  assign new_n10186_ = new_n10176_ & new_n10185_;
  assign new_n10187_ = new_n10164_ & new_n10186_;
  assign new_n10188_ = new_n4969_ & new_n8617_;
  assign new_n10189_ = new_n296_ & new_n10165_;
  assign new_n10190_ = new_n4968_ & new_n10189_;
  assign new_n10191_ = new_n10146_ & new_n10190_;
  assign new_n10192_ = new_n10151_ & new_n10190_;
  assign new_n10193_ = ~new_n10191_ & ~new_n10192_;
  assign new_n10194_ = ~new_n10188_ & new_n10193_;
  assign new_n10195_ = new_n4969_ & new_n8625_;
  assign new_n10196_ = new_n4969_ & new_n8628_;
  assign new_n10197_ = new_n4969_ & new_n8630_;
  assign new_n10198_ = ~new_n10196_ & ~new_n10197_;
  assign new_n10199_ = ~new_n10195_ & new_n10198_;
  assign new_n10200_ = new_n10194_ & new_n10199_;
  assign new_n10201_ = new_n4969_ & new_n8635_;
  assign new_n10202_ = new_n4969_ & new_n8637_;
  assign new_n10203_ = new_n4969_ & new_n8639_;
  assign new_n10204_ = ~new_n10202_ & ~new_n10203_;
  assign new_n10205_ = ~new_n10201_ & new_n10204_;
  assign new_n10206_ = new_n4969_ & new_n8648_;
  assign new_n10207_ = new_n4969_ & new_n8650_;
  assign new_n10208_ = ~new_n10206_ & ~new_n10207_;
  assign new_n10209_ = new_n10205_ & new_n10208_;
  assign new_n10210_ = new_n10200_ & new_n10209_;
  assign new_n10211_ = new_n10187_ & new_n10210_;
  assign new_n10212_ = new_n4969_ & new_n8659_;
  assign new_n10213_ = new_n4969_ & new_n8646_;
  assign new_n10214_ = new_n4969_ & new_n8657_;
  assign new_n10215_ = ~new_n10213_ & ~new_n10214_;
  assign new_n10216_ = ~new_n10212_ & new_n10215_;
  assign new_n10217_ = new_n4969_ & new_n8670_;
  assign new_n10218_ = new_n4969_ & new_n8655_;
  assign new_n10219_ = new_n4969_ & new_n8667_;
  assign new_n10220_ = ~new_n10218_ & ~new_n10219_;
  assign new_n10221_ = ~new_n10217_ & new_n10220_;
  assign new_n10222_ = new_n10216_ & new_n10221_;
  assign new_n10223_ = new_n4969_ & new_n8681_;
  assign new_n10224_ = new_n4969_ & new_n8665_;
  assign new_n10225_ = new_n4969_ & new_n8678_;
  assign new_n10226_ = ~new_n10224_ & ~new_n10225_;
  assign new_n10227_ = ~new_n10223_ & new_n10226_;
  assign new_n10228_ = new_n4969_ & new_n8694_;
  assign new_n10229_ = new_n4969_ & new_n8675_;
  assign new_n10230_ = new_n4969_ & new_n8692_;
  assign new_n10231_ = ~new_n10229_ & ~new_n10230_;
  assign new_n10232_ = ~new_n10228_ & new_n10231_;
  assign new_n10233_ = new_n10227_ & new_n10232_;
  assign new_n10234_ = new_n10222_ & new_n10233_;
  assign new_n10235_ = new_n4969_ & new_n8701_;
  assign new_n10236_ = new_n4969_ & new_n8689_;
  assign new_n10237_ = new_n4969_ & new_n8699_;
  assign new_n10238_ = ~new_n10236_ & ~new_n10237_;
  assign new_n10239_ = ~new_n10235_ & new_n10238_;
  assign new_n10240_ = ~A232 & A200;
  assign new_n10241_ = new_n4700_ & new_n10240_;
  assign new_n10242_ = new_n4983_ & new_n10241_;
  assign new_n10243_ = new_n10146_ & new_n10242_;
  assign new_n10244_ = new_n4623_ & new_n10240_;
  assign new_n10245_ = new_n4983_ & new_n10244_;
  assign new_n10246_ = new_n10125_ & new_n10245_;
  assign new_n10247_ = new_n4629_ & new_n10240_;
  assign new_n10248_ = new_n4983_ & new_n10247_;
  assign new_n10249_ = new_n10131_ & new_n10248_;
  assign new_n10250_ = ~new_n10246_ & ~new_n10249_;
  assign new_n10251_ = ~new_n10243_ & new_n10250_;
  assign new_n10252_ = new_n10239_ & new_n10251_;
  assign new_n10253_ = A232 & A200;
  assign new_n10254_ = new_n4710_ & new_n10253_;
  assign new_n10255_ = new_n4983_ & new_n10254_;
  assign new_n10256_ = new_n10131_ & new_n10255_;
  assign new_n10257_ = new_n10151_ & new_n10242_;
  assign new_n10258_ = new_n4725_ & new_n10253_;
  assign new_n10259_ = new_n4983_ & new_n10258_;
  assign new_n10260_ = new_n10125_ & new_n10259_;
  assign new_n10261_ = ~new_n10257_ & ~new_n10260_;
  assign new_n10262_ = ~new_n10256_ & new_n10261_;
  assign new_n10263_ = new_n4789_ & new_n10253_;
  assign new_n10264_ = new_n4983_ & new_n10263_;
  assign new_n10265_ = new_n10146_ & new_n10264_;
  assign new_n10266_ = new_n10151_ & new_n10264_;
  assign new_n10267_ = ~new_n10265_ & ~new_n10266_;
  assign new_n10268_ = new_n10262_ & new_n10267_;
  assign new_n10269_ = new_n10252_ & new_n10268_;
  assign new_n10270_ = new_n10234_ & new_n10269_;
  assign new_n10271_ = new_n10211_ & new_n10270_;
  assign new_n10272_ = ~A234 & A200;
  assign new_n10273_ = new_n261_ & new_n10272_;
  assign new_n10274_ = new_n4983_ & new_n10273_;
  assign new_n10275_ = new_n10146_ & new_n10274_;
  assign new_n10276_ = new_n268_ & new_n10272_;
  assign new_n10277_ = new_n4983_ & new_n10276_;
  assign new_n10278_ = new_n10125_ & new_n10277_;
  assign new_n10279_ = new_n272_ & new_n10272_;
  assign new_n10280_ = new_n4983_ & new_n10279_;
  assign new_n10281_ = new_n10131_ & new_n10280_;
  assign new_n10282_ = ~new_n10278_ & ~new_n10281_;
  assign new_n10283_ = ~new_n10275_ & new_n10282_;
  assign new_n10284_ = new_n280_ & new_n10272_;
  assign new_n10285_ = new_n4983_ & new_n10284_;
  assign new_n10286_ = new_n10131_ & new_n10285_;
  assign new_n10287_ = new_n10151_ & new_n10274_;
  assign new_n10288_ = new_n286_ & new_n10272_;
  assign new_n10289_ = new_n4983_ & new_n10288_;
  assign new_n10290_ = new_n10125_ & new_n10289_;
  assign new_n10291_ = ~new_n10287_ & ~new_n10290_;
  assign new_n10292_ = ~new_n10286_ & new_n10291_;
  assign new_n10293_ = new_n10283_ & new_n10292_;
  assign new_n10294_ = new_n4984_ & new_n8617_;
  assign new_n10295_ = new_n296_ & new_n10272_;
  assign new_n10296_ = new_n4983_ & new_n10295_;
  assign new_n10297_ = new_n10146_ & new_n10296_;
  assign new_n10298_ = new_n10151_ & new_n10296_;
  assign new_n10299_ = ~new_n10297_ & ~new_n10298_;
  assign new_n10300_ = ~new_n10294_ & new_n10299_;
  assign new_n10301_ = new_n4984_ & new_n8625_;
  assign new_n10302_ = new_n4984_ & new_n8628_;
  assign new_n10303_ = new_n4984_ & new_n8630_;
  assign new_n10304_ = ~new_n10302_ & ~new_n10303_;
  assign new_n10305_ = ~new_n10301_ & new_n10304_;
  assign new_n10306_ = new_n10300_ & new_n10305_;
  assign new_n10307_ = new_n10293_ & new_n10306_;
  assign new_n10308_ = new_n4984_ & new_n8635_;
  assign new_n10309_ = new_n4984_ & new_n8637_;
  assign new_n10310_ = new_n4984_ & new_n8639_;
  assign new_n10311_ = ~new_n10309_ & ~new_n10310_;
  assign new_n10312_ = ~new_n10308_ & new_n10311_;
  assign new_n10313_ = new_n4984_ & new_n8646_;
  assign new_n10314_ = new_n4984_ & new_n8648_;
  assign new_n10315_ = new_n4984_ & new_n8650_;
  assign new_n10316_ = ~new_n10314_ & ~new_n10315_;
  assign new_n10317_ = ~new_n10313_ & new_n10316_;
  assign new_n10318_ = new_n10312_ & new_n10317_;
  assign new_n10319_ = new_n4984_ & new_n8655_;
  assign new_n10320_ = new_n4984_ & new_n8657_;
  assign new_n10321_ = new_n4984_ & new_n8659_;
  assign new_n10322_ = ~new_n10320_ & ~new_n10321_;
  assign new_n10323_ = ~new_n10319_ & new_n10322_;
  assign new_n10324_ = new_n4984_ & new_n8667_;
  assign new_n10325_ = new_n4984_ & new_n8670_;
  assign new_n10326_ = ~new_n10324_ & ~new_n10325_;
  assign new_n10327_ = new_n10323_ & new_n10326_;
  assign new_n10328_ = new_n10318_ & new_n10327_;
  assign new_n10329_ = new_n10307_ & new_n10328_;
  assign new_n10330_ = new_n4984_ & new_n8681_;
  assign new_n10331_ = new_n4984_ & new_n8665_;
  assign new_n10332_ = new_n4984_ & new_n8678_;
  assign new_n10333_ = ~new_n10331_ & ~new_n10332_;
  assign new_n10334_ = ~new_n10330_ & new_n10333_;
  assign new_n10335_ = new_n4984_ & new_n8694_;
  assign new_n10336_ = new_n4984_ & new_n8675_;
  assign new_n10337_ = new_n4984_ & new_n8692_;
  assign new_n10338_ = ~new_n10336_ & ~new_n10337_;
  assign new_n10339_ = ~new_n10335_ & new_n10338_;
  assign new_n10340_ = new_n10334_ & new_n10339_;
  assign new_n10341_ = new_n4984_ & new_n8701_;
  assign new_n10342_ = new_n4984_ & new_n8689_;
  assign new_n10343_ = new_n4984_ & new_n8699_;
  assign new_n10344_ = ~new_n10342_ & ~new_n10343_;
  assign new_n10345_ = ~new_n10341_ & new_n10344_;
  assign new_n10346_ = new_n4700_ & new_n7214_;
  assign new_n10347_ = new_n4992_ & new_n10346_;
  assign new_n10348_ = new_n10146_ & new_n10347_;
  assign new_n10349_ = new_n4623_ & new_n7214_;
  assign new_n10350_ = new_n4992_ & new_n10349_;
  assign new_n10351_ = new_n10125_ & new_n10350_;
  assign new_n10352_ = new_n4629_ & new_n7214_;
  assign new_n10353_ = new_n4992_ & new_n10352_;
  assign new_n10354_ = new_n10131_ & new_n10353_;
  assign new_n10355_ = ~new_n10351_ & ~new_n10354_;
  assign new_n10356_ = ~new_n10348_ & new_n10355_;
  assign new_n10357_ = new_n10345_ & new_n10356_;
  assign new_n10358_ = new_n10340_ & new_n10357_;
  assign new_n10359_ = new_n4710_ & new_n7045_;
  assign new_n10360_ = new_n4992_ & new_n10359_;
  assign new_n10361_ = new_n10131_ & new_n10360_;
  assign new_n10362_ = new_n10151_ & new_n10347_;
  assign new_n10363_ = new_n4725_ & new_n7045_;
  assign new_n10364_ = new_n4992_ & new_n10363_;
  assign new_n10365_ = new_n10125_ & new_n10364_;
  assign new_n10366_ = ~new_n10362_ & ~new_n10365_;
  assign new_n10367_ = ~new_n10361_ & new_n10366_;
  assign new_n10368_ = ~A234 & ~A203;
  assign new_n10369_ = new_n268_ & new_n10368_;
  assign new_n10370_ = new_n4992_ & new_n10369_;
  assign new_n10371_ = new_n10125_ & new_n10370_;
  assign new_n10372_ = new_n4789_ & new_n7045_;
  assign new_n10373_ = new_n4992_ & new_n10372_;
  assign new_n10374_ = new_n10146_ & new_n10373_;
  assign new_n10375_ = new_n10151_ & new_n10373_;
  assign new_n10376_ = ~new_n10374_ & ~new_n10375_;
  assign new_n10377_ = ~new_n10371_ & new_n10376_;
  assign new_n10378_ = new_n10367_ & new_n10377_;
  assign new_n10379_ = new_n261_ & new_n10368_;
  assign new_n10380_ = new_n4992_ & new_n10379_;
  assign new_n10381_ = new_n10151_ & new_n10380_;
  assign new_n10382_ = new_n272_ & new_n10368_;
  assign new_n10383_ = new_n4992_ & new_n10382_;
  assign new_n10384_ = new_n10131_ & new_n10383_;
  assign new_n10385_ = new_n10146_ & new_n10380_;
  assign new_n10386_ = ~new_n10384_ & ~new_n10385_;
  assign new_n10387_ = ~new_n10381_ & new_n10386_;
  assign new_n10388_ = new_n286_ & new_n10368_;
  assign new_n10389_ = new_n4992_ & new_n10388_;
  assign new_n10390_ = new_n10125_ & new_n10389_;
  assign new_n10391_ = new_n280_ & new_n10368_;
  assign new_n10392_ = new_n4992_ & new_n10391_;
  assign new_n10393_ = new_n10131_ & new_n10392_;
  assign new_n10394_ = ~new_n10390_ & ~new_n10393_;
  assign new_n10395_ = new_n10387_ & new_n10394_;
  assign new_n10396_ = new_n10378_ & new_n10395_;
  assign new_n10397_ = new_n10358_ & new_n10396_;
  assign new_n10398_ = new_n10329_ & new_n10397_;
  assign new_n10399_ = new_n10271_ & new_n10398_;
  assign new_n10400_ = new_n10140_ & new_n10399_;
  assign new_n10401_ = new_n4993_ & new_n8617_;
  assign new_n10402_ = new_n296_ & new_n10368_;
  assign new_n10403_ = new_n4992_ & new_n10402_;
  assign new_n10404_ = new_n10146_ & new_n10403_;
  assign new_n10405_ = new_n10151_ & new_n10403_;
  assign new_n10406_ = ~new_n10404_ & ~new_n10405_;
  assign new_n10407_ = ~new_n10401_ & new_n10406_;
  assign new_n10408_ = new_n4993_ & new_n8625_;
  assign new_n10409_ = new_n4993_ & new_n8628_;
  assign new_n10410_ = new_n4993_ & new_n8630_;
  assign new_n10411_ = ~new_n10409_ & ~new_n10410_;
  assign new_n10412_ = ~new_n10408_ & new_n10411_;
  assign new_n10413_ = new_n10407_ & new_n10412_;
  assign new_n10414_ = new_n4993_ & new_n8635_;
  assign new_n10415_ = new_n4993_ & new_n8637_;
  assign new_n10416_ = new_n4993_ & new_n8639_;
  assign new_n10417_ = ~new_n10415_ & ~new_n10416_;
  assign new_n10418_ = ~new_n10414_ & new_n10417_;
  assign new_n10419_ = new_n4993_ & new_n8646_;
  assign new_n10420_ = new_n4993_ & new_n8648_;
  assign new_n10421_ = new_n4993_ & new_n8650_;
  assign new_n10422_ = ~new_n10420_ & ~new_n10421_;
  assign new_n10423_ = ~new_n10419_ & new_n10422_;
  assign new_n10424_ = new_n10418_ & new_n10423_;
  assign new_n10425_ = new_n10413_ & new_n10424_;
  assign new_n10426_ = new_n4993_ & new_n8655_;
  assign new_n10427_ = new_n4993_ & new_n8657_;
  assign new_n10428_ = new_n4993_ & new_n8659_;
  assign new_n10429_ = ~new_n10427_ & ~new_n10428_;
  assign new_n10430_ = ~new_n10426_ & new_n10429_;
  assign new_n10431_ = new_n4993_ & new_n8665_;
  assign new_n10432_ = new_n4993_ & new_n8667_;
  assign new_n10433_ = new_n4993_ & new_n8670_;
  assign new_n10434_ = ~new_n10432_ & ~new_n10433_;
  assign new_n10435_ = ~new_n10431_ & new_n10434_;
  assign new_n10436_ = new_n10430_ & new_n10435_;
  assign new_n10437_ = new_n4993_ & new_n8675_;
  assign new_n10438_ = new_n4993_ & new_n8678_;
  assign new_n10439_ = new_n4993_ & new_n8681_;
  assign new_n10440_ = ~new_n10438_ & ~new_n10439_;
  assign new_n10441_ = ~new_n10437_ & new_n10440_;
  assign new_n10442_ = new_n4993_ & new_n8689_;
  assign new_n10443_ = new_n4993_ & new_n8692_;
  assign new_n10444_ = new_n4993_ & new_n8694_;
  assign new_n10445_ = ~new_n10443_ & ~new_n10444_;
  assign new_n10446_ = ~new_n10442_ & new_n10445_;
  assign new_n10447_ = new_n10441_ & new_n10446_;
  assign new_n10448_ = new_n10436_ & new_n10447_;
  assign new_n10449_ = new_n10425_ & new_n10448_;
  assign new_n10450_ = new_n4623_ & new_n7543_;
  assign new_n10451_ = new_n4992_ & new_n10450_;
  assign new_n10452_ = new_n10125_ & new_n10451_;
  assign new_n10453_ = new_n4993_ & new_n8699_;
  assign new_n10454_ = new_n4993_ & new_n8701_;
  assign new_n10455_ = ~new_n10453_ & ~new_n10454_;
  assign new_n10456_ = ~new_n10452_ & new_n10455_;
  assign new_n10457_ = new_n4700_ & new_n7543_;
  assign new_n10458_ = new_n4992_ & new_n10457_;
  assign new_n10459_ = new_n10151_ & new_n10458_;
  assign new_n10460_ = new_n4629_ & new_n7543_;
  assign new_n10461_ = new_n4992_ & new_n10460_;
  assign new_n10462_ = new_n10131_ & new_n10461_;
  assign new_n10463_ = new_n10146_ & new_n10458_;
  assign new_n10464_ = ~new_n10462_ & ~new_n10463_;
  assign new_n10465_ = ~new_n10459_ & new_n10464_;
  assign new_n10466_ = new_n10456_ & new_n10465_;
  assign new_n10467_ = new_n4789_ & new_n7374_;
  assign new_n10468_ = new_n4992_ & new_n10467_;
  assign new_n10469_ = new_n10146_ & new_n10468_;
  assign new_n10470_ = new_n4725_ & new_n7374_;
  assign new_n10471_ = new_n4992_ & new_n10470_;
  assign new_n10472_ = new_n10125_ & new_n10471_;
  assign new_n10473_ = new_n4710_ & new_n7374_;
  assign new_n10474_ = new_n4992_ & new_n10473_;
  assign new_n10475_ = new_n10131_ & new_n10474_;
  assign new_n10476_ = ~new_n10472_ & ~new_n10475_;
  assign new_n10477_ = ~new_n10469_ & new_n10476_;
  assign new_n10478_ = ~A234 & A202;
  assign new_n10479_ = new_n272_ & new_n10478_;
  assign new_n10480_ = new_n4992_ & new_n10479_;
  assign new_n10481_ = new_n10131_ & new_n10480_;
  assign new_n10482_ = new_n10151_ & new_n10468_;
  assign new_n10483_ = new_n268_ & new_n10478_;
  assign new_n10484_ = new_n4992_ & new_n10483_;
  assign new_n10485_ = new_n10125_ & new_n10484_;
  assign new_n10486_ = ~new_n10482_ & ~new_n10485_;
  assign new_n10487_ = ~new_n10481_ & new_n10486_;
  assign new_n10488_ = new_n10477_ & new_n10487_;
  assign new_n10489_ = new_n10466_ & new_n10488_;
  assign new_n10490_ = new_n286_ & new_n10478_;
  assign new_n10491_ = new_n4992_ & new_n10490_;
  assign new_n10492_ = new_n10125_ & new_n10491_;
  assign new_n10493_ = new_n261_ & new_n10478_;
  assign new_n10494_ = new_n4992_ & new_n10493_;
  assign new_n10495_ = new_n10146_ & new_n10494_;
  assign new_n10496_ = new_n10151_ & new_n10494_;
  assign new_n10497_ = ~new_n10495_ & ~new_n10496_;
  assign new_n10498_ = ~new_n10492_ & new_n10497_;
  assign new_n10499_ = new_n296_ & new_n10478_;
  assign new_n10500_ = new_n4992_ & new_n10499_;
  assign new_n10501_ = new_n10151_ & new_n10500_;
  assign new_n10502_ = new_n280_ & new_n10478_;
  assign new_n10503_ = new_n4992_ & new_n10502_;
  assign new_n10504_ = new_n10131_ & new_n10503_;
  assign new_n10505_ = new_n10146_ & new_n10500_;
  assign new_n10506_ = ~new_n10504_ & ~new_n10505_;
  assign new_n10507_ = ~new_n10501_ & new_n10506_;
  assign new_n10508_ = new_n10498_ & new_n10507_;
  assign new_n10509_ = new_n4999_ & new_n8630_;
  assign new_n10510_ = new_n4999_ & new_n8617_;
  assign new_n10511_ = new_n4999_ & new_n8628_;
  assign new_n10512_ = ~new_n10510_ & ~new_n10511_;
  assign new_n10513_ = ~new_n10509_ & new_n10512_;
  assign new_n10514_ = new_n4999_ & new_n8625_;
  assign new_n10515_ = new_n4999_ & new_n8637_;
  assign new_n10516_ = ~new_n10514_ & ~new_n10515_;
  assign new_n10517_ = new_n10513_ & new_n10516_;
  assign new_n10518_ = new_n10508_ & new_n10517_;
  assign new_n10519_ = new_n10489_ & new_n10518_;
  assign new_n10520_ = new_n10449_ & new_n10519_;
  assign new_n10521_ = new_n4999_ & new_n8648_;
  assign new_n10522_ = new_n4999_ & new_n8639_;
  assign new_n10523_ = new_n4999_ & new_n8635_;
  assign new_n10524_ = ~new_n10522_ & ~new_n10523_;
  assign new_n10525_ = ~new_n10521_ & new_n10524_;
  assign new_n10526_ = new_n4999_ & new_n8657_;
  assign new_n10527_ = new_n4999_ & new_n8650_;
  assign new_n10528_ = new_n4999_ & new_n8646_;
  assign new_n10529_ = ~new_n10527_ & ~new_n10528_;
  assign new_n10530_ = ~new_n10526_ & new_n10529_;
  assign new_n10531_ = new_n10525_ & new_n10530_;
  assign new_n10532_ = new_n4999_ & new_n8667_;
  assign new_n10533_ = new_n4999_ & new_n8659_;
  assign new_n10534_ = new_n4999_ & new_n8655_;
  assign new_n10535_ = ~new_n10533_ & ~new_n10534_;
  assign new_n10536_ = ~new_n10532_ & new_n10535_;
  assign new_n10537_ = new_n4999_ & new_n8678_;
  assign new_n10538_ = new_n4999_ & new_n8670_;
  assign new_n10539_ = new_n4999_ & new_n8665_;
  assign new_n10540_ = ~new_n10538_ & ~new_n10539_;
  assign new_n10541_ = ~new_n10537_ & new_n10540_;
  assign new_n10542_ = new_n10536_ & new_n10541_;
  assign new_n10543_ = new_n10531_ & new_n10542_;
  assign new_n10544_ = new_n4999_ & new_n8692_;
  assign new_n10545_ = new_n4999_ & new_n8681_;
  assign new_n10546_ = new_n4999_ & new_n8675_;
  assign new_n10547_ = ~new_n10545_ & ~new_n10546_;
  assign new_n10548_ = ~new_n10544_ & new_n10547_;
  assign new_n10549_ = new_n4999_ & new_n8699_;
  assign new_n10550_ = new_n4999_ & new_n8694_;
  assign new_n10551_ = new_n4999_ & new_n8689_;
  assign new_n10552_ = ~new_n10550_ & ~new_n10551_;
  assign new_n10553_ = ~new_n10549_ & new_n10552_;
  assign new_n10554_ = new_n10548_ & new_n10553_;
  assign new_n10555_ = new_n5014_ & new_n8628_;
  assign new_n10556_ = new_n4999_ & new_n8701_;
  assign new_n10557_ = new_n5014_ & new_n8617_;
  assign new_n10558_ = ~new_n10556_ & ~new_n10557_;
  assign new_n10559_ = ~new_n10555_ & new_n10558_;
  assign new_n10560_ = new_n5014_ & new_n8630_;
  assign new_n10561_ = new_n5014_ & new_n8625_;
  assign new_n10562_ = ~new_n10560_ & ~new_n10561_;
  assign new_n10563_ = new_n10559_ & new_n10562_;
  assign new_n10564_ = new_n10554_ & new_n10563_;
  assign new_n10565_ = new_n10543_ & new_n10564_;
  assign new_n10566_ = new_n5014_ & new_n8635_;
  assign new_n10567_ = new_n5014_ & new_n8637_;
  assign new_n10568_ = new_n5014_ & new_n8639_;
  assign new_n10569_ = ~new_n10567_ & ~new_n10568_;
  assign new_n10570_ = ~new_n10566_ & new_n10569_;
  assign new_n10571_ = new_n5014_ & new_n8646_;
  assign new_n10572_ = new_n5014_ & new_n8648_;
  assign new_n10573_ = new_n5014_ & new_n8650_;
  assign new_n10574_ = ~new_n10572_ & ~new_n10573_;
  assign new_n10575_ = ~new_n10571_ & new_n10574_;
  assign new_n10576_ = new_n10570_ & new_n10575_;
  assign new_n10577_ = new_n5014_ & new_n8655_;
  assign new_n10578_ = new_n5014_ & new_n8657_;
  assign new_n10579_ = new_n5014_ & new_n8659_;
  assign new_n10580_ = ~new_n10578_ & ~new_n10579_;
  assign new_n10581_ = ~new_n10577_ & new_n10580_;
  assign new_n10582_ = new_n5014_ & new_n8665_;
  assign new_n10583_ = new_n5014_ & new_n8667_;
  assign new_n10584_ = new_n5014_ & new_n8670_;
  assign new_n10585_ = ~new_n10583_ & ~new_n10584_;
  assign new_n10586_ = ~new_n10582_ & new_n10585_;
  assign new_n10587_ = new_n10581_ & new_n10586_;
  assign new_n10588_ = new_n10576_ & new_n10587_;
  assign new_n10589_ = new_n5014_ & new_n8675_;
  assign new_n10590_ = new_n5014_ & new_n8678_;
  assign new_n10591_ = new_n5014_ & new_n8681_;
  assign new_n10592_ = ~new_n10590_ & ~new_n10591_;
  assign new_n10593_ = ~new_n10589_ & new_n10592_;
  assign new_n10594_ = new_n5014_ & new_n8689_;
  assign new_n10595_ = new_n5014_ & new_n8692_;
  assign new_n10596_ = new_n5014_ & new_n8694_;
  assign new_n10597_ = ~new_n10595_ & ~new_n10596_;
  assign new_n10598_ = ~new_n10594_ & new_n10597_;
  assign new_n10599_ = new_n10593_ & new_n10598_;
  assign new_n10600_ = new_n5021_ & new_n8617_;
  assign new_n10601_ = new_n5014_ & new_n8699_;
  assign new_n10602_ = new_n5014_ & new_n8701_;
  assign new_n10603_ = ~new_n10601_ & ~new_n10602_;
  assign new_n10604_ = ~new_n10600_ & new_n10603_;
  assign new_n10605_ = new_n5021_ & new_n8628_;
  assign new_n10606_ = new_n5021_ & new_n8630_;
  assign new_n10607_ = ~new_n10605_ & ~new_n10606_;
  assign new_n10608_ = new_n10604_ & new_n10607_;
  assign new_n10609_ = new_n10599_ & new_n10608_;
  assign new_n10610_ = new_n10588_ & new_n10609_;
  assign new_n10611_ = new_n10565_ & new_n10610_;
  assign new_n10612_ = new_n10520_ & new_n10611_;
  assign new_n10613_ = new_n5021_ & new_n8639_;
  assign new_n10614_ = new_n5021_ & new_n8625_;
  assign new_n10615_ = new_n5021_ & new_n8637_;
  assign new_n10616_ = ~new_n10614_ & ~new_n10615_;
  assign new_n10617_ = ~new_n10613_ & new_n10616_;
  assign new_n10618_ = new_n5021_ & new_n8650_;
  assign new_n10619_ = new_n5021_ & new_n8635_;
  assign new_n10620_ = new_n5021_ & new_n8648_;
  assign new_n10621_ = ~new_n10619_ & ~new_n10620_;
  assign new_n10622_ = ~new_n10618_ & new_n10621_;
  assign new_n10623_ = new_n10617_ & new_n10622_;
  assign new_n10624_ = new_n5021_ & new_n8659_;
  assign new_n10625_ = new_n5021_ & new_n8646_;
  assign new_n10626_ = new_n5021_ & new_n8657_;
  assign new_n10627_ = ~new_n10625_ & ~new_n10626_;
  assign new_n10628_ = ~new_n10624_ & new_n10627_;
  assign new_n10629_ = new_n5021_ & new_n8670_;
  assign new_n10630_ = new_n5021_ & new_n8655_;
  assign new_n10631_ = new_n5021_ & new_n8667_;
  assign new_n10632_ = ~new_n10630_ & ~new_n10631_;
  assign new_n10633_ = ~new_n10629_ & new_n10632_;
  assign new_n10634_ = new_n10628_ & new_n10633_;
  assign new_n10635_ = new_n10623_ & new_n10634_;
  assign new_n10636_ = new_n5021_ & new_n8681_;
  assign new_n10637_ = new_n5021_ & new_n8665_;
  assign new_n10638_ = new_n5021_ & new_n8678_;
  assign new_n10639_ = ~new_n10637_ & ~new_n10638_;
  assign new_n10640_ = ~new_n10636_ & new_n10639_;
  assign new_n10641_ = new_n5021_ & new_n8694_;
  assign new_n10642_ = new_n5021_ & new_n8675_;
  assign new_n10643_ = new_n5021_ & new_n8692_;
  assign new_n10644_ = ~new_n10642_ & ~new_n10643_;
  assign new_n10645_ = ~new_n10641_ & new_n10644_;
  assign new_n10646_ = new_n10640_ & new_n10645_;
  assign new_n10647_ = new_n5021_ & new_n8701_;
  assign new_n10648_ = new_n5021_ & new_n8689_;
  assign new_n10649_ = new_n5021_ & new_n8699_;
  assign new_n10650_ = ~new_n10648_ & ~new_n10649_;
  assign new_n10651_ = ~new_n10647_ & new_n10650_;
  assign new_n10652_ = new_n5033_ & new_n8617_;
  assign new_n10653_ = new_n5033_ & new_n8628_;
  assign new_n10654_ = ~new_n10652_ & ~new_n10653_;
  assign new_n10655_ = new_n10651_ & new_n10654_;
  assign new_n10656_ = new_n10646_ & new_n10655_;
  assign new_n10657_ = new_n10635_ & new_n10656_;
  assign new_n10658_ = new_n5033_ & new_n8637_;
  assign new_n10659_ = new_n5033_ & new_n8630_;
  assign new_n10660_ = new_n5033_ & new_n8625_;
  assign new_n10661_ = ~new_n10659_ & ~new_n10660_;
  assign new_n10662_ = ~new_n10658_ & new_n10661_;
  assign new_n10663_ = new_n5033_ & new_n8648_;
  assign new_n10664_ = new_n5033_ & new_n8639_;
  assign new_n10665_ = new_n5033_ & new_n8635_;
  assign new_n10666_ = ~new_n10664_ & ~new_n10665_;
  assign new_n10667_ = ~new_n10663_ & new_n10666_;
  assign new_n10668_ = new_n10662_ & new_n10667_;
  assign new_n10669_ = new_n5033_ & new_n8657_;
  assign new_n10670_ = new_n5033_ & new_n8650_;
  assign new_n10671_ = new_n5033_ & new_n8646_;
  assign new_n10672_ = ~new_n10670_ & ~new_n10671_;
  assign new_n10673_ = ~new_n10669_ & new_n10672_;
  assign new_n10674_ = new_n5033_ & new_n8667_;
  assign new_n10675_ = new_n5033_ & new_n8659_;
  assign new_n10676_ = new_n5033_ & new_n8655_;
  assign new_n10677_ = ~new_n10675_ & ~new_n10676_;
  assign new_n10678_ = ~new_n10674_ & new_n10677_;
  assign new_n10679_ = new_n10673_ & new_n10678_;
  assign new_n10680_ = new_n10668_ & new_n10679_;
  assign new_n10681_ = new_n5033_ & new_n8678_;
  assign new_n10682_ = new_n5033_ & new_n8670_;
  assign new_n10683_ = new_n5033_ & new_n8665_;
  assign new_n10684_ = ~new_n10682_ & ~new_n10683_;
  assign new_n10685_ = ~new_n10681_ & new_n10684_;
  assign new_n10686_ = new_n5033_ & new_n8692_;
  assign new_n10687_ = new_n5033_ & new_n8681_;
  assign new_n10688_ = new_n5033_ & new_n8675_;
  assign new_n10689_ = ~new_n10687_ & ~new_n10688_;
  assign new_n10690_ = ~new_n10686_ & new_n10689_;
  assign new_n10691_ = new_n10685_ & new_n10690_;
  assign new_n10692_ = new_n5033_ & new_n8699_;
  assign new_n10693_ = new_n5033_ & new_n8694_;
  assign new_n10694_ = new_n5033_ & new_n8689_;
  assign new_n10695_ = ~new_n10693_ & ~new_n10694_;
  assign new_n10696_ = ~new_n10692_ & new_n10695_;
  assign new_n10697_ = new_n5033_ & new_n8701_;
  assign new_n10698_ = new_n5039_ & new_n8617_;
  assign new_n10699_ = ~new_n10697_ & ~new_n10698_;
  assign new_n10700_ = new_n10696_ & new_n10699_;
  assign new_n10701_ = new_n10691_ & new_n10700_;
  assign new_n10702_ = new_n10680_ & new_n10701_;
  assign new_n10703_ = new_n10657_ & new_n10702_;
  assign new_n10704_ = new_n5039_ & new_n8625_;
  assign new_n10705_ = new_n5039_ & new_n8628_;
  assign new_n10706_ = new_n5039_ & new_n8630_;
  assign new_n10707_ = ~new_n10705_ & ~new_n10706_;
  assign new_n10708_ = ~new_n10704_ & new_n10707_;
  assign new_n10709_ = new_n5039_ & new_n8635_;
  assign new_n10710_ = new_n5039_ & new_n8637_;
  assign new_n10711_ = new_n5039_ & new_n8639_;
  assign new_n10712_ = ~new_n10710_ & ~new_n10711_;
  assign new_n10713_ = ~new_n10709_ & new_n10712_;
  assign new_n10714_ = new_n10708_ & new_n10713_;
  assign new_n10715_ = new_n5039_ & new_n8646_;
  assign new_n10716_ = new_n5039_ & new_n8648_;
  assign new_n10717_ = new_n5039_ & new_n8650_;
  assign new_n10718_ = ~new_n10716_ & ~new_n10717_;
  assign new_n10719_ = ~new_n10715_ & new_n10718_;
  assign new_n10720_ = new_n5039_ & new_n8655_;
  assign new_n10721_ = new_n5039_ & new_n8657_;
  assign new_n10722_ = new_n5039_ & new_n8659_;
  assign new_n10723_ = ~new_n10721_ & ~new_n10722_;
  assign new_n10724_ = ~new_n10720_ & new_n10723_;
  assign new_n10725_ = new_n10719_ & new_n10724_;
  assign new_n10726_ = new_n10714_ & new_n10725_;
  assign new_n10727_ = new_n5039_ & new_n8665_;
  assign new_n10728_ = new_n5039_ & new_n8667_;
  assign new_n10729_ = new_n5039_ & new_n8670_;
  assign new_n10730_ = ~new_n10728_ & ~new_n10729_;
  assign new_n10731_ = ~new_n10727_ & new_n10730_;
  assign new_n10732_ = new_n5039_ & new_n8675_;
  assign new_n10733_ = new_n5039_ & new_n8678_;
  assign new_n10734_ = new_n5039_ & new_n8681_;
  assign new_n10735_ = ~new_n10733_ & ~new_n10734_;
  assign new_n10736_ = ~new_n10732_ & new_n10735_;
  assign new_n10737_ = new_n10731_ & new_n10736_;
  assign new_n10738_ = new_n5039_ & new_n8689_;
  assign new_n10739_ = new_n5039_ & new_n8692_;
  assign new_n10740_ = new_n5039_ & new_n8694_;
  assign new_n10741_ = ~new_n10739_ & ~new_n10740_;
  assign new_n10742_ = ~new_n10738_ & new_n10741_;
  assign new_n10743_ = new_n5039_ & new_n8699_;
  assign new_n10744_ = new_n5039_ & new_n8701_;
  assign new_n10745_ = ~new_n10743_ & ~new_n10744_;
  assign new_n10746_ = new_n10742_ & new_n10745_;
  assign new_n10747_ = new_n10737_ & new_n10746_;
  assign new_n10748_ = new_n10726_ & new_n10747_;
  assign new_n10749_ = new_n5046_ & new_n8855_;
  assign new_n10750_ = new_n5046_ & new_n8845_;
  assign new_n10751_ = new_n5046_ & new_n8853_;
  assign new_n10752_ = ~new_n10750_ & ~new_n10751_;
  assign new_n10753_ = ~new_n10749_ & new_n10752_;
  assign new_n10754_ = new_n5046_ & new_n8866_;
  assign new_n10755_ = new_n5046_ & new_n8851_;
  assign new_n10756_ = new_n5046_ & new_n8864_;
  assign new_n10757_ = ~new_n10755_ & ~new_n10756_;
  assign new_n10758_ = ~new_n10754_ & new_n10757_;
  assign new_n10759_ = new_n10753_ & new_n10758_;
  assign new_n10760_ = new_n5046_ & new_n8874_;
  assign new_n10761_ = new_n5046_ & new_n8862_;
  assign new_n10762_ = new_n5046_ & new_n8872_;
  assign new_n10763_ = ~new_n10761_ & ~new_n10762_;
  assign new_n10764_ = ~new_n10760_ & new_n10763_;
  assign new_n10765_ = new_n5046_ & new_n8884_;
  assign new_n10766_ = new_n5046_ & new_n8870_;
  assign new_n10767_ = new_n5046_ & new_n8882_;
  assign new_n10768_ = ~new_n10766_ & ~new_n10767_;
  assign new_n10769_ = ~new_n10765_ & new_n10768_;
  assign new_n10770_ = new_n10764_ & new_n10769_;
  assign new_n10771_ = new_n10759_ & new_n10770_;
  assign new_n10772_ = new_n5046_ & new_n8890_;
  assign new_n10773_ = new_n5046_ & new_n8880_;
  assign new_n10774_ = new_n5046_ & new_n8888_;
  assign new_n10775_ = ~new_n10773_ & ~new_n10774_;
  assign new_n10776_ = ~new_n10772_ & new_n10775_;
  assign new_n10777_ = new_n5046_ & new_n8896_;
  assign new_n10778_ = new_n5046_ & new_n8898_;
  assign new_n10779_ = new_n5046_ & new_n8900_;
  assign new_n10780_ = ~new_n10778_ & ~new_n10779_;
  assign new_n10781_ = ~new_n10777_ & new_n10780_;
  assign new_n10782_ = new_n10776_ & new_n10781_;
  assign new_n10783_ = new_n5046_ & new_n8905_;
  assign new_n10784_ = new_n5046_ & new_n8907_;
  assign new_n10785_ = new_n5046_ & new_n8909_;
  assign new_n10786_ = ~new_n10784_ & ~new_n10785_;
  assign new_n10787_ = ~new_n10783_ & new_n10786_;
  assign new_n10788_ = new_n5046_ & new_n8916_;
  assign new_n10789_ = new_n5046_ & new_n8918_;
  assign new_n10790_ = ~new_n10788_ & ~new_n10789_;
  assign new_n10791_ = new_n10787_ & new_n10790_;
  assign new_n10792_ = new_n10782_ & new_n10791_;
  assign new_n10793_ = new_n10771_ & new_n10792_;
  assign new_n10794_ = new_n10748_ & new_n10793_;
  assign new_n10795_ = new_n10703_ & new_n10794_;
  assign new_n10796_ = new_n10612_ & new_n10795_;
  assign new_n10797_ = new_n10400_ & new_n10796_;
  assign new_n10798_ = new_n5046_ & new_n8927_;
  assign new_n10799_ = new_n5046_ & new_n8914_;
  assign new_n10800_ = new_n5046_ & new_n8925_;
  assign new_n10801_ = ~new_n10799_ & ~new_n10800_;
  assign new_n10802_ = ~new_n10798_ & new_n10801_;
  assign new_n10803_ = new_n5046_ & new_n8938_;
  assign new_n10804_ = new_n5046_ & new_n8923_;
  assign new_n10805_ = new_n5046_ & new_n8936_;
  assign new_n10806_ = ~new_n10804_ & ~new_n10805_;
  assign new_n10807_ = ~new_n10803_ & new_n10806_;
  assign new_n10808_ = new_n10802_ & new_n10807_;
  assign new_n10809_ = new_n5046_ & new_n8945_;
  assign new_n10810_ = new_n5046_ & new_n8934_;
  assign new_n10811_ = new_n5046_ & new_n8943_;
  assign new_n10812_ = ~new_n10810_ & ~new_n10811_;
  assign new_n10813_ = ~new_n10809_ & new_n10812_;
  assign new_n10814_ = new_n5164_ & new_n9924_;
  assign new_n10815_ = new_n5164_ & new_n9926_;
  assign new_n10816_ = new_n5164_ & new_n9928_;
  assign new_n10817_ = ~new_n10815_ & ~new_n10816_;
  assign new_n10818_ = ~new_n10814_ & new_n10817_;
  assign new_n10819_ = new_n10813_ & new_n10818_;
  assign new_n10820_ = new_n10808_ & new_n10819_;
  assign new_n10821_ = new_n5164_ & new_n9934_;
  assign new_n10822_ = new_n5164_ & new_n9936_;
  assign new_n10823_ = new_n5164_ & new_n9938_;
  assign new_n10824_ = ~new_n10822_ & ~new_n10823_;
  assign new_n10825_ = ~new_n10821_ & new_n10824_;
  assign new_n10826_ = new_n5164_ & new_n9942_;
  assign new_n10827_ = new_n5164_ & new_n9944_;
  assign new_n10828_ = new_n5164_ & new_n9946_;
  assign new_n10829_ = ~new_n10827_ & ~new_n10828_;
  assign new_n10830_ = ~new_n10826_ & new_n10829_;
  assign new_n10831_ = new_n10825_ & new_n10830_;
  assign new_n10832_ = new_n5164_ & new_n9952_;
  assign new_n10833_ = new_n5164_ & new_n9954_;
  assign new_n10834_ = new_n5164_ & new_n9956_;
  assign new_n10835_ = ~new_n10833_ & ~new_n10834_;
  assign new_n10836_ = ~new_n10832_ & new_n10835_;
  assign new_n10837_ = new_n5164_ & new_n9961_;
  assign new_n10838_ = new_n5164_ & new_n9963_;
  assign new_n10839_ = new_n5164_ & new_n9965_;
  assign new_n10840_ = ~new_n10838_ & ~new_n10839_;
  assign new_n10841_ = ~new_n10837_ & new_n10840_;
  assign new_n10842_ = new_n10836_ & new_n10841_;
  assign new_n10843_ = new_n10831_ & new_n10842_;
  assign new_n10844_ = new_n10820_ & new_n10843_;
  assign new_n10845_ = new_n5164_ & new_n9970_;
  assign new_n10846_ = new_n5164_ & new_n9972_;
  assign new_n10847_ = new_n5164_ & new_n9974_;
  assign new_n10848_ = ~new_n10846_ & ~new_n10847_;
  assign new_n10849_ = ~new_n10845_ & new_n10848_;
  assign new_n10850_ = new_n5164_ & new_n9990_;
  assign new_n10851_ = new_n5164_ & new_n9978_;
  assign new_n10852_ = new_n5164_ & new_n9980_;
  assign new_n10853_ = ~new_n10851_ & ~new_n10852_;
  assign new_n10854_ = ~new_n10850_ & new_n10853_;
  assign new_n10855_ = new_n10849_ & new_n10854_;
  assign new_n10856_ = new_n5164_ & new_n9999_;
  assign new_n10857_ = new_n5164_ & new_n9992_;
  assign new_n10858_ = new_n5164_ & new_n9988_;
  assign new_n10859_ = ~new_n10857_ & ~new_n10858_;
  assign new_n10860_ = ~new_n10856_ & new_n10859_;
  assign new_n10861_ = new_n5164_ & new_n10009_;
  assign new_n10862_ = new_n5164_ & new_n10001_;
  assign new_n10863_ = new_n5164_ & new_n9997_;
  assign new_n10864_ = ~new_n10862_ & ~new_n10863_;
  assign new_n10865_ = ~new_n10861_ & new_n10864_;
  assign new_n10866_ = new_n10860_ & new_n10865_;
  assign new_n10867_ = new_n10855_ & new_n10866_;
  assign new_n10868_ = new_n5164_ & new_n10017_;
  assign new_n10869_ = new_n5164_ & new_n10011_;
  assign new_n10870_ = new_n5164_ & new_n10007_;
  assign new_n10871_ = ~new_n10869_ & ~new_n10870_;
  assign new_n10872_ = ~new_n10868_ & new_n10871_;
  assign new_n10873_ = new_n5164_ & new_n10028_;
  assign new_n10874_ = new_n5164_ & new_n10019_;
  assign new_n10875_ = new_n5164_ & new_n10015_;
  assign new_n10876_ = ~new_n10874_ & ~new_n10875_;
  assign new_n10877_ = ~new_n10873_ & new_n10876_;
  assign new_n10878_ = new_n10872_ & new_n10877_;
  assign new_n10879_ = new_n5164_ & new_n10037_;
  assign new_n10880_ = new_n5164_ & new_n10030_;
  assign new_n10881_ = new_n5164_ & new_n10026_;
  assign new_n10882_ = ~new_n10880_ & ~new_n10881_;
  assign new_n10883_ = ~new_n10879_ & new_n10882_;
  assign new_n10884_ = new_n5164_ & new_n10039_;
  assign new_n10885_ = new_n5164_ & new_n10035_;
  assign new_n10886_ = ~new_n10884_ & ~new_n10885_;
  assign new_n10887_ = new_n10883_ & new_n10886_;
  assign new_n10888_ = new_n10878_ & new_n10887_;
  assign new_n10889_ = new_n10867_ & new_n10888_;
  assign new_n10890_ = new_n10844_ & new_n10889_;
  assign new_n10891_ = new_n5164_ & new_n10044_;
  assign new_n10892_ = new_n5164_ & new_n10046_;
  assign new_n10893_ = new_n5164_ & new_n10048_;
  assign new_n10894_ = ~new_n10892_ & ~new_n10893_;
  assign new_n10895_ = ~new_n10891_ & new_n10894_;
  assign new_n10896_ = new_n5164_ & new_n10063_;
  assign new_n10897_ = new_n5164_ & new_n10052_;
  assign new_n10898_ = new_n5164_ & new_n10054_;
  assign new_n10899_ = ~new_n10897_ & ~new_n10898_;
  assign new_n10900_ = ~new_n10896_ & new_n10899_;
  assign new_n10901_ = new_n10895_ & new_n10900_;
  assign new_n10902_ = new_n5164_ & new_n10071_;
  assign new_n10903_ = new_n5164_ & new_n10065_;
  assign new_n10904_ = new_n5164_ & new_n10061_;
  assign new_n10905_ = ~new_n10903_ & ~new_n10904_;
  assign new_n10906_ = ~new_n10902_ & new_n10905_;
  assign new_n10907_ = new_n5164_ & new_n10080_;
  assign new_n10908_ = new_n5164_ & new_n10073_;
  assign new_n10909_ = new_n5164_ & new_n10069_;
  assign new_n10910_ = ~new_n10908_ & ~new_n10909_;
  assign new_n10911_ = ~new_n10907_ & new_n10910_;
  assign new_n10912_ = new_n10906_ & new_n10911_;
  assign new_n10913_ = new_n10901_ & new_n10912_;
  assign new_n10914_ = new_n5164_ & new_n10089_;
  assign new_n10915_ = new_n5164_ & new_n10082_;
  assign new_n10916_ = new_n5164_ & new_n10078_;
  assign new_n10917_ = ~new_n10915_ & ~new_n10916_;
  assign new_n10918_ = ~new_n10914_ & new_n10917_;
  assign new_n10919_ = new_n5164_ & new_n10100_;
  assign new_n10920_ = new_n5164_ & new_n10091_;
  assign new_n10921_ = new_n5164_ & new_n10087_;
  assign new_n10922_ = ~new_n10920_ & ~new_n10921_;
  assign new_n10923_ = ~new_n10919_ & new_n10922_;
  assign new_n10924_ = new_n10918_ & new_n10923_;
  assign new_n10925_ = new_n5164_ & new_n10109_;
  assign new_n10926_ = new_n5164_ & new_n10102_;
  assign new_n10927_ = new_n5164_ & new_n10098_;
  assign new_n10928_ = ~new_n10926_ & ~new_n10927_;
  assign new_n10929_ = ~new_n10925_ & new_n10928_;
  assign new_n10930_ = new_n5164_ & new_n10111_;
  assign new_n10931_ = new_n5164_ & new_n10107_;
  assign new_n10932_ = ~new_n10930_ & ~new_n10931_;
  assign new_n10933_ = new_n10929_ & new_n10932_;
  assign new_n10934_ = new_n10924_ & new_n10933_;
  assign new_n10935_ = new_n10913_ & new_n10934_;
  assign new_n10936_ = new_n5164_ & new_n10116_;
  assign new_n10937_ = new_n5164_ & new_n10118_;
  assign new_n10938_ = new_n5164_ & new_n10120_;
  assign new_n10939_ = ~new_n10937_ & ~new_n10938_;
  assign new_n10940_ = ~new_n10936_ & new_n10939_;
  assign new_n10941_ = new_n5325_ & new_n9924_;
  assign new_n10942_ = new_n5325_ & new_n9926_;
  assign new_n10943_ = new_n5325_ & new_n9928_;
  assign new_n10944_ = ~new_n10942_ & ~new_n10943_;
  assign new_n10945_ = ~new_n10941_ & new_n10944_;
  assign new_n10946_ = new_n10940_ & new_n10945_;
  assign new_n10947_ = new_n5325_ & new_n9934_;
  assign new_n10948_ = new_n5325_ & new_n9936_;
  assign new_n10949_ = new_n5325_ & new_n9938_;
  assign new_n10950_ = ~new_n10948_ & ~new_n10949_;
  assign new_n10951_ = ~new_n10947_ & new_n10950_;
  assign new_n10952_ = new_n5325_ & new_n9942_;
  assign new_n10953_ = new_n5325_ & new_n9944_;
  assign new_n10954_ = new_n5325_ & new_n9946_;
  assign new_n10955_ = ~new_n10953_ & ~new_n10954_;
  assign new_n10956_ = ~new_n10952_ & new_n10955_;
  assign new_n10957_ = new_n10951_ & new_n10956_;
  assign new_n10958_ = new_n10946_ & new_n10957_;
  assign new_n10959_ = new_n5325_ & new_n9952_;
  assign new_n10960_ = new_n5325_ & new_n9954_;
  assign new_n10961_ = new_n5325_ & new_n9956_;
  assign new_n10962_ = ~new_n10960_ & ~new_n10961_;
  assign new_n10963_ = ~new_n10959_ & new_n10962_;
  assign new_n10964_ = new_n5325_ & new_n9961_;
  assign new_n10965_ = new_n5325_ & new_n9963_;
  assign new_n10966_ = new_n5325_ & new_n9965_;
  assign new_n10967_ = ~new_n10965_ & ~new_n10966_;
  assign new_n10968_ = ~new_n10964_ & new_n10967_;
  assign new_n10969_ = new_n10963_ & new_n10968_;
  assign new_n10970_ = new_n5325_ & new_n9970_;
  assign new_n10971_ = new_n5325_ & new_n9972_;
  assign new_n10972_ = new_n5325_ & new_n9974_;
  assign new_n10973_ = ~new_n10971_ & ~new_n10972_;
  assign new_n10974_ = ~new_n10970_ & new_n10973_;
  assign new_n10975_ = new_n5325_ & new_n9978_;
  assign new_n10976_ = new_n5325_ & new_n9980_;
  assign new_n10977_ = ~new_n10975_ & ~new_n10976_;
  assign new_n10978_ = new_n10974_ & new_n10977_;
  assign new_n10979_ = new_n10969_ & new_n10978_;
  assign new_n10980_ = new_n10958_ & new_n10979_;
  assign new_n10981_ = new_n10935_ & new_n10980_;
  assign new_n10982_ = new_n10890_ & new_n10981_;
  assign new_n10983_ = new_n5325_ & new_n9988_;
  assign new_n10984_ = new_n5325_ & new_n9990_;
  assign new_n10985_ = new_n5325_ & new_n9992_;
  assign new_n10986_ = ~new_n10984_ & ~new_n10985_;
  assign new_n10987_ = ~new_n10983_ & new_n10986_;
  assign new_n10988_ = new_n5325_ & new_n9997_;
  assign new_n10989_ = new_n5325_ & new_n9999_;
  assign new_n10990_ = new_n5325_ & new_n10001_;
  assign new_n10991_ = ~new_n10989_ & ~new_n10990_;
  assign new_n10992_ = ~new_n10988_ & new_n10991_;
  assign new_n10993_ = new_n10987_ & new_n10992_;
  assign new_n10994_ = new_n5325_ & new_n10007_;
  assign new_n10995_ = new_n5325_ & new_n10009_;
  assign new_n10996_ = new_n5325_ & new_n10011_;
  assign new_n10997_ = ~new_n10995_ & ~new_n10996_;
  assign new_n10998_ = ~new_n10994_ & new_n10997_;
  assign new_n10999_ = new_n5325_ & new_n10015_;
  assign new_n11000_ = new_n5325_ & new_n10017_;
  assign new_n11001_ = new_n5325_ & new_n10019_;
  assign new_n11002_ = ~new_n11000_ & ~new_n11001_;
  assign new_n11003_ = ~new_n10999_ & new_n11002_;
  assign new_n11004_ = new_n10998_ & new_n11003_;
  assign new_n11005_ = new_n10993_ & new_n11004_;
  assign new_n11006_ = new_n5325_ & new_n10026_;
  assign new_n11007_ = new_n5325_ & new_n10028_;
  assign new_n11008_ = new_n5325_ & new_n10030_;
  assign new_n11009_ = ~new_n11007_ & ~new_n11008_;
  assign new_n11010_ = ~new_n11006_ & new_n11009_;
  assign new_n11011_ = new_n5325_ & new_n10035_;
  assign new_n11012_ = new_n5325_ & new_n10037_;
  assign new_n11013_ = new_n5325_ & new_n10039_;
  assign new_n11014_ = ~new_n11012_ & ~new_n11013_;
  assign new_n11015_ = ~new_n11011_ & new_n11014_;
  assign new_n11016_ = new_n11010_ & new_n11015_;
  assign new_n11017_ = new_n5325_ & new_n10044_;
  assign new_n11018_ = new_n5325_ & new_n10046_;
  assign new_n11019_ = new_n5325_ & new_n10048_;
  assign new_n11020_ = ~new_n11018_ & ~new_n11019_;
  assign new_n11021_ = ~new_n11017_ & new_n11020_;
  assign new_n11022_ = new_n5325_ & new_n10052_;
  assign new_n11023_ = new_n5325_ & new_n10054_;
  assign new_n11024_ = ~new_n11022_ & ~new_n11023_;
  assign new_n11025_ = new_n11021_ & new_n11024_;
  assign new_n11026_ = new_n11016_ & new_n11025_;
  assign new_n11027_ = new_n11005_ & new_n11026_;
  assign new_n11028_ = new_n5325_ & new_n10061_;
  assign new_n11029_ = new_n5325_ & new_n10063_;
  assign new_n11030_ = new_n5325_ & new_n10065_;
  assign new_n11031_ = ~new_n11029_ & ~new_n11030_;
  assign new_n11032_ = ~new_n11028_ & new_n11031_;
  assign new_n11033_ = new_n5325_ & new_n10069_;
  assign new_n11034_ = new_n5325_ & new_n10071_;
  assign new_n11035_ = new_n5325_ & new_n10073_;
  assign new_n11036_ = ~new_n11034_ & ~new_n11035_;
  assign new_n11037_ = ~new_n11033_ & new_n11036_;
  assign new_n11038_ = new_n11032_ & new_n11037_;
  assign new_n11039_ = new_n5325_ & new_n10078_;
  assign new_n11040_ = new_n5325_ & new_n10080_;
  assign new_n11041_ = new_n5325_ & new_n10082_;
  assign new_n11042_ = ~new_n11040_ & ~new_n11041_;
  assign new_n11043_ = ~new_n11039_ & new_n11042_;
  assign new_n11044_ = new_n5325_ & new_n10087_;
  assign new_n11045_ = new_n5325_ & new_n10089_;
  assign new_n11046_ = new_n5325_ & new_n10091_;
  assign new_n11047_ = ~new_n11045_ & ~new_n11046_;
  assign new_n11048_ = ~new_n11044_ & new_n11047_;
  assign new_n11049_ = new_n11043_ & new_n11048_;
  assign new_n11050_ = new_n11038_ & new_n11049_;
  assign new_n11051_ = new_n5325_ & new_n10098_;
  assign new_n11052_ = new_n5325_ & new_n10100_;
  assign new_n11053_ = new_n5325_ & new_n10102_;
  assign new_n11054_ = ~new_n11052_ & ~new_n11053_;
  assign new_n11055_ = ~new_n11051_ & new_n11054_;
  assign new_n11056_ = new_n5325_ & new_n10107_;
  assign new_n11057_ = new_n5325_ & new_n10109_;
  assign new_n11058_ = new_n5325_ & new_n10111_;
  assign new_n11059_ = ~new_n11057_ & ~new_n11058_;
  assign new_n11060_ = ~new_n11056_ & new_n11059_;
  assign new_n11061_ = new_n11055_ & new_n11060_;
  assign new_n11062_ = new_n5325_ & new_n10116_;
  assign new_n11063_ = new_n5325_ & new_n10118_;
  assign new_n11064_ = new_n5325_ & new_n10120_;
  assign new_n11065_ = ~new_n11063_ & ~new_n11064_;
  assign new_n11066_ = ~new_n11062_ & new_n11065_;
  assign new_n11067_ = new_n5490_ & new_n9926_;
  assign new_n11068_ = new_n5490_ & new_n9928_;
  assign new_n11069_ = ~new_n11067_ & ~new_n11068_;
  assign new_n11070_ = new_n11066_ & new_n11069_;
  assign new_n11071_ = new_n11061_ & new_n11070_;
  assign new_n11072_ = new_n11050_ & new_n11071_;
  assign new_n11073_ = new_n11027_ & new_n11072_;
  assign new_n11074_ = new_n5490_ & new_n9938_;
  assign new_n11075_ = new_n5490_ & new_n9924_;
  assign new_n11076_ = new_n5490_ & new_n9936_;
  assign new_n11077_ = ~new_n11075_ & ~new_n11076_;
  assign new_n11078_ = ~new_n11074_ & new_n11077_;
  assign new_n11079_ = new_n5490_ & new_n9946_;
  assign new_n11080_ = new_n5490_ & new_n9934_;
  assign new_n11081_ = new_n5490_ & new_n9944_;
  assign new_n11082_ = ~new_n11080_ & ~new_n11081_;
  assign new_n11083_ = ~new_n11079_ & new_n11082_;
  assign new_n11084_ = new_n11078_ & new_n11083_;
  assign new_n11085_ = new_n5490_ & new_n9956_;
  assign new_n11086_ = new_n5490_ & new_n9942_;
  assign new_n11087_ = new_n5490_ & new_n9954_;
  assign new_n11088_ = ~new_n11086_ & ~new_n11087_;
  assign new_n11089_ = ~new_n11085_ & new_n11088_;
  assign new_n11090_ = new_n5490_ & new_n9965_;
  assign new_n11091_ = new_n5490_ & new_n9952_;
  assign new_n11092_ = new_n5490_ & new_n9963_;
  assign new_n11093_ = ~new_n11091_ & ~new_n11092_;
  assign new_n11094_ = ~new_n11090_ & new_n11093_;
  assign new_n11095_ = new_n11089_ & new_n11094_;
  assign new_n11096_ = new_n11084_ & new_n11095_;
  assign new_n11097_ = new_n5490_ & new_n9974_;
  assign new_n11098_ = new_n5490_ & new_n9961_;
  assign new_n11099_ = new_n5490_ & new_n9972_;
  assign new_n11100_ = ~new_n11098_ & ~new_n11099_;
  assign new_n11101_ = ~new_n11097_ & new_n11100_;
  assign new_n11102_ = new_n5490_ & new_n9980_;
  assign new_n11103_ = new_n5490_ & new_n9970_;
  assign new_n11104_ = new_n5490_ & new_n9978_;
  assign new_n11105_ = ~new_n11103_ & ~new_n11104_;
  assign new_n11106_ = ~new_n11102_ & new_n11105_;
  assign new_n11107_ = new_n11101_ & new_n11106_;
  assign new_n11108_ = new_n5490_ & new_n9988_;
  assign new_n11109_ = new_n5490_ & new_n9990_;
  assign new_n11110_ = new_n5490_ & new_n9992_;
  assign new_n11111_ = ~new_n11109_ & ~new_n11110_;
  assign new_n11112_ = ~new_n11108_ & new_n11111_;
  assign new_n11113_ = new_n5490_ & new_n9999_;
  assign new_n11114_ = new_n5490_ & new_n10001_;
  assign new_n11115_ = ~new_n11113_ & ~new_n11114_;
  assign new_n11116_ = new_n11112_ & new_n11115_;
  assign new_n11117_ = new_n11107_ & new_n11116_;
  assign new_n11118_ = new_n11096_ & new_n11117_;
  assign new_n11119_ = new_n5490_ & new_n10011_;
  assign new_n11120_ = new_n5490_ & new_n9997_;
  assign new_n11121_ = new_n5490_ & new_n10009_;
  assign new_n11122_ = ~new_n11120_ & ~new_n11121_;
  assign new_n11123_ = ~new_n11119_ & new_n11122_;
  assign new_n11124_ = new_n5490_ & new_n10019_;
  assign new_n11125_ = new_n5490_ & new_n10007_;
  assign new_n11126_ = new_n5490_ & new_n10017_;
  assign new_n11127_ = ~new_n11125_ & ~new_n11126_;
  assign new_n11128_ = ~new_n11124_ & new_n11127_;
  assign new_n11129_ = new_n11123_ & new_n11128_;
  assign new_n11130_ = new_n5490_ & new_n10030_;
  assign new_n11131_ = new_n5490_ & new_n10015_;
  assign new_n11132_ = new_n5490_ & new_n10028_;
  assign new_n11133_ = ~new_n11131_ & ~new_n11132_;
  assign new_n11134_ = ~new_n11130_ & new_n11133_;
  assign new_n11135_ = new_n5490_ & new_n10039_;
  assign new_n11136_ = new_n5490_ & new_n10026_;
  assign new_n11137_ = new_n5490_ & new_n10037_;
  assign new_n11138_ = ~new_n11136_ & ~new_n11137_;
  assign new_n11139_ = ~new_n11135_ & new_n11138_;
  assign new_n11140_ = new_n11134_ & new_n11139_;
  assign new_n11141_ = new_n11129_ & new_n11140_;
  assign new_n11142_ = new_n5490_ & new_n10048_;
  assign new_n11143_ = new_n5490_ & new_n10035_;
  assign new_n11144_ = new_n5490_ & new_n10046_;
  assign new_n11145_ = ~new_n11143_ & ~new_n11144_;
  assign new_n11146_ = ~new_n11142_ & new_n11145_;
  assign new_n11147_ = new_n5490_ & new_n10054_;
  assign new_n11148_ = new_n5490_ & new_n10044_;
  assign new_n11149_ = new_n5490_ & new_n10052_;
  assign new_n11150_ = ~new_n11148_ & ~new_n11149_;
  assign new_n11151_ = ~new_n11147_ & new_n11150_;
  assign new_n11152_ = new_n11146_ & new_n11151_;
  assign new_n11153_ = new_n5490_ & new_n10061_;
  assign new_n11154_ = new_n5490_ & new_n10063_;
  assign new_n11155_ = new_n5490_ & new_n10065_;
  assign new_n11156_ = ~new_n11154_ & ~new_n11155_;
  assign new_n11157_ = ~new_n11153_ & new_n11156_;
  assign new_n11158_ = new_n5490_ & new_n10071_;
  assign new_n11159_ = new_n5490_ & new_n10073_;
  assign new_n11160_ = ~new_n11158_ & ~new_n11159_;
  assign new_n11161_ = new_n11157_ & new_n11160_;
  assign new_n11162_ = new_n11152_ & new_n11161_;
  assign new_n11163_ = new_n11141_ & new_n11162_;
  assign new_n11164_ = new_n11118_ & new_n11163_;
  assign new_n11165_ = new_n11073_ & new_n11164_;
  assign new_n11166_ = new_n10982_ & new_n11165_;
  assign new_n11167_ = new_n5490_ & new_n10082_;
  assign new_n11168_ = new_n5490_ & new_n10069_;
  assign new_n11169_ = new_n5490_ & new_n10080_;
  assign new_n11170_ = ~new_n11168_ & ~new_n11169_;
  assign new_n11171_ = ~new_n11167_ & new_n11170_;
  assign new_n11172_ = new_n5490_ & new_n10091_;
  assign new_n11173_ = new_n5490_ & new_n10078_;
  assign new_n11174_ = new_n5490_ & new_n10089_;
  assign new_n11175_ = ~new_n11173_ & ~new_n11174_;
  assign new_n11176_ = ~new_n11172_ & new_n11175_;
  assign new_n11177_ = new_n11171_ & new_n11176_;
  assign new_n11178_ = new_n5490_ & new_n10102_;
  assign new_n11179_ = new_n5490_ & new_n10087_;
  assign new_n11180_ = new_n5490_ & new_n10100_;
  assign new_n11181_ = ~new_n11179_ & ~new_n11180_;
  assign new_n11182_ = ~new_n11178_ & new_n11181_;
  assign new_n11183_ = new_n5490_ & new_n10111_;
  assign new_n11184_ = new_n5490_ & new_n10098_;
  assign new_n11185_ = new_n5490_ & new_n10109_;
  assign new_n11186_ = ~new_n11184_ & ~new_n11185_;
  assign new_n11187_ = ~new_n11183_ & new_n11186_;
  assign new_n11188_ = new_n11182_ & new_n11187_;
  assign new_n11189_ = new_n11177_ & new_n11188_;
  assign new_n11190_ = new_n5490_ & new_n10120_;
  assign new_n11191_ = new_n5490_ & new_n10107_;
  assign new_n11192_ = new_n5490_ & new_n10118_;
  assign new_n11193_ = ~new_n11191_ & ~new_n11192_;
  assign new_n11194_ = ~new_n11190_ & new_n11193_;
  assign new_n11195_ = new_n5653_ & new_n9928_;
  assign new_n11196_ = new_n5490_ & new_n10116_;
  assign new_n11197_ = new_n5653_ & new_n9926_;
  assign new_n11198_ = ~new_n11196_ & ~new_n11197_;
  assign new_n11199_ = ~new_n11195_ & new_n11198_;
  assign new_n11200_ = new_n11194_ & new_n11199_;
  assign new_n11201_ = new_n5653_ & new_n9938_;
  assign new_n11202_ = new_n5653_ & new_n9924_;
  assign new_n11203_ = new_n5653_ & new_n9936_;
  assign new_n11204_ = ~new_n11202_ & ~new_n11203_;
  assign new_n11205_ = ~new_n11201_ & new_n11204_;
  assign new_n11206_ = new_n5653_ & new_n9934_;
  assign new_n11207_ = new_n5653_ & new_n9944_;
  assign new_n11208_ = ~new_n11206_ & ~new_n11207_;
  assign new_n11209_ = new_n11205_ & new_n11208_;
  assign new_n11210_ = new_n11200_ & new_n11209_;
  assign new_n11211_ = new_n11189_ & new_n11210_;
  assign new_n11212_ = new_n5653_ & new_n9954_;
  assign new_n11213_ = new_n5653_ & new_n9946_;
  assign new_n11214_ = new_n5653_ & new_n9942_;
  assign new_n11215_ = ~new_n11213_ & ~new_n11214_;
  assign new_n11216_ = ~new_n11212_ & new_n11215_;
  assign new_n11217_ = new_n5653_ & new_n9963_;
  assign new_n11218_ = new_n5653_ & new_n9956_;
  assign new_n11219_ = new_n5653_ & new_n9952_;
  assign new_n11220_ = ~new_n11218_ & ~new_n11219_;
  assign new_n11221_ = ~new_n11217_ & new_n11220_;
  assign new_n11222_ = new_n11216_ & new_n11221_;
  assign new_n11223_ = new_n5653_ & new_n9972_;
  assign new_n11224_ = new_n5653_ & new_n9965_;
  assign new_n11225_ = new_n5653_ & new_n9961_;
  assign new_n11226_ = ~new_n11224_ & ~new_n11225_;
  assign new_n11227_ = ~new_n11223_ & new_n11226_;
  assign new_n11228_ = new_n5653_ & new_n9978_;
  assign new_n11229_ = new_n5653_ & new_n9974_;
  assign new_n11230_ = new_n5653_ & new_n9970_;
  assign new_n11231_ = ~new_n11229_ & ~new_n11230_;
  assign new_n11232_ = ~new_n11228_ & new_n11231_;
  assign new_n11233_ = new_n11227_ & new_n11232_;
  assign new_n11234_ = new_n11222_ & new_n11233_;
  assign new_n11235_ = new_n5653_ & new_n9992_;
  assign new_n11236_ = new_n5653_ & new_n9980_;
  assign new_n11237_ = new_n5653_ & new_n9990_;
  assign new_n11238_ = ~new_n11236_ & ~new_n11237_;
  assign new_n11239_ = ~new_n11235_ & new_n11238_;
  assign new_n11240_ = new_n5653_ & new_n10001_;
  assign new_n11241_ = new_n5653_ & new_n9988_;
  assign new_n11242_ = new_n5653_ & new_n9999_;
  assign new_n11243_ = ~new_n11241_ & ~new_n11242_;
  assign new_n11244_ = ~new_n11240_ & new_n11243_;
  assign new_n11245_ = new_n11239_ & new_n11244_;
  assign new_n11246_ = new_n5653_ & new_n10011_;
  assign new_n11247_ = new_n5653_ & new_n9997_;
  assign new_n11248_ = new_n5653_ & new_n10009_;
  assign new_n11249_ = ~new_n11247_ & ~new_n11248_;
  assign new_n11250_ = ~new_n11246_ & new_n11249_;
  assign new_n11251_ = new_n5653_ & new_n10007_;
  assign new_n11252_ = new_n5653_ & new_n10017_;
  assign new_n11253_ = ~new_n11251_ & ~new_n11252_;
  assign new_n11254_ = new_n11250_ & new_n11253_;
  assign new_n11255_ = new_n11245_ & new_n11254_;
  assign new_n11256_ = new_n11234_ & new_n11255_;
  assign new_n11257_ = new_n11211_ & new_n11256_;
  assign new_n11258_ = new_n5653_ & new_n10028_;
  assign new_n11259_ = new_n5653_ & new_n10019_;
  assign new_n11260_ = new_n5653_ & new_n10015_;
  assign new_n11261_ = ~new_n11259_ & ~new_n11260_;
  assign new_n11262_ = ~new_n11258_ & new_n11261_;
  assign new_n11263_ = new_n5653_ & new_n10037_;
  assign new_n11264_ = new_n5653_ & new_n10030_;
  assign new_n11265_ = new_n5653_ & new_n10026_;
  assign new_n11266_ = ~new_n11264_ & ~new_n11265_;
  assign new_n11267_ = ~new_n11263_ & new_n11266_;
  assign new_n11268_ = new_n11262_ & new_n11267_;
  assign new_n11269_ = new_n5653_ & new_n10046_;
  assign new_n11270_ = new_n5653_ & new_n10039_;
  assign new_n11271_ = new_n5653_ & new_n10035_;
  assign new_n11272_ = ~new_n11270_ & ~new_n11271_;
  assign new_n11273_ = ~new_n11269_ & new_n11272_;
  assign new_n11274_ = new_n5653_ & new_n10052_;
  assign new_n11275_ = new_n5653_ & new_n10048_;
  assign new_n11276_ = new_n5653_ & new_n10044_;
  assign new_n11277_ = ~new_n11275_ & ~new_n11276_;
  assign new_n11278_ = ~new_n11274_ & new_n11277_;
  assign new_n11279_ = new_n11273_ & new_n11278_;
  assign new_n11280_ = new_n11268_ & new_n11279_;
  assign new_n11281_ = new_n5653_ & new_n10065_;
  assign new_n11282_ = new_n5653_ & new_n10054_;
  assign new_n11283_ = new_n5653_ & new_n10063_;
  assign new_n11284_ = ~new_n11282_ & ~new_n11283_;
  assign new_n11285_ = ~new_n11281_ & new_n11284_;
  assign new_n11286_ = new_n5653_ & new_n10073_;
  assign new_n11287_ = new_n5653_ & new_n10061_;
  assign new_n11288_ = new_n5653_ & new_n10071_;
  assign new_n11289_ = ~new_n11287_ & ~new_n11288_;
  assign new_n11290_ = ~new_n11286_ & new_n11289_;
  assign new_n11291_ = new_n11285_ & new_n11290_;
  assign new_n11292_ = new_n5653_ & new_n10082_;
  assign new_n11293_ = new_n5653_ & new_n10069_;
  assign new_n11294_ = new_n5653_ & new_n10080_;
  assign new_n11295_ = ~new_n11293_ & ~new_n11294_;
  assign new_n11296_ = ~new_n11292_ & new_n11295_;
  assign new_n11297_ = new_n5653_ & new_n10078_;
  assign new_n11298_ = new_n5653_ & new_n10089_;
  assign new_n11299_ = ~new_n11297_ & ~new_n11298_;
  assign new_n11300_ = new_n11296_ & new_n11299_;
  assign new_n11301_ = new_n11291_ & new_n11300_;
  assign new_n11302_ = new_n11280_ & new_n11301_;
  assign new_n11303_ = new_n5653_ & new_n10100_;
  assign new_n11304_ = new_n5653_ & new_n10091_;
  assign new_n11305_ = new_n5653_ & new_n10087_;
  assign new_n11306_ = ~new_n11304_ & ~new_n11305_;
  assign new_n11307_ = ~new_n11303_ & new_n11306_;
  assign new_n11308_ = new_n5653_ & new_n10109_;
  assign new_n11309_ = new_n5653_ & new_n10102_;
  assign new_n11310_ = new_n5653_ & new_n10098_;
  assign new_n11311_ = ~new_n11309_ & ~new_n11310_;
  assign new_n11312_ = ~new_n11308_ & new_n11311_;
  assign new_n11313_ = new_n11307_ & new_n11312_;
  assign new_n11314_ = new_n5653_ & new_n10118_;
  assign new_n11315_ = new_n5653_ & new_n10111_;
  assign new_n11316_ = new_n5653_ & new_n10107_;
  assign new_n11317_ = ~new_n11315_ & ~new_n11316_;
  assign new_n11318_ = ~new_n11314_ & new_n11317_;
  assign new_n11319_ = new_n5752_ & new_n10127_;
  assign new_n11320_ = new_n10125_ & new_n11319_;
  assign new_n11321_ = new_n5653_ & new_n10120_;
  assign new_n11322_ = new_n5653_ & new_n10116_;
  assign new_n11323_ = ~new_n11321_ & ~new_n11322_;
  assign new_n11324_ = ~new_n11320_ & new_n11323_;
  assign new_n11325_ = new_n11318_ & new_n11324_;
  assign new_n11326_ = new_n11313_ & new_n11325_;
  assign new_n11327_ = new_n5752_ & new_n10147_;
  assign new_n11328_ = new_n10151_ & new_n11327_;
  assign new_n11329_ = new_n5752_ & new_n10132_;
  assign new_n11330_ = new_n10131_ & new_n11329_;
  assign new_n11331_ = new_n10146_ & new_n11327_;
  assign new_n11332_ = ~new_n11330_ & ~new_n11331_;
  assign new_n11333_ = ~new_n11328_ & new_n11332_;
  assign new_n11334_ = new_n5752_ & new_n10155_;
  assign new_n11335_ = new_n10146_ & new_n11334_;
  assign new_n11336_ = new_n5752_ & new_n10142_;
  assign new_n11337_ = new_n10125_ & new_n11336_;
  assign new_n11338_ = new_n5752_ & new_n10158_;
  assign new_n11339_ = new_n10131_ & new_n11338_;
  assign new_n11340_ = ~new_n11337_ & ~new_n11339_;
  assign new_n11341_ = ~new_n11335_ & new_n11340_;
  assign new_n11342_ = new_n11333_ & new_n11341_;
  assign new_n11343_ = new_n5752_ & new_n10172_;
  assign new_n11344_ = new_n10131_ & new_n11343_;
  assign new_n11345_ = new_n10151_ & new_n11334_;
  assign new_n11346_ = new_n5752_ & new_n10169_;
  assign new_n11347_ = new_n10125_ & new_n11346_;
  assign new_n11348_ = ~new_n11345_ & ~new_n11347_;
  assign new_n11349_ = ~new_n11344_ & new_n11348_;
  assign new_n11350_ = new_n5752_ & new_n10166_;
  assign new_n11351_ = new_n10146_ & new_n11350_;
  assign new_n11352_ = new_n10151_ & new_n11350_;
  assign new_n11353_ = ~new_n11351_ & ~new_n11352_;
  assign new_n11354_ = new_n11349_ & new_n11353_;
  assign new_n11355_ = new_n11342_ & new_n11354_;
  assign new_n11356_ = new_n11326_ & new_n11355_;
  assign new_n11357_ = new_n11302_ & new_n11356_;
  assign new_n11358_ = new_n11257_ & new_n11357_;
  assign new_n11359_ = new_n5752_ & new_n10189_;
  assign new_n11360_ = new_n10146_ & new_n11359_;
  assign new_n11361_ = new_n5752_ & new_n10181_;
  assign new_n11362_ = new_n10125_ & new_n11361_;
  assign new_n11363_ = new_n5752_ & new_n10177_;
  assign new_n11364_ = new_n10131_ & new_n11363_;
  assign new_n11365_ = ~new_n11362_ & ~new_n11364_;
  assign new_n11366_ = ~new_n11360_ & new_n11365_;
  assign new_n11367_ = new_n5753_ & new_n8628_;
  assign new_n11368_ = new_n10151_ & new_n11359_;
  assign new_n11369_ = new_n5753_ & new_n8617_;
  assign new_n11370_ = ~new_n11368_ & ~new_n11369_;
  assign new_n11371_ = ~new_n11367_ & new_n11370_;
  assign new_n11372_ = new_n11366_ & new_n11371_;
  assign new_n11373_ = new_n5753_ & new_n8637_;
  assign new_n11374_ = new_n5753_ & new_n8630_;
  assign new_n11375_ = new_n5753_ & new_n8625_;
  assign new_n11376_ = ~new_n11374_ & ~new_n11375_;
  assign new_n11377_ = ~new_n11373_ & new_n11376_;
  assign new_n11378_ = new_n5753_ & new_n8648_;
  assign new_n11379_ = new_n5753_ & new_n8639_;
  assign new_n11380_ = new_n5753_ & new_n8635_;
  assign new_n11381_ = ~new_n11379_ & ~new_n11380_;
  assign new_n11382_ = ~new_n11378_ & new_n11381_;
  assign new_n11383_ = new_n11377_ & new_n11382_;
  assign new_n11384_ = new_n11372_ & new_n11383_;
  assign new_n11385_ = new_n5753_ & new_n8657_;
  assign new_n11386_ = new_n5753_ & new_n8650_;
  assign new_n11387_ = new_n5753_ & new_n8646_;
  assign new_n11388_ = ~new_n11386_ & ~new_n11387_;
  assign new_n11389_ = ~new_n11385_ & new_n11388_;
  assign new_n11390_ = new_n5753_ & new_n8667_;
  assign new_n11391_ = new_n5753_ & new_n8659_;
  assign new_n11392_ = new_n5753_ & new_n8655_;
  assign new_n11393_ = ~new_n11391_ & ~new_n11392_;
  assign new_n11394_ = ~new_n11390_ & new_n11393_;
  assign new_n11395_ = new_n11389_ & new_n11394_;
  assign new_n11396_ = new_n5753_ & new_n8678_;
  assign new_n11397_ = new_n5753_ & new_n8670_;
  assign new_n11398_ = new_n5753_ & new_n8665_;
  assign new_n11399_ = ~new_n11397_ & ~new_n11398_;
  assign new_n11400_ = ~new_n11396_ & new_n11399_;
  assign new_n11401_ = new_n5753_ & new_n8681_;
  assign new_n11402_ = new_n5753_ & new_n8675_;
  assign new_n11403_ = ~new_n11401_ & ~new_n11402_;
  assign new_n11404_ = new_n11400_ & new_n11403_;
  assign new_n11405_ = new_n11395_ & new_n11404_;
  assign new_n11406_ = new_n11384_ & new_n11405_;
  assign new_n11407_ = new_n5753_ & new_n8689_;
  assign new_n11408_ = new_n5753_ & new_n8692_;
  assign new_n11409_ = new_n5753_ & new_n8694_;
  assign new_n11410_ = ~new_n11408_ & ~new_n11409_;
  assign new_n11411_ = ~new_n11407_ & new_n11410_;
  assign new_n11412_ = new_n5759_ & new_n10244_;
  assign new_n11413_ = new_n10125_ & new_n11412_;
  assign new_n11414_ = new_n5753_ & new_n8699_;
  assign new_n11415_ = new_n5753_ & new_n8701_;
  assign new_n11416_ = ~new_n11414_ & ~new_n11415_;
  assign new_n11417_ = ~new_n11413_ & new_n11416_;
  assign new_n11418_ = new_n11411_ & new_n11417_;
  assign new_n11419_ = new_n5759_ & new_n10241_;
  assign new_n11420_ = new_n10151_ & new_n11419_;
  assign new_n11421_ = new_n5759_ & new_n10247_;
  assign new_n11422_ = new_n10131_ & new_n11421_;
  assign new_n11423_ = new_n10146_ & new_n11419_;
  assign new_n11424_ = ~new_n11422_ & ~new_n11423_;
  assign new_n11425_ = ~new_n11420_ & new_n11424_;
  assign new_n11426_ = new_n5759_ & new_n10263_;
  assign new_n11427_ = new_n10146_ & new_n11426_;
  assign new_n11428_ = new_n5759_ & new_n10258_;
  assign new_n11429_ = new_n10125_ & new_n11428_;
  assign new_n11430_ = new_n5759_ & new_n10254_;
  assign new_n11431_ = new_n10131_ & new_n11430_;
  assign new_n11432_ = ~new_n11429_ & ~new_n11431_;
  assign new_n11433_ = ~new_n11427_ & new_n11432_;
  assign new_n11434_ = new_n11425_ & new_n11433_;
  assign new_n11435_ = new_n11418_ & new_n11434_;
  assign new_n11436_ = new_n5759_ & new_n10279_;
  assign new_n11437_ = new_n10131_ & new_n11436_;
  assign new_n11438_ = new_n10151_ & new_n11426_;
  assign new_n11439_ = new_n5759_ & new_n10276_;
  assign new_n11440_ = new_n10125_ & new_n11439_;
  assign new_n11441_ = ~new_n11438_ & ~new_n11440_;
  assign new_n11442_ = ~new_n11437_ & new_n11441_;
  assign new_n11443_ = new_n5759_ & new_n10288_;
  assign new_n11444_ = new_n10125_ & new_n11443_;
  assign new_n11445_ = new_n5759_ & new_n10273_;
  assign new_n11446_ = new_n10146_ & new_n11445_;
  assign new_n11447_ = new_n10151_ & new_n11445_;
  assign new_n11448_ = ~new_n11446_ & ~new_n11447_;
  assign new_n11449_ = ~new_n11444_ & new_n11448_;
  assign new_n11450_ = new_n11442_ & new_n11449_;
  assign new_n11451_ = new_n5759_ & new_n10295_;
  assign new_n11452_ = new_n10151_ & new_n11451_;
  assign new_n11453_ = new_n5759_ & new_n10284_;
  assign new_n11454_ = new_n10131_ & new_n11453_;
  assign new_n11455_ = new_n10146_ & new_n11451_;
  assign new_n11456_ = ~new_n11454_ & ~new_n11455_;
  assign new_n11457_ = ~new_n11452_ & new_n11456_;
  assign new_n11458_ = new_n5760_ & new_n8617_;
  assign new_n11459_ = new_n5760_ & new_n8628_;
  assign new_n11460_ = ~new_n11458_ & ~new_n11459_;
  assign new_n11461_ = new_n11457_ & new_n11460_;
  assign new_n11462_ = new_n11450_ & new_n11461_;
  assign new_n11463_ = new_n11435_ & new_n11462_;
  assign new_n11464_ = new_n11406_ & new_n11463_;
  assign new_n11465_ = new_n5760_ & new_n8637_;
  assign new_n11466_ = new_n5760_ & new_n8630_;
  assign new_n11467_ = new_n5760_ & new_n8625_;
  assign new_n11468_ = ~new_n11466_ & ~new_n11467_;
  assign new_n11469_ = ~new_n11465_ & new_n11468_;
  assign new_n11470_ = new_n5760_ & new_n8648_;
  assign new_n11471_ = new_n5760_ & new_n8639_;
  assign new_n11472_ = new_n5760_ & new_n8635_;
  assign new_n11473_ = ~new_n11471_ & ~new_n11472_;
  assign new_n11474_ = ~new_n11470_ & new_n11473_;
  assign new_n11475_ = new_n11469_ & new_n11474_;
  assign new_n11476_ = new_n5760_ & new_n8657_;
  assign new_n11477_ = new_n5760_ & new_n8650_;
  assign new_n11478_ = new_n5760_ & new_n8646_;
  assign new_n11479_ = ~new_n11477_ & ~new_n11478_;
  assign new_n11480_ = ~new_n11476_ & new_n11479_;
  assign new_n11481_ = new_n5760_ & new_n8667_;
  assign new_n11482_ = new_n5760_ & new_n8659_;
  assign new_n11483_ = new_n5760_ & new_n8655_;
  assign new_n11484_ = ~new_n11482_ & ~new_n11483_;
  assign new_n11485_ = ~new_n11481_ & new_n11484_;
  assign new_n11486_ = new_n11480_ & new_n11485_;
  assign new_n11487_ = new_n11475_ & new_n11486_;
  assign new_n11488_ = new_n5760_ & new_n8678_;
  assign new_n11489_ = new_n5760_ & new_n8670_;
  assign new_n11490_ = new_n5760_ & new_n8665_;
  assign new_n11491_ = ~new_n11489_ & ~new_n11490_;
  assign new_n11492_ = ~new_n11488_ & new_n11491_;
  assign new_n11493_ = new_n5760_ & new_n8692_;
  assign new_n11494_ = new_n5760_ & new_n8681_;
  assign new_n11495_ = new_n5760_ & new_n8675_;
  assign new_n11496_ = ~new_n11494_ & ~new_n11495_;
  assign new_n11497_ = ~new_n11493_ & new_n11496_;
  assign new_n11498_ = new_n11492_ & new_n11497_;
  assign new_n11499_ = new_n5760_ & new_n8699_;
  assign new_n11500_ = new_n5760_ & new_n8694_;
  assign new_n11501_ = new_n5760_ & new_n8689_;
  assign new_n11502_ = ~new_n11500_ & ~new_n11501_;
  assign new_n11503_ = ~new_n11499_ & new_n11502_;
  assign new_n11504_ = new_n5760_ & new_n8701_;
  assign new_n11505_ = new_n5768_ & new_n10349_;
  assign new_n11506_ = new_n10125_ & new_n11505_;
  assign new_n11507_ = ~new_n11504_ & ~new_n11506_;
  assign new_n11508_ = new_n11503_ & new_n11507_;
  assign new_n11509_ = new_n11498_ & new_n11508_;
  assign new_n11510_ = new_n11487_ & new_n11509_;
  assign new_n11511_ = new_n5768_ & new_n10346_;
  assign new_n11512_ = new_n10151_ & new_n11511_;
  assign new_n11513_ = new_n5768_ & new_n10352_;
  assign new_n11514_ = new_n10131_ & new_n11513_;
  assign new_n11515_ = new_n10146_ & new_n11511_;
  assign new_n11516_ = ~new_n11514_ & ~new_n11515_;
  assign new_n11517_ = ~new_n11512_ & new_n11516_;
  assign new_n11518_ = new_n5768_ & new_n10372_;
  assign new_n11519_ = new_n10146_ & new_n11518_;
  assign new_n11520_ = new_n5768_ & new_n10363_;
  assign new_n11521_ = new_n10125_ & new_n11520_;
  assign new_n11522_ = new_n5768_ & new_n10359_;
  assign new_n11523_ = new_n10131_ & new_n11522_;
  assign new_n11524_ = ~new_n11521_ & ~new_n11523_;
  assign new_n11525_ = ~new_n11519_ & new_n11524_;
  assign new_n11526_ = new_n11517_ & new_n11525_;
  assign new_n11527_ = new_n5768_ & new_n10382_;
  assign new_n11528_ = new_n10131_ & new_n11527_;
  assign new_n11529_ = new_n10151_ & new_n11518_;
  assign new_n11530_ = new_n5768_ & new_n10369_;
  assign new_n11531_ = new_n10125_ & new_n11530_;
  assign new_n11532_ = ~new_n11529_ & ~new_n11531_;
  assign new_n11533_ = ~new_n11528_ & new_n11532_;
  assign new_n11534_ = new_n5768_ & new_n10388_;
  assign new_n11535_ = new_n10125_ & new_n11534_;
  assign new_n11536_ = new_n5768_ & new_n10379_;
  assign new_n11537_ = new_n10146_ & new_n11536_;
  assign new_n11538_ = new_n10151_ & new_n11536_;
  assign new_n11539_ = ~new_n11537_ & ~new_n11538_;
  assign new_n11540_ = ~new_n11535_ & new_n11539_;
  assign new_n11541_ = new_n11533_ & new_n11540_;
  assign new_n11542_ = new_n11526_ & new_n11541_;
  assign new_n11543_ = new_n5768_ & new_n10402_;
  assign new_n11544_ = new_n10151_ & new_n11543_;
  assign new_n11545_ = new_n5768_ & new_n10391_;
  assign new_n11546_ = new_n10131_ & new_n11545_;
  assign new_n11547_ = new_n10146_ & new_n11543_;
  assign new_n11548_ = ~new_n11546_ & ~new_n11547_;
  assign new_n11549_ = ~new_n11544_ & new_n11548_;
  assign new_n11550_ = new_n5769_ & new_n8630_;
  assign new_n11551_ = new_n5769_ & new_n8617_;
  assign new_n11552_ = new_n5769_ & new_n8628_;
  assign new_n11553_ = ~new_n11551_ & ~new_n11552_;
  assign new_n11554_ = ~new_n11550_ & new_n11553_;
  assign new_n11555_ = new_n11549_ & new_n11554_;
  assign new_n11556_ = new_n5769_ & new_n8639_;
  assign new_n11557_ = new_n5769_ & new_n8625_;
  assign new_n11558_ = new_n5769_ & new_n8637_;
  assign new_n11559_ = ~new_n11557_ & ~new_n11558_;
  assign new_n11560_ = ~new_n11556_ & new_n11559_;
  assign new_n11561_ = new_n5769_ & new_n8635_;
  assign new_n11562_ = new_n5769_ & new_n8648_;
  assign new_n11563_ = ~new_n11561_ & ~new_n11562_;
  assign new_n11564_ = new_n11560_ & new_n11563_;
  assign new_n11565_ = new_n11555_ & new_n11564_;
  assign new_n11566_ = new_n11542_ & new_n11565_;
  assign new_n11567_ = new_n11510_ & new_n11566_;
  assign new_n11568_ = new_n11464_ & new_n11567_;
  assign new_n11569_ = new_n11358_ & new_n11568_;
  assign new_n11570_ = new_n11166_ & new_n11569_;
  assign new_n11571_ = new_n10797_ & new_n11570_;
  assign new_n11572_ = new_n5769_ & new_n8657_;
  assign new_n11573_ = new_n5769_ & new_n8650_;
  assign new_n11574_ = new_n5769_ & new_n8646_;
  assign new_n11575_ = ~new_n11573_ & ~new_n11574_;
  assign new_n11576_ = ~new_n11572_ & new_n11575_;
  assign new_n11577_ = new_n5769_ & new_n8667_;
  assign new_n11578_ = new_n5769_ & new_n8659_;
  assign new_n11579_ = new_n5769_ & new_n8655_;
  assign new_n11580_ = ~new_n11578_ & ~new_n11579_;
  assign new_n11581_ = ~new_n11577_ & new_n11580_;
  assign new_n11582_ = new_n11576_ & new_n11581_;
  assign new_n11583_ = new_n5769_ & new_n8678_;
  assign new_n11584_ = new_n5769_ & new_n8670_;
  assign new_n11585_ = new_n5769_ & new_n8665_;
  assign new_n11586_ = ~new_n11584_ & ~new_n11585_;
  assign new_n11587_ = ~new_n11583_ & new_n11586_;
  assign new_n11588_ = new_n5769_ & new_n8692_;
  assign new_n11589_ = new_n5769_ & new_n8681_;
  assign new_n11590_ = new_n5769_ & new_n8675_;
  assign new_n11591_ = ~new_n11589_ & ~new_n11590_;
  assign new_n11592_ = ~new_n11588_ & new_n11591_;
  assign new_n11593_ = new_n11587_ & new_n11592_;
  assign new_n11594_ = new_n11582_ & new_n11593_;
  assign new_n11595_ = new_n5769_ & new_n8699_;
  assign new_n11596_ = new_n5769_ & new_n8694_;
  assign new_n11597_ = new_n5769_ & new_n8689_;
  assign new_n11598_ = ~new_n11596_ & ~new_n11597_;
  assign new_n11599_ = ~new_n11595_ & new_n11598_;
  assign new_n11600_ = new_n5768_ & new_n10460_;
  assign new_n11601_ = new_n10131_ & new_n11600_;
  assign new_n11602_ = new_n5769_ & new_n8701_;
  assign new_n11603_ = new_n5768_ & new_n10450_;
  assign new_n11604_ = new_n10125_ & new_n11603_;
  assign new_n11605_ = ~new_n11602_ & ~new_n11604_;
  assign new_n11606_ = ~new_n11601_ & new_n11605_;
  assign new_n11607_ = new_n11599_ & new_n11606_;
  assign new_n11608_ = new_n5768_ & new_n10470_;
  assign new_n11609_ = new_n10125_ & new_n11608_;
  assign new_n11610_ = new_n5768_ & new_n10457_;
  assign new_n11611_ = new_n10146_ & new_n11610_;
  assign new_n11612_ = new_n10151_ & new_n11610_;
  assign new_n11613_ = ~new_n11611_ & ~new_n11612_;
  assign new_n11614_ = ~new_n11609_ & new_n11613_;
  assign new_n11615_ = new_n5768_ & new_n10467_;
  assign new_n11616_ = new_n10151_ & new_n11615_;
  assign new_n11617_ = new_n5768_ & new_n10473_;
  assign new_n11618_ = new_n10131_ & new_n11617_;
  assign new_n11619_ = new_n10146_ & new_n11615_;
  assign new_n11620_ = ~new_n11618_ & ~new_n11619_;
  assign new_n11621_ = ~new_n11616_ & new_n11620_;
  assign new_n11622_ = new_n11614_ & new_n11621_;
  assign new_n11623_ = new_n11607_ & new_n11622_;
  assign new_n11624_ = new_n11594_ & new_n11623_;
  assign new_n11625_ = new_n5768_ & new_n10493_;
  assign new_n11626_ = new_n10146_ & new_n11625_;
  assign new_n11627_ = new_n5768_ & new_n10483_;
  assign new_n11628_ = new_n10125_ & new_n11627_;
  assign new_n11629_ = new_n5768_ & new_n10479_;
  assign new_n11630_ = new_n10131_ & new_n11629_;
  assign new_n11631_ = ~new_n11628_ & ~new_n11630_;
  assign new_n11632_ = ~new_n11626_ & new_n11631_;
  assign new_n11633_ = new_n5768_ & new_n10502_;
  assign new_n11634_ = new_n10131_ & new_n11633_;
  assign new_n11635_ = new_n10151_ & new_n11625_;
  assign new_n11636_ = new_n5768_ & new_n10490_;
  assign new_n11637_ = new_n10125_ & new_n11636_;
  assign new_n11638_ = ~new_n11635_ & ~new_n11637_;
  assign new_n11639_ = ~new_n11634_ & new_n11638_;
  assign new_n11640_ = new_n11632_ & new_n11639_;
  assign new_n11641_ = new_n5781_ & new_n8617_;
  assign new_n11642_ = new_n5768_ & new_n10499_;
  assign new_n11643_ = new_n10146_ & new_n11642_;
  assign new_n11644_ = new_n10151_ & new_n11642_;
  assign new_n11645_ = ~new_n11643_ & ~new_n11644_;
  assign new_n11646_ = ~new_n11641_ & new_n11645_;
  assign new_n11647_ = new_n5781_ & new_n8625_;
  assign new_n11648_ = new_n5781_ & new_n8628_;
  assign new_n11649_ = new_n5781_ & new_n8630_;
  assign new_n11650_ = ~new_n11648_ & ~new_n11649_;
  assign new_n11651_ = ~new_n11647_ & new_n11650_;
  assign new_n11652_ = new_n11646_ & new_n11651_;
  assign new_n11653_ = new_n11640_ & new_n11652_;
  assign new_n11654_ = new_n5781_ & new_n8635_;
  assign new_n11655_ = new_n5781_ & new_n8637_;
  assign new_n11656_ = new_n5781_ & new_n8639_;
  assign new_n11657_ = ~new_n11655_ & ~new_n11656_;
  assign new_n11658_ = ~new_n11654_ & new_n11657_;
  assign new_n11659_ = new_n5781_ & new_n8646_;
  assign new_n11660_ = new_n5781_ & new_n8648_;
  assign new_n11661_ = new_n5781_ & new_n8650_;
  assign new_n11662_ = ~new_n11660_ & ~new_n11661_;
  assign new_n11663_ = ~new_n11659_ & new_n11662_;
  assign new_n11664_ = new_n11658_ & new_n11663_;
  assign new_n11665_ = new_n5781_ & new_n8655_;
  assign new_n11666_ = new_n5781_ & new_n8657_;
  assign new_n11667_ = new_n5781_ & new_n8659_;
  assign new_n11668_ = ~new_n11666_ & ~new_n11667_;
  assign new_n11669_ = ~new_n11665_ & new_n11668_;
  assign new_n11670_ = new_n5781_ & new_n8667_;
  assign new_n11671_ = new_n5781_ & new_n8670_;
  assign new_n11672_ = ~new_n11670_ & ~new_n11671_;
  assign new_n11673_ = new_n11669_ & new_n11672_;
  assign new_n11674_ = new_n11664_ & new_n11673_;
  assign new_n11675_ = new_n11653_ & new_n11674_;
  assign new_n11676_ = new_n11624_ & new_n11675_;
  assign new_n11677_ = new_n5781_ & new_n8681_;
  assign new_n11678_ = new_n5781_ & new_n8665_;
  assign new_n11679_ = new_n5781_ & new_n8678_;
  assign new_n11680_ = ~new_n11678_ & ~new_n11679_;
  assign new_n11681_ = ~new_n11677_ & new_n11680_;
  assign new_n11682_ = new_n5781_ & new_n8694_;
  assign new_n11683_ = new_n5781_ & new_n8675_;
  assign new_n11684_ = new_n5781_ & new_n8692_;
  assign new_n11685_ = ~new_n11683_ & ~new_n11684_;
  assign new_n11686_ = ~new_n11682_ & new_n11685_;
  assign new_n11687_ = new_n11681_ & new_n11686_;
  assign new_n11688_ = new_n5781_ & new_n8701_;
  assign new_n11689_ = new_n5781_ & new_n8689_;
  assign new_n11690_ = new_n5781_ & new_n8699_;
  assign new_n11691_ = ~new_n11689_ & ~new_n11690_;
  assign new_n11692_ = ~new_n11688_ & new_n11691_;
  assign new_n11693_ = new_n5789_ & new_n8630_;
  assign new_n11694_ = new_n5789_ & new_n8617_;
  assign new_n11695_ = new_n5789_ & new_n8628_;
  assign new_n11696_ = ~new_n11694_ & ~new_n11695_;
  assign new_n11697_ = ~new_n11693_ & new_n11696_;
  assign new_n11698_ = new_n11692_ & new_n11697_;
  assign new_n11699_ = new_n11687_ & new_n11698_;
  assign new_n11700_ = new_n5789_ & new_n8639_;
  assign new_n11701_ = new_n5789_ & new_n8625_;
  assign new_n11702_ = new_n5789_ & new_n8637_;
  assign new_n11703_ = ~new_n11701_ & ~new_n11702_;
  assign new_n11704_ = ~new_n11700_ & new_n11703_;
  assign new_n11705_ = new_n5789_ & new_n8650_;
  assign new_n11706_ = new_n5789_ & new_n8635_;
  assign new_n11707_ = new_n5789_ & new_n8648_;
  assign new_n11708_ = ~new_n11706_ & ~new_n11707_;
  assign new_n11709_ = ~new_n11705_ & new_n11708_;
  assign new_n11710_ = new_n11704_ & new_n11709_;
  assign new_n11711_ = new_n5789_ & new_n8659_;
  assign new_n11712_ = new_n5789_ & new_n8646_;
  assign new_n11713_ = new_n5789_ & new_n8657_;
  assign new_n11714_ = ~new_n11712_ & ~new_n11713_;
  assign new_n11715_ = ~new_n11711_ & new_n11714_;
  assign new_n11716_ = new_n5789_ & new_n8655_;
  assign new_n11717_ = new_n5789_ & new_n8667_;
  assign new_n11718_ = ~new_n11716_ & ~new_n11717_;
  assign new_n11719_ = new_n11715_ & new_n11718_;
  assign new_n11720_ = new_n11710_ & new_n11719_;
  assign new_n11721_ = new_n11699_ & new_n11720_;
  assign new_n11722_ = new_n5789_ & new_n8678_;
  assign new_n11723_ = new_n5789_ & new_n8670_;
  assign new_n11724_ = new_n5789_ & new_n8665_;
  assign new_n11725_ = ~new_n11723_ & ~new_n11724_;
  assign new_n11726_ = ~new_n11722_ & new_n11725_;
  assign new_n11727_ = new_n5789_ & new_n8692_;
  assign new_n11728_ = new_n5789_ & new_n8681_;
  assign new_n11729_ = new_n5789_ & new_n8675_;
  assign new_n11730_ = ~new_n11728_ & ~new_n11729_;
  assign new_n11731_ = ~new_n11727_ & new_n11730_;
  assign new_n11732_ = new_n11726_ & new_n11731_;
  assign new_n11733_ = new_n5789_ & new_n8699_;
  assign new_n11734_ = new_n5789_ & new_n8694_;
  assign new_n11735_ = new_n5789_ & new_n8689_;
  assign new_n11736_ = ~new_n11734_ & ~new_n11735_;
  assign new_n11737_ = ~new_n11733_ & new_n11736_;
  assign new_n11738_ = new_n5800_ & new_n8628_;
  assign new_n11739_ = new_n5789_ & new_n8701_;
  assign new_n11740_ = new_n5800_ & new_n8617_;
  assign new_n11741_ = ~new_n11739_ & ~new_n11740_;
  assign new_n11742_ = ~new_n11738_ & new_n11741_;
  assign new_n11743_ = new_n11737_ & new_n11742_;
  assign new_n11744_ = new_n11732_ & new_n11743_;
  assign new_n11745_ = new_n5800_ & new_n8637_;
  assign new_n11746_ = new_n5800_ & new_n8630_;
  assign new_n11747_ = new_n5800_ & new_n8625_;
  assign new_n11748_ = ~new_n11746_ & ~new_n11747_;
  assign new_n11749_ = ~new_n11745_ & new_n11748_;
  assign new_n11750_ = new_n5800_ & new_n8648_;
  assign new_n11751_ = new_n5800_ & new_n8639_;
  assign new_n11752_ = new_n5800_ & new_n8635_;
  assign new_n11753_ = ~new_n11751_ & ~new_n11752_;
  assign new_n11754_ = ~new_n11750_ & new_n11753_;
  assign new_n11755_ = new_n11749_ & new_n11754_;
  assign new_n11756_ = new_n5800_ & new_n8657_;
  assign new_n11757_ = new_n5800_ & new_n8650_;
  assign new_n11758_ = new_n5800_ & new_n8646_;
  assign new_n11759_ = ~new_n11757_ & ~new_n11758_;
  assign new_n11760_ = ~new_n11756_ & new_n11759_;
  assign new_n11761_ = new_n5800_ & new_n8659_;
  assign new_n11762_ = new_n5800_ & new_n8655_;
  assign new_n11763_ = ~new_n11761_ & ~new_n11762_;
  assign new_n11764_ = new_n11760_ & new_n11763_;
  assign new_n11765_ = new_n11755_ & new_n11764_;
  assign new_n11766_ = new_n11744_ & new_n11765_;
  assign new_n11767_ = new_n11721_ & new_n11766_;
  assign new_n11768_ = new_n11676_ & new_n11767_;
  assign new_n11769_ = new_n5800_ & new_n8665_;
  assign new_n11770_ = new_n5800_ & new_n8667_;
  assign new_n11771_ = new_n5800_ & new_n8670_;
  assign new_n11772_ = ~new_n11770_ & ~new_n11771_;
  assign new_n11773_ = ~new_n11769_ & new_n11772_;
  assign new_n11774_ = new_n5800_ & new_n8675_;
  assign new_n11775_ = new_n5800_ & new_n8678_;
  assign new_n11776_ = new_n5800_ & new_n8681_;
  assign new_n11777_ = ~new_n11775_ & ~new_n11776_;
  assign new_n11778_ = ~new_n11774_ & new_n11777_;
  assign new_n11779_ = new_n11773_ & new_n11778_;
  assign new_n11780_ = new_n5800_ & new_n8689_;
  assign new_n11781_ = new_n5800_ & new_n8692_;
  assign new_n11782_ = new_n5800_ & new_n8694_;
  assign new_n11783_ = ~new_n11781_ & ~new_n11782_;
  assign new_n11784_ = ~new_n11780_ & new_n11783_;
  assign new_n11785_ = new_n5807_ & new_n8617_;
  assign new_n11786_ = new_n5800_ & new_n8699_;
  assign new_n11787_ = new_n5800_ & new_n8701_;
  assign new_n11788_ = ~new_n11786_ & ~new_n11787_;
  assign new_n11789_ = ~new_n11785_ & new_n11788_;
  assign new_n11790_ = new_n11784_ & new_n11789_;
  assign new_n11791_ = new_n11779_ & new_n11790_;
  assign new_n11792_ = new_n5807_ & new_n8625_;
  assign new_n11793_ = new_n5807_ & new_n8628_;
  assign new_n11794_ = new_n5807_ & new_n8630_;
  assign new_n11795_ = ~new_n11793_ & ~new_n11794_;
  assign new_n11796_ = ~new_n11792_ & new_n11795_;
  assign new_n11797_ = new_n5807_ & new_n8635_;
  assign new_n11798_ = new_n5807_ & new_n8637_;
  assign new_n11799_ = new_n5807_ & new_n8639_;
  assign new_n11800_ = ~new_n11798_ & ~new_n11799_;
  assign new_n11801_ = ~new_n11797_ & new_n11800_;
  assign new_n11802_ = new_n11796_ & new_n11801_;
  assign new_n11803_ = new_n5807_ & new_n8646_;
  assign new_n11804_ = new_n5807_ & new_n8648_;
  assign new_n11805_ = new_n5807_ & new_n8650_;
  assign new_n11806_ = ~new_n11804_ & ~new_n11805_;
  assign new_n11807_ = ~new_n11803_ & new_n11806_;
  assign new_n11808_ = new_n5807_ & new_n8657_;
  assign new_n11809_ = new_n5807_ & new_n8659_;
  assign new_n11810_ = ~new_n11808_ & ~new_n11809_;
  assign new_n11811_ = new_n11807_ & new_n11810_;
  assign new_n11812_ = new_n11802_ & new_n11811_;
  assign new_n11813_ = new_n11791_ & new_n11812_;
  assign new_n11814_ = new_n5807_ & new_n8670_;
  assign new_n11815_ = new_n5807_ & new_n8655_;
  assign new_n11816_ = new_n5807_ & new_n8667_;
  assign new_n11817_ = ~new_n11815_ & ~new_n11816_;
  assign new_n11818_ = ~new_n11814_ & new_n11817_;
  assign new_n11819_ = new_n5807_ & new_n8681_;
  assign new_n11820_ = new_n5807_ & new_n8665_;
  assign new_n11821_ = new_n5807_ & new_n8678_;
  assign new_n11822_ = ~new_n11820_ & ~new_n11821_;
  assign new_n11823_ = ~new_n11819_ & new_n11822_;
  assign new_n11824_ = new_n11818_ & new_n11823_;
  assign new_n11825_ = new_n5807_ & new_n8694_;
  assign new_n11826_ = new_n5807_ & new_n8675_;
  assign new_n11827_ = new_n5807_ & new_n8692_;
  assign new_n11828_ = ~new_n11826_ & ~new_n11827_;
  assign new_n11829_ = ~new_n11825_ & new_n11828_;
  assign new_n11830_ = new_n5807_ & new_n8701_;
  assign new_n11831_ = new_n5807_ & new_n8689_;
  assign new_n11832_ = new_n5807_ & new_n8699_;
  assign new_n11833_ = ~new_n11831_ & ~new_n11832_;
  assign new_n11834_ = ~new_n11830_ & new_n11833_;
  assign new_n11835_ = new_n11829_ & new_n11834_;
  assign new_n11836_ = new_n11824_ & new_n11835_;
  assign new_n11837_ = new_n5813_ & new_n8630_;
  assign new_n11838_ = new_n5813_ & new_n8617_;
  assign new_n11839_ = new_n5813_ & new_n8628_;
  assign new_n11840_ = ~new_n11838_ & ~new_n11839_;
  assign new_n11841_ = ~new_n11837_ & new_n11840_;
  assign new_n11842_ = new_n5813_ & new_n8639_;
  assign new_n11843_ = new_n5813_ & new_n8625_;
  assign new_n11844_ = new_n5813_ & new_n8637_;
  assign new_n11845_ = ~new_n11843_ & ~new_n11844_;
  assign new_n11846_ = ~new_n11842_ & new_n11845_;
  assign new_n11847_ = new_n11841_ & new_n11846_;
  assign new_n11848_ = new_n5813_ & new_n8650_;
  assign new_n11849_ = new_n5813_ & new_n8635_;
  assign new_n11850_ = new_n5813_ & new_n8648_;
  assign new_n11851_ = ~new_n11849_ & ~new_n11850_;
  assign new_n11852_ = ~new_n11848_ & new_n11851_;
  assign new_n11853_ = new_n5813_ & new_n8646_;
  assign new_n11854_ = new_n5813_ & new_n8657_;
  assign new_n11855_ = ~new_n11853_ & ~new_n11854_;
  assign new_n11856_ = new_n11852_ & new_n11855_;
  assign new_n11857_ = new_n11847_ & new_n11856_;
  assign new_n11858_ = new_n11836_ & new_n11857_;
  assign new_n11859_ = new_n11813_ & new_n11858_;
  assign new_n11860_ = new_n5813_ & new_n8667_;
  assign new_n11861_ = new_n5813_ & new_n8659_;
  assign new_n11862_ = new_n5813_ & new_n8655_;
  assign new_n11863_ = ~new_n11861_ & ~new_n11862_;
  assign new_n11864_ = ~new_n11860_ & new_n11863_;
  assign new_n11865_ = new_n5813_ & new_n8678_;
  assign new_n11866_ = new_n5813_ & new_n8670_;
  assign new_n11867_ = new_n5813_ & new_n8665_;
  assign new_n11868_ = ~new_n11866_ & ~new_n11867_;
  assign new_n11869_ = ~new_n11865_ & new_n11868_;
  assign new_n11870_ = new_n11864_ & new_n11869_;
  assign new_n11871_ = new_n5813_ & new_n8692_;
  assign new_n11872_ = new_n5813_ & new_n8681_;
  assign new_n11873_ = new_n5813_ & new_n8675_;
  assign new_n11874_ = ~new_n11872_ & ~new_n11873_;
  assign new_n11875_ = ~new_n11871_ & new_n11874_;
  assign new_n11876_ = new_n5813_ & new_n8699_;
  assign new_n11877_ = new_n5813_ & new_n8694_;
  assign new_n11878_ = new_n5813_ & new_n8689_;
  assign new_n11879_ = ~new_n11877_ & ~new_n11878_;
  assign new_n11880_ = ~new_n11876_ & new_n11879_;
  assign new_n11881_ = new_n11875_ & new_n11880_;
  assign new_n11882_ = new_n11870_ & new_n11881_;
  assign new_n11883_ = new_n5826_ & new_n8853_;
  assign new_n11884_ = new_n5813_ & new_n8701_;
  assign new_n11885_ = new_n5826_ & new_n8845_;
  assign new_n11886_ = ~new_n11884_ & ~new_n11885_;
  assign new_n11887_ = ~new_n11883_ & new_n11886_;
  assign new_n11888_ = new_n5826_ & new_n8864_;
  assign new_n11889_ = new_n5826_ & new_n8855_;
  assign new_n11890_ = new_n5826_ & new_n8851_;
  assign new_n11891_ = ~new_n11889_ & ~new_n11890_;
  assign new_n11892_ = ~new_n11888_ & new_n11891_;
  assign new_n11893_ = new_n11887_ & new_n11892_;
  assign new_n11894_ = new_n5826_ & new_n8872_;
  assign new_n11895_ = new_n5826_ & new_n8866_;
  assign new_n11896_ = new_n5826_ & new_n8862_;
  assign new_n11897_ = ~new_n11895_ & ~new_n11896_;
  assign new_n11898_ = ~new_n11894_ & new_n11897_;
  assign new_n11899_ = new_n5826_ & new_n8874_;
  assign new_n11900_ = new_n5826_ & new_n8870_;
  assign new_n11901_ = ~new_n11899_ & ~new_n11900_;
  assign new_n11902_ = new_n11898_ & new_n11901_;
  assign new_n11903_ = new_n11893_ & new_n11902_;
  assign new_n11904_ = new_n11882_ & new_n11903_;
  assign new_n11905_ = new_n5826_ & new_n8880_;
  assign new_n11906_ = new_n5826_ & new_n8882_;
  assign new_n11907_ = new_n5826_ & new_n8884_;
  assign new_n11908_ = ~new_n11906_ & ~new_n11907_;
  assign new_n11909_ = ~new_n11905_ & new_n11908_;
  assign new_n11910_ = new_n5826_ & new_n8898_;
  assign new_n11911_ = new_n5826_ & new_n8888_;
  assign new_n11912_ = new_n5826_ & new_n8890_;
  assign new_n11913_ = ~new_n11911_ & ~new_n11912_;
  assign new_n11914_ = ~new_n11910_ & new_n11913_;
  assign new_n11915_ = new_n11909_ & new_n11914_;
  assign new_n11916_ = new_n5826_ & new_n8907_;
  assign new_n11917_ = new_n5826_ & new_n8900_;
  assign new_n11918_ = new_n5826_ & new_n8896_;
  assign new_n11919_ = ~new_n11917_ & ~new_n11918_;
  assign new_n11920_ = ~new_n11916_ & new_n11919_;
  assign new_n11921_ = new_n5826_ & new_n8916_;
  assign new_n11922_ = new_n5826_ & new_n8909_;
  assign new_n11923_ = new_n5826_ & new_n8905_;
  assign new_n11924_ = ~new_n11922_ & ~new_n11923_;
  assign new_n11925_ = ~new_n11921_ & new_n11924_;
  assign new_n11926_ = new_n11920_ & new_n11925_;
  assign new_n11927_ = new_n11915_ & new_n11926_;
  assign new_n11928_ = new_n5826_ & new_n8925_;
  assign new_n11929_ = new_n5826_ & new_n8918_;
  assign new_n11930_ = new_n5826_ & new_n8914_;
  assign new_n11931_ = ~new_n11929_ & ~new_n11930_;
  assign new_n11932_ = ~new_n11928_ & new_n11931_;
  assign new_n11933_ = new_n5826_ & new_n8936_;
  assign new_n11934_ = new_n5826_ & new_n8927_;
  assign new_n11935_ = new_n5826_ & new_n8923_;
  assign new_n11936_ = ~new_n11934_ & ~new_n11935_;
  assign new_n11937_ = ~new_n11933_ & new_n11936_;
  assign new_n11938_ = new_n11932_ & new_n11937_;
  assign new_n11939_ = new_n5826_ & new_n8943_;
  assign new_n11940_ = new_n5826_ & new_n8938_;
  assign new_n11941_ = new_n5826_ & new_n8934_;
  assign new_n11942_ = ~new_n11940_ & ~new_n11941_;
  assign new_n11943_ = ~new_n11939_ & new_n11942_;
  assign new_n11944_ = new_n5826_ & new_n8945_;
  assign new_n11945_ = new_n5941_ & new_n9926_;
  assign new_n11946_ = ~new_n11944_ & ~new_n11945_;
  assign new_n11947_ = new_n11943_ & new_n11946_;
  assign new_n11948_ = new_n11938_ & new_n11947_;
  assign new_n11949_ = new_n11927_ & new_n11948_;
  assign new_n11950_ = new_n11904_ & new_n11949_;
  assign new_n11951_ = new_n11859_ & new_n11950_;
  assign new_n11952_ = new_n11768_ & new_n11951_;
  assign new_n11953_ = new_n5941_ & new_n9936_;
  assign new_n11954_ = new_n5941_ & new_n9928_;
  assign new_n11955_ = new_n5941_ & new_n9924_;
  assign new_n11956_ = ~new_n11954_ & ~new_n11955_;
  assign new_n11957_ = ~new_n11953_ & new_n11956_;
  assign new_n11958_ = new_n5941_ & new_n9944_;
  assign new_n11959_ = new_n5941_ & new_n9938_;
  assign new_n11960_ = new_n5941_ & new_n9934_;
  assign new_n11961_ = ~new_n11959_ & ~new_n11960_;
  assign new_n11962_ = ~new_n11958_ & new_n11961_;
  assign new_n11963_ = new_n11957_ & new_n11962_;
  assign new_n11964_ = new_n5941_ & new_n9954_;
  assign new_n11965_ = new_n5941_ & new_n9946_;
  assign new_n11966_ = new_n5941_ & new_n9942_;
  assign new_n11967_ = ~new_n11965_ & ~new_n11966_;
  assign new_n11968_ = ~new_n11964_ & new_n11967_;
  assign new_n11969_ = new_n5941_ & new_n9963_;
  assign new_n11970_ = new_n5941_ & new_n9956_;
  assign new_n11971_ = new_n5941_ & new_n9952_;
  assign new_n11972_ = ~new_n11970_ & ~new_n11971_;
  assign new_n11973_ = ~new_n11969_ & new_n11972_;
  assign new_n11974_ = new_n11968_ & new_n11973_;
  assign new_n11975_ = new_n11963_ & new_n11974_;
  assign new_n11976_ = new_n5941_ & new_n9972_;
  assign new_n11977_ = new_n5941_ & new_n9965_;
  assign new_n11978_ = new_n5941_ & new_n9961_;
  assign new_n11979_ = ~new_n11977_ & ~new_n11978_;
  assign new_n11980_ = ~new_n11976_ & new_n11979_;
  assign new_n11981_ = new_n5941_ & new_n9978_;
  assign new_n11982_ = new_n5941_ & new_n9974_;
  assign new_n11983_ = new_n5941_ & new_n9970_;
  assign new_n11984_ = ~new_n11982_ & ~new_n11983_;
  assign new_n11985_ = ~new_n11981_ & new_n11984_;
  assign new_n11986_ = new_n11980_ & new_n11985_;
  assign new_n11987_ = new_n5941_ & new_n9992_;
  assign new_n11988_ = new_n5941_ & new_n9980_;
  assign new_n11989_ = new_n5941_ & new_n9990_;
  assign new_n11990_ = ~new_n11988_ & ~new_n11989_;
  assign new_n11991_ = ~new_n11987_ & new_n11990_;
  assign new_n11992_ = new_n5941_ & new_n9988_;
  assign new_n11993_ = new_n5941_ & new_n9999_;
  assign new_n11994_ = ~new_n11992_ & ~new_n11993_;
  assign new_n11995_ = new_n11991_ & new_n11994_;
  assign new_n11996_ = new_n11986_ & new_n11995_;
  assign new_n11997_ = new_n11975_ & new_n11996_;
  assign new_n11998_ = new_n5941_ & new_n10009_;
  assign new_n11999_ = new_n5941_ & new_n10001_;
  assign new_n12000_ = new_n5941_ & new_n9997_;
  assign new_n12001_ = ~new_n11999_ & ~new_n12000_;
  assign new_n12002_ = ~new_n11998_ & new_n12001_;
  assign new_n12003_ = new_n5941_ & new_n10017_;
  assign new_n12004_ = new_n5941_ & new_n10011_;
  assign new_n12005_ = new_n5941_ & new_n10007_;
  assign new_n12006_ = ~new_n12004_ & ~new_n12005_;
  assign new_n12007_ = ~new_n12003_ & new_n12006_;
  assign new_n12008_ = new_n12002_ & new_n12007_;
  assign new_n12009_ = new_n5941_ & new_n10028_;
  assign new_n12010_ = new_n5941_ & new_n10019_;
  assign new_n12011_ = new_n5941_ & new_n10015_;
  assign new_n12012_ = ~new_n12010_ & ~new_n12011_;
  assign new_n12013_ = ~new_n12009_ & new_n12012_;
  assign new_n12014_ = new_n5941_ & new_n10037_;
  assign new_n12015_ = new_n5941_ & new_n10030_;
  assign new_n12016_ = new_n5941_ & new_n10026_;
  assign new_n12017_ = ~new_n12015_ & ~new_n12016_;
  assign new_n12018_ = ~new_n12014_ & new_n12017_;
  assign new_n12019_ = new_n12013_ & new_n12018_;
  assign new_n12020_ = new_n12008_ & new_n12019_;
  assign new_n12021_ = new_n5941_ & new_n10046_;
  assign new_n12022_ = new_n5941_ & new_n10039_;
  assign new_n12023_ = new_n5941_ & new_n10035_;
  assign new_n12024_ = ~new_n12022_ & ~new_n12023_;
  assign new_n12025_ = ~new_n12021_ & new_n12024_;
  assign new_n12026_ = new_n5941_ & new_n10052_;
  assign new_n12027_ = new_n5941_ & new_n10048_;
  assign new_n12028_ = new_n5941_ & new_n10044_;
  assign new_n12029_ = ~new_n12027_ & ~new_n12028_;
  assign new_n12030_ = ~new_n12026_ & new_n12029_;
  assign new_n12031_ = new_n12025_ & new_n12030_;
  assign new_n12032_ = new_n5941_ & new_n10065_;
  assign new_n12033_ = new_n5941_ & new_n10054_;
  assign new_n12034_ = new_n5941_ & new_n10063_;
  assign new_n12035_ = ~new_n12033_ & ~new_n12034_;
  assign new_n12036_ = ~new_n12032_ & new_n12035_;
  assign new_n12037_ = new_n5941_ & new_n10061_;
  assign new_n12038_ = new_n5941_ & new_n10071_;
  assign new_n12039_ = ~new_n12037_ & ~new_n12038_;
  assign new_n12040_ = new_n12036_ & new_n12039_;
  assign new_n12041_ = new_n12031_ & new_n12040_;
  assign new_n12042_ = new_n12020_ & new_n12041_;
  assign new_n12043_ = new_n11997_ & new_n12042_;
  assign new_n12044_ = new_n5941_ & new_n10080_;
  assign new_n12045_ = new_n5941_ & new_n10073_;
  assign new_n12046_ = new_n5941_ & new_n10069_;
  assign new_n12047_ = ~new_n12045_ & ~new_n12046_;
  assign new_n12048_ = ~new_n12044_ & new_n12047_;
  assign new_n12049_ = new_n5941_ & new_n10089_;
  assign new_n12050_ = new_n5941_ & new_n10082_;
  assign new_n12051_ = new_n5941_ & new_n10078_;
  assign new_n12052_ = ~new_n12050_ & ~new_n12051_;
  assign new_n12053_ = ~new_n12049_ & new_n12052_;
  assign new_n12054_ = new_n12048_ & new_n12053_;
  assign new_n12055_ = new_n5941_ & new_n10100_;
  assign new_n12056_ = new_n5941_ & new_n10091_;
  assign new_n12057_ = new_n5941_ & new_n10087_;
  assign new_n12058_ = ~new_n12056_ & ~new_n12057_;
  assign new_n12059_ = ~new_n12055_ & new_n12058_;
  assign new_n12060_ = new_n5941_ & new_n10109_;
  assign new_n12061_ = new_n5941_ & new_n10102_;
  assign new_n12062_ = new_n5941_ & new_n10098_;
  assign new_n12063_ = ~new_n12061_ & ~new_n12062_;
  assign new_n12064_ = ~new_n12060_ & new_n12063_;
  assign new_n12065_ = new_n12059_ & new_n12064_;
  assign new_n12066_ = new_n12054_ & new_n12065_;
  assign new_n12067_ = new_n5941_ & new_n10118_;
  assign new_n12068_ = new_n5941_ & new_n10111_;
  assign new_n12069_ = new_n5941_ & new_n10107_;
  assign new_n12070_ = ~new_n12068_ & ~new_n12069_;
  assign new_n12071_ = ~new_n12067_ & new_n12070_;
  assign new_n12072_ = new_n6104_ & new_n9926_;
  assign new_n12073_ = new_n5941_ & new_n10120_;
  assign new_n12074_ = new_n5941_ & new_n10116_;
  assign new_n12075_ = ~new_n12073_ & ~new_n12074_;
  assign new_n12076_ = ~new_n12072_ & new_n12075_;
  assign new_n12077_ = new_n12071_ & new_n12076_;
  assign new_n12078_ = new_n6104_ & new_n9936_;
  assign new_n12079_ = new_n6104_ & new_n9928_;
  assign new_n12080_ = new_n6104_ & new_n9924_;
  assign new_n12081_ = ~new_n12079_ & ~new_n12080_;
  assign new_n12082_ = ~new_n12078_ & new_n12081_;
  assign new_n12083_ = new_n6104_ & new_n9938_;
  assign new_n12084_ = new_n6104_ & new_n9934_;
  assign new_n12085_ = ~new_n12083_ & ~new_n12084_;
  assign new_n12086_ = new_n12082_ & new_n12085_;
  assign new_n12087_ = new_n12077_ & new_n12086_;
  assign new_n12088_ = new_n12066_ & new_n12087_;
  assign new_n12089_ = new_n6104_ & new_n9942_;
  assign new_n12090_ = new_n6104_ & new_n9944_;
  assign new_n12091_ = new_n6104_ & new_n9946_;
  assign new_n12092_ = ~new_n12090_ & ~new_n12091_;
  assign new_n12093_ = ~new_n12089_ & new_n12092_;
  assign new_n12094_ = new_n6104_ & new_n9952_;
  assign new_n12095_ = new_n6104_ & new_n9954_;
  assign new_n12096_ = new_n6104_ & new_n9956_;
  assign new_n12097_ = ~new_n12095_ & ~new_n12096_;
  assign new_n12098_ = ~new_n12094_ & new_n12097_;
  assign new_n12099_ = new_n12093_ & new_n12098_;
  assign new_n12100_ = new_n6104_ & new_n9961_;
  assign new_n12101_ = new_n6104_ & new_n9963_;
  assign new_n12102_ = new_n6104_ & new_n9965_;
  assign new_n12103_ = ~new_n12101_ & ~new_n12102_;
  assign new_n12104_ = ~new_n12100_ & new_n12103_;
  assign new_n12105_ = new_n6104_ & new_n9970_;
  assign new_n12106_ = new_n6104_ & new_n9972_;
  assign new_n12107_ = new_n6104_ & new_n9974_;
  assign new_n12108_ = ~new_n12106_ & ~new_n12107_;
  assign new_n12109_ = ~new_n12105_ & new_n12108_;
  assign new_n12110_ = new_n12104_ & new_n12109_;
  assign new_n12111_ = new_n12099_ & new_n12110_;
  assign new_n12112_ = new_n6104_ & new_n9990_;
  assign new_n12113_ = new_n6104_ & new_n9978_;
  assign new_n12114_ = new_n6104_ & new_n9980_;
  assign new_n12115_ = ~new_n12113_ & ~new_n12114_;
  assign new_n12116_ = ~new_n12112_ & new_n12115_;
  assign new_n12117_ = new_n6104_ & new_n9999_;
  assign new_n12118_ = new_n6104_ & new_n9992_;
  assign new_n12119_ = new_n6104_ & new_n9988_;
  assign new_n12120_ = ~new_n12118_ & ~new_n12119_;
  assign new_n12121_ = ~new_n12117_ & new_n12120_;
  assign new_n12122_ = new_n12116_ & new_n12121_;
  assign new_n12123_ = new_n6104_ & new_n10009_;
  assign new_n12124_ = new_n6104_ & new_n10001_;
  assign new_n12125_ = new_n6104_ & new_n9997_;
  assign new_n12126_ = ~new_n12124_ & ~new_n12125_;
  assign new_n12127_ = ~new_n12123_ & new_n12126_;
  assign new_n12128_ = new_n6104_ & new_n10011_;
  assign new_n12129_ = new_n6104_ & new_n10007_;
  assign new_n12130_ = ~new_n12128_ & ~new_n12129_;
  assign new_n12131_ = new_n12127_ & new_n12130_;
  assign new_n12132_ = new_n12122_ & new_n12131_;
  assign new_n12133_ = new_n12111_ & new_n12132_;
  assign new_n12134_ = new_n12088_ & new_n12133_;
  assign new_n12135_ = new_n12043_ & new_n12134_;
  assign new_n12136_ = new_n6104_ & new_n10015_;
  assign new_n12137_ = new_n6104_ & new_n10017_;
  assign new_n12138_ = new_n6104_ & new_n10019_;
  assign new_n12139_ = ~new_n12137_ & ~new_n12138_;
  assign new_n12140_ = ~new_n12136_ & new_n12139_;
  assign new_n12141_ = new_n6104_ & new_n10026_;
  assign new_n12142_ = new_n6104_ & new_n10028_;
  assign new_n12143_ = new_n6104_ & new_n10030_;
  assign new_n12144_ = ~new_n12142_ & ~new_n12143_;
  assign new_n12145_ = ~new_n12141_ & new_n12144_;
  assign new_n12146_ = new_n12140_ & new_n12145_;
  assign new_n12147_ = new_n6104_ & new_n10035_;
  assign new_n12148_ = new_n6104_ & new_n10037_;
  assign new_n12149_ = new_n6104_ & new_n10039_;
  assign new_n12150_ = ~new_n12148_ & ~new_n12149_;
  assign new_n12151_ = ~new_n12147_ & new_n12150_;
  assign new_n12152_ = new_n6104_ & new_n10044_;
  assign new_n12153_ = new_n6104_ & new_n10046_;
  assign new_n12154_ = new_n6104_ & new_n10048_;
  assign new_n12155_ = ~new_n12153_ & ~new_n12154_;
  assign new_n12156_ = ~new_n12152_ & new_n12155_;
  assign new_n12157_ = new_n12151_ & new_n12156_;
  assign new_n12158_ = new_n12146_ & new_n12157_;
  assign new_n12159_ = new_n6104_ & new_n10063_;
  assign new_n12160_ = new_n6104_ & new_n10052_;
  assign new_n12161_ = new_n6104_ & new_n10054_;
  assign new_n12162_ = ~new_n12160_ & ~new_n12161_;
  assign new_n12163_ = ~new_n12159_ & new_n12162_;
  assign new_n12164_ = new_n6104_ & new_n10071_;
  assign new_n12165_ = new_n6104_ & new_n10065_;
  assign new_n12166_ = new_n6104_ & new_n10061_;
  assign new_n12167_ = ~new_n12165_ & ~new_n12166_;
  assign new_n12168_ = ~new_n12164_ & new_n12167_;
  assign new_n12169_ = new_n12163_ & new_n12168_;
  assign new_n12170_ = new_n6104_ & new_n10080_;
  assign new_n12171_ = new_n6104_ & new_n10073_;
  assign new_n12172_ = new_n6104_ & new_n10069_;
  assign new_n12173_ = ~new_n12171_ & ~new_n12172_;
  assign new_n12174_ = ~new_n12170_ & new_n12173_;
  assign new_n12175_ = new_n6104_ & new_n10082_;
  assign new_n12176_ = new_n6104_ & new_n10078_;
  assign new_n12177_ = ~new_n12175_ & ~new_n12176_;
  assign new_n12178_ = new_n12174_ & new_n12177_;
  assign new_n12179_ = new_n12169_ & new_n12178_;
  assign new_n12180_ = new_n12158_ & new_n12179_;
  assign new_n12181_ = new_n6104_ & new_n10087_;
  assign new_n12182_ = new_n6104_ & new_n10089_;
  assign new_n12183_ = new_n6104_ & new_n10091_;
  assign new_n12184_ = ~new_n12182_ & ~new_n12183_;
  assign new_n12185_ = ~new_n12181_ & new_n12184_;
  assign new_n12186_ = new_n6104_ & new_n10098_;
  assign new_n12187_ = new_n6104_ & new_n10100_;
  assign new_n12188_ = new_n6104_ & new_n10102_;
  assign new_n12189_ = ~new_n12187_ & ~new_n12188_;
  assign new_n12190_ = ~new_n12186_ & new_n12189_;
  assign new_n12191_ = new_n12185_ & new_n12190_;
  assign new_n12192_ = new_n6104_ & new_n10107_;
  assign new_n12193_ = new_n6104_ & new_n10109_;
  assign new_n12194_ = new_n6104_ & new_n10111_;
  assign new_n12195_ = ~new_n12193_ & ~new_n12194_;
  assign new_n12196_ = ~new_n12192_ & new_n12195_;
  assign new_n12197_ = new_n6104_ & new_n10116_;
  assign new_n12198_ = new_n6104_ & new_n10118_;
  assign new_n12199_ = new_n6104_ & new_n10120_;
  assign new_n12200_ = ~new_n12198_ & ~new_n12199_;
  assign new_n12201_ = ~new_n12197_ & new_n12200_;
  assign new_n12202_ = new_n12196_ & new_n12201_;
  assign new_n12203_ = new_n12191_ & new_n12202_;
  assign new_n12204_ = new_n6267_ & new_n9924_;
  assign new_n12205_ = new_n6267_ & new_n9926_;
  assign new_n12206_ = new_n6267_ & new_n9928_;
  assign new_n12207_ = ~new_n12205_ & ~new_n12206_;
  assign new_n12208_ = ~new_n12204_ & new_n12207_;
  assign new_n12209_ = new_n6267_ & new_n9934_;
  assign new_n12210_ = new_n6267_ & new_n9936_;
  assign new_n12211_ = new_n6267_ & new_n9938_;
  assign new_n12212_ = ~new_n12210_ & ~new_n12211_;
  assign new_n12213_ = ~new_n12209_ & new_n12212_;
  assign new_n12214_ = new_n12208_ & new_n12213_;
  assign new_n12215_ = new_n6267_ & new_n9942_;
  assign new_n12216_ = new_n6267_ & new_n9944_;
  assign new_n12217_ = new_n6267_ & new_n9946_;
  assign new_n12218_ = ~new_n12216_ & ~new_n12217_;
  assign new_n12219_ = ~new_n12215_ & new_n12218_;
  assign new_n12220_ = new_n6267_ & new_n9954_;
  assign new_n12221_ = new_n6267_ & new_n9956_;
  assign new_n12222_ = ~new_n12220_ & ~new_n12221_;
  assign new_n12223_ = new_n12219_ & new_n12222_;
  assign new_n12224_ = new_n12214_ & new_n12223_;
  assign new_n12225_ = new_n12203_ & new_n12224_;
  assign new_n12226_ = new_n12180_ & new_n12225_;
  assign new_n12227_ = new_n6267_ & new_n9965_;
  assign new_n12228_ = new_n6267_ & new_n9952_;
  assign new_n12229_ = new_n6267_ & new_n9963_;
  assign new_n12230_ = ~new_n12228_ & ~new_n12229_;
  assign new_n12231_ = ~new_n12227_ & new_n12230_;
  assign new_n12232_ = new_n6267_ & new_n9974_;
  assign new_n12233_ = new_n6267_ & new_n9961_;
  assign new_n12234_ = new_n6267_ & new_n9972_;
  assign new_n12235_ = ~new_n12233_ & ~new_n12234_;
  assign new_n12236_ = ~new_n12232_ & new_n12235_;
  assign new_n12237_ = new_n12231_ & new_n12236_;
  assign new_n12238_ = new_n6267_ & new_n9980_;
  assign new_n12239_ = new_n6267_ & new_n9970_;
  assign new_n12240_ = new_n6267_ & new_n9978_;
  assign new_n12241_ = ~new_n12239_ & ~new_n12240_;
  assign new_n12242_ = ~new_n12238_ & new_n12241_;
  assign new_n12243_ = new_n6267_ & new_n9988_;
  assign new_n12244_ = new_n6267_ & new_n9990_;
  assign new_n12245_ = new_n6267_ & new_n9992_;
  assign new_n12246_ = ~new_n12244_ & ~new_n12245_;
  assign new_n12247_ = ~new_n12243_ & new_n12246_;
  assign new_n12248_ = new_n12242_ & new_n12247_;
  assign new_n12249_ = new_n12237_ & new_n12248_;
  assign new_n12250_ = new_n6267_ & new_n9997_;
  assign new_n12251_ = new_n6267_ & new_n9999_;
  assign new_n12252_ = new_n6267_ & new_n10001_;
  assign new_n12253_ = ~new_n12251_ & ~new_n12252_;
  assign new_n12254_ = ~new_n12250_ & new_n12253_;
  assign new_n12255_ = new_n6267_ & new_n10007_;
  assign new_n12256_ = new_n6267_ & new_n10009_;
  assign new_n12257_ = new_n6267_ & new_n10011_;
  assign new_n12258_ = ~new_n12256_ & ~new_n12257_;
  assign new_n12259_ = ~new_n12255_ & new_n12258_;
  assign new_n12260_ = new_n12254_ & new_n12259_;
  assign new_n12261_ = new_n6267_ & new_n10015_;
  assign new_n12262_ = new_n6267_ & new_n10017_;
  assign new_n12263_ = new_n6267_ & new_n10019_;
  assign new_n12264_ = ~new_n12262_ & ~new_n12263_;
  assign new_n12265_ = ~new_n12261_ & new_n12264_;
  assign new_n12266_ = new_n6267_ & new_n10028_;
  assign new_n12267_ = new_n6267_ & new_n10030_;
  assign new_n12268_ = ~new_n12266_ & ~new_n12267_;
  assign new_n12269_ = new_n12265_ & new_n12268_;
  assign new_n12270_ = new_n12260_ & new_n12269_;
  assign new_n12271_ = new_n12249_ & new_n12270_;
  assign new_n12272_ = new_n6267_ & new_n10039_;
  assign new_n12273_ = new_n6267_ & new_n10026_;
  assign new_n12274_ = new_n6267_ & new_n10037_;
  assign new_n12275_ = ~new_n12273_ & ~new_n12274_;
  assign new_n12276_ = ~new_n12272_ & new_n12275_;
  assign new_n12277_ = new_n6267_ & new_n10048_;
  assign new_n12278_ = new_n6267_ & new_n10035_;
  assign new_n12279_ = new_n6267_ & new_n10046_;
  assign new_n12280_ = ~new_n12278_ & ~new_n12279_;
  assign new_n12281_ = ~new_n12277_ & new_n12280_;
  assign new_n12282_ = new_n12276_ & new_n12281_;
  assign new_n12283_ = new_n6267_ & new_n10054_;
  assign new_n12284_ = new_n6267_ & new_n10044_;
  assign new_n12285_ = new_n6267_ & new_n10052_;
  assign new_n12286_ = ~new_n12284_ & ~new_n12285_;
  assign new_n12287_ = ~new_n12283_ & new_n12286_;
  assign new_n12288_ = new_n6267_ & new_n10061_;
  assign new_n12289_ = new_n6267_ & new_n10063_;
  assign new_n12290_ = new_n6267_ & new_n10065_;
  assign new_n12291_ = ~new_n12289_ & ~new_n12290_;
  assign new_n12292_ = ~new_n12288_ & new_n12291_;
  assign new_n12293_ = new_n12287_ & new_n12292_;
  assign new_n12294_ = new_n12282_ & new_n12293_;
  assign new_n12295_ = new_n6267_ & new_n10069_;
  assign new_n12296_ = new_n6267_ & new_n10071_;
  assign new_n12297_ = new_n6267_ & new_n10073_;
  assign new_n12298_ = ~new_n12296_ & ~new_n12297_;
  assign new_n12299_ = ~new_n12295_ & new_n12298_;
  assign new_n12300_ = new_n6267_ & new_n10078_;
  assign new_n12301_ = new_n6267_ & new_n10080_;
  assign new_n12302_ = new_n6267_ & new_n10082_;
  assign new_n12303_ = ~new_n12301_ & ~new_n12302_;
  assign new_n12304_ = ~new_n12300_ & new_n12303_;
  assign new_n12305_ = new_n12299_ & new_n12304_;
  assign new_n12306_ = new_n6267_ & new_n10087_;
  assign new_n12307_ = new_n6267_ & new_n10089_;
  assign new_n12308_ = new_n6267_ & new_n10091_;
  assign new_n12309_ = ~new_n12307_ & ~new_n12308_;
  assign new_n12310_ = ~new_n12306_ & new_n12309_;
  assign new_n12311_ = new_n6267_ & new_n10100_;
  assign new_n12312_ = new_n6267_ & new_n10102_;
  assign new_n12313_ = ~new_n12311_ & ~new_n12312_;
  assign new_n12314_ = new_n12310_ & new_n12313_;
  assign new_n12315_ = new_n12305_ & new_n12314_;
  assign new_n12316_ = new_n12294_ & new_n12315_;
  assign new_n12317_ = new_n12271_ & new_n12316_;
  assign new_n12318_ = new_n12226_ & new_n12317_;
  assign new_n12319_ = new_n12135_ & new_n12318_;
  assign new_n12320_ = new_n11952_ & new_n12319_;
  assign new_n12321_ = new_n6267_ & new_n10111_;
  assign new_n12322_ = new_n6267_ & new_n10098_;
  assign new_n12323_ = new_n6267_ & new_n10109_;
  assign new_n12324_ = ~new_n12322_ & ~new_n12323_;
  assign new_n12325_ = ~new_n12321_ & new_n12324_;
  assign new_n12326_ = new_n6267_ & new_n10120_;
  assign new_n12327_ = new_n6267_ & new_n10107_;
  assign new_n12328_ = new_n6267_ & new_n10118_;
  assign new_n12329_ = ~new_n12327_ & ~new_n12328_;
  assign new_n12330_ = ~new_n12326_ & new_n12329_;
  assign new_n12331_ = new_n12325_ & new_n12330_;
  assign new_n12332_ = new_n6424_ & new_n9928_;
  assign new_n12333_ = new_n6267_ & new_n10116_;
  assign new_n12334_ = new_n6424_ & new_n9926_;
  assign new_n12335_ = ~new_n12333_ & ~new_n12334_;
  assign new_n12336_ = ~new_n12332_ & new_n12335_;
  assign new_n12337_ = new_n6424_ & new_n9938_;
  assign new_n12338_ = new_n6424_ & new_n9924_;
  assign new_n12339_ = new_n6424_ & new_n9936_;
  assign new_n12340_ = ~new_n12338_ & ~new_n12339_;
  assign new_n12341_ = ~new_n12337_ & new_n12340_;
  assign new_n12342_ = new_n12336_ & new_n12341_;
  assign new_n12343_ = new_n12331_ & new_n12342_;
  assign new_n12344_ = new_n6424_ & new_n9946_;
  assign new_n12345_ = new_n6424_ & new_n9934_;
  assign new_n12346_ = new_n6424_ & new_n9944_;
  assign new_n12347_ = ~new_n12345_ & ~new_n12346_;
  assign new_n12348_ = ~new_n12344_ & new_n12347_;
  assign new_n12349_ = new_n6424_ & new_n9956_;
  assign new_n12350_ = new_n6424_ & new_n9942_;
  assign new_n12351_ = new_n6424_ & new_n9954_;
  assign new_n12352_ = ~new_n12350_ & ~new_n12351_;
  assign new_n12353_ = ~new_n12349_ & new_n12352_;
  assign new_n12354_ = new_n12348_ & new_n12353_;
  assign new_n12355_ = new_n6424_ & new_n9965_;
  assign new_n12356_ = new_n6424_ & new_n9952_;
  assign new_n12357_ = new_n6424_ & new_n9963_;
  assign new_n12358_ = ~new_n12356_ & ~new_n12357_;
  assign new_n12359_ = ~new_n12355_ & new_n12358_;
  assign new_n12360_ = new_n6424_ & new_n9974_;
  assign new_n12361_ = new_n6424_ & new_n9961_;
  assign new_n12362_ = new_n6424_ & new_n9972_;
  assign new_n12363_ = ~new_n12361_ & ~new_n12362_;
  assign new_n12364_ = ~new_n12360_ & new_n12363_;
  assign new_n12365_ = new_n12359_ & new_n12364_;
  assign new_n12366_ = new_n12354_ & new_n12365_;
  assign new_n12367_ = new_n12343_ & new_n12366_;
  assign new_n12368_ = new_n6424_ & new_n9980_;
  assign new_n12369_ = new_n6424_ & new_n9970_;
  assign new_n12370_ = new_n6424_ & new_n9978_;
  assign new_n12371_ = ~new_n12369_ & ~new_n12370_;
  assign new_n12372_ = ~new_n12368_ & new_n12371_;
  assign new_n12373_ = new_n6424_ & new_n9988_;
  assign new_n12374_ = new_n6424_ & new_n9990_;
  assign new_n12375_ = new_n6424_ & new_n9992_;
  assign new_n12376_ = ~new_n12374_ & ~new_n12375_;
  assign new_n12377_ = ~new_n12373_ & new_n12376_;
  assign new_n12378_ = new_n12372_ & new_n12377_;
  assign new_n12379_ = new_n6424_ & new_n9997_;
  assign new_n12380_ = new_n6424_ & new_n9999_;
  assign new_n12381_ = new_n6424_ & new_n10001_;
  assign new_n12382_ = ~new_n12380_ & ~new_n12381_;
  assign new_n12383_ = ~new_n12379_ & new_n12382_;
  assign new_n12384_ = new_n6424_ & new_n10007_;
  assign new_n12385_ = new_n6424_ & new_n10009_;
  assign new_n12386_ = new_n6424_ & new_n10011_;
  assign new_n12387_ = ~new_n12385_ & ~new_n12386_;
  assign new_n12388_ = ~new_n12384_ & new_n12387_;
  assign new_n12389_ = new_n12383_ & new_n12388_;
  assign new_n12390_ = new_n12378_ & new_n12389_;
  assign new_n12391_ = new_n6424_ & new_n10015_;
  assign new_n12392_ = new_n6424_ & new_n10017_;
  assign new_n12393_ = new_n6424_ & new_n10019_;
  assign new_n12394_ = ~new_n12392_ & ~new_n12393_;
  assign new_n12395_ = ~new_n12391_ & new_n12394_;
  assign new_n12396_ = new_n6424_ & new_n10026_;
  assign new_n12397_ = new_n6424_ & new_n10028_;
  assign new_n12398_ = new_n6424_ & new_n10030_;
  assign new_n12399_ = ~new_n12397_ & ~new_n12398_;
  assign new_n12400_ = ~new_n12396_ & new_n12399_;
  assign new_n12401_ = new_n12395_ & new_n12400_;
  assign new_n12402_ = new_n6424_ & new_n10035_;
  assign new_n12403_ = new_n6424_ & new_n10037_;
  assign new_n12404_ = new_n6424_ & new_n10039_;
  assign new_n12405_ = ~new_n12403_ & ~new_n12404_;
  assign new_n12406_ = ~new_n12402_ & new_n12405_;
  assign new_n12407_ = new_n6424_ & new_n10046_;
  assign new_n12408_ = new_n6424_ & new_n10048_;
  assign new_n12409_ = ~new_n12407_ & ~new_n12408_;
  assign new_n12410_ = new_n12406_ & new_n12409_;
  assign new_n12411_ = new_n12401_ & new_n12410_;
  assign new_n12412_ = new_n12390_ & new_n12411_;
  assign new_n12413_ = new_n12367_ & new_n12412_;
  assign new_n12414_ = new_n6424_ & new_n10054_;
  assign new_n12415_ = new_n6424_ & new_n10044_;
  assign new_n12416_ = new_n6424_ & new_n10052_;
  assign new_n12417_ = ~new_n12415_ & ~new_n12416_;
  assign new_n12418_ = ~new_n12414_ & new_n12417_;
  assign new_n12419_ = new_n6424_ & new_n10061_;
  assign new_n12420_ = new_n6424_ & new_n10063_;
  assign new_n12421_ = new_n6424_ & new_n10065_;
  assign new_n12422_ = ~new_n12420_ & ~new_n12421_;
  assign new_n12423_ = ~new_n12419_ & new_n12422_;
  assign new_n12424_ = new_n12418_ & new_n12423_;
  assign new_n12425_ = new_n6424_ & new_n10069_;
  assign new_n12426_ = new_n6424_ & new_n10071_;
  assign new_n12427_ = new_n6424_ & new_n10073_;
  assign new_n12428_ = ~new_n12426_ & ~new_n12427_;
  assign new_n12429_ = ~new_n12425_ & new_n12428_;
  assign new_n12430_ = new_n6424_ & new_n10078_;
  assign new_n12431_ = new_n6424_ & new_n10080_;
  assign new_n12432_ = new_n6424_ & new_n10082_;
  assign new_n12433_ = ~new_n12431_ & ~new_n12432_;
  assign new_n12434_ = ~new_n12430_ & new_n12433_;
  assign new_n12435_ = new_n12429_ & new_n12434_;
  assign new_n12436_ = new_n12424_ & new_n12435_;
  assign new_n12437_ = new_n6424_ & new_n10087_;
  assign new_n12438_ = new_n6424_ & new_n10089_;
  assign new_n12439_ = new_n6424_ & new_n10091_;
  assign new_n12440_ = ~new_n12438_ & ~new_n12439_;
  assign new_n12441_ = ~new_n12437_ & new_n12440_;
  assign new_n12442_ = new_n6424_ & new_n10098_;
  assign new_n12443_ = new_n6424_ & new_n10100_;
  assign new_n12444_ = new_n6424_ & new_n10102_;
  assign new_n12445_ = ~new_n12443_ & ~new_n12444_;
  assign new_n12446_ = ~new_n12442_ & new_n12445_;
  assign new_n12447_ = new_n12441_ & new_n12446_;
  assign new_n12448_ = new_n6424_ & new_n10107_;
  assign new_n12449_ = new_n6424_ & new_n10109_;
  assign new_n12450_ = new_n6424_ & new_n10111_;
  assign new_n12451_ = ~new_n12449_ & ~new_n12450_;
  assign new_n12452_ = ~new_n12448_ & new_n12451_;
  assign new_n12453_ = new_n6424_ & new_n10118_;
  assign new_n12454_ = new_n6424_ & new_n10120_;
  assign new_n12455_ = ~new_n12453_ & ~new_n12454_;
  assign new_n12456_ = new_n12452_ & new_n12455_;
  assign new_n12457_ = new_n12447_ & new_n12456_;
  assign new_n12458_ = new_n12436_ & new_n12457_;
  assign new_n12459_ = new_n6525_ & new_n10132_;
  assign new_n12460_ = new_n10131_ & new_n12459_;
  assign new_n12461_ = new_n6424_ & new_n10116_;
  assign new_n12462_ = new_n6525_ & new_n10127_;
  assign new_n12463_ = new_n10125_ & new_n12462_;
  assign new_n12464_ = ~new_n12461_ & ~new_n12463_;
  assign new_n12465_ = ~new_n12460_ & new_n12464_;
  assign new_n12466_ = new_n6525_ & new_n10142_;
  assign new_n12467_ = new_n10125_ & new_n12466_;
  assign new_n12468_ = new_n6525_ & new_n10147_;
  assign new_n12469_ = new_n10146_ & new_n12468_;
  assign new_n12470_ = new_n10151_ & new_n12468_;
  assign new_n12471_ = ~new_n12469_ & ~new_n12470_;
  assign new_n12472_ = ~new_n12467_ & new_n12471_;
  assign new_n12473_ = new_n12465_ & new_n12472_;
  assign new_n12474_ = new_n6525_ & new_n10155_;
  assign new_n12475_ = new_n10151_ & new_n12474_;
  assign new_n12476_ = new_n6525_ & new_n10158_;
  assign new_n12477_ = new_n10131_ & new_n12476_;
  assign new_n12478_ = new_n10146_ & new_n12474_;
  assign new_n12479_ = ~new_n12477_ & ~new_n12478_;
  assign new_n12480_ = ~new_n12475_ & new_n12479_;
  assign new_n12481_ = new_n6525_ & new_n10166_;
  assign new_n12482_ = new_n10146_ & new_n12481_;
  assign new_n12483_ = new_n6525_ & new_n10169_;
  assign new_n12484_ = new_n10125_ & new_n12483_;
  assign new_n12485_ = new_n6525_ & new_n10172_;
  assign new_n12486_ = new_n10131_ & new_n12485_;
  assign new_n12487_ = ~new_n12484_ & ~new_n12486_;
  assign new_n12488_ = ~new_n12482_ & new_n12487_;
  assign new_n12489_ = new_n12480_ & new_n12488_;
  assign new_n12490_ = new_n12473_ & new_n12489_;
  assign new_n12491_ = new_n6525_ & new_n10177_;
  assign new_n12492_ = new_n10131_ & new_n12491_;
  assign new_n12493_ = new_n10151_ & new_n12481_;
  assign new_n12494_ = new_n6525_ & new_n10181_;
  assign new_n12495_ = new_n10125_ & new_n12494_;
  assign new_n12496_ = ~new_n12493_ & ~new_n12495_;
  assign new_n12497_ = ~new_n12492_ & new_n12496_;
  assign new_n12498_ = new_n6526_ & new_n8617_;
  assign new_n12499_ = new_n6525_ & new_n10189_;
  assign new_n12500_ = new_n10146_ & new_n12499_;
  assign new_n12501_ = new_n10151_ & new_n12499_;
  assign new_n12502_ = ~new_n12500_ & ~new_n12501_;
  assign new_n12503_ = ~new_n12498_ & new_n12502_;
  assign new_n12504_ = new_n12497_ & new_n12503_;
  assign new_n12505_ = new_n6526_ & new_n8625_;
  assign new_n12506_ = new_n6526_ & new_n8628_;
  assign new_n12507_ = new_n6526_ & new_n8630_;
  assign new_n12508_ = ~new_n12506_ & ~new_n12507_;
  assign new_n12509_ = ~new_n12505_ & new_n12508_;
  assign new_n12510_ = new_n6526_ & new_n8637_;
  assign new_n12511_ = new_n6526_ & new_n8639_;
  assign new_n12512_ = ~new_n12510_ & ~new_n12511_;
  assign new_n12513_ = new_n12509_ & new_n12512_;
  assign new_n12514_ = new_n12504_ & new_n12513_;
  assign new_n12515_ = new_n12490_ & new_n12514_;
  assign new_n12516_ = new_n12458_ & new_n12515_;
  assign new_n12517_ = new_n12413_ & new_n12516_;
  assign new_n12518_ = new_n6526_ & new_n8650_;
  assign new_n12519_ = new_n6526_ & new_n8635_;
  assign new_n12520_ = new_n6526_ & new_n8648_;
  assign new_n12521_ = ~new_n12519_ & ~new_n12520_;
  assign new_n12522_ = ~new_n12518_ & new_n12521_;
  assign new_n12523_ = new_n6526_ & new_n8659_;
  assign new_n12524_ = new_n6526_ & new_n8646_;
  assign new_n12525_ = new_n6526_ & new_n8657_;
  assign new_n12526_ = ~new_n12524_ & ~new_n12525_;
  assign new_n12527_ = ~new_n12523_ & new_n12526_;
  assign new_n12528_ = new_n12522_ & new_n12527_;
  assign new_n12529_ = new_n6526_ & new_n8670_;
  assign new_n12530_ = new_n6526_ & new_n8655_;
  assign new_n12531_ = new_n6526_ & new_n8667_;
  assign new_n12532_ = ~new_n12530_ & ~new_n12531_;
  assign new_n12533_ = ~new_n12529_ & new_n12532_;
  assign new_n12534_ = new_n6526_ & new_n8681_;
  assign new_n12535_ = new_n6526_ & new_n8665_;
  assign new_n12536_ = new_n6526_ & new_n8678_;
  assign new_n12537_ = ~new_n12535_ & ~new_n12536_;
  assign new_n12538_ = ~new_n12534_ & new_n12537_;
  assign new_n12539_ = new_n12533_ & new_n12538_;
  assign new_n12540_ = new_n12528_ & new_n12539_;
  assign new_n12541_ = new_n6526_ & new_n8694_;
  assign new_n12542_ = new_n6526_ & new_n8675_;
  assign new_n12543_ = new_n6526_ & new_n8692_;
  assign new_n12544_ = ~new_n12542_ & ~new_n12543_;
  assign new_n12545_ = ~new_n12541_ & new_n12544_;
  assign new_n12546_ = new_n6526_ & new_n8701_;
  assign new_n12547_ = new_n6526_ & new_n8689_;
  assign new_n12548_ = new_n6526_ & new_n8699_;
  assign new_n12549_ = ~new_n12547_ & ~new_n12548_;
  assign new_n12550_ = ~new_n12546_ & new_n12549_;
  assign new_n12551_ = new_n12545_ & new_n12550_;
  assign new_n12552_ = new_n6533_ & new_n10241_;
  assign new_n12553_ = new_n10146_ & new_n12552_;
  assign new_n12554_ = new_n6533_ & new_n10244_;
  assign new_n12555_ = new_n10125_ & new_n12554_;
  assign new_n12556_ = new_n6533_ & new_n10247_;
  assign new_n12557_ = new_n10131_ & new_n12556_;
  assign new_n12558_ = ~new_n12555_ & ~new_n12557_;
  assign new_n12559_ = ~new_n12553_ & new_n12558_;
  assign new_n12560_ = new_n10151_ & new_n12552_;
  assign new_n12561_ = new_n6533_ & new_n10258_;
  assign new_n12562_ = new_n10125_ & new_n12561_;
  assign new_n12563_ = ~new_n12560_ & ~new_n12562_;
  assign new_n12564_ = new_n12559_ & new_n12563_;
  assign new_n12565_ = new_n12551_ & new_n12564_;
  assign new_n12566_ = new_n12540_ & new_n12565_;
  assign new_n12567_ = new_n6533_ & new_n10263_;
  assign new_n12568_ = new_n10151_ & new_n12567_;
  assign new_n12569_ = new_n6533_ & new_n10254_;
  assign new_n12570_ = new_n10131_ & new_n12569_;
  assign new_n12571_ = new_n10146_ & new_n12567_;
  assign new_n12572_ = ~new_n12570_ & ~new_n12571_;
  assign new_n12573_ = ~new_n12568_ & new_n12572_;
  assign new_n12574_ = new_n6533_ & new_n10273_;
  assign new_n12575_ = new_n10146_ & new_n12574_;
  assign new_n12576_ = new_n6533_ & new_n10276_;
  assign new_n12577_ = new_n10125_ & new_n12576_;
  assign new_n12578_ = new_n6533_ & new_n10279_;
  assign new_n12579_ = new_n10131_ & new_n12578_;
  assign new_n12580_ = ~new_n12577_ & ~new_n12579_;
  assign new_n12581_ = ~new_n12575_ & new_n12580_;
  assign new_n12582_ = new_n12573_ & new_n12581_;
  assign new_n12583_ = new_n6533_ & new_n10284_;
  assign new_n12584_ = new_n10131_ & new_n12583_;
  assign new_n12585_ = new_n10151_ & new_n12574_;
  assign new_n12586_ = new_n6533_ & new_n10288_;
  assign new_n12587_ = new_n10125_ & new_n12586_;
  assign new_n12588_ = ~new_n12585_ & ~new_n12587_;
  assign new_n12589_ = ~new_n12584_ & new_n12588_;
  assign new_n12590_ = new_n6534_ & new_n8617_;
  assign new_n12591_ = new_n6533_ & new_n10295_;
  assign new_n12592_ = new_n10146_ & new_n12591_;
  assign new_n12593_ = new_n10151_ & new_n12591_;
  assign new_n12594_ = ~new_n12592_ & ~new_n12593_;
  assign new_n12595_ = ~new_n12590_ & new_n12594_;
  assign new_n12596_ = new_n12589_ & new_n12595_;
  assign new_n12597_ = new_n12582_ & new_n12596_;
  assign new_n12598_ = new_n6534_ & new_n8625_;
  assign new_n12599_ = new_n6534_ & new_n8628_;
  assign new_n12600_ = new_n6534_ & new_n8630_;
  assign new_n12601_ = ~new_n12599_ & ~new_n12600_;
  assign new_n12602_ = ~new_n12598_ & new_n12601_;
  assign new_n12603_ = new_n6534_ & new_n8635_;
  assign new_n12604_ = new_n6534_ & new_n8637_;
  assign new_n12605_ = new_n6534_ & new_n8639_;
  assign new_n12606_ = ~new_n12604_ & ~new_n12605_;
  assign new_n12607_ = ~new_n12603_ & new_n12606_;
  assign new_n12608_ = new_n12602_ & new_n12607_;
  assign new_n12609_ = new_n6534_ & new_n8646_;
  assign new_n12610_ = new_n6534_ & new_n8648_;
  assign new_n12611_ = new_n6534_ & new_n8650_;
  assign new_n12612_ = ~new_n12610_ & ~new_n12611_;
  assign new_n12613_ = ~new_n12609_ & new_n12612_;
  assign new_n12614_ = new_n6534_ & new_n8657_;
  assign new_n12615_ = new_n6534_ & new_n8659_;
  assign new_n12616_ = ~new_n12614_ & ~new_n12615_;
  assign new_n12617_ = new_n12613_ & new_n12616_;
  assign new_n12618_ = new_n12608_ & new_n12617_;
  assign new_n12619_ = new_n12597_ & new_n12618_;
  assign new_n12620_ = new_n12566_ & new_n12619_;
  assign new_n12621_ = new_n6534_ & new_n8670_;
  assign new_n12622_ = new_n6534_ & new_n8655_;
  assign new_n12623_ = new_n6534_ & new_n8667_;
  assign new_n12624_ = ~new_n12622_ & ~new_n12623_;
  assign new_n12625_ = ~new_n12621_ & new_n12624_;
  assign new_n12626_ = new_n6534_ & new_n8681_;
  assign new_n12627_ = new_n6534_ & new_n8665_;
  assign new_n12628_ = new_n6534_ & new_n8678_;
  assign new_n12629_ = ~new_n12627_ & ~new_n12628_;
  assign new_n12630_ = ~new_n12626_ & new_n12629_;
  assign new_n12631_ = new_n12625_ & new_n12630_;
  assign new_n12632_ = new_n6534_ & new_n8694_;
  assign new_n12633_ = new_n6534_ & new_n8675_;
  assign new_n12634_ = new_n6534_ & new_n8692_;
  assign new_n12635_ = ~new_n12633_ & ~new_n12634_;
  assign new_n12636_ = ~new_n12632_ & new_n12635_;
  assign new_n12637_ = new_n6534_ & new_n8701_;
  assign new_n12638_ = new_n6534_ & new_n8689_;
  assign new_n12639_ = new_n6534_ & new_n8699_;
  assign new_n12640_ = ~new_n12638_ & ~new_n12639_;
  assign new_n12641_ = ~new_n12637_ & new_n12640_;
  assign new_n12642_ = new_n12636_ & new_n12641_;
  assign new_n12643_ = new_n12631_ & new_n12642_;
  assign new_n12644_ = new_n6547_ & new_n10346_;
  assign new_n12645_ = new_n10146_ & new_n12644_;
  assign new_n12646_ = new_n6547_ & new_n10349_;
  assign new_n12647_ = new_n10125_ & new_n12646_;
  assign new_n12648_ = new_n6547_ & new_n10352_;
  assign new_n12649_ = new_n10131_ & new_n12648_;
  assign new_n12650_ = ~new_n12647_ & ~new_n12649_;
  assign new_n12651_ = ~new_n12645_ & new_n12650_;
  assign new_n12652_ = new_n6547_ & new_n10359_;
  assign new_n12653_ = new_n10131_ & new_n12652_;
  assign new_n12654_ = new_n10151_ & new_n12644_;
  assign new_n12655_ = new_n6547_ & new_n10363_;
  assign new_n12656_ = new_n10125_ & new_n12655_;
  assign new_n12657_ = ~new_n12654_ & ~new_n12656_;
  assign new_n12658_ = ~new_n12653_ & new_n12657_;
  assign new_n12659_ = new_n12651_ & new_n12658_;
  assign new_n12660_ = new_n6547_ & new_n10369_;
  assign new_n12661_ = new_n10125_ & new_n12660_;
  assign new_n12662_ = new_n6547_ & new_n10372_;
  assign new_n12663_ = new_n10146_ & new_n12662_;
  assign new_n12664_ = new_n10151_ & new_n12662_;
  assign new_n12665_ = ~new_n12663_ & ~new_n12664_;
  assign new_n12666_ = ~new_n12661_ & new_n12665_;
  assign new_n12667_ = new_n6547_ & new_n10382_;
  assign new_n12668_ = new_n10131_ & new_n12667_;
  assign new_n12669_ = new_n6547_ & new_n10379_;
  assign new_n12670_ = new_n10146_ & new_n12669_;
  assign new_n12671_ = ~new_n12668_ & ~new_n12670_;
  assign new_n12672_ = new_n12666_ & new_n12671_;
  assign new_n12673_ = new_n12659_ & new_n12672_;
  assign new_n12674_ = new_n12643_ & new_n12673_;
  assign new_n12675_ = new_n6547_ & new_n10391_;
  assign new_n12676_ = new_n10131_ & new_n12675_;
  assign new_n12677_ = new_n10151_ & new_n12669_;
  assign new_n12678_ = new_n6547_ & new_n10388_;
  assign new_n12679_ = new_n10125_ & new_n12678_;
  assign new_n12680_ = ~new_n12677_ & ~new_n12679_;
  assign new_n12681_ = ~new_n12676_ & new_n12680_;
  assign new_n12682_ = new_n6548_ & new_n8617_;
  assign new_n12683_ = new_n6547_ & new_n10402_;
  assign new_n12684_ = new_n10146_ & new_n12683_;
  assign new_n12685_ = new_n10151_ & new_n12683_;
  assign new_n12686_ = ~new_n12684_ & ~new_n12685_;
  assign new_n12687_ = ~new_n12682_ & new_n12686_;
  assign new_n12688_ = new_n12681_ & new_n12687_;
  assign new_n12689_ = new_n6548_ & new_n8625_;
  assign new_n12690_ = new_n6548_ & new_n8628_;
  assign new_n12691_ = new_n6548_ & new_n8630_;
  assign new_n12692_ = ~new_n12690_ & ~new_n12691_;
  assign new_n12693_ = ~new_n12689_ & new_n12692_;
  assign new_n12694_ = new_n6548_ & new_n8635_;
  assign new_n12695_ = new_n6548_ & new_n8637_;
  assign new_n12696_ = new_n6548_ & new_n8639_;
  assign new_n12697_ = ~new_n12695_ & ~new_n12696_;
  assign new_n12698_ = ~new_n12694_ & new_n12697_;
  assign new_n12699_ = new_n12693_ & new_n12698_;
  assign new_n12700_ = new_n12688_ & new_n12699_;
  assign new_n12701_ = new_n6548_ & new_n8646_;
  assign new_n12702_ = new_n6548_ & new_n8648_;
  assign new_n12703_ = new_n6548_ & new_n8650_;
  assign new_n12704_ = ~new_n12702_ & ~new_n12703_;
  assign new_n12705_ = ~new_n12701_ & new_n12704_;
  assign new_n12706_ = new_n6548_ & new_n8655_;
  assign new_n12707_ = new_n6548_ & new_n8657_;
  assign new_n12708_ = new_n6548_ & new_n8659_;
  assign new_n12709_ = ~new_n12707_ & ~new_n12708_;
  assign new_n12710_ = ~new_n12706_ & new_n12709_;
  assign new_n12711_ = new_n12705_ & new_n12710_;
  assign new_n12712_ = new_n6548_ & new_n8665_;
  assign new_n12713_ = new_n6548_ & new_n8667_;
  assign new_n12714_ = new_n6548_ & new_n8670_;
  assign new_n12715_ = ~new_n12713_ & ~new_n12714_;
  assign new_n12716_ = ~new_n12712_ & new_n12715_;
  assign new_n12717_ = new_n6548_ & new_n8678_;
  assign new_n12718_ = new_n6548_ & new_n8681_;
  assign new_n12719_ = ~new_n12717_ & ~new_n12718_;
  assign new_n12720_ = new_n12716_ & new_n12719_;
  assign new_n12721_ = new_n12711_ & new_n12720_;
  assign new_n12722_ = new_n12700_ & new_n12721_;
  assign new_n12723_ = new_n12674_ & new_n12722_;
  assign new_n12724_ = new_n12620_ & new_n12723_;
  assign new_n12725_ = new_n12517_ & new_n12724_;
  assign new_n12726_ = new_n6548_ & new_n8694_;
  assign new_n12727_ = new_n6548_ & new_n8675_;
  assign new_n12728_ = new_n6548_ & new_n8692_;
  assign new_n12729_ = ~new_n12727_ & ~new_n12728_;
  assign new_n12730_ = ~new_n12726_ & new_n12729_;
  assign new_n12731_ = new_n6548_ & new_n8701_;
  assign new_n12732_ = new_n6548_ & new_n8689_;
  assign new_n12733_ = new_n6548_ & new_n8699_;
  assign new_n12734_ = ~new_n12732_ & ~new_n12733_;
  assign new_n12735_ = ~new_n12731_ & new_n12734_;
  assign new_n12736_ = new_n12730_ & new_n12735_;
  assign new_n12737_ = new_n6547_ & new_n10457_;
  assign new_n12738_ = new_n10146_ & new_n12737_;
  assign new_n12739_ = new_n6547_ & new_n10450_;
  assign new_n12740_ = new_n10125_ & new_n12739_;
  assign new_n12741_ = new_n6547_ & new_n10460_;
  assign new_n12742_ = new_n10131_ & new_n12741_;
  assign new_n12743_ = ~new_n12740_ & ~new_n12742_;
  assign new_n12744_ = ~new_n12738_ & new_n12743_;
  assign new_n12745_ = new_n6547_ & new_n10473_;
  assign new_n12746_ = new_n10131_ & new_n12745_;
  assign new_n12747_ = new_n10151_ & new_n12737_;
  assign new_n12748_ = new_n6547_ & new_n10470_;
  assign new_n12749_ = new_n10125_ & new_n12748_;
  assign new_n12750_ = ~new_n12747_ & ~new_n12749_;
  assign new_n12751_ = ~new_n12746_ & new_n12750_;
  assign new_n12752_ = new_n12744_ & new_n12751_;
  assign new_n12753_ = new_n12736_ & new_n12752_;
  assign new_n12754_ = new_n6547_ & new_n10483_;
  assign new_n12755_ = new_n10125_ & new_n12754_;
  assign new_n12756_ = new_n6547_ & new_n10467_;
  assign new_n12757_ = new_n10146_ & new_n12756_;
  assign new_n12758_ = new_n10151_ & new_n12756_;
  assign new_n12759_ = ~new_n12757_ & ~new_n12758_;
  assign new_n12760_ = ~new_n12755_ & new_n12759_;
  assign new_n12761_ = new_n6547_ & new_n10493_;
  assign new_n12762_ = new_n10151_ & new_n12761_;
  assign new_n12763_ = new_n6547_ & new_n10479_;
  assign new_n12764_ = new_n10131_ & new_n12763_;
  assign new_n12765_ = new_n10146_ & new_n12761_;
  assign new_n12766_ = ~new_n12764_ & ~new_n12765_;
  assign new_n12767_ = ~new_n12762_ & new_n12766_;
  assign new_n12768_ = new_n12760_ & new_n12767_;
  assign new_n12769_ = new_n6547_ & new_n10499_;
  assign new_n12770_ = new_n10146_ & new_n12769_;
  assign new_n12771_ = new_n6547_ & new_n10490_;
  assign new_n12772_ = new_n10125_ & new_n12771_;
  assign new_n12773_ = new_n6547_ & new_n10502_;
  assign new_n12774_ = new_n10131_ & new_n12773_;
  assign new_n12775_ = ~new_n12772_ & ~new_n12774_;
  assign new_n12776_ = ~new_n12770_ & new_n12775_;
  assign new_n12777_ = new_n10151_ & new_n12769_;
  assign new_n12778_ = new_n6555_ & new_n8617_;
  assign new_n12779_ = ~new_n12777_ & ~new_n12778_;
  assign new_n12780_ = new_n12776_ & new_n12779_;
  assign new_n12781_ = new_n12768_ & new_n12780_;
  assign new_n12782_ = new_n12753_ & new_n12781_;
  assign new_n12783_ = new_n6555_ & new_n8625_;
  assign new_n12784_ = new_n6555_ & new_n8628_;
  assign new_n12785_ = new_n6555_ & new_n8630_;
  assign new_n12786_ = ~new_n12784_ & ~new_n12785_;
  assign new_n12787_ = ~new_n12783_ & new_n12786_;
  assign new_n12788_ = new_n6555_ & new_n8635_;
  assign new_n12789_ = new_n6555_ & new_n8637_;
  assign new_n12790_ = new_n6555_ & new_n8639_;
  assign new_n12791_ = ~new_n12789_ & ~new_n12790_;
  assign new_n12792_ = ~new_n12788_ & new_n12791_;
  assign new_n12793_ = new_n12787_ & new_n12792_;
  assign new_n12794_ = new_n6555_ & new_n8646_;
  assign new_n12795_ = new_n6555_ & new_n8648_;
  assign new_n12796_ = new_n6555_ & new_n8650_;
  assign new_n12797_ = ~new_n12795_ & ~new_n12796_;
  assign new_n12798_ = ~new_n12794_ & new_n12797_;
  assign new_n12799_ = new_n6555_ & new_n8655_;
  assign new_n12800_ = new_n6555_ & new_n8657_;
  assign new_n12801_ = new_n6555_ & new_n8659_;
  assign new_n12802_ = ~new_n12800_ & ~new_n12801_;
  assign new_n12803_ = ~new_n12799_ & new_n12802_;
  assign new_n12804_ = new_n12798_ & new_n12803_;
  assign new_n12805_ = new_n12793_ & new_n12804_;
  assign new_n12806_ = new_n6555_ & new_n8665_;
  assign new_n12807_ = new_n6555_ & new_n8667_;
  assign new_n12808_ = new_n6555_ & new_n8670_;
  assign new_n12809_ = ~new_n12807_ & ~new_n12808_;
  assign new_n12810_ = ~new_n12806_ & new_n12809_;
  assign new_n12811_ = new_n6555_ & new_n8675_;
  assign new_n12812_ = new_n6555_ & new_n8678_;
  assign new_n12813_ = new_n6555_ & new_n8681_;
  assign new_n12814_ = ~new_n12812_ & ~new_n12813_;
  assign new_n12815_ = ~new_n12811_ & new_n12814_;
  assign new_n12816_ = new_n12810_ & new_n12815_;
  assign new_n12817_ = new_n6555_ & new_n8689_;
  assign new_n12818_ = new_n6555_ & new_n8692_;
  assign new_n12819_ = new_n6555_ & new_n8694_;
  assign new_n12820_ = ~new_n12818_ & ~new_n12819_;
  assign new_n12821_ = ~new_n12817_ & new_n12820_;
  assign new_n12822_ = new_n6555_ & new_n8699_;
  assign new_n12823_ = new_n6555_ & new_n8701_;
  assign new_n12824_ = ~new_n12822_ & ~new_n12823_;
  assign new_n12825_ = new_n12821_ & new_n12824_;
  assign new_n12826_ = new_n12816_ & new_n12825_;
  assign new_n12827_ = new_n12805_ & new_n12826_;
  assign new_n12828_ = new_n12782_ & new_n12827_;
  assign new_n12829_ = new_n6569_ & new_n8630_;
  assign new_n12830_ = new_n6569_ & new_n8617_;
  assign new_n12831_ = new_n6569_ & new_n8628_;
  assign new_n12832_ = ~new_n12830_ & ~new_n12831_;
  assign new_n12833_ = ~new_n12829_ & new_n12832_;
  assign new_n12834_ = new_n6569_ & new_n8639_;
  assign new_n12835_ = new_n6569_ & new_n8625_;
  assign new_n12836_ = new_n6569_ & new_n8637_;
  assign new_n12837_ = ~new_n12835_ & ~new_n12836_;
  assign new_n12838_ = ~new_n12834_ & new_n12837_;
  assign new_n12839_ = new_n12833_ & new_n12838_;
  assign new_n12840_ = new_n6569_ & new_n8650_;
  assign new_n12841_ = new_n6569_ & new_n8635_;
  assign new_n12842_ = new_n6569_ & new_n8648_;
  assign new_n12843_ = ~new_n12841_ & ~new_n12842_;
  assign new_n12844_ = ~new_n12840_ & new_n12843_;
  assign new_n12845_ = new_n6569_ & new_n8659_;
  assign new_n12846_ = new_n6569_ & new_n8646_;
  assign new_n12847_ = new_n6569_ & new_n8657_;
  assign new_n12848_ = ~new_n12846_ & ~new_n12847_;
  assign new_n12849_ = ~new_n12845_ & new_n12848_;
  assign new_n12850_ = new_n12844_ & new_n12849_;
  assign new_n12851_ = new_n12839_ & new_n12850_;
  assign new_n12852_ = new_n6569_ & new_n8670_;
  assign new_n12853_ = new_n6569_ & new_n8655_;
  assign new_n12854_ = new_n6569_ & new_n8667_;
  assign new_n12855_ = ~new_n12853_ & ~new_n12854_;
  assign new_n12856_ = ~new_n12852_ & new_n12855_;
  assign new_n12857_ = new_n6569_ & new_n8681_;
  assign new_n12858_ = new_n6569_ & new_n8665_;
  assign new_n12859_ = new_n6569_ & new_n8678_;
  assign new_n12860_ = ~new_n12858_ & ~new_n12859_;
  assign new_n12861_ = ~new_n12857_ & new_n12860_;
  assign new_n12862_ = new_n12856_ & new_n12861_;
  assign new_n12863_ = new_n6569_ & new_n8694_;
  assign new_n12864_ = new_n6569_ & new_n8675_;
  assign new_n12865_ = new_n6569_ & new_n8692_;
  assign new_n12866_ = ~new_n12864_ & ~new_n12865_;
  assign new_n12867_ = ~new_n12863_ & new_n12866_;
  assign new_n12868_ = new_n6569_ & new_n8689_;
  assign new_n12869_ = new_n6569_ & new_n8699_;
  assign new_n12870_ = ~new_n12868_ & ~new_n12869_;
  assign new_n12871_ = new_n12867_ & new_n12870_;
  assign new_n12872_ = new_n12862_ & new_n12871_;
  assign new_n12873_ = new_n12851_ & new_n12872_;
  assign new_n12874_ = new_n6575_ & new_n8628_;
  assign new_n12875_ = new_n6569_ & new_n8701_;
  assign new_n12876_ = new_n6575_ & new_n8617_;
  assign new_n12877_ = ~new_n12875_ & ~new_n12876_;
  assign new_n12878_ = ~new_n12874_ & new_n12877_;
  assign new_n12879_ = new_n6575_ & new_n8637_;
  assign new_n12880_ = new_n6575_ & new_n8630_;
  assign new_n12881_ = new_n6575_ & new_n8625_;
  assign new_n12882_ = ~new_n12880_ & ~new_n12881_;
  assign new_n12883_ = ~new_n12879_ & new_n12882_;
  assign new_n12884_ = new_n12878_ & new_n12883_;
  assign new_n12885_ = new_n6575_ & new_n8648_;
  assign new_n12886_ = new_n6575_ & new_n8639_;
  assign new_n12887_ = new_n6575_ & new_n8635_;
  assign new_n12888_ = ~new_n12886_ & ~new_n12887_;
  assign new_n12889_ = ~new_n12885_ & new_n12888_;
  assign new_n12890_ = new_n6575_ & new_n8657_;
  assign new_n12891_ = new_n6575_ & new_n8650_;
  assign new_n12892_ = new_n6575_ & new_n8646_;
  assign new_n12893_ = ~new_n12891_ & ~new_n12892_;
  assign new_n12894_ = ~new_n12890_ & new_n12893_;
  assign new_n12895_ = new_n12889_ & new_n12894_;
  assign new_n12896_ = new_n12884_ & new_n12895_;
  assign new_n12897_ = new_n6575_ & new_n8667_;
  assign new_n12898_ = new_n6575_ & new_n8659_;
  assign new_n12899_ = new_n6575_ & new_n8655_;
  assign new_n12900_ = ~new_n12898_ & ~new_n12899_;
  assign new_n12901_ = ~new_n12897_ & new_n12900_;
  assign new_n12902_ = new_n6575_ & new_n8678_;
  assign new_n12903_ = new_n6575_ & new_n8670_;
  assign new_n12904_ = new_n6575_ & new_n8665_;
  assign new_n12905_ = ~new_n12903_ & ~new_n12904_;
  assign new_n12906_ = ~new_n12902_ & new_n12905_;
  assign new_n12907_ = new_n12901_ & new_n12906_;
  assign new_n12908_ = new_n6575_ & new_n8692_;
  assign new_n12909_ = new_n6575_ & new_n8681_;
  assign new_n12910_ = new_n6575_ & new_n8675_;
  assign new_n12911_ = ~new_n12909_ & ~new_n12910_;
  assign new_n12912_ = ~new_n12908_ & new_n12911_;
  assign new_n12913_ = new_n6575_ & new_n8694_;
  assign new_n12914_ = new_n6575_ & new_n8689_;
  assign new_n12915_ = ~new_n12913_ & ~new_n12914_;
  assign new_n12916_ = new_n12912_ & new_n12915_;
  assign new_n12917_ = new_n12907_ & new_n12916_;
  assign new_n12918_ = new_n12896_ & new_n12917_;
  assign new_n12919_ = new_n12873_ & new_n12918_;
  assign new_n12920_ = new_n12828_ & new_n12919_;
  assign new_n12921_ = new_n6583_ & new_n8617_;
  assign new_n12922_ = new_n6575_ & new_n8699_;
  assign new_n12923_ = new_n6575_ & new_n8701_;
  assign new_n12924_ = ~new_n12922_ & ~new_n12923_;
  assign new_n12925_ = ~new_n12921_ & new_n12924_;
  assign new_n12926_ = new_n6583_ & new_n8625_;
  assign new_n12927_ = new_n6583_ & new_n8628_;
  assign new_n12928_ = new_n6583_ & new_n8630_;
  assign new_n12929_ = ~new_n12927_ & ~new_n12928_;
  assign new_n12930_ = ~new_n12926_ & new_n12929_;
  assign new_n12931_ = new_n12925_ & new_n12930_;
  assign new_n12932_ = new_n6583_ & new_n8635_;
  assign new_n12933_ = new_n6583_ & new_n8637_;
  assign new_n12934_ = new_n6583_ & new_n8639_;
  assign new_n12935_ = ~new_n12933_ & ~new_n12934_;
  assign new_n12936_ = ~new_n12932_ & new_n12935_;
  assign new_n12937_ = new_n6583_ & new_n8646_;
  assign new_n12938_ = new_n6583_ & new_n8648_;
  assign new_n12939_ = new_n6583_ & new_n8650_;
  assign new_n12940_ = ~new_n12938_ & ~new_n12939_;
  assign new_n12941_ = ~new_n12937_ & new_n12940_;
  assign new_n12942_ = new_n12936_ & new_n12941_;
  assign new_n12943_ = new_n12931_ & new_n12942_;
  assign new_n12944_ = new_n6583_ & new_n8655_;
  assign new_n12945_ = new_n6583_ & new_n8657_;
  assign new_n12946_ = new_n6583_ & new_n8659_;
  assign new_n12947_ = ~new_n12945_ & ~new_n12946_;
  assign new_n12948_ = ~new_n12944_ & new_n12947_;
  assign new_n12949_ = new_n6583_ & new_n8665_;
  assign new_n12950_ = new_n6583_ & new_n8667_;
  assign new_n12951_ = new_n6583_ & new_n8670_;
  assign new_n12952_ = ~new_n12950_ & ~new_n12951_;
  assign new_n12953_ = ~new_n12949_ & new_n12952_;
  assign new_n12954_ = new_n12948_ & new_n12953_;
  assign new_n12955_ = new_n6583_ & new_n8675_;
  assign new_n12956_ = new_n6583_ & new_n8678_;
  assign new_n12957_ = new_n6583_ & new_n8681_;
  assign new_n12958_ = ~new_n12956_ & ~new_n12957_;
  assign new_n12959_ = ~new_n12955_ & new_n12958_;
  assign new_n12960_ = new_n6583_ & new_n8692_;
  assign new_n12961_ = new_n6583_ & new_n8694_;
  assign new_n12962_ = ~new_n12960_ & ~new_n12961_;
  assign new_n12963_ = new_n12959_ & new_n12962_;
  assign new_n12964_ = new_n12954_ & new_n12963_;
  assign new_n12965_ = new_n12943_ & new_n12964_;
  assign new_n12966_ = new_n6583_ & new_n8701_;
  assign new_n12967_ = new_n6583_ & new_n8689_;
  assign new_n12968_ = new_n6583_ & new_n8699_;
  assign new_n12969_ = ~new_n12967_ & ~new_n12968_;
  assign new_n12970_ = ~new_n12966_ & new_n12969_;
  assign new_n12971_ = new_n6595_ & new_n8630_;
  assign new_n12972_ = new_n6595_ & new_n8617_;
  assign new_n12973_ = new_n6595_ & new_n8628_;
  assign new_n12974_ = ~new_n12972_ & ~new_n12973_;
  assign new_n12975_ = ~new_n12971_ & new_n12974_;
  assign new_n12976_ = new_n12970_ & new_n12975_;
  assign new_n12977_ = new_n6595_ & new_n8639_;
  assign new_n12978_ = new_n6595_ & new_n8625_;
  assign new_n12979_ = new_n6595_ & new_n8637_;
  assign new_n12980_ = ~new_n12978_ & ~new_n12979_;
  assign new_n12981_ = ~new_n12977_ & new_n12980_;
  assign new_n12982_ = new_n6595_ & new_n8650_;
  assign new_n12983_ = new_n6595_ & new_n8635_;
  assign new_n12984_ = new_n6595_ & new_n8648_;
  assign new_n12985_ = ~new_n12983_ & ~new_n12984_;
  assign new_n12986_ = ~new_n12982_ & new_n12985_;
  assign new_n12987_ = new_n12981_ & new_n12986_;
  assign new_n12988_ = new_n12976_ & new_n12987_;
  assign new_n12989_ = new_n6595_ & new_n8659_;
  assign new_n12990_ = new_n6595_ & new_n8646_;
  assign new_n12991_ = new_n6595_ & new_n8657_;
  assign new_n12992_ = ~new_n12990_ & ~new_n12991_;
  assign new_n12993_ = ~new_n12989_ & new_n12992_;
  assign new_n12994_ = new_n6595_ & new_n8670_;
  assign new_n12995_ = new_n6595_ & new_n8655_;
  assign new_n12996_ = new_n6595_ & new_n8667_;
  assign new_n12997_ = ~new_n12995_ & ~new_n12996_;
  assign new_n12998_ = ~new_n12994_ & new_n12997_;
  assign new_n12999_ = new_n12993_ & new_n12998_;
  assign new_n13000_ = new_n6595_ & new_n8681_;
  assign new_n13001_ = new_n6595_ & new_n8665_;
  assign new_n13002_ = new_n6595_ & new_n8678_;
  assign new_n13003_ = ~new_n13001_ & ~new_n13002_;
  assign new_n13004_ = ~new_n13000_ & new_n13003_;
  assign new_n13005_ = new_n6595_ & new_n8675_;
  assign new_n13006_ = new_n6595_ & new_n8692_;
  assign new_n13007_ = ~new_n13005_ & ~new_n13006_;
  assign new_n13008_ = new_n13004_ & new_n13007_;
  assign new_n13009_ = new_n12999_ & new_n13008_;
  assign new_n13010_ = new_n12988_ & new_n13009_;
  assign new_n13011_ = new_n12965_ & new_n13010_;
  assign new_n13012_ = new_n6595_ & new_n8699_;
  assign new_n13013_ = new_n6595_ & new_n8694_;
  assign new_n13014_ = new_n6595_ & new_n8689_;
  assign new_n13015_ = ~new_n13013_ & ~new_n13014_;
  assign new_n13016_ = ~new_n13012_ & new_n13015_;
  assign new_n13017_ = new_n6602_ & new_n8853_;
  assign new_n13018_ = new_n6595_ & new_n8701_;
  assign new_n13019_ = new_n6602_ & new_n8845_;
  assign new_n13020_ = ~new_n13018_ & ~new_n13019_;
  assign new_n13021_ = ~new_n13017_ & new_n13020_;
  assign new_n13022_ = new_n13016_ & new_n13021_;
  assign new_n13023_ = new_n6602_ & new_n8864_;
  assign new_n13024_ = new_n6602_ & new_n8855_;
  assign new_n13025_ = new_n6602_ & new_n8851_;
  assign new_n13026_ = ~new_n13024_ & ~new_n13025_;
  assign new_n13027_ = ~new_n13023_ & new_n13026_;
  assign new_n13028_ = new_n6602_ & new_n8872_;
  assign new_n13029_ = new_n6602_ & new_n8866_;
  assign new_n13030_ = new_n6602_ & new_n8862_;
  assign new_n13031_ = ~new_n13029_ & ~new_n13030_;
  assign new_n13032_ = ~new_n13028_ & new_n13031_;
  assign new_n13033_ = new_n13027_ & new_n13032_;
  assign new_n13034_ = new_n13022_ & new_n13033_;
  assign new_n13035_ = new_n6602_ & new_n8882_;
  assign new_n13036_ = new_n6602_ & new_n8874_;
  assign new_n13037_ = new_n6602_ & new_n8870_;
  assign new_n13038_ = ~new_n13036_ & ~new_n13037_;
  assign new_n13039_ = ~new_n13035_ & new_n13038_;
  assign new_n13040_ = new_n6602_ & new_n8888_;
  assign new_n13041_ = new_n6602_ & new_n8884_;
  assign new_n13042_ = new_n6602_ & new_n8880_;
  assign new_n13043_ = ~new_n13041_ & ~new_n13042_;
  assign new_n13044_ = ~new_n13040_ & new_n13043_;
  assign new_n13045_ = new_n13039_ & new_n13044_;
  assign new_n13046_ = new_n6602_ & new_n8900_;
  assign new_n13047_ = new_n6602_ & new_n8890_;
  assign new_n13048_ = new_n6602_ & new_n8898_;
  assign new_n13049_ = ~new_n13047_ & ~new_n13048_;
  assign new_n13050_ = ~new_n13046_ & new_n13049_;
  assign new_n13051_ = new_n6602_ & new_n8896_;
  assign new_n13052_ = new_n6602_ & new_n8907_;
  assign new_n13053_ = ~new_n13051_ & ~new_n13052_;
  assign new_n13054_ = new_n13050_ & new_n13053_;
  assign new_n13055_ = new_n13045_ & new_n13054_;
  assign new_n13056_ = new_n13034_ & new_n13055_;
  assign new_n13057_ = new_n6602_ & new_n8916_;
  assign new_n13058_ = new_n6602_ & new_n8909_;
  assign new_n13059_ = new_n6602_ & new_n8905_;
  assign new_n13060_ = ~new_n13058_ & ~new_n13059_;
  assign new_n13061_ = ~new_n13057_ & new_n13060_;
  assign new_n13062_ = new_n6602_ & new_n8925_;
  assign new_n13063_ = new_n6602_ & new_n8918_;
  assign new_n13064_ = new_n6602_ & new_n8914_;
  assign new_n13065_ = ~new_n13063_ & ~new_n13064_;
  assign new_n13066_ = ~new_n13062_ & new_n13065_;
  assign new_n13067_ = new_n13061_ & new_n13066_;
  assign new_n13068_ = new_n6602_ & new_n8936_;
  assign new_n13069_ = new_n6602_ & new_n8927_;
  assign new_n13070_ = new_n6602_ & new_n8923_;
  assign new_n13071_ = ~new_n13069_ & ~new_n13070_;
  assign new_n13072_ = ~new_n13068_ & new_n13071_;
  assign new_n13073_ = new_n6602_ & new_n8943_;
  assign new_n13074_ = new_n6602_ & new_n8938_;
  assign new_n13075_ = new_n6602_ & new_n8934_;
  assign new_n13076_ = ~new_n13074_ & ~new_n13075_;
  assign new_n13077_ = ~new_n13073_ & new_n13076_;
  assign new_n13078_ = new_n13072_ & new_n13077_;
  assign new_n13079_ = new_n13067_ & new_n13078_;
  assign new_n13080_ = new_n6655_ & new_n10132_;
  assign new_n13081_ = new_n10131_ & new_n13080_;
  assign new_n13082_ = new_n6602_ & new_n8945_;
  assign new_n13083_ = new_n6655_ & new_n10127_;
  assign new_n13084_ = new_n10125_ & new_n13083_;
  assign new_n13085_ = ~new_n13082_ & ~new_n13084_;
  assign new_n13086_ = ~new_n13081_ & new_n13085_;
  assign new_n13087_ = new_n6655_ & new_n10142_;
  assign new_n13088_ = new_n10125_ & new_n13087_;
  assign new_n13089_ = new_n6655_ & new_n10147_;
  assign new_n13090_ = new_n10146_ & new_n13089_;
  assign new_n13091_ = new_n10151_ & new_n13089_;
  assign new_n13092_ = ~new_n13090_ & ~new_n13091_;
  assign new_n13093_ = ~new_n13088_ & new_n13092_;
  assign new_n13094_ = new_n13086_ & new_n13093_;
  assign new_n13095_ = new_n6655_ & new_n10155_;
  assign new_n13096_ = new_n10151_ & new_n13095_;
  assign new_n13097_ = new_n6655_ & new_n10158_;
  assign new_n13098_ = new_n10131_ & new_n13097_;
  assign new_n13099_ = new_n10146_ & new_n13095_;
  assign new_n13100_ = ~new_n13098_ & ~new_n13099_;
  assign new_n13101_ = ~new_n13096_ & new_n13100_;
  assign new_n13102_ = new_n6655_ & new_n10169_;
  assign new_n13103_ = new_n10125_ & new_n13102_;
  assign new_n13104_ = new_n6655_ & new_n10172_;
  assign new_n13105_ = new_n10131_ & new_n13104_;
  assign new_n13106_ = ~new_n13103_ & ~new_n13105_;
  assign new_n13107_ = new_n13101_ & new_n13106_;
  assign new_n13108_ = new_n13094_ & new_n13107_;
  assign new_n13109_ = new_n13079_ & new_n13108_;
  assign new_n13110_ = new_n13056_ & new_n13109_;
  assign new_n13111_ = new_n13011_ & new_n13110_;
  assign new_n13112_ = new_n12920_ & new_n13111_;
  assign new_n13113_ = new_n12725_ & new_n13112_;
  assign new_n13114_ = new_n12320_ & new_n13113_;
  assign new_n13115_ = new_n11571_ & new_n13114_;
  assign new_n13116_ = new_n9839_ & new_n13115_;
  assign new_n13117_ = new_n6719_ & new_n13116_;
  assign new_n13118_ = new_n6655_ & new_n10181_;
  assign new_n13119_ = new_n10125_ & new_n13118_;
  assign new_n13120_ = new_n6655_ & new_n10166_;
  assign new_n13121_ = new_n10146_ & new_n13120_;
  assign new_n13122_ = new_n10151_ & new_n13120_;
  assign new_n13123_ = ~new_n13121_ & ~new_n13122_;
  assign new_n13124_ = ~new_n13119_ & new_n13123_;
  assign new_n13125_ = new_n6655_ & new_n10189_;
  assign new_n13126_ = new_n10151_ & new_n13125_;
  assign new_n13127_ = new_n6655_ & new_n10177_;
  assign new_n13128_ = new_n10131_ & new_n13127_;
  assign new_n13129_ = new_n10146_ & new_n13125_;
  assign new_n13130_ = ~new_n13128_ & ~new_n13129_;
  assign new_n13131_ = ~new_n13126_ & new_n13130_;
  assign new_n13132_ = new_n13124_ & new_n13131_;
  assign new_n13133_ = new_n6656_ & new_n8630_;
  assign new_n13134_ = new_n6656_ & new_n8617_;
  assign new_n13135_ = new_n6656_ & new_n8628_;
  assign new_n13136_ = ~new_n13134_ & ~new_n13135_;
  assign new_n13137_ = ~new_n13133_ & new_n13136_;
  assign new_n13138_ = new_n6656_ & new_n8639_;
  assign new_n13139_ = new_n6656_ & new_n8625_;
  assign new_n13140_ = new_n6656_ & new_n8637_;
  assign new_n13141_ = ~new_n13139_ & ~new_n13140_;
  assign new_n13142_ = ~new_n13138_ & new_n13141_;
  assign new_n13143_ = new_n13137_ & new_n13142_;
  assign new_n13144_ = new_n13132_ & new_n13143_;
  assign new_n13145_ = new_n6656_ & new_n8650_;
  assign new_n13146_ = new_n6656_ & new_n8635_;
  assign new_n13147_ = new_n6656_ & new_n8648_;
  assign new_n13148_ = ~new_n13146_ & ~new_n13147_;
  assign new_n13149_ = ~new_n13145_ & new_n13148_;
  assign new_n13150_ = new_n6656_ & new_n8659_;
  assign new_n13151_ = new_n6656_ & new_n8646_;
  assign new_n13152_ = new_n6656_ & new_n8657_;
  assign new_n13153_ = ~new_n13151_ & ~new_n13152_;
  assign new_n13154_ = ~new_n13150_ & new_n13153_;
  assign new_n13155_ = new_n13149_ & new_n13154_;
  assign new_n13156_ = new_n6656_ & new_n8670_;
  assign new_n13157_ = new_n6656_ & new_n8655_;
  assign new_n13158_ = new_n6656_ & new_n8667_;
  assign new_n13159_ = ~new_n13157_ & ~new_n13158_;
  assign new_n13160_ = ~new_n13156_ & new_n13159_;
  assign new_n13161_ = new_n6656_ & new_n8681_;
  assign new_n13162_ = new_n6656_ & new_n8665_;
  assign new_n13163_ = new_n6656_ & new_n8678_;
  assign new_n13164_ = ~new_n13162_ & ~new_n13163_;
  assign new_n13165_ = ~new_n13161_ & new_n13164_;
  assign new_n13166_ = new_n13160_ & new_n13165_;
  assign new_n13167_ = new_n13155_ & new_n13166_;
  assign new_n13168_ = new_n13144_ & new_n13167_;
  assign new_n13169_ = new_n6656_ & new_n8694_;
  assign new_n13170_ = new_n6656_ & new_n8675_;
  assign new_n13171_ = new_n6656_ & new_n8692_;
  assign new_n13172_ = ~new_n13170_ & ~new_n13171_;
  assign new_n13173_ = ~new_n13169_ & new_n13172_;
  assign new_n13174_ = new_n6656_ & new_n8701_;
  assign new_n13175_ = new_n6656_ & new_n8689_;
  assign new_n13176_ = new_n6656_ & new_n8699_;
  assign new_n13177_ = ~new_n13175_ & ~new_n13176_;
  assign new_n13178_ = ~new_n13174_ & new_n13177_;
  assign new_n13179_ = new_n13173_ & new_n13178_;
  assign new_n13180_ = new_n6663_ & new_n10241_;
  assign new_n13181_ = new_n10146_ & new_n13180_;
  assign new_n13182_ = new_n6663_ & new_n10244_;
  assign new_n13183_ = new_n10125_ & new_n13182_;
  assign new_n13184_ = new_n6663_ & new_n10247_;
  assign new_n13185_ = new_n10131_ & new_n13184_;
  assign new_n13186_ = ~new_n13183_ & ~new_n13185_;
  assign new_n13187_ = ~new_n13181_ & new_n13186_;
  assign new_n13188_ = new_n6663_ & new_n10254_;
  assign new_n13189_ = new_n10131_ & new_n13188_;
  assign new_n13190_ = new_n10151_ & new_n13180_;
  assign new_n13191_ = new_n6663_ & new_n10258_;
  assign new_n13192_ = new_n10125_ & new_n13191_;
  assign new_n13193_ = ~new_n13190_ & ~new_n13192_;
  assign new_n13194_ = ~new_n13189_ & new_n13193_;
  assign new_n13195_ = new_n13187_ & new_n13194_;
  assign new_n13196_ = new_n13179_ & new_n13195_;
  assign new_n13197_ = new_n6663_ & new_n10276_;
  assign new_n13198_ = new_n10125_ & new_n13197_;
  assign new_n13199_ = new_n6663_ & new_n10263_;
  assign new_n13200_ = new_n10146_ & new_n13199_;
  assign new_n13201_ = new_n10151_ & new_n13199_;
  assign new_n13202_ = ~new_n13200_ & ~new_n13201_;
  assign new_n13203_ = ~new_n13198_ & new_n13202_;
  assign new_n13204_ = new_n6663_ & new_n10273_;
  assign new_n13205_ = new_n10151_ & new_n13204_;
  assign new_n13206_ = new_n6663_ & new_n10279_;
  assign new_n13207_ = new_n10131_ & new_n13206_;
  assign new_n13208_ = new_n10146_ & new_n13204_;
  assign new_n13209_ = ~new_n13207_ & ~new_n13208_;
  assign new_n13210_ = ~new_n13205_ & new_n13209_;
  assign new_n13211_ = new_n13203_ & new_n13210_;
  assign new_n13212_ = new_n6663_ & new_n10295_;
  assign new_n13213_ = new_n10146_ & new_n13212_;
  assign new_n13214_ = new_n6663_ & new_n10288_;
  assign new_n13215_ = new_n10125_ & new_n13214_;
  assign new_n13216_ = new_n6663_ & new_n10284_;
  assign new_n13217_ = new_n10131_ & new_n13216_;
  assign new_n13218_ = ~new_n13215_ & ~new_n13217_;
  assign new_n13219_ = ~new_n13213_ & new_n13218_;
  assign new_n13220_ = new_n10151_ & new_n13212_;
  assign new_n13221_ = new_n6664_ & new_n8617_;
  assign new_n13222_ = ~new_n13220_ & ~new_n13221_;
  assign new_n13223_ = new_n13219_ & new_n13222_;
  assign new_n13224_ = new_n13211_ & new_n13223_;
  assign new_n13225_ = new_n13196_ & new_n13224_;
  assign new_n13226_ = new_n13168_ & new_n13225_;
  assign new_n13227_ = new_n6664_ & new_n8625_;
  assign new_n13228_ = new_n6664_ & new_n8628_;
  assign new_n13229_ = new_n6664_ & new_n8630_;
  assign new_n13230_ = ~new_n13228_ & ~new_n13229_;
  assign new_n13231_ = ~new_n13227_ & new_n13230_;
  assign new_n13232_ = new_n6664_ & new_n8635_;
  assign new_n13233_ = new_n6664_ & new_n8637_;
  assign new_n13234_ = new_n6664_ & new_n8639_;
  assign new_n13235_ = ~new_n13233_ & ~new_n13234_;
  assign new_n13236_ = ~new_n13232_ & new_n13235_;
  assign new_n13237_ = new_n13231_ & new_n13236_;
  assign new_n13238_ = new_n6664_ & new_n8646_;
  assign new_n13239_ = new_n6664_ & new_n8648_;
  assign new_n13240_ = new_n6664_ & new_n8650_;
  assign new_n13241_ = ~new_n13239_ & ~new_n13240_;
  assign new_n13242_ = ~new_n13238_ & new_n13241_;
  assign new_n13243_ = new_n6664_ & new_n8655_;
  assign new_n13244_ = new_n6664_ & new_n8657_;
  assign new_n13245_ = new_n6664_ & new_n8659_;
  assign new_n13246_ = ~new_n13244_ & ~new_n13245_;
  assign new_n13247_ = ~new_n13243_ & new_n13246_;
  assign new_n13248_ = new_n13242_ & new_n13247_;
  assign new_n13249_ = new_n13237_ & new_n13248_;
  assign new_n13250_ = new_n6664_ & new_n8665_;
  assign new_n13251_ = new_n6664_ & new_n8667_;
  assign new_n13252_ = new_n6664_ & new_n8670_;
  assign new_n13253_ = ~new_n13251_ & ~new_n13252_;
  assign new_n13254_ = ~new_n13250_ & new_n13253_;
  assign new_n13255_ = new_n6664_ & new_n8675_;
  assign new_n13256_ = new_n6664_ & new_n8678_;
  assign new_n13257_ = new_n6664_ & new_n8681_;
  assign new_n13258_ = ~new_n13256_ & ~new_n13257_;
  assign new_n13259_ = ~new_n13255_ & new_n13258_;
  assign new_n13260_ = new_n13254_ & new_n13259_;
  assign new_n13261_ = new_n6664_ & new_n8689_;
  assign new_n13262_ = new_n6664_ & new_n8692_;
  assign new_n13263_ = new_n6664_ & new_n8694_;
  assign new_n13264_ = ~new_n13262_ & ~new_n13263_;
  assign new_n13265_ = ~new_n13261_ & new_n13264_;
  assign new_n13266_ = new_n6664_ & new_n8699_;
  assign new_n13267_ = new_n6664_ & new_n8701_;
  assign new_n13268_ = ~new_n13266_ & ~new_n13267_;
  assign new_n13269_ = new_n13265_ & new_n13268_;
  assign new_n13270_ = new_n13260_ & new_n13269_;
  assign new_n13271_ = new_n13249_ & new_n13270_;
  assign new_n13272_ = new_n6672_ & new_n10346_;
  assign new_n13273_ = new_n10146_ & new_n13272_;
  assign new_n13274_ = new_n6672_ & new_n10349_;
  assign new_n13275_ = new_n10125_ & new_n13274_;
  assign new_n13276_ = new_n6672_ & new_n10352_;
  assign new_n13277_ = new_n10131_ & new_n13276_;
  assign new_n13278_ = ~new_n13275_ & ~new_n13277_;
  assign new_n13279_ = ~new_n13273_ & new_n13278_;
  assign new_n13280_ = new_n6672_ & new_n10359_;
  assign new_n13281_ = new_n10131_ & new_n13280_;
  assign new_n13282_ = new_n10151_ & new_n13272_;
  assign new_n13283_ = new_n6672_ & new_n10363_;
  assign new_n13284_ = new_n10125_ & new_n13283_;
  assign new_n13285_ = ~new_n13282_ & ~new_n13284_;
  assign new_n13286_ = ~new_n13281_ & new_n13285_;
  assign new_n13287_ = new_n13279_ & new_n13286_;
  assign new_n13288_ = new_n6672_ & new_n10369_;
  assign new_n13289_ = new_n10125_ & new_n13288_;
  assign new_n13290_ = new_n6672_ & new_n10372_;
  assign new_n13291_ = new_n10146_ & new_n13290_;
  assign new_n13292_ = new_n10151_ & new_n13290_;
  assign new_n13293_ = ~new_n13291_ & ~new_n13292_;
  assign new_n13294_ = ~new_n13289_ & new_n13293_;
  assign new_n13295_ = new_n6672_ & new_n10379_;
  assign new_n13296_ = new_n10151_ & new_n13295_;
  assign new_n13297_ = new_n6672_ & new_n10382_;
  assign new_n13298_ = new_n10131_ & new_n13297_;
  assign new_n13299_ = new_n10146_ & new_n13295_;
  assign new_n13300_ = ~new_n13298_ & ~new_n13299_;
  assign new_n13301_ = ~new_n13296_ & new_n13300_;
  assign new_n13302_ = new_n13294_ & new_n13301_;
  assign new_n13303_ = new_n13287_ & new_n13302_;
  assign new_n13304_ = new_n6672_ & new_n10402_;
  assign new_n13305_ = new_n10146_ & new_n13304_;
  assign new_n13306_ = new_n6672_ & new_n10388_;
  assign new_n13307_ = new_n10125_ & new_n13306_;
  assign new_n13308_ = new_n6672_ & new_n10391_;
  assign new_n13309_ = new_n10131_ & new_n13308_;
  assign new_n13310_ = ~new_n13307_ & ~new_n13309_;
  assign new_n13311_ = ~new_n13305_ & new_n13310_;
  assign new_n13312_ = new_n6673_ & new_n8628_;
  assign new_n13313_ = new_n10151_ & new_n13304_;
  assign new_n13314_ = new_n6673_ & new_n8617_;
  assign new_n13315_ = ~new_n13313_ & ~new_n13314_;
  assign new_n13316_ = ~new_n13312_ & new_n13315_;
  assign new_n13317_ = new_n13311_ & new_n13316_;
  assign new_n13318_ = new_n6673_ & new_n8637_;
  assign new_n13319_ = new_n6673_ & new_n8630_;
  assign new_n13320_ = new_n6673_ & new_n8625_;
  assign new_n13321_ = ~new_n13319_ & ~new_n13320_;
  assign new_n13322_ = ~new_n13318_ & new_n13321_;
  assign new_n13323_ = new_n6673_ & new_n8639_;
  assign new_n13324_ = new_n6673_ & new_n8635_;
  assign new_n13325_ = ~new_n13323_ & ~new_n13324_;
  assign new_n13326_ = new_n13322_ & new_n13325_;
  assign new_n13327_ = new_n13317_ & new_n13326_;
  assign new_n13328_ = new_n13303_ & new_n13327_;
  assign new_n13329_ = new_n13271_ & new_n13328_;
  assign new_n13330_ = new_n13226_ & new_n13329_;
  assign new_n13331_ = new_n6673_ & new_n8646_;
  assign new_n13332_ = new_n6673_ & new_n8648_;
  assign new_n13333_ = new_n6673_ & new_n8650_;
  assign new_n13334_ = ~new_n13332_ & ~new_n13333_;
  assign new_n13335_ = ~new_n13331_ & new_n13334_;
  assign new_n13336_ = new_n6673_ & new_n8655_;
  assign new_n13337_ = new_n6673_ & new_n8657_;
  assign new_n13338_ = new_n6673_ & new_n8659_;
  assign new_n13339_ = ~new_n13337_ & ~new_n13338_;
  assign new_n13340_ = ~new_n13336_ & new_n13339_;
  assign new_n13341_ = new_n13335_ & new_n13340_;
  assign new_n13342_ = new_n6673_ & new_n8665_;
  assign new_n13343_ = new_n6673_ & new_n8667_;
  assign new_n13344_ = new_n6673_ & new_n8670_;
  assign new_n13345_ = ~new_n13343_ & ~new_n13344_;
  assign new_n13346_ = ~new_n13342_ & new_n13345_;
  assign new_n13347_ = new_n6673_ & new_n8675_;
  assign new_n13348_ = new_n6673_ & new_n8678_;
  assign new_n13349_ = new_n6673_ & new_n8681_;
  assign new_n13350_ = ~new_n13348_ & ~new_n13349_;
  assign new_n13351_ = ~new_n13347_ & new_n13350_;
  assign new_n13352_ = new_n13346_ & new_n13351_;
  assign new_n13353_ = new_n13341_ & new_n13352_;
  assign new_n13354_ = new_n6673_ & new_n8689_;
  assign new_n13355_ = new_n6673_ & new_n8692_;
  assign new_n13356_ = new_n6673_ & new_n8694_;
  assign new_n13357_ = ~new_n13355_ & ~new_n13356_;
  assign new_n13358_ = ~new_n13354_ & new_n13357_;
  assign new_n13359_ = new_n6672_ & new_n10450_;
  assign new_n13360_ = new_n10125_ & new_n13359_;
  assign new_n13361_ = new_n6673_ & new_n8699_;
  assign new_n13362_ = new_n6673_ & new_n8701_;
  assign new_n13363_ = ~new_n13361_ & ~new_n13362_;
  assign new_n13364_ = ~new_n13360_ & new_n13363_;
  assign new_n13365_ = new_n13358_ & new_n13364_;
  assign new_n13366_ = new_n6672_ & new_n10457_;
  assign new_n13367_ = new_n10151_ & new_n13366_;
  assign new_n13368_ = new_n6672_ & new_n10460_;
  assign new_n13369_ = new_n10131_ & new_n13368_;
  assign new_n13370_ = new_n10146_ & new_n13366_;
  assign new_n13371_ = ~new_n13369_ & ~new_n13370_;
  assign new_n13372_ = ~new_n13367_ & new_n13371_;
  assign new_n13373_ = new_n6672_ & new_n10470_;
  assign new_n13374_ = new_n10125_ & new_n13373_;
  assign new_n13375_ = new_n6672_ & new_n10473_;
  assign new_n13376_ = new_n10131_ & new_n13375_;
  assign new_n13377_ = ~new_n13374_ & ~new_n13376_;
  assign new_n13378_ = new_n13372_ & new_n13377_;
  assign new_n13379_ = new_n13365_ & new_n13378_;
  assign new_n13380_ = new_n13353_ & new_n13379_;
  assign new_n13381_ = new_n6672_ & new_n10483_;
  assign new_n13382_ = new_n10125_ & new_n13381_;
  assign new_n13383_ = new_n6672_ & new_n10467_;
  assign new_n13384_ = new_n10146_ & new_n13383_;
  assign new_n13385_ = new_n10151_ & new_n13383_;
  assign new_n13386_ = ~new_n13384_ & ~new_n13385_;
  assign new_n13387_ = ~new_n13382_ & new_n13386_;
  assign new_n13388_ = new_n6672_ & new_n10493_;
  assign new_n13389_ = new_n10151_ & new_n13388_;
  assign new_n13390_ = new_n6672_ & new_n10479_;
  assign new_n13391_ = new_n10131_ & new_n13390_;
  assign new_n13392_ = new_n10146_ & new_n13388_;
  assign new_n13393_ = ~new_n13391_ & ~new_n13392_;
  assign new_n13394_ = ~new_n13389_ & new_n13393_;
  assign new_n13395_ = new_n13387_ & new_n13394_;
  assign new_n13396_ = new_n6672_ & new_n10499_;
  assign new_n13397_ = new_n10146_ & new_n13396_;
  assign new_n13398_ = new_n6672_ & new_n10490_;
  assign new_n13399_ = new_n10125_ & new_n13398_;
  assign new_n13400_ = new_n6672_ & new_n10502_;
  assign new_n13401_ = new_n10131_ & new_n13400_;
  assign new_n13402_ = ~new_n13399_ & ~new_n13401_;
  assign new_n13403_ = ~new_n13397_ & new_n13402_;
  assign new_n13404_ = new_n6686_ & new_n8628_;
  assign new_n13405_ = new_n10151_ & new_n13396_;
  assign new_n13406_ = new_n6686_ & new_n8617_;
  assign new_n13407_ = ~new_n13405_ & ~new_n13406_;
  assign new_n13408_ = ~new_n13404_ & new_n13407_;
  assign new_n13409_ = new_n13403_ & new_n13408_;
  assign new_n13410_ = new_n13395_ & new_n13409_;
  assign new_n13411_ = new_n6686_ & new_n8637_;
  assign new_n13412_ = new_n6686_ & new_n8630_;
  assign new_n13413_ = new_n6686_ & new_n8625_;
  assign new_n13414_ = ~new_n13412_ & ~new_n13413_;
  assign new_n13415_ = ~new_n13411_ & new_n13414_;
  assign new_n13416_ = new_n6686_ & new_n8648_;
  assign new_n13417_ = new_n6686_ & new_n8639_;
  assign new_n13418_ = new_n6686_ & new_n8635_;
  assign new_n13419_ = ~new_n13417_ & ~new_n13418_;
  assign new_n13420_ = ~new_n13416_ & new_n13419_;
  assign new_n13421_ = new_n13415_ & new_n13420_;
  assign new_n13422_ = new_n6686_ & new_n8657_;
  assign new_n13423_ = new_n6686_ & new_n8650_;
  assign new_n13424_ = new_n6686_ & new_n8646_;
  assign new_n13425_ = ~new_n13423_ & ~new_n13424_;
  assign new_n13426_ = ~new_n13422_ & new_n13425_;
  assign new_n13427_ = new_n6686_ & new_n8659_;
  assign new_n13428_ = new_n6686_ & new_n8655_;
  assign new_n13429_ = ~new_n13427_ & ~new_n13428_;
  assign new_n13430_ = new_n13426_ & new_n13429_;
  assign new_n13431_ = new_n13421_ & new_n13430_;
  assign new_n13432_ = new_n13410_ & new_n13431_;
  assign new_n13433_ = new_n13380_ & new_n13432_;
  assign new_n13434_ = new_n6686_ & new_n8665_;
  assign new_n13435_ = new_n6686_ & new_n8667_;
  assign new_n13436_ = new_n6686_ & new_n8670_;
  assign new_n13437_ = ~new_n13435_ & ~new_n13436_;
  assign new_n13438_ = ~new_n13434_ & new_n13437_;
  assign new_n13439_ = new_n6686_ & new_n8675_;
  assign new_n13440_ = new_n6686_ & new_n8678_;
  assign new_n13441_ = new_n6686_ & new_n8681_;
  assign new_n13442_ = ~new_n13440_ & ~new_n13441_;
  assign new_n13443_ = ~new_n13439_ & new_n13442_;
  assign new_n13444_ = new_n13438_ & new_n13443_;
  assign new_n13445_ = new_n6686_ & new_n8689_;
  assign new_n13446_ = new_n6686_ & new_n8692_;
  assign new_n13447_ = new_n6686_ & new_n8694_;
  assign new_n13448_ = ~new_n13446_ & ~new_n13447_;
  assign new_n13449_ = ~new_n13445_ & new_n13448_;
  assign new_n13450_ = new_n6694_ & new_n8617_;
  assign new_n13451_ = new_n6686_ & new_n8699_;
  assign new_n13452_ = new_n6686_ & new_n8701_;
  assign new_n13453_ = ~new_n13451_ & ~new_n13452_;
  assign new_n13454_ = ~new_n13450_ & new_n13453_;
  assign new_n13455_ = new_n13449_ & new_n13454_;
  assign new_n13456_ = new_n13444_ & new_n13455_;
  assign new_n13457_ = new_n6694_ & new_n8625_;
  assign new_n13458_ = new_n6694_ & new_n8628_;
  assign new_n13459_ = new_n6694_ & new_n8630_;
  assign new_n13460_ = ~new_n13458_ & ~new_n13459_;
  assign new_n13461_ = ~new_n13457_ & new_n13460_;
  assign new_n13462_ = new_n6694_ & new_n8635_;
  assign new_n13463_ = new_n6694_ & new_n8637_;
  assign new_n13464_ = new_n6694_ & new_n8639_;
  assign new_n13465_ = ~new_n13463_ & ~new_n13464_;
  assign new_n13466_ = ~new_n13462_ & new_n13465_;
  assign new_n13467_ = new_n13461_ & new_n13466_;
  assign new_n13468_ = new_n6694_ & new_n8646_;
  assign new_n13469_ = new_n6694_ & new_n8648_;
  assign new_n13470_ = new_n6694_ & new_n8650_;
  assign new_n13471_ = ~new_n13469_ & ~new_n13470_;
  assign new_n13472_ = ~new_n13468_ & new_n13471_;
  assign new_n13473_ = new_n6694_ & new_n8657_;
  assign new_n13474_ = new_n6694_ & new_n8659_;
  assign new_n13475_ = ~new_n13473_ & ~new_n13474_;
  assign new_n13476_ = new_n13472_ & new_n13475_;
  assign new_n13477_ = new_n13467_ & new_n13476_;
  assign new_n13478_ = new_n13456_ & new_n13477_;
  assign new_n13479_ = new_n6694_ & new_n8670_;
  assign new_n13480_ = new_n6694_ & new_n8655_;
  assign new_n13481_ = new_n6694_ & new_n8667_;
  assign new_n13482_ = ~new_n13480_ & ~new_n13481_;
  assign new_n13483_ = ~new_n13479_ & new_n13482_;
  assign new_n13484_ = new_n6694_ & new_n8681_;
  assign new_n13485_ = new_n6694_ & new_n8665_;
  assign new_n13486_ = new_n6694_ & new_n8678_;
  assign new_n13487_ = ~new_n13485_ & ~new_n13486_;
  assign new_n13488_ = ~new_n13484_ & new_n13487_;
  assign new_n13489_ = new_n13483_ & new_n13488_;
  assign new_n13490_ = new_n6694_ & new_n8694_;
  assign new_n13491_ = new_n6694_ & new_n8675_;
  assign new_n13492_ = new_n6694_ & new_n8692_;
  assign new_n13493_ = ~new_n13491_ & ~new_n13492_;
  assign new_n13494_ = ~new_n13490_ & new_n13493_;
  assign new_n13495_ = new_n6694_ & new_n8701_;
  assign new_n13496_ = new_n6694_ & new_n8689_;
  assign new_n13497_ = new_n6694_ & new_n8699_;
  assign new_n13498_ = ~new_n13496_ & ~new_n13497_;
  assign new_n13499_ = ~new_n13495_ & new_n13498_;
  assign new_n13500_ = new_n13494_ & new_n13499_;
  assign new_n13501_ = new_n13489_ & new_n13500_;
  assign new_n13502_ = new_n6701_ & new_n8630_;
  assign new_n13503_ = new_n6701_ & new_n8617_;
  assign new_n13504_ = new_n6701_ & new_n8628_;
  assign new_n13505_ = ~new_n13503_ & ~new_n13504_;
  assign new_n13506_ = ~new_n13502_ & new_n13505_;
  assign new_n13507_ = new_n6701_ & new_n8639_;
  assign new_n13508_ = new_n6701_ & new_n8625_;
  assign new_n13509_ = new_n6701_ & new_n8637_;
  assign new_n13510_ = ~new_n13508_ & ~new_n13509_;
  assign new_n13511_ = ~new_n13507_ & new_n13510_;
  assign new_n13512_ = new_n13506_ & new_n13511_;
  assign new_n13513_ = new_n6701_ & new_n8650_;
  assign new_n13514_ = new_n6701_ & new_n8635_;
  assign new_n13515_ = new_n6701_ & new_n8648_;
  assign new_n13516_ = ~new_n13514_ & ~new_n13515_;
  assign new_n13517_ = ~new_n13513_ & new_n13516_;
  assign new_n13518_ = new_n6701_ & new_n8646_;
  assign new_n13519_ = new_n6701_ & new_n8657_;
  assign new_n13520_ = ~new_n13518_ & ~new_n13519_;
  assign new_n13521_ = new_n13517_ & new_n13520_;
  assign new_n13522_ = new_n13512_ & new_n13521_;
  assign new_n13523_ = new_n13501_ & new_n13522_;
  assign new_n13524_ = new_n13478_ & new_n13523_;
  assign new_n13525_ = new_n13433_ & new_n13524_;
  assign new_n13526_ = new_n13330_ & new_n13525_;
  assign new_n13527_ = new_n6701_ & new_n8667_;
  assign new_n13528_ = new_n6701_ & new_n8659_;
  assign new_n13529_ = new_n6701_ & new_n8655_;
  assign new_n13530_ = ~new_n13528_ & ~new_n13529_;
  assign new_n13531_ = ~new_n13527_ & new_n13530_;
  assign new_n13532_ = new_n6701_ & new_n8678_;
  assign new_n13533_ = new_n6701_ & new_n8670_;
  assign new_n13534_ = new_n6701_ & new_n8665_;
  assign new_n13535_ = ~new_n13533_ & ~new_n13534_;
  assign new_n13536_ = ~new_n13532_ & new_n13535_;
  assign new_n13537_ = new_n13531_ & new_n13536_;
  assign new_n13538_ = new_n6701_ & new_n8692_;
  assign new_n13539_ = new_n6701_ & new_n8681_;
  assign new_n13540_ = new_n6701_ & new_n8675_;
  assign new_n13541_ = ~new_n13539_ & ~new_n13540_;
  assign new_n13542_ = ~new_n13538_ & new_n13541_;
  assign new_n13543_ = new_n6701_ & new_n8699_;
  assign new_n13544_ = new_n6701_ & new_n8694_;
  assign new_n13545_ = new_n6701_ & new_n8689_;
  assign new_n13546_ = ~new_n13544_ & ~new_n13545_;
  assign new_n13547_ = ~new_n13543_ & new_n13546_;
  assign new_n13548_ = new_n13542_ & new_n13547_;
  assign new_n13549_ = new_n13537_ & new_n13548_;
  assign new_n13550_ = new_n6720_ & new_n8628_;
  assign new_n13551_ = new_n6701_ & new_n8701_;
  assign new_n13552_ = new_n6720_ & new_n8617_;
  assign new_n13553_ = ~new_n13551_ & ~new_n13552_;
  assign new_n13554_ = ~new_n13550_ & new_n13553_;
  assign new_n13555_ = new_n6720_ & new_n8637_;
  assign new_n13556_ = new_n6720_ & new_n8630_;
  assign new_n13557_ = new_n6720_ & new_n8625_;
  assign new_n13558_ = ~new_n13556_ & ~new_n13557_;
  assign new_n13559_ = ~new_n13555_ & new_n13558_;
  assign new_n13560_ = new_n13554_ & new_n13559_;
  assign new_n13561_ = new_n6720_ & new_n8648_;
  assign new_n13562_ = new_n6720_ & new_n8639_;
  assign new_n13563_ = new_n6720_ & new_n8635_;
  assign new_n13564_ = ~new_n13562_ & ~new_n13563_;
  assign new_n13565_ = ~new_n13561_ & new_n13564_;
  assign new_n13566_ = new_n6720_ & new_n8657_;
  assign new_n13567_ = new_n6720_ & new_n8650_;
  assign new_n13568_ = new_n6720_ & new_n8646_;
  assign new_n13569_ = ~new_n13567_ & ~new_n13568_;
  assign new_n13570_ = ~new_n13566_ & new_n13569_;
  assign new_n13571_ = new_n13565_ & new_n13570_;
  assign new_n13572_ = new_n13560_ & new_n13571_;
  assign new_n13573_ = new_n13549_ & new_n13572_;
  assign new_n13574_ = new_n6720_ & new_n8667_;
  assign new_n13575_ = new_n6720_ & new_n8659_;
  assign new_n13576_ = new_n6720_ & new_n8655_;
  assign new_n13577_ = ~new_n13575_ & ~new_n13576_;
  assign new_n13578_ = ~new_n13574_ & new_n13577_;
  assign new_n13579_ = new_n6720_ & new_n8678_;
  assign new_n13580_ = new_n6720_ & new_n8670_;
  assign new_n13581_ = new_n6720_ & new_n8665_;
  assign new_n13582_ = ~new_n13580_ & ~new_n13581_;
  assign new_n13583_ = ~new_n13579_ & new_n13582_;
  assign new_n13584_ = new_n13578_ & new_n13583_;
  assign new_n13585_ = new_n6720_ & new_n8692_;
  assign new_n13586_ = new_n6720_ & new_n8681_;
  assign new_n13587_ = new_n6720_ & new_n8675_;
  assign new_n13588_ = ~new_n13586_ & ~new_n13587_;
  assign new_n13589_ = ~new_n13585_ & new_n13588_;
  assign new_n13590_ = new_n6720_ & new_n8699_;
  assign new_n13591_ = new_n6720_ & new_n8694_;
  assign new_n13592_ = new_n6720_ & new_n8689_;
  assign new_n13593_ = ~new_n13591_ & ~new_n13592_;
  assign new_n13594_ = ~new_n13590_ & new_n13593_;
  assign new_n13595_ = new_n13589_ & new_n13594_;
  assign new_n13596_ = new_n13584_ & new_n13595_;
  assign new_n13597_ = new_n6726_ & new_n8628_;
  assign new_n13598_ = new_n6720_ & new_n8701_;
  assign new_n13599_ = new_n6726_ & new_n8617_;
  assign new_n13600_ = ~new_n13598_ & ~new_n13599_;
  assign new_n13601_ = ~new_n13597_ & new_n13600_;
  assign new_n13602_ = new_n6726_ & new_n8637_;
  assign new_n13603_ = new_n6726_ & new_n8630_;
  assign new_n13604_ = new_n6726_ & new_n8625_;
  assign new_n13605_ = ~new_n13603_ & ~new_n13604_;
  assign new_n13606_ = ~new_n13602_ & new_n13605_;
  assign new_n13607_ = new_n13601_ & new_n13606_;
  assign new_n13608_ = new_n6726_ & new_n8648_;
  assign new_n13609_ = new_n6726_ & new_n8639_;
  assign new_n13610_ = new_n6726_ & new_n8635_;
  assign new_n13611_ = ~new_n13609_ & ~new_n13610_;
  assign new_n13612_ = ~new_n13608_ & new_n13611_;
  assign new_n13613_ = new_n6726_ & new_n8650_;
  assign new_n13614_ = new_n6726_ & new_n8646_;
  assign new_n13615_ = ~new_n13613_ & ~new_n13614_;
  assign new_n13616_ = new_n13612_ & new_n13615_;
  assign new_n13617_ = new_n13607_ & new_n13616_;
  assign new_n13618_ = new_n13596_ & new_n13617_;
  assign new_n13619_ = new_n13573_ & new_n13618_;
  assign new_n13620_ = new_n6726_ & new_n8655_;
  assign new_n13621_ = new_n6726_ & new_n8657_;
  assign new_n13622_ = new_n6726_ & new_n8659_;
  assign new_n13623_ = ~new_n13621_ & ~new_n13622_;
  assign new_n13624_ = ~new_n13620_ & new_n13623_;
  assign new_n13625_ = new_n6726_ & new_n8665_;
  assign new_n13626_ = new_n6726_ & new_n8667_;
  assign new_n13627_ = new_n6726_ & new_n8670_;
  assign new_n13628_ = ~new_n13626_ & ~new_n13627_;
  assign new_n13629_ = ~new_n13625_ & new_n13628_;
  assign new_n13630_ = new_n13624_ & new_n13629_;
  assign new_n13631_ = new_n6726_ & new_n8675_;
  assign new_n13632_ = new_n6726_ & new_n8678_;
  assign new_n13633_ = new_n6726_ & new_n8681_;
  assign new_n13634_ = ~new_n13632_ & ~new_n13633_;
  assign new_n13635_ = ~new_n13631_ & new_n13634_;
  assign new_n13636_ = new_n6726_ & new_n8689_;
  assign new_n13637_ = new_n6726_ & new_n8692_;
  assign new_n13638_ = new_n6726_ & new_n8694_;
  assign new_n13639_ = ~new_n13637_ & ~new_n13638_;
  assign new_n13640_ = ~new_n13636_ & new_n13639_;
  assign new_n13641_ = new_n13635_ & new_n13640_;
  assign new_n13642_ = new_n13630_ & new_n13641_;
  assign new_n13643_ = new_n6738_ & new_n8845_;
  assign new_n13644_ = new_n6726_ & new_n8699_;
  assign new_n13645_ = new_n6726_ & new_n8701_;
  assign new_n13646_ = ~new_n13644_ & ~new_n13645_;
  assign new_n13647_ = ~new_n13643_ & new_n13646_;
  assign new_n13648_ = new_n6738_ & new_n8851_;
  assign new_n13649_ = new_n6738_ & new_n8853_;
  assign new_n13650_ = new_n6738_ & new_n8855_;
  assign new_n13651_ = ~new_n13649_ & ~new_n13650_;
  assign new_n13652_ = ~new_n13648_ & new_n13651_;
  assign new_n13653_ = new_n13647_ & new_n13652_;
  assign new_n13654_ = new_n6738_ & new_n8862_;
  assign new_n13655_ = new_n6738_ & new_n8864_;
  assign new_n13656_ = new_n6738_ & new_n8866_;
  assign new_n13657_ = ~new_n13655_ & ~new_n13656_;
  assign new_n13658_ = ~new_n13654_ & new_n13657_;
  assign new_n13659_ = new_n6738_ & new_n8872_;
  assign new_n13660_ = new_n6738_ & new_n8874_;
  assign new_n13661_ = ~new_n13659_ & ~new_n13660_;
  assign new_n13662_ = new_n13658_ & new_n13661_;
  assign new_n13663_ = new_n13653_ & new_n13662_;
  assign new_n13664_ = new_n13642_ & new_n13663_;
  assign new_n13665_ = new_n6738_ & new_n8884_;
  assign new_n13666_ = new_n6738_ & new_n8870_;
  assign new_n13667_ = new_n6738_ & new_n8882_;
  assign new_n13668_ = ~new_n13666_ & ~new_n13667_;
  assign new_n13669_ = ~new_n13665_ & new_n13668_;
  assign new_n13670_ = new_n6738_ & new_n8890_;
  assign new_n13671_ = new_n6738_ & new_n8880_;
  assign new_n13672_ = new_n6738_ & new_n8888_;
  assign new_n13673_ = ~new_n13671_ & ~new_n13672_;
  assign new_n13674_ = ~new_n13670_ & new_n13673_;
  assign new_n13675_ = new_n13669_ & new_n13674_;
  assign new_n13676_ = new_n6738_ & new_n8896_;
  assign new_n13677_ = new_n6738_ & new_n8898_;
  assign new_n13678_ = new_n6738_ & new_n8900_;
  assign new_n13679_ = ~new_n13677_ & ~new_n13678_;
  assign new_n13680_ = ~new_n13676_ & new_n13679_;
  assign new_n13681_ = new_n6738_ & new_n8905_;
  assign new_n13682_ = new_n6738_ & new_n8907_;
  assign new_n13683_ = new_n6738_ & new_n8909_;
  assign new_n13684_ = ~new_n13682_ & ~new_n13683_;
  assign new_n13685_ = ~new_n13681_ & new_n13684_;
  assign new_n13686_ = new_n13680_ & new_n13685_;
  assign new_n13687_ = new_n13675_ & new_n13686_;
  assign new_n13688_ = new_n6738_ & new_n8914_;
  assign new_n13689_ = new_n6738_ & new_n8916_;
  assign new_n13690_ = new_n6738_ & new_n8918_;
  assign new_n13691_ = ~new_n13689_ & ~new_n13690_;
  assign new_n13692_ = ~new_n13688_ & new_n13691_;
  assign new_n13693_ = new_n6738_ & new_n8923_;
  assign new_n13694_ = new_n6738_ & new_n8925_;
  assign new_n13695_ = new_n6738_ & new_n8927_;
  assign new_n13696_ = ~new_n13694_ & ~new_n13695_;
  assign new_n13697_ = ~new_n13693_ & new_n13696_;
  assign new_n13698_ = new_n13692_ & new_n13697_;
  assign new_n13699_ = new_n6738_ & new_n8934_;
  assign new_n13700_ = new_n6738_ & new_n8936_;
  assign new_n13701_ = new_n6738_ & new_n8938_;
  assign new_n13702_ = ~new_n13700_ & ~new_n13701_;
  assign new_n13703_ = ~new_n13699_ & new_n13702_;
  assign new_n13704_ = new_n6738_ & new_n8943_;
  assign new_n13705_ = new_n6738_ & new_n8945_;
  assign new_n13706_ = ~new_n13704_ & ~new_n13705_;
  assign new_n13707_ = new_n13703_ & new_n13706_;
  assign new_n13708_ = new_n13698_ & new_n13707_;
  assign new_n13709_ = new_n13687_ & new_n13708_;
  assign new_n13710_ = new_n13664_ & new_n13709_;
  assign new_n13711_ = new_n13619_ & new_n13710_;
  assign new_n13712_ = new_n7115_ & new_n9924_;
  assign new_n13713_ = new_n7115_ & new_n9926_;
  assign new_n13714_ = new_n7115_ & new_n9928_;
  assign new_n13715_ = ~new_n13713_ & ~new_n13714_;
  assign new_n13716_ = ~new_n13712_ & new_n13715_;
  assign new_n13717_ = new_n7115_ & new_n9934_;
  assign new_n13718_ = new_n7115_ & new_n9936_;
  assign new_n13719_ = new_n7115_ & new_n9938_;
  assign new_n13720_ = ~new_n13718_ & ~new_n13719_;
  assign new_n13721_ = ~new_n13717_ & new_n13720_;
  assign new_n13722_ = new_n13716_ & new_n13721_;
  assign new_n13723_ = new_n7115_ & new_n9942_;
  assign new_n13724_ = new_n7115_ & new_n9944_;
  assign new_n13725_ = new_n7115_ & new_n9946_;
  assign new_n13726_ = ~new_n13724_ & ~new_n13725_;
  assign new_n13727_ = ~new_n13723_ & new_n13726_;
  assign new_n13728_ = new_n7115_ & new_n9952_;
  assign new_n13729_ = new_n7115_ & new_n9954_;
  assign new_n13730_ = new_n7115_ & new_n9956_;
  assign new_n13731_ = ~new_n13729_ & ~new_n13730_;
  assign new_n13732_ = ~new_n13728_ & new_n13731_;
  assign new_n13733_ = new_n13727_ & new_n13732_;
  assign new_n13734_ = new_n13722_ & new_n13733_;
  assign new_n13735_ = new_n7115_ & new_n9961_;
  assign new_n13736_ = new_n7115_ & new_n9963_;
  assign new_n13737_ = new_n7115_ & new_n9965_;
  assign new_n13738_ = ~new_n13736_ & ~new_n13737_;
  assign new_n13739_ = ~new_n13735_ & new_n13738_;
  assign new_n13740_ = new_n7115_ & new_n9970_;
  assign new_n13741_ = new_n7115_ & new_n9972_;
  assign new_n13742_ = new_n7115_ & new_n9974_;
  assign new_n13743_ = ~new_n13741_ & ~new_n13742_;
  assign new_n13744_ = ~new_n13740_ & new_n13743_;
  assign new_n13745_ = new_n13739_ & new_n13744_;
  assign new_n13746_ = new_n7115_ & new_n9990_;
  assign new_n13747_ = new_n7115_ & new_n9978_;
  assign new_n13748_ = new_n7115_ & new_n9980_;
  assign new_n13749_ = ~new_n13747_ & ~new_n13748_;
  assign new_n13750_ = ~new_n13746_ & new_n13749_;
  assign new_n13751_ = new_n7115_ & new_n9992_;
  assign new_n13752_ = new_n7115_ & new_n9988_;
  assign new_n13753_ = ~new_n13751_ & ~new_n13752_;
  assign new_n13754_ = new_n13750_ & new_n13753_;
  assign new_n13755_ = new_n13745_ & new_n13754_;
  assign new_n13756_ = new_n13734_ & new_n13755_;
  assign new_n13757_ = new_n7115_ & new_n9997_;
  assign new_n13758_ = new_n7115_ & new_n9999_;
  assign new_n13759_ = new_n7115_ & new_n10001_;
  assign new_n13760_ = ~new_n13758_ & ~new_n13759_;
  assign new_n13761_ = ~new_n13757_ & new_n13760_;
  assign new_n13762_ = new_n7115_ & new_n10007_;
  assign new_n13763_ = new_n7115_ & new_n10009_;
  assign new_n13764_ = new_n7115_ & new_n10011_;
  assign new_n13765_ = ~new_n13763_ & ~new_n13764_;
  assign new_n13766_ = ~new_n13762_ & new_n13765_;
  assign new_n13767_ = new_n13761_ & new_n13766_;
  assign new_n13768_ = new_n7115_ & new_n10015_;
  assign new_n13769_ = new_n7115_ & new_n10017_;
  assign new_n13770_ = new_n7115_ & new_n10019_;
  assign new_n13771_ = ~new_n13769_ & ~new_n13770_;
  assign new_n13772_ = ~new_n13768_ & new_n13771_;
  assign new_n13773_ = new_n7115_ & new_n10026_;
  assign new_n13774_ = new_n7115_ & new_n10028_;
  assign new_n13775_ = new_n7115_ & new_n10030_;
  assign new_n13776_ = ~new_n13774_ & ~new_n13775_;
  assign new_n13777_ = ~new_n13773_ & new_n13776_;
  assign new_n13778_ = new_n13772_ & new_n13777_;
  assign new_n13779_ = new_n13767_ & new_n13778_;
  assign new_n13780_ = new_n7115_ & new_n10035_;
  assign new_n13781_ = new_n7115_ & new_n10037_;
  assign new_n13782_ = new_n7115_ & new_n10039_;
  assign new_n13783_ = ~new_n13781_ & ~new_n13782_;
  assign new_n13784_ = ~new_n13780_ & new_n13783_;
  assign new_n13785_ = new_n7115_ & new_n10044_;
  assign new_n13786_ = new_n7115_ & new_n10046_;
  assign new_n13787_ = new_n7115_ & new_n10048_;
  assign new_n13788_ = ~new_n13786_ & ~new_n13787_;
  assign new_n13789_ = ~new_n13785_ & new_n13788_;
  assign new_n13790_ = new_n13784_ & new_n13789_;
  assign new_n13791_ = new_n7115_ & new_n10063_;
  assign new_n13792_ = new_n7115_ & new_n10052_;
  assign new_n13793_ = new_n7115_ & new_n10054_;
  assign new_n13794_ = ~new_n13792_ & ~new_n13793_;
  assign new_n13795_ = ~new_n13791_ & new_n13794_;
  assign new_n13796_ = new_n7115_ & new_n10065_;
  assign new_n13797_ = new_n7115_ & new_n10061_;
  assign new_n13798_ = ~new_n13796_ & ~new_n13797_;
  assign new_n13799_ = new_n13795_ & new_n13798_;
  assign new_n13800_ = new_n13790_ & new_n13799_;
  assign new_n13801_ = new_n13779_ & new_n13800_;
  assign new_n13802_ = new_n13756_ & new_n13801_;
  assign new_n13803_ = new_n7115_ & new_n10069_;
  assign new_n13804_ = new_n7115_ & new_n10071_;
  assign new_n13805_ = new_n7115_ & new_n10073_;
  assign new_n13806_ = ~new_n13804_ & ~new_n13805_;
  assign new_n13807_ = ~new_n13803_ & new_n13806_;
  assign new_n13808_ = new_n7115_ & new_n10078_;
  assign new_n13809_ = new_n7115_ & new_n10080_;
  assign new_n13810_ = new_n7115_ & new_n10082_;
  assign new_n13811_ = ~new_n13809_ & ~new_n13810_;
  assign new_n13812_ = ~new_n13808_ & new_n13811_;
  assign new_n13813_ = new_n13807_ & new_n13812_;
  assign new_n13814_ = new_n7115_ & new_n10087_;
  assign new_n13815_ = new_n7115_ & new_n10089_;
  assign new_n13816_ = new_n7115_ & new_n10091_;
  assign new_n13817_ = ~new_n13815_ & ~new_n13816_;
  assign new_n13818_ = ~new_n13814_ & new_n13817_;
  assign new_n13819_ = new_n7115_ & new_n10098_;
  assign new_n13820_ = new_n7115_ & new_n10100_;
  assign new_n13821_ = new_n7115_ & new_n10102_;
  assign new_n13822_ = ~new_n13820_ & ~new_n13821_;
  assign new_n13823_ = ~new_n13819_ & new_n13822_;
  assign new_n13824_ = new_n13818_ & new_n13823_;
  assign new_n13825_ = new_n13813_ & new_n13824_;
  assign new_n13826_ = new_n7115_ & new_n10107_;
  assign new_n13827_ = new_n7115_ & new_n10109_;
  assign new_n13828_ = new_n7115_ & new_n10111_;
  assign new_n13829_ = ~new_n13827_ & ~new_n13828_;
  assign new_n13830_ = ~new_n13826_ & new_n13829_;
  assign new_n13831_ = new_n7115_ & new_n10116_;
  assign new_n13832_ = new_n7115_ & new_n10118_;
  assign new_n13833_ = new_n7115_ & new_n10120_;
  assign new_n13834_ = ~new_n13832_ & ~new_n13833_;
  assign new_n13835_ = ~new_n13831_ & new_n13834_;
  assign new_n13836_ = new_n13830_ & new_n13835_;
  assign new_n13837_ = new_n7281_ & new_n9924_;
  assign new_n13838_ = new_n7281_ & new_n9926_;
  assign new_n13839_ = new_n7281_ & new_n9928_;
  assign new_n13840_ = ~new_n13838_ & ~new_n13839_;
  assign new_n13841_ = ~new_n13837_ & new_n13840_;
  assign new_n13842_ = new_n7281_ & new_n9936_;
  assign new_n13843_ = new_n7281_ & new_n9938_;
  assign new_n13844_ = ~new_n13842_ & ~new_n13843_;
  assign new_n13845_ = new_n13841_ & new_n13844_;
  assign new_n13846_ = new_n13836_ & new_n13845_;
  assign new_n13847_ = new_n13825_ & new_n13846_;
  assign new_n13848_ = new_n7281_ & new_n9946_;
  assign new_n13849_ = new_n7281_ & new_n9934_;
  assign new_n13850_ = new_n7281_ & new_n9944_;
  assign new_n13851_ = ~new_n13849_ & ~new_n13850_;
  assign new_n13852_ = ~new_n13848_ & new_n13851_;
  assign new_n13853_ = new_n7281_ & new_n9956_;
  assign new_n13854_ = new_n7281_ & new_n9942_;
  assign new_n13855_ = new_n7281_ & new_n9954_;
  assign new_n13856_ = ~new_n13854_ & ~new_n13855_;
  assign new_n13857_ = ~new_n13853_ & new_n13856_;
  assign new_n13858_ = new_n13852_ & new_n13857_;
  assign new_n13859_ = new_n7281_ & new_n9965_;
  assign new_n13860_ = new_n7281_ & new_n9952_;
  assign new_n13861_ = new_n7281_ & new_n9963_;
  assign new_n13862_ = ~new_n13860_ & ~new_n13861_;
  assign new_n13863_ = ~new_n13859_ & new_n13862_;
  assign new_n13864_ = new_n7281_ & new_n9974_;
  assign new_n13865_ = new_n7281_ & new_n9961_;
  assign new_n13866_ = new_n7281_ & new_n9972_;
  assign new_n13867_ = ~new_n13865_ & ~new_n13866_;
  assign new_n13868_ = ~new_n13864_ & new_n13867_;
  assign new_n13869_ = new_n13863_ & new_n13868_;
  assign new_n13870_ = new_n13858_ & new_n13869_;
  assign new_n13871_ = new_n7281_ & new_n9980_;
  assign new_n13872_ = new_n7281_ & new_n9970_;
  assign new_n13873_ = new_n7281_ & new_n9978_;
  assign new_n13874_ = ~new_n13872_ & ~new_n13873_;
  assign new_n13875_ = ~new_n13871_ & new_n13874_;
  assign new_n13876_ = new_n7281_ & new_n9988_;
  assign new_n13877_ = new_n7281_ & new_n9990_;
  assign new_n13878_ = new_n7281_ & new_n9992_;
  assign new_n13879_ = ~new_n13877_ & ~new_n13878_;
  assign new_n13880_ = ~new_n13876_ & new_n13879_;
  assign new_n13881_ = new_n13875_ & new_n13880_;
  assign new_n13882_ = new_n7281_ & new_n9997_;
  assign new_n13883_ = new_n7281_ & new_n9999_;
  assign new_n13884_ = new_n7281_ & new_n10001_;
  assign new_n13885_ = ~new_n13883_ & ~new_n13884_;
  assign new_n13886_ = ~new_n13882_ & new_n13885_;
  assign new_n13887_ = new_n7281_ & new_n10009_;
  assign new_n13888_ = new_n7281_ & new_n10011_;
  assign new_n13889_ = ~new_n13887_ & ~new_n13888_;
  assign new_n13890_ = new_n13886_ & new_n13889_;
  assign new_n13891_ = new_n13881_ & new_n13890_;
  assign new_n13892_ = new_n13870_ & new_n13891_;
  assign new_n13893_ = new_n13847_ & new_n13892_;
  assign new_n13894_ = new_n13802_ & new_n13893_;
  assign new_n13895_ = new_n13711_ & new_n13894_;
  assign new_n13896_ = new_n13526_ & new_n13895_;
  assign new_n13897_ = new_n7281_ & new_n10019_;
  assign new_n13898_ = new_n7281_ & new_n10007_;
  assign new_n13899_ = new_n7281_ & new_n10017_;
  assign new_n13900_ = ~new_n13898_ & ~new_n13899_;
  assign new_n13901_ = ~new_n13897_ & new_n13900_;
  assign new_n13902_ = new_n7281_ & new_n10030_;
  assign new_n13903_ = new_n7281_ & new_n10015_;
  assign new_n13904_ = new_n7281_ & new_n10028_;
  assign new_n13905_ = ~new_n13903_ & ~new_n13904_;
  assign new_n13906_ = ~new_n13902_ & new_n13905_;
  assign new_n13907_ = new_n13901_ & new_n13906_;
  assign new_n13908_ = new_n7281_ & new_n10039_;
  assign new_n13909_ = new_n7281_ & new_n10026_;
  assign new_n13910_ = new_n7281_ & new_n10037_;
  assign new_n13911_ = ~new_n13909_ & ~new_n13910_;
  assign new_n13912_ = ~new_n13908_ & new_n13911_;
  assign new_n13913_ = new_n7281_ & new_n10048_;
  assign new_n13914_ = new_n7281_ & new_n10035_;
  assign new_n13915_ = new_n7281_ & new_n10046_;
  assign new_n13916_ = ~new_n13914_ & ~new_n13915_;
  assign new_n13917_ = ~new_n13913_ & new_n13916_;
  assign new_n13918_ = new_n13912_ & new_n13917_;
  assign new_n13919_ = new_n13907_ & new_n13918_;
  assign new_n13920_ = new_n7281_ & new_n10054_;
  assign new_n13921_ = new_n7281_ & new_n10044_;
  assign new_n13922_ = new_n7281_ & new_n10052_;
  assign new_n13923_ = ~new_n13921_ & ~new_n13922_;
  assign new_n13924_ = ~new_n13920_ & new_n13923_;
  assign new_n13925_ = new_n7281_ & new_n10061_;
  assign new_n13926_ = new_n7281_ & new_n10063_;
  assign new_n13927_ = new_n7281_ & new_n10065_;
  assign new_n13928_ = ~new_n13926_ & ~new_n13927_;
  assign new_n13929_ = ~new_n13925_ & new_n13928_;
  assign new_n13930_ = new_n13924_ & new_n13929_;
  assign new_n13931_ = new_n7281_ & new_n10069_;
  assign new_n13932_ = new_n7281_ & new_n10071_;
  assign new_n13933_ = new_n7281_ & new_n10073_;
  assign new_n13934_ = ~new_n13932_ & ~new_n13933_;
  assign new_n13935_ = ~new_n13931_ & new_n13934_;
  assign new_n13936_ = new_n7281_ & new_n10078_;
  assign new_n13937_ = new_n7281_ & new_n10080_;
  assign new_n13938_ = new_n7281_ & new_n10082_;
  assign new_n13939_ = ~new_n13937_ & ~new_n13938_;
  assign new_n13940_ = ~new_n13936_ & new_n13939_;
  assign new_n13941_ = new_n13935_ & new_n13940_;
  assign new_n13942_ = new_n13930_ & new_n13941_;
  assign new_n13943_ = new_n13919_ & new_n13942_;
  assign new_n13944_ = new_n7281_ & new_n10087_;
  assign new_n13945_ = new_n7281_ & new_n10089_;
  assign new_n13946_ = new_n7281_ & new_n10091_;
  assign new_n13947_ = ~new_n13945_ & ~new_n13946_;
  assign new_n13948_ = ~new_n13944_ & new_n13947_;
  assign new_n13949_ = new_n7281_ & new_n10098_;
  assign new_n13950_ = new_n7281_ & new_n10100_;
  assign new_n13951_ = new_n7281_ & new_n10102_;
  assign new_n13952_ = ~new_n13950_ & ~new_n13951_;
  assign new_n13953_ = ~new_n13949_ & new_n13952_;
  assign new_n13954_ = new_n13948_ & new_n13953_;
  assign new_n13955_ = new_n7281_ & new_n10107_;
  assign new_n13956_ = new_n7281_ & new_n10109_;
  assign new_n13957_ = new_n7281_ & new_n10111_;
  assign new_n13958_ = ~new_n13956_ & ~new_n13957_;
  assign new_n13959_ = ~new_n13955_ & new_n13958_;
  assign new_n13960_ = new_n7281_ & new_n10116_;
  assign new_n13961_ = new_n7281_ & new_n10118_;
  assign new_n13962_ = new_n7281_ & new_n10120_;
  assign new_n13963_ = ~new_n13961_ & ~new_n13962_;
  assign new_n13964_ = ~new_n13960_ & new_n13963_;
  assign new_n13965_ = new_n13959_ & new_n13964_;
  assign new_n13966_ = new_n13954_ & new_n13965_;
  assign new_n13967_ = new_n7446_ & new_n9924_;
  assign new_n13968_ = new_n7446_ & new_n9926_;
  assign new_n13969_ = new_n7446_ & new_n9928_;
  assign new_n13970_ = ~new_n13968_ & ~new_n13969_;
  assign new_n13971_ = ~new_n13967_ & new_n13970_;
  assign new_n13972_ = new_n7446_ & new_n9934_;
  assign new_n13973_ = new_n7446_ & new_n9936_;
  assign new_n13974_ = new_n7446_ & new_n9938_;
  assign new_n13975_ = ~new_n13973_ & ~new_n13974_;
  assign new_n13976_ = ~new_n13972_ & new_n13975_;
  assign new_n13977_ = new_n13971_ & new_n13976_;
  assign new_n13978_ = new_n7446_ & new_n9942_;
  assign new_n13979_ = new_n7446_ & new_n9944_;
  assign new_n13980_ = new_n7446_ & new_n9946_;
  assign new_n13981_ = ~new_n13979_ & ~new_n13980_;
  assign new_n13982_ = ~new_n13978_ & new_n13981_;
  assign new_n13983_ = new_n7446_ & new_n9954_;
  assign new_n13984_ = new_n7446_ & new_n9956_;
  assign new_n13985_ = ~new_n13983_ & ~new_n13984_;
  assign new_n13986_ = new_n13982_ & new_n13985_;
  assign new_n13987_ = new_n13977_ & new_n13986_;
  assign new_n13988_ = new_n13966_ & new_n13987_;
  assign new_n13989_ = new_n13943_ & new_n13988_;
  assign new_n13990_ = new_n7446_ & new_n9965_;
  assign new_n13991_ = new_n7446_ & new_n9952_;
  assign new_n13992_ = new_n7446_ & new_n9963_;
  assign new_n13993_ = ~new_n13991_ & ~new_n13992_;
  assign new_n13994_ = ~new_n13990_ & new_n13993_;
  assign new_n13995_ = new_n7446_ & new_n9974_;
  assign new_n13996_ = new_n7446_ & new_n9961_;
  assign new_n13997_ = new_n7446_ & new_n9972_;
  assign new_n13998_ = ~new_n13996_ & ~new_n13997_;
  assign new_n13999_ = ~new_n13995_ & new_n13998_;
  assign new_n14000_ = new_n13994_ & new_n13999_;
  assign new_n14001_ = new_n7446_ & new_n9980_;
  assign new_n14002_ = new_n7446_ & new_n9970_;
  assign new_n14003_ = new_n7446_ & new_n9978_;
  assign new_n14004_ = ~new_n14002_ & ~new_n14003_;
  assign new_n14005_ = ~new_n14001_ & new_n14004_;
  assign new_n14006_ = new_n7446_ & new_n9988_;
  assign new_n14007_ = new_n7446_ & new_n9990_;
  assign new_n14008_ = new_n7446_ & new_n9992_;
  assign new_n14009_ = ~new_n14007_ & ~new_n14008_;
  assign new_n14010_ = ~new_n14006_ & new_n14009_;
  assign new_n14011_ = new_n14005_ & new_n14010_;
  assign new_n14012_ = new_n14000_ & new_n14011_;
  assign new_n14013_ = new_n7446_ & new_n9997_;
  assign new_n14014_ = new_n7446_ & new_n9999_;
  assign new_n14015_ = new_n7446_ & new_n10001_;
  assign new_n14016_ = ~new_n14014_ & ~new_n14015_;
  assign new_n14017_ = ~new_n14013_ & new_n14016_;
  assign new_n14018_ = new_n7446_ & new_n10007_;
  assign new_n14019_ = new_n7446_ & new_n10009_;
  assign new_n14020_ = new_n7446_ & new_n10011_;
  assign new_n14021_ = ~new_n14019_ & ~new_n14020_;
  assign new_n14022_ = ~new_n14018_ & new_n14021_;
  assign new_n14023_ = new_n14017_ & new_n14022_;
  assign new_n14024_ = new_n7446_ & new_n10015_;
  assign new_n14025_ = new_n7446_ & new_n10017_;
  assign new_n14026_ = new_n7446_ & new_n10019_;
  assign new_n14027_ = ~new_n14025_ & ~new_n14026_;
  assign new_n14028_ = ~new_n14024_ & new_n14027_;
  assign new_n14029_ = new_n7446_ & new_n10028_;
  assign new_n14030_ = new_n7446_ & new_n10030_;
  assign new_n14031_ = ~new_n14029_ & ~new_n14030_;
  assign new_n14032_ = new_n14028_ & new_n14031_;
  assign new_n14033_ = new_n14023_ & new_n14032_;
  assign new_n14034_ = new_n14012_ & new_n14033_;
  assign new_n14035_ = new_n7446_ & new_n10039_;
  assign new_n14036_ = new_n7446_ & new_n10026_;
  assign new_n14037_ = new_n7446_ & new_n10037_;
  assign new_n14038_ = ~new_n14036_ & ~new_n14037_;
  assign new_n14039_ = ~new_n14035_ & new_n14038_;
  assign new_n14040_ = new_n7446_ & new_n10048_;
  assign new_n14041_ = new_n7446_ & new_n10035_;
  assign new_n14042_ = new_n7446_ & new_n10046_;
  assign new_n14043_ = ~new_n14041_ & ~new_n14042_;
  assign new_n14044_ = ~new_n14040_ & new_n14043_;
  assign new_n14045_ = new_n14039_ & new_n14044_;
  assign new_n14046_ = new_n7446_ & new_n10054_;
  assign new_n14047_ = new_n7446_ & new_n10044_;
  assign new_n14048_ = new_n7446_ & new_n10052_;
  assign new_n14049_ = ~new_n14047_ & ~new_n14048_;
  assign new_n14050_ = ~new_n14046_ & new_n14049_;
  assign new_n14051_ = new_n7446_ & new_n10061_;
  assign new_n14052_ = new_n7446_ & new_n10063_;
  assign new_n14053_ = new_n7446_ & new_n10065_;
  assign new_n14054_ = ~new_n14052_ & ~new_n14053_;
  assign new_n14055_ = ~new_n14051_ & new_n14054_;
  assign new_n14056_ = new_n14050_ & new_n14055_;
  assign new_n14057_ = new_n14045_ & new_n14056_;
  assign new_n14058_ = new_n7446_ & new_n10069_;
  assign new_n14059_ = new_n7446_ & new_n10071_;
  assign new_n14060_ = new_n7446_ & new_n10073_;
  assign new_n14061_ = ~new_n14059_ & ~new_n14060_;
  assign new_n14062_ = ~new_n14058_ & new_n14061_;
  assign new_n14063_ = new_n7446_ & new_n10078_;
  assign new_n14064_ = new_n7446_ & new_n10080_;
  assign new_n14065_ = new_n7446_ & new_n10082_;
  assign new_n14066_ = ~new_n14064_ & ~new_n14065_;
  assign new_n14067_ = ~new_n14063_ & new_n14066_;
  assign new_n14068_ = new_n14062_ & new_n14067_;
  assign new_n14069_ = new_n7446_ & new_n10087_;
  assign new_n14070_ = new_n7446_ & new_n10089_;
  assign new_n14071_ = new_n7446_ & new_n10091_;
  assign new_n14072_ = ~new_n14070_ & ~new_n14071_;
  assign new_n14073_ = ~new_n14069_ & new_n14072_;
  assign new_n14074_ = new_n7446_ & new_n10100_;
  assign new_n14075_ = new_n7446_ & new_n10102_;
  assign new_n14076_ = ~new_n14074_ & ~new_n14075_;
  assign new_n14077_ = new_n14073_ & new_n14076_;
  assign new_n14078_ = new_n14068_ & new_n14077_;
  assign new_n14079_ = new_n14057_ & new_n14078_;
  assign new_n14080_ = new_n14034_ & new_n14079_;
  assign new_n14081_ = new_n13989_ & new_n14080_;
  assign new_n14082_ = new_n7446_ & new_n10111_;
  assign new_n14083_ = new_n7446_ & new_n10098_;
  assign new_n14084_ = new_n7446_ & new_n10109_;
  assign new_n14085_ = ~new_n14083_ & ~new_n14084_;
  assign new_n14086_ = ~new_n14082_ & new_n14085_;
  assign new_n14087_ = new_n7446_ & new_n10120_;
  assign new_n14088_ = new_n7446_ & new_n10107_;
  assign new_n14089_ = new_n7446_ & new_n10118_;
  assign new_n14090_ = ~new_n14088_ & ~new_n14089_;
  assign new_n14091_ = ~new_n14087_ & new_n14090_;
  assign new_n14092_ = new_n14086_ & new_n14091_;
  assign new_n14093_ = new_n7610_ & new_n9928_;
  assign new_n14094_ = new_n7446_ & new_n10116_;
  assign new_n14095_ = new_n7610_ & new_n9926_;
  assign new_n14096_ = ~new_n14094_ & ~new_n14095_;
  assign new_n14097_ = ~new_n14093_ & new_n14096_;
  assign new_n14098_ = new_n7610_ & new_n9938_;
  assign new_n14099_ = new_n7610_ & new_n9924_;
  assign new_n14100_ = new_n7610_ & new_n9936_;
  assign new_n14101_ = ~new_n14099_ & ~new_n14100_;
  assign new_n14102_ = ~new_n14098_ & new_n14101_;
  assign new_n14103_ = new_n14097_ & new_n14102_;
  assign new_n14104_ = new_n14092_ & new_n14103_;
  assign new_n14105_ = new_n7610_ & new_n9946_;
  assign new_n14106_ = new_n7610_ & new_n9934_;
  assign new_n14107_ = new_n7610_ & new_n9944_;
  assign new_n14108_ = ~new_n14106_ & ~new_n14107_;
  assign new_n14109_ = ~new_n14105_ & new_n14108_;
  assign new_n14110_ = new_n7610_ & new_n9956_;
  assign new_n14111_ = new_n7610_ & new_n9942_;
  assign new_n14112_ = new_n7610_ & new_n9954_;
  assign new_n14113_ = ~new_n14111_ & ~new_n14112_;
  assign new_n14114_ = ~new_n14110_ & new_n14113_;
  assign new_n14115_ = new_n14109_ & new_n14114_;
  assign new_n14116_ = new_n7610_ & new_n9965_;
  assign new_n14117_ = new_n7610_ & new_n9952_;
  assign new_n14118_ = new_n7610_ & new_n9963_;
  assign new_n14119_ = ~new_n14117_ & ~new_n14118_;
  assign new_n14120_ = ~new_n14116_ & new_n14119_;
  assign new_n14121_ = new_n7610_ & new_n9961_;
  assign new_n14122_ = new_n7610_ & new_n9972_;
  assign new_n14123_ = ~new_n14121_ & ~new_n14122_;
  assign new_n14124_ = new_n14120_ & new_n14123_;
  assign new_n14125_ = new_n14115_ & new_n14124_;
  assign new_n14126_ = new_n14104_ & new_n14125_;
  assign new_n14127_ = new_n7610_ & new_n9978_;
  assign new_n14128_ = new_n7610_ & new_n9974_;
  assign new_n14129_ = new_n7610_ & new_n9970_;
  assign new_n14130_ = ~new_n14128_ & ~new_n14129_;
  assign new_n14131_ = ~new_n14127_ & new_n14130_;
  assign new_n14132_ = new_n7610_ & new_n9992_;
  assign new_n14133_ = new_n7610_ & new_n9980_;
  assign new_n14134_ = new_n7610_ & new_n9990_;
  assign new_n14135_ = ~new_n14133_ & ~new_n14134_;
  assign new_n14136_ = ~new_n14132_ & new_n14135_;
  assign new_n14137_ = new_n14131_ & new_n14136_;
  assign new_n14138_ = new_n7610_ & new_n10001_;
  assign new_n14139_ = new_n7610_ & new_n9988_;
  assign new_n14140_ = new_n7610_ & new_n9999_;
  assign new_n14141_ = ~new_n14139_ & ~new_n14140_;
  assign new_n14142_ = ~new_n14138_ & new_n14141_;
  assign new_n14143_ = new_n7610_ & new_n10011_;
  assign new_n14144_ = new_n7610_ & new_n9997_;
  assign new_n14145_ = new_n7610_ & new_n10009_;
  assign new_n14146_ = ~new_n14144_ & ~new_n14145_;
  assign new_n14147_ = ~new_n14143_ & new_n14146_;
  assign new_n14148_ = new_n14142_ & new_n14147_;
  assign new_n14149_ = new_n14137_ & new_n14148_;
  assign new_n14150_ = new_n7610_ & new_n10019_;
  assign new_n14151_ = new_n7610_ & new_n10007_;
  assign new_n14152_ = new_n7610_ & new_n10017_;
  assign new_n14153_ = ~new_n14151_ & ~new_n14152_;
  assign new_n14154_ = ~new_n14150_ & new_n14153_;
  assign new_n14155_ = new_n7610_ & new_n10030_;
  assign new_n14156_ = new_n7610_ & new_n10015_;
  assign new_n14157_ = new_n7610_ & new_n10028_;
  assign new_n14158_ = ~new_n14156_ & ~new_n14157_;
  assign new_n14159_ = ~new_n14155_ & new_n14158_;
  assign new_n14160_ = new_n14154_ & new_n14159_;
  assign new_n14161_ = new_n7610_ & new_n10039_;
  assign new_n14162_ = new_n7610_ & new_n10026_;
  assign new_n14163_ = new_n7610_ & new_n10037_;
  assign new_n14164_ = ~new_n14162_ & ~new_n14163_;
  assign new_n14165_ = ~new_n14161_ & new_n14164_;
  assign new_n14166_ = new_n7610_ & new_n10035_;
  assign new_n14167_ = new_n7610_ & new_n10046_;
  assign new_n14168_ = ~new_n14166_ & ~new_n14167_;
  assign new_n14169_ = new_n14165_ & new_n14168_;
  assign new_n14170_ = new_n14160_ & new_n14169_;
  assign new_n14171_ = new_n14149_ & new_n14170_;
  assign new_n14172_ = new_n14126_ & new_n14171_;
  assign new_n14173_ = new_n7610_ & new_n10052_;
  assign new_n14174_ = new_n7610_ & new_n10048_;
  assign new_n14175_ = new_n7610_ & new_n10044_;
  assign new_n14176_ = ~new_n14174_ & ~new_n14175_;
  assign new_n14177_ = ~new_n14173_ & new_n14176_;
  assign new_n14178_ = new_n7610_ & new_n10065_;
  assign new_n14179_ = new_n7610_ & new_n10054_;
  assign new_n14180_ = new_n7610_ & new_n10063_;
  assign new_n14181_ = ~new_n14179_ & ~new_n14180_;
  assign new_n14182_ = ~new_n14178_ & new_n14181_;
  assign new_n14183_ = new_n14177_ & new_n14182_;
  assign new_n14184_ = new_n7610_ & new_n10073_;
  assign new_n14185_ = new_n7610_ & new_n10061_;
  assign new_n14186_ = new_n7610_ & new_n10071_;
  assign new_n14187_ = ~new_n14185_ & ~new_n14186_;
  assign new_n14188_ = ~new_n14184_ & new_n14187_;
  assign new_n14189_ = new_n7610_ & new_n10082_;
  assign new_n14190_ = new_n7610_ & new_n10069_;
  assign new_n14191_ = new_n7610_ & new_n10080_;
  assign new_n14192_ = ~new_n14190_ & ~new_n14191_;
  assign new_n14193_ = ~new_n14189_ & new_n14192_;
  assign new_n14194_ = new_n14188_ & new_n14193_;
  assign new_n14195_ = new_n14183_ & new_n14194_;
  assign new_n14196_ = new_n7610_ & new_n10091_;
  assign new_n14197_ = new_n7610_ & new_n10078_;
  assign new_n14198_ = new_n7610_ & new_n10089_;
  assign new_n14199_ = ~new_n14197_ & ~new_n14198_;
  assign new_n14200_ = ~new_n14196_ & new_n14199_;
  assign new_n14201_ = new_n7610_ & new_n10102_;
  assign new_n14202_ = new_n7610_ & new_n10087_;
  assign new_n14203_ = new_n7610_ & new_n10100_;
  assign new_n14204_ = ~new_n14202_ & ~new_n14203_;
  assign new_n14205_ = ~new_n14201_ & new_n14204_;
  assign new_n14206_ = new_n14200_ & new_n14205_;
  assign new_n14207_ = new_n7610_ & new_n10111_;
  assign new_n14208_ = new_n7610_ & new_n10098_;
  assign new_n14209_ = new_n7610_ & new_n10109_;
  assign new_n14210_ = ~new_n14208_ & ~new_n14209_;
  assign new_n14211_ = ~new_n14207_ & new_n14210_;
  assign new_n14212_ = new_n7610_ & new_n10107_;
  assign new_n14213_ = new_n7610_ & new_n10118_;
  assign new_n14214_ = ~new_n14212_ & ~new_n14213_;
  assign new_n14215_ = new_n14211_ & new_n14214_;
  assign new_n14216_ = new_n14206_ & new_n14215_;
  assign new_n14217_ = new_n14195_ & new_n14216_;
  assign new_n14218_ = new_n8030_ & new_n9926_;
  assign new_n14219_ = new_n7610_ & new_n10120_;
  assign new_n14220_ = new_n7610_ & new_n10116_;
  assign new_n14221_ = ~new_n14219_ & ~new_n14220_;
  assign new_n14222_ = ~new_n14218_ & new_n14221_;
  assign new_n14223_ = new_n8030_ & new_n9936_;
  assign new_n14224_ = new_n8030_ & new_n9928_;
  assign new_n14225_ = new_n8030_ & new_n9924_;
  assign new_n14226_ = ~new_n14224_ & ~new_n14225_;
  assign new_n14227_ = ~new_n14223_ & new_n14226_;
  assign new_n14228_ = new_n14222_ & new_n14227_;
  assign new_n14229_ = new_n8030_ & new_n9944_;
  assign new_n14230_ = new_n8030_ & new_n9938_;
  assign new_n14231_ = new_n8030_ & new_n9934_;
  assign new_n14232_ = ~new_n14230_ & ~new_n14231_;
  assign new_n14233_ = ~new_n14229_ & new_n14232_;
  assign new_n14234_ = new_n8030_ & new_n9954_;
  assign new_n14235_ = new_n8030_ & new_n9946_;
  assign new_n14236_ = new_n8030_ & new_n9942_;
  assign new_n14237_ = ~new_n14235_ & ~new_n14236_;
  assign new_n14238_ = ~new_n14234_ & new_n14237_;
  assign new_n14239_ = new_n14233_ & new_n14238_;
  assign new_n14240_ = new_n14228_ & new_n14239_;
  assign new_n14241_ = new_n8030_ & new_n9963_;
  assign new_n14242_ = new_n8030_ & new_n9956_;
  assign new_n14243_ = new_n8030_ & new_n9952_;
  assign new_n14244_ = ~new_n14242_ & ~new_n14243_;
  assign new_n14245_ = ~new_n14241_ & new_n14244_;
  assign new_n14246_ = new_n8030_ & new_n9972_;
  assign new_n14247_ = new_n8030_ & new_n9965_;
  assign new_n14248_ = new_n8030_ & new_n9961_;
  assign new_n14249_ = ~new_n14247_ & ~new_n14248_;
  assign new_n14250_ = ~new_n14246_ & new_n14249_;
  assign new_n14251_ = new_n14245_ & new_n14250_;
  assign new_n14252_ = new_n8030_ & new_n9978_;
  assign new_n14253_ = new_n8030_ & new_n9974_;
  assign new_n14254_ = new_n8030_ & new_n9970_;
  assign new_n14255_ = ~new_n14253_ & ~new_n14254_;
  assign new_n14256_ = ~new_n14252_ & new_n14255_;
  assign new_n14257_ = new_n8030_ & new_n9980_;
  assign new_n14258_ = new_n8030_ & new_n9990_;
  assign new_n14259_ = ~new_n14257_ & ~new_n14258_;
  assign new_n14260_ = new_n14256_ & new_n14259_;
  assign new_n14261_ = new_n14251_ & new_n14260_;
  assign new_n14262_ = new_n14240_ & new_n14261_;
  assign new_n14263_ = new_n14217_ & new_n14262_;
  assign new_n14264_ = new_n14172_ & new_n14263_;
  assign new_n14265_ = new_n14081_ & new_n14264_;
  assign new_n14266_ = new_n8030_ & new_n9999_;
  assign new_n14267_ = new_n8030_ & new_n9992_;
  assign new_n14268_ = new_n8030_ & new_n9988_;
  assign new_n14269_ = ~new_n14267_ & ~new_n14268_;
  assign new_n14270_ = ~new_n14266_ & new_n14269_;
  assign new_n14271_ = new_n8030_ & new_n10009_;
  assign new_n14272_ = new_n8030_ & new_n10001_;
  assign new_n14273_ = new_n8030_ & new_n9997_;
  assign new_n14274_ = ~new_n14272_ & ~new_n14273_;
  assign new_n14275_ = ~new_n14271_ & new_n14274_;
  assign new_n14276_ = new_n14270_ & new_n14275_;
  assign new_n14277_ = new_n8030_ & new_n10017_;
  assign new_n14278_ = new_n8030_ & new_n10011_;
  assign new_n14279_ = new_n8030_ & new_n10007_;
  assign new_n14280_ = ~new_n14278_ & ~new_n14279_;
  assign new_n14281_ = ~new_n14277_ & new_n14280_;
  assign new_n14282_ = new_n8030_ & new_n10028_;
  assign new_n14283_ = new_n8030_ & new_n10019_;
  assign new_n14284_ = new_n8030_ & new_n10015_;
  assign new_n14285_ = ~new_n14283_ & ~new_n14284_;
  assign new_n14286_ = ~new_n14282_ & new_n14285_;
  assign new_n14287_ = new_n14281_ & new_n14286_;
  assign new_n14288_ = new_n14276_ & new_n14287_;
  assign new_n14289_ = new_n8030_ & new_n10037_;
  assign new_n14290_ = new_n8030_ & new_n10030_;
  assign new_n14291_ = new_n8030_ & new_n10026_;
  assign new_n14292_ = ~new_n14290_ & ~new_n14291_;
  assign new_n14293_ = ~new_n14289_ & new_n14292_;
  assign new_n14294_ = new_n8030_ & new_n10046_;
  assign new_n14295_ = new_n8030_ & new_n10039_;
  assign new_n14296_ = new_n8030_ & new_n10035_;
  assign new_n14297_ = ~new_n14295_ & ~new_n14296_;
  assign new_n14298_ = ~new_n14294_ & new_n14297_;
  assign new_n14299_ = new_n14293_ & new_n14298_;
  assign new_n14300_ = new_n8030_ & new_n10052_;
  assign new_n14301_ = new_n8030_ & new_n10048_;
  assign new_n14302_ = new_n8030_ & new_n10044_;
  assign new_n14303_ = ~new_n14301_ & ~new_n14302_;
  assign new_n14304_ = ~new_n14300_ & new_n14303_;
  assign new_n14305_ = new_n8030_ & new_n10054_;
  assign new_n14306_ = new_n8030_ & new_n10063_;
  assign new_n14307_ = ~new_n14305_ & ~new_n14306_;
  assign new_n14308_ = new_n14304_ & new_n14307_;
  assign new_n14309_ = new_n14299_ & new_n14308_;
  assign new_n14310_ = new_n14288_ & new_n14309_;
  assign new_n14311_ = new_n8030_ & new_n10071_;
  assign new_n14312_ = new_n8030_ & new_n10065_;
  assign new_n14313_ = new_n8030_ & new_n10061_;
  assign new_n14314_ = ~new_n14312_ & ~new_n14313_;
  assign new_n14315_ = ~new_n14311_ & new_n14314_;
  assign new_n14316_ = new_n8030_ & new_n10080_;
  assign new_n14317_ = new_n8030_ & new_n10073_;
  assign new_n14318_ = new_n8030_ & new_n10069_;
  assign new_n14319_ = ~new_n14317_ & ~new_n14318_;
  assign new_n14320_ = ~new_n14316_ & new_n14319_;
  assign new_n14321_ = new_n14315_ & new_n14320_;
  assign new_n14322_ = new_n8030_ & new_n10089_;
  assign new_n14323_ = new_n8030_ & new_n10082_;
  assign new_n14324_ = new_n8030_ & new_n10078_;
  assign new_n14325_ = ~new_n14323_ & ~new_n14324_;
  assign new_n14326_ = ~new_n14322_ & new_n14325_;
  assign new_n14327_ = new_n8030_ & new_n10100_;
  assign new_n14328_ = new_n8030_ & new_n10091_;
  assign new_n14329_ = new_n8030_ & new_n10087_;
  assign new_n14330_ = ~new_n14328_ & ~new_n14329_;
  assign new_n14331_ = ~new_n14327_ & new_n14330_;
  assign new_n14332_ = new_n14326_ & new_n14331_;
  assign new_n14333_ = new_n14321_ & new_n14332_;
  assign new_n14334_ = new_n8030_ & new_n10109_;
  assign new_n14335_ = new_n8030_ & new_n10102_;
  assign new_n14336_ = new_n8030_ & new_n10098_;
  assign new_n14337_ = ~new_n14335_ & ~new_n14336_;
  assign new_n14338_ = ~new_n14334_ & new_n14337_;
  assign new_n14339_ = new_n8030_ & new_n10118_;
  assign new_n14340_ = new_n8030_ & new_n10111_;
  assign new_n14341_ = new_n8030_ & new_n10107_;
  assign new_n14342_ = ~new_n14340_ & ~new_n14341_;
  assign new_n14343_ = ~new_n14339_ & new_n14342_;
  assign new_n14344_ = new_n14338_ & new_n14343_;
  assign new_n14345_ = new_n8192_ & new_n9926_;
  assign new_n14346_ = new_n8030_ & new_n10120_;
  assign new_n14347_ = new_n8030_ & new_n10116_;
  assign new_n14348_ = ~new_n14346_ & ~new_n14347_;
  assign new_n14349_ = ~new_n14345_ & new_n14348_;
  assign new_n14350_ = new_n8192_ & new_n9928_;
  assign new_n14351_ = new_n8192_ & new_n9924_;
  assign new_n14352_ = ~new_n14350_ & ~new_n14351_;
  assign new_n14353_ = new_n14349_ & new_n14352_;
  assign new_n14354_ = new_n14344_ & new_n14353_;
  assign new_n14355_ = new_n14333_ & new_n14354_;
  assign new_n14356_ = new_n14310_ & new_n14355_;
  assign new_n14357_ = new_n8192_ & new_n9934_;
  assign new_n14358_ = new_n8192_ & new_n9936_;
  assign new_n14359_ = new_n8192_ & new_n9938_;
  assign new_n14360_ = ~new_n14358_ & ~new_n14359_;
  assign new_n14361_ = ~new_n14357_ & new_n14360_;
  assign new_n14362_ = new_n8192_ & new_n9942_;
  assign new_n14363_ = new_n8192_ & new_n9944_;
  assign new_n14364_ = new_n8192_ & new_n9946_;
  assign new_n14365_ = ~new_n14363_ & ~new_n14364_;
  assign new_n14366_ = ~new_n14362_ & new_n14365_;
  assign new_n14367_ = new_n14361_ & new_n14366_;
  assign new_n14368_ = new_n8192_ & new_n9952_;
  assign new_n14369_ = new_n8192_ & new_n9954_;
  assign new_n14370_ = new_n8192_ & new_n9956_;
  assign new_n14371_ = ~new_n14369_ & ~new_n14370_;
  assign new_n14372_ = ~new_n14368_ & new_n14371_;
  assign new_n14373_ = new_n8192_ & new_n9961_;
  assign new_n14374_ = new_n8192_ & new_n9963_;
  assign new_n14375_ = new_n8192_ & new_n9965_;
  assign new_n14376_ = ~new_n14374_ & ~new_n14375_;
  assign new_n14377_ = ~new_n14373_ & new_n14376_;
  assign new_n14378_ = new_n14372_ & new_n14377_;
  assign new_n14379_ = new_n14367_ & new_n14378_;
  assign new_n14380_ = new_n8192_ & new_n9970_;
  assign new_n14381_ = new_n8192_ & new_n9972_;
  assign new_n14382_ = new_n8192_ & new_n9974_;
  assign new_n14383_ = ~new_n14381_ & ~new_n14382_;
  assign new_n14384_ = ~new_n14380_ & new_n14383_;
  assign new_n14385_ = new_n8192_ & new_n9990_;
  assign new_n14386_ = new_n8192_ & new_n9978_;
  assign new_n14387_ = new_n8192_ & new_n9980_;
  assign new_n14388_ = ~new_n14386_ & ~new_n14387_;
  assign new_n14389_ = ~new_n14385_ & new_n14388_;
  assign new_n14390_ = new_n14384_ & new_n14389_;
  assign new_n14391_ = new_n8192_ & new_n9999_;
  assign new_n14392_ = new_n8192_ & new_n9992_;
  assign new_n14393_ = new_n8192_ & new_n9988_;
  assign new_n14394_ = ~new_n14392_ & ~new_n14393_;
  assign new_n14395_ = ~new_n14391_ & new_n14394_;
  assign new_n14396_ = new_n8192_ & new_n10001_;
  assign new_n14397_ = new_n8192_ & new_n9997_;
  assign new_n14398_ = ~new_n14396_ & ~new_n14397_;
  assign new_n14399_ = new_n14395_ & new_n14398_;
  assign new_n14400_ = new_n14390_ & new_n14399_;
  assign new_n14401_ = new_n14379_ & new_n14400_;
  assign new_n14402_ = new_n8192_ & new_n10007_;
  assign new_n14403_ = new_n8192_ & new_n10009_;
  assign new_n14404_ = new_n8192_ & new_n10011_;
  assign new_n14405_ = ~new_n14403_ & ~new_n14404_;
  assign new_n14406_ = ~new_n14402_ & new_n14405_;
  assign new_n14407_ = new_n8192_ & new_n10015_;
  assign new_n14408_ = new_n8192_ & new_n10017_;
  assign new_n14409_ = new_n8192_ & new_n10019_;
  assign new_n14410_ = ~new_n14408_ & ~new_n14409_;
  assign new_n14411_ = ~new_n14407_ & new_n14410_;
  assign new_n14412_ = new_n14406_ & new_n14411_;
  assign new_n14413_ = new_n8192_ & new_n10026_;
  assign new_n14414_ = new_n8192_ & new_n10028_;
  assign new_n14415_ = new_n8192_ & new_n10030_;
  assign new_n14416_ = ~new_n14414_ & ~new_n14415_;
  assign new_n14417_ = ~new_n14413_ & new_n14416_;
  assign new_n14418_ = new_n8192_ & new_n10035_;
  assign new_n14419_ = new_n8192_ & new_n10037_;
  assign new_n14420_ = new_n8192_ & new_n10039_;
  assign new_n14421_ = ~new_n14419_ & ~new_n14420_;
  assign new_n14422_ = ~new_n14418_ & new_n14421_;
  assign new_n14423_ = new_n14417_ & new_n14422_;
  assign new_n14424_ = new_n14412_ & new_n14423_;
  assign new_n14425_ = new_n8192_ & new_n10044_;
  assign new_n14426_ = new_n8192_ & new_n10046_;
  assign new_n14427_ = new_n8192_ & new_n10048_;
  assign new_n14428_ = ~new_n14426_ & ~new_n14427_;
  assign new_n14429_ = ~new_n14425_ & new_n14428_;
  assign new_n14430_ = new_n8192_ & new_n10063_;
  assign new_n14431_ = new_n8192_ & new_n10052_;
  assign new_n14432_ = new_n8192_ & new_n10054_;
  assign new_n14433_ = ~new_n14431_ & ~new_n14432_;
  assign new_n14434_ = ~new_n14430_ & new_n14433_;
  assign new_n14435_ = new_n14429_ & new_n14434_;
  assign new_n14436_ = new_n8192_ & new_n10071_;
  assign new_n14437_ = new_n8192_ & new_n10065_;
  assign new_n14438_ = new_n8192_ & new_n10061_;
  assign new_n14439_ = ~new_n14437_ & ~new_n14438_;
  assign new_n14440_ = ~new_n14436_ & new_n14439_;
  assign new_n14441_ = new_n8192_ & new_n10073_;
  assign new_n14442_ = new_n8192_ & new_n10069_;
  assign new_n14443_ = ~new_n14441_ & ~new_n14442_;
  assign new_n14444_ = new_n14440_ & new_n14443_;
  assign new_n14445_ = new_n14435_ & new_n14444_;
  assign new_n14446_ = new_n14424_ & new_n14445_;
  assign new_n14447_ = new_n14401_ & new_n14446_;
  assign new_n14448_ = new_n14356_ & new_n14447_;
  assign new_n14449_ = new_n8192_ & new_n10078_;
  assign new_n14450_ = new_n8192_ & new_n10080_;
  assign new_n14451_ = new_n8192_ & new_n10082_;
  assign new_n14452_ = ~new_n14450_ & ~new_n14451_;
  assign new_n14453_ = ~new_n14449_ & new_n14452_;
  assign new_n14454_ = new_n8192_ & new_n10087_;
  assign new_n14455_ = new_n8192_ & new_n10089_;
  assign new_n14456_ = new_n8192_ & new_n10091_;
  assign new_n14457_ = ~new_n14455_ & ~new_n14456_;
  assign new_n14458_ = ~new_n14454_ & new_n14457_;
  assign new_n14459_ = new_n14453_ & new_n14458_;
  assign new_n14460_ = new_n8192_ & new_n10098_;
  assign new_n14461_ = new_n8192_ & new_n10100_;
  assign new_n14462_ = new_n8192_ & new_n10102_;
  assign new_n14463_ = ~new_n14461_ & ~new_n14462_;
  assign new_n14464_ = ~new_n14460_ & new_n14463_;
  assign new_n14465_ = new_n8192_ & new_n10107_;
  assign new_n14466_ = new_n8192_ & new_n10109_;
  assign new_n14467_ = new_n8192_ & new_n10111_;
  assign new_n14468_ = ~new_n14466_ & ~new_n14467_;
  assign new_n14469_ = ~new_n14465_ & new_n14468_;
  assign new_n14470_ = new_n14464_ & new_n14469_;
  assign new_n14471_ = new_n14459_ & new_n14470_;
  assign new_n14472_ = new_n8192_ & new_n10116_;
  assign new_n14473_ = new_n8192_ & new_n10118_;
  assign new_n14474_ = new_n8192_ & new_n10120_;
  assign new_n14475_ = ~new_n14473_ & ~new_n14474_;
  assign new_n14476_ = ~new_n14472_ & new_n14475_;
  assign new_n14477_ = new_n8360_ & new_n9924_;
  assign new_n14478_ = new_n8360_ & new_n9926_;
  assign new_n14479_ = new_n8360_ & new_n9928_;
  assign new_n14480_ = ~new_n14478_ & ~new_n14479_;
  assign new_n14481_ = ~new_n14477_ & new_n14480_;
  assign new_n14482_ = new_n14476_ & new_n14481_;
  assign new_n14483_ = new_n8360_ & new_n9934_;
  assign new_n14484_ = new_n8360_ & new_n9936_;
  assign new_n14485_ = new_n8360_ & new_n9938_;
  assign new_n14486_ = ~new_n14484_ & ~new_n14485_;
  assign new_n14487_ = ~new_n14483_ & new_n14486_;
  assign new_n14488_ = new_n8360_ & new_n9944_;
  assign new_n14489_ = new_n8360_ & new_n9946_;
  assign new_n14490_ = ~new_n14488_ & ~new_n14489_;
  assign new_n14491_ = new_n14487_ & new_n14490_;
  assign new_n14492_ = new_n14482_ & new_n14491_;
  assign new_n14493_ = new_n14471_ & new_n14492_;
  assign new_n14494_ = new_n8360_ & new_n9956_;
  assign new_n14495_ = new_n8360_ & new_n9942_;
  assign new_n14496_ = new_n8360_ & new_n9954_;
  assign new_n14497_ = ~new_n14495_ & ~new_n14496_;
  assign new_n14498_ = ~new_n14494_ & new_n14497_;
  assign new_n14499_ = new_n8360_ & new_n9965_;
  assign new_n14500_ = new_n8360_ & new_n9952_;
  assign new_n14501_ = new_n8360_ & new_n9963_;
  assign new_n14502_ = ~new_n14500_ & ~new_n14501_;
  assign new_n14503_ = ~new_n14499_ & new_n14502_;
  assign new_n14504_ = new_n14498_ & new_n14503_;
  assign new_n14505_ = new_n8360_ & new_n9974_;
  assign new_n14506_ = new_n8360_ & new_n9961_;
  assign new_n14507_ = new_n8360_ & new_n9972_;
  assign new_n14508_ = ~new_n14506_ & ~new_n14507_;
  assign new_n14509_ = ~new_n14505_ & new_n14508_;
  assign new_n14510_ = new_n8360_ & new_n9980_;
  assign new_n14511_ = new_n8360_ & new_n9970_;
  assign new_n14512_ = new_n8360_ & new_n9978_;
  assign new_n14513_ = ~new_n14511_ & ~new_n14512_;
  assign new_n14514_ = ~new_n14510_ & new_n14513_;
  assign new_n14515_ = new_n14509_ & new_n14514_;
  assign new_n14516_ = new_n14504_ & new_n14515_;
  assign new_n14517_ = new_n8360_ & new_n9988_;
  assign new_n14518_ = new_n8360_ & new_n9990_;
  assign new_n14519_ = new_n8360_ & new_n9992_;
  assign new_n14520_ = ~new_n14518_ & ~new_n14519_;
  assign new_n14521_ = ~new_n14517_ & new_n14520_;
  assign new_n14522_ = new_n8360_ & new_n9997_;
  assign new_n14523_ = new_n8360_ & new_n9999_;
  assign new_n14524_ = new_n8360_ & new_n10001_;
  assign new_n14525_ = ~new_n14523_ & ~new_n14524_;
  assign new_n14526_ = ~new_n14522_ & new_n14525_;
  assign new_n14527_ = new_n14521_ & new_n14526_;
  assign new_n14528_ = new_n8360_ & new_n10007_;
  assign new_n14529_ = new_n8360_ & new_n10009_;
  assign new_n14530_ = new_n8360_ & new_n10011_;
  assign new_n14531_ = ~new_n14529_ & ~new_n14530_;
  assign new_n14532_ = ~new_n14528_ & new_n14531_;
  assign new_n14533_ = new_n8360_ & new_n10017_;
  assign new_n14534_ = new_n8360_ & new_n10019_;
  assign new_n14535_ = ~new_n14533_ & ~new_n14534_;
  assign new_n14536_ = new_n14532_ & new_n14535_;
  assign new_n14537_ = new_n14527_ & new_n14536_;
  assign new_n14538_ = new_n14516_ & new_n14537_;
  assign new_n14539_ = new_n14493_ & new_n14538_;
  assign new_n14540_ = new_n8360_ & new_n10030_;
  assign new_n14541_ = new_n8360_ & new_n10015_;
  assign new_n14542_ = new_n8360_ & new_n10028_;
  assign new_n14543_ = ~new_n14541_ & ~new_n14542_;
  assign new_n14544_ = ~new_n14540_ & new_n14543_;
  assign new_n14545_ = new_n8360_ & new_n10039_;
  assign new_n14546_ = new_n8360_ & new_n10026_;
  assign new_n14547_ = new_n8360_ & new_n10037_;
  assign new_n14548_ = ~new_n14546_ & ~new_n14547_;
  assign new_n14549_ = ~new_n14545_ & new_n14548_;
  assign new_n14550_ = new_n14544_ & new_n14549_;
  assign new_n14551_ = new_n8360_ & new_n10048_;
  assign new_n14552_ = new_n8360_ & new_n10035_;
  assign new_n14553_ = new_n8360_ & new_n10046_;
  assign new_n14554_ = ~new_n14552_ & ~new_n14553_;
  assign new_n14555_ = ~new_n14551_ & new_n14554_;
  assign new_n14556_ = new_n8360_ & new_n10054_;
  assign new_n14557_ = new_n8360_ & new_n10044_;
  assign new_n14558_ = new_n8360_ & new_n10052_;
  assign new_n14559_ = ~new_n14557_ & ~new_n14558_;
  assign new_n14560_ = ~new_n14556_ & new_n14559_;
  assign new_n14561_ = new_n14555_ & new_n14560_;
  assign new_n14562_ = new_n14550_ & new_n14561_;
  assign new_n14563_ = new_n8360_ & new_n10061_;
  assign new_n14564_ = new_n8360_ & new_n10063_;
  assign new_n14565_ = new_n8360_ & new_n10065_;
  assign new_n14566_ = ~new_n14564_ & ~new_n14565_;
  assign new_n14567_ = ~new_n14563_ & new_n14566_;
  assign new_n14568_ = new_n8360_ & new_n10069_;
  assign new_n14569_ = new_n8360_ & new_n10071_;
  assign new_n14570_ = new_n8360_ & new_n10073_;
  assign new_n14571_ = ~new_n14569_ & ~new_n14570_;
  assign new_n14572_ = ~new_n14568_ & new_n14571_;
  assign new_n14573_ = new_n14567_ & new_n14572_;
  assign new_n14574_ = new_n8360_ & new_n10078_;
  assign new_n14575_ = new_n8360_ & new_n10080_;
  assign new_n14576_ = new_n8360_ & new_n10082_;
  assign new_n14577_ = ~new_n14575_ & ~new_n14576_;
  assign new_n14578_ = ~new_n14574_ & new_n14577_;
  assign new_n14579_ = new_n8360_ & new_n10089_;
  assign new_n14580_ = new_n8360_ & new_n10091_;
  assign new_n14581_ = ~new_n14579_ & ~new_n14580_;
  assign new_n14582_ = new_n14578_ & new_n14581_;
  assign new_n14583_ = new_n14573_ & new_n14582_;
  assign new_n14584_ = new_n14562_ & new_n14583_;
  assign new_n14585_ = new_n8360_ & new_n10102_;
  assign new_n14586_ = new_n8360_ & new_n10087_;
  assign new_n14587_ = new_n8360_ & new_n10100_;
  assign new_n14588_ = ~new_n14586_ & ~new_n14587_;
  assign new_n14589_ = ~new_n14585_ & new_n14588_;
  assign new_n14590_ = new_n8360_ & new_n10111_;
  assign new_n14591_ = new_n8360_ & new_n10098_;
  assign new_n14592_ = new_n8360_ & new_n10109_;
  assign new_n14593_ = ~new_n14591_ & ~new_n14592_;
  assign new_n14594_ = ~new_n14590_ & new_n14593_;
  assign new_n14595_ = new_n14589_ & new_n14594_;
  assign new_n14596_ = new_n8360_ & new_n10120_;
  assign new_n14597_ = new_n8360_ & new_n10107_;
  assign new_n14598_ = new_n8360_ & new_n10118_;
  assign new_n14599_ = ~new_n14597_ & ~new_n14598_;
  assign new_n14600_ = ~new_n14596_ & new_n14599_;
  assign new_n14601_ = new_n8522_ & new_n9928_;
  assign new_n14602_ = new_n8360_ & new_n10116_;
  assign new_n14603_ = new_n8522_ & new_n9926_;
  assign new_n14604_ = ~new_n14602_ & ~new_n14603_;
  assign new_n14605_ = ~new_n14601_ & new_n14604_;
  assign new_n14606_ = new_n14600_ & new_n14605_;
  assign new_n14607_ = new_n14595_ & new_n14606_;
  assign new_n14608_ = new_n8522_ & new_n9938_;
  assign new_n14609_ = new_n8522_ & new_n9924_;
  assign new_n14610_ = new_n8522_ & new_n9936_;
  assign new_n14611_ = ~new_n14609_ & ~new_n14610_;
  assign new_n14612_ = ~new_n14608_ & new_n14611_;
  assign new_n14613_ = new_n8522_ & new_n9946_;
  assign new_n14614_ = new_n8522_ & new_n9934_;
  assign new_n14615_ = new_n8522_ & new_n9944_;
  assign new_n14616_ = ~new_n14614_ & ~new_n14615_;
  assign new_n14617_ = ~new_n14613_ & new_n14616_;
  assign new_n14618_ = new_n14612_ & new_n14617_;
  assign new_n14619_ = new_n8522_ & new_n9956_;
  assign new_n14620_ = new_n8522_ & new_n9942_;
  assign new_n14621_ = new_n8522_ & new_n9954_;
  assign new_n14622_ = ~new_n14620_ & ~new_n14621_;
  assign new_n14623_ = ~new_n14619_ & new_n14622_;
  assign new_n14624_ = new_n8522_ & new_n9952_;
  assign new_n14625_ = new_n8522_ & new_n9963_;
  assign new_n14626_ = ~new_n14624_ & ~new_n14625_;
  assign new_n14627_ = new_n14623_ & new_n14626_;
  assign new_n14628_ = new_n14618_ & new_n14627_;
  assign new_n14629_ = new_n14607_ & new_n14628_;
  assign new_n14630_ = new_n14584_ & new_n14629_;
  assign new_n14631_ = new_n14539_ & new_n14630_;
  assign new_n14632_ = new_n14448_ & new_n14631_;
  assign new_n14633_ = new_n14265_ & new_n14632_;
  assign new_n14634_ = new_n13896_ & new_n14633_;
  assign new_n14635_ = new_n8522_ & new_n9972_;
  assign new_n14636_ = new_n8522_ & new_n9965_;
  assign new_n14637_ = new_n8522_ & new_n9961_;
  assign new_n14638_ = ~new_n14636_ & ~new_n14637_;
  assign new_n14639_ = ~new_n14635_ & new_n14638_;
  assign new_n14640_ = new_n8522_ & new_n9978_;
  assign new_n14641_ = new_n8522_ & new_n9974_;
  assign new_n14642_ = new_n8522_ & new_n9970_;
  assign new_n14643_ = ~new_n14641_ & ~new_n14642_;
  assign new_n14644_ = ~new_n14640_ & new_n14643_;
  assign new_n14645_ = new_n14639_ & new_n14644_;
  assign new_n14646_ = new_n8522_ & new_n9992_;
  assign new_n14647_ = new_n8522_ & new_n9980_;
  assign new_n14648_ = new_n8522_ & new_n9990_;
  assign new_n14649_ = ~new_n14647_ & ~new_n14648_;
  assign new_n14650_ = ~new_n14646_ & new_n14649_;
  assign new_n14651_ = new_n8522_ & new_n10001_;
  assign new_n14652_ = new_n8522_ & new_n9988_;
  assign new_n14653_ = new_n8522_ & new_n9999_;
  assign new_n14654_ = ~new_n14652_ & ~new_n14653_;
  assign new_n14655_ = ~new_n14651_ & new_n14654_;
  assign new_n14656_ = new_n14650_ & new_n14655_;
  assign new_n14657_ = new_n14645_ & new_n14656_;
  assign new_n14658_ = new_n8522_ & new_n10011_;
  assign new_n14659_ = new_n8522_ & new_n9997_;
  assign new_n14660_ = new_n8522_ & new_n10009_;
  assign new_n14661_ = ~new_n14659_ & ~new_n14660_;
  assign new_n14662_ = ~new_n14658_ & new_n14661_;
  assign new_n14663_ = new_n8522_ & new_n10019_;
  assign new_n14664_ = new_n8522_ & new_n10007_;
  assign new_n14665_ = new_n8522_ & new_n10017_;
  assign new_n14666_ = ~new_n14664_ & ~new_n14665_;
  assign new_n14667_ = ~new_n14663_ & new_n14666_;
  assign new_n14668_ = new_n14662_ & new_n14667_;
  assign new_n14669_ = new_n8522_ & new_n10030_;
  assign new_n14670_ = new_n8522_ & new_n10015_;
  assign new_n14671_ = new_n8522_ & new_n10028_;
  assign new_n14672_ = ~new_n14670_ & ~new_n14671_;
  assign new_n14673_ = ~new_n14669_ & new_n14672_;
  assign new_n14674_ = new_n8522_ & new_n10039_;
  assign new_n14675_ = new_n8522_ & new_n10026_;
  assign new_n14676_ = new_n8522_ & new_n10037_;
  assign new_n14677_ = ~new_n14675_ & ~new_n14676_;
  assign new_n14678_ = ~new_n14674_ & new_n14677_;
  assign new_n14679_ = new_n14673_ & new_n14678_;
  assign new_n14680_ = new_n14668_ & new_n14679_;
  assign new_n14681_ = new_n14657_ & new_n14680_;
  assign new_n14682_ = new_n8522_ & new_n10048_;
  assign new_n14683_ = new_n8522_ & new_n10035_;
  assign new_n14684_ = new_n8522_ & new_n10046_;
  assign new_n14685_ = ~new_n14683_ & ~new_n14684_;
  assign new_n14686_ = ~new_n14682_ & new_n14685_;
  assign new_n14687_ = new_n8522_ & new_n10054_;
  assign new_n14688_ = new_n8522_ & new_n10044_;
  assign new_n14689_ = new_n8522_ & new_n10052_;
  assign new_n14690_ = ~new_n14688_ & ~new_n14689_;
  assign new_n14691_ = ~new_n14687_ & new_n14690_;
  assign new_n14692_ = new_n14686_ & new_n14691_;
  assign new_n14693_ = new_n8522_ & new_n10061_;
  assign new_n14694_ = new_n8522_ & new_n10063_;
  assign new_n14695_ = new_n8522_ & new_n10065_;
  assign new_n14696_ = ~new_n14694_ & ~new_n14695_;
  assign new_n14697_ = ~new_n14693_ & new_n14696_;
  assign new_n14698_ = new_n8522_ & new_n10069_;
  assign new_n14699_ = new_n8522_ & new_n10071_;
  assign new_n14700_ = new_n8522_ & new_n10073_;
  assign new_n14701_ = ~new_n14699_ & ~new_n14700_;
  assign new_n14702_ = ~new_n14698_ & new_n14701_;
  assign new_n14703_ = new_n14697_ & new_n14702_;
  assign new_n14704_ = new_n14692_ & new_n14703_;
  assign new_n14705_ = new_n8522_ & new_n10078_;
  assign new_n14706_ = new_n8522_ & new_n10080_;
  assign new_n14707_ = new_n8522_ & new_n10082_;
  assign new_n14708_ = ~new_n14706_ & ~new_n14707_;
  assign new_n14709_ = ~new_n14705_ & new_n14708_;
  assign new_n14710_ = new_n8522_ & new_n10087_;
  assign new_n14711_ = new_n8522_ & new_n10089_;
  assign new_n14712_ = new_n8522_ & new_n10091_;
  assign new_n14713_ = ~new_n14711_ & ~new_n14712_;
  assign new_n14714_ = ~new_n14710_ & new_n14713_;
  assign new_n14715_ = new_n14709_ & new_n14714_;
  assign new_n14716_ = new_n8522_ & new_n10098_;
  assign new_n14717_ = new_n8522_ & new_n10100_;
  assign new_n14718_ = new_n8522_ & new_n10102_;
  assign new_n14719_ = ~new_n14717_ & ~new_n14718_;
  assign new_n14720_ = ~new_n14716_ & new_n14719_;
  assign new_n14721_ = new_n8522_ & new_n10109_;
  assign new_n14722_ = new_n8522_ & new_n10111_;
  assign new_n14723_ = ~new_n14721_ & ~new_n14722_;
  assign new_n14724_ = new_n14720_ & new_n14723_;
  assign new_n14725_ = new_n14715_ & new_n14724_;
  assign new_n14726_ = new_n14704_ & new_n14725_;
  assign new_n14727_ = new_n14681_ & new_n14726_;
  assign new_n14728_ = new_n8522_ & new_n10120_;
  assign new_n14729_ = new_n8522_ & new_n10107_;
  assign new_n14730_ = new_n8522_ & new_n10118_;
  assign new_n14731_ = ~new_n14729_ & ~new_n14730_;
  assign new_n14732_ = ~new_n14728_ & new_n14731_;
  assign new_n14733_ = ~A199 & new_n10126_;
  assign new_n14734_ = new_n4255_ & new_n14733_;
  assign new_n14735_ = new_n9720_ & new_n14734_;
  assign new_n14736_ = new_n8522_ & new_n10116_;
  assign new_n14737_ = new_n9718_ & new_n14734_;
  assign new_n14738_ = ~new_n14736_ & ~new_n14737_;
  assign new_n14739_ = ~new_n14735_ & new_n14738_;
  assign new_n14740_ = new_n14732_ & new_n14739_;
  assign new_n14741_ = new_n9731_ & new_n14734_;
  assign new_n14742_ = new_n9716_ & new_n14734_;
  assign new_n14743_ = new_n9729_ & new_n14734_;
  assign new_n14744_ = ~new_n14742_ & ~new_n14743_;
  assign new_n14745_ = ~new_n14741_ & new_n14744_;
  assign new_n14746_ = new_n9739_ & new_n14734_;
  assign new_n14747_ = new_n9727_ & new_n14734_;
  assign new_n14748_ = new_n9737_ & new_n14734_;
  assign new_n14749_ = ~new_n14747_ & ~new_n14748_;
  assign new_n14750_ = ~new_n14746_ & new_n14749_;
  assign new_n14751_ = new_n14745_ & new_n14750_;
  assign new_n14752_ = new_n14740_ & new_n14751_;
  assign new_n14753_ = new_n9748_ & new_n14734_;
  assign new_n14754_ = new_n9735_ & new_n14734_;
  assign new_n14755_ = new_n9746_ & new_n14734_;
  assign new_n14756_ = ~new_n14754_ & ~new_n14755_;
  assign new_n14757_ = ~new_n14753_ & new_n14756_;
  assign new_n14758_ = new_n9755_ & new_n14734_;
  assign new_n14759_ = new_n9744_ & new_n14734_;
  assign new_n14760_ = new_n9753_ & new_n14734_;
  assign new_n14761_ = ~new_n14759_ & ~new_n14760_;
  assign new_n14762_ = ~new_n14758_ & new_n14761_;
  assign new_n14763_ = new_n14757_ & new_n14762_;
  assign new_n14764_ = new_n9761_ & new_n14734_;
  assign new_n14765_ = new_n9763_ & new_n14734_;
  assign new_n14766_ = new_n9765_ & new_n14734_;
  assign new_n14767_ = ~new_n14765_ & ~new_n14766_;
  assign new_n14768_ = ~new_n14764_ & new_n14767_;
  assign new_n14769_ = new_n9771_ & new_n14734_;
  assign new_n14770_ = new_n9773_ & new_n14734_;
  assign new_n14771_ = ~new_n14769_ & ~new_n14770_;
  assign new_n14772_ = new_n14768_ & new_n14771_;
  assign new_n14773_ = new_n14763_ & new_n14772_;
  assign new_n14774_ = new_n14752_ & new_n14773_;
  assign new_n14775_ = new_n9783_ & new_n14734_;
  assign new_n14776_ = new_n9769_ & new_n14734_;
  assign new_n14777_ = new_n9781_ & new_n14734_;
  assign new_n14778_ = ~new_n14776_ & ~new_n14777_;
  assign new_n14779_ = ~new_n14775_ & new_n14778_;
  assign new_n14780_ = new_n9792_ & new_n14734_;
  assign new_n14781_ = new_n9779_ & new_n14734_;
  assign new_n14782_ = new_n9790_ & new_n14734_;
  assign new_n14783_ = ~new_n14781_ & ~new_n14782_;
  assign new_n14784_ = ~new_n14780_ & new_n14783_;
  assign new_n14785_ = new_n14779_ & new_n14784_;
  assign new_n14786_ = new_n9803_ & new_n14734_;
  assign new_n14787_ = new_n9788_ & new_n14734_;
  assign new_n14788_ = new_n9801_ & new_n14734_;
  assign new_n14789_ = ~new_n14787_ & ~new_n14788_;
  assign new_n14790_ = ~new_n14786_ & new_n14789_;
  assign new_n14791_ = new_n9811_ & new_n14734_;
  assign new_n14792_ = new_n9799_ & new_n14734_;
  assign new_n14793_ = new_n9809_ & new_n14734_;
  assign new_n14794_ = ~new_n14792_ & ~new_n14793_;
  assign new_n14795_ = ~new_n14791_ & new_n14794_;
  assign new_n14796_ = new_n14790_ & new_n14795_;
  assign new_n14797_ = new_n14785_ & new_n14796_;
  assign new_n14798_ = ~A199 & new_n10141_;
  assign new_n14799_ = new_n4255_ & new_n14798_;
  assign new_n14800_ = new_n9821_ & new_n14799_;
  assign new_n14801_ = new_n9807_ & new_n14734_;
  assign new_n14802_ = new_n9819_ & new_n14799_;
  assign new_n14803_ = ~new_n14801_ & ~new_n14802_;
  assign new_n14804_ = ~new_n14800_ & new_n14803_;
  assign new_n14805_ = new_n9828_ & new_n14799_;
  assign new_n14806_ = new_n9817_ & new_n14799_;
  assign new_n14807_ = new_n9825_ & new_n14799_;
  assign new_n14808_ = ~new_n14806_ & ~new_n14807_;
  assign new_n14809_ = ~new_n14805_ & new_n14808_;
  assign new_n14810_ = new_n14804_ & new_n14809_;
  assign new_n14811_ = new_n9840_ & new_n14799_;
  assign new_n14812_ = new_n9842_ & new_n14799_;
  assign new_n14813_ = new_n9844_ & new_n14799_;
  assign new_n14814_ = ~new_n14812_ & ~new_n14813_;
  assign new_n14815_ = ~new_n14811_ & new_n14814_;
  assign new_n14816_ = new_n9850_ & new_n14799_;
  assign new_n14817_ = new_n9852_ & new_n14799_;
  assign new_n14818_ = ~new_n14816_ & ~new_n14817_;
  assign new_n14819_ = new_n14815_ & new_n14818_;
  assign new_n14820_ = new_n14810_ & new_n14819_;
  assign new_n14821_ = new_n14797_ & new_n14820_;
  assign new_n14822_ = new_n14774_ & new_n14821_;
  assign new_n14823_ = new_n14727_ & new_n14822_;
  assign new_n14824_ = new_n9862_ & new_n14799_;
  assign new_n14825_ = new_n9848_ & new_n14799_;
  assign new_n14826_ = new_n9860_ & new_n14799_;
  assign new_n14827_ = ~new_n14825_ & ~new_n14826_;
  assign new_n14828_ = ~new_n14824_ & new_n14827_;
  assign new_n14829_ = new_n9870_ & new_n14799_;
  assign new_n14830_ = new_n9858_ & new_n14799_;
  assign new_n14831_ = new_n9868_ & new_n14799_;
  assign new_n14832_ = ~new_n14830_ & ~new_n14831_;
  assign new_n14833_ = ~new_n14829_ & new_n14832_;
  assign new_n14834_ = new_n14828_ & new_n14833_;
  assign new_n14835_ = new_n9880_ & new_n14799_;
  assign new_n14836_ = new_n9866_ & new_n14799_;
  assign new_n14837_ = new_n9878_ & new_n14799_;
  assign new_n14838_ = ~new_n14836_ & ~new_n14837_;
  assign new_n14839_ = ~new_n14835_ & new_n14838_;
  assign new_n14840_ = new_n9889_ & new_n14799_;
  assign new_n14841_ = new_n9876_ & new_n14799_;
  assign new_n14842_ = new_n9887_ & new_n14799_;
  assign new_n14843_ = ~new_n14841_ & ~new_n14842_;
  assign new_n14844_ = ~new_n14840_ & new_n14843_;
  assign new_n14845_ = new_n14839_ & new_n14844_;
  assign new_n14846_ = new_n14834_ & new_n14845_;
  assign new_n14847_ = new_n9899_ & new_n14799_;
  assign new_n14848_ = new_n9885_ & new_n14799_;
  assign new_n14849_ = new_n9897_ & new_n14799_;
  assign new_n14850_ = ~new_n14848_ & ~new_n14849_;
  assign new_n14851_ = ~new_n14847_ & new_n14850_;
  assign new_n14852_ = new_n9908_ & new_n14799_;
  assign new_n14853_ = new_n9895_ & new_n14799_;
  assign new_n14854_ = new_n9906_ & new_n14799_;
  assign new_n14855_ = ~new_n14853_ & ~new_n14854_;
  assign new_n14856_ = ~new_n14852_ & new_n14855_;
  assign new_n14857_ = new_n14851_ & new_n14856_;
  assign new_n14858_ = new_n9919_ & new_n14799_;
  assign new_n14859_ = new_n9904_ & new_n14799_;
  assign new_n14860_ = new_n9917_ & new_n14799_;
  assign new_n14861_ = ~new_n14859_ & ~new_n14860_;
  assign new_n14862_ = ~new_n14858_ & new_n14861_;
  assign new_n14863_ = new_n9915_ & new_n14799_;
  assign new_n14864_ = ~A199 & new_n10165_;
  assign new_n14865_ = new_n4255_ & new_n14864_;
  assign new_n14866_ = new_n9926_ & new_n14865_;
  assign new_n14867_ = ~new_n14863_ & ~new_n14866_;
  assign new_n14868_ = new_n14862_ & new_n14867_;
  assign new_n14869_ = new_n14857_ & new_n14868_;
  assign new_n14870_ = new_n14846_ & new_n14869_;
  assign new_n14871_ = new_n9936_ & new_n14865_;
  assign new_n14872_ = new_n9928_ & new_n14865_;
  assign new_n14873_ = new_n9924_ & new_n14865_;
  assign new_n14874_ = ~new_n14872_ & ~new_n14873_;
  assign new_n14875_ = ~new_n14871_ & new_n14874_;
  assign new_n14876_ = new_n9944_ & new_n14865_;
  assign new_n14877_ = new_n9938_ & new_n14865_;
  assign new_n14878_ = new_n9934_ & new_n14865_;
  assign new_n14879_ = ~new_n14877_ & ~new_n14878_;
  assign new_n14880_ = ~new_n14876_ & new_n14879_;
  assign new_n14881_ = new_n14875_ & new_n14880_;
  assign new_n14882_ = new_n9954_ & new_n14865_;
  assign new_n14883_ = new_n9946_ & new_n14865_;
  assign new_n14884_ = new_n9942_ & new_n14865_;
  assign new_n14885_ = ~new_n14883_ & ~new_n14884_;
  assign new_n14886_ = ~new_n14882_ & new_n14885_;
  assign new_n14887_ = new_n9963_ & new_n14865_;
  assign new_n14888_ = new_n9956_ & new_n14865_;
  assign new_n14889_ = new_n9952_ & new_n14865_;
  assign new_n14890_ = ~new_n14888_ & ~new_n14889_;
  assign new_n14891_ = ~new_n14887_ & new_n14890_;
  assign new_n14892_ = new_n14886_ & new_n14891_;
  assign new_n14893_ = new_n14881_ & new_n14892_;
  assign new_n14894_ = new_n9972_ & new_n14865_;
  assign new_n14895_ = new_n9965_ & new_n14865_;
  assign new_n14896_ = new_n9961_ & new_n14865_;
  assign new_n14897_ = ~new_n14895_ & ~new_n14896_;
  assign new_n14898_ = ~new_n14894_ & new_n14897_;
  assign new_n14899_ = new_n9978_ & new_n14865_;
  assign new_n14900_ = new_n9974_ & new_n14865_;
  assign new_n14901_ = new_n9970_ & new_n14865_;
  assign new_n14902_ = ~new_n14900_ & ~new_n14901_;
  assign new_n14903_ = ~new_n14899_ & new_n14902_;
  assign new_n14904_ = new_n14898_ & new_n14903_;
  assign new_n14905_ = new_n9992_ & new_n14865_;
  assign new_n14906_ = new_n9980_ & new_n14865_;
  assign new_n14907_ = new_n9990_ & new_n14865_;
  assign new_n14908_ = ~new_n14906_ & ~new_n14907_;
  assign new_n14909_ = ~new_n14905_ & new_n14908_;
  assign new_n14910_ = new_n9988_ & new_n14865_;
  assign new_n14911_ = new_n9999_ & new_n14865_;
  assign new_n14912_ = ~new_n14910_ & ~new_n14911_;
  assign new_n14913_ = new_n14909_ & new_n14912_;
  assign new_n14914_ = new_n14904_ & new_n14913_;
  assign new_n14915_ = new_n14893_ & new_n14914_;
  assign new_n14916_ = new_n14870_ & new_n14915_;
  assign new_n14917_ = new_n10009_ & new_n14865_;
  assign new_n14918_ = new_n10001_ & new_n14865_;
  assign new_n14919_ = new_n9997_ & new_n14865_;
  assign new_n14920_ = ~new_n14918_ & ~new_n14919_;
  assign new_n14921_ = ~new_n14917_ & new_n14920_;
  assign new_n14922_ = new_n10017_ & new_n14865_;
  assign new_n14923_ = new_n10011_ & new_n14865_;
  assign new_n14924_ = new_n10007_ & new_n14865_;
  assign new_n14925_ = ~new_n14923_ & ~new_n14924_;
  assign new_n14926_ = ~new_n14922_ & new_n14925_;
  assign new_n14927_ = new_n14921_ & new_n14926_;
  assign new_n14928_ = new_n10028_ & new_n14865_;
  assign new_n14929_ = new_n10019_ & new_n14865_;
  assign new_n14930_ = new_n10015_ & new_n14865_;
  assign new_n14931_ = ~new_n14929_ & ~new_n14930_;
  assign new_n14932_ = ~new_n14928_ & new_n14931_;
  assign new_n14933_ = new_n10037_ & new_n14865_;
  assign new_n14934_ = new_n10030_ & new_n14865_;
  assign new_n14935_ = new_n10026_ & new_n14865_;
  assign new_n14936_ = ~new_n14934_ & ~new_n14935_;
  assign new_n14937_ = ~new_n14933_ & new_n14936_;
  assign new_n14938_ = new_n14932_ & new_n14937_;
  assign new_n14939_ = new_n14927_ & new_n14938_;
  assign new_n14940_ = new_n10046_ & new_n14865_;
  assign new_n14941_ = new_n10039_ & new_n14865_;
  assign new_n14942_ = new_n10035_ & new_n14865_;
  assign new_n14943_ = ~new_n14941_ & ~new_n14942_;
  assign new_n14944_ = ~new_n14940_ & new_n14943_;
  assign new_n14945_ = new_n10052_ & new_n14865_;
  assign new_n14946_ = new_n10048_ & new_n14865_;
  assign new_n14947_ = new_n10044_ & new_n14865_;
  assign new_n14948_ = ~new_n14946_ & ~new_n14947_;
  assign new_n14949_ = ~new_n14945_ & new_n14948_;
  assign new_n14950_ = new_n14944_ & new_n14949_;
  assign new_n14951_ = new_n10065_ & new_n14865_;
  assign new_n14952_ = new_n10054_ & new_n14865_;
  assign new_n14953_ = new_n10063_ & new_n14865_;
  assign new_n14954_ = ~new_n14952_ & ~new_n14953_;
  assign new_n14955_ = ~new_n14951_ & new_n14954_;
  assign new_n14956_ = new_n10061_ & new_n14865_;
  assign new_n14957_ = new_n10071_ & new_n14865_;
  assign new_n14958_ = ~new_n14956_ & ~new_n14957_;
  assign new_n14959_ = new_n14955_ & new_n14958_;
  assign new_n14960_ = new_n14950_ & new_n14959_;
  assign new_n14961_ = new_n14939_ & new_n14960_;
  assign new_n14962_ = new_n10080_ & new_n14865_;
  assign new_n14963_ = new_n10073_ & new_n14865_;
  assign new_n14964_ = new_n10069_ & new_n14865_;
  assign new_n14965_ = ~new_n14963_ & ~new_n14964_;
  assign new_n14966_ = ~new_n14962_ & new_n14965_;
  assign new_n14967_ = new_n10089_ & new_n14865_;
  assign new_n14968_ = new_n10082_ & new_n14865_;
  assign new_n14969_ = new_n10078_ & new_n14865_;
  assign new_n14970_ = ~new_n14968_ & ~new_n14969_;
  assign new_n14971_ = ~new_n14967_ & new_n14970_;
  assign new_n14972_ = new_n14966_ & new_n14971_;
  assign new_n14973_ = new_n10100_ & new_n14865_;
  assign new_n14974_ = new_n10091_ & new_n14865_;
  assign new_n14975_ = new_n10087_ & new_n14865_;
  assign new_n14976_ = ~new_n14974_ & ~new_n14975_;
  assign new_n14977_ = ~new_n14973_ & new_n14976_;
  assign new_n14978_ = new_n10109_ & new_n14865_;
  assign new_n14979_ = new_n10102_ & new_n14865_;
  assign new_n14980_ = new_n10098_ & new_n14865_;
  assign new_n14981_ = ~new_n14979_ & ~new_n14980_;
  assign new_n14982_ = ~new_n14978_ & new_n14981_;
  assign new_n14983_ = new_n14977_ & new_n14982_;
  assign new_n14984_ = new_n14972_ & new_n14983_;
  assign new_n14985_ = new_n10118_ & new_n14865_;
  assign new_n14986_ = new_n10111_ & new_n14865_;
  assign new_n14987_ = new_n10107_ & new_n14865_;
  assign new_n14988_ = ~new_n14986_ & ~new_n14987_;
  assign new_n14989_ = ~new_n14985_ & new_n14988_;
  assign new_n14990_ = A199 & new_n10240_;
  assign new_n14991_ = new_n4255_ & new_n14990_;
  assign new_n14992_ = new_n9718_ & new_n14991_;
  assign new_n14993_ = new_n10120_ & new_n14865_;
  assign new_n14994_ = new_n10116_ & new_n14865_;
  assign new_n14995_ = ~new_n14993_ & ~new_n14994_;
  assign new_n14996_ = ~new_n14992_ & new_n14995_;
  assign new_n14997_ = new_n14989_ & new_n14996_;
  assign new_n14998_ = new_n9729_ & new_n14991_;
  assign new_n14999_ = new_n9720_ & new_n14991_;
  assign new_n15000_ = new_n9716_ & new_n14991_;
  assign new_n15001_ = ~new_n14999_ & ~new_n15000_;
  assign new_n15002_ = ~new_n14998_ & new_n15001_;
  assign new_n15003_ = new_n9731_ & new_n14991_;
  assign new_n15004_ = new_n9727_ & new_n14991_;
  assign new_n15005_ = ~new_n15003_ & ~new_n15004_;
  assign new_n15006_ = new_n15002_ & new_n15005_;
  assign new_n15007_ = new_n14997_ & new_n15006_;
  assign new_n15008_ = new_n14984_ & new_n15007_;
  assign new_n15009_ = new_n14961_ & new_n15008_;
  assign new_n15010_ = new_n14916_ & new_n15009_;
  assign new_n15011_ = new_n14823_ & new_n15010_;
  assign new_n15012_ = new_n9735_ & new_n14991_;
  assign new_n15013_ = new_n9737_ & new_n14991_;
  assign new_n15014_ = new_n9739_ & new_n14991_;
  assign new_n15015_ = ~new_n15013_ & ~new_n15014_;
  assign new_n15016_ = ~new_n15012_ & new_n15015_;
  assign new_n15017_ = new_n9744_ & new_n14991_;
  assign new_n15018_ = new_n9746_ & new_n14991_;
  assign new_n15019_ = new_n9748_ & new_n14991_;
  assign new_n15020_ = ~new_n15018_ & ~new_n15019_;
  assign new_n15021_ = ~new_n15017_ & new_n15020_;
  assign new_n15022_ = new_n15016_ & new_n15021_;
  assign new_n15023_ = new_n9763_ & new_n14991_;
  assign new_n15024_ = new_n9753_ & new_n14991_;
  assign new_n15025_ = new_n9755_ & new_n14991_;
  assign new_n15026_ = ~new_n15024_ & ~new_n15025_;
  assign new_n15027_ = ~new_n15023_ & new_n15026_;
  assign new_n15028_ = new_n9771_ & new_n14991_;
  assign new_n15029_ = new_n9765_ & new_n14991_;
  assign new_n15030_ = new_n9761_ & new_n14991_;
  assign new_n15031_ = ~new_n15029_ & ~new_n15030_;
  assign new_n15032_ = ~new_n15028_ & new_n15031_;
  assign new_n15033_ = new_n15027_ & new_n15032_;
  assign new_n15034_ = new_n15022_ & new_n15033_;
  assign new_n15035_ = new_n9781_ & new_n14991_;
  assign new_n15036_ = new_n9773_ & new_n14991_;
  assign new_n15037_ = new_n9769_ & new_n14991_;
  assign new_n15038_ = ~new_n15036_ & ~new_n15037_;
  assign new_n15039_ = ~new_n15035_ & new_n15038_;
  assign new_n15040_ = new_n9790_ & new_n14991_;
  assign new_n15041_ = new_n9783_ & new_n14991_;
  assign new_n15042_ = new_n9779_ & new_n14991_;
  assign new_n15043_ = ~new_n15041_ & ~new_n15042_;
  assign new_n15044_ = ~new_n15040_ & new_n15043_;
  assign new_n15045_ = new_n15039_ & new_n15044_;
  assign new_n15046_ = new_n9801_ & new_n14991_;
  assign new_n15047_ = new_n9792_ & new_n14991_;
  assign new_n15048_ = new_n9788_ & new_n14991_;
  assign new_n15049_ = ~new_n15047_ & ~new_n15048_;
  assign new_n15050_ = ~new_n15046_ & new_n15049_;
  assign new_n15051_ = new_n9809_ & new_n14991_;
  assign new_n15052_ = new_n9803_ & new_n14991_;
  assign new_n15053_ = new_n9799_ & new_n14991_;
  assign new_n15054_ = ~new_n15052_ & ~new_n15053_;
  assign new_n15055_ = ~new_n15051_ & new_n15054_;
  assign new_n15056_ = new_n15050_ & new_n15055_;
  assign new_n15057_ = new_n15045_ & new_n15056_;
  assign new_n15058_ = new_n15034_ & new_n15057_;
  assign new_n15059_ = A199 & new_n10253_;
  assign new_n15060_ = new_n4255_ & new_n15059_;
  assign new_n15061_ = new_n9819_ & new_n15060_;
  assign new_n15062_ = new_n9811_ & new_n14991_;
  assign new_n15063_ = new_n9807_ & new_n14991_;
  assign new_n15064_ = ~new_n15062_ & ~new_n15063_;
  assign new_n15065_ = ~new_n15061_ & new_n15064_;
  assign new_n15066_ = new_n9825_ & new_n15060_;
  assign new_n15067_ = new_n9821_ & new_n15060_;
  assign new_n15068_ = new_n9817_ & new_n15060_;
  assign new_n15069_ = ~new_n15067_ & ~new_n15068_;
  assign new_n15070_ = ~new_n15066_ & new_n15069_;
  assign new_n15071_ = new_n15065_ & new_n15070_;
  assign new_n15072_ = new_n9844_ & new_n15060_;
  assign new_n15073_ = new_n9828_ & new_n15060_;
  assign new_n15074_ = new_n9842_ & new_n15060_;
  assign new_n15075_ = ~new_n15073_ & ~new_n15074_;
  assign new_n15076_ = ~new_n15072_ & new_n15075_;
  assign new_n15077_ = new_n9852_ & new_n15060_;
  assign new_n15078_ = new_n9840_ & new_n15060_;
  assign new_n15079_ = new_n9850_ & new_n15060_;
  assign new_n15080_ = ~new_n15078_ & ~new_n15079_;
  assign new_n15081_ = ~new_n15077_ & new_n15080_;
  assign new_n15082_ = new_n15076_ & new_n15081_;
  assign new_n15083_ = new_n15071_ & new_n15082_;
  assign new_n15084_ = new_n9862_ & new_n15060_;
  assign new_n15085_ = new_n9848_ & new_n15060_;
  assign new_n15086_ = new_n9860_ & new_n15060_;
  assign new_n15087_ = ~new_n15085_ & ~new_n15086_;
  assign new_n15088_ = ~new_n15084_ & new_n15087_;
  assign new_n15089_ = new_n9870_ & new_n15060_;
  assign new_n15090_ = new_n9858_ & new_n15060_;
  assign new_n15091_ = new_n9868_ & new_n15060_;
  assign new_n15092_ = ~new_n15090_ & ~new_n15091_;
  assign new_n15093_ = ~new_n15089_ & new_n15092_;
  assign new_n15094_ = new_n15088_ & new_n15093_;
  assign new_n15095_ = new_n9880_ & new_n15060_;
  assign new_n15096_ = new_n9866_ & new_n15060_;
  assign new_n15097_ = new_n9878_ & new_n15060_;
  assign new_n15098_ = ~new_n15096_ & ~new_n15097_;
  assign new_n15099_ = ~new_n15095_ & new_n15098_;
  assign new_n15100_ = new_n9876_ & new_n15060_;
  assign new_n15101_ = new_n9887_ & new_n15060_;
  assign new_n15102_ = ~new_n15100_ & ~new_n15101_;
  assign new_n15103_ = new_n15099_ & new_n15102_;
  assign new_n15104_ = new_n15094_ & new_n15103_;
  assign new_n15105_ = new_n15083_ & new_n15104_;
  assign new_n15106_ = new_n15058_ & new_n15105_;
  assign new_n15107_ = new_n9897_ & new_n15060_;
  assign new_n15108_ = new_n9889_ & new_n15060_;
  assign new_n15109_ = new_n9885_ & new_n15060_;
  assign new_n15110_ = ~new_n15108_ & ~new_n15109_;
  assign new_n15111_ = ~new_n15107_ & new_n15110_;
  assign new_n15112_ = new_n9906_ & new_n15060_;
  assign new_n15113_ = new_n9899_ & new_n15060_;
  assign new_n15114_ = new_n9895_ & new_n15060_;
  assign new_n15115_ = ~new_n15113_ & ~new_n15114_;
  assign new_n15116_ = ~new_n15112_ & new_n15115_;
  assign new_n15117_ = new_n15111_ & new_n15116_;
  assign new_n15118_ = new_n9917_ & new_n15060_;
  assign new_n15119_ = new_n9908_ & new_n15060_;
  assign new_n15120_ = new_n9904_ & new_n15060_;
  assign new_n15121_ = ~new_n15119_ & ~new_n15120_;
  assign new_n15122_ = ~new_n15118_ & new_n15121_;
  assign new_n15123_ = A199 & new_n10272_;
  assign new_n15124_ = new_n4255_ & new_n15123_;
  assign new_n15125_ = new_n9926_ & new_n15124_;
  assign new_n15126_ = new_n9919_ & new_n15060_;
  assign new_n15127_ = new_n9915_ & new_n15060_;
  assign new_n15128_ = ~new_n15126_ & ~new_n15127_;
  assign new_n15129_ = ~new_n15125_ & new_n15128_;
  assign new_n15130_ = new_n15122_ & new_n15129_;
  assign new_n15131_ = new_n15117_ & new_n15130_;
  assign new_n15132_ = new_n9936_ & new_n15124_;
  assign new_n15133_ = new_n9928_ & new_n15124_;
  assign new_n15134_ = new_n9924_ & new_n15124_;
  assign new_n15135_ = ~new_n15133_ & ~new_n15134_;
  assign new_n15136_ = ~new_n15132_ & new_n15135_;
  assign new_n15137_ = new_n9944_ & new_n15124_;
  assign new_n15138_ = new_n9938_ & new_n15124_;
  assign new_n15139_ = new_n9934_ & new_n15124_;
  assign new_n15140_ = ~new_n15138_ & ~new_n15139_;
  assign new_n15141_ = ~new_n15137_ & new_n15140_;
  assign new_n15142_ = new_n15136_ & new_n15141_;
  assign new_n15143_ = new_n9954_ & new_n15124_;
  assign new_n15144_ = new_n9946_ & new_n15124_;
  assign new_n15145_ = new_n9942_ & new_n15124_;
  assign new_n15146_ = ~new_n15144_ & ~new_n15145_;
  assign new_n15147_ = ~new_n15143_ & new_n15146_;
  assign new_n15148_ = new_n9956_ & new_n15124_;
  assign new_n15149_ = new_n9952_ & new_n15124_;
  assign new_n15150_ = ~new_n15148_ & ~new_n15149_;
  assign new_n15151_ = new_n15147_ & new_n15150_;
  assign new_n15152_ = new_n15142_ & new_n15151_;
  assign new_n15153_ = new_n15131_ & new_n15152_;
  assign new_n15154_ = new_n9961_ & new_n15124_;
  assign new_n15155_ = new_n9963_ & new_n15124_;
  assign new_n15156_ = new_n9965_ & new_n15124_;
  assign new_n15157_ = ~new_n15155_ & ~new_n15156_;
  assign new_n15158_ = ~new_n15154_ & new_n15157_;
  assign new_n15159_ = new_n9970_ & new_n15124_;
  assign new_n15160_ = new_n9972_ & new_n15124_;
  assign new_n15161_ = new_n9974_ & new_n15124_;
  assign new_n15162_ = ~new_n15160_ & ~new_n15161_;
  assign new_n15163_ = ~new_n15159_ & new_n15162_;
  assign new_n15164_ = new_n15158_ & new_n15163_;
  assign new_n15165_ = new_n9990_ & new_n15124_;
  assign new_n15166_ = new_n9978_ & new_n15124_;
  assign new_n15167_ = new_n9980_ & new_n15124_;
  assign new_n15168_ = ~new_n15166_ & ~new_n15167_;
  assign new_n15169_ = ~new_n15165_ & new_n15168_;
  assign new_n15170_ = new_n9999_ & new_n15124_;
  assign new_n15171_ = new_n9992_ & new_n15124_;
  assign new_n15172_ = new_n9988_ & new_n15124_;
  assign new_n15173_ = ~new_n15171_ & ~new_n15172_;
  assign new_n15174_ = ~new_n15170_ & new_n15173_;
  assign new_n15175_ = new_n15169_ & new_n15174_;
  assign new_n15176_ = new_n15164_ & new_n15175_;
  assign new_n15177_ = new_n10009_ & new_n15124_;
  assign new_n15178_ = new_n10001_ & new_n15124_;
  assign new_n15179_ = new_n9997_ & new_n15124_;
  assign new_n15180_ = ~new_n15178_ & ~new_n15179_;
  assign new_n15181_ = ~new_n15177_ & new_n15180_;
  assign new_n15182_ = new_n10017_ & new_n15124_;
  assign new_n15183_ = new_n10011_ & new_n15124_;
  assign new_n15184_ = new_n10007_ & new_n15124_;
  assign new_n15185_ = ~new_n15183_ & ~new_n15184_;
  assign new_n15186_ = ~new_n15182_ & new_n15185_;
  assign new_n15187_ = new_n15181_ & new_n15186_;
  assign new_n15188_ = new_n10028_ & new_n15124_;
  assign new_n15189_ = new_n10019_ & new_n15124_;
  assign new_n15190_ = new_n10015_ & new_n15124_;
  assign new_n15191_ = ~new_n15189_ & ~new_n15190_;
  assign new_n15192_ = ~new_n15188_ & new_n15191_;
  assign new_n15193_ = new_n10030_ & new_n15124_;
  assign new_n15194_ = new_n10026_ & new_n15124_;
  assign new_n15195_ = ~new_n15193_ & ~new_n15194_;
  assign new_n15196_ = new_n15192_ & new_n15195_;
  assign new_n15197_ = new_n15187_ & new_n15196_;
  assign new_n15198_ = new_n15176_ & new_n15197_;
  assign new_n15199_ = new_n15153_ & new_n15198_;
  assign new_n15200_ = new_n15106_ & new_n15199_;
  assign new_n15201_ = new_n10035_ & new_n15124_;
  assign new_n15202_ = new_n10037_ & new_n15124_;
  assign new_n15203_ = new_n10039_ & new_n15124_;
  assign new_n15204_ = ~new_n15202_ & ~new_n15203_;
  assign new_n15205_ = ~new_n15201_ & new_n15204_;
  assign new_n15206_ = new_n10044_ & new_n15124_;
  assign new_n15207_ = new_n10046_ & new_n15124_;
  assign new_n15208_ = new_n10048_ & new_n15124_;
  assign new_n15209_ = ~new_n15207_ & ~new_n15208_;
  assign new_n15210_ = ~new_n15206_ & new_n15209_;
  assign new_n15211_ = new_n15205_ & new_n15210_;
  assign new_n15212_ = new_n10063_ & new_n15124_;
  assign new_n15213_ = new_n10052_ & new_n15124_;
  assign new_n15214_ = new_n10054_ & new_n15124_;
  assign new_n15215_ = ~new_n15213_ & ~new_n15214_;
  assign new_n15216_ = ~new_n15212_ & new_n15215_;
  assign new_n15217_ = new_n10071_ & new_n15124_;
  assign new_n15218_ = new_n10065_ & new_n15124_;
  assign new_n15219_ = new_n10061_ & new_n15124_;
  assign new_n15220_ = ~new_n15218_ & ~new_n15219_;
  assign new_n15221_ = ~new_n15217_ & new_n15220_;
  assign new_n15222_ = new_n15216_ & new_n15221_;
  assign new_n15223_ = new_n15211_ & new_n15222_;
  assign new_n15224_ = new_n10080_ & new_n15124_;
  assign new_n15225_ = new_n10073_ & new_n15124_;
  assign new_n15226_ = new_n10069_ & new_n15124_;
  assign new_n15227_ = ~new_n15225_ & ~new_n15226_;
  assign new_n15228_ = ~new_n15224_ & new_n15227_;
  assign new_n15229_ = new_n10089_ & new_n15124_;
  assign new_n15230_ = new_n10082_ & new_n15124_;
  assign new_n15231_ = new_n10078_ & new_n15124_;
  assign new_n15232_ = ~new_n15230_ & ~new_n15231_;
  assign new_n15233_ = ~new_n15229_ & new_n15232_;
  assign new_n15234_ = new_n15228_ & new_n15233_;
  assign new_n15235_ = new_n10100_ & new_n15124_;
  assign new_n15236_ = new_n10091_ & new_n15124_;
  assign new_n15237_ = new_n10087_ & new_n15124_;
  assign new_n15238_ = ~new_n15236_ & ~new_n15237_;
  assign new_n15239_ = ~new_n15235_ & new_n15238_;
  assign new_n15240_ = new_n10102_ & new_n15124_;
  assign new_n15241_ = new_n10098_ & new_n15124_;
  assign new_n15242_ = ~new_n15240_ & ~new_n15241_;
  assign new_n15243_ = new_n15239_ & new_n15242_;
  assign new_n15244_ = new_n15234_ & new_n15243_;
  assign new_n15245_ = new_n15223_ & new_n15244_;
  assign new_n15246_ = new_n10107_ & new_n15124_;
  assign new_n15247_ = new_n10109_ & new_n15124_;
  assign new_n15248_ = new_n10111_ & new_n15124_;
  assign new_n15249_ = ~new_n15247_ & ~new_n15248_;
  assign new_n15250_ = ~new_n15246_ & new_n15249_;
  assign new_n15251_ = new_n10116_ & new_n15124_;
  assign new_n15252_ = new_n10118_ & new_n15124_;
  assign new_n15253_ = new_n10120_ & new_n15124_;
  assign new_n15254_ = ~new_n15252_ & ~new_n15253_;
  assign new_n15255_ = ~new_n15251_ & new_n15254_;
  assign new_n15256_ = new_n15250_ & new_n15255_;
  assign new_n15257_ = ~A201 & new_n7214_;
  assign new_n15258_ = new_n4255_ & new_n15257_;
  assign new_n15259_ = new_n9716_ & new_n15258_;
  assign new_n15260_ = new_n9718_ & new_n15258_;
  assign new_n15261_ = new_n9720_ & new_n15258_;
  assign new_n15262_ = ~new_n15260_ & ~new_n15261_;
  assign new_n15263_ = ~new_n15259_ & new_n15262_;
  assign new_n15264_ = new_n9727_ & new_n15258_;
  assign new_n15265_ = new_n9729_ & new_n15258_;
  assign new_n15266_ = new_n9731_ & new_n15258_;
  assign new_n15267_ = ~new_n15265_ & ~new_n15266_;
  assign new_n15268_ = ~new_n15264_ & new_n15267_;
  assign new_n15269_ = new_n15263_ & new_n15268_;
  assign new_n15270_ = new_n15256_ & new_n15269_;
  assign new_n15271_ = new_n9735_ & new_n15258_;
  assign new_n15272_ = new_n9737_ & new_n15258_;
  assign new_n15273_ = new_n9739_ & new_n15258_;
  assign new_n15274_ = ~new_n15272_ & ~new_n15273_;
  assign new_n15275_ = ~new_n15271_ & new_n15274_;
  assign new_n15276_ = new_n9744_ & new_n15258_;
  assign new_n15277_ = new_n9746_ & new_n15258_;
  assign new_n15278_ = new_n9748_ & new_n15258_;
  assign new_n15279_ = ~new_n15277_ & ~new_n15278_;
  assign new_n15280_ = ~new_n15276_ & new_n15279_;
  assign new_n15281_ = new_n15275_ & new_n15280_;
  assign new_n15282_ = new_n9763_ & new_n15258_;
  assign new_n15283_ = new_n9753_ & new_n15258_;
  assign new_n15284_ = new_n9755_ & new_n15258_;
  assign new_n15285_ = ~new_n15283_ & ~new_n15284_;
  assign new_n15286_ = ~new_n15282_ & new_n15285_;
  assign new_n15287_ = new_n9765_ & new_n15258_;
  assign new_n15288_ = new_n9761_ & new_n15258_;
  assign new_n15289_ = ~new_n15287_ & ~new_n15288_;
  assign new_n15290_ = new_n15286_ & new_n15289_;
  assign new_n15291_ = new_n15281_ & new_n15290_;
  assign new_n15292_ = new_n15270_ & new_n15291_;
  assign new_n15293_ = new_n15245_ & new_n15292_;
  assign new_n15294_ = new_n9769_ & new_n15258_;
  assign new_n15295_ = new_n9771_ & new_n15258_;
  assign new_n15296_ = new_n9773_ & new_n15258_;
  assign new_n15297_ = ~new_n15295_ & ~new_n15296_;
  assign new_n15298_ = ~new_n15294_ & new_n15297_;
  assign new_n15299_ = new_n9779_ & new_n15258_;
  assign new_n15300_ = new_n9781_ & new_n15258_;
  assign new_n15301_ = new_n9783_ & new_n15258_;
  assign new_n15302_ = ~new_n15300_ & ~new_n15301_;
  assign new_n15303_ = ~new_n15299_ & new_n15302_;
  assign new_n15304_ = new_n15298_ & new_n15303_;
  assign new_n15305_ = new_n9788_ & new_n15258_;
  assign new_n15306_ = new_n9790_ & new_n15258_;
  assign new_n15307_ = new_n9792_ & new_n15258_;
  assign new_n15308_ = ~new_n15306_ & ~new_n15307_;
  assign new_n15309_ = ~new_n15305_ & new_n15308_;
  assign new_n15310_ = new_n9799_ & new_n15258_;
  assign new_n15311_ = new_n9801_ & new_n15258_;
  assign new_n15312_ = new_n9803_ & new_n15258_;
  assign new_n15313_ = ~new_n15311_ & ~new_n15312_;
  assign new_n15314_ = ~new_n15310_ & new_n15313_;
  assign new_n15315_ = new_n15309_ & new_n15314_;
  assign new_n15316_ = new_n15304_ & new_n15315_;
  assign new_n15317_ = new_n9807_ & new_n15258_;
  assign new_n15318_ = new_n9809_ & new_n15258_;
  assign new_n15319_ = new_n9811_ & new_n15258_;
  assign new_n15320_ = ~new_n15318_ & ~new_n15319_;
  assign new_n15321_ = ~new_n15317_ & new_n15320_;
  assign new_n15322_ = ~A201 & new_n7045_;
  assign new_n15323_ = new_n4255_ & new_n15322_;
  assign new_n15324_ = new_n9817_ & new_n15323_;
  assign new_n15325_ = new_n9819_ & new_n15323_;
  assign new_n15326_ = new_n9821_ & new_n15323_;
  assign new_n15327_ = ~new_n15325_ & ~new_n15326_;
  assign new_n15328_ = ~new_n15324_ & new_n15327_;
  assign new_n15329_ = new_n15321_ & new_n15328_;
  assign new_n15330_ = new_n9842_ & new_n15323_;
  assign new_n15331_ = new_n9825_ & new_n15323_;
  assign new_n15332_ = new_n9828_ & new_n15323_;
  assign new_n15333_ = ~new_n15331_ & ~new_n15332_;
  assign new_n15334_ = ~new_n15330_ & new_n15333_;
  assign new_n15335_ = new_n9844_ & new_n15323_;
  assign new_n15336_ = new_n9840_ & new_n15323_;
  assign new_n15337_ = ~new_n15335_ & ~new_n15336_;
  assign new_n15338_ = new_n15334_ & new_n15337_;
  assign new_n15339_ = new_n15329_ & new_n15338_;
  assign new_n15340_ = new_n15316_ & new_n15339_;
  assign new_n15341_ = new_n9848_ & new_n15323_;
  assign new_n15342_ = new_n9850_ & new_n15323_;
  assign new_n15343_ = new_n9852_ & new_n15323_;
  assign new_n15344_ = ~new_n15342_ & ~new_n15343_;
  assign new_n15345_ = ~new_n15341_ & new_n15344_;
  assign new_n15346_ = new_n9858_ & new_n15323_;
  assign new_n15347_ = new_n9860_ & new_n15323_;
  assign new_n15348_ = new_n9862_ & new_n15323_;
  assign new_n15349_ = ~new_n15347_ & ~new_n15348_;
  assign new_n15350_ = ~new_n15346_ & new_n15349_;
  assign new_n15351_ = new_n15345_ & new_n15350_;
  assign new_n15352_ = new_n9866_ & new_n15323_;
  assign new_n15353_ = new_n9868_ & new_n15323_;
  assign new_n15354_ = new_n9870_ & new_n15323_;
  assign new_n15355_ = ~new_n15353_ & ~new_n15354_;
  assign new_n15356_ = ~new_n15352_ & new_n15355_;
  assign new_n15357_ = new_n9876_ & new_n15323_;
  assign new_n15358_ = new_n9878_ & new_n15323_;
  assign new_n15359_ = new_n9880_ & new_n15323_;
  assign new_n15360_ = ~new_n15358_ & ~new_n15359_;
  assign new_n15361_ = ~new_n15357_ & new_n15360_;
  assign new_n15362_ = new_n15356_ & new_n15361_;
  assign new_n15363_ = new_n15351_ & new_n15362_;
  assign new_n15364_ = new_n9885_ & new_n15323_;
  assign new_n15365_ = new_n9887_ & new_n15323_;
  assign new_n15366_ = new_n9889_ & new_n15323_;
  assign new_n15367_ = ~new_n15365_ & ~new_n15366_;
  assign new_n15368_ = ~new_n15364_ & new_n15367_;
  assign new_n15369_ = new_n9895_ & new_n15323_;
  assign new_n15370_ = new_n9897_ & new_n15323_;
  assign new_n15371_ = new_n9899_ & new_n15323_;
  assign new_n15372_ = ~new_n15370_ & ~new_n15371_;
  assign new_n15373_ = ~new_n15369_ & new_n15372_;
  assign new_n15374_ = new_n15368_ & new_n15373_;
  assign new_n15375_ = new_n9904_ & new_n15323_;
  assign new_n15376_ = new_n9906_ & new_n15323_;
  assign new_n15377_ = new_n9908_ & new_n15323_;
  assign new_n15378_ = ~new_n15376_ & ~new_n15377_;
  assign new_n15379_ = ~new_n15375_ & new_n15378_;
  assign new_n15380_ = new_n9917_ & new_n15323_;
  assign new_n15381_ = new_n9919_ & new_n15323_;
  assign new_n15382_ = ~new_n15380_ & ~new_n15381_;
  assign new_n15383_ = new_n15379_ & new_n15382_;
  assign new_n15384_ = new_n15374_ & new_n15383_;
  assign new_n15385_ = new_n15363_ & new_n15384_;
  assign new_n15386_ = new_n15340_ & new_n15385_;
  assign new_n15387_ = new_n15293_ & new_n15386_;
  assign new_n15388_ = new_n15200_ & new_n15387_;
  assign new_n15389_ = new_n15011_ & new_n15388_;
  assign new_n15390_ = ~A201 & new_n10368_;
  assign new_n15391_ = new_n4255_ & new_n15390_;
  assign new_n15392_ = new_n9928_ & new_n15391_;
  assign new_n15393_ = new_n9915_ & new_n15323_;
  assign new_n15394_ = new_n9926_ & new_n15391_;
  assign new_n15395_ = ~new_n15393_ & ~new_n15394_;
  assign new_n15396_ = ~new_n15392_ & new_n15395_;
  assign new_n15397_ = new_n9938_ & new_n15391_;
  assign new_n15398_ = new_n9924_ & new_n15391_;
  assign new_n15399_ = new_n9936_ & new_n15391_;
  assign new_n15400_ = ~new_n15398_ & ~new_n15399_;
  assign new_n15401_ = ~new_n15397_ & new_n15400_;
  assign new_n15402_ = new_n15396_ & new_n15401_;
  assign new_n15403_ = new_n9946_ & new_n15391_;
  assign new_n15404_ = new_n9934_ & new_n15391_;
  assign new_n15405_ = new_n9944_ & new_n15391_;
  assign new_n15406_ = ~new_n15404_ & ~new_n15405_;
  assign new_n15407_ = ~new_n15403_ & new_n15406_;
  assign new_n15408_ = new_n9956_ & new_n15391_;
  assign new_n15409_ = new_n9942_ & new_n15391_;
  assign new_n15410_ = new_n9954_ & new_n15391_;
  assign new_n15411_ = ~new_n15409_ & ~new_n15410_;
  assign new_n15412_ = ~new_n15408_ & new_n15411_;
  assign new_n15413_ = new_n15407_ & new_n15412_;
  assign new_n15414_ = new_n15402_ & new_n15413_;
  assign new_n15415_ = new_n9965_ & new_n15391_;
  assign new_n15416_ = new_n9952_ & new_n15391_;
  assign new_n15417_ = new_n9963_ & new_n15391_;
  assign new_n15418_ = ~new_n15416_ & ~new_n15417_;
  assign new_n15419_ = ~new_n15415_ & new_n15418_;
  assign new_n15420_ = new_n9974_ & new_n15391_;
  assign new_n15421_ = new_n9961_ & new_n15391_;
  assign new_n15422_ = new_n9972_ & new_n15391_;
  assign new_n15423_ = ~new_n15421_ & ~new_n15422_;
  assign new_n15424_ = ~new_n15420_ & new_n15423_;
  assign new_n15425_ = new_n15419_ & new_n15424_;
  assign new_n15426_ = new_n9980_ & new_n15391_;
  assign new_n15427_ = new_n9970_ & new_n15391_;
  assign new_n15428_ = new_n9978_ & new_n15391_;
  assign new_n15429_ = ~new_n15427_ & ~new_n15428_;
  assign new_n15430_ = ~new_n15426_ & new_n15429_;
  assign new_n15431_ = new_n9988_ & new_n15391_;
  assign new_n15432_ = new_n9990_ & new_n15391_;
  assign new_n15433_ = new_n9992_ & new_n15391_;
  assign new_n15434_ = ~new_n15432_ & ~new_n15433_;
  assign new_n15435_ = ~new_n15431_ & new_n15434_;
  assign new_n15436_ = new_n15430_ & new_n15435_;
  assign new_n15437_ = new_n15425_ & new_n15436_;
  assign new_n15438_ = new_n15414_ & new_n15437_;
  assign new_n15439_ = new_n9997_ & new_n15391_;
  assign new_n15440_ = new_n9999_ & new_n15391_;
  assign new_n15441_ = new_n10001_ & new_n15391_;
  assign new_n15442_ = ~new_n15440_ & ~new_n15441_;
  assign new_n15443_ = ~new_n15439_ & new_n15442_;
  assign new_n15444_ = new_n10007_ & new_n15391_;
  assign new_n15445_ = new_n10009_ & new_n15391_;
  assign new_n15446_ = new_n10011_ & new_n15391_;
  assign new_n15447_ = ~new_n15445_ & ~new_n15446_;
  assign new_n15448_ = ~new_n15444_ & new_n15447_;
  assign new_n15449_ = new_n15443_ & new_n15448_;
  assign new_n15450_ = new_n10015_ & new_n15391_;
  assign new_n15451_ = new_n10017_ & new_n15391_;
  assign new_n15452_ = new_n10019_ & new_n15391_;
  assign new_n15453_ = ~new_n15451_ & ~new_n15452_;
  assign new_n15454_ = ~new_n15450_ & new_n15453_;
  assign new_n15455_ = new_n10026_ & new_n15391_;
  assign new_n15456_ = new_n10028_ & new_n15391_;
  assign new_n15457_ = new_n10030_ & new_n15391_;
  assign new_n15458_ = ~new_n15456_ & ~new_n15457_;
  assign new_n15459_ = ~new_n15455_ & new_n15458_;
  assign new_n15460_ = new_n15454_ & new_n15459_;
  assign new_n15461_ = new_n15449_ & new_n15460_;
  assign new_n15462_ = new_n10035_ & new_n15391_;
  assign new_n15463_ = new_n10037_ & new_n15391_;
  assign new_n15464_ = new_n10039_ & new_n15391_;
  assign new_n15465_ = ~new_n15463_ & ~new_n15464_;
  assign new_n15466_ = ~new_n15462_ & new_n15465_;
  assign new_n15467_ = new_n10044_ & new_n15391_;
  assign new_n15468_ = new_n10046_ & new_n15391_;
  assign new_n15469_ = new_n10048_ & new_n15391_;
  assign new_n15470_ = ~new_n15468_ & ~new_n15469_;
  assign new_n15471_ = ~new_n15467_ & new_n15470_;
  assign new_n15472_ = new_n15466_ & new_n15471_;
  assign new_n15473_ = new_n10063_ & new_n15391_;
  assign new_n15474_ = new_n10052_ & new_n15391_;
  assign new_n15475_ = new_n10054_ & new_n15391_;
  assign new_n15476_ = ~new_n15474_ & ~new_n15475_;
  assign new_n15477_ = ~new_n15473_ & new_n15476_;
  assign new_n15478_ = new_n10065_ & new_n15391_;
  assign new_n15479_ = new_n10061_ & new_n15391_;
  assign new_n15480_ = ~new_n15478_ & ~new_n15479_;
  assign new_n15481_ = new_n15477_ & new_n15480_;
  assign new_n15482_ = new_n15472_ & new_n15481_;
  assign new_n15483_ = new_n15461_ & new_n15482_;
  assign new_n15484_ = new_n15438_ & new_n15483_;
  assign new_n15485_ = new_n10069_ & new_n15391_;
  assign new_n15486_ = new_n10071_ & new_n15391_;
  assign new_n15487_ = new_n10073_ & new_n15391_;
  assign new_n15488_ = ~new_n15486_ & ~new_n15487_;
  assign new_n15489_ = ~new_n15485_ & new_n15488_;
  assign new_n15490_ = new_n10078_ & new_n15391_;
  assign new_n15491_ = new_n10080_ & new_n15391_;
  assign new_n15492_ = new_n10082_ & new_n15391_;
  assign new_n15493_ = ~new_n15491_ & ~new_n15492_;
  assign new_n15494_ = ~new_n15490_ & new_n15493_;
  assign new_n15495_ = new_n15489_ & new_n15494_;
  assign new_n15496_ = new_n10087_ & new_n15391_;
  assign new_n15497_ = new_n10089_ & new_n15391_;
  assign new_n15498_ = new_n10091_ & new_n15391_;
  assign new_n15499_ = ~new_n15497_ & ~new_n15498_;
  assign new_n15500_ = ~new_n15496_ & new_n15499_;
  assign new_n15501_ = new_n10098_ & new_n15391_;
  assign new_n15502_ = new_n10100_ & new_n15391_;
  assign new_n15503_ = new_n10102_ & new_n15391_;
  assign new_n15504_ = ~new_n15502_ & ~new_n15503_;
  assign new_n15505_ = ~new_n15501_ & new_n15504_;
  assign new_n15506_ = new_n15500_ & new_n15505_;
  assign new_n15507_ = new_n15495_ & new_n15506_;
  assign new_n15508_ = new_n10107_ & new_n15391_;
  assign new_n15509_ = new_n10109_ & new_n15391_;
  assign new_n15510_ = new_n10111_ & new_n15391_;
  assign new_n15511_ = ~new_n15509_ & ~new_n15510_;
  assign new_n15512_ = ~new_n15508_ & new_n15511_;
  assign new_n15513_ = new_n10116_ & new_n15391_;
  assign new_n15514_ = new_n10118_ & new_n15391_;
  assign new_n15515_ = new_n10120_ & new_n15391_;
  assign new_n15516_ = ~new_n15514_ & ~new_n15515_;
  assign new_n15517_ = ~new_n15513_ & new_n15516_;
  assign new_n15518_ = new_n15512_ & new_n15517_;
  assign new_n15519_ = ~A201 & new_n7543_;
  assign new_n15520_ = new_n4255_ & new_n15519_;
  assign new_n15521_ = new_n9716_ & new_n15520_;
  assign new_n15522_ = new_n9718_ & new_n15520_;
  assign new_n15523_ = new_n9720_ & new_n15520_;
  assign new_n15524_ = ~new_n15522_ & ~new_n15523_;
  assign new_n15525_ = ~new_n15521_ & new_n15524_;
  assign new_n15526_ = new_n9729_ & new_n15520_;
  assign new_n15527_ = new_n9731_ & new_n15520_;
  assign new_n15528_ = ~new_n15526_ & ~new_n15527_;
  assign new_n15529_ = new_n15525_ & new_n15528_;
  assign new_n15530_ = new_n15518_ & new_n15529_;
  assign new_n15531_ = new_n15507_ & new_n15530_;
  assign new_n15532_ = new_n9739_ & new_n15520_;
  assign new_n15533_ = new_n9727_ & new_n15520_;
  assign new_n15534_ = new_n9737_ & new_n15520_;
  assign new_n15535_ = ~new_n15533_ & ~new_n15534_;
  assign new_n15536_ = ~new_n15532_ & new_n15535_;
  assign new_n15537_ = new_n9748_ & new_n15520_;
  assign new_n15538_ = new_n9735_ & new_n15520_;
  assign new_n15539_ = new_n9746_ & new_n15520_;
  assign new_n15540_ = ~new_n15538_ & ~new_n15539_;
  assign new_n15541_ = ~new_n15537_ & new_n15540_;
  assign new_n15542_ = new_n15536_ & new_n15541_;
  assign new_n15543_ = new_n9755_ & new_n15520_;
  assign new_n15544_ = new_n9744_ & new_n15520_;
  assign new_n15545_ = new_n9753_ & new_n15520_;
  assign new_n15546_ = ~new_n15544_ & ~new_n15545_;
  assign new_n15547_ = ~new_n15543_ & new_n15546_;
  assign new_n15548_ = new_n9761_ & new_n15520_;
  assign new_n15549_ = new_n9763_ & new_n15520_;
  assign new_n15550_ = new_n9765_ & new_n15520_;
  assign new_n15551_ = ~new_n15549_ & ~new_n15550_;
  assign new_n15552_ = ~new_n15548_ & new_n15551_;
  assign new_n15553_ = new_n15547_ & new_n15552_;
  assign new_n15554_ = new_n15542_ & new_n15553_;
  assign new_n15555_ = new_n9769_ & new_n15520_;
  assign new_n15556_ = new_n9771_ & new_n15520_;
  assign new_n15557_ = new_n9773_ & new_n15520_;
  assign new_n15558_ = ~new_n15556_ & ~new_n15557_;
  assign new_n15559_ = ~new_n15555_ & new_n15558_;
  assign new_n15560_ = new_n9779_ & new_n15520_;
  assign new_n15561_ = new_n9781_ & new_n15520_;
  assign new_n15562_ = new_n9783_ & new_n15520_;
  assign new_n15563_ = ~new_n15561_ & ~new_n15562_;
  assign new_n15564_ = ~new_n15560_ & new_n15563_;
  assign new_n15565_ = new_n15559_ & new_n15564_;
  assign new_n15566_ = new_n9788_ & new_n15520_;
  assign new_n15567_ = new_n9790_ & new_n15520_;
  assign new_n15568_ = new_n9792_ & new_n15520_;
  assign new_n15569_ = ~new_n15567_ & ~new_n15568_;
  assign new_n15570_ = ~new_n15566_ & new_n15569_;
  assign new_n15571_ = new_n9801_ & new_n15520_;
  assign new_n15572_ = new_n9803_ & new_n15520_;
  assign new_n15573_ = ~new_n15571_ & ~new_n15572_;
  assign new_n15574_ = new_n15570_ & new_n15573_;
  assign new_n15575_ = new_n15565_ & new_n15574_;
  assign new_n15576_ = new_n15554_ & new_n15575_;
  assign new_n15577_ = new_n15531_ & new_n15576_;
  assign new_n15578_ = new_n15484_ & new_n15577_;
  assign new_n15579_ = new_n9811_ & new_n15520_;
  assign new_n15580_ = new_n9799_ & new_n15520_;
  assign new_n15581_ = new_n9809_ & new_n15520_;
  assign new_n15582_ = ~new_n15580_ & ~new_n15581_;
  assign new_n15583_ = ~new_n15579_ & new_n15582_;
  assign new_n15584_ = ~A201 & new_n7374_;
  assign new_n15585_ = new_n4255_ & new_n15584_;
  assign new_n15586_ = new_n9821_ & new_n15585_;
  assign new_n15587_ = new_n9807_ & new_n15520_;
  assign new_n15588_ = new_n9819_ & new_n15585_;
  assign new_n15589_ = ~new_n15587_ & ~new_n15588_;
  assign new_n15590_ = ~new_n15586_ & new_n15589_;
  assign new_n15591_ = new_n15583_ & new_n15590_;
  assign new_n15592_ = new_n9828_ & new_n15585_;
  assign new_n15593_ = new_n9817_ & new_n15585_;
  assign new_n15594_ = new_n9825_ & new_n15585_;
  assign new_n15595_ = ~new_n15593_ & ~new_n15594_;
  assign new_n15596_ = ~new_n15592_ & new_n15595_;
  assign new_n15597_ = new_n9840_ & new_n15585_;
  assign new_n15598_ = new_n9842_ & new_n15585_;
  assign new_n15599_ = new_n9844_ & new_n15585_;
  assign new_n15600_ = ~new_n15598_ & ~new_n15599_;
  assign new_n15601_ = ~new_n15597_ & new_n15600_;
  assign new_n15602_ = new_n15596_ & new_n15601_;
  assign new_n15603_ = new_n15591_ & new_n15602_;
  assign new_n15604_ = new_n9848_ & new_n15585_;
  assign new_n15605_ = new_n9850_ & new_n15585_;
  assign new_n15606_ = new_n9852_ & new_n15585_;
  assign new_n15607_ = ~new_n15605_ & ~new_n15606_;
  assign new_n15608_ = ~new_n15604_ & new_n15607_;
  assign new_n15609_ = new_n9858_ & new_n15585_;
  assign new_n15610_ = new_n9860_ & new_n15585_;
  assign new_n15611_ = new_n9862_ & new_n15585_;
  assign new_n15612_ = ~new_n15610_ & ~new_n15611_;
  assign new_n15613_ = ~new_n15609_ & new_n15612_;
  assign new_n15614_ = new_n15608_ & new_n15613_;
  assign new_n15615_ = new_n9866_ & new_n15585_;
  assign new_n15616_ = new_n9868_ & new_n15585_;
  assign new_n15617_ = new_n9870_ & new_n15585_;
  assign new_n15618_ = ~new_n15616_ & ~new_n15617_;
  assign new_n15619_ = ~new_n15615_ & new_n15618_;
  assign new_n15620_ = new_n9878_ & new_n15585_;
  assign new_n15621_ = new_n9880_ & new_n15585_;
  assign new_n15622_ = ~new_n15620_ & ~new_n15621_;
  assign new_n15623_ = new_n15619_ & new_n15622_;
  assign new_n15624_ = new_n15614_ & new_n15623_;
  assign new_n15625_ = new_n15603_ & new_n15624_;
  assign new_n15626_ = new_n9889_ & new_n15585_;
  assign new_n15627_ = new_n9876_ & new_n15585_;
  assign new_n15628_ = new_n9887_ & new_n15585_;
  assign new_n15629_ = ~new_n15627_ & ~new_n15628_;
  assign new_n15630_ = ~new_n15626_ & new_n15629_;
  assign new_n15631_ = new_n9899_ & new_n15585_;
  assign new_n15632_ = new_n9885_ & new_n15585_;
  assign new_n15633_ = new_n9897_ & new_n15585_;
  assign new_n15634_ = ~new_n15632_ & ~new_n15633_;
  assign new_n15635_ = ~new_n15631_ & new_n15634_;
  assign new_n15636_ = new_n15630_ & new_n15635_;
  assign new_n15637_ = new_n9908_ & new_n15585_;
  assign new_n15638_ = new_n9895_ & new_n15585_;
  assign new_n15639_ = new_n9906_ & new_n15585_;
  assign new_n15640_ = ~new_n15638_ & ~new_n15639_;
  assign new_n15641_ = ~new_n15637_ & new_n15640_;
  assign new_n15642_ = new_n9919_ & new_n15585_;
  assign new_n15643_ = new_n9904_ & new_n15585_;
  assign new_n15644_ = new_n9917_ & new_n15585_;
  assign new_n15645_ = ~new_n15643_ & ~new_n15644_;
  assign new_n15646_ = ~new_n15642_ & new_n15645_;
  assign new_n15647_ = new_n15641_ & new_n15646_;
  assign new_n15648_ = new_n15636_ & new_n15647_;
  assign new_n15649_ = ~A201 & new_n10478_;
  assign new_n15650_ = new_n4255_ & new_n15649_;
  assign new_n15651_ = new_n9928_ & new_n15650_;
  assign new_n15652_ = new_n9915_ & new_n15585_;
  assign new_n15653_ = new_n9926_ & new_n15650_;
  assign new_n15654_ = ~new_n15652_ & ~new_n15653_;
  assign new_n15655_ = ~new_n15651_ & new_n15654_;
  assign new_n15656_ = new_n9938_ & new_n15650_;
  assign new_n15657_ = new_n9924_ & new_n15650_;
  assign new_n15658_ = new_n9936_ & new_n15650_;
  assign new_n15659_ = ~new_n15657_ & ~new_n15658_;
  assign new_n15660_ = ~new_n15656_ & new_n15659_;
  assign new_n15661_ = new_n15655_ & new_n15660_;
  assign new_n15662_ = new_n9946_ & new_n15650_;
  assign new_n15663_ = new_n9934_ & new_n15650_;
  assign new_n15664_ = new_n9944_ & new_n15650_;
  assign new_n15665_ = ~new_n15663_ & ~new_n15664_;
  assign new_n15666_ = ~new_n15662_ & new_n15665_;
  assign new_n15667_ = new_n9942_ & new_n15650_;
  assign new_n15668_ = new_n9954_ & new_n15650_;
  assign new_n15669_ = ~new_n15667_ & ~new_n15668_;
  assign new_n15670_ = new_n15666_ & new_n15669_;
  assign new_n15671_ = new_n15661_ & new_n15670_;
  assign new_n15672_ = new_n15648_ & new_n15671_;
  assign new_n15673_ = new_n15625_ & new_n15672_;
  assign new_n15674_ = new_n9963_ & new_n15650_;
  assign new_n15675_ = new_n9956_ & new_n15650_;
  assign new_n15676_ = new_n9952_ & new_n15650_;
  assign new_n15677_ = ~new_n15675_ & ~new_n15676_;
  assign new_n15678_ = ~new_n15674_ & new_n15677_;
  assign new_n15679_ = new_n9972_ & new_n15650_;
  assign new_n15680_ = new_n9965_ & new_n15650_;
  assign new_n15681_ = new_n9961_ & new_n15650_;
  assign new_n15682_ = ~new_n15680_ & ~new_n15681_;
  assign new_n15683_ = ~new_n15679_ & new_n15682_;
  assign new_n15684_ = new_n15678_ & new_n15683_;
  assign new_n15685_ = new_n9978_ & new_n15650_;
  assign new_n15686_ = new_n9974_ & new_n15650_;
  assign new_n15687_ = new_n9970_ & new_n15650_;
  assign new_n15688_ = ~new_n15686_ & ~new_n15687_;
  assign new_n15689_ = ~new_n15685_ & new_n15688_;
  assign new_n15690_ = new_n9992_ & new_n15650_;
  assign new_n15691_ = new_n9980_ & new_n15650_;
  assign new_n15692_ = new_n9990_ & new_n15650_;
  assign new_n15693_ = ~new_n15691_ & ~new_n15692_;
  assign new_n15694_ = ~new_n15690_ & new_n15693_;
  assign new_n15695_ = new_n15689_ & new_n15694_;
  assign new_n15696_ = new_n15684_ & new_n15695_;
  assign new_n15697_ = new_n10001_ & new_n15650_;
  assign new_n15698_ = new_n9988_ & new_n15650_;
  assign new_n15699_ = new_n9999_ & new_n15650_;
  assign new_n15700_ = ~new_n15698_ & ~new_n15699_;
  assign new_n15701_ = ~new_n15697_ & new_n15700_;
  assign new_n15702_ = new_n10011_ & new_n15650_;
  assign new_n15703_ = new_n9997_ & new_n15650_;
  assign new_n15704_ = new_n10009_ & new_n15650_;
  assign new_n15705_ = ~new_n15703_ & ~new_n15704_;
  assign new_n15706_ = ~new_n15702_ & new_n15705_;
  assign new_n15707_ = new_n15701_ & new_n15706_;
  assign new_n15708_ = new_n10019_ & new_n15650_;
  assign new_n15709_ = new_n10007_ & new_n15650_;
  assign new_n15710_ = new_n10017_ & new_n15650_;
  assign new_n15711_ = ~new_n15709_ & ~new_n15710_;
  assign new_n15712_ = ~new_n15708_ & new_n15711_;
  assign new_n15713_ = new_n10015_ & new_n15650_;
  assign new_n15714_ = new_n10028_ & new_n15650_;
  assign new_n15715_ = ~new_n15713_ & ~new_n15714_;
  assign new_n15716_ = new_n15712_ & new_n15715_;
  assign new_n15717_ = new_n15707_ & new_n15716_;
  assign new_n15718_ = new_n15696_ & new_n15717_;
  assign new_n15719_ = new_n10037_ & new_n15650_;
  assign new_n15720_ = new_n10030_ & new_n15650_;
  assign new_n15721_ = new_n10026_ & new_n15650_;
  assign new_n15722_ = ~new_n15720_ & ~new_n15721_;
  assign new_n15723_ = ~new_n15719_ & new_n15722_;
  assign new_n15724_ = new_n10046_ & new_n15650_;
  assign new_n15725_ = new_n10039_ & new_n15650_;
  assign new_n15726_ = new_n10035_ & new_n15650_;
  assign new_n15727_ = ~new_n15725_ & ~new_n15726_;
  assign new_n15728_ = ~new_n15724_ & new_n15727_;
  assign new_n15729_ = new_n15723_ & new_n15728_;
  assign new_n15730_ = new_n10052_ & new_n15650_;
  assign new_n15731_ = new_n10048_ & new_n15650_;
  assign new_n15732_ = new_n10044_ & new_n15650_;
  assign new_n15733_ = ~new_n15731_ & ~new_n15732_;
  assign new_n15734_ = ~new_n15730_ & new_n15733_;
  assign new_n15735_ = new_n10065_ & new_n15650_;
  assign new_n15736_ = new_n10054_ & new_n15650_;
  assign new_n15737_ = new_n10063_ & new_n15650_;
  assign new_n15738_ = ~new_n15736_ & ~new_n15737_;
  assign new_n15739_ = ~new_n15735_ & new_n15738_;
  assign new_n15740_ = new_n15734_ & new_n15739_;
  assign new_n15741_ = new_n15729_ & new_n15740_;
  assign new_n15742_ = new_n10073_ & new_n15650_;
  assign new_n15743_ = new_n10061_ & new_n15650_;
  assign new_n15744_ = new_n10071_ & new_n15650_;
  assign new_n15745_ = ~new_n15743_ & ~new_n15744_;
  assign new_n15746_ = ~new_n15742_ & new_n15745_;
  assign new_n15747_ = new_n10082_ & new_n15650_;
  assign new_n15748_ = new_n10069_ & new_n15650_;
  assign new_n15749_ = new_n10080_ & new_n15650_;
  assign new_n15750_ = ~new_n15748_ & ~new_n15749_;
  assign new_n15751_ = ~new_n15747_ & new_n15750_;
  assign new_n15752_ = new_n15746_ & new_n15751_;
  assign new_n15753_ = new_n10091_ & new_n15650_;
  assign new_n15754_ = new_n10078_ & new_n15650_;
  assign new_n15755_ = new_n10089_ & new_n15650_;
  assign new_n15756_ = ~new_n15754_ & ~new_n15755_;
  assign new_n15757_ = ~new_n15753_ & new_n15756_;
  assign new_n15758_ = new_n10087_ & new_n15650_;
  assign new_n15759_ = new_n10100_ & new_n15650_;
  assign new_n15760_ = ~new_n15758_ & ~new_n15759_;
  assign new_n15761_ = new_n15757_ & new_n15760_;
  assign new_n15762_ = new_n15752_ & new_n15761_;
  assign new_n15763_ = new_n15741_ & new_n15762_;
  assign new_n15764_ = new_n15718_ & new_n15763_;
  assign new_n15765_ = new_n15673_ & new_n15764_;
  assign new_n15766_ = new_n15578_ & new_n15765_;
  assign new_n15767_ = new_n10109_ & new_n15650_;
  assign new_n15768_ = new_n10102_ & new_n15650_;
  assign new_n15769_ = new_n10098_ & new_n15650_;
  assign new_n15770_ = ~new_n15768_ & ~new_n15769_;
  assign new_n15771_ = ~new_n15767_ & new_n15770_;
  assign new_n15772_ = new_n10118_ & new_n15650_;
  assign new_n15773_ = new_n10111_ & new_n15650_;
  assign new_n15774_ = new_n10107_ & new_n15650_;
  assign new_n15775_ = ~new_n15773_ & ~new_n15774_;
  assign new_n15776_ = ~new_n15772_ & new_n15775_;
  assign new_n15777_ = new_n15771_ & new_n15776_;
  assign new_n15778_ = ~A200 & new_n1781_;
  assign new_n15779_ = new_n4968_ & new_n15778_;
  assign new_n15780_ = new_n8617_ & new_n15779_;
  assign new_n15781_ = new_n10120_ & new_n15650_;
  assign new_n15782_ = new_n10116_ & new_n15650_;
  assign new_n15783_ = ~new_n15781_ & ~new_n15782_;
  assign new_n15784_ = ~new_n15780_ & new_n15783_;
  assign new_n15785_ = new_n8625_ & new_n15779_;
  assign new_n15786_ = new_n8628_ & new_n15779_;
  assign new_n15787_ = new_n8630_ & new_n15779_;
  assign new_n15788_ = ~new_n15786_ & ~new_n15787_;
  assign new_n15789_ = ~new_n15785_ & new_n15788_;
  assign new_n15790_ = new_n15784_ & new_n15789_;
  assign new_n15791_ = new_n15777_ & new_n15790_;
  assign new_n15792_ = new_n8635_ & new_n15779_;
  assign new_n15793_ = new_n8637_ & new_n15779_;
  assign new_n15794_ = new_n8639_ & new_n15779_;
  assign new_n15795_ = ~new_n15793_ & ~new_n15794_;
  assign new_n15796_ = ~new_n15792_ & new_n15795_;
  assign new_n15797_ = new_n8646_ & new_n15779_;
  assign new_n15798_ = new_n8648_ & new_n15779_;
  assign new_n15799_ = new_n8650_ & new_n15779_;
  assign new_n15800_ = ~new_n15798_ & ~new_n15799_;
  assign new_n15801_ = ~new_n15797_ & new_n15800_;
  assign new_n15802_ = new_n15796_ & new_n15801_;
  assign new_n15803_ = new_n8655_ & new_n15779_;
  assign new_n15804_ = new_n8657_ & new_n15779_;
  assign new_n15805_ = new_n8659_ & new_n15779_;
  assign new_n15806_ = ~new_n15804_ & ~new_n15805_;
  assign new_n15807_ = ~new_n15803_ & new_n15806_;
  assign new_n15808_ = new_n8667_ & new_n15779_;
  assign new_n15809_ = new_n8670_ & new_n15779_;
  assign new_n15810_ = ~new_n15808_ & ~new_n15809_;
  assign new_n15811_ = new_n15807_ & new_n15810_;
  assign new_n15812_ = new_n15802_ & new_n15811_;
  assign new_n15813_ = new_n15791_ & new_n15812_;
  assign new_n15814_ = new_n8681_ & new_n15779_;
  assign new_n15815_ = new_n8665_ & new_n15779_;
  assign new_n15816_ = new_n8678_ & new_n15779_;
  assign new_n15817_ = ~new_n15815_ & ~new_n15816_;
  assign new_n15818_ = ~new_n15814_ & new_n15817_;
  assign new_n15819_ = new_n8694_ & new_n15779_;
  assign new_n15820_ = new_n8675_ & new_n15779_;
  assign new_n15821_ = new_n8692_ & new_n15779_;
  assign new_n15822_ = ~new_n15820_ & ~new_n15821_;
  assign new_n15823_ = ~new_n15819_ & new_n15822_;
  assign new_n15824_ = new_n15818_ & new_n15823_;
  assign new_n15825_ = new_n8701_ & new_n15779_;
  assign new_n15826_ = new_n8689_ & new_n15779_;
  assign new_n15827_ = new_n8699_ & new_n15779_;
  assign new_n15828_ = ~new_n15826_ & ~new_n15827_;
  assign new_n15829_ = ~new_n15825_ & new_n15828_;
  assign new_n15830_ = ~A200 & new_n1795_;
  assign new_n15831_ = new_n4968_ & new_n15830_;
  assign new_n15832_ = new_n8630_ & new_n15831_;
  assign new_n15833_ = new_n8617_ & new_n15831_;
  assign new_n15834_ = new_n8628_ & new_n15831_;
  assign new_n15835_ = ~new_n15833_ & ~new_n15834_;
  assign new_n15836_ = ~new_n15832_ & new_n15835_;
  assign new_n15837_ = new_n15829_ & new_n15836_;
  assign new_n15838_ = new_n15824_ & new_n15837_;
  assign new_n15839_ = new_n8639_ & new_n15831_;
  assign new_n15840_ = new_n8625_ & new_n15831_;
  assign new_n15841_ = new_n8637_ & new_n15831_;
  assign new_n15842_ = ~new_n15840_ & ~new_n15841_;
  assign new_n15843_ = ~new_n15839_ & new_n15842_;
  assign new_n15844_ = new_n8650_ & new_n15831_;
  assign new_n15845_ = new_n8635_ & new_n15831_;
  assign new_n15846_ = new_n8648_ & new_n15831_;
  assign new_n15847_ = ~new_n15845_ & ~new_n15846_;
  assign new_n15848_ = ~new_n15844_ & new_n15847_;
  assign new_n15849_ = new_n15843_ & new_n15848_;
  assign new_n15850_ = new_n8659_ & new_n15831_;
  assign new_n15851_ = new_n8646_ & new_n15831_;
  assign new_n15852_ = new_n8657_ & new_n15831_;
  assign new_n15853_ = ~new_n15851_ & ~new_n15852_;
  assign new_n15854_ = ~new_n15850_ & new_n15853_;
  assign new_n15855_ = new_n8655_ & new_n15831_;
  assign new_n15856_ = new_n8667_ & new_n15831_;
  assign new_n15857_ = ~new_n15855_ & ~new_n15856_;
  assign new_n15858_ = new_n15854_ & new_n15857_;
  assign new_n15859_ = new_n15849_ & new_n15858_;
  assign new_n15860_ = new_n15838_ & new_n15859_;
  assign new_n15861_ = new_n15813_ & new_n15860_;
  assign new_n15862_ = new_n8678_ & new_n15831_;
  assign new_n15863_ = new_n8670_ & new_n15831_;
  assign new_n15864_ = new_n8665_ & new_n15831_;
  assign new_n15865_ = ~new_n15863_ & ~new_n15864_;
  assign new_n15866_ = ~new_n15862_ & new_n15865_;
  assign new_n15867_ = new_n8692_ & new_n15831_;
  assign new_n15868_ = new_n8681_ & new_n15831_;
  assign new_n15869_ = new_n8675_ & new_n15831_;
  assign new_n15870_ = ~new_n15868_ & ~new_n15869_;
  assign new_n15871_ = ~new_n15867_ & new_n15870_;
  assign new_n15872_ = new_n15866_ & new_n15871_;
  assign new_n15873_ = new_n8699_ & new_n15831_;
  assign new_n15874_ = new_n8694_ & new_n15831_;
  assign new_n15875_ = new_n8689_ & new_n15831_;
  assign new_n15876_ = ~new_n15874_ & ~new_n15875_;
  assign new_n15877_ = ~new_n15873_ & new_n15876_;
  assign new_n15878_ = ~A200 & new_n1804_;
  assign new_n15879_ = new_n4968_ & new_n15878_;
  assign new_n15880_ = new_n8628_ & new_n15879_;
  assign new_n15881_ = new_n8701_ & new_n15831_;
  assign new_n15882_ = new_n8617_ & new_n15879_;
  assign new_n15883_ = ~new_n15881_ & ~new_n15882_;
  assign new_n15884_ = ~new_n15880_ & new_n15883_;
  assign new_n15885_ = new_n15877_ & new_n15884_;
  assign new_n15886_ = new_n15872_ & new_n15885_;
  assign new_n15887_ = new_n8637_ & new_n15879_;
  assign new_n15888_ = new_n8630_ & new_n15879_;
  assign new_n15889_ = new_n8625_ & new_n15879_;
  assign new_n15890_ = ~new_n15888_ & ~new_n15889_;
  assign new_n15891_ = ~new_n15887_ & new_n15890_;
  assign new_n15892_ = new_n8648_ & new_n15879_;
  assign new_n15893_ = new_n8639_ & new_n15879_;
  assign new_n15894_ = new_n8635_ & new_n15879_;
  assign new_n15895_ = ~new_n15893_ & ~new_n15894_;
  assign new_n15896_ = ~new_n15892_ & new_n15895_;
  assign new_n15897_ = new_n15891_ & new_n15896_;
  assign new_n15898_ = new_n8657_ & new_n15879_;
  assign new_n15899_ = new_n8650_ & new_n15879_;
  assign new_n15900_ = new_n8646_ & new_n15879_;
  assign new_n15901_ = ~new_n15899_ & ~new_n15900_;
  assign new_n15902_ = ~new_n15898_ & new_n15901_;
  assign new_n15903_ = new_n8659_ & new_n15879_;
  assign new_n15904_ = new_n8655_ & new_n15879_;
  assign new_n15905_ = ~new_n15903_ & ~new_n15904_;
  assign new_n15906_ = new_n15902_ & new_n15905_;
  assign new_n15907_ = new_n15897_ & new_n15906_;
  assign new_n15908_ = new_n15886_ & new_n15907_;
  assign new_n15909_ = new_n8665_ & new_n15879_;
  assign new_n15910_ = new_n8667_ & new_n15879_;
  assign new_n15911_ = new_n8670_ & new_n15879_;
  assign new_n15912_ = ~new_n15910_ & ~new_n15911_;
  assign new_n15913_ = ~new_n15909_ & new_n15912_;
  assign new_n15914_ = new_n8675_ & new_n15879_;
  assign new_n15915_ = new_n8678_ & new_n15879_;
  assign new_n15916_ = new_n8681_ & new_n15879_;
  assign new_n15917_ = ~new_n15915_ & ~new_n15916_;
  assign new_n15918_ = ~new_n15914_ & new_n15917_;
  assign new_n15919_ = new_n15913_ & new_n15918_;
  assign new_n15920_ = new_n8689_ & new_n15879_;
  assign new_n15921_ = new_n8692_ & new_n15879_;
  assign new_n15922_ = new_n8694_ & new_n15879_;
  assign new_n15923_ = ~new_n15921_ & ~new_n15922_;
  assign new_n15924_ = ~new_n15920_ & new_n15923_;
  assign new_n15925_ = ~A200 & new_n1812_;
  assign new_n15926_ = new_n4968_ & new_n15925_;
  assign new_n15927_ = new_n8617_ & new_n15926_;
  assign new_n15928_ = new_n8699_ & new_n15879_;
  assign new_n15929_ = new_n8701_ & new_n15879_;
  assign new_n15930_ = ~new_n15928_ & ~new_n15929_;
  assign new_n15931_ = ~new_n15927_ & new_n15930_;
  assign new_n15932_ = new_n15924_ & new_n15931_;
  assign new_n15933_ = new_n15919_ & new_n15932_;
  assign new_n15934_ = new_n8625_ & new_n15926_;
  assign new_n15935_ = new_n8628_ & new_n15926_;
  assign new_n15936_ = new_n8630_ & new_n15926_;
  assign new_n15937_ = ~new_n15935_ & ~new_n15936_;
  assign new_n15938_ = ~new_n15934_ & new_n15937_;
  assign new_n15939_ = new_n8635_ & new_n15926_;
  assign new_n15940_ = new_n8637_ & new_n15926_;
  assign new_n15941_ = new_n8639_ & new_n15926_;
  assign new_n15942_ = ~new_n15940_ & ~new_n15941_;
  assign new_n15943_ = ~new_n15939_ & new_n15942_;
  assign new_n15944_ = new_n15938_ & new_n15943_;
  assign new_n15945_ = new_n8646_ & new_n15926_;
  assign new_n15946_ = new_n8648_ & new_n15926_;
  assign new_n15947_ = new_n8650_ & new_n15926_;
  assign new_n15948_ = ~new_n15946_ & ~new_n15947_;
  assign new_n15949_ = ~new_n15945_ & new_n15948_;
  assign new_n15950_ = new_n8657_ & new_n15926_;
  assign new_n15951_ = new_n8659_ & new_n15926_;
  assign new_n15952_ = ~new_n15950_ & ~new_n15951_;
  assign new_n15953_ = new_n15949_ & new_n15952_;
  assign new_n15954_ = new_n15944_ & new_n15953_;
  assign new_n15955_ = new_n15933_ & new_n15954_;
  assign new_n15956_ = new_n15908_ & new_n15955_;
  assign new_n15957_ = new_n15861_ & new_n15956_;
  assign new_n15958_ = new_n8670_ & new_n15926_;
  assign new_n15959_ = new_n8655_ & new_n15926_;
  assign new_n15960_ = new_n8667_ & new_n15926_;
  assign new_n15961_ = ~new_n15959_ & ~new_n15960_;
  assign new_n15962_ = ~new_n15958_ & new_n15961_;
  assign new_n15963_ = new_n8681_ & new_n15926_;
  assign new_n15964_ = new_n8665_ & new_n15926_;
  assign new_n15965_ = new_n8678_ & new_n15926_;
  assign new_n15966_ = ~new_n15964_ & ~new_n15965_;
  assign new_n15967_ = ~new_n15963_ & new_n15966_;
  assign new_n15968_ = new_n15962_ & new_n15967_;
  assign new_n15969_ = new_n8694_ & new_n15926_;
  assign new_n15970_ = new_n8675_ & new_n15926_;
  assign new_n15971_ = new_n8692_ & new_n15926_;
  assign new_n15972_ = ~new_n15970_ & ~new_n15971_;
  assign new_n15973_ = ~new_n15969_ & new_n15972_;
  assign new_n15974_ = new_n8701_ & new_n15926_;
  assign new_n15975_ = new_n8689_ & new_n15926_;
  assign new_n15976_ = new_n8699_ & new_n15926_;
  assign new_n15977_ = ~new_n15975_ & ~new_n15976_;
  assign new_n15978_ = ~new_n15974_ & new_n15977_;
  assign new_n15979_ = new_n15973_ & new_n15978_;
  assign new_n15980_ = new_n15968_ & new_n15979_;
  assign new_n15981_ = ~A200 & new_n504_;
  assign new_n15982_ = new_n4968_ & new_n15981_;
  assign new_n15983_ = new_n8855_ & new_n15982_;
  assign new_n15984_ = new_n8845_ & new_n15982_;
  assign new_n15985_ = new_n8853_ & new_n15982_;
  assign new_n15986_ = ~new_n15984_ & ~new_n15985_;
  assign new_n15987_ = ~new_n15983_ & new_n15986_;
  assign new_n15988_ = new_n8866_ & new_n15982_;
  assign new_n15989_ = new_n8851_ & new_n15982_;
  assign new_n15990_ = new_n8864_ & new_n15982_;
  assign new_n15991_ = ~new_n15989_ & ~new_n15990_;
  assign new_n15992_ = ~new_n15988_ & new_n15991_;
  assign new_n15993_ = new_n15987_ & new_n15992_;
  assign new_n15994_ = new_n8874_ & new_n15982_;
  assign new_n15995_ = new_n8862_ & new_n15982_;
  assign new_n15996_ = new_n8872_ & new_n15982_;
  assign new_n15997_ = ~new_n15995_ & ~new_n15996_;
  assign new_n15998_ = ~new_n15994_ & new_n15997_;
  assign new_n15999_ = new_n8870_ & new_n15982_;
  assign new_n16000_ = new_n8882_ & new_n15982_;
  assign new_n16001_ = ~new_n15999_ & ~new_n16000_;
  assign new_n16002_ = new_n15998_ & new_n16001_;
  assign new_n16003_ = new_n15993_ & new_n16002_;
  assign new_n16004_ = new_n15980_ & new_n16003_;
  assign new_n16005_ = new_n8888_ & new_n15982_;
  assign new_n16006_ = new_n8884_ & new_n15982_;
  assign new_n16007_ = new_n8880_ & new_n15982_;
  assign new_n16008_ = ~new_n16006_ & ~new_n16007_;
  assign new_n16009_ = ~new_n16005_ & new_n16008_;
  assign new_n16010_ = new_n8900_ & new_n15982_;
  assign new_n16011_ = new_n8890_ & new_n15982_;
  assign new_n16012_ = new_n8898_ & new_n15982_;
  assign new_n16013_ = ~new_n16011_ & ~new_n16012_;
  assign new_n16014_ = ~new_n16010_ & new_n16013_;
  assign new_n16015_ = new_n16009_ & new_n16014_;
  assign new_n16016_ = new_n8909_ & new_n15982_;
  assign new_n16017_ = new_n8896_ & new_n15982_;
  assign new_n16018_ = new_n8907_ & new_n15982_;
  assign new_n16019_ = ~new_n16017_ & ~new_n16018_;
  assign new_n16020_ = ~new_n16016_ & new_n16019_;
  assign new_n16021_ = new_n8918_ & new_n15982_;
  assign new_n16022_ = new_n8905_ & new_n15982_;
  assign new_n16023_ = new_n8916_ & new_n15982_;
  assign new_n16024_ = ~new_n16022_ & ~new_n16023_;
  assign new_n16025_ = ~new_n16021_ & new_n16024_;
  assign new_n16026_ = new_n16020_ & new_n16025_;
  assign new_n16027_ = new_n16015_ & new_n16026_;
  assign new_n16028_ = new_n8927_ & new_n15982_;
  assign new_n16029_ = new_n8914_ & new_n15982_;
  assign new_n16030_ = new_n8925_ & new_n15982_;
  assign new_n16031_ = ~new_n16029_ & ~new_n16030_;
  assign new_n16032_ = ~new_n16028_ & new_n16031_;
  assign new_n16033_ = new_n8938_ & new_n15982_;
  assign new_n16034_ = new_n8923_ & new_n15982_;
  assign new_n16035_ = new_n8936_ & new_n15982_;
  assign new_n16036_ = ~new_n16034_ & ~new_n16035_;
  assign new_n16037_ = ~new_n16033_ & new_n16036_;
  assign new_n16038_ = new_n16032_ & new_n16037_;
  assign new_n16039_ = new_n8945_ & new_n15982_;
  assign new_n16040_ = new_n8934_ & new_n15982_;
  assign new_n16041_ = new_n8943_ & new_n15982_;
  assign new_n16042_ = ~new_n16040_ & ~new_n16041_;
  assign new_n16043_ = ~new_n16039_ & new_n16042_;
  assign new_n16044_ = A200 & new_n1781_;
  assign new_n16045_ = new_n4983_ & new_n16044_;
  assign new_n16046_ = new_n8617_ & new_n16045_;
  assign new_n16047_ = new_n8628_ & new_n16045_;
  assign new_n16048_ = ~new_n16046_ & ~new_n16047_;
  assign new_n16049_ = new_n16043_ & new_n16048_;
  assign new_n16050_ = new_n16038_ & new_n16049_;
  assign new_n16051_ = new_n16027_ & new_n16050_;
  assign new_n16052_ = new_n16004_ & new_n16051_;
  assign new_n16053_ = new_n8637_ & new_n16045_;
  assign new_n16054_ = new_n8630_ & new_n16045_;
  assign new_n16055_ = new_n8625_ & new_n16045_;
  assign new_n16056_ = ~new_n16054_ & ~new_n16055_;
  assign new_n16057_ = ~new_n16053_ & new_n16056_;
  assign new_n16058_ = new_n8648_ & new_n16045_;
  assign new_n16059_ = new_n8639_ & new_n16045_;
  assign new_n16060_ = new_n8635_ & new_n16045_;
  assign new_n16061_ = ~new_n16059_ & ~new_n16060_;
  assign new_n16062_ = ~new_n16058_ & new_n16061_;
  assign new_n16063_ = new_n16057_ & new_n16062_;
  assign new_n16064_ = new_n8657_ & new_n16045_;
  assign new_n16065_ = new_n8650_ & new_n16045_;
  assign new_n16066_ = new_n8646_ & new_n16045_;
  assign new_n16067_ = ~new_n16065_ & ~new_n16066_;
  assign new_n16068_ = ~new_n16064_ & new_n16067_;
  assign new_n16069_ = new_n8667_ & new_n16045_;
  assign new_n16070_ = new_n8659_ & new_n16045_;
  assign new_n16071_ = new_n8655_ & new_n16045_;
  assign new_n16072_ = ~new_n16070_ & ~new_n16071_;
  assign new_n16073_ = ~new_n16069_ & new_n16072_;
  assign new_n16074_ = new_n16068_ & new_n16073_;
  assign new_n16075_ = new_n16063_ & new_n16074_;
  assign new_n16076_ = new_n8678_ & new_n16045_;
  assign new_n16077_ = new_n8670_ & new_n16045_;
  assign new_n16078_ = new_n8665_ & new_n16045_;
  assign new_n16079_ = ~new_n16077_ & ~new_n16078_;
  assign new_n16080_ = ~new_n16076_ & new_n16079_;
  assign new_n16081_ = new_n8692_ & new_n16045_;
  assign new_n16082_ = new_n8681_ & new_n16045_;
  assign new_n16083_ = new_n8675_ & new_n16045_;
  assign new_n16084_ = ~new_n16082_ & ~new_n16083_;
  assign new_n16085_ = ~new_n16081_ & new_n16084_;
  assign new_n16086_ = new_n16080_ & new_n16085_;
  assign new_n16087_ = new_n8699_ & new_n16045_;
  assign new_n16088_ = new_n8694_ & new_n16045_;
  assign new_n16089_ = new_n8689_ & new_n16045_;
  assign new_n16090_ = ~new_n16088_ & ~new_n16089_;
  assign new_n16091_ = ~new_n16087_ & new_n16090_;
  assign new_n16092_ = new_n8701_ & new_n16045_;
  assign new_n16093_ = A200 & new_n1795_;
  assign new_n16094_ = new_n4983_ & new_n16093_;
  assign new_n16095_ = new_n8617_ & new_n16094_;
  assign new_n16096_ = ~new_n16092_ & ~new_n16095_;
  assign new_n16097_ = new_n16091_ & new_n16096_;
  assign new_n16098_ = new_n16086_ & new_n16097_;
  assign new_n16099_ = new_n16075_ & new_n16098_;
  assign new_n16100_ = new_n8625_ & new_n16094_;
  assign new_n16101_ = new_n8628_ & new_n16094_;
  assign new_n16102_ = new_n8630_ & new_n16094_;
  assign new_n16103_ = ~new_n16101_ & ~new_n16102_;
  assign new_n16104_ = ~new_n16100_ & new_n16103_;
  assign new_n16105_ = new_n8635_ & new_n16094_;
  assign new_n16106_ = new_n8637_ & new_n16094_;
  assign new_n16107_ = new_n8639_ & new_n16094_;
  assign new_n16108_ = ~new_n16106_ & ~new_n16107_;
  assign new_n16109_ = ~new_n16105_ & new_n16108_;
  assign new_n16110_ = new_n16104_ & new_n16109_;
  assign new_n16111_ = new_n8646_ & new_n16094_;
  assign new_n16112_ = new_n8648_ & new_n16094_;
  assign new_n16113_ = new_n8650_ & new_n16094_;
  assign new_n16114_ = ~new_n16112_ & ~new_n16113_;
  assign new_n16115_ = ~new_n16111_ & new_n16114_;
  assign new_n16116_ = new_n8655_ & new_n16094_;
  assign new_n16117_ = new_n8657_ & new_n16094_;
  assign new_n16118_ = new_n8659_ & new_n16094_;
  assign new_n16119_ = ~new_n16117_ & ~new_n16118_;
  assign new_n16120_ = ~new_n16116_ & new_n16119_;
  assign new_n16121_ = new_n16115_ & new_n16120_;
  assign new_n16122_ = new_n16110_ & new_n16121_;
  assign new_n16123_ = new_n8665_ & new_n16094_;
  assign new_n16124_ = new_n8667_ & new_n16094_;
  assign new_n16125_ = new_n8670_ & new_n16094_;
  assign new_n16126_ = ~new_n16124_ & ~new_n16125_;
  assign new_n16127_ = ~new_n16123_ & new_n16126_;
  assign new_n16128_ = new_n8675_ & new_n16094_;
  assign new_n16129_ = new_n8678_ & new_n16094_;
  assign new_n16130_ = new_n8681_ & new_n16094_;
  assign new_n16131_ = ~new_n16129_ & ~new_n16130_;
  assign new_n16132_ = ~new_n16128_ & new_n16131_;
  assign new_n16133_ = new_n16127_ & new_n16132_;
  assign new_n16134_ = new_n8689_ & new_n16094_;
  assign new_n16135_ = new_n8692_ & new_n16094_;
  assign new_n16136_ = new_n8694_ & new_n16094_;
  assign new_n16137_ = ~new_n16135_ & ~new_n16136_;
  assign new_n16138_ = ~new_n16134_ & new_n16137_;
  assign new_n16139_ = new_n8699_ & new_n16094_;
  assign new_n16140_ = new_n8701_ & new_n16094_;
  assign new_n16141_ = ~new_n16139_ & ~new_n16140_;
  assign new_n16142_ = new_n16138_ & new_n16141_;
  assign new_n16143_ = new_n16133_ & new_n16142_;
  assign new_n16144_ = new_n16122_ & new_n16143_;
  assign new_n16145_ = new_n16099_ & new_n16144_;
  assign new_n16146_ = new_n16052_ & new_n16145_;
  assign new_n16147_ = new_n15957_ & new_n16146_;
  assign new_n16148_ = new_n15766_ & new_n16147_;
  assign new_n16149_ = new_n15389_ & new_n16148_;
  assign new_n16150_ = new_n14634_ & new_n16149_;
  assign new_n16151_ = A200 & new_n1804_;
  assign new_n16152_ = new_n4983_ & new_n16151_;
  assign new_n16153_ = new_n8630_ & new_n16152_;
  assign new_n16154_ = new_n8617_ & new_n16152_;
  assign new_n16155_ = new_n8628_ & new_n16152_;
  assign new_n16156_ = ~new_n16154_ & ~new_n16155_;
  assign new_n16157_ = ~new_n16153_ & new_n16156_;
  assign new_n16158_ = new_n8639_ & new_n16152_;
  assign new_n16159_ = new_n8625_ & new_n16152_;
  assign new_n16160_ = new_n8637_ & new_n16152_;
  assign new_n16161_ = ~new_n16159_ & ~new_n16160_;
  assign new_n16162_ = ~new_n16158_ & new_n16161_;
  assign new_n16163_ = new_n16157_ & new_n16162_;
  assign new_n16164_ = new_n8650_ & new_n16152_;
  assign new_n16165_ = new_n8635_ & new_n16152_;
  assign new_n16166_ = new_n8648_ & new_n16152_;
  assign new_n16167_ = ~new_n16165_ & ~new_n16166_;
  assign new_n16168_ = ~new_n16164_ & new_n16167_;
  assign new_n16169_ = new_n8659_ & new_n16152_;
  assign new_n16170_ = new_n8646_ & new_n16152_;
  assign new_n16171_ = new_n8657_ & new_n16152_;
  assign new_n16172_ = ~new_n16170_ & ~new_n16171_;
  assign new_n16173_ = ~new_n16169_ & new_n16172_;
  assign new_n16174_ = new_n16168_ & new_n16173_;
  assign new_n16175_ = new_n16163_ & new_n16174_;
  assign new_n16176_ = new_n8670_ & new_n16152_;
  assign new_n16177_ = new_n8655_ & new_n16152_;
  assign new_n16178_ = new_n8667_ & new_n16152_;
  assign new_n16179_ = ~new_n16177_ & ~new_n16178_;
  assign new_n16180_ = ~new_n16176_ & new_n16179_;
  assign new_n16181_ = new_n8681_ & new_n16152_;
  assign new_n16182_ = new_n8665_ & new_n16152_;
  assign new_n16183_ = new_n8678_ & new_n16152_;
  assign new_n16184_ = ~new_n16182_ & ~new_n16183_;
  assign new_n16185_ = ~new_n16181_ & new_n16184_;
  assign new_n16186_ = new_n16180_ & new_n16185_;
  assign new_n16187_ = new_n8694_ & new_n16152_;
  assign new_n16188_ = new_n8675_ & new_n16152_;
  assign new_n16189_ = new_n8692_ & new_n16152_;
  assign new_n16190_ = ~new_n16188_ & ~new_n16189_;
  assign new_n16191_ = ~new_n16187_ & new_n16190_;
  assign new_n16192_ = new_n8701_ & new_n16152_;
  assign new_n16193_ = new_n8689_ & new_n16152_;
  assign new_n16194_ = new_n8699_ & new_n16152_;
  assign new_n16195_ = ~new_n16193_ & ~new_n16194_;
  assign new_n16196_ = ~new_n16192_ & new_n16195_;
  assign new_n16197_ = new_n16191_ & new_n16196_;
  assign new_n16198_ = new_n16186_ & new_n16197_;
  assign new_n16199_ = new_n16175_ & new_n16198_;
  assign new_n16200_ = A200 & new_n1812_;
  assign new_n16201_ = new_n4983_ & new_n16200_;
  assign new_n16202_ = new_n8630_ & new_n16201_;
  assign new_n16203_ = new_n8617_ & new_n16201_;
  assign new_n16204_ = new_n8628_ & new_n16201_;
  assign new_n16205_ = ~new_n16203_ & ~new_n16204_;
  assign new_n16206_ = ~new_n16202_ & new_n16205_;
  assign new_n16207_ = new_n8639_ & new_n16201_;
  assign new_n16208_ = new_n8625_ & new_n16201_;
  assign new_n16209_ = new_n8637_ & new_n16201_;
  assign new_n16210_ = ~new_n16208_ & ~new_n16209_;
  assign new_n16211_ = ~new_n16207_ & new_n16210_;
  assign new_n16212_ = new_n16206_ & new_n16211_;
  assign new_n16213_ = new_n8650_ & new_n16201_;
  assign new_n16214_ = new_n8635_ & new_n16201_;
  assign new_n16215_ = new_n8648_ & new_n16201_;
  assign new_n16216_ = ~new_n16214_ & ~new_n16215_;
  assign new_n16217_ = ~new_n16213_ & new_n16216_;
  assign new_n16218_ = new_n8659_ & new_n16201_;
  assign new_n16219_ = new_n8646_ & new_n16201_;
  assign new_n16220_ = new_n8657_ & new_n16201_;
  assign new_n16221_ = ~new_n16219_ & ~new_n16220_;
  assign new_n16222_ = ~new_n16218_ & new_n16221_;
  assign new_n16223_ = new_n16217_ & new_n16222_;
  assign new_n16224_ = new_n16212_ & new_n16223_;
  assign new_n16225_ = new_n8670_ & new_n16201_;
  assign new_n16226_ = new_n8655_ & new_n16201_;
  assign new_n16227_ = new_n8667_ & new_n16201_;
  assign new_n16228_ = ~new_n16226_ & ~new_n16227_;
  assign new_n16229_ = ~new_n16225_ & new_n16228_;
  assign new_n16230_ = new_n8681_ & new_n16201_;
  assign new_n16231_ = new_n8665_ & new_n16201_;
  assign new_n16232_ = new_n8678_ & new_n16201_;
  assign new_n16233_ = ~new_n16231_ & ~new_n16232_;
  assign new_n16234_ = ~new_n16230_ & new_n16233_;
  assign new_n16235_ = new_n16229_ & new_n16234_;
  assign new_n16236_ = new_n8694_ & new_n16201_;
  assign new_n16237_ = new_n8675_ & new_n16201_;
  assign new_n16238_ = new_n8692_ & new_n16201_;
  assign new_n16239_ = ~new_n16237_ & ~new_n16238_;
  assign new_n16240_ = ~new_n16236_ & new_n16239_;
  assign new_n16241_ = new_n8689_ & new_n16201_;
  assign new_n16242_ = new_n8699_ & new_n16201_;
  assign new_n16243_ = ~new_n16241_ & ~new_n16242_;
  assign new_n16244_ = new_n16240_ & new_n16243_;
  assign new_n16245_ = new_n16235_ & new_n16244_;
  assign new_n16246_ = new_n16224_ & new_n16245_;
  assign new_n16247_ = new_n16199_ & new_n16246_;
  assign new_n16248_ = A200 & new_n504_;
  assign new_n16249_ = new_n4983_ & new_n16248_;
  assign new_n16250_ = new_n8853_ & new_n16249_;
  assign new_n16251_ = new_n8701_ & new_n16201_;
  assign new_n16252_ = new_n8845_ & new_n16249_;
  assign new_n16253_ = ~new_n16251_ & ~new_n16252_;
  assign new_n16254_ = ~new_n16250_ & new_n16253_;
  assign new_n16255_ = new_n8864_ & new_n16249_;
  assign new_n16256_ = new_n8855_ & new_n16249_;
  assign new_n16257_ = new_n8851_ & new_n16249_;
  assign new_n16258_ = ~new_n16256_ & ~new_n16257_;
  assign new_n16259_ = ~new_n16255_ & new_n16258_;
  assign new_n16260_ = new_n16254_ & new_n16259_;
  assign new_n16261_ = new_n8872_ & new_n16249_;
  assign new_n16262_ = new_n8866_ & new_n16249_;
  assign new_n16263_ = new_n8862_ & new_n16249_;
  assign new_n16264_ = ~new_n16262_ & ~new_n16263_;
  assign new_n16265_ = ~new_n16261_ & new_n16264_;
  assign new_n16266_ = new_n8882_ & new_n16249_;
  assign new_n16267_ = new_n8874_ & new_n16249_;
  assign new_n16268_ = new_n8870_ & new_n16249_;
  assign new_n16269_ = ~new_n16267_ & ~new_n16268_;
  assign new_n16270_ = ~new_n16266_ & new_n16269_;
  assign new_n16271_ = new_n16265_ & new_n16270_;
  assign new_n16272_ = new_n16260_ & new_n16271_;
  assign new_n16273_ = new_n8888_ & new_n16249_;
  assign new_n16274_ = new_n8884_ & new_n16249_;
  assign new_n16275_ = new_n8880_ & new_n16249_;
  assign new_n16276_ = ~new_n16274_ & ~new_n16275_;
  assign new_n16277_ = ~new_n16273_ & new_n16276_;
  assign new_n16278_ = new_n8900_ & new_n16249_;
  assign new_n16279_ = new_n8890_ & new_n16249_;
  assign new_n16280_ = new_n8898_ & new_n16249_;
  assign new_n16281_ = ~new_n16279_ & ~new_n16280_;
  assign new_n16282_ = ~new_n16278_ & new_n16281_;
  assign new_n16283_ = new_n16277_ & new_n16282_;
  assign new_n16284_ = new_n8909_ & new_n16249_;
  assign new_n16285_ = new_n8896_ & new_n16249_;
  assign new_n16286_ = new_n8907_ & new_n16249_;
  assign new_n16287_ = ~new_n16285_ & ~new_n16286_;
  assign new_n16288_ = ~new_n16284_ & new_n16287_;
  assign new_n16289_ = new_n8905_ & new_n16249_;
  assign new_n16290_ = new_n8916_ & new_n16249_;
  assign new_n16291_ = ~new_n16289_ & ~new_n16290_;
  assign new_n16292_ = new_n16288_ & new_n16291_;
  assign new_n16293_ = new_n16283_ & new_n16292_;
  assign new_n16294_ = new_n16272_ & new_n16293_;
  assign new_n16295_ = new_n8925_ & new_n16249_;
  assign new_n16296_ = new_n8918_ & new_n16249_;
  assign new_n16297_ = new_n8914_ & new_n16249_;
  assign new_n16298_ = ~new_n16296_ & ~new_n16297_;
  assign new_n16299_ = ~new_n16295_ & new_n16298_;
  assign new_n16300_ = new_n8936_ & new_n16249_;
  assign new_n16301_ = new_n8927_ & new_n16249_;
  assign new_n16302_ = new_n8923_ & new_n16249_;
  assign new_n16303_ = ~new_n16301_ & ~new_n16302_;
  assign new_n16304_ = ~new_n16300_ & new_n16303_;
  assign new_n16305_ = new_n16299_ & new_n16304_;
  assign new_n16306_ = new_n8943_ & new_n16249_;
  assign new_n16307_ = new_n8938_ & new_n16249_;
  assign new_n16308_ = new_n8934_ & new_n16249_;
  assign new_n16309_ = ~new_n16307_ & ~new_n16308_;
  assign new_n16310_ = ~new_n16306_ & new_n16309_;
  assign new_n16311_ = ~A203 & new_n1781_;
  assign new_n16312_ = new_n4992_ & new_n16311_;
  assign new_n16313_ = new_n8628_ & new_n16312_;
  assign new_n16314_ = new_n8945_ & new_n16249_;
  assign new_n16315_ = new_n8617_ & new_n16312_;
  assign new_n16316_ = ~new_n16314_ & ~new_n16315_;
  assign new_n16317_ = ~new_n16313_ & new_n16316_;
  assign new_n16318_ = new_n16310_ & new_n16317_;
  assign new_n16319_ = new_n16305_ & new_n16318_;
  assign new_n16320_ = new_n8637_ & new_n16312_;
  assign new_n16321_ = new_n8630_ & new_n16312_;
  assign new_n16322_ = new_n8625_ & new_n16312_;
  assign new_n16323_ = ~new_n16321_ & ~new_n16322_;
  assign new_n16324_ = ~new_n16320_ & new_n16323_;
  assign new_n16325_ = new_n8648_ & new_n16312_;
  assign new_n16326_ = new_n8639_ & new_n16312_;
  assign new_n16327_ = new_n8635_ & new_n16312_;
  assign new_n16328_ = ~new_n16326_ & ~new_n16327_;
  assign new_n16329_ = ~new_n16325_ & new_n16328_;
  assign new_n16330_ = new_n16324_ & new_n16329_;
  assign new_n16331_ = new_n8657_ & new_n16312_;
  assign new_n16332_ = new_n8650_ & new_n16312_;
  assign new_n16333_ = new_n8646_ & new_n16312_;
  assign new_n16334_ = ~new_n16332_ & ~new_n16333_;
  assign new_n16335_ = ~new_n16331_ & new_n16334_;
  assign new_n16336_ = new_n8659_ & new_n16312_;
  assign new_n16337_ = new_n8655_ & new_n16312_;
  assign new_n16338_ = ~new_n16336_ & ~new_n16337_;
  assign new_n16339_ = new_n16335_ & new_n16338_;
  assign new_n16340_ = new_n16330_ & new_n16339_;
  assign new_n16341_ = new_n16319_ & new_n16340_;
  assign new_n16342_ = new_n16294_ & new_n16341_;
  assign new_n16343_ = new_n16247_ & new_n16342_;
  assign new_n16344_ = new_n8665_ & new_n16312_;
  assign new_n16345_ = new_n8667_ & new_n16312_;
  assign new_n16346_ = new_n8670_ & new_n16312_;
  assign new_n16347_ = ~new_n16345_ & ~new_n16346_;
  assign new_n16348_ = ~new_n16344_ & new_n16347_;
  assign new_n16349_ = new_n8675_ & new_n16312_;
  assign new_n16350_ = new_n8678_ & new_n16312_;
  assign new_n16351_ = new_n8681_ & new_n16312_;
  assign new_n16352_ = ~new_n16350_ & ~new_n16351_;
  assign new_n16353_ = ~new_n16349_ & new_n16352_;
  assign new_n16354_ = new_n16348_ & new_n16353_;
  assign new_n16355_ = new_n8689_ & new_n16312_;
  assign new_n16356_ = new_n8692_ & new_n16312_;
  assign new_n16357_ = new_n8694_ & new_n16312_;
  assign new_n16358_ = ~new_n16356_ & ~new_n16357_;
  assign new_n16359_ = ~new_n16355_ & new_n16358_;
  assign new_n16360_ = ~A203 & new_n1795_;
  assign new_n16361_ = new_n4992_ & new_n16360_;
  assign new_n16362_ = new_n8617_ & new_n16361_;
  assign new_n16363_ = new_n8699_ & new_n16312_;
  assign new_n16364_ = new_n8701_ & new_n16312_;
  assign new_n16365_ = ~new_n16363_ & ~new_n16364_;
  assign new_n16366_ = ~new_n16362_ & new_n16365_;
  assign new_n16367_ = new_n16359_ & new_n16366_;
  assign new_n16368_ = new_n16354_ & new_n16367_;
  assign new_n16369_ = new_n8625_ & new_n16361_;
  assign new_n16370_ = new_n8628_ & new_n16361_;
  assign new_n16371_ = new_n8630_ & new_n16361_;
  assign new_n16372_ = ~new_n16370_ & ~new_n16371_;
  assign new_n16373_ = ~new_n16369_ & new_n16372_;
  assign new_n16374_ = new_n8635_ & new_n16361_;
  assign new_n16375_ = new_n8637_ & new_n16361_;
  assign new_n16376_ = new_n8639_ & new_n16361_;
  assign new_n16377_ = ~new_n16375_ & ~new_n16376_;
  assign new_n16378_ = ~new_n16374_ & new_n16377_;
  assign new_n16379_ = new_n16373_ & new_n16378_;
  assign new_n16380_ = new_n8646_ & new_n16361_;
  assign new_n16381_ = new_n8648_ & new_n16361_;
  assign new_n16382_ = new_n8650_ & new_n16361_;
  assign new_n16383_ = ~new_n16381_ & ~new_n16382_;
  assign new_n16384_ = ~new_n16380_ & new_n16383_;
  assign new_n16385_ = new_n8657_ & new_n16361_;
  assign new_n16386_ = new_n8659_ & new_n16361_;
  assign new_n16387_ = ~new_n16385_ & ~new_n16386_;
  assign new_n16388_ = new_n16384_ & new_n16387_;
  assign new_n16389_ = new_n16379_ & new_n16388_;
  assign new_n16390_ = new_n16368_ & new_n16389_;
  assign new_n16391_ = new_n8670_ & new_n16361_;
  assign new_n16392_ = new_n8655_ & new_n16361_;
  assign new_n16393_ = new_n8667_ & new_n16361_;
  assign new_n16394_ = ~new_n16392_ & ~new_n16393_;
  assign new_n16395_ = ~new_n16391_ & new_n16394_;
  assign new_n16396_ = new_n8681_ & new_n16361_;
  assign new_n16397_ = new_n8665_ & new_n16361_;
  assign new_n16398_ = new_n8678_ & new_n16361_;
  assign new_n16399_ = ~new_n16397_ & ~new_n16398_;
  assign new_n16400_ = ~new_n16396_ & new_n16399_;
  assign new_n16401_ = new_n16395_ & new_n16400_;
  assign new_n16402_ = new_n8694_ & new_n16361_;
  assign new_n16403_ = new_n8675_ & new_n16361_;
  assign new_n16404_ = new_n8692_ & new_n16361_;
  assign new_n16405_ = ~new_n16403_ & ~new_n16404_;
  assign new_n16406_ = ~new_n16402_ & new_n16405_;
  assign new_n16407_ = new_n8701_ & new_n16361_;
  assign new_n16408_ = new_n8689_ & new_n16361_;
  assign new_n16409_ = new_n8699_ & new_n16361_;
  assign new_n16410_ = ~new_n16408_ & ~new_n16409_;
  assign new_n16411_ = ~new_n16407_ & new_n16410_;
  assign new_n16412_ = new_n16406_ & new_n16411_;
  assign new_n16413_ = new_n16401_ & new_n16412_;
  assign new_n16414_ = ~A203 & new_n1804_;
  assign new_n16415_ = new_n4992_ & new_n16414_;
  assign new_n16416_ = new_n8630_ & new_n16415_;
  assign new_n16417_ = new_n8617_ & new_n16415_;
  assign new_n16418_ = new_n8628_ & new_n16415_;
  assign new_n16419_ = ~new_n16417_ & ~new_n16418_;
  assign new_n16420_ = ~new_n16416_ & new_n16419_;
  assign new_n16421_ = new_n8639_ & new_n16415_;
  assign new_n16422_ = new_n8625_ & new_n16415_;
  assign new_n16423_ = new_n8637_ & new_n16415_;
  assign new_n16424_ = ~new_n16422_ & ~new_n16423_;
  assign new_n16425_ = ~new_n16421_ & new_n16424_;
  assign new_n16426_ = new_n16420_ & new_n16425_;
  assign new_n16427_ = new_n8650_ & new_n16415_;
  assign new_n16428_ = new_n8635_ & new_n16415_;
  assign new_n16429_ = new_n8648_ & new_n16415_;
  assign new_n16430_ = ~new_n16428_ & ~new_n16429_;
  assign new_n16431_ = ~new_n16427_ & new_n16430_;
  assign new_n16432_ = new_n8646_ & new_n16415_;
  assign new_n16433_ = new_n8657_ & new_n16415_;
  assign new_n16434_ = ~new_n16432_ & ~new_n16433_;
  assign new_n16435_ = new_n16431_ & new_n16434_;
  assign new_n16436_ = new_n16426_ & new_n16435_;
  assign new_n16437_ = new_n16413_ & new_n16436_;
  assign new_n16438_ = new_n16390_ & new_n16437_;
  assign new_n16439_ = new_n8667_ & new_n16415_;
  assign new_n16440_ = new_n8659_ & new_n16415_;
  assign new_n16441_ = new_n8655_ & new_n16415_;
  assign new_n16442_ = ~new_n16440_ & ~new_n16441_;
  assign new_n16443_ = ~new_n16439_ & new_n16442_;
  assign new_n16444_ = new_n8678_ & new_n16415_;
  assign new_n16445_ = new_n8670_ & new_n16415_;
  assign new_n16446_ = new_n8665_ & new_n16415_;
  assign new_n16447_ = ~new_n16445_ & ~new_n16446_;
  assign new_n16448_ = ~new_n16444_ & new_n16447_;
  assign new_n16449_ = new_n16443_ & new_n16448_;
  assign new_n16450_ = new_n8692_ & new_n16415_;
  assign new_n16451_ = new_n8681_ & new_n16415_;
  assign new_n16452_ = new_n8675_ & new_n16415_;
  assign new_n16453_ = ~new_n16451_ & ~new_n16452_;
  assign new_n16454_ = ~new_n16450_ & new_n16453_;
  assign new_n16455_ = new_n8699_ & new_n16415_;
  assign new_n16456_ = new_n8694_ & new_n16415_;
  assign new_n16457_ = new_n8689_ & new_n16415_;
  assign new_n16458_ = ~new_n16456_ & ~new_n16457_;
  assign new_n16459_ = ~new_n16455_ & new_n16458_;
  assign new_n16460_ = new_n16454_ & new_n16459_;
  assign new_n16461_ = new_n16449_ & new_n16460_;
  assign new_n16462_ = ~A203 & new_n1812_;
  assign new_n16463_ = new_n4992_ & new_n16462_;
  assign new_n16464_ = new_n8628_ & new_n16463_;
  assign new_n16465_ = new_n8701_ & new_n16415_;
  assign new_n16466_ = new_n8617_ & new_n16463_;
  assign new_n16467_ = ~new_n16465_ & ~new_n16466_;
  assign new_n16468_ = ~new_n16464_ & new_n16467_;
  assign new_n16469_ = new_n8637_ & new_n16463_;
  assign new_n16470_ = new_n8630_ & new_n16463_;
  assign new_n16471_ = new_n8625_ & new_n16463_;
  assign new_n16472_ = ~new_n16470_ & ~new_n16471_;
  assign new_n16473_ = ~new_n16469_ & new_n16472_;
  assign new_n16474_ = new_n16468_ & new_n16473_;
  assign new_n16475_ = new_n8648_ & new_n16463_;
  assign new_n16476_ = new_n8639_ & new_n16463_;
  assign new_n16477_ = new_n8635_ & new_n16463_;
  assign new_n16478_ = ~new_n16476_ & ~new_n16477_;
  assign new_n16479_ = ~new_n16475_ & new_n16478_;
  assign new_n16480_ = new_n8650_ & new_n16463_;
  assign new_n16481_ = new_n8646_ & new_n16463_;
  assign new_n16482_ = ~new_n16480_ & ~new_n16481_;
  assign new_n16483_ = new_n16479_ & new_n16482_;
  assign new_n16484_ = new_n16474_ & new_n16483_;
  assign new_n16485_ = new_n16461_ & new_n16484_;
  assign new_n16486_ = new_n8655_ & new_n16463_;
  assign new_n16487_ = new_n8657_ & new_n16463_;
  assign new_n16488_ = new_n8659_ & new_n16463_;
  assign new_n16489_ = ~new_n16487_ & ~new_n16488_;
  assign new_n16490_ = ~new_n16486_ & new_n16489_;
  assign new_n16491_ = new_n8665_ & new_n16463_;
  assign new_n16492_ = new_n8667_ & new_n16463_;
  assign new_n16493_ = new_n8670_ & new_n16463_;
  assign new_n16494_ = ~new_n16492_ & ~new_n16493_;
  assign new_n16495_ = ~new_n16491_ & new_n16494_;
  assign new_n16496_ = new_n16490_ & new_n16495_;
  assign new_n16497_ = new_n8675_ & new_n16463_;
  assign new_n16498_ = new_n8678_ & new_n16463_;
  assign new_n16499_ = new_n8681_ & new_n16463_;
  assign new_n16500_ = ~new_n16498_ & ~new_n16499_;
  assign new_n16501_ = ~new_n16497_ & new_n16500_;
  assign new_n16502_ = new_n8689_ & new_n16463_;
  assign new_n16503_ = new_n8692_ & new_n16463_;
  assign new_n16504_ = new_n8694_ & new_n16463_;
  assign new_n16505_ = ~new_n16503_ & ~new_n16504_;
  assign new_n16506_ = ~new_n16502_ & new_n16505_;
  assign new_n16507_ = new_n16501_ & new_n16506_;
  assign new_n16508_ = new_n16496_ & new_n16507_;
  assign new_n16509_ = ~A203 & new_n504_;
  assign new_n16510_ = new_n4992_ & new_n16509_;
  assign new_n16511_ = new_n8845_ & new_n16510_;
  assign new_n16512_ = new_n8699_ & new_n16463_;
  assign new_n16513_ = new_n8701_ & new_n16463_;
  assign new_n16514_ = ~new_n16512_ & ~new_n16513_;
  assign new_n16515_ = ~new_n16511_ & new_n16514_;
  assign new_n16516_ = new_n8851_ & new_n16510_;
  assign new_n16517_ = new_n8853_ & new_n16510_;
  assign new_n16518_ = new_n8855_ & new_n16510_;
  assign new_n16519_ = ~new_n16517_ & ~new_n16518_;
  assign new_n16520_ = ~new_n16516_ & new_n16519_;
  assign new_n16521_ = new_n16515_ & new_n16520_;
  assign new_n16522_ = new_n8862_ & new_n16510_;
  assign new_n16523_ = new_n8864_ & new_n16510_;
  assign new_n16524_ = new_n8866_ & new_n16510_;
  assign new_n16525_ = ~new_n16523_ & ~new_n16524_;
  assign new_n16526_ = ~new_n16522_ & new_n16525_;
  assign new_n16527_ = new_n8872_ & new_n16510_;
  assign new_n16528_ = new_n8874_ & new_n16510_;
  assign new_n16529_ = ~new_n16527_ & ~new_n16528_;
  assign new_n16530_ = new_n16526_ & new_n16529_;
  assign new_n16531_ = new_n16521_ & new_n16530_;
  assign new_n16532_ = new_n16508_ & new_n16531_;
  assign new_n16533_ = new_n16485_ & new_n16532_;
  assign new_n16534_ = new_n16438_ & new_n16533_;
  assign new_n16535_ = new_n16343_ & new_n16534_;
  assign new_n16536_ = new_n8884_ & new_n16510_;
  assign new_n16537_ = new_n8870_ & new_n16510_;
  assign new_n16538_ = new_n8882_ & new_n16510_;
  assign new_n16539_ = ~new_n16537_ & ~new_n16538_;
  assign new_n16540_ = ~new_n16536_ & new_n16539_;
  assign new_n16541_ = new_n8890_ & new_n16510_;
  assign new_n16542_ = new_n8880_ & new_n16510_;
  assign new_n16543_ = new_n8888_ & new_n16510_;
  assign new_n16544_ = ~new_n16542_ & ~new_n16543_;
  assign new_n16545_ = ~new_n16541_ & new_n16544_;
  assign new_n16546_ = new_n16540_ & new_n16545_;
  assign new_n16547_ = new_n8896_ & new_n16510_;
  assign new_n16548_ = new_n8898_ & new_n16510_;
  assign new_n16549_ = new_n8900_ & new_n16510_;
  assign new_n16550_ = ~new_n16548_ & ~new_n16549_;
  assign new_n16551_ = ~new_n16547_ & new_n16550_;
  assign new_n16552_ = new_n8905_ & new_n16510_;
  assign new_n16553_ = new_n8907_ & new_n16510_;
  assign new_n16554_ = new_n8909_ & new_n16510_;
  assign new_n16555_ = ~new_n16553_ & ~new_n16554_;
  assign new_n16556_ = ~new_n16552_ & new_n16555_;
  assign new_n16557_ = new_n16551_ & new_n16556_;
  assign new_n16558_ = new_n16546_ & new_n16557_;
  assign new_n16559_ = new_n8914_ & new_n16510_;
  assign new_n16560_ = new_n8916_ & new_n16510_;
  assign new_n16561_ = new_n8918_ & new_n16510_;
  assign new_n16562_ = ~new_n16560_ & ~new_n16561_;
  assign new_n16563_ = ~new_n16559_ & new_n16562_;
  assign new_n16564_ = new_n8923_ & new_n16510_;
  assign new_n16565_ = new_n8925_ & new_n16510_;
  assign new_n16566_ = new_n8927_ & new_n16510_;
  assign new_n16567_ = ~new_n16565_ & ~new_n16566_;
  assign new_n16568_ = ~new_n16564_ & new_n16567_;
  assign new_n16569_ = new_n16563_ & new_n16568_;
  assign new_n16570_ = new_n8934_ & new_n16510_;
  assign new_n16571_ = new_n8936_ & new_n16510_;
  assign new_n16572_ = new_n8938_ & new_n16510_;
  assign new_n16573_ = ~new_n16571_ & ~new_n16572_;
  assign new_n16574_ = ~new_n16570_ & new_n16573_;
  assign new_n16575_ = A202 & new_n1781_;
  assign new_n16576_ = new_n4992_ & new_n16575_;
  assign new_n16577_ = new_n8617_ & new_n16576_;
  assign new_n16578_ = new_n8943_ & new_n16510_;
  assign new_n16579_ = new_n8945_ & new_n16510_;
  assign new_n16580_ = ~new_n16578_ & ~new_n16579_;
  assign new_n16581_ = ~new_n16577_ & new_n16580_;
  assign new_n16582_ = new_n16574_ & new_n16581_;
  assign new_n16583_ = new_n16569_ & new_n16582_;
  assign new_n16584_ = new_n16558_ & new_n16583_;
  assign new_n16585_ = new_n8625_ & new_n16576_;
  assign new_n16586_ = new_n8628_ & new_n16576_;
  assign new_n16587_ = new_n8630_ & new_n16576_;
  assign new_n16588_ = ~new_n16586_ & ~new_n16587_;
  assign new_n16589_ = ~new_n16585_ & new_n16588_;
  assign new_n16590_ = new_n8635_ & new_n16576_;
  assign new_n16591_ = new_n8637_ & new_n16576_;
  assign new_n16592_ = new_n8639_ & new_n16576_;
  assign new_n16593_ = ~new_n16591_ & ~new_n16592_;
  assign new_n16594_ = ~new_n16590_ & new_n16593_;
  assign new_n16595_ = new_n16589_ & new_n16594_;
  assign new_n16596_ = new_n8646_ & new_n16576_;
  assign new_n16597_ = new_n8648_ & new_n16576_;
  assign new_n16598_ = new_n8650_ & new_n16576_;
  assign new_n16599_ = ~new_n16597_ & ~new_n16598_;
  assign new_n16600_ = ~new_n16596_ & new_n16599_;
  assign new_n16601_ = new_n8655_ & new_n16576_;
  assign new_n16602_ = new_n8657_ & new_n16576_;
  assign new_n16603_ = new_n8659_ & new_n16576_;
  assign new_n16604_ = ~new_n16602_ & ~new_n16603_;
  assign new_n16605_ = ~new_n16601_ & new_n16604_;
  assign new_n16606_ = new_n16600_ & new_n16605_;
  assign new_n16607_ = new_n16595_ & new_n16606_;
  assign new_n16608_ = new_n8665_ & new_n16576_;
  assign new_n16609_ = new_n8667_ & new_n16576_;
  assign new_n16610_ = new_n8670_ & new_n16576_;
  assign new_n16611_ = ~new_n16609_ & ~new_n16610_;
  assign new_n16612_ = ~new_n16608_ & new_n16611_;
  assign new_n16613_ = new_n8675_ & new_n16576_;
  assign new_n16614_ = new_n8678_ & new_n16576_;
  assign new_n16615_ = new_n8681_ & new_n16576_;
  assign new_n16616_ = ~new_n16614_ & ~new_n16615_;
  assign new_n16617_ = ~new_n16613_ & new_n16616_;
  assign new_n16618_ = new_n16612_ & new_n16617_;
  assign new_n16619_ = new_n8689_ & new_n16576_;
  assign new_n16620_ = new_n8692_ & new_n16576_;
  assign new_n16621_ = new_n8694_ & new_n16576_;
  assign new_n16622_ = ~new_n16620_ & ~new_n16621_;
  assign new_n16623_ = ~new_n16619_ & new_n16622_;
  assign new_n16624_ = new_n8699_ & new_n16576_;
  assign new_n16625_ = new_n8701_ & new_n16576_;
  assign new_n16626_ = ~new_n16624_ & ~new_n16625_;
  assign new_n16627_ = new_n16623_ & new_n16626_;
  assign new_n16628_ = new_n16618_ & new_n16627_;
  assign new_n16629_ = new_n16607_ & new_n16628_;
  assign new_n16630_ = new_n16584_ & new_n16629_;
  assign new_n16631_ = A202 & new_n1795_;
  assign new_n16632_ = new_n4992_ & new_n16631_;
  assign new_n16633_ = new_n8630_ & new_n16632_;
  assign new_n16634_ = new_n8617_ & new_n16632_;
  assign new_n16635_ = new_n8628_ & new_n16632_;
  assign new_n16636_ = ~new_n16634_ & ~new_n16635_;
  assign new_n16637_ = ~new_n16633_ & new_n16636_;
  assign new_n16638_ = new_n8639_ & new_n16632_;
  assign new_n16639_ = new_n8625_ & new_n16632_;
  assign new_n16640_ = new_n8637_ & new_n16632_;
  assign new_n16641_ = ~new_n16639_ & ~new_n16640_;
  assign new_n16642_ = ~new_n16638_ & new_n16641_;
  assign new_n16643_ = new_n16637_ & new_n16642_;
  assign new_n16644_ = new_n8650_ & new_n16632_;
  assign new_n16645_ = new_n8635_ & new_n16632_;
  assign new_n16646_ = new_n8648_ & new_n16632_;
  assign new_n16647_ = ~new_n16645_ & ~new_n16646_;
  assign new_n16648_ = ~new_n16644_ & new_n16647_;
  assign new_n16649_ = new_n8659_ & new_n16632_;
  assign new_n16650_ = new_n8646_ & new_n16632_;
  assign new_n16651_ = new_n8657_ & new_n16632_;
  assign new_n16652_ = ~new_n16650_ & ~new_n16651_;
  assign new_n16653_ = ~new_n16649_ & new_n16652_;
  assign new_n16654_ = new_n16648_ & new_n16653_;
  assign new_n16655_ = new_n16643_ & new_n16654_;
  assign new_n16656_ = new_n8670_ & new_n16632_;
  assign new_n16657_ = new_n8655_ & new_n16632_;
  assign new_n16658_ = new_n8667_ & new_n16632_;
  assign new_n16659_ = ~new_n16657_ & ~new_n16658_;
  assign new_n16660_ = ~new_n16656_ & new_n16659_;
  assign new_n16661_ = new_n8681_ & new_n16632_;
  assign new_n16662_ = new_n8665_ & new_n16632_;
  assign new_n16663_ = new_n8678_ & new_n16632_;
  assign new_n16664_ = ~new_n16662_ & ~new_n16663_;
  assign new_n16665_ = ~new_n16661_ & new_n16664_;
  assign new_n16666_ = new_n16660_ & new_n16665_;
  assign new_n16667_ = new_n8694_ & new_n16632_;
  assign new_n16668_ = new_n8675_ & new_n16632_;
  assign new_n16669_ = new_n8692_ & new_n16632_;
  assign new_n16670_ = ~new_n16668_ & ~new_n16669_;
  assign new_n16671_ = ~new_n16667_ & new_n16670_;
  assign new_n16672_ = new_n8689_ & new_n16632_;
  assign new_n16673_ = new_n8699_ & new_n16632_;
  assign new_n16674_ = ~new_n16672_ & ~new_n16673_;
  assign new_n16675_ = new_n16671_ & new_n16674_;
  assign new_n16676_ = new_n16666_ & new_n16675_;
  assign new_n16677_ = new_n16655_ & new_n16676_;
  assign new_n16678_ = A202 & new_n1804_;
  assign new_n16679_ = new_n4992_ & new_n16678_;
  assign new_n16680_ = new_n8628_ & new_n16679_;
  assign new_n16681_ = new_n8701_ & new_n16632_;
  assign new_n16682_ = new_n8617_ & new_n16679_;
  assign new_n16683_ = ~new_n16681_ & ~new_n16682_;
  assign new_n16684_ = ~new_n16680_ & new_n16683_;
  assign new_n16685_ = new_n8637_ & new_n16679_;
  assign new_n16686_ = new_n8630_ & new_n16679_;
  assign new_n16687_ = new_n8625_ & new_n16679_;
  assign new_n16688_ = ~new_n16686_ & ~new_n16687_;
  assign new_n16689_ = ~new_n16685_ & new_n16688_;
  assign new_n16690_ = new_n16684_ & new_n16689_;
  assign new_n16691_ = new_n8648_ & new_n16679_;
  assign new_n16692_ = new_n8639_ & new_n16679_;
  assign new_n16693_ = new_n8635_ & new_n16679_;
  assign new_n16694_ = ~new_n16692_ & ~new_n16693_;
  assign new_n16695_ = ~new_n16691_ & new_n16694_;
  assign new_n16696_ = new_n8657_ & new_n16679_;
  assign new_n16697_ = new_n8650_ & new_n16679_;
  assign new_n16698_ = new_n8646_ & new_n16679_;
  assign new_n16699_ = ~new_n16697_ & ~new_n16698_;
  assign new_n16700_ = ~new_n16696_ & new_n16699_;
  assign new_n16701_ = new_n16695_ & new_n16700_;
  assign new_n16702_ = new_n16690_ & new_n16701_;
  assign new_n16703_ = new_n8667_ & new_n16679_;
  assign new_n16704_ = new_n8659_ & new_n16679_;
  assign new_n16705_ = new_n8655_ & new_n16679_;
  assign new_n16706_ = ~new_n16704_ & ~new_n16705_;
  assign new_n16707_ = ~new_n16703_ & new_n16706_;
  assign new_n16708_ = new_n8678_ & new_n16679_;
  assign new_n16709_ = new_n8670_ & new_n16679_;
  assign new_n16710_ = new_n8665_ & new_n16679_;
  assign new_n16711_ = ~new_n16709_ & ~new_n16710_;
  assign new_n16712_ = ~new_n16708_ & new_n16711_;
  assign new_n16713_ = new_n16707_ & new_n16712_;
  assign new_n16714_ = new_n8692_ & new_n16679_;
  assign new_n16715_ = new_n8681_ & new_n16679_;
  assign new_n16716_ = new_n8675_ & new_n16679_;
  assign new_n16717_ = ~new_n16715_ & ~new_n16716_;
  assign new_n16718_ = ~new_n16714_ & new_n16717_;
  assign new_n16719_ = new_n8694_ & new_n16679_;
  assign new_n16720_ = new_n8689_ & new_n16679_;
  assign new_n16721_ = ~new_n16719_ & ~new_n16720_;
  assign new_n16722_ = new_n16718_ & new_n16721_;
  assign new_n16723_ = new_n16713_ & new_n16722_;
  assign new_n16724_ = new_n16702_ & new_n16723_;
  assign new_n16725_ = new_n16677_ & new_n16724_;
  assign new_n16726_ = new_n16630_ & new_n16725_;
  assign new_n16727_ = A202 & new_n1812_;
  assign new_n16728_ = new_n4992_ & new_n16727_;
  assign new_n16729_ = new_n8617_ & new_n16728_;
  assign new_n16730_ = new_n8699_ & new_n16679_;
  assign new_n16731_ = new_n8701_ & new_n16679_;
  assign new_n16732_ = ~new_n16730_ & ~new_n16731_;
  assign new_n16733_ = ~new_n16729_ & new_n16732_;
  assign new_n16734_ = new_n8625_ & new_n16728_;
  assign new_n16735_ = new_n8628_ & new_n16728_;
  assign new_n16736_ = new_n8630_ & new_n16728_;
  assign new_n16737_ = ~new_n16735_ & ~new_n16736_;
  assign new_n16738_ = ~new_n16734_ & new_n16737_;
  assign new_n16739_ = new_n16733_ & new_n16738_;
  assign new_n16740_ = new_n8635_ & new_n16728_;
  assign new_n16741_ = new_n8637_ & new_n16728_;
  assign new_n16742_ = new_n8639_ & new_n16728_;
  assign new_n16743_ = ~new_n16741_ & ~new_n16742_;
  assign new_n16744_ = ~new_n16740_ & new_n16743_;
  assign new_n16745_ = new_n8646_ & new_n16728_;
  assign new_n16746_ = new_n8648_ & new_n16728_;
  assign new_n16747_ = new_n8650_ & new_n16728_;
  assign new_n16748_ = ~new_n16746_ & ~new_n16747_;
  assign new_n16749_ = ~new_n16745_ & new_n16748_;
  assign new_n16750_ = new_n16744_ & new_n16749_;
  assign new_n16751_ = new_n16739_ & new_n16750_;
  assign new_n16752_ = new_n8655_ & new_n16728_;
  assign new_n16753_ = new_n8657_ & new_n16728_;
  assign new_n16754_ = new_n8659_ & new_n16728_;
  assign new_n16755_ = ~new_n16753_ & ~new_n16754_;
  assign new_n16756_ = ~new_n16752_ & new_n16755_;
  assign new_n16757_ = new_n8665_ & new_n16728_;
  assign new_n16758_ = new_n8667_ & new_n16728_;
  assign new_n16759_ = new_n8670_ & new_n16728_;
  assign new_n16760_ = ~new_n16758_ & ~new_n16759_;
  assign new_n16761_ = ~new_n16757_ & new_n16760_;
  assign new_n16762_ = new_n16756_ & new_n16761_;
  assign new_n16763_ = new_n8675_ & new_n16728_;
  assign new_n16764_ = new_n8678_ & new_n16728_;
  assign new_n16765_ = new_n8681_ & new_n16728_;
  assign new_n16766_ = ~new_n16764_ & ~new_n16765_;
  assign new_n16767_ = ~new_n16763_ & new_n16766_;
  assign new_n16768_ = new_n8692_ & new_n16728_;
  assign new_n16769_ = new_n8694_ & new_n16728_;
  assign new_n16770_ = ~new_n16768_ & ~new_n16769_;
  assign new_n16771_ = new_n16767_ & new_n16770_;
  assign new_n16772_ = new_n16762_ & new_n16771_;
  assign new_n16773_ = new_n16751_ & new_n16772_;
  assign new_n16774_ = new_n8701_ & new_n16728_;
  assign new_n16775_ = new_n8689_ & new_n16728_;
  assign new_n16776_ = new_n8699_ & new_n16728_;
  assign new_n16777_ = ~new_n16775_ & ~new_n16776_;
  assign new_n16778_ = ~new_n16774_ & new_n16777_;
  assign new_n16779_ = A202 & new_n504_;
  assign new_n16780_ = new_n4992_ & new_n16779_;
  assign new_n16781_ = new_n8855_ & new_n16780_;
  assign new_n16782_ = new_n8845_ & new_n16780_;
  assign new_n16783_ = new_n8853_ & new_n16780_;
  assign new_n16784_ = ~new_n16782_ & ~new_n16783_;
  assign new_n16785_ = ~new_n16781_ & new_n16784_;
  assign new_n16786_ = new_n16778_ & new_n16785_;
  assign new_n16787_ = new_n8866_ & new_n16780_;
  assign new_n16788_ = new_n8851_ & new_n16780_;
  assign new_n16789_ = new_n8864_ & new_n16780_;
  assign new_n16790_ = ~new_n16788_ & ~new_n16789_;
  assign new_n16791_ = ~new_n16787_ & new_n16790_;
  assign new_n16792_ = new_n8874_ & new_n16780_;
  assign new_n16793_ = new_n8862_ & new_n16780_;
  assign new_n16794_ = new_n8872_ & new_n16780_;
  assign new_n16795_ = ~new_n16793_ & ~new_n16794_;
  assign new_n16796_ = ~new_n16792_ & new_n16795_;
  assign new_n16797_ = new_n16791_ & new_n16796_;
  assign new_n16798_ = new_n16786_ & new_n16797_;
  assign new_n16799_ = new_n8884_ & new_n16780_;
  assign new_n16800_ = new_n8870_ & new_n16780_;
  assign new_n16801_ = new_n8882_ & new_n16780_;
  assign new_n16802_ = ~new_n16800_ & ~new_n16801_;
  assign new_n16803_ = ~new_n16799_ & new_n16802_;
  assign new_n16804_ = new_n8890_ & new_n16780_;
  assign new_n16805_ = new_n8880_ & new_n16780_;
  assign new_n16806_ = new_n8888_ & new_n16780_;
  assign new_n16807_ = ~new_n16805_ & ~new_n16806_;
  assign new_n16808_ = ~new_n16804_ & new_n16807_;
  assign new_n16809_ = new_n16803_ & new_n16808_;
  assign new_n16810_ = new_n8896_ & new_n16780_;
  assign new_n16811_ = new_n8898_ & new_n16780_;
  assign new_n16812_ = new_n8900_ & new_n16780_;
  assign new_n16813_ = ~new_n16811_ & ~new_n16812_;
  assign new_n16814_ = ~new_n16810_ & new_n16813_;
  assign new_n16815_ = new_n8907_ & new_n16780_;
  assign new_n16816_ = new_n8909_ & new_n16780_;
  assign new_n16817_ = ~new_n16815_ & ~new_n16816_;
  assign new_n16818_ = new_n16814_ & new_n16817_;
  assign new_n16819_ = new_n16809_ & new_n16818_;
  assign new_n16820_ = new_n16798_ & new_n16819_;
  assign new_n16821_ = new_n16773_ & new_n16820_;
  assign new_n16822_ = new_n8918_ & new_n16780_;
  assign new_n16823_ = new_n8905_ & new_n16780_;
  assign new_n16824_ = new_n8916_ & new_n16780_;
  assign new_n16825_ = ~new_n16823_ & ~new_n16824_;
  assign new_n16826_ = ~new_n16822_ & new_n16825_;
  assign new_n16827_ = new_n8927_ & new_n16780_;
  assign new_n16828_ = new_n8914_ & new_n16780_;
  assign new_n16829_ = new_n8925_ & new_n16780_;
  assign new_n16830_ = ~new_n16828_ & ~new_n16829_;
  assign new_n16831_ = ~new_n16827_ & new_n16830_;
  assign new_n16832_ = new_n16826_ & new_n16831_;
  assign new_n16833_ = new_n8938_ & new_n16780_;
  assign new_n16834_ = new_n8923_ & new_n16780_;
  assign new_n16835_ = new_n8936_ & new_n16780_;
  assign new_n16836_ = ~new_n16834_ & ~new_n16835_;
  assign new_n16837_ = ~new_n16833_ & new_n16836_;
  assign new_n16838_ = new_n8945_ & new_n16780_;
  assign new_n16839_ = new_n8934_ & new_n16780_;
  assign new_n16840_ = new_n8943_ & new_n16780_;
  assign new_n16841_ = ~new_n16839_ & ~new_n16840_;
  assign new_n16842_ = ~new_n16838_ & new_n16841_;
  assign new_n16843_ = new_n16837_ & new_n16842_;
  assign new_n16844_ = new_n16832_ & new_n16843_;
  assign new_n16845_ = ~A202 & new_n108_;
  assign new_n16846_ = new_n5013_ & new_n16845_;
  assign new_n16847_ = new_n9716_ & new_n16846_;
  assign new_n16848_ = new_n9718_ & new_n16846_;
  assign new_n16849_ = new_n9720_ & new_n16846_;
  assign new_n16850_ = ~new_n16848_ & ~new_n16849_;
  assign new_n16851_ = ~new_n16847_ & new_n16850_;
  assign new_n16852_ = new_n9727_ & new_n16846_;
  assign new_n16853_ = new_n9729_ & new_n16846_;
  assign new_n16854_ = new_n9731_ & new_n16846_;
  assign new_n16855_ = ~new_n16853_ & ~new_n16854_;
  assign new_n16856_ = ~new_n16852_ & new_n16855_;
  assign new_n16857_ = new_n16851_ & new_n16856_;
  assign new_n16858_ = new_n9735_ & new_n16846_;
  assign new_n16859_ = new_n9737_ & new_n16846_;
  assign new_n16860_ = new_n9739_ & new_n16846_;
  assign new_n16861_ = ~new_n16859_ & ~new_n16860_;
  assign new_n16862_ = ~new_n16858_ & new_n16861_;
  assign new_n16863_ = new_n9746_ & new_n16846_;
  assign new_n16864_ = new_n9748_ & new_n16846_;
  assign new_n16865_ = ~new_n16863_ & ~new_n16864_;
  assign new_n16866_ = new_n16862_ & new_n16865_;
  assign new_n16867_ = new_n16857_ & new_n16866_;
  assign new_n16868_ = new_n16844_ & new_n16867_;
  assign new_n16869_ = new_n9755_ & new_n16846_;
  assign new_n16870_ = new_n9744_ & new_n16846_;
  assign new_n16871_ = new_n9753_ & new_n16846_;
  assign new_n16872_ = ~new_n16870_ & ~new_n16871_;
  assign new_n16873_ = ~new_n16869_ & new_n16872_;
  assign new_n16874_ = new_n9761_ & new_n16846_;
  assign new_n16875_ = new_n9763_ & new_n16846_;
  assign new_n16876_ = new_n9765_ & new_n16846_;
  assign new_n16877_ = ~new_n16875_ & ~new_n16876_;
  assign new_n16878_ = ~new_n16874_ & new_n16877_;
  assign new_n16879_ = new_n16873_ & new_n16878_;
  assign new_n16880_ = new_n9769_ & new_n16846_;
  assign new_n16881_ = new_n9771_ & new_n16846_;
  assign new_n16882_ = new_n9773_ & new_n16846_;
  assign new_n16883_ = ~new_n16881_ & ~new_n16882_;
  assign new_n16884_ = ~new_n16880_ & new_n16883_;
  assign new_n16885_ = new_n9779_ & new_n16846_;
  assign new_n16886_ = new_n9781_ & new_n16846_;
  assign new_n16887_ = new_n9783_ & new_n16846_;
  assign new_n16888_ = ~new_n16886_ & ~new_n16887_;
  assign new_n16889_ = ~new_n16885_ & new_n16888_;
  assign new_n16890_ = new_n16884_ & new_n16889_;
  assign new_n16891_ = new_n16879_ & new_n16890_;
  assign new_n16892_ = new_n9788_ & new_n16846_;
  assign new_n16893_ = new_n9790_ & new_n16846_;
  assign new_n16894_ = new_n9792_ & new_n16846_;
  assign new_n16895_ = ~new_n16893_ & ~new_n16894_;
  assign new_n16896_ = ~new_n16892_ & new_n16895_;
  assign new_n16897_ = new_n9799_ & new_n16846_;
  assign new_n16898_ = new_n9801_ & new_n16846_;
  assign new_n16899_ = new_n9803_ & new_n16846_;
  assign new_n16900_ = ~new_n16898_ & ~new_n16899_;
  assign new_n16901_ = ~new_n16897_ & new_n16900_;
  assign new_n16902_ = new_n16896_ & new_n16901_;
  assign new_n16903_ = new_n9807_ & new_n16846_;
  assign new_n16904_ = new_n9809_ & new_n16846_;
  assign new_n16905_ = new_n9811_ & new_n16846_;
  assign new_n16906_ = ~new_n16904_ & ~new_n16905_;
  assign new_n16907_ = ~new_n16903_ & new_n16906_;
  assign new_n16908_ = ~A202 & new_n96_;
  assign new_n16909_ = new_n5013_ & new_n16908_;
  assign new_n16910_ = new_n9819_ & new_n16909_;
  assign new_n16911_ = new_n9821_ & new_n16909_;
  assign new_n16912_ = ~new_n16910_ & ~new_n16911_;
  assign new_n16913_ = new_n16907_ & new_n16912_;
  assign new_n16914_ = new_n16902_ & new_n16913_;
  assign new_n16915_ = new_n16891_ & new_n16914_;
  assign new_n16916_ = new_n16868_ & new_n16915_;
  assign new_n16917_ = new_n16821_ & new_n16916_;
  assign new_n16918_ = new_n16726_ & new_n16917_;
  assign new_n16919_ = new_n16535_ & new_n16918_;
  assign new_n16920_ = new_n9828_ & new_n16909_;
  assign new_n16921_ = new_n9817_ & new_n16909_;
  assign new_n16922_ = new_n9825_ & new_n16909_;
  assign new_n16923_ = ~new_n16921_ & ~new_n16922_;
  assign new_n16924_ = ~new_n16920_ & new_n16923_;
  assign new_n16925_ = new_n9840_ & new_n16909_;
  assign new_n16926_ = new_n9842_ & new_n16909_;
  assign new_n16927_ = new_n9844_ & new_n16909_;
  assign new_n16928_ = ~new_n16926_ & ~new_n16927_;
  assign new_n16929_ = ~new_n16925_ & new_n16928_;
  assign new_n16930_ = new_n16924_ & new_n16929_;
  assign new_n16931_ = new_n9848_ & new_n16909_;
  assign new_n16932_ = new_n9850_ & new_n16909_;
  assign new_n16933_ = new_n9852_ & new_n16909_;
  assign new_n16934_ = ~new_n16932_ & ~new_n16933_;
  assign new_n16935_ = ~new_n16931_ & new_n16934_;
  assign new_n16936_ = new_n9858_ & new_n16909_;
  assign new_n16937_ = new_n9860_ & new_n16909_;
  assign new_n16938_ = new_n9862_ & new_n16909_;
  assign new_n16939_ = ~new_n16937_ & ~new_n16938_;
  assign new_n16940_ = ~new_n16936_ & new_n16939_;
  assign new_n16941_ = new_n16935_ & new_n16940_;
  assign new_n16942_ = new_n16930_ & new_n16941_;
  assign new_n16943_ = new_n9866_ & new_n16909_;
  assign new_n16944_ = new_n9868_ & new_n16909_;
  assign new_n16945_ = new_n9870_ & new_n16909_;
  assign new_n16946_ = ~new_n16944_ & ~new_n16945_;
  assign new_n16947_ = ~new_n16943_ & new_n16946_;
  assign new_n16948_ = new_n9876_ & new_n16909_;
  assign new_n16949_ = new_n9878_ & new_n16909_;
  assign new_n16950_ = new_n9880_ & new_n16909_;
  assign new_n16951_ = ~new_n16949_ & ~new_n16950_;
  assign new_n16952_ = ~new_n16948_ & new_n16951_;
  assign new_n16953_ = new_n16947_ & new_n16952_;
  assign new_n16954_ = new_n9885_ & new_n16909_;
  assign new_n16955_ = new_n9887_ & new_n16909_;
  assign new_n16956_ = new_n9889_ & new_n16909_;
  assign new_n16957_ = ~new_n16955_ & ~new_n16956_;
  assign new_n16958_ = ~new_n16954_ & new_n16957_;
  assign new_n16959_ = new_n9895_ & new_n16909_;
  assign new_n16960_ = new_n9897_ & new_n16909_;
  assign new_n16961_ = new_n9899_ & new_n16909_;
  assign new_n16962_ = ~new_n16960_ & ~new_n16961_;
  assign new_n16963_ = ~new_n16959_ & new_n16962_;
  assign new_n16964_ = new_n16958_ & new_n16963_;
  assign new_n16965_ = new_n16953_ & new_n16964_;
  assign new_n16966_ = new_n16942_ & new_n16965_;
  assign new_n16967_ = new_n9904_ & new_n16909_;
  assign new_n16968_ = new_n9906_ & new_n16909_;
  assign new_n16969_ = new_n9908_ & new_n16909_;
  assign new_n16970_ = ~new_n16968_ & ~new_n16969_;
  assign new_n16971_ = ~new_n16967_ & new_n16970_;
  assign new_n16972_ = new_n9915_ & new_n16909_;
  assign new_n16973_ = new_n9917_ & new_n16909_;
  assign new_n16974_ = new_n9919_ & new_n16909_;
  assign new_n16975_ = ~new_n16973_ & ~new_n16974_;
  assign new_n16976_ = ~new_n16972_ & new_n16975_;
  assign new_n16977_ = new_n16971_ & new_n16976_;
  assign new_n16978_ = ~A202 & new_n4800_;
  assign new_n16979_ = new_n5013_ & new_n16978_;
  assign new_n16980_ = new_n9924_ & new_n16979_;
  assign new_n16981_ = new_n9926_ & new_n16979_;
  assign new_n16982_ = new_n9928_ & new_n16979_;
  assign new_n16983_ = ~new_n16981_ & ~new_n16982_;
  assign new_n16984_ = ~new_n16980_ & new_n16983_;
  assign new_n16985_ = new_n9934_ & new_n16979_;
  assign new_n16986_ = new_n9936_ & new_n16979_;
  assign new_n16987_ = new_n9938_ & new_n16979_;
  assign new_n16988_ = ~new_n16986_ & ~new_n16987_;
  assign new_n16989_ = ~new_n16985_ & new_n16988_;
  assign new_n16990_ = new_n16984_ & new_n16989_;
  assign new_n16991_ = new_n16977_ & new_n16990_;
  assign new_n16992_ = new_n9942_ & new_n16979_;
  assign new_n16993_ = new_n9944_ & new_n16979_;
  assign new_n16994_ = new_n9946_ & new_n16979_;
  assign new_n16995_ = ~new_n16993_ & ~new_n16994_;
  assign new_n16996_ = ~new_n16992_ & new_n16995_;
  assign new_n16997_ = new_n9952_ & new_n16979_;
  assign new_n16998_ = new_n9954_ & new_n16979_;
  assign new_n16999_ = new_n9956_ & new_n16979_;
  assign new_n17000_ = ~new_n16998_ & ~new_n16999_;
  assign new_n17001_ = ~new_n16997_ & new_n17000_;
  assign new_n17002_ = new_n16996_ & new_n17001_;
  assign new_n17003_ = new_n9961_ & new_n16979_;
  assign new_n17004_ = new_n9963_ & new_n16979_;
  assign new_n17005_ = new_n9965_ & new_n16979_;
  assign new_n17006_ = ~new_n17004_ & ~new_n17005_;
  assign new_n17007_ = ~new_n17003_ & new_n17006_;
  assign new_n17008_ = new_n9972_ & new_n16979_;
  assign new_n17009_ = new_n9974_ & new_n16979_;
  assign new_n17010_ = ~new_n17008_ & ~new_n17009_;
  assign new_n17011_ = new_n17007_ & new_n17010_;
  assign new_n17012_ = new_n17002_ & new_n17011_;
  assign new_n17013_ = new_n16991_ & new_n17012_;
  assign new_n17014_ = new_n16966_ & new_n17013_;
  assign new_n17015_ = new_n9980_ & new_n16979_;
  assign new_n17016_ = new_n9970_ & new_n16979_;
  assign new_n17017_ = new_n9978_ & new_n16979_;
  assign new_n17018_ = ~new_n17016_ & ~new_n17017_;
  assign new_n17019_ = ~new_n17015_ & new_n17018_;
  assign new_n17020_ = new_n9988_ & new_n16979_;
  assign new_n17021_ = new_n9990_ & new_n16979_;
  assign new_n17022_ = new_n9992_ & new_n16979_;
  assign new_n17023_ = ~new_n17021_ & ~new_n17022_;
  assign new_n17024_ = ~new_n17020_ & new_n17023_;
  assign new_n17025_ = new_n17019_ & new_n17024_;
  assign new_n17026_ = new_n9997_ & new_n16979_;
  assign new_n17027_ = new_n9999_ & new_n16979_;
  assign new_n17028_ = new_n10001_ & new_n16979_;
  assign new_n17029_ = ~new_n17027_ & ~new_n17028_;
  assign new_n17030_ = ~new_n17026_ & new_n17029_;
  assign new_n17031_ = new_n10007_ & new_n16979_;
  assign new_n17032_ = new_n10009_ & new_n16979_;
  assign new_n17033_ = new_n10011_ & new_n16979_;
  assign new_n17034_ = ~new_n17032_ & ~new_n17033_;
  assign new_n17035_ = ~new_n17031_ & new_n17034_;
  assign new_n17036_ = new_n17030_ & new_n17035_;
  assign new_n17037_ = new_n17025_ & new_n17036_;
  assign new_n17038_ = new_n10015_ & new_n16979_;
  assign new_n17039_ = new_n10017_ & new_n16979_;
  assign new_n17040_ = new_n10019_ & new_n16979_;
  assign new_n17041_ = ~new_n17039_ & ~new_n17040_;
  assign new_n17042_ = ~new_n17038_ & new_n17041_;
  assign new_n17043_ = new_n10026_ & new_n16979_;
  assign new_n17044_ = new_n10028_ & new_n16979_;
  assign new_n17045_ = new_n10030_ & new_n16979_;
  assign new_n17046_ = ~new_n17044_ & ~new_n17045_;
  assign new_n17047_ = ~new_n17043_ & new_n17046_;
  assign new_n17048_ = new_n17042_ & new_n17047_;
  assign new_n17049_ = new_n10035_ & new_n16979_;
  assign new_n17050_ = new_n10037_ & new_n16979_;
  assign new_n17051_ = new_n10039_ & new_n16979_;
  assign new_n17052_ = ~new_n17050_ & ~new_n17051_;
  assign new_n17053_ = ~new_n17049_ & new_n17052_;
  assign new_n17054_ = new_n10046_ & new_n16979_;
  assign new_n17055_ = new_n10048_ & new_n16979_;
  assign new_n17056_ = ~new_n17054_ & ~new_n17055_;
  assign new_n17057_ = new_n17053_ & new_n17056_;
  assign new_n17058_ = new_n17048_ & new_n17057_;
  assign new_n17059_ = new_n17037_ & new_n17058_;
  assign new_n17060_ = new_n10054_ & new_n16979_;
  assign new_n17061_ = new_n10044_ & new_n16979_;
  assign new_n17062_ = new_n10052_ & new_n16979_;
  assign new_n17063_ = ~new_n17061_ & ~new_n17062_;
  assign new_n17064_ = ~new_n17060_ & new_n17063_;
  assign new_n17065_ = new_n10061_ & new_n16979_;
  assign new_n17066_ = new_n10063_ & new_n16979_;
  assign new_n17067_ = new_n10065_ & new_n16979_;
  assign new_n17068_ = ~new_n17066_ & ~new_n17067_;
  assign new_n17069_ = ~new_n17065_ & new_n17068_;
  assign new_n17070_ = new_n17064_ & new_n17069_;
  assign new_n17071_ = new_n10069_ & new_n16979_;
  assign new_n17072_ = new_n10071_ & new_n16979_;
  assign new_n17073_ = new_n10073_ & new_n16979_;
  assign new_n17074_ = ~new_n17072_ & ~new_n17073_;
  assign new_n17075_ = ~new_n17071_ & new_n17074_;
  assign new_n17076_ = new_n10078_ & new_n16979_;
  assign new_n17077_ = new_n10080_ & new_n16979_;
  assign new_n17078_ = new_n10082_ & new_n16979_;
  assign new_n17079_ = ~new_n17077_ & ~new_n17078_;
  assign new_n17080_ = ~new_n17076_ & new_n17079_;
  assign new_n17081_ = new_n17075_ & new_n17080_;
  assign new_n17082_ = new_n17070_ & new_n17081_;
  assign new_n17083_ = new_n10087_ & new_n16979_;
  assign new_n17084_ = new_n10089_ & new_n16979_;
  assign new_n17085_ = new_n10091_ & new_n16979_;
  assign new_n17086_ = ~new_n17084_ & ~new_n17085_;
  assign new_n17087_ = ~new_n17083_ & new_n17086_;
  assign new_n17088_ = new_n10098_ & new_n16979_;
  assign new_n17089_ = new_n10100_ & new_n16979_;
  assign new_n17090_ = new_n10102_ & new_n16979_;
  assign new_n17091_ = ~new_n17089_ & ~new_n17090_;
  assign new_n17092_ = ~new_n17088_ & new_n17091_;
  assign new_n17093_ = new_n17087_ & new_n17092_;
  assign new_n17094_ = new_n10107_ & new_n16979_;
  assign new_n17095_ = new_n10109_ & new_n16979_;
  assign new_n17096_ = new_n10111_ & new_n16979_;
  assign new_n17097_ = ~new_n17095_ & ~new_n17096_;
  assign new_n17098_ = ~new_n17094_ & new_n17097_;
  assign new_n17099_ = new_n10118_ & new_n16979_;
  assign new_n17100_ = new_n10120_ & new_n16979_;
  assign new_n17101_ = ~new_n17099_ & ~new_n17100_;
  assign new_n17102_ = new_n17098_ & new_n17101_;
  assign new_n17103_ = new_n17093_ & new_n17102_;
  assign new_n17104_ = new_n17082_ & new_n17103_;
  assign new_n17105_ = new_n17059_ & new_n17104_;
  assign new_n17106_ = new_n17014_ & new_n17105_;
  assign new_n17107_ = new_n5752_ & new_n15778_;
  assign new_n17108_ = new_n8628_ & new_n17107_;
  assign new_n17109_ = new_n10116_ & new_n16979_;
  assign new_n17110_ = new_n8617_ & new_n17107_;
  assign new_n17111_ = ~new_n17109_ & ~new_n17110_;
  assign new_n17112_ = ~new_n17108_ & new_n17111_;
  assign new_n17113_ = new_n8637_ & new_n17107_;
  assign new_n17114_ = new_n8630_ & new_n17107_;
  assign new_n17115_ = new_n8625_ & new_n17107_;
  assign new_n17116_ = ~new_n17114_ & ~new_n17115_;
  assign new_n17117_ = ~new_n17113_ & new_n17116_;
  assign new_n17118_ = new_n17112_ & new_n17117_;
  assign new_n17119_ = new_n8648_ & new_n17107_;
  assign new_n17120_ = new_n8639_ & new_n17107_;
  assign new_n17121_ = new_n8635_ & new_n17107_;
  assign new_n17122_ = ~new_n17120_ & ~new_n17121_;
  assign new_n17123_ = ~new_n17119_ & new_n17122_;
  assign new_n17124_ = new_n8657_ & new_n17107_;
  assign new_n17125_ = new_n8650_ & new_n17107_;
  assign new_n17126_ = new_n8646_ & new_n17107_;
  assign new_n17127_ = ~new_n17125_ & ~new_n17126_;
  assign new_n17128_ = ~new_n17124_ & new_n17127_;
  assign new_n17129_ = new_n17123_ & new_n17128_;
  assign new_n17130_ = new_n17118_ & new_n17129_;
  assign new_n17131_ = new_n8667_ & new_n17107_;
  assign new_n17132_ = new_n8659_ & new_n17107_;
  assign new_n17133_ = new_n8655_ & new_n17107_;
  assign new_n17134_ = ~new_n17132_ & ~new_n17133_;
  assign new_n17135_ = ~new_n17131_ & new_n17134_;
  assign new_n17136_ = new_n8678_ & new_n17107_;
  assign new_n17137_ = new_n8670_ & new_n17107_;
  assign new_n17138_ = new_n8665_ & new_n17107_;
  assign new_n17139_ = ~new_n17137_ & ~new_n17138_;
  assign new_n17140_ = ~new_n17136_ & new_n17139_;
  assign new_n17141_ = new_n17135_ & new_n17140_;
  assign new_n17142_ = new_n8692_ & new_n17107_;
  assign new_n17143_ = new_n8681_ & new_n17107_;
  assign new_n17144_ = new_n8675_ & new_n17107_;
  assign new_n17145_ = ~new_n17143_ & ~new_n17144_;
  assign new_n17146_ = ~new_n17142_ & new_n17145_;
  assign new_n17147_ = new_n8694_ & new_n17107_;
  assign new_n17148_ = new_n8689_ & new_n17107_;
  assign new_n17149_ = ~new_n17147_ & ~new_n17148_;
  assign new_n17150_ = new_n17146_ & new_n17149_;
  assign new_n17151_ = new_n17141_ & new_n17150_;
  assign new_n17152_ = new_n17130_ & new_n17151_;
  assign new_n17153_ = new_n5752_ & new_n15830_;
  assign new_n17154_ = new_n8617_ & new_n17153_;
  assign new_n17155_ = new_n8699_ & new_n17107_;
  assign new_n17156_ = new_n8701_ & new_n17107_;
  assign new_n17157_ = ~new_n17155_ & ~new_n17156_;
  assign new_n17158_ = ~new_n17154_ & new_n17157_;
  assign new_n17159_ = new_n8625_ & new_n17153_;
  assign new_n17160_ = new_n8628_ & new_n17153_;
  assign new_n17161_ = new_n8630_ & new_n17153_;
  assign new_n17162_ = ~new_n17160_ & ~new_n17161_;
  assign new_n17163_ = ~new_n17159_ & new_n17162_;
  assign new_n17164_ = new_n17158_ & new_n17163_;
  assign new_n17165_ = new_n8635_ & new_n17153_;
  assign new_n17166_ = new_n8637_ & new_n17153_;
  assign new_n17167_ = new_n8639_ & new_n17153_;
  assign new_n17168_ = ~new_n17166_ & ~new_n17167_;
  assign new_n17169_ = ~new_n17165_ & new_n17168_;
  assign new_n17170_ = new_n8646_ & new_n17153_;
  assign new_n17171_ = new_n8648_ & new_n17153_;
  assign new_n17172_ = new_n8650_ & new_n17153_;
  assign new_n17173_ = ~new_n17171_ & ~new_n17172_;
  assign new_n17174_ = ~new_n17170_ & new_n17173_;
  assign new_n17175_ = new_n17169_ & new_n17174_;
  assign new_n17176_ = new_n17164_ & new_n17175_;
  assign new_n17177_ = new_n8655_ & new_n17153_;
  assign new_n17178_ = new_n8657_ & new_n17153_;
  assign new_n17179_ = new_n8659_ & new_n17153_;
  assign new_n17180_ = ~new_n17178_ & ~new_n17179_;
  assign new_n17181_ = ~new_n17177_ & new_n17180_;
  assign new_n17182_ = new_n8665_ & new_n17153_;
  assign new_n17183_ = new_n8667_ & new_n17153_;
  assign new_n17184_ = new_n8670_ & new_n17153_;
  assign new_n17185_ = ~new_n17183_ & ~new_n17184_;
  assign new_n17186_ = ~new_n17182_ & new_n17185_;
  assign new_n17187_ = new_n17181_ & new_n17186_;
  assign new_n17188_ = new_n8675_ & new_n17153_;
  assign new_n17189_ = new_n8678_ & new_n17153_;
  assign new_n17190_ = new_n8681_ & new_n17153_;
  assign new_n17191_ = ~new_n17189_ & ~new_n17190_;
  assign new_n17192_ = ~new_n17188_ & new_n17191_;
  assign new_n17193_ = new_n8692_ & new_n17153_;
  assign new_n17194_ = new_n8694_ & new_n17153_;
  assign new_n17195_ = ~new_n17193_ & ~new_n17194_;
  assign new_n17196_ = new_n17192_ & new_n17195_;
  assign new_n17197_ = new_n17187_ & new_n17196_;
  assign new_n17198_ = new_n17176_ & new_n17197_;
  assign new_n17199_ = new_n17152_ & new_n17198_;
  assign new_n17200_ = new_n8701_ & new_n17153_;
  assign new_n17201_ = new_n8689_ & new_n17153_;
  assign new_n17202_ = new_n8699_ & new_n17153_;
  assign new_n17203_ = ~new_n17201_ & ~new_n17202_;
  assign new_n17204_ = ~new_n17200_ & new_n17203_;
  assign new_n17205_ = new_n5752_ & new_n15878_;
  assign new_n17206_ = new_n8630_ & new_n17205_;
  assign new_n17207_ = new_n8617_ & new_n17205_;
  assign new_n17208_ = new_n8628_ & new_n17205_;
  assign new_n17209_ = ~new_n17207_ & ~new_n17208_;
  assign new_n17210_ = ~new_n17206_ & new_n17209_;
  assign new_n17211_ = new_n17204_ & new_n17210_;
  assign new_n17212_ = new_n8639_ & new_n17205_;
  assign new_n17213_ = new_n8625_ & new_n17205_;
  assign new_n17214_ = new_n8637_ & new_n17205_;
  assign new_n17215_ = ~new_n17213_ & ~new_n17214_;
  assign new_n17216_ = ~new_n17212_ & new_n17215_;
  assign new_n17217_ = new_n8650_ & new_n17205_;
  assign new_n17218_ = new_n8635_ & new_n17205_;
  assign new_n17219_ = new_n8648_ & new_n17205_;
  assign new_n17220_ = ~new_n17218_ & ~new_n17219_;
  assign new_n17221_ = ~new_n17217_ & new_n17220_;
  assign new_n17222_ = new_n17216_ & new_n17221_;
  assign new_n17223_ = new_n17211_ & new_n17222_;
  assign new_n17224_ = new_n8659_ & new_n17205_;
  assign new_n17225_ = new_n8646_ & new_n17205_;
  assign new_n17226_ = new_n8657_ & new_n17205_;
  assign new_n17227_ = ~new_n17225_ & ~new_n17226_;
  assign new_n17228_ = ~new_n17224_ & new_n17227_;
  assign new_n17229_ = new_n8670_ & new_n17205_;
  assign new_n17230_ = new_n8655_ & new_n17205_;
  assign new_n17231_ = new_n8667_ & new_n17205_;
  assign new_n17232_ = ~new_n17230_ & ~new_n17231_;
  assign new_n17233_ = ~new_n17229_ & new_n17232_;
  assign new_n17234_ = new_n17228_ & new_n17233_;
  assign new_n17235_ = new_n8681_ & new_n17205_;
  assign new_n17236_ = new_n8665_ & new_n17205_;
  assign new_n17237_ = new_n8678_ & new_n17205_;
  assign new_n17238_ = ~new_n17236_ & ~new_n17237_;
  assign new_n17239_ = ~new_n17235_ & new_n17238_;
  assign new_n17240_ = new_n8675_ & new_n17205_;
  assign new_n17241_ = new_n8692_ & new_n17205_;
  assign new_n17242_ = ~new_n17240_ & ~new_n17241_;
  assign new_n17243_ = new_n17239_ & new_n17242_;
  assign new_n17244_ = new_n17234_ & new_n17243_;
  assign new_n17245_ = new_n17223_ & new_n17244_;
  assign new_n17246_ = new_n8699_ & new_n17205_;
  assign new_n17247_ = new_n8694_ & new_n17205_;
  assign new_n17248_ = new_n8689_ & new_n17205_;
  assign new_n17249_ = ~new_n17247_ & ~new_n17248_;
  assign new_n17250_ = ~new_n17246_ & new_n17249_;
  assign new_n17251_ = new_n5752_ & new_n15925_;
  assign new_n17252_ = new_n8628_ & new_n17251_;
  assign new_n17253_ = new_n8701_ & new_n17205_;
  assign new_n17254_ = new_n8617_ & new_n17251_;
  assign new_n17255_ = ~new_n17253_ & ~new_n17254_;
  assign new_n17256_ = ~new_n17252_ & new_n17255_;
  assign new_n17257_ = new_n17250_ & new_n17256_;
  assign new_n17258_ = new_n8637_ & new_n17251_;
  assign new_n17259_ = new_n8630_ & new_n17251_;
  assign new_n17260_ = new_n8625_ & new_n17251_;
  assign new_n17261_ = ~new_n17259_ & ~new_n17260_;
  assign new_n17262_ = ~new_n17258_ & new_n17261_;
  assign new_n17263_ = new_n8648_ & new_n17251_;
  assign new_n17264_ = new_n8639_ & new_n17251_;
  assign new_n17265_ = new_n8635_ & new_n17251_;
  assign new_n17266_ = ~new_n17264_ & ~new_n17265_;
  assign new_n17267_ = ~new_n17263_ & new_n17266_;
  assign new_n17268_ = new_n17262_ & new_n17267_;
  assign new_n17269_ = new_n17257_ & new_n17268_;
  assign new_n17270_ = new_n8657_ & new_n17251_;
  assign new_n17271_ = new_n8650_ & new_n17251_;
  assign new_n17272_ = new_n8646_ & new_n17251_;
  assign new_n17273_ = ~new_n17271_ & ~new_n17272_;
  assign new_n17274_ = ~new_n17270_ & new_n17273_;
  assign new_n17275_ = new_n8667_ & new_n17251_;
  assign new_n17276_ = new_n8659_ & new_n17251_;
  assign new_n17277_ = new_n8655_ & new_n17251_;
  assign new_n17278_ = ~new_n17276_ & ~new_n17277_;
  assign new_n17279_ = ~new_n17275_ & new_n17278_;
  assign new_n17280_ = new_n17274_ & new_n17279_;
  assign new_n17281_ = new_n8678_ & new_n17251_;
  assign new_n17282_ = new_n8670_ & new_n17251_;
  assign new_n17283_ = new_n8665_ & new_n17251_;
  assign new_n17284_ = ~new_n17282_ & ~new_n17283_;
  assign new_n17285_ = ~new_n17281_ & new_n17284_;
  assign new_n17286_ = new_n8681_ & new_n17251_;
  assign new_n17287_ = new_n8675_ & new_n17251_;
  assign new_n17288_ = ~new_n17286_ & ~new_n17287_;
  assign new_n17289_ = new_n17285_ & new_n17288_;
  assign new_n17290_ = new_n17280_ & new_n17289_;
  assign new_n17291_ = new_n17269_ & new_n17290_;
  assign new_n17292_ = new_n17245_ & new_n17291_;
  assign new_n17293_ = new_n17199_ & new_n17292_;
  assign new_n17294_ = new_n17106_ & new_n17293_;
  assign new_n17295_ = new_n8689_ & new_n17251_;
  assign new_n17296_ = new_n8692_ & new_n17251_;
  assign new_n17297_ = new_n8694_ & new_n17251_;
  assign new_n17298_ = ~new_n17296_ & ~new_n17297_;
  assign new_n17299_ = ~new_n17295_ & new_n17298_;
  assign new_n17300_ = new_n5752_ & new_n15981_;
  assign new_n17301_ = new_n8845_ & new_n17300_;
  assign new_n17302_ = new_n8699_ & new_n17251_;
  assign new_n17303_ = new_n8701_ & new_n17251_;
  assign new_n17304_ = ~new_n17302_ & ~new_n17303_;
  assign new_n17305_ = ~new_n17301_ & new_n17304_;
  assign new_n17306_ = new_n17299_ & new_n17305_;
  assign new_n17307_ = new_n8851_ & new_n17300_;
  assign new_n17308_ = new_n8853_ & new_n17300_;
  assign new_n17309_ = new_n8855_ & new_n17300_;
  assign new_n17310_ = ~new_n17308_ & ~new_n17309_;
  assign new_n17311_ = ~new_n17307_ & new_n17310_;
  assign new_n17312_ = new_n8862_ & new_n17300_;
  assign new_n17313_ = new_n8864_ & new_n17300_;
  assign new_n17314_ = new_n8866_ & new_n17300_;
  assign new_n17315_ = ~new_n17313_ & ~new_n17314_;
  assign new_n17316_ = ~new_n17312_ & new_n17315_;
  assign new_n17317_ = new_n17311_ & new_n17316_;
  assign new_n17318_ = new_n17306_ & new_n17317_;
  assign new_n17319_ = new_n8870_ & new_n17300_;
  assign new_n17320_ = new_n8872_ & new_n17300_;
  assign new_n17321_ = new_n8874_ & new_n17300_;
  assign new_n17322_ = ~new_n17320_ & ~new_n17321_;
  assign new_n17323_ = ~new_n17319_ & new_n17322_;
  assign new_n17324_ = new_n8880_ & new_n17300_;
  assign new_n17325_ = new_n8882_ & new_n17300_;
  assign new_n17326_ = new_n8884_ & new_n17300_;
  assign new_n17327_ = ~new_n17325_ & ~new_n17326_;
  assign new_n17328_ = ~new_n17324_ & new_n17327_;
  assign new_n17329_ = new_n17323_ & new_n17328_;
  assign new_n17330_ = new_n8898_ & new_n17300_;
  assign new_n17331_ = new_n8888_ & new_n17300_;
  assign new_n17332_ = new_n8890_ & new_n17300_;
  assign new_n17333_ = ~new_n17331_ & ~new_n17332_;
  assign new_n17334_ = ~new_n17330_ & new_n17333_;
  assign new_n17335_ = new_n8900_ & new_n17300_;
  assign new_n17336_ = new_n8896_ & new_n17300_;
  assign new_n17337_ = ~new_n17335_ & ~new_n17336_;
  assign new_n17338_ = new_n17334_ & new_n17337_;
  assign new_n17339_ = new_n17329_ & new_n17338_;
  assign new_n17340_ = new_n17318_ & new_n17339_;
  assign new_n17341_ = new_n8905_ & new_n17300_;
  assign new_n17342_ = new_n8907_ & new_n17300_;
  assign new_n17343_ = new_n8909_ & new_n17300_;
  assign new_n17344_ = ~new_n17342_ & ~new_n17343_;
  assign new_n17345_ = ~new_n17341_ & new_n17344_;
  assign new_n17346_ = new_n8914_ & new_n17300_;
  assign new_n17347_ = new_n8916_ & new_n17300_;
  assign new_n17348_ = new_n8918_ & new_n17300_;
  assign new_n17349_ = ~new_n17347_ & ~new_n17348_;
  assign new_n17350_ = ~new_n17346_ & new_n17349_;
  assign new_n17351_ = new_n17345_ & new_n17350_;
  assign new_n17352_ = new_n8923_ & new_n17300_;
  assign new_n17353_ = new_n8925_ & new_n17300_;
  assign new_n17354_ = new_n8927_ & new_n17300_;
  assign new_n17355_ = ~new_n17353_ & ~new_n17354_;
  assign new_n17356_ = ~new_n17352_ & new_n17355_;
  assign new_n17357_ = new_n8934_ & new_n17300_;
  assign new_n17358_ = new_n8936_ & new_n17300_;
  assign new_n17359_ = new_n8938_ & new_n17300_;
  assign new_n17360_ = ~new_n17358_ & ~new_n17359_;
  assign new_n17361_ = ~new_n17357_ & new_n17360_;
  assign new_n17362_ = new_n17356_ & new_n17361_;
  assign new_n17363_ = new_n17351_ & new_n17362_;
  assign new_n17364_ = new_n5759_ & new_n16044_;
  assign new_n17365_ = new_n8617_ & new_n17364_;
  assign new_n17366_ = new_n8943_ & new_n17300_;
  assign new_n17367_ = new_n8945_ & new_n17300_;
  assign new_n17368_ = ~new_n17366_ & ~new_n17367_;
  assign new_n17369_ = ~new_n17365_ & new_n17368_;
  assign new_n17370_ = new_n8625_ & new_n17364_;
  assign new_n17371_ = new_n8628_ & new_n17364_;
  assign new_n17372_ = new_n8630_ & new_n17364_;
  assign new_n17373_ = ~new_n17371_ & ~new_n17372_;
  assign new_n17374_ = ~new_n17370_ & new_n17373_;
  assign new_n17375_ = new_n17369_ & new_n17374_;
  assign new_n17376_ = new_n8635_ & new_n17364_;
  assign new_n17377_ = new_n8637_ & new_n17364_;
  assign new_n17378_ = new_n8639_ & new_n17364_;
  assign new_n17379_ = ~new_n17377_ & ~new_n17378_;
  assign new_n17380_ = ~new_n17376_ & new_n17379_;
  assign new_n17381_ = new_n8648_ & new_n17364_;
  assign new_n17382_ = new_n8650_ & new_n17364_;
  assign new_n17383_ = ~new_n17381_ & ~new_n17382_;
  assign new_n17384_ = new_n17380_ & new_n17383_;
  assign new_n17385_ = new_n17375_ & new_n17384_;
  assign new_n17386_ = new_n17363_ & new_n17385_;
  assign new_n17387_ = new_n17340_ & new_n17386_;
  assign new_n17388_ = new_n8659_ & new_n17364_;
  assign new_n17389_ = new_n8646_ & new_n17364_;
  assign new_n17390_ = new_n8657_ & new_n17364_;
  assign new_n17391_ = ~new_n17389_ & ~new_n17390_;
  assign new_n17392_ = ~new_n17388_ & new_n17391_;
  assign new_n17393_ = new_n8670_ & new_n17364_;
  assign new_n17394_ = new_n8655_ & new_n17364_;
  assign new_n17395_ = new_n8667_ & new_n17364_;
  assign new_n17396_ = ~new_n17394_ & ~new_n17395_;
  assign new_n17397_ = ~new_n17393_ & new_n17396_;
  assign new_n17398_ = new_n17392_ & new_n17397_;
  assign new_n17399_ = new_n8681_ & new_n17364_;
  assign new_n17400_ = new_n8665_ & new_n17364_;
  assign new_n17401_ = new_n8678_ & new_n17364_;
  assign new_n17402_ = ~new_n17400_ & ~new_n17401_;
  assign new_n17403_ = ~new_n17399_ & new_n17402_;
  assign new_n17404_ = new_n8694_ & new_n17364_;
  assign new_n17405_ = new_n8675_ & new_n17364_;
  assign new_n17406_ = new_n8692_ & new_n17364_;
  assign new_n17407_ = ~new_n17405_ & ~new_n17406_;
  assign new_n17408_ = ~new_n17404_ & new_n17407_;
  assign new_n17409_ = new_n17403_ & new_n17408_;
  assign new_n17410_ = new_n17398_ & new_n17409_;
  assign new_n17411_ = new_n8701_ & new_n17364_;
  assign new_n17412_ = new_n8689_ & new_n17364_;
  assign new_n17413_ = new_n8699_ & new_n17364_;
  assign new_n17414_ = ~new_n17412_ & ~new_n17413_;
  assign new_n17415_ = ~new_n17411_ & new_n17414_;
  assign new_n17416_ = new_n5759_ & new_n16093_;
  assign new_n17417_ = new_n8630_ & new_n17416_;
  assign new_n17418_ = new_n8617_ & new_n17416_;
  assign new_n17419_ = new_n8628_ & new_n17416_;
  assign new_n17420_ = ~new_n17418_ & ~new_n17419_;
  assign new_n17421_ = ~new_n17417_ & new_n17420_;
  assign new_n17422_ = new_n17415_ & new_n17421_;
  assign new_n17423_ = new_n8639_ & new_n17416_;
  assign new_n17424_ = new_n8625_ & new_n17416_;
  assign new_n17425_ = new_n8637_ & new_n17416_;
  assign new_n17426_ = ~new_n17424_ & ~new_n17425_;
  assign new_n17427_ = ~new_n17423_ & new_n17426_;
  assign new_n17428_ = new_n8635_ & new_n17416_;
  assign new_n17429_ = new_n8648_ & new_n17416_;
  assign new_n17430_ = ~new_n17428_ & ~new_n17429_;
  assign new_n17431_ = new_n17427_ & new_n17430_;
  assign new_n17432_ = new_n17422_ & new_n17431_;
  assign new_n17433_ = new_n17410_ & new_n17432_;
  assign new_n17434_ = new_n8657_ & new_n17416_;
  assign new_n17435_ = new_n8650_ & new_n17416_;
  assign new_n17436_ = new_n8646_ & new_n17416_;
  assign new_n17437_ = ~new_n17435_ & ~new_n17436_;
  assign new_n17438_ = ~new_n17434_ & new_n17437_;
  assign new_n17439_ = new_n8667_ & new_n17416_;
  assign new_n17440_ = new_n8659_ & new_n17416_;
  assign new_n17441_ = new_n8655_ & new_n17416_;
  assign new_n17442_ = ~new_n17440_ & ~new_n17441_;
  assign new_n17443_ = ~new_n17439_ & new_n17442_;
  assign new_n17444_ = new_n17438_ & new_n17443_;
  assign new_n17445_ = new_n8678_ & new_n17416_;
  assign new_n17446_ = new_n8670_ & new_n17416_;
  assign new_n17447_ = new_n8665_ & new_n17416_;
  assign new_n17448_ = ~new_n17446_ & ~new_n17447_;
  assign new_n17449_ = ~new_n17445_ & new_n17448_;
  assign new_n17450_ = new_n8692_ & new_n17416_;
  assign new_n17451_ = new_n8681_ & new_n17416_;
  assign new_n17452_ = new_n8675_ & new_n17416_;
  assign new_n17453_ = ~new_n17451_ & ~new_n17452_;
  assign new_n17454_ = ~new_n17450_ & new_n17453_;
  assign new_n17455_ = new_n17449_ & new_n17454_;
  assign new_n17456_ = new_n17444_ & new_n17455_;
  assign new_n17457_ = new_n8699_ & new_n17416_;
  assign new_n17458_ = new_n8694_ & new_n17416_;
  assign new_n17459_ = new_n8689_ & new_n17416_;
  assign new_n17460_ = ~new_n17458_ & ~new_n17459_;
  assign new_n17461_ = ~new_n17457_ & new_n17460_;
  assign new_n17462_ = new_n5759_ & new_n16151_;
  assign new_n17463_ = new_n8628_ & new_n17462_;
  assign new_n17464_ = new_n8701_ & new_n17416_;
  assign new_n17465_ = new_n8617_ & new_n17462_;
  assign new_n17466_ = ~new_n17464_ & ~new_n17465_;
  assign new_n17467_ = ~new_n17463_ & new_n17466_;
  assign new_n17468_ = new_n17461_ & new_n17467_;
  assign new_n17469_ = new_n8637_ & new_n17462_;
  assign new_n17470_ = new_n8630_ & new_n17462_;
  assign new_n17471_ = new_n8625_ & new_n17462_;
  assign new_n17472_ = ~new_n17470_ & ~new_n17471_;
  assign new_n17473_ = ~new_n17469_ & new_n17472_;
  assign new_n17474_ = new_n8639_ & new_n17462_;
  assign new_n17475_ = new_n8635_ & new_n17462_;
  assign new_n17476_ = ~new_n17474_ & ~new_n17475_;
  assign new_n17477_ = new_n17473_ & new_n17476_;
  assign new_n17478_ = new_n17468_ & new_n17477_;
  assign new_n17479_ = new_n17456_ & new_n17478_;
  assign new_n17480_ = new_n17433_ & new_n17479_;
  assign new_n17481_ = new_n17387_ & new_n17480_;
  assign new_n17482_ = new_n8646_ & new_n17462_;
  assign new_n17483_ = new_n8648_ & new_n17462_;
  assign new_n17484_ = new_n8650_ & new_n17462_;
  assign new_n17485_ = ~new_n17483_ & ~new_n17484_;
  assign new_n17486_ = ~new_n17482_ & new_n17485_;
  assign new_n17487_ = new_n8655_ & new_n17462_;
  assign new_n17488_ = new_n8657_ & new_n17462_;
  assign new_n17489_ = new_n8659_ & new_n17462_;
  assign new_n17490_ = ~new_n17488_ & ~new_n17489_;
  assign new_n17491_ = ~new_n17487_ & new_n17490_;
  assign new_n17492_ = new_n17486_ & new_n17491_;
  assign new_n17493_ = new_n8665_ & new_n17462_;
  assign new_n17494_ = new_n8667_ & new_n17462_;
  assign new_n17495_ = new_n8670_ & new_n17462_;
  assign new_n17496_ = ~new_n17494_ & ~new_n17495_;
  assign new_n17497_ = ~new_n17493_ & new_n17496_;
  assign new_n17498_ = new_n8675_ & new_n17462_;
  assign new_n17499_ = new_n8678_ & new_n17462_;
  assign new_n17500_ = new_n8681_ & new_n17462_;
  assign new_n17501_ = ~new_n17499_ & ~new_n17500_;
  assign new_n17502_ = ~new_n17498_ & new_n17501_;
  assign new_n17503_ = new_n17497_ & new_n17502_;
  assign new_n17504_ = new_n17492_ & new_n17503_;
  assign new_n17505_ = new_n8689_ & new_n17462_;
  assign new_n17506_ = new_n8692_ & new_n17462_;
  assign new_n17507_ = new_n8694_ & new_n17462_;
  assign new_n17508_ = ~new_n17506_ & ~new_n17507_;
  assign new_n17509_ = ~new_n17505_ & new_n17508_;
  assign new_n17510_ = new_n5759_ & new_n16200_;
  assign new_n17511_ = new_n8617_ & new_n17510_;
  assign new_n17512_ = new_n8699_ & new_n17462_;
  assign new_n17513_ = new_n8701_ & new_n17462_;
  assign new_n17514_ = ~new_n17512_ & ~new_n17513_;
  assign new_n17515_ = ~new_n17511_ & new_n17514_;
  assign new_n17516_ = new_n17509_ & new_n17515_;
  assign new_n17517_ = new_n8625_ & new_n17510_;
  assign new_n17518_ = new_n8628_ & new_n17510_;
  assign new_n17519_ = new_n8630_ & new_n17510_;
  assign new_n17520_ = ~new_n17518_ & ~new_n17519_;
  assign new_n17521_ = ~new_n17517_ & new_n17520_;
  assign new_n17522_ = new_n8637_ & new_n17510_;
  assign new_n17523_ = new_n8639_ & new_n17510_;
  assign new_n17524_ = ~new_n17522_ & ~new_n17523_;
  assign new_n17525_ = new_n17521_ & new_n17524_;
  assign new_n17526_ = new_n17516_ & new_n17525_;
  assign new_n17527_ = new_n17504_ & new_n17526_;
  assign new_n17528_ = new_n8650_ & new_n17510_;
  assign new_n17529_ = new_n8635_ & new_n17510_;
  assign new_n17530_ = new_n8648_ & new_n17510_;
  assign new_n17531_ = ~new_n17529_ & ~new_n17530_;
  assign new_n17532_ = ~new_n17528_ & new_n17531_;
  assign new_n17533_ = new_n8659_ & new_n17510_;
  assign new_n17534_ = new_n8646_ & new_n17510_;
  assign new_n17535_ = new_n8657_ & new_n17510_;
  assign new_n17536_ = ~new_n17534_ & ~new_n17535_;
  assign new_n17537_ = ~new_n17533_ & new_n17536_;
  assign new_n17538_ = new_n17532_ & new_n17537_;
  assign new_n17539_ = new_n8670_ & new_n17510_;
  assign new_n17540_ = new_n8655_ & new_n17510_;
  assign new_n17541_ = new_n8667_ & new_n17510_;
  assign new_n17542_ = ~new_n17540_ & ~new_n17541_;
  assign new_n17543_ = ~new_n17539_ & new_n17542_;
  assign new_n17544_ = new_n8681_ & new_n17510_;
  assign new_n17545_ = new_n8665_ & new_n17510_;
  assign new_n17546_ = new_n8678_ & new_n17510_;
  assign new_n17547_ = ~new_n17545_ & ~new_n17546_;
  assign new_n17548_ = ~new_n17544_ & new_n17547_;
  assign new_n17549_ = new_n17543_ & new_n17548_;
  assign new_n17550_ = new_n17538_ & new_n17549_;
  assign new_n17551_ = new_n8694_ & new_n17510_;
  assign new_n17552_ = new_n8675_ & new_n17510_;
  assign new_n17553_ = new_n8692_ & new_n17510_;
  assign new_n17554_ = ~new_n17552_ & ~new_n17553_;
  assign new_n17555_ = ~new_n17551_ & new_n17554_;
  assign new_n17556_ = new_n8701_ & new_n17510_;
  assign new_n17557_ = new_n8689_ & new_n17510_;
  assign new_n17558_ = new_n8699_ & new_n17510_;
  assign new_n17559_ = ~new_n17557_ & ~new_n17558_;
  assign new_n17560_ = ~new_n17556_ & new_n17559_;
  assign new_n17561_ = new_n17555_ & new_n17560_;
  assign new_n17562_ = new_n5759_ & new_n16248_;
  assign new_n17563_ = new_n8855_ & new_n17562_;
  assign new_n17564_ = new_n8845_ & new_n17562_;
  assign new_n17565_ = new_n8853_ & new_n17562_;
  assign new_n17566_ = ~new_n17564_ & ~new_n17565_;
  assign new_n17567_ = ~new_n17563_ & new_n17566_;
  assign new_n17568_ = new_n8851_ & new_n17562_;
  assign new_n17569_ = new_n8864_ & new_n17562_;
  assign new_n17570_ = ~new_n17568_ & ~new_n17569_;
  assign new_n17571_ = new_n17567_ & new_n17570_;
  assign new_n17572_ = new_n17561_ & new_n17571_;
  assign new_n17573_ = new_n17550_ & new_n17572_;
  assign new_n17574_ = new_n17527_ & new_n17573_;
  assign new_n17575_ = new_n8872_ & new_n17562_;
  assign new_n17576_ = new_n8866_ & new_n17562_;
  assign new_n17577_ = new_n8862_ & new_n17562_;
  assign new_n17578_ = ~new_n17576_ & ~new_n17577_;
  assign new_n17579_ = ~new_n17575_ & new_n17578_;
  assign new_n17580_ = new_n8882_ & new_n17562_;
  assign new_n17581_ = new_n8874_ & new_n17562_;
  assign new_n17582_ = new_n8870_ & new_n17562_;
  assign new_n17583_ = ~new_n17581_ & ~new_n17582_;
  assign new_n17584_ = ~new_n17580_ & new_n17583_;
  assign new_n17585_ = new_n17579_ & new_n17584_;
  assign new_n17586_ = new_n8888_ & new_n17562_;
  assign new_n17587_ = new_n8884_ & new_n17562_;
  assign new_n17588_ = new_n8880_ & new_n17562_;
  assign new_n17589_ = ~new_n17587_ & ~new_n17588_;
  assign new_n17590_ = ~new_n17586_ & new_n17589_;
  assign new_n17591_ = new_n8900_ & new_n17562_;
  assign new_n17592_ = new_n8890_ & new_n17562_;
  assign new_n17593_ = new_n8898_ & new_n17562_;
  assign new_n17594_ = ~new_n17592_ & ~new_n17593_;
  assign new_n17595_ = ~new_n17591_ & new_n17594_;
  assign new_n17596_ = new_n17590_ & new_n17595_;
  assign new_n17597_ = new_n17585_ & new_n17596_;
  assign new_n17598_ = new_n8909_ & new_n17562_;
  assign new_n17599_ = new_n8896_ & new_n17562_;
  assign new_n17600_ = new_n8907_ & new_n17562_;
  assign new_n17601_ = ~new_n17599_ & ~new_n17600_;
  assign new_n17602_ = ~new_n17598_ & new_n17601_;
  assign new_n17603_ = new_n8918_ & new_n17562_;
  assign new_n17604_ = new_n8905_ & new_n17562_;
  assign new_n17605_ = new_n8916_ & new_n17562_;
  assign new_n17606_ = ~new_n17604_ & ~new_n17605_;
  assign new_n17607_ = ~new_n17603_ & new_n17606_;
  assign new_n17608_ = new_n17602_ & new_n17607_;
  assign new_n17609_ = new_n8927_ & new_n17562_;
  assign new_n17610_ = new_n8914_ & new_n17562_;
  assign new_n17611_ = new_n8925_ & new_n17562_;
  assign new_n17612_ = ~new_n17610_ & ~new_n17611_;
  assign new_n17613_ = ~new_n17609_ & new_n17612_;
  assign new_n17614_ = new_n8923_ & new_n17562_;
  assign new_n17615_ = new_n8936_ & new_n17562_;
  assign new_n17616_ = ~new_n17614_ & ~new_n17615_;
  assign new_n17617_ = new_n17613_ & new_n17616_;
  assign new_n17618_ = new_n17608_ & new_n17617_;
  assign new_n17619_ = new_n17597_ & new_n17618_;
  assign new_n17620_ = new_n8943_ & new_n17562_;
  assign new_n17621_ = new_n8938_ & new_n17562_;
  assign new_n17622_ = new_n8934_ & new_n17562_;
  assign new_n17623_ = ~new_n17621_ & ~new_n17622_;
  assign new_n17624_ = ~new_n17620_ & new_n17623_;
  assign new_n17625_ = new_n5768_ & new_n16311_;
  assign new_n17626_ = new_n8628_ & new_n17625_;
  assign new_n17627_ = new_n8945_ & new_n17562_;
  assign new_n17628_ = new_n8617_ & new_n17625_;
  assign new_n17629_ = ~new_n17627_ & ~new_n17628_;
  assign new_n17630_ = ~new_n17626_ & new_n17629_;
  assign new_n17631_ = new_n17624_ & new_n17630_;
  assign new_n17632_ = new_n8637_ & new_n17625_;
  assign new_n17633_ = new_n8630_ & new_n17625_;
  assign new_n17634_ = new_n8625_ & new_n17625_;
  assign new_n17635_ = ~new_n17633_ & ~new_n17634_;
  assign new_n17636_ = ~new_n17632_ & new_n17635_;
  assign new_n17637_ = new_n8648_ & new_n17625_;
  assign new_n17638_ = new_n8639_ & new_n17625_;
  assign new_n17639_ = new_n8635_ & new_n17625_;
  assign new_n17640_ = ~new_n17638_ & ~new_n17639_;
  assign new_n17641_ = ~new_n17637_ & new_n17640_;
  assign new_n17642_ = new_n17636_ & new_n17641_;
  assign new_n17643_ = new_n17631_ & new_n17642_;
  assign new_n17644_ = new_n8657_ & new_n17625_;
  assign new_n17645_ = new_n8650_ & new_n17625_;
  assign new_n17646_ = new_n8646_ & new_n17625_;
  assign new_n17647_ = ~new_n17645_ & ~new_n17646_;
  assign new_n17648_ = ~new_n17644_ & new_n17647_;
  assign new_n17649_ = new_n8667_ & new_n17625_;
  assign new_n17650_ = new_n8659_ & new_n17625_;
  assign new_n17651_ = new_n8655_ & new_n17625_;
  assign new_n17652_ = ~new_n17650_ & ~new_n17651_;
  assign new_n17653_ = ~new_n17649_ & new_n17652_;
  assign new_n17654_ = new_n17648_ & new_n17653_;
  assign new_n17655_ = new_n8678_ & new_n17625_;
  assign new_n17656_ = new_n8670_ & new_n17625_;
  assign new_n17657_ = new_n8665_ & new_n17625_;
  assign new_n17658_ = ~new_n17656_ & ~new_n17657_;
  assign new_n17659_ = ~new_n17655_ & new_n17658_;
  assign new_n17660_ = new_n8681_ & new_n17625_;
  assign new_n17661_ = new_n8675_ & new_n17625_;
  assign new_n17662_ = ~new_n17660_ & ~new_n17661_;
  assign new_n17663_ = new_n17659_ & new_n17662_;
  assign new_n17664_ = new_n17654_ & new_n17663_;
  assign new_n17665_ = new_n17643_ & new_n17664_;
  assign new_n17666_ = new_n17619_ & new_n17665_;
  assign new_n17667_ = new_n17574_ & new_n17666_;
  assign new_n17668_ = new_n17481_ & new_n17667_;
  assign new_n17669_ = new_n17294_ & new_n17668_;
  assign new_n17670_ = new_n16919_ & new_n17669_;
  assign new_n17671_ = new_n8689_ & new_n17625_;
  assign new_n17672_ = new_n8692_ & new_n17625_;
  assign new_n17673_ = new_n8694_ & new_n17625_;
  assign new_n17674_ = ~new_n17672_ & ~new_n17673_;
  assign new_n17675_ = ~new_n17671_ & new_n17674_;
  assign new_n17676_ = new_n5768_ & new_n16360_;
  assign new_n17677_ = new_n8617_ & new_n17676_;
  assign new_n17678_ = new_n8699_ & new_n17625_;
  assign new_n17679_ = new_n8701_ & new_n17625_;
  assign new_n17680_ = ~new_n17678_ & ~new_n17679_;
  assign new_n17681_ = ~new_n17677_ & new_n17680_;
  assign new_n17682_ = new_n17675_ & new_n17681_;
  assign new_n17683_ = new_n8625_ & new_n17676_;
  assign new_n17684_ = new_n8628_ & new_n17676_;
  assign new_n17685_ = new_n8630_ & new_n17676_;
  assign new_n17686_ = ~new_n17684_ & ~new_n17685_;
  assign new_n17687_ = ~new_n17683_ & new_n17686_;
  assign new_n17688_ = new_n8635_ & new_n17676_;
  assign new_n17689_ = new_n8637_ & new_n17676_;
  assign new_n17690_ = new_n8639_ & new_n17676_;
  assign new_n17691_ = ~new_n17689_ & ~new_n17690_;
  assign new_n17692_ = ~new_n17688_ & new_n17691_;
  assign new_n17693_ = new_n17687_ & new_n17692_;
  assign new_n17694_ = new_n17682_ & new_n17693_;
  assign new_n17695_ = new_n8646_ & new_n17676_;
  assign new_n17696_ = new_n8648_ & new_n17676_;
  assign new_n17697_ = new_n8650_ & new_n17676_;
  assign new_n17698_ = ~new_n17696_ & ~new_n17697_;
  assign new_n17699_ = ~new_n17695_ & new_n17698_;
  assign new_n17700_ = new_n8655_ & new_n17676_;
  assign new_n17701_ = new_n8657_ & new_n17676_;
  assign new_n17702_ = new_n8659_ & new_n17676_;
  assign new_n17703_ = ~new_n17701_ & ~new_n17702_;
  assign new_n17704_ = ~new_n17700_ & new_n17703_;
  assign new_n17705_ = new_n17699_ & new_n17704_;
  assign new_n17706_ = new_n8665_ & new_n17676_;
  assign new_n17707_ = new_n8667_ & new_n17676_;
  assign new_n17708_ = new_n8670_ & new_n17676_;
  assign new_n17709_ = ~new_n17707_ & ~new_n17708_;
  assign new_n17710_ = ~new_n17706_ & new_n17709_;
  assign new_n17711_ = new_n8675_ & new_n17676_;
  assign new_n17712_ = new_n8678_ & new_n17676_;
  assign new_n17713_ = new_n8681_ & new_n17676_;
  assign new_n17714_ = ~new_n17712_ & ~new_n17713_;
  assign new_n17715_ = ~new_n17711_ & new_n17714_;
  assign new_n17716_ = new_n17710_ & new_n17715_;
  assign new_n17717_ = new_n17705_ & new_n17716_;
  assign new_n17718_ = new_n17694_ & new_n17717_;
  assign new_n17719_ = new_n8689_ & new_n17676_;
  assign new_n17720_ = new_n8692_ & new_n17676_;
  assign new_n17721_ = new_n8694_ & new_n17676_;
  assign new_n17722_ = ~new_n17720_ & ~new_n17721_;
  assign new_n17723_ = ~new_n17719_ & new_n17722_;
  assign new_n17724_ = new_n5768_ & new_n16414_;
  assign new_n17725_ = new_n8617_ & new_n17724_;
  assign new_n17726_ = new_n8699_ & new_n17676_;
  assign new_n17727_ = new_n8701_ & new_n17676_;
  assign new_n17728_ = ~new_n17726_ & ~new_n17727_;
  assign new_n17729_ = ~new_n17725_ & new_n17728_;
  assign new_n17730_ = new_n17723_ & new_n17729_;
  assign new_n17731_ = new_n8625_ & new_n17724_;
  assign new_n17732_ = new_n8628_ & new_n17724_;
  assign new_n17733_ = new_n8630_ & new_n17724_;
  assign new_n17734_ = ~new_n17732_ & ~new_n17733_;
  assign new_n17735_ = ~new_n17731_ & new_n17734_;
  assign new_n17736_ = new_n8635_ & new_n17724_;
  assign new_n17737_ = new_n8637_ & new_n17724_;
  assign new_n17738_ = new_n8639_ & new_n17724_;
  assign new_n17739_ = ~new_n17737_ & ~new_n17738_;
  assign new_n17740_ = ~new_n17736_ & new_n17739_;
  assign new_n17741_ = new_n17735_ & new_n17740_;
  assign new_n17742_ = new_n17730_ & new_n17741_;
  assign new_n17743_ = new_n8646_ & new_n17724_;
  assign new_n17744_ = new_n8648_ & new_n17724_;
  assign new_n17745_ = new_n8650_ & new_n17724_;
  assign new_n17746_ = ~new_n17744_ & ~new_n17745_;
  assign new_n17747_ = ~new_n17743_ & new_n17746_;
  assign new_n17748_ = new_n8655_ & new_n17724_;
  assign new_n17749_ = new_n8657_ & new_n17724_;
  assign new_n17750_ = new_n8659_ & new_n17724_;
  assign new_n17751_ = ~new_n17749_ & ~new_n17750_;
  assign new_n17752_ = ~new_n17748_ & new_n17751_;
  assign new_n17753_ = new_n17747_ & new_n17752_;
  assign new_n17754_ = new_n8665_ & new_n17724_;
  assign new_n17755_ = new_n8667_ & new_n17724_;
  assign new_n17756_ = new_n8670_ & new_n17724_;
  assign new_n17757_ = ~new_n17755_ & ~new_n17756_;
  assign new_n17758_ = ~new_n17754_ & new_n17757_;
  assign new_n17759_ = new_n8678_ & new_n17724_;
  assign new_n17760_ = new_n8681_ & new_n17724_;
  assign new_n17761_ = ~new_n17759_ & ~new_n17760_;
  assign new_n17762_ = new_n17758_ & new_n17761_;
  assign new_n17763_ = new_n17753_ & new_n17762_;
  assign new_n17764_ = new_n17742_ & new_n17763_;
  assign new_n17765_ = new_n17718_ & new_n17764_;
  assign new_n17766_ = new_n8694_ & new_n17724_;
  assign new_n17767_ = new_n8675_ & new_n17724_;
  assign new_n17768_ = new_n8692_ & new_n17724_;
  assign new_n17769_ = ~new_n17767_ & ~new_n17768_;
  assign new_n17770_ = ~new_n17766_ & new_n17769_;
  assign new_n17771_ = new_n8701_ & new_n17724_;
  assign new_n17772_ = new_n8689_ & new_n17724_;
  assign new_n17773_ = new_n8699_ & new_n17724_;
  assign new_n17774_ = ~new_n17772_ & ~new_n17773_;
  assign new_n17775_ = ~new_n17771_ & new_n17774_;
  assign new_n17776_ = new_n17770_ & new_n17775_;
  assign new_n17777_ = new_n5768_ & new_n16462_;
  assign new_n17778_ = new_n8630_ & new_n17777_;
  assign new_n17779_ = new_n8617_ & new_n17777_;
  assign new_n17780_ = new_n8628_ & new_n17777_;
  assign new_n17781_ = ~new_n17779_ & ~new_n17780_;
  assign new_n17782_ = ~new_n17778_ & new_n17781_;
  assign new_n17783_ = new_n8639_ & new_n17777_;
  assign new_n17784_ = new_n8625_ & new_n17777_;
  assign new_n17785_ = new_n8637_ & new_n17777_;
  assign new_n17786_ = ~new_n17784_ & ~new_n17785_;
  assign new_n17787_ = ~new_n17783_ & new_n17786_;
  assign new_n17788_ = new_n17782_ & new_n17787_;
  assign new_n17789_ = new_n17776_ & new_n17788_;
  assign new_n17790_ = new_n8650_ & new_n17777_;
  assign new_n17791_ = new_n8635_ & new_n17777_;
  assign new_n17792_ = new_n8648_ & new_n17777_;
  assign new_n17793_ = ~new_n17791_ & ~new_n17792_;
  assign new_n17794_ = ~new_n17790_ & new_n17793_;
  assign new_n17795_ = new_n8659_ & new_n17777_;
  assign new_n17796_ = new_n8646_ & new_n17777_;
  assign new_n17797_ = new_n8657_ & new_n17777_;
  assign new_n17798_ = ~new_n17796_ & ~new_n17797_;
  assign new_n17799_ = ~new_n17795_ & new_n17798_;
  assign new_n17800_ = new_n17794_ & new_n17799_;
  assign new_n17801_ = new_n8670_ & new_n17777_;
  assign new_n17802_ = new_n8655_ & new_n17777_;
  assign new_n17803_ = new_n8667_ & new_n17777_;
  assign new_n17804_ = ~new_n17802_ & ~new_n17803_;
  assign new_n17805_ = ~new_n17801_ & new_n17804_;
  assign new_n17806_ = new_n8665_ & new_n17777_;
  assign new_n17807_ = new_n8678_ & new_n17777_;
  assign new_n17808_ = ~new_n17806_ & ~new_n17807_;
  assign new_n17809_ = new_n17805_ & new_n17808_;
  assign new_n17810_ = new_n17800_ & new_n17809_;
  assign new_n17811_ = new_n17789_ & new_n17810_;
  assign new_n17812_ = new_n8692_ & new_n17777_;
  assign new_n17813_ = new_n8681_ & new_n17777_;
  assign new_n17814_ = new_n8675_ & new_n17777_;
  assign new_n17815_ = ~new_n17813_ & ~new_n17814_;
  assign new_n17816_ = ~new_n17812_ & new_n17815_;
  assign new_n17817_ = new_n8699_ & new_n17777_;
  assign new_n17818_ = new_n8694_ & new_n17777_;
  assign new_n17819_ = new_n8689_ & new_n17777_;
  assign new_n17820_ = ~new_n17818_ & ~new_n17819_;
  assign new_n17821_ = ~new_n17817_ & new_n17820_;
  assign new_n17822_ = new_n17816_ & new_n17821_;
  assign new_n17823_ = new_n5768_ & new_n16509_;
  assign new_n17824_ = new_n8853_ & new_n17823_;
  assign new_n17825_ = new_n8701_ & new_n17777_;
  assign new_n17826_ = new_n8845_ & new_n17823_;
  assign new_n17827_ = ~new_n17825_ & ~new_n17826_;
  assign new_n17828_ = ~new_n17824_ & new_n17827_;
  assign new_n17829_ = new_n8864_ & new_n17823_;
  assign new_n17830_ = new_n8855_ & new_n17823_;
  assign new_n17831_ = new_n8851_ & new_n17823_;
  assign new_n17832_ = ~new_n17830_ & ~new_n17831_;
  assign new_n17833_ = ~new_n17829_ & new_n17832_;
  assign new_n17834_ = new_n17828_ & new_n17833_;
  assign new_n17835_ = new_n17822_ & new_n17834_;
  assign new_n17836_ = new_n8872_ & new_n17823_;
  assign new_n17837_ = new_n8866_ & new_n17823_;
  assign new_n17838_ = new_n8862_ & new_n17823_;
  assign new_n17839_ = ~new_n17837_ & ~new_n17838_;
  assign new_n17840_ = ~new_n17836_ & new_n17839_;
  assign new_n17841_ = new_n8882_ & new_n17823_;
  assign new_n17842_ = new_n8874_ & new_n17823_;
  assign new_n17843_ = new_n8870_ & new_n17823_;
  assign new_n17844_ = ~new_n17842_ & ~new_n17843_;
  assign new_n17845_ = ~new_n17841_ & new_n17844_;
  assign new_n17846_ = new_n17840_ & new_n17845_;
  assign new_n17847_ = new_n8888_ & new_n17823_;
  assign new_n17848_ = new_n8884_ & new_n17823_;
  assign new_n17849_ = new_n8880_ & new_n17823_;
  assign new_n17850_ = ~new_n17848_ & ~new_n17849_;
  assign new_n17851_ = ~new_n17847_ & new_n17850_;
  assign new_n17852_ = new_n8890_ & new_n17823_;
  assign new_n17853_ = new_n8898_ & new_n17823_;
  assign new_n17854_ = ~new_n17852_ & ~new_n17853_;
  assign new_n17855_ = new_n17851_ & new_n17854_;
  assign new_n17856_ = new_n17846_ & new_n17855_;
  assign new_n17857_ = new_n17835_ & new_n17856_;
  assign new_n17858_ = new_n17811_ & new_n17857_;
  assign new_n17859_ = new_n17765_ & new_n17858_;
  assign new_n17860_ = new_n8907_ & new_n17823_;
  assign new_n17861_ = new_n8900_ & new_n17823_;
  assign new_n17862_ = new_n8896_ & new_n17823_;
  assign new_n17863_ = ~new_n17861_ & ~new_n17862_;
  assign new_n17864_ = ~new_n17860_ & new_n17863_;
  assign new_n17865_ = new_n8916_ & new_n17823_;
  assign new_n17866_ = new_n8909_ & new_n17823_;
  assign new_n17867_ = new_n8905_ & new_n17823_;
  assign new_n17868_ = ~new_n17866_ & ~new_n17867_;
  assign new_n17869_ = ~new_n17865_ & new_n17868_;
  assign new_n17870_ = new_n17864_ & new_n17869_;
  assign new_n17871_ = new_n8925_ & new_n17823_;
  assign new_n17872_ = new_n8918_ & new_n17823_;
  assign new_n17873_ = new_n8914_ & new_n17823_;
  assign new_n17874_ = ~new_n17872_ & ~new_n17873_;
  assign new_n17875_ = ~new_n17871_ & new_n17874_;
  assign new_n17876_ = new_n8936_ & new_n17823_;
  assign new_n17877_ = new_n8927_ & new_n17823_;
  assign new_n17878_ = new_n8923_ & new_n17823_;
  assign new_n17879_ = ~new_n17877_ & ~new_n17878_;
  assign new_n17880_ = ~new_n17876_ & new_n17879_;
  assign new_n17881_ = new_n17875_ & new_n17880_;
  assign new_n17882_ = new_n17870_ & new_n17881_;
  assign new_n17883_ = new_n8943_ & new_n17823_;
  assign new_n17884_ = new_n8938_ & new_n17823_;
  assign new_n17885_ = new_n8934_ & new_n17823_;
  assign new_n17886_ = ~new_n17884_ & ~new_n17885_;
  assign new_n17887_ = ~new_n17883_ & new_n17886_;
  assign new_n17888_ = new_n5768_ & new_n16575_;
  assign new_n17889_ = new_n8628_ & new_n17888_;
  assign new_n17890_ = new_n8945_ & new_n17823_;
  assign new_n17891_ = new_n8617_ & new_n17888_;
  assign new_n17892_ = ~new_n17890_ & ~new_n17891_;
  assign new_n17893_ = ~new_n17889_ & new_n17892_;
  assign new_n17894_ = new_n17887_ & new_n17893_;
  assign new_n17895_ = new_n8637_ & new_n17888_;
  assign new_n17896_ = new_n8630_ & new_n17888_;
  assign new_n17897_ = new_n8625_ & new_n17888_;
  assign new_n17898_ = ~new_n17896_ & ~new_n17897_;
  assign new_n17899_ = ~new_n17895_ & new_n17898_;
  assign new_n17900_ = new_n8639_ & new_n17888_;
  assign new_n17901_ = new_n8635_ & new_n17888_;
  assign new_n17902_ = ~new_n17900_ & ~new_n17901_;
  assign new_n17903_ = new_n17899_ & new_n17902_;
  assign new_n17904_ = new_n17894_ & new_n17903_;
  assign new_n17905_ = new_n17882_ & new_n17904_;
  assign new_n17906_ = new_n8646_ & new_n17888_;
  assign new_n17907_ = new_n8648_ & new_n17888_;
  assign new_n17908_ = new_n8650_ & new_n17888_;
  assign new_n17909_ = ~new_n17907_ & ~new_n17908_;
  assign new_n17910_ = ~new_n17906_ & new_n17909_;
  assign new_n17911_ = new_n8655_ & new_n17888_;
  assign new_n17912_ = new_n8657_ & new_n17888_;
  assign new_n17913_ = new_n8659_ & new_n17888_;
  assign new_n17914_ = ~new_n17912_ & ~new_n17913_;
  assign new_n17915_ = ~new_n17911_ & new_n17914_;
  assign new_n17916_ = new_n17910_ & new_n17915_;
  assign new_n17917_ = new_n8665_ & new_n17888_;
  assign new_n17918_ = new_n8667_ & new_n17888_;
  assign new_n17919_ = new_n8670_ & new_n17888_;
  assign new_n17920_ = ~new_n17918_ & ~new_n17919_;
  assign new_n17921_ = ~new_n17917_ & new_n17920_;
  assign new_n17922_ = new_n8675_ & new_n17888_;
  assign new_n17923_ = new_n8678_ & new_n17888_;
  assign new_n17924_ = new_n8681_ & new_n17888_;
  assign new_n17925_ = ~new_n17923_ & ~new_n17924_;
  assign new_n17926_ = ~new_n17922_ & new_n17925_;
  assign new_n17927_ = new_n17921_ & new_n17926_;
  assign new_n17928_ = new_n17916_ & new_n17927_;
  assign new_n17929_ = new_n8689_ & new_n17888_;
  assign new_n17930_ = new_n8692_ & new_n17888_;
  assign new_n17931_ = new_n8694_ & new_n17888_;
  assign new_n17932_ = ~new_n17930_ & ~new_n17931_;
  assign new_n17933_ = ~new_n17929_ & new_n17932_;
  assign new_n17934_ = new_n5768_ & new_n16631_;
  assign new_n17935_ = new_n8617_ & new_n17934_;
  assign new_n17936_ = new_n8699_ & new_n17888_;
  assign new_n17937_ = new_n8701_ & new_n17888_;
  assign new_n17938_ = ~new_n17936_ & ~new_n17937_;
  assign new_n17939_ = ~new_n17935_ & new_n17938_;
  assign new_n17940_ = new_n17933_ & new_n17939_;
  assign new_n17941_ = new_n8625_ & new_n17934_;
  assign new_n17942_ = new_n8628_ & new_n17934_;
  assign new_n17943_ = new_n8630_ & new_n17934_;
  assign new_n17944_ = ~new_n17942_ & ~new_n17943_;
  assign new_n17945_ = ~new_n17941_ & new_n17944_;
  assign new_n17946_ = new_n8637_ & new_n17934_;
  assign new_n17947_ = new_n8639_ & new_n17934_;
  assign new_n17948_ = ~new_n17946_ & ~new_n17947_;
  assign new_n17949_ = new_n17945_ & new_n17948_;
  assign new_n17950_ = new_n17940_ & new_n17949_;
  assign new_n17951_ = new_n17928_ & new_n17950_;
  assign new_n17952_ = new_n17905_ & new_n17951_;
  assign new_n17953_ = new_n8650_ & new_n17934_;
  assign new_n17954_ = new_n8635_ & new_n17934_;
  assign new_n17955_ = new_n8648_ & new_n17934_;
  assign new_n17956_ = ~new_n17954_ & ~new_n17955_;
  assign new_n17957_ = ~new_n17953_ & new_n17956_;
  assign new_n17958_ = new_n8659_ & new_n17934_;
  assign new_n17959_ = new_n8646_ & new_n17934_;
  assign new_n17960_ = new_n8657_ & new_n17934_;
  assign new_n17961_ = ~new_n17959_ & ~new_n17960_;
  assign new_n17962_ = ~new_n17958_ & new_n17961_;
  assign new_n17963_ = new_n17957_ & new_n17962_;
  assign new_n17964_ = new_n8670_ & new_n17934_;
  assign new_n17965_ = new_n8655_ & new_n17934_;
  assign new_n17966_ = new_n8667_ & new_n17934_;
  assign new_n17967_ = ~new_n17965_ & ~new_n17966_;
  assign new_n17968_ = ~new_n17964_ & new_n17967_;
  assign new_n17969_ = new_n8681_ & new_n17934_;
  assign new_n17970_ = new_n8665_ & new_n17934_;
  assign new_n17971_ = new_n8678_ & new_n17934_;
  assign new_n17972_ = ~new_n17970_ & ~new_n17971_;
  assign new_n17973_ = ~new_n17969_ & new_n17972_;
  assign new_n17974_ = new_n17968_ & new_n17973_;
  assign new_n17975_ = new_n17963_ & new_n17974_;
  assign new_n17976_ = new_n8694_ & new_n17934_;
  assign new_n17977_ = new_n8675_ & new_n17934_;
  assign new_n17978_ = new_n8692_ & new_n17934_;
  assign new_n17979_ = ~new_n17977_ & ~new_n17978_;
  assign new_n17980_ = ~new_n17976_ & new_n17979_;
  assign new_n17981_ = new_n8701_ & new_n17934_;
  assign new_n17982_ = new_n8689_ & new_n17934_;
  assign new_n17983_ = new_n8699_ & new_n17934_;
  assign new_n17984_ = ~new_n17982_ & ~new_n17983_;
  assign new_n17985_ = ~new_n17981_ & new_n17984_;
  assign new_n17986_ = new_n17980_ & new_n17985_;
  assign new_n17987_ = new_n5768_ & new_n16678_;
  assign new_n17988_ = new_n8630_ & new_n17987_;
  assign new_n17989_ = new_n8617_ & new_n17987_;
  assign new_n17990_ = new_n8628_ & new_n17987_;
  assign new_n17991_ = ~new_n17989_ & ~new_n17990_;
  assign new_n17992_ = ~new_n17988_ & new_n17991_;
  assign new_n17993_ = new_n8625_ & new_n17987_;
  assign new_n17994_ = new_n8637_ & new_n17987_;
  assign new_n17995_ = ~new_n17993_ & ~new_n17994_;
  assign new_n17996_ = new_n17992_ & new_n17995_;
  assign new_n17997_ = new_n17986_ & new_n17996_;
  assign new_n17998_ = new_n17975_ & new_n17997_;
  assign new_n17999_ = new_n8648_ & new_n17987_;
  assign new_n18000_ = new_n8639_ & new_n17987_;
  assign new_n18001_ = new_n8635_ & new_n17987_;
  assign new_n18002_ = ~new_n18000_ & ~new_n18001_;
  assign new_n18003_ = ~new_n17999_ & new_n18002_;
  assign new_n18004_ = new_n8657_ & new_n17987_;
  assign new_n18005_ = new_n8650_ & new_n17987_;
  assign new_n18006_ = new_n8646_ & new_n17987_;
  assign new_n18007_ = ~new_n18005_ & ~new_n18006_;
  assign new_n18008_ = ~new_n18004_ & new_n18007_;
  assign new_n18009_ = new_n18003_ & new_n18008_;
  assign new_n18010_ = new_n8667_ & new_n17987_;
  assign new_n18011_ = new_n8659_ & new_n17987_;
  assign new_n18012_ = new_n8655_ & new_n17987_;
  assign new_n18013_ = ~new_n18011_ & ~new_n18012_;
  assign new_n18014_ = ~new_n18010_ & new_n18013_;
  assign new_n18015_ = new_n8678_ & new_n17987_;
  assign new_n18016_ = new_n8670_ & new_n17987_;
  assign new_n18017_ = new_n8665_ & new_n17987_;
  assign new_n18018_ = ~new_n18016_ & ~new_n18017_;
  assign new_n18019_ = ~new_n18015_ & new_n18018_;
  assign new_n18020_ = new_n18014_ & new_n18019_;
  assign new_n18021_ = new_n18009_ & new_n18020_;
  assign new_n18022_ = new_n8692_ & new_n17987_;
  assign new_n18023_ = new_n8681_ & new_n17987_;
  assign new_n18024_ = new_n8675_ & new_n17987_;
  assign new_n18025_ = ~new_n18023_ & ~new_n18024_;
  assign new_n18026_ = ~new_n18022_ & new_n18025_;
  assign new_n18027_ = new_n8699_ & new_n17987_;
  assign new_n18028_ = new_n8694_ & new_n17987_;
  assign new_n18029_ = new_n8689_ & new_n17987_;
  assign new_n18030_ = ~new_n18028_ & ~new_n18029_;
  assign new_n18031_ = ~new_n18027_ & new_n18030_;
  assign new_n18032_ = new_n18026_ & new_n18031_;
  assign new_n18033_ = new_n5768_ & new_n16727_;
  assign new_n18034_ = new_n8628_ & new_n18033_;
  assign new_n18035_ = new_n8701_ & new_n17987_;
  assign new_n18036_ = new_n8617_ & new_n18033_;
  assign new_n18037_ = ~new_n18035_ & ~new_n18036_;
  assign new_n18038_ = ~new_n18034_ & new_n18037_;
  assign new_n18039_ = new_n8630_ & new_n18033_;
  assign new_n18040_ = new_n8625_ & new_n18033_;
  assign new_n18041_ = ~new_n18039_ & ~new_n18040_;
  assign new_n18042_ = new_n18038_ & new_n18041_;
  assign new_n18043_ = new_n18032_ & new_n18042_;
  assign new_n18044_ = new_n18021_ & new_n18043_;
  assign new_n18045_ = new_n17998_ & new_n18044_;
  assign new_n18046_ = new_n17952_ & new_n18045_;
  assign new_n18047_ = new_n17859_ & new_n18046_;
  assign new_n18048_ = new_n8635_ & new_n18033_;
  assign new_n18049_ = new_n8637_ & new_n18033_;
  assign new_n18050_ = new_n8639_ & new_n18033_;
  assign new_n18051_ = ~new_n18049_ & ~new_n18050_;
  assign new_n18052_ = ~new_n18048_ & new_n18051_;
  assign new_n18053_ = new_n8646_ & new_n18033_;
  assign new_n18054_ = new_n8648_ & new_n18033_;
  assign new_n18055_ = new_n8650_ & new_n18033_;
  assign new_n18056_ = ~new_n18054_ & ~new_n18055_;
  assign new_n18057_ = ~new_n18053_ & new_n18056_;
  assign new_n18058_ = new_n18052_ & new_n18057_;
  assign new_n18059_ = new_n8655_ & new_n18033_;
  assign new_n18060_ = new_n8657_ & new_n18033_;
  assign new_n18061_ = new_n8659_ & new_n18033_;
  assign new_n18062_ = ~new_n18060_ & ~new_n18061_;
  assign new_n18063_ = ~new_n18059_ & new_n18062_;
  assign new_n18064_ = new_n8665_ & new_n18033_;
  assign new_n18065_ = new_n8667_ & new_n18033_;
  assign new_n18066_ = new_n8670_ & new_n18033_;
  assign new_n18067_ = ~new_n18065_ & ~new_n18066_;
  assign new_n18068_ = ~new_n18064_ & new_n18067_;
  assign new_n18069_ = new_n18063_ & new_n18068_;
  assign new_n18070_ = new_n18058_ & new_n18069_;
  assign new_n18071_ = new_n8675_ & new_n18033_;
  assign new_n18072_ = new_n8678_ & new_n18033_;
  assign new_n18073_ = new_n8681_ & new_n18033_;
  assign new_n18074_ = ~new_n18072_ & ~new_n18073_;
  assign new_n18075_ = ~new_n18071_ & new_n18074_;
  assign new_n18076_ = new_n8689_ & new_n18033_;
  assign new_n18077_ = new_n8692_ & new_n18033_;
  assign new_n18078_ = new_n8694_ & new_n18033_;
  assign new_n18079_ = ~new_n18077_ & ~new_n18078_;
  assign new_n18080_ = ~new_n18076_ & new_n18079_;
  assign new_n18081_ = new_n18075_ & new_n18080_;
  assign new_n18082_ = new_n5768_ & new_n16779_;
  assign new_n18083_ = new_n8845_ & new_n18082_;
  assign new_n18084_ = new_n8699_ & new_n18033_;
  assign new_n18085_ = new_n8701_ & new_n18033_;
  assign new_n18086_ = ~new_n18084_ & ~new_n18085_;
  assign new_n18087_ = ~new_n18083_ & new_n18086_;
  assign new_n18088_ = new_n8853_ & new_n18082_;
  assign new_n18089_ = new_n8855_ & new_n18082_;
  assign new_n18090_ = ~new_n18088_ & ~new_n18089_;
  assign new_n18091_ = new_n18087_ & new_n18090_;
  assign new_n18092_ = new_n18081_ & new_n18091_;
  assign new_n18093_ = new_n18070_ & new_n18092_;
  assign new_n18094_ = new_n8866_ & new_n18082_;
  assign new_n18095_ = new_n8851_ & new_n18082_;
  assign new_n18096_ = new_n8864_ & new_n18082_;
  assign new_n18097_ = ~new_n18095_ & ~new_n18096_;
  assign new_n18098_ = ~new_n18094_ & new_n18097_;
  assign new_n18099_ = new_n8874_ & new_n18082_;
  assign new_n18100_ = new_n8862_ & new_n18082_;
  assign new_n18101_ = new_n8872_ & new_n18082_;
  assign new_n18102_ = ~new_n18100_ & ~new_n18101_;
  assign new_n18103_ = ~new_n18099_ & new_n18102_;
  assign new_n18104_ = new_n18098_ & new_n18103_;
  assign new_n18105_ = new_n8884_ & new_n18082_;
  assign new_n18106_ = new_n8870_ & new_n18082_;
  assign new_n18107_ = new_n8882_ & new_n18082_;
  assign new_n18108_ = ~new_n18106_ & ~new_n18107_;
  assign new_n18109_ = ~new_n18105_ & new_n18108_;
  assign new_n18110_ = new_n8890_ & new_n18082_;
  assign new_n18111_ = new_n8880_ & new_n18082_;
  assign new_n18112_ = new_n8888_ & new_n18082_;
  assign new_n18113_ = ~new_n18111_ & ~new_n18112_;
  assign new_n18114_ = ~new_n18110_ & new_n18113_;
  assign new_n18115_ = new_n18109_ & new_n18114_;
  assign new_n18116_ = new_n18104_ & new_n18115_;
  assign new_n18117_ = new_n8896_ & new_n18082_;
  assign new_n18118_ = new_n8898_ & new_n18082_;
  assign new_n18119_ = new_n8900_ & new_n18082_;
  assign new_n18120_ = ~new_n18118_ & ~new_n18119_;
  assign new_n18121_ = ~new_n18117_ & new_n18120_;
  assign new_n18122_ = new_n8905_ & new_n18082_;
  assign new_n18123_ = new_n8907_ & new_n18082_;
  assign new_n18124_ = new_n8909_ & new_n18082_;
  assign new_n18125_ = ~new_n18123_ & ~new_n18124_;
  assign new_n18126_ = ~new_n18122_ & new_n18125_;
  assign new_n18127_ = new_n18121_ & new_n18126_;
  assign new_n18128_ = new_n8914_ & new_n18082_;
  assign new_n18129_ = new_n8916_ & new_n18082_;
  assign new_n18130_ = new_n8918_ & new_n18082_;
  assign new_n18131_ = ~new_n18129_ & ~new_n18130_;
  assign new_n18132_ = ~new_n18128_ & new_n18131_;
  assign new_n18133_ = new_n8925_ & new_n18082_;
  assign new_n18134_ = new_n8927_ & new_n18082_;
  assign new_n18135_ = ~new_n18133_ & ~new_n18134_;
  assign new_n18136_ = new_n18132_ & new_n18135_;
  assign new_n18137_ = new_n18127_ & new_n18136_;
  assign new_n18138_ = new_n18116_ & new_n18137_;
  assign new_n18139_ = new_n18093_ & new_n18138_;
  assign new_n18140_ = new_n8938_ & new_n18082_;
  assign new_n18141_ = new_n8923_ & new_n18082_;
  assign new_n18142_ = new_n8936_ & new_n18082_;
  assign new_n18143_ = ~new_n18141_ & ~new_n18142_;
  assign new_n18144_ = ~new_n18140_ & new_n18143_;
  assign new_n18145_ = new_n8945_ & new_n18082_;
  assign new_n18146_ = new_n8934_ & new_n18082_;
  assign new_n18147_ = new_n8943_ & new_n18082_;
  assign new_n18148_ = ~new_n18146_ & ~new_n18147_;
  assign new_n18149_ = ~new_n18145_ & new_n18148_;
  assign new_n18150_ = new_n18144_ & new_n18149_;
  assign new_n18151_ = new_n5788_ & new_n16845_;
  assign new_n18152_ = new_n9716_ & new_n18151_;
  assign new_n18153_ = new_n9718_ & new_n18151_;
  assign new_n18154_ = new_n9720_ & new_n18151_;
  assign new_n18155_ = ~new_n18153_ & ~new_n18154_;
  assign new_n18156_ = ~new_n18152_ & new_n18155_;
  assign new_n18157_ = new_n9727_ & new_n18151_;
  assign new_n18158_ = new_n9729_ & new_n18151_;
  assign new_n18159_ = new_n9731_ & new_n18151_;
  assign new_n18160_ = ~new_n18158_ & ~new_n18159_;
  assign new_n18161_ = ~new_n18157_ & new_n18160_;
  assign new_n18162_ = new_n18156_ & new_n18161_;
  assign new_n18163_ = new_n18150_ & new_n18162_;
  assign new_n18164_ = new_n9735_ & new_n18151_;
  assign new_n18165_ = new_n9737_ & new_n18151_;
  assign new_n18166_ = new_n9739_ & new_n18151_;
  assign new_n18167_ = ~new_n18165_ & ~new_n18166_;
  assign new_n18168_ = ~new_n18164_ & new_n18167_;
  assign new_n18169_ = new_n9744_ & new_n18151_;
  assign new_n18170_ = new_n9746_ & new_n18151_;
  assign new_n18171_ = new_n9748_ & new_n18151_;
  assign new_n18172_ = ~new_n18170_ & ~new_n18171_;
  assign new_n18173_ = ~new_n18169_ & new_n18172_;
  assign new_n18174_ = new_n18168_ & new_n18173_;
  assign new_n18175_ = new_n9763_ & new_n18151_;
  assign new_n18176_ = new_n9753_ & new_n18151_;
  assign new_n18177_ = new_n9755_ & new_n18151_;
  assign new_n18178_ = ~new_n18176_ & ~new_n18177_;
  assign new_n18179_ = ~new_n18175_ & new_n18178_;
  assign new_n18180_ = new_n9765_ & new_n18151_;
  assign new_n18181_ = new_n9761_ & new_n18151_;
  assign new_n18182_ = ~new_n18180_ & ~new_n18181_;
  assign new_n18183_ = new_n18179_ & new_n18182_;
  assign new_n18184_ = new_n18174_ & new_n18183_;
  assign new_n18185_ = new_n18163_ & new_n18184_;
  assign new_n18186_ = new_n9769_ & new_n18151_;
  assign new_n18187_ = new_n9771_ & new_n18151_;
  assign new_n18188_ = new_n9773_ & new_n18151_;
  assign new_n18189_ = ~new_n18187_ & ~new_n18188_;
  assign new_n18190_ = ~new_n18186_ & new_n18189_;
  assign new_n18191_ = new_n9779_ & new_n18151_;
  assign new_n18192_ = new_n9781_ & new_n18151_;
  assign new_n18193_ = new_n9783_ & new_n18151_;
  assign new_n18194_ = ~new_n18192_ & ~new_n18193_;
  assign new_n18195_ = ~new_n18191_ & new_n18194_;
  assign new_n18196_ = new_n18190_ & new_n18195_;
  assign new_n18197_ = new_n9788_ & new_n18151_;
  assign new_n18198_ = new_n9790_ & new_n18151_;
  assign new_n18199_ = new_n9792_ & new_n18151_;
  assign new_n18200_ = ~new_n18198_ & ~new_n18199_;
  assign new_n18201_ = ~new_n18197_ & new_n18200_;
  assign new_n18202_ = new_n9799_ & new_n18151_;
  assign new_n18203_ = new_n9801_ & new_n18151_;
  assign new_n18204_ = new_n9803_ & new_n18151_;
  assign new_n18205_ = ~new_n18203_ & ~new_n18204_;
  assign new_n18206_ = ~new_n18202_ & new_n18205_;
  assign new_n18207_ = new_n18201_ & new_n18206_;
  assign new_n18208_ = new_n18196_ & new_n18207_;
  assign new_n18209_ = new_n9807_ & new_n18151_;
  assign new_n18210_ = new_n9809_ & new_n18151_;
  assign new_n18211_ = new_n9811_ & new_n18151_;
  assign new_n18212_ = ~new_n18210_ & ~new_n18211_;
  assign new_n18213_ = ~new_n18209_ & new_n18212_;
  assign new_n18214_ = new_n5788_ & new_n16908_;
  assign new_n18215_ = new_n9817_ & new_n18214_;
  assign new_n18216_ = new_n9819_ & new_n18214_;
  assign new_n18217_ = new_n9821_ & new_n18214_;
  assign new_n18218_ = ~new_n18216_ & ~new_n18217_;
  assign new_n18219_ = ~new_n18215_ & new_n18218_;
  assign new_n18220_ = new_n18213_ & new_n18219_;
  assign new_n18221_ = new_n9842_ & new_n18214_;
  assign new_n18222_ = new_n9825_ & new_n18214_;
  assign new_n18223_ = new_n9828_ & new_n18214_;
  assign new_n18224_ = ~new_n18222_ & ~new_n18223_;
  assign new_n18225_ = ~new_n18221_ & new_n18224_;
  assign new_n18226_ = new_n9844_ & new_n18214_;
  assign new_n18227_ = new_n9840_ & new_n18214_;
  assign new_n18228_ = ~new_n18226_ & ~new_n18227_;
  assign new_n18229_ = new_n18225_ & new_n18228_;
  assign new_n18230_ = new_n18220_ & new_n18229_;
  assign new_n18231_ = new_n18208_ & new_n18230_;
  assign new_n18232_ = new_n18185_ & new_n18231_;
  assign new_n18233_ = new_n18139_ & new_n18232_;
  assign new_n18234_ = new_n9848_ & new_n18214_;
  assign new_n18235_ = new_n9850_ & new_n18214_;
  assign new_n18236_ = new_n9852_ & new_n18214_;
  assign new_n18237_ = ~new_n18235_ & ~new_n18236_;
  assign new_n18238_ = ~new_n18234_ & new_n18237_;
  assign new_n18239_ = new_n9858_ & new_n18214_;
  assign new_n18240_ = new_n9860_ & new_n18214_;
  assign new_n18241_ = new_n9862_ & new_n18214_;
  assign new_n18242_ = ~new_n18240_ & ~new_n18241_;
  assign new_n18243_ = ~new_n18239_ & new_n18242_;
  assign new_n18244_ = new_n18238_ & new_n18243_;
  assign new_n18245_ = new_n9866_ & new_n18214_;
  assign new_n18246_ = new_n9868_ & new_n18214_;
  assign new_n18247_ = new_n9870_ & new_n18214_;
  assign new_n18248_ = ~new_n18246_ & ~new_n18247_;
  assign new_n18249_ = ~new_n18245_ & new_n18248_;
  assign new_n18250_ = new_n9876_ & new_n18214_;
  assign new_n18251_ = new_n9878_ & new_n18214_;
  assign new_n18252_ = new_n9880_ & new_n18214_;
  assign new_n18253_ = ~new_n18251_ & ~new_n18252_;
  assign new_n18254_ = ~new_n18250_ & new_n18253_;
  assign new_n18255_ = new_n18249_ & new_n18254_;
  assign new_n18256_ = new_n18244_ & new_n18255_;
  assign new_n18257_ = new_n9885_ & new_n18214_;
  assign new_n18258_ = new_n9887_ & new_n18214_;
  assign new_n18259_ = new_n9889_ & new_n18214_;
  assign new_n18260_ = ~new_n18258_ & ~new_n18259_;
  assign new_n18261_ = ~new_n18257_ & new_n18260_;
  assign new_n18262_ = new_n9895_ & new_n18214_;
  assign new_n18263_ = new_n9897_ & new_n18214_;
  assign new_n18264_ = new_n9899_ & new_n18214_;
  assign new_n18265_ = ~new_n18263_ & ~new_n18264_;
  assign new_n18266_ = ~new_n18262_ & new_n18265_;
  assign new_n18267_ = new_n18261_ & new_n18266_;
  assign new_n18268_ = new_n9904_ & new_n18214_;
  assign new_n18269_ = new_n9906_ & new_n18214_;
  assign new_n18270_ = new_n9908_ & new_n18214_;
  assign new_n18271_ = ~new_n18269_ & ~new_n18270_;
  assign new_n18272_ = ~new_n18268_ & new_n18271_;
  assign new_n18273_ = new_n9917_ & new_n18214_;
  assign new_n18274_ = new_n9919_ & new_n18214_;
  assign new_n18275_ = ~new_n18273_ & ~new_n18274_;
  assign new_n18276_ = new_n18272_ & new_n18275_;
  assign new_n18277_ = new_n18267_ & new_n18276_;
  assign new_n18278_ = new_n18256_ & new_n18277_;
  assign new_n18279_ = new_n5788_ & new_n16978_;
  assign new_n18280_ = new_n9928_ & new_n18279_;
  assign new_n18281_ = new_n9915_ & new_n18214_;
  assign new_n18282_ = new_n9926_ & new_n18279_;
  assign new_n18283_ = ~new_n18281_ & ~new_n18282_;
  assign new_n18284_ = ~new_n18280_ & new_n18283_;
  assign new_n18285_ = new_n9938_ & new_n18279_;
  assign new_n18286_ = new_n9924_ & new_n18279_;
  assign new_n18287_ = new_n9936_ & new_n18279_;
  assign new_n18288_ = ~new_n18286_ & ~new_n18287_;
  assign new_n18289_ = ~new_n18285_ & new_n18288_;
  assign new_n18290_ = new_n18284_ & new_n18289_;
  assign new_n18291_ = new_n9946_ & new_n18279_;
  assign new_n18292_ = new_n9934_ & new_n18279_;
  assign new_n18293_ = new_n9944_ & new_n18279_;
  assign new_n18294_ = ~new_n18292_ & ~new_n18293_;
  assign new_n18295_ = ~new_n18291_ & new_n18294_;
  assign new_n18296_ = new_n9956_ & new_n18279_;
  assign new_n18297_ = new_n9942_ & new_n18279_;
  assign new_n18298_ = new_n9954_ & new_n18279_;
  assign new_n18299_ = ~new_n18297_ & ~new_n18298_;
  assign new_n18300_ = ~new_n18296_ & new_n18299_;
  assign new_n18301_ = new_n18295_ & new_n18300_;
  assign new_n18302_ = new_n18290_ & new_n18301_;
  assign new_n18303_ = new_n9965_ & new_n18279_;
  assign new_n18304_ = new_n9952_ & new_n18279_;
  assign new_n18305_ = new_n9963_ & new_n18279_;
  assign new_n18306_ = ~new_n18304_ & ~new_n18305_;
  assign new_n18307_ = ~new_n18303_ & new_n18306_;
  assign new_n18308_ = new_n9974_ & new_n18279_;
  assign new_n18309_ = new_n9961_ & new_n18279_;
  assign new_n18310_ = new_n9972_ & new_n18279_;
  assign new_n18311_ = ~new_n18309_ & ~new_n18310_;
  assign new_n18312_ = ~new_n18308_ & new_n18311_;
  assign new_n18313_ = new_n18307_ & new_n18312_;
  assign new_n18314_ = new_n9980_ & new_n18279_;
  assign new_n18315_ = new_n9970_ & new_n18279_;
  assign new_n18316_ = new_n9978_ & new_n18279_;
  assign new_n18317_ = ~new_n18315_ & ~new_n18316_;
  assign new_n18318_ = ~new_n18314_ & new_n18317_;
  assign new_n18319_ = new_n9990_ & new_n18279_;
  assign new_n18320_ = new_n9992_ & new_n18279_;
  assign new_n18321_ = ~new_n18319_ & ~new_n18320_;
  assign new_n18322_ = new_n18318_ & new_n18321_;
  assign new_n18323_ = new_n18313_ & new_n18322_;
  assign new_n18324_ = new_n18302_ & new_n18323_;
  assign new_n18325_ = new_n18278_ & new_n18324_;
  assign new_n18326_ = new_n10001_ & new_n18279_;
  assign new_n18327_ = new_n9988_ & new_n18279_;
  assign new_n18328_ = new_n9999_ & new_n18279_;
  assign new_n18329_ = ~new_n18327_ & ~new_n18328_;
  assign new_n18330_ = ~new_n18326_ & new_n18329_;
  assign new_n18331_ = new_n10011_ & new_n18279_;
  assign new_n18332_ = new_n9997_ & new_n18279_;
  assign new_n18333_ = new_n10009_ & new_n18279_;
  assign new_n18334_ = ~new_n18332_ & ~new_n18333_;
  assign new_n18335_ = ~new_n18331_ & new_n18334_;
  assign new_n18336_ = new_n18330_ & new_n18335_;
  assign new_n18337_ = new_n10019_ & new_n18279_;
  assign new_n18338_ = new_n10007_ & new_n18279_;
  assign new_n18339_ = new_n10017_ & new_n18279_;
  assign new_n18340_ = ~new_n18338_ & ~new_n18339_;
  assign new_n18341_ = ~new_n18337_ & new_n18340_;
  assign new_n18342_ = new_n10030_ & new_n18279_;
  assign new_n18343_ = new_n10015_ & new_n18279_;
  assign new_n18344_ = new_n10028_ & new_n18279_;
  assign new_n18345_ = ~new_n18343_ & ~new_n18344_;
  assign new_n18346_ = ~new_n18342_ & new_n18345_;
  assign new_n18347_ = new_n18341_ & new_n18346_;
  assign new_n18348_ = new_n18336_ & new_n18347_;
  assign new_n18349_ = new_n10039_ & new_n18279_;
  assign new_n18350_ = new_n10026_ & new_n18279_;
  assign new_n18351_ = new_n10037_ & new_n18279_;
  assign new_n18352_ = ~new_n18350_ & ~new_n18351_;
  assign new_n18353_ = ~new_n18349_ & new_n18352_;
  assign new_n18354_ = new_n10048_ & new_n18279_;
  assign new_n18355_ = new_n10035_ & new_n18279_;
  assign new_n18356_ = new_n10046_ & new_n18279_;
  assign new_n18357_ = ~new_n18355_ & ~new_n18356_;
  assign new_n18358_ = ~new_n18354_ & new_n18357_;
  assign new_n18359_ = new_n18353_ & new_n18358_;
  assign new_n18360_ = new_n10054_ & new_n18279_;
  assign new_n18361_ = new_n10044_ & new_n18279_;
  assign new_n18362_ = new_n10052_ & new_n18279_;
  assign new_n18363_ = ~new_n18361_ & ~new_n18362_;
  assign new_n18364_ = ~new_n18360_ & new_n18363_;
  assign new_n18365_ = new_n10063_ & new_n18279_;
  assign new_n18366_ = new_n10065_ & new_n18279_;
  assign new_n18367_ = ~new_n18365_ & ~new_n18366_;
  assign new_n18368_ = new_n18364_ & new_n18367_;
  assign new_n18369_ = new_n18359_ & new_n18368_;
  assign new_n18370_ = new_n18348_ & new_n18369_;
  assign new_n18371_ = new_n10073_ & new_n18279_;
  assign new_n18372_ = new_n10061_ & new_n18279_;
  assign new_n18373_ = new_n10071_ & new_n18279_;
  assign new_n18374_ = ~new_n18372_ & ~new_n18373_;
  assign new_n18375_ = ~new_n18371_ & new_n18374_;
  assign new_n18376_ = new_n10082_ & new_n18279_;
  assign new_n18377_ = new_n10069_ & new_n18279_;
  assign new_n18378_ = new_n10080_ & new_n18279_;
  assign new_n18379_ = ~new_n18377_ & ~new_n18378_;
  assign new_n18380_ = ~new_n18376_ & new_n18379_;
  assign new_n18381_ = new_n18375_ & new_n18380_;
  assign new_n18382_ = new_n10091_ & new_n18279_;
  assign new_n18383_ = new_n10078_ & new_n18279_;
  assign new_n18384_ = new_n10089_ & new_n18279_;
  assign new_n18385_ = ~new_n18383_ & ~new_n18384_;
  assign new_n18386_ = ~new_n18382_ & new_n18385_;
  assign new_n18387_ = new_n10102_ & new_n18279_;
  assign new_n18388_ = new_n10087_ & new_n18279_;
  assign new_n18389_ = new_n10100_ & new_n18279_;
  assign new_n18390_ = ~new_n18388_ & ~new_n18389_;
  assign new_n18391_ = ~new_n18387_ & new_n18390_;
  assign new_n18392_ = new_n18386_ & new_n18391_;
  assign new_n18393_ = new_n18381_ & new_n18392_;
  assign new_n18394_ = new_n10111_ & new_n18279_;
  assign new_n18395_ = new_n10098_ & new_n18279_;
  assign new_n18396_ = new_n10109_ & new_n18279_;
  assign new_n18397_ = ~new_n18395_ & ~new_n18396_;
  assign new_n18398_ = ~new_n18394_ & new_n18397_;
  assign new_n18399_ = new_n10120_ & new_n18279_;
  assign new_n18400_ = new_n10107_ & new_n18279_;
  assign new_n18401_ = new_n10118_ & new_n18279_;
  assign new_n18402_ = ~new_n18400_ & ~new_n18401_;
  assign new_n18403_ = ~new_n18399_ & new_n18402_;
  assign new_n18404_ = new_n18398_ & new_n18403_;
  assign new_n18405_ = new_n6525_ & new_n15778_;
  assign new_n18406_ = new_n8628_ & new_n18405_;
  assign new_n18407_ = new_n10116_ & new_n18279_;
  assign new_n18408_ = new_n8617_ & new_n18405_;
  assign new_n18409_ = ~new_n18407_ & ~new_n18408_;
  assign new_n18410_ = ~new_n18406_ & new_n18409_;
  assign new_n18411_ = new_n8630_ & new_n18405_;
  assign new_n18412_ = new_n8625_ & new_n18405_;
  assign new_n18413_ = ~new_n18411_ & ~new_n18412_;
  assign new_n18414_ = new_n18410_ & new_n18413_;
  assign new_n18415_ = new_n18404_ & new_n18414_;
  assign new_n18416_ = new_n18393_ & new_n18415_;
  assign new_n18417_ = new_n18370_ & new_n18416_;
  assign new_n18418_ = new_n18325_ & new_n18417_;
  assign new_n18419_ = new_n18233_ & new_n18418_;
  assign new_n18420_ = new_n18047_ & new_n18419_;
  assign new_n18421_ = new_n8635_ & new_n18405_;
  assign new_n18422_ = new_n8637_ & new_n18405_;
  assign new_n18423_ = new_n8639_ & new_n18405_;
  assign new_n18424_ = ~new_n18422_ & ~new_n18423_;
  assign new_n18425_ = ~new_n18421_ & new_n18424_;
  assign new_n18426_ = new_n8646_ & new_n18405_;
  assign new_n18427_ = new_n8648_ & new_n18405_;
  assign new_n18428_ = new_n8650_ & new_n18405_;
  assign new_n18429_ = ~new_n18427_ & ~new_n18428_;
  assign new_n18430_ = ~new_n18426_ & new_n18429_;
  assign new_n18431_ = new_n18425_ & new_n18430_;
  assign new_n18432_ = new_n8655_ & new_n18405_;
  assign new_n18433_ = new_n8657_ & new_n18405_;
  assign new_n18434_ = new_n8659_ & new_n18405_;
  assign new_n18435_ = ~new_n18433_ & ~new_n18434_;
  assign new_n18436_ = ~new_n18432_ & new_n18435_;
  assign new_n18437_ = new_n8665_ & new_n18405_;
  assign new_n18438_ = new_n8667_ & new_n18405_;
  assign new_n18439_ = new_n8670_ & new_n18405_;
  assign new_n18440_ = ~new_n18438_ & ~new_n18439_;
  assign new_n18441_ = ~new_n18437_ & new_n18440_;
  assign new_n18442_ = new_n18436_ & new_n18441_;
  assign new_n18443_ = new_n18431_ & new_n18442_;
  assign new_n18444_ = new_n8675_ & new_n18405_;
  assign new_n18445_ = new_n8678_ & new_n18405_;
  assign new_n18446_ = new_n8681_ & new_n18405_;
  assign new_n18447_ = ~new_n18445_ & ~new_n18446_;
  assign new_n18448_ = ~new_n18444_ & new_n18447_;
  assign new_n18449_ = new_n8689_ & new_n18405_;
  assign new_n18450_ = new_n8692_ & new_n18405_;
  assign new_n18451_ = new_n8694_ & new_n18405_;
  assign new_n18452_ = ~new_n18450_ & ~new_n18451_;
  assign new_n18453_ = ~new_n18449_ & new_n18452_;
  assign new_n18454_ = new_n18448_ & new_n18453_;
  assign new_n18455_ = new_n6525_ & new_n15830_;
  assign new_n18456_ = new_n8617_ & new_n18455_;
  assign new_n18457_ = new_n8699_ & new_n18405_;
  assign new_n18458_ = new_n8701_ & new_n18405_;
  assign new_n18459_ = ~new_n18457_ & ~new_n18458_;
  assign new_n18460_ = ~new_n18456_ & new_n18459_;
  assign new_n18461_ = new_n8625_ & new_n18455_;
  assign new_n18462_ = new_n8628_ & new_n18455_;
  assign new_n18463_ = new_n8630_ & new_n18455_;
  assign new_n18464_ = ~new_n18462_ & ~new_n18463_;
  assign new_n18465_ = ~new_n18461_ & new_n18464_;
  assign new_n18466_ = new_n18460_ & new_n18465_;
  assign new_n18467_ = new_n18454_ & new_n18466_;
  assign new_n18468_ = new_n18443_ & new_n18467_;
  assign new_n18469_ = new_n8635_ & new_n18455_;
  assign new_n18470_ = new_n8637_ & new_n18455_;
  assign new_n18471_ = new_n8639_ & new_n18455_;
  assign new_n18472_ = ~new_n18470_ & ~new_n18471_;
  assign new_n18473_ = ~new_n18469_ & new_n18472_;
  assign new_n18474_ = new_n8646_ & new_n18455_;
  assign new_n18475_ = new_n8648_ & new_n18455_;
  assign new_n18476_ = new_n8650_ & new_n18455_;
  assign new_n18477_ = ~new_n18475_ & ~new_n18476_;
  assign new_n18478_ = ~new_n18474_ & new_n18477_;
  assign new_n18479_ = new_n18473_ & new_n18478_;
  assign new_n18480_ = new_n8655_ & new_n18455_;
  assign new_n18481_ = new_n8657_ & new_n18455_;
  assign new_n18482_ = new_n8659_ & new_n18455_;
  assign new_n18483_ = ~new_n18481_ & ~new_n18482_;
  assign new_n18484_ = ~new_n18480_ & new_n18483_;
  assign new_n18485_ = new_n8665_ & new_n18455_;
  assign new_n18486_ = new_n8667_ & new_n18455_;
  assign new_n18487_ = new_n8670_ & new_n18455_;
  assign new_n18488_ = ~new_n18486_ & ~new_n18487_;
  assign new_n18489_ = ~new_n18485_ & new_n18488_;
  assign new_n18490_ = new_n18484_ & new_n18489_;
  assign new_n18491_ = new_n18479_ & new_n18490_;
  assign new_n18492_ = new_n8675_ & new_n18455_;
  assign new_n18493_ = new_n8678_ & new_n18455_;
  assign new_n18494_ = new_n8681_ & new_n18455_;
  assign new_n18495_ = ~new_n18493_ & ~new_n18494_;
  assign new_n18496_ = ~new_n18492_ & new_n18495_;
  assign new_n18497_ = new_n8689_ & new_n18455_;
  assign new_n18498_ = new_n8692_ & new_n18455_;
  assign new_n18499_ = new_n8694_ & new_n18455_;
  assign new_n18500_ = ~new_n18498_ & ~new_n18499_;
  assign new_n18501_ = ~new_n18497_ & new_n18500_;
  assign new_n18502_ = new_n18496_ & new_n18501_;
  assign new_n18503_ = new_n6525_ & new_n15878_;
  assign new_n18504_ = new_n8617_ & new_n18503_;
  assign new_n18505_ = new_n8699_ & new_n18455_;
  assign new_n18506_ = new_n8701_ & new_n18455_;
  assign new_n18507_ = ~new_n18505_ & ~new_n18506_;
  assign new_n18508_ = ~new_n18504_ & new_n18507_;
  assign new_n18509_ = new_n8628_ & new_n18503_;
  assign new_n18510_ = new_n8630_ & new_n18503_;
  assign new_n18511_ = ~new_n18509_ & ~new_n18510_;
  assign new_n18512_ = new_n18508_ & new_n18511_;
  assign new_n18513_ = new_n18502_ & new_n18512_;
  assign new_n18514_ = new_n18491_ & new_n18513_;
  assign new_n18515_ = new_n18468_ & new_n18514_;
  assign new_n18516_ = new_n8639_ & new_n18503_;
  assign new_n18517_ = new_n8625_ & new_n18503_;
  assign new_n18518_ = new_n8637_ & new_n18503_;
  assign new_n18519_ = ~new_n18517_ & ~new_n18518_;
  assign new_n18520_ = ~new_n18516_ & new_n18519_;
  assign new_n18521_ = new_n8650_ & new_n18503_;
  assign new_n18522_ = new_n8635_ & new_n18503_;
  assign new_n18523_ = new_n8648_ & new_n18503_;
  assign new_n18524_ = ~new_n18522_ & ~new_n18523_;
  assign new_n18525_ = ~new_n18521_ & new_n18524_;
  assign new_n18526_ = new_n18520_ & new_n18525_;
  assign new_n18527_ = new_n8659_ & new_n18503_;
  assign new_n18528_ = new_n8646_ & new_n18503_;
  assign new_n18529_ = new_n8657_ & new_n18503_;
  assign new_n18530_ = ~new_n18528_ & ~new_n18529_;
  assign new_n18531_ = ~new_n18527_ & new_n18530_;
  assign new_n18532_ = new_n8670_ & new_n18503_;
  assign new_n18533_ = new_n8655_ & new_n18503_;
  assign new_n18534_ = new_n8667_ & new_n18503_;
  assign new_n18535_ = ~new_n18533_ & ~new_n18534_;
  assign new_n18536_ = ~new_n18532_ & new_n18535_;
  assign new_n18537_ = new_n18531_ & new_n18536_;
  assign new_n18538_ = new_n18526_ & new_n18537_;
  assign new_n18539_ = new_n8681_ & new_n18503_;
  assign new_n18540_ = new_n8665_ & new_n18503_;
  assign new_n18541_ = new_n8678_ & new_n18503_;
  assign new_n18542_ = ~new_n18540_ & ~new_n18541_;
  assign new_n18543_ = ~new_n18539_ & new_n18542_;
  assign new_n18544_ = new_n8694_ & new_n18503_;
  assign new_n18545_ = new_n8675_ & new_n18503_;
  assign new_n18546_ = new_n8692_ & new_n18503_;
  assign new_n18547_ = ~new_n18545_ & ~new_n18546_;
  assign new_n18548_ = ~new_n18544_ & new_n18547_;
  assign new_n18549_ = new_n18543_ & new_n18548_;
  assign new_n18550_ = new_n8701_ & new_n18503_;
  assign new_n18551_ = new_n8689_ & new_n18503_;
  assign new_n18552_ = new_n8699_ & new_n18503_;
  assign new_n18553_ = ~new_n18551_ & ~new_n18552_;
  assign new_n18554_ = ~new_n18550_ & new_n18553_;
  assign new_n18555_ = new_n6525_ & new_n15925_;
  assign new_n18556_ = new_n8617_ & new_n18555_;
  assign new_n18557_ = new_n8628_ & new_n18555_;
  assign new_n18558_ = ~new_n18556_ & ~new_n18557_;
  assign new_n18559_ = new_n18554_ & new_n18558_;
  assign new_n18560_ = new_n18549_ & new_n18559_;
  assign new_n18561_ = new_n18538_ & new_n18560_;
  assign new_n18562_ = new_n8637_ & new_n18555_;
  assign new_n18563_ = new_n8630_ & new_n18555_;
  assign new_n18564_ = new_n8625_ & new_n18555_;
  assign new_n18565_ = ~new_n18563_ & ~new_n18564_;
  assign new_n18566_ = ~new_n18562_ & new_n18565_;
  assign new_n18567_ = new_n8648_ & new_n18555_;
  assign new_n18568_ = new_n8639_ & new_n18555_;
  assign new_n18569_ = new_n8635_ & new_n18555_;
  assign new_n18570_ = ~new_n18568_ & ~new_n18569_;
  assign new_n18571_ = ~new_n18567_ & new_n18570_;
  assign new_n18572_ = new_n18566_ & new_n18571_;
  assign new_n18573_ = new_n8657_ & new_n18555_;
  assign new_n18574_ = new_n8650_ & new_n18555_;
  assign new_n18575_ = new_n8646_ & new_n18555_;
  assign new_n18576_ = ~new_n18574_ & ~new_n18575_;
  assign new_n18577_ = ~new_n18573_ & new_n18576_;
  assign new_n18578_ = new_n8667_ & new_n18555_;
  assign new_n18579_ = new_n8659_ & new_n18555_;
  assign new_n18580_ = new_n8655_ & new_n18555_;
  assign new_n18581_ = ~new_n18579_ & ~new_n18580_;
  assign new_n18582_ = ~new_n18578_ & new_n18581_;
  assign new_n18583_ = new_n18577_ & new_n18582_;
  assign new_n18584_ = new_n18572_ & new_n18583_;
  assign new_n18585_ = new_n8678_ & new_n18555_;
  assign new_n18586_ = new_n8670_ & new_n18555_;
  assign new_n18587_ = new_n8665_ & new_n18555_;
  assign new_n18588_ = ~new_n18586_ & ~new_n18587_;
  assign new_n18589_ = ~new_n18585_ & new_n18588_;
  assign new_n18590_ = new_n8692_ & new_n18555_;
  assign new_n18591_ = new_n8681_ & new_n18555_;
  assign new_n18592_ = new_n8675_ & new_n18555_;
  assign new_n18593_ = ~new_n18591_ & ~new_n18592_;
  assign new_n18594_ = ~new_n18590_ & new_n18593_;
  assign new_n18595_ = new_n18589_ & new_n18594_;
  assign new_n18596_ = new_n8699_ & new_n18555_;
  assign new_n18597_ = new_n8694_ & new_n18555_;
  assign new_n18598_ = new_n8689_ & new_n18555_;
  assign new_n18599_ = ~new_n18597_ & ~new_n18598_;
  assign new_n18600_ = ~new_n18596_ & new_n18599_;
  assign new_n18601_ = new_n8701_ & new_n18555_;
  assign new_n18602_ = new_n6525_ & new_n15981_;
  assign new_n18603_ = new_n8845_ & new_n18602_;
  assign new_n18604_ = ~new_n18601_ & ~new_n18603_;
  assign new_n18605_ = new_n18600_ & new_n18604_;
  assign new_n18606_ = new_n18595_ & new_n18605_;
  assign new_n18607_ = new_n18584_ & new_n18606_;
  assign new_n18608_ = new_n18561_ & new_n18607_;
  assign new_n18609_ = new_n18515_ & new_n18608_;
  assign new_n18610_ = new_n8851_ & new_n18602_;
  assign new_n18611_ = new_n8853_ & new_n18602_;
  assign new_n18612_ = new_n8855_ & new_n18602_;
  assign new_n18613_ = ~new_n18611_ & ~new_n18612_;
  assign new_n18614_ = ~new_n18610_ & new_n18613_;
  assign new_n18615_ = new_n8862_ & new_n18602_;
  assign new_n18616_ = new_n8864_ & new_n18602_;
  assign new_n18617_ = new_n8866_ & new_n18602_;
  assign new_n18618_ = ~new_n18616_ & ~new_n18617_;
  assign new_n18619_ = ~new_n18615_ & new_n18618_;
  assign new_n18620_ = new_n18614_ & new_n18619_;
  assign new_n18621_ = new_n8870_ & new_n18602_;
  assign new_n18622_ = new_n8872_ & new_n18602_;
  assign new_n18623_ = new_n8874_ & new_n18602_;
  assign new_n18624_ = ~new_n18622_ & ~new_n18623_;
  assign new_n18625_ = ~new_n18621_ & new_n18624_;
  assign new_n18626_ = new_n8880_ & new_n18602_;
  assign new_n18627_ = new_n8882_ & new_n18602_;
  assign new_n18628_ = new_n8884_ & new_n18602_;
  assign new_n18629_ = ~new_n18627_ & ~new_n18628_;
  assign new_n18630_ = ~new_n18626_ & new_n18629_;
  assign new_n18631_ = new_n18625_ & new_n18630_;
  assign new_n18632_ = new_n18620_ & new_n18631_;
  assign new_n18633_ = new_n8898_ & new_n18602_;
  assign new_n18634_ = new_n8888_ & new_n18602_;
  assign new_n18635_ = new_n8890_ & new_n18602_;
  assign new_n18636_ = ~new_n18634_ & ~new_n18635_;
  assign new_n18637_ = ~new_n18633_ & new_n18636_;
  assign new_n18638_ = new_n8907_ & new_n18602_;
  assign new_n18639_ = new_n8900_ & new_n18602_;
  assign new_n18640_ = new_n8896_ & new_n18602_;
  assign new_n18641_ = ~new_n18639_ & ~new_n18640_;
  assign new_n18642_ = ~new_n18638_ & new_n18641_;
  assign new_n18643_ = new_n18637_ & new_n18642_;
  assign new_n18644_ = new_n8916_ & new_n18602_;
  assign new_n18645_ = new_n8909_ & new_n18602_;
  assign new_n18646_ = new_n8905_ & new_n18602_;
  assign new_n18647_ = ~new_n18645_ & ~new_n18646_;
  assign new_n18648_ = ~new_n18644_ & new_n18647_;
  assign new_n18649_ = new_n8918_ & new_n18602_;
  assign new_n18650_ = new_n8914_ & new_n18602_;
  assign new_n18651_ = ~new_n18649_ & ~new_n18650_;
  assign new_n18652_ = new_n18648_ & new_n18651_;
  assign new_n18653_ = new_n18643_ & new_n18652_;
  assign new_n18654_ = new_n18632_ & new_n18653_;
  assign new_n18655_ = new_n8923_ & new_n18602_;
  assign new_n18656_ = new_n8925_ & new_n18602_;
  assign new_n18657_ = new_n8927_ & new_n18602_;
  assign new_n18658_ = ~new_n18656_ & ~new_n18657_;
  assign new_n18659_ = ~new_n18655_ & new_n18658_;
  assign new_n18660_ = new_n8934_ & new_n18602_;
  assign new_n18661_ = new_n8936_ & new_n18602_;
  assign new_n18662_ = new_n8938_ & new_n18602_;
  assign new_n18663_ = ~new_n18661_ & ~new_n18662_;
  assign new_n18664_ = ~new_n18660_ & new_n18663_;
  assign new_n18665_ = new_n18659_ & new_n18664_;
  assign new_n18666_ = new_n6533_ & new_n16044_;
  assign new_n18667_ = new_n8617_ & new_n18666_;
  assign new_n18668_ = new_n8943_ & new_n18602_;
  assign new_n18669_ = new_n8945_ & new_n18602_;
  assign new_n18670_ = ~new_n18668_ & ~new_n18669_;
  assign new_n18671_ = ~new_n18667_ & new_n18670_;
  assign new_n18672_ = new_n8625_ & new_n18666_;
  assign new_n18673_ = new_n8628_ & new_n18666_;
  assign new_n18674_ = new_n8630_ & new_n18666_;
  assign new_n18675_ = ~new_n18673_ & ~new_n18674_;
  assign new_n18676_ = ~new_n18672_ & new_n18675_;
  assign new_n18677_ = new_n18671_ & new_n18676_;
  assign new_n18678_ = new_n18665_ & new_n18677_;
  assign new_n18679_ = new_n8635_ & new_n18666_;
  assign new_n18680_ = new_n8637_ & new_n18666_;
  assign new_n18681_ = new_n8639_ & new_n18666_;
  assign new_n18682_ = ~new_n18680_ & ~new_n18681_;
  assign new_n18683_ = ~new_n18679_ & new_n18682_;
  assign new_n18684_ = new_n8646_ & new_n18666_;
  assign new_n18685_ = new_n8648_ & new_n18666_;
  assign new_n18686_ = new_n8650_ & new_n18666_;
  assign new_n18687_ = ~new_n18685_ & ~new_n18686_;
  assign new_n18688_ = ~new_n18684_ & new_n18687_;
  assign new_n18689_ = new_n18683_ & new_n18688_;
  assign new_n18690_ = new_n8655_ & new_n18666_;
  assign new_n18691_ = new_n8657_ & new_n18666_;
  assign new_n18692_ = new_n8659_ & new_n18666_;
  assign new_n18693_ = ~new_n18691_ & ~new_n18692_;
  assign new_n18694_ = ~new_n18690_ & new_n18693_;
  assign new_n18695_ = new_n8667_ & new_n18666_;
  assign new_n18696_ = new_n8670_ & new_n18666_;
  assign new_n18697_ = ~new_n18695_ & ~new_n18696_;
  assign new_n18698_ = new_n18694_ & new_n18697_;
  assign new_n18699_ = new_n18689_ & new_n18698_;
  assign new_n18700_ = new_n18678_ & new_n18699_;
  assign new_n18701_ = new_n18654_ & new_n18700_;
  assign new_n18702_ = new_n8681_ & new_n18666_;
  assign new_n18703_ = new_n8665_ & new_n18666_;
  assign new_n18704_ = new_n8678_ & new_n18666_;
  assign new_n18705_ = ~new_n18703_ & ~new_n18704_;
  assign new_n18706_ = ~new_n18702_ & new_n18705_;
  assign new_n18707_ = new_n8694_ & new_n18666_;
  assign new_n18708_ = new_n8675_ & new_n18666_;
  assign new_n18709_ = new_n8692_ & new_n18666_;
  assign new_n18710_ = ~new_n18708_ & ~new_n18709_;
  assign new_n18711_ = ~new_n18707_ & new_n18710_;
  assign new_n18712_ = new_n18706_ & new_n18711_;
  assign new_n18713_ = new_n8701_ & new_n18666_;
  assign new_n18714_ = new_n8689_ & new_n18666_;
  assign new_n18715_ = new_n8699_ & new_n18666_;
  assign new_n18716_ = ~new_n18714_ & ~new_n18715_;
  assign new_n18717_ = ~new_n18713_ & new_n18716_;
  assign new_n18718_ = new_n6533_ & new_n16093_;
  assign new_n18719_ = new_n8630_ & new_n18718_;
  assign new_n18720_ = new_n8617_ & new_n18718_;
  assign new_n18721_ = new_n8628_ & new_n18718_;
  assign new_n18722_ = ~new_n18720_ & ~new_n18721_;
  assign new_n18723_ = ~new_n18719_ & new_n18722_;
  assign new_n18724_ = new_n18717_ & new_n18723_;
  assign new_n18725_ = new_n18712_ & new_n18724_;
  assign new_n18726_ = new_n8639_ & new_n18718_;
  assign new_n18727_ = new_n8625_ & new_n18718_;
  assign new_n18728_ = new_n8637_ & new_n18718_;
  assign new_n18729_ = ~new_n18727_ & ~new_n18728_;
  assign new_n18730_ = ~new_n18726_ & new_n18729_;
  assign new_n18731_ = new_n8650_ & new_n18718_;
  assign new_n18732_ = new_n8635_ & new_n18718_;
  assign new_n18733_ = new_n8648_ & new_n18718_;
  assign new_n18734_ = ~new_n18732_ & ~new_n18733_;
  assign new_n18735_ = ~new_n18731_ & new_n18734_;
  assign new_n18736_ = new_n18730_ & new_n18735_;
  assign new_n18737_ = new_n8659_ & new_n18718_;
  assign new_n18738_ = new_n8646_ & new_n18718_;
  assign new_n18739_ = new_n8657_ & new_n18718_;
  assign new_n18740_ = ~new_n18738_ & ~new_n18739_;
  assign new_n18741_ = ~new_n18737_ & new_n18740_;
  assign new_n18742_ = new_n8655_ & new_n18718_;
  assign new_n18743_ = new_n8667_ & new_n18718_;
  assign new_n18744_ = ~new_n18742_ & ~new_n18743_;
  assign new_n18745_ = new_n18741_ & new_n18744_;
  assign new_n18746_ = new_n18736_ & new_n18745_;
  assign new_n18747_ = new_n18725_ & new_n18746_;
  assign new_n18748_ = new_n8678_ & new_n18718_;
  assign new_n18749_ = new_n8670_ & new_n18718_;
  assign new_n18750_ = new_n8665_ & new_n18718_;
  assign new_n18751_ = ~new_n18749_ & ~new_n18750_;
  assign new_n18752_ = ~new_n18748_ & new_n18751_;
  assign new_n18753_ = new_n8692_ & new_n18718_;
  assign new_n18754_ = new_n8681_ & new_n18718_;
  assign new_n18755_ = new_n8675_ & new_n18718_;
  assign new_n18756_ = ~new_n18754_ & ~new_n18755_;
  assign new_n18757_ = ~new_n18753_ & new_n18756_;
  assign new_n18758_ = new_n18752_ & new_n18757_;
  assign new_n18759_ = new_n8699_ & new_n18718_;
  assign new_n18760_ = new_n8694_ & new_n18718_;
  assign new_n18761_ = new_n8689_ & new_n18718_;
  assign new_n18762_ = ~new_n18760_ & ~new_n18761_;
  assign new_n18763_ = ~new_n18759_ & new_n18762_;
  assign new_n18764_ = new_n6533_ & new_n16151_;
  assign new_n18765_ = new_n8628_ & new_n18764_;
  assign new_n18766_ = new_n8701_ & new_n18718_;
  assign new_n18767_ = new_n8617_ & new_n18764_;
  assign new_n18768_ = ~new_n18766_ & ~new_n18767_;
  assign new_n18769_ = ~new_n18765_ & new_n18768_;
  assign new_n18770_ = new_n18763_ & new_n18769_;
  assign new_n18771_ = new_n18758_ & new_n18770_;
  assign new_n18772_ = new_n8637_ & new_n18764_;
  assign new_n18773_ = new_n8630_ & new_n18764_;
  assign new_n18774_ = new_n8625_ & new_n18764_;
  assign new_n18775_ = ~new_n18773_ & ~new_n18774_;
  assign new_n18776_ = ~new_n18772_ & new_n18775_;
  assign new_n18777_ = new_n8648_ & new_n18764_;
  assign new_n18778_ = new_n8639_ & new_n18764_;
  assign new_n18779_ = new_n8635_ & new_n18764_;
  assign new_n18780_ = ~new_n18778_ & ~new_n18779_;
  assign new_n18781_ = ~new_n18777_ & new_n18780_;
  assign new_n18782_ = new_n18776_ & new_n18781_;
  assign new_n18783_ = new_n8657_ & new_n18764_;
  assign new_n18784_ = new_n8650_ & new_n18764_;
  assign new_n18785_ = new_n8646_ & new_n18764_;
  assign new_n18786_ = ~new_n18784_ & ~new_n18785_;
  assign new_n18787_ = ~new_n18783_ & new_n18786_;
  assign new_n18788_ = new_n8659_ & new_n18764_;
  assign new_n18789_ = new_n8655_ & new_n18764_;
  assign new_n18790_ = ~new_n18788_ & ~new_n18789_;
  assign new_n18791_ = new_n18787_ & new_n18790_;
  assign new_n18792_ = new_n18782_ & new_n18791_;
  assign new_n18793_ = new_n18771_ & new_n18792_;
  assign new_n18794_ = new_n18747_ & new_n18793_;
  assign new_n18795_ = new_n18701_ & new_n18794_;
  assign new_n18796_ = new_n18609_ & new_n18795_;
  assign new_n18797_ = new_n8665_ & new_n18764_;
  assign new_n18798_ = new_n8667_ & new_n18764_;
  assign new_n18799_ = new_n8670_ & new_n18764_;
  assign new_n18800_ = ~new_n18798_ & ~new_n18799_;
  assign new_n18801_ = ~new_n18797_ & new_n18800_;
  assign new_n18802_ = new_n8675_ & new_n18764_;
  assign new_n18803_ = new_n8678_ & new_n18764_;
  assign new_n18804_ = new_n8681_ & new_n18764_;
  assign new_n18805_ = ~new_n18803_ & ~new_n18804_;
  assign new_n18806_ = ~new_n18802_ & new_n18805_;
  assign new_n18807_ = new_n18801_ & new_n18806_;
  assign new_n18808_ = new_n8689_ & new_n18764_;
  assign new_n18809_ = new_n8692_ & new_n18764_;
  assign new_n18810_ = new_n8694_ & new_n18764_;
  assign new_n18811_ = ~new_n18809_ & ~new_n18810_;
  assign new_n18812_ = ~new_n18808_ & new_n18811_;
  assign new_n18813_ = new_n6533_ & new_n16200_;
  assign new_n18814_ = new_n8617_ & new_n18813_;
  assign new_n18815_ = new_n8699_ & new_n18764_;
  assign new_n18816_ = new_n8701_ & new_n18764_;
  assign new_n18817_ = ~new_n18815_ & ~new_n18816_;
  assign new_n18818_ = ~new_n18814_ & new_n18817_;
  assign new_n18819_ = new_n18812_ & new_n18818_;
  assign new_n18820_ = new_n18807_ & new_n18819_;
  assign new_n18821_ = new_n8625_ & new_n18813_;
  assign new_n18822_ = new_n8628_ & new_n18813_;
  assign new_n18823_ = new_n8630_ & new_n18813_;
  assign new_n18824_ = ~new_n18822_ & ~new_n18823_;
  assign new_n18825_ = ~new_n18821_ & new_n18824_;
  assign new_n18826_ = new_n8635_ & new_n18813_;
  assign new_n18827_ = new_n8637_ & new_n18813_;
  assign new_n18828_ = new_n8639_ & new_n18813_;
  assign new_n18829_ = ~new_n18827_ & ~new_n18828_;
  assign new_n18830_ = ~new_n18826_ & new_n18829_;
  assign new_n18831_ = new_n18825_ & new_n18830_;
  assign new_n18832_ = new_n8646_ & new_n18813_;
  assign new_n18833_ = new_n8648_ & new_n18813_;
  assign new_n18834_ = new_n8650_ & new_n18813_;
  assign new_n18835_ = ~new_n18833_ & ~new_n18834_;
  assign new_n18836_ = ~new_n18832_ & new_n18835_;
  assign new_n18837_ = new_n8657_ & new_n18813_;
  assign new_n18838_ = new_n8659_ & new_n18813_;
  assign new_n18839_ = ~new_n18837_ & ~new_n18838_;
  assign new_n18840_ = new_n18836_ & new_n18839_;
  assign new_n18841_ = new_n18831_ & new_n18840_;
  assign new_n18842_ = new_n18820_ & new_n18841_;
  assign new_n18843_ = new_n8670_ & new_n18813_;
  assign new_n18844_ = new_n8655_ & new_n18813_;
  assign new_n18845_ = new_n8667_ & new_n18813_;
  assign new_n18846_ = ~new_n18844_ & ~new_n18845_;
  assign new_n18847_ = ~new_n18843_ & new_n18846_;
  assign new_n18848_ = new_n8681_ & new_n18813_;
  assign new_n18849_ = new_n8665_ & new_n18813_;
  assign new_n18850_ = new_n8678_ & new_n18813_;
  assign new_n18851_ = ~new_n18849_ & ~new_n18850_;
  assign new_n18852_ = ~new_n18848_ & new_n18851_;
  assign new_n18853_ = new_n18847_ & new_n18852_;
  assign new_n18854_ = new_n8694_ & new_n18813_;
  assign new_n18855_ = new_n8675_ & new_n18813_;
  assign new_n18856_ = new_n8692_ & new_n18813_;
  assign new_n18857_ = ~new_n18855_ & ~new_n18856_;
  assign new_n18858_ = ~new_n18854_ & new_n18857_;
  assign new_n18859_ = new_n8701_ & new_n18813_;
  assign new_n18860_ = new_n8689_ & new_n18813_;
  assign new_n18861_ = new_n8699_ & new_n18813_;
  assign new_n18862_ = ~new_n18860_ & ~new_n18861_;
  assign new_n18863_ = ~new_n18859_ & new_n18862_;
  assign new_n18864_ = new_n18858_ & new_n18863_;
  assign new_n18865_ = new_n18853_ & new_n18864_;
  assign new_n18866_ = new_n6533_ & new_n16248_;
  assign new_n18867_ = new_n8855_ & new_n18866_;
  assign new_n18868_ = new_n8845_ & new_n18866_;
  assign new_n18869_ = new_n8853_ & new_n18866_;
  assign new_n18870_ = ~new_n18868_ & ~new_n18869_;
  assign new_n18871_ = ~new_n18867_ & new_n18870_;
  assign new_n18872_ = new_n8866_ & new_n18866_;
  assign new_n18873_ = new_n8851_ & new_n18866_;
  assign new_n18874_ = new_n8864_ & new_n18866_;
  assign new_n18875_ = ~new_n18873_ & ~new_n18874_;
  assign new_n18876_ = ~new_n18872_ & new_n18875_;
  assign new_n18877_ = new_n18871_ & new_n18876_;
  assign new_n18878_ = new_n8874_ & new_n18866_;
  assign new_n18879_ = new_n8862_ & new_n18866_;
  assign new_n18880_ = new_n8872_ & new_n18866_;
  assign new_n18881_ = ~new_n18879_ & ~new_n18880_;
  assign new_n18882_ = ~new_n18878_ & new_n18881_;
  assign new_n18883_ = new_n8870_ & new_n18866_;
  assign new_n18884_ = new_n8882_ & new_n18866_;
  assign new_n18885_ = ~new_n18883_ & ~new_n18884_;
  assign new_n18886_ = new_n18882_ & new_n18885_;
  assign new_n18887_ = new_n18877_ & new_n18886_;
  assign new_n18888_ = new_n18865_ & new_n18887_;
  assign new_n18889_ = new_n18842_ & new_n18888_;
  assign new_n18890_ = new_n8888_ & new_n18866_;
  assign new_n18891_ = new_n8884_ & new_n18866_;
  assign new_n18892_ = new_n8880_ & new_n18866_;
  assign new_n18893_ = ~new_n18891_ & ~new_n18892_;
  assign new_n18894_ = ~new_n18890_ & new_n18893_;
  assign new_n18895_ = new_n8900_ & new_n18866_;
  assign new_n18896_ = new_n8890_ & new_n18866_;
  assign new_n18897_ = new_n8898_ & new_n18866_;
  assign new_n18898_ = ~new_n18896_ & ~new_n18897_;
  assign new_n18899_ = ~new_n18895_ & new_n18898_;
  assign new_n18900_ = new_n18894_ & new_n18899_;
  assign new_n18901_ = new_n8909_ & new_n18866_;
  assign new_n18902_ = new_n8896_ & new_n18866_;
  assign new_n18903_ = new_n8907_ & new_n18866_;
  assign new_n18904_ = ~new_n18902_ & ~new_n18903_;
  assign new_n18905_ = ~new_n18901_ & new_n18904_;
  assign new_n18906_ = new_n8918_ & new_n18866_;
  assign new_n18907_ = new_n8905_ & new_n18866_;
  assign new_n18908_ = new_n8916_ & new_n18866_;
  assign new_n18909_ = ~new_n18907_ & ~new_n18908_;
  assign new_n18910_ = ~new_n18906_ & new_n18909_;
  assign new_n18911_ = new_n18905_ & new_n18910_;
  assign new_n18912_ = new_n18900_ & new_n18911_;
  assign new_n18913_ = new_n8927_ & new_n18866_;
  assign new_n18914_ = new_n8914_ & new_n18866_;
  assign new_n18915_ = new_n8925_ & new_n18866_;
  assign new_n18916_ = ~new_n18914_ & ~new_n18915_;
  assign new_n18917_ = ~new_n18913_ & new_n18916_;
  assign new_n18918_ = new_n8938_ & new_n18866_;
  assign new_n18919_ = new_n8923_ & new_n18866_;
  assign new_n18920_ = new_n8936_ & new_n18866_;
  assign new_n18921_ = ~new_n18919_ & ~new_n18920_;
  assign new_n18922_ = ~new_n18918_ & new_n18921_;
  assign new_n18923_ = new_n18917_ & new_n18922_;
  assign new_n18924_ = new_n8945_ & new_n18866_;
  assign new_n18925_ = new_n8934_ & new_n18866_;
  assign new_n18926_ = new_n8943_ & new_n18866_;
  assign new_n18927_ = ~new_n18925_ & ~new_n18926_;
  assign new_n18928_ = ~new_n18924_ & new_n18927_;
  assign new_n18929_ = new_n6547_ & new_n16311_;
  assign new_n18930_ = new_n8617_ & new_n18929_;
  assign new_n18931_ = new_n8628_ & new_n18929_;
  assign new_n18932_ = ~new_n18930_ & ~new_n18931_;
  assign new_n18933_ = new_n18928_ & new_n18932_;
  assign new_n18934_ = new_n18923_ & new_n18933_;
  assign new_n18935_ = new_n18912_ & new_n18934_;
  assign new_n18936_ = new_n8637_ & new_n18929_;
  assign new_n18937_ = new_n8630_ & new_n18929_;
  assign new_n18938_ = new_n8625_ & new_n18929_;
  assign new_n18939_ = ~new_n18937_ & ~new_n18938_;
  assign new_n18940_ = ~new_n18936_ & new_n18939_;
  assign new_n18941_ = new_n8648_ & new_n18929_;
  assign new_n18942_ = new_n8639_ & new_n18929_;
  assign new_n18943_ = new_n8635_ & new_n18929_;
  assign new_n18944_ = ~new_n18942_ & ~new_n18943_;
  assign new_n18945_ = ~new_n18941_ & new_n18944_;
  assign new_n18946_ = new_n18940_ & new_n18945_;
  assign new_n18947_ = new_n8657_ & new_n18929_;
  assign new_n18948_ = new_n8650_ & new_n18929_;
  assign new_n18949_ = new_n8646_ & new_n18929_;
  assign new_n18950_ = ~new_n18948_ & ~new_n18949_;
  assign new_n18951_ = ~new_n18947_ & new_n18950_;
  assign new_n18952_ = new_n8667_ & new_n18929_;
  assign new_n18953_ = new_n8659_ & new_n18929_;
  assign new_n18954_ = new_n8655_ & new_n18929_;
  assign new_n18955_ = ~new_n18953_ & ~new_n18954_;
  assign new_n18956_ = ~new_n18952_ & new_n18955_;
  assign new_n18957_ = new_n18951_ & new_n18956_;
  assign new_n18958_ = new_n18946_ & new_n18957_;
  assign new_n18959_ = new_n8678_ & new_n18929_;
  assign new_n18960_ = new_n8670_ & new_n18929_;
  assign new_n18961_ = new_n8665_ & new_n18929_;
  assign new_n18962_ = ~new_n18960_ & ~new_n18961_;
  assign new_n18963_ = ~new_n18959_ & new_n18962_;
  assign new_n18964_ = new_n8692_ & new_n18929_;
  assign new_n18965_ = new_n8681_ & new_n18929_;
  assign new_n18966_ = new_n8675_ & new_n18929_;
  assign new_n18967_ = ~new_n18965_ & ~new_n18966_;
  assign new_n18968_ = ~new_n18964_ & new_n18967_;
  assign new_n18969_ = new_n18963_ & new_n18968_;
  assign new_n18970_ = new_n8699_ & new_n18929_;
  assign new_n18971_ = new_n8694_ & new_n18929_;
  assign new_n18972_ = new_n8689_ & new_n18929_;
  assign new_n18973_ = ~new_n18971_ & ~new_n18972_;
  assign new_n18974_ = ~new_n18970_ & new_n18973_;
  assign new_n18975_ = new_n8701_ & new_n18929_;
  assign new_n18976_ = new_n6547_ & new_n16360_;
  assign new_n18977_ = new_n8617_ & new_n18976_;
  assign new_n18978_ = ~new_n18975_ & ~new_n18977_;
  assign new_n18979_ = new_n18974_ & new_n18978_;
  assign new_n18980_ = new_n18969_ & new_n18979_;
  assign new_n18981_ = new_n18958_ & new_n18980_;
  assign new_n18982_ = new_n18935_ & new_n18981_;
  assign new_n18983_ = new_n18889_ & new_n18982_;
  assign new_n18984_ = new_n8625_ & new_n18976_;
  assign new_n18985_ = new_n8628_ & new_n18976_;
  assign new_n18986_ = new_n8630_ & new_n18976_;
  assign new_n18987_ = ~new_n18985_ & ~new_n18986_;
  assign new_n18988_ = ~new_n18984_ & new_n18987_;
  assign new_n18989_ = new_n8635_ & new_n18976_;
  assign new_n18990_ = new_n8637_ & new_n18976_;
  assign new_n18991_ = new_n8639_ & new_n18976_;
  assign new_n18992_ = ~new_n18990_ & ~new_n18991_;
  assign new_n18993_ = ~new_n18989_ & new_n18992_;
  assign new_n18994_ = new_n18988_ & new_n18993_;
  assign new_n18995_ = new_n8646_ & new_n18976_;
  assign new_n18996_ = new_n8648_ & new_n18976_;
  assign new_n18997_ = new_n8650_ & new_n18976_;
  assign new_n18998_ = ~new_n18996_ & ~new_n18997_;
  assign new_n18999_ = ~new_n18995_ & new_n18998_;
  assign new_n19000_ = new_n8655_ & new_n18976_;
  assign new_n19001_ = new_n8657_ & new_n18976_;
  assign new_n19002_ = new_n8659_ & new_n18976_;
  assign new_n19003_ = ~new_n19001_ & ~new_n19002_;
  assign new_n19004_ = ~new_n19000_ & new_n19003_;
  assign new_n19005_ = new_n18999_ & new_n19004_;
  assign new_n19006_ = new_n18994_ & new_n19005_;
  assign new_n19007_ = new_n8665_ & new_n18976_;
  assign new_n19008_ = new_n8667_ & new_n18976_;
  assign new_n19009_ = new_n8670_ & new_n18976_;
  assign new_n19010_ = ~new_n19008_ & ~new_n19009_;
  assign new_n19011_ = ~new_n19007_ & new_n19010_;
  assign new_n19012_ = new_n8675_ & new_n18976_;
  assign new_n19013_ = new_n8678_ & new_n18976_;
  assign new_n19014_ = new_n8681_ & new_n18976_;
  assign new_n19015_ = ~new_n19013_ & ~new_n19014_;
  assign new_n19016_ = ~new_n19012_ & new_n19015_;
  assign new_n19017_ = new_n19011_ & new_n19016_;
  assign new_n19018_ = new_n8689_ & new_n18976_;
  assign new_n19019_ = new_n8692_ & new_n18976_;
  assign new_n19020_ = new_n8694_ & new_n18976_;
  assign new_n19021_ = ~new_n19019_ & ~new_n19020_;
  assign new_n19022_ = ~new_n19018_ & new_n19021_;
  assign new_n19023_ = new_n8699_ & new_n18976_;
  assign new_n19024_ = new_n8701_ & new_n18976_;
  assign new_n19025_ = ~new_n19023_ & ~new_n19024_;
  assign new_n19026_ = new_n19022_ & new_n19025_;
  assign new_n19027_ = new_n19017_ & new_n19026_;
  assign new_n19028_ = new_n19006_ & new_n19027_;
  assign new_n19029_ = new_n6547_ & new_n16414_;
  assign new_n19030_ = new_n8630_ & new_n19029_;
  assign new_n19031_ = new_n8617_ & new_n19029_;
  assign new_n19032_ = new_n8628_ & new_n19029_;
  assign new_n19033_ = ~new_n19031_ & ~new_n19032_;
  assign new_n19034_ = ~new_n19030_ & new_n19033_;
  assign new_n19035_ = new_n8639_ & new_n19029_;
  assign new_n19036_ = new_n8625_ & new_n19029_;
  assign new_n19037_ = new_n8637_ & new_n19029_;
  assign new_n19038_ = ~new_n19036_ & ~new_n19037_;
  assign new_n19039_ = ~new_n19035_ & new_n19038_;
  assign new_n19040_ = new_n19034_ & new_n19039_;
  assign new_n19041_ = new_n8650_ & new_n19029_;
  assign new_n19042_ = new_n8635_ & new_n19029_;
  assign new_n19043_ = new_n8648_ & new_n19029_;
  assign new_n19044_ = ~new_n19042_ & ~new_n19043_;
  assign new_n19045_ = ~new_n19041_ & new_n19044_;
  assign new_n19046_ = new_n8659_ & new_n19029_;
  assign new_n19047_ = new_n8646_ & new_n19029_;
  assign new_n19048_ = new_n8657_ & new_n19029_;
  assign new_n19049_ = ~new_n19047_ & ~new_n19048_;
  assign new_n19050_ = ~new_n19046_ & new_n19049_;
  assign new_n19051_ = new_n19045_ & new_n19050_;
  assign new_n19052_ = new_n19040_ & new_n19051_;
  assign new_n19053_ = new_n8670_ & new_n19029_;
  assign new_n19054_ = new_n8655_ & new_n19029_;
  assign new_n19055_ = new_n8667_ & new_n19029_;
  assign new_n19056_ = ~new_n19054_ & ~new_n19055_;
  assign new_n19057_ = ~new_n19053_ & new_n19056_;
  assign new_n19058_ = new_n8681_ & new_n19029_;
  assign new_n19059_ = new_n8665_ & new_n19029_;
  assign new_n19060_ = new_n8678_ & new_n19029_;
  assign new_n19061_ = ~new_n19059_ & ~new_n19060_;
  assign new_n19062_ = ~new_n19058_ & new_n19061_;
  assign new_n19063_ = new_n19057_ & new_n19062_;
  assign new_n19064_ = new_n8694_ & new_n19029_;
  assign new_n19065_ = new_n8675_ & new_n19029_;
  assign new_n19066_ = new_n8692_ & new_n19029_;
  assign new_n19067_ = ~new_n19065_ & ~new_n19066_;
  assign new_n19068_ = ~new_n19064_ & new_n19067_;
  assign new_n19069_ = new_n8689_ & new_n19029_;
  assign new_n19070_ = new_n8699_ & new_n19029_;
  assign new_n19071_ = ~new_n19069_ & ~new_n19070_;
  assign new_n19072_ = new_n19068_ & new_n19071_;
  assign new_n19073_ = new_n19063_ & new_n19072_;
  assign new_n19074_ = new_n19052_ & new_n19073_;
  assign new_n19075_ = new_n19028_ & new_n19074_;
  assign new_n19076_ = new_n6547_ & new_n16462_;
  assign new_n19077_ = new_n8628_ & new_n19076_;
  assign new_n19078_ = new_n8701_ & new_n19029_;
  assign new_n19079_ = new_n8617_ & new_n19076_;
  assign new_n19080_ = ~new_n19078_ & ~new_n19079_;
  assign new_n19081_ = ~new_n19077_ & new_n19080_;
  assign new_n19082_ = new_n8637_ & new_n19076_;
  assign new_n19083_ = new_n8630_ & new_n19076_;
  assign new_n19084_ = new_n8625_ & new_n19076_;
  assign new_n19085_ = ~new_n19083_ & ~new_n19084_;
  assign new_n19086_ = ~new_n19082_ & new_n19085_;
  assign new_n19087_ = new_n19081_ & new_n19086_;
  assign new_n19088_ = new_n8648_ & new_n19076_;
  assign new_n19089_ = new_n8639_ & new_n19076_;
  assign new_n19090_ = new_n8635_ & new_n19076_;
  assign new_n19091_ = ~new_n19089_ & ~new_n19090_;
  assign new_n19092_ = ~new_n19088_ & new_n19091_;
  assign new_n19093_ = new_n8657_ & new_n19076_;
  assign new_n19094_ = new_n8650_ & new_n19076_;
  assign new_n19095_ = new_n8646_ & new_n19076_;
  assign new_n19096_ = ~new_n19094_ & ~new_n19095_;
  assign new_n19097_ = ~new_n19093_ & new_n19096_;
  assign new_n19098_ = new_n19092_ & new_n19097_;
  assign new_n19099_ = new_n19087_ & new_n19098_;
  assign new_n19100_ = new_n8667_ & new_n19076_;
  assign new_n19101_ = new_n8659_ & new_n19076_;
  assign new_n19102_ = new_n8655_ & new_n19076_;
  assign new_n19103_ = ~new_n19101_ & ~new_n19102_;
  assign new_n19104_ = ~new_n19100_ & new_n19103_;
  assign new_n19105_ = new_n8678_ & new_n19076_;
  assign new_n19106_ = new_n8670_ & new_n19076_;
  assign new_n19107_ = new_n8665_ & new_n19076_;
  assign new_n19108_ = ~new_n19106_ & ~new_n19107_;
  assign new_n19109_ = ~new_n19105_ & new_n19108_;
  assign new_n19110_ = new_n19104_ & new_n19109_;
  assign new_n19111_ = new_n8692_ & new_n19076_;
  assign new_n19112_ = new_n8681_ & new_n19076_;
  assign new_n19113_ = new_n8675_ & new_n19076_;
  assign new_n19114_ = ~new_n19112_ & ~new_n19113_;
  assign new_n19115_ = ~new_n19111_ & new_n19114_;
  assign new_n19116_ = new_n8694_ & new_n19076_;
  assign new_n19117_ = new_n8689_ & new_n19076_;
  assign new_n19118_ = ~new_n19116_ & ~new_n19117_;
  assign new_n19119_ = new_n19115_ & new_n19118_;
  assign new_n19120_ = new_n19110_ & new_n19119_;
  assign new_n19121_ = new_n19099_ & new_n19120_;
  assign new_n19122_ = new_n6547_ & new_n16509_;
  assign new_n19123_ = new_n8845_ & new_n19122_;
  assign new_n19124_ = new_n8699_ & new_n19076_;
  assign new_n19125_ = new_n8701_ & new_n19076_;
  assign new_n19126_ = ~new_n19124_ & ~new_n19125_;
  assign new_n19127_ = ~new_n19123_ & new_n19126_;
  assign new_n19128_ = new_n8851_ & new_n19122_;
  assign new_n19129_ = new_n8853_ & new_n19122_;
  assign new_n19130_ = new_n8855_ & new_n19122_;
  assign new_n19131_ = ~new_n19129_ & ~new_n19130_;
  assign new_n19132_ = ~new_n19128_ & new_n19131_;
  assign new_n19133_ = new_n19127_ & new_n19132_;
  assign new_n19134_ = new_n8862_ & new_n19122_;
  assign new_n19135_ = new_n8864_ & new_n19122_;
  assign new_n19136_ = new_n8866_ & new_n19122_;
  assign new_n19137_ = ~new_n19135_ & ~new_n19136_;
  assign new_n19138_ = ~new_n19134_ & new_n19137_;
  assign new_n19139_ = new_n8870_ & new_n19122_;
  assign new_n19140_ = new_n8872_ & new_n19122_;
  assign new_n19141_ = new_n8874_ & new_n19122_;
  assign new_n19142_ = ~new_n19140_ & ~new_n19141_;
  assign new_n19143_ = ~new_n19139_ & new_n19142_;
  assign new_n19144_ = new_n19138_ & new_n19143_;
  assign new_n19145_ = new_n19133_ & new_n19144_;
  assign new_n19146_ = new_n8880_ & new_n19122_;
  assign new_n19147_ = new_n8882_ & new_n19122_;
  assign new_n19148_ = new_n8884_ & new_n19122_;
  assign new_n19149_ = ~new_n19147_ & ~new_n19148_;
  assign new_n19150_ = ~new_n19146_ & new_n19149_;
  assign new_n19151_ = new_n8898_ & new_n19122_;
  assign new_n19152_ = new_n8888_ & new_n19122_;
  assign new_n19153_ = new_n8890_ & new_n19122_;
  assign new_n19154_ = ~new_n19152_ & ~new_n19153_;
  assign new_n19155_ = ~new_n19151_ & new_n19154_;
  assign new_n19156_ = new_n19150_ & new_n19155_;
  assign new_n19157_ = new_n8907_ & new_n19122_;
  assign new_n19158_ = new_n8900_ & new_n19122_;
  assign new_n19159_ = new_n8896_ & new_n19122_;
  assign new_n19160_ = ~new_n19158_ & ~new_n19159_;
  assign new_n19161_ = ~new_n19157_ & new_n19160_;
  assign new_n19162_ = new_n8909_ & new_n19122_;
  assign new_n19163_ = new_n8905_ & new_n19122_;
  assign new_n19164_ = ~new_n19162_ & ~new_n19163_;
  assign new_n19165_ = new_n19161_ & new_n19164_;
  assign new_n19166_ = new_n19156_ & new_n19165_;
  assign new_n19167_ = new_n19145_ & new_n19166_;
  assign new_n19168_ = new_n19121_ & new_n19167_;
  assign new_n19169_ = new_n19075_ & new_n19168_;
  assign new_n19170_ = new_n18983_ & new_n19169_;
  assign new_n19171_ = new_n18796_ & new_n19170_;
  assign new_n19172_ = new_n18420_ & new_n19171_;
  assign new_n19173_ = new_n17670_ & new_n19172_;
  assign new_n19174_ = new_n16150_ & new_n19173_;
  assign new_n19175_ = new_n8914_ & new_n19122_;
  assign new_n19176_ = new_n8916_ & new_n19122_;
  assign new_n19177_ = new_n8918_ & new_n19122_;
  assign new_n19178_ = ~new_n19176_ & ~new_n19177_;
  assign new_n19179_ = ~new_n19175_ & new_n19178_;
  assign new_n19180_ = new_n8923_ & new_n19122_;
  assign new_n19181_ = new_n8925_ & new_n19122_;
  assign new_n19182_ = new_n8927_ & new_n19122_;
  assign new_n19183_ = ~new_n19181_ & ~new_n19182_;
  assign new_n19184_ = ~new_n19180_ & new_n19183_;
  assign new_n19185_ = new_n19179_ & new_n19184_;
  assign new_n19186_ = new_n8934_ & new_n19122_;
  assign new_n19187_ = new_n8936_ & new_n19122_;
  assign new_n19188_ = new_n8938_ & new_n19122_;
  assign new_n19189_ = ~new_n19187_ & ~new_n19188_;
  assign new_n19190_ = ~new_n19186_ & new_n19189_;
  assign new_n19191_ = new_n6547_ & new_n16575_;
  assign new_n19192_ = new_n8617_ & new_n19191_;
  assign new_n19193_ = new_n8943_ & new_n19122_;
  assign new_n19194_ = new_n8945_ & new_n19122_;
  assign new_n19195_ = ~new_n19193_ & ~new_n19194_;
  assign new_n19196_ = ~new_n19192_ & new_n19195_;
  assign new_n19197_ = new_n19190_ & new_n19196_;
  assign new_n19198_ = new_n19185_ & new_n19197_;
  assign new_n19199_ = new_n8625_ & new_n19191_;
  assign new_n19200_ = new_n8628_ & new_n19191_;
  assign new_n19201_ = new_n8630_ & new_n19191_;
  assign new_n19202_ = ~new_n19200_ & ~new_n19201_;
  assign new_n19203_ = ~new_n19199_ & new_n19202_;
  assign new_n19204_ = new_n8635_ & new_n19191_;
  assign new_n19205_ = new_n8637_ & new_n19191_;
  assign new_n19206_ = new_n8639_ & new_n19191_;
  assign new_n19207_ = ~new_n19205_ & ~new_n19206_;
  assign new_n19208_ = ~new_n19204_ & new_n19207_;
  assign new_n19209_ = new_n19203_ & new_n19208_;
  assign new_n19210_ = new_n8646_ & new_n19191_;
  assign new_n19211_ = new_n8648_ & new_n19191_;
  assign new_n19212_ = new_n8650_ & new_n19191_;
  assign new_n19213_ = ~new_n19211_ & ~new_n19212_;
  assign new_n19214_ = ~new_n19210_ & new_n19213_;
  assign new_n19215_ = new_n8655_ & new_n19191_;
  assign new_n19216_ = new_n8657_ & new_n19191_;
  assign new_n19217_ = new_n8659_ & new_n19191_;
  assign new_n19218_ = ~new_n19216_ & ~new_n19217_;
  assign new_n19219_ = ~new_n19215_ & new_n19218_;
  assign new_n19220_ = new_n19214_ & new_n19219_;
  assign new_n19221_ = new_n19209_ & new_n19220_;
  assign new_n19222_ = new_n19198_ & new_n19221_;
  assign new_n19223_ = new_n8665_ & new_n19191_;
  assign new_n19224_ = new_n8667_ & new_n19191_;
  assign new_n19225_ = new_n8670_ & new_n19191_;
  assign new_n19226_ = ~new_n19224_ & ~new_n19225_;
  assign new_n19227_ = ~new_n19223_ & new_n19226_;
  assign new_n19228_ = new_n8675_ & new_n19191_;
  assign new_n19229_ = new_n8678_ & new_n19191_;
  assign new_n19230_ = new_n8681_ & new_n19191_;
  assign new_n19231_ = ~new_n19229_ & ~new_n19230_;
  assign new_n19232_ = ~new_n19228_ & new_n19231_;
  assign new_n19233_ = new_n19227_ & new_n19232_;
  assign new_n19234_ = new_n8689_ & new_n19191_;
  assign new_n19235_ = new_n8692_ & new_n19191_;
  assign new_n19236_ = new_n8694_ & new_n19191_;
  assign new_n19237_ = ~new_n19235_ & ~new_n19236_;
  assign new_n19238_ = ~new_n19234_ & new_n19237_;
  assign new_n19239_ = new_n6547_ & new_n16631_;
  assign new_n19240_ = new_n8617_ & new_n19239_;
  assign new_n19241_ = new_n8699_ & new_n19191_;
  assign new_n19242_ = new_n8701_ & new_n19191_;
  assign new_n19243_ = ~new_n19241_ & ~new_n19242_;
  assign new_n19244_ = ~new_n19240_ & new_n19243_;
  assign new_n19245_ = new_n19238_ & new_n19244_;
  assign new_n19246_ = new_n19233_ & new_n19245_;
  assign new_n19247_ = new_n8625_ & new_n19239_;
  assign new_n19248_ = new_n8628_ & new_n19239_;
  assign new_n19249_ = new_n8630_ & new_n19239_;
  assign new_n19250_ = ~new_n19248_ & ~new_n19249_;
  assign new_n19251_ = ~new_n19247_ & new_n19250_;
  assign new_n19252_ = new_n8635_ & new_n19239_;
  assign new_n19253_ = new_n8637_ & new_n19239_;
  assign new_n19254_ = new_n8639_ & new_n19239_;
  assign new_n19255_ = ~new_n19253_ & ~new_n19254_;
  assign new_n19256_ = ~new_n19252_ & new_n19255_;
  assign new_n19257_ = new_n19251_ & new_n19256_;
  assign new_n19258_ = new_n8646_ & new_n19239_;
  assign new_n19259_ = new_n8648_ & new_n19239_;
  assign new_n19260_ = new_n8650_ & new_n19239_;
  assign new_n19261_ = ~new_n19259_ & ~new_n19260_;
  assign new_n19262_ = ~new_n19258_ & new_n19261_;
  assign new_n19263_ = new_n8657_ & new_n19239_;
  assign new_n19264_ = new_n8659_ & new_n19239_;
  assign new_n19265_ = ~new_n19263_ & ~new_n19264_;
  assign new_n19266_ = new_n19262_ & new_n19265_;
  assign new_n19267_ = new_n19257_ & new_n19266_;
  assign new_n19268_ = new_n19246_ & new_n19267_;
  assign new_n19269_ = new_n19222_ & new_n19268_;
  assign new_n19270_ = new_n8670_ & new_n19239_;
  assign new_n19271_ = new_n8655_ & new_n19239_;
  assign new_n19272_ = new_n8667_ & new_n19239_;
  assign new_n19273_ = ~new_n19271_ & ~new_n19272_;
  assign new_n19274_ = ~new_n19270_ & new_n19273_;
  assign new_n19275_ = new_n8681_ & new_n19239_;
  assign new_n19276_ = new_n8665_ & new_n19239_;
  assign new_n19277_ = new_n8678_ & new_n19239_;
  assign new_n19278_ = ~new_n19276_ & ~new_n19277_;
  assign new_n19279_ = ~new_n19275_ & new_n19278_;
  assign new_n19280_ = new_n19274_ & new_n19279_;
  assign new_n19281_ = new_n8694_ & new_n19239_;
  assign new_n19282_ = new_n8675_ & new_n19239_;
  assign new_n19283_ = new_n8692_ & new_n19239_;
  assign new_n19284_ = ~new_n19282_ & ~new_n19283_;
  assign new_n19285_ = ~new_n19281_ & new_n19284_;
  assign new_n19286_ = new_n8701_ & new_n19239_;
  assign new_n19287_ = new_n8689_ & new_n19239_;
  assign new_n19288_ = new_n8699_ & new_n19239_;
  assign new_n19289_ = ~new_n19287_ & ~new_n19288_;
  assign new_n19290_ = ~new_n19286_ & new_n19289_;
  assign new_n19291_ = new_n19285_ & new_n19290_;
  assign new_n19292_ = new_n19280_ & new_n19291_;
  assign new_n19293_ = new_n6547_ & new_n16678_;
  assign new_n19294_ = new_n8630_ & new_n19293_;
  assign new_n19295_ = new_n8617_ & new_n19293_;
  assign new_n19296_ = new_n8628_ & new_n19293_;
  assign new_n19297_ = ~new_n19295_ & ~new_n19296_;
  assign new_n19298_ = ~new_n19294_ & new_n19297_;
  assign new_n19299_ = new_n8639_ & new_n19293_;
  assign new_n19300_ = new_n8625_ & new_n19293_;
  assign new_n19301_ = new_n8637_ & new_n19293_;
  assign new_n19302_ = ~new_n19300_ & ~new_n19301_;
  assign new_n19303_ = ~new_n19299_ & new_n19302_;
  assign new_n19304_ = new_n19298_ & new_n19303_;
  assign new_n19305_ = new_n8650_ & new_n19293_;
  assign new_n19306_ = new_n8635_ & new_n19293_;
  assign new_n19307_ = new_n8648_ & new_n19293_;
  assign new_n19308_ = ~new_n19306_ & ~new_n19307_;
  assign new_n19309_ = ~new_n19305_ & new_n19308_;
  assign new_n19310_ = new_n8646_ & new_n19293_;
  assign new_n19311_ = new_n8657_ & new_n19293_;
  assign new_n19312_ = ~new_n19310_ & ~new_n19311_;
  assign new_n19313_ = new_n19309_ & new_n19312_;
  assign new_n19314_ = new_n19304_ & new_n19313_;
  assign new_n19315_ = new_n19292_ & new_n19314_;
  assign new_n19316_ = new_n8667_ & new_n19293_;
  assign new_n19317_ = new_n8659_ & new_n19293_;
  assign new_n19318_ = new_n8655_ & new_n19293_;
  assign new_n19319_ = ~new_n19317_ & ~new_n19318_;
  assign new_n19320_ = ~new_n19316_ & new_n19319_;
  assign new_n19321_ = new_n8678_ & new_n19293_;
  assign new_n19322_ = new_n8670_ & new_n19293_;
  assign new_n19323_ = new_n8665_ & new_n19293_;
  assign new_n19324_ = ~new_n19322_ & ~new_n19323_;
  assign new_n19325_ = ~new_n19321_ & new_n19324_;
  assign new_n19326_ = new_n19320_ & new_n19325_;
  assign new_n19327_ = new_n8692_ & new_n19293_;
  assign new_n19328_ = new_n8681_ & new_n19293_;
  assign new_n19329_ = new_n8675_ & new_n19293_;
  assign new_n19330_ = ~new_n19328_ & ~new_n19329_;
  assign new_n19331_ = ~new_n19327_ & new_n19330_;
  assign new_n19332_ = new_n8699_ & new_n19293_;
  assign new_n19333_ = new_n8694_ & new_n19293_;
  assign new_n19334_ = new_n8689_ & new_n19293_;
  assign new_n19335_ = ~new_n19333_ & ~new_n19334_;
  assign new_n19336_ = ~new_n19332_ & new_n19335_;
  assign new_n19337_ = new_n19331_ & new_n19336_;
  assign new_n19338_ = new_n19326_ & new_n19337_;
  assign new_n19339_ = new_n6547_ & new_n16727_;
  assign new_n19340_ = new_n8628_ & new_n19339_;
  assign new_n19341_ = new_n8701_ & new_n19293_;
  assign new_n19342_ = new_n8617_ & new_n19339_;
  assign new_n19343_ = ~new_n19341_ & ~new_n19342_;
  assign new_n19344_ = ~new_n19340_ & new_n19343_;
  assign new_n19345_ = new_n8637_ & new_n19339_;
  assign new_n19346_ = new_n8630_ & new_n19339_;
  assign new_n19347_ = new_n8625_ & new_n19339_;
  assign new_n19348_ = ~new_n19346_ & ~new_n19347_;
  assign new_n19349_ = ~new_n19345_ & new_n19348_;
  assign new_n19350_ = new_n19344_ & new_n19349_;
  assign new_n19351_ = new_n8648_ & new_n19339_;
  assign new_n19352_ = new_n8639_ & new_n19339_;
  assign new_n19353_ = new_n8635_ & new_n19339_;
  assign new_n19354_ = ~new_n19352_ & ~new_n19353_;
  assign new_n19355_ = ~new_n19351_ & new_n19354_;
  assign new_n19356_ = new_n8650_ & new_n19339_;
  assign new_n19357_ = new_n8646_ & new_n19339_;
  assign new_n19358_ = ~new_n19356_ & ~new_n19357_;
  assign new_n19359_ = new_n19355_ & new_n19358_;
  assign new_n19360_ = new_n19350_ & new_n19359_;
  assign new_n19361_ = new_n19338_ & new_n19360_;
  assign new_n19362_ = new_n19315_ & new_n19361_;
  assign new_n19363_ = new_n19269_ & new_n19362_;
  assign new_n19364_ = new_n8655_ & new_n19339_;
  assign new_n19365_ = new_n8657_ & new_n19339_;
  assign new_n19366_ = new_n8659_ & new_n19339_;
  assign new_n19367_ = ~new_n19365_ & ~new_n19366_;
  assign new_n19368_ = ~new_n19364_ & new_n19367_;
  assign new_n19369_ = new_n8665_ & new_n19339_;
  assign new_n19370_ = new_n8667_ & new_n19339_;
  assign new_n19371_ = new_n8670_ & new_n19339_;
  assign new_n19372_ = ~new_n19370_ & ~new_n19371_;
  assign new_n19373_ = ~new_n19369_ & new_n19372_;
  assign new_n19374_ = new_n19368_ & new_n19373_;
  assign new_n19375_ = new_n8675_ & new_n19339_;
  assign new_n19376_ = new_n8678_ & new_n19339_;
  assign new_n19377_ = new_n8681_ & new_n19339_;
  assign new_n19378_ = ~new_n19376_ & ~new_n19377_;
  assign new_n19379_ = ~new_n19375_ & new_n19378_;
  assign new_n19380_ = new_n8689_ & new_n19339_;
  assign new_n19381_ = new_n8692_ & new_n19339_;
  assign new_n19382_ = new_n8694_ & new_n19339_;
  assign new_n19383_ = ~new_n19381_ & ~new_n19382_;
  assign new_n19384_ = ~new_n19380_ & new_n19383_;
  assign new_n19385_ = new_n19379_ & new_n19384_;
  assign new_n19386_ = new_n19374_ & new_n19385_;
  assign new_n19387_ = new_n6547_ & new_n16779_;
  assign new_n19388_ = new_n8845_ & new_n19387_;
  assign new_n19389_ = new_n8699_ & new_n19339_;
  assign new_n19390_ = new_n8701_ & new_n19339_;
  assign new_n19391_ = ~new_n19389_ & ~new_n19390_;
  assign new_n19392_ = ~new_n19388_ & new_n19391_;
  assign new_n19393_ = new_n8851_ & new_n19387_;
  assign new_n19394_ = new_n8853_ & new_n19387_;
  assign new_n19395_ = new_n8855_ & new_n19387_;
  assign new_n19396_ = ~new_n19394_ & ~new_n19395_;
  assign new_n19397_ = ~new_n19393_ & new_n19396_;
  assign new_n19398_ = new_n19392_ & new_n19397_;
  assign new_n19399_ = new_n8862_ & new_n19387_;
  assign new_n19400_ = new_n8864_ & new_n19387_;
  assign new_n19401_ = new_n8866_ & new_n19387_;
  assign new_n19402_ = ~new_n19400_ & ~new_n19401_;
  assign new_n19403_ = ~new_n19399_ & new_n19402_;
  assign new_n19404_ = new_n8872_ & new_n19387_;
  assign new_n19405_ = new_n8874_ & new_n19387_;
  assign new_n19406_ = ~new_n19404_ & ~new_n19405_;
  assign new_n19407_ = new_n19403_ & new_n19406_;
  assign new_n19408_ = new_n19398_ & new_n19407_;
  assign new_n19409_ = new_n19386_ & new_n19408_;
  assign new_n19410_ = new_n8884_ & new_n19387_;
  assign new_n19411_ = new_n8870_ & new_n19387_;
  assign new_n19412_ = new_n8882_ & new_n19387_;
  assign new_n19413_ = ~new_n19411_ & ~new_n19412_;
  assign new_n19414_ = ~new_n19410_ & new_n19413_;
  assign new_n19415_ = new_n8890_ & new_n19387_;
  assign new_n19416_ = new_n8880_ & new_n19387_;
  assign new_n19417_ = new_n8888_ & new_n19387_;
  assign new_n19418_ = ~new_n19416_ & ~new_n19417_;
  assign new_n19419_ = ~new_n19415_ & new_n19418_;
  assign new_n19420_ = new_n19414_ & new_n19419_;
  assign new_n19421_ = new_n8896_ & new_n19387_;
  assign new_n19422_ = new_n8898_ & new_n19387_;
  assign new_n19423_ = new_n8900_ & new_n19387_;
  assign new_n19424_ = ~new_n19422_ & ~new_n19423_;
  assign new_n19425_ = ~new_n19421_ & new_n19424_;
  assign new_n19426_ = new_n8905_ & new_n19387_;
  assign new_n19427_ = new_n8907_ & new_n19387_;
  assign new_n19428_ = new_n8909_ & new_n19387_;
  assign new_n19429_ = ~new_n19427_ & ~new_n19428_;
  assign new_n19430_ = ~new_n19426_ & new_n19429_;
  assign new_n19431_ = new_n19425_ & new_n19430_;
  assign new_n19432_ = new_n19420_ & new_n19431_;
  assign new_n19433_ = new_n8914_ & new_n19387_;
  assign new_n19434_ = new_n8916_ & new_n19387_;
  assign new_n19435_ = new_n8918_ & new_n19387_;
  assign new_n19436_ = ~new_n19434_ & ~new_n19435_;
  assign new_n19437_ = ~new_n19433_ & new_n19436_;
  assign new_n19438_ = new_n8923_ & new_n19387_;
  assign new_n19439_ = new_n8925_ & new_n19387_;
  assign new_n19440_ = new_n8927_ & new_n19387_;
  assign new_n19441_ = ~new_n19439_ & ~new_n19440_;
  assign new_n19442_ = ~new_n19438_ & new_n19441_;
  assign new_n19443_ = new_n19437_ & new_n19442_;
  assign new_n19444_ = new_n8934_ & new_n19387_;
  assign new_n19445_ = new_n8936_ & new_n19387_;
  assign new_n19446_ = new_n8938_ & new_n19387_;
  assign new_n19447_ = ~new_n19445_ & ~new_n19446_;
  assign new_n19448_ = ~new_n19444_ & new_n19447_;
  assign new_n19449_ = new_n8943_ & new_n19387_;
  assign new_n19450_ = new_n8945_ & new_n19387_;
  assign new_n19451_ = ~new_n19449_ & ~new_n19450_;
  assign new_n19452_ = new_n19448_ & new_n19451_;
  assign new_n19453_ = new_n19443_ & new_n19452_;
  assign new_n19454_ = new_n19432_ & new_n19453_;
  assign new_n19455_ = new_n19409_ & new_n19454_;
  assign new_n19456_ = new_n6568_ & new_n16845_;
  assign new_n19457_ = new_n9716_ & new_n19456_;
  assign new_n19458_ = new_n9718_ & new_n19456_;
  assign new_n19459_ = new_n9720_ & new_n19456_;
  assign new_n19460_ = ~new_n19458_ & ~new_n19459_;
  assign new_n19461_ = ~new_n19457_ & new_n19460_;
  assign new_n19462_ = new_n9727_ & new_n19456_;
  assign new_n19463_ = new_n9729_ & new_n19456_;
  assign new_n19464_ = new_n9731_ & new_n19456_;
  assign new_n19465_ = ~new_n19463_ & ~new_n19464_;
  assign new_n19466_ = ~new_n19462_ & new_n19465_;
  assign new_n19467_ = new_n19461_ & new_n19466_;
  assign new_n19468_ = new_n9735_ & new_n19456_;
  assign new_n19469_ = new_n9737_ & new_n19456_;
  assign new_n19470_ = new_n9739_ & new_n19456_;
  assign new_n19471_ = ~new_n19469_ & ~new_n19470_;
  assign new_n19472_ = ~new_n19468_ & new_n19471_;
  assign new_n19473_ = new_n9744_ & new_n19456_;
  assign new_n19474_ = new_n9746_ & new_n19456_;
  assign new_n19475_ = new_n9748_ & new_n19456_;
  assign new_n19476_ = ~new_n19474_ & ~new_n19475_;
  assign new_n19477_ = ~new_n19473_ & new_n19476_;
  assign new_n19478_ = new_n19472_ & new_n19477_;
  assign new_n19479_ = new_n19467_ & new_n19478_;
  assign new_n19480_ = new_n9763_ & new_n19456_;
  assign new_n19481_ = new_n9753_ & new_n19456_;
  assign new_n19482_ = new_n9755_ & new_n19456_;
  assign new_n19483_ = ~new_n19481_ & ~new_n19482_;
  assign new_n19484_ = ~new_n19480_ & new_n19483_;
  assign new_n19485_ = new_n9771_ & new_n19456_;
  assign new_n19486_ = new_n9765_ & new_n19456_;
  assign new_n19487_ = new_n9761_ & new_n19456_;
  assign new_n19488_ = ~new_n19486_ & ~new_n19487_;
  assign new_n19489_ = ~new_n19485_ & new_n19488_;
  assign new_n19490_ = new_n19484_ & new_n19489_;
  assign new_n19491_ = new_n9781_ & new_n19456_;
  assign new_n19492_ = new_n9773_ & new_n19456_;
  assign new_n19493_ = new_n9769_ & new_n19456_;
  assign new_n19494_ = ~new_n19492_ & ~new_n19493_;
  assign new_n19495_ = ~new_n19491_ & new_n19494_;
  assign new_n19496_ = new_n9783_ & new_n19456_;
  assign new_n19497_ = new_n9779_ & new_n19456_;
  assign new_n19498_ = ~new_n19496_ & ~new_n19497_;
  assign new_n19499_ = new_n19495_ & new_n19498_;
  assign new_n19500_ = new_n19490_ & new_n19499_;
  assign new_n19501_ = new_n19479_ & new_n19500_;
  assign new_n19502_ = new_n9788_ & new_n19456_;
  assign new_n19503_ = new_n9790_ & new_n19456_;
  assign new_n19504_ = new_n9792_ & new_n19456_;
  assign new_n19505_ = ~new_n19503_ & ~new_n19504_;
  assign new_n19506_ = ~new_n19502_ & new_n19505_;
  assign new_n19507_ = new_n9799_ & new_n19456_;
  assign new_n19508_ = new_n9801_ & new_n19456_;
  assign new_n19509_ = new_n9803_ & new_n19456_;
  assign new_n19510_ = ~new_n19508_ & ~new_n19509_;
  assign new_n19511_ = ~new_n19507_ & new_n19510_;
  assign new_n19512_ = new_n19506_ & new_n19511_;
  assign new_n19513_ = new_n9807_ & new_n19456_;
  assign new_n19514_ = new_n9809_ & new_n19456_;
  assign new_n19515_ = new_n9811_ & new_n19456_;
  assign new_n19516_ = ~new_n19514_ & ~new_n19515_;
  assign new_n19517_ = ~new_n19513_ & new_n19516_;
  assign new_n19518_ = new_n6568_ & new_n16908_;
  assign new_n19519_ = new_n9817_ & new_n19518_;
  assign new_n19520_ = new_n9819_ & new_n19518_;
  assign new_n19521_ = new_n9821_ & new_n19518_;
  assign new_n19522_ = ~new_n19520_ & ~new_n19521_;
  assign new_n19523_ = ~new_n19519_ & new_n19522_;
  assign new_n19524_ = new_n19517_ & new_n19523_;
  assign new_n19525_ = new_n19512_ & new_n19524_;
  assign new_n19526_ = new_n9842_ & new_n19518_;
  assign new_n19527_ = new_n9825_ & new_n19518_;
  assign new_n19528_ = new_n9828_ & new_n19518_;
  assign new_n19529_ = ~new_n19527_ & ~new_n19528_;
  assign new_n19530_ = ~new_n19526_ & new_n19529_;
  assign new_n19531_ = new_n9850_ & new_n19518_;
  assign new_n19532_ = new_n9844_ & new_n19518_;
  assign new_n19533_ = new_n9840_ & new_n19518_;
  assign new_n19534_ = ~new_n19532_ & ~new_n19533_;
  assign new_n19535_ = ~new_n19531_ & new_n19534_;
  assign new_n19536_ = new_n19530_ & new_n19535_;
  assign new_n19537_ = new_n9860_ & new_n19518_;
  assign new_n19538_ = new_n9852_ & new_n19518_;
  assign new_n19539_ = new_n9848_ & new_n19518_;
  assign new_n19540_ = ~new_n19538_ & ~new_n19539_;
  assign new_n19541_ = ~new_n19537_ & new_n19540_;
  assign new_n19542_ = new_n9862_ & new_n19518_;
  assign new_n19543_ = new_n9858_ & new_n19518_;
  assign new_n19544_ = ~new_n19542_ & ~new_n19543_;
  assign new_n19545_ = new_n19541_ & new_n19544_;
  assign new_n19546_ = new_n19536_ & new_n19545_;
  assign new_n19547_ = new_n19525_ & new_n19546_;
  assign new_n19548_ = new_n19501_ & new_n19547_;
  assign new_n19549_ = new_n19455_ & new_n19548_;
  assign new_n19550_ = new_n19363_ & new_n19549_;
  assign new_n19551_ = new_n9866_ & new_n19518_;
  assign new_n19552_ = new_n9868_ & new_n19518_;
  assign new_n19553_ = new_n9870_ & new_n19518_;
  assign new_n19554_ = ~new_n19552_ & ~new_n19553_;
  assign new_n19555_ = ~new_n19551_ & new_n19554_;
  assign new_n19556_ = new_n9876_ & new_n19518_;
  assign new_n19557_ = new_n9878_ & new_n19518_;
  assign new_n19558_ = new_n9880_ & new_n19518_;
  assign new_n19559_ = ~new_n19557_ & ~new_n19558_;
  assign new_n19560_ = ~new_n19556_ & new_n19559_;
  assign new_n19561_ = new_n19555_ & new_n19560_;
  assign new_n19562_ = new_n9885_ & new_n19518_;
  assign new_n19563_ = new_n9887_ & new_n19518_;
  assign new_n19564_ = new_n9889_ & new_n19518_;
  assign new_n19565_ = ~new_n19563_ & ~new_n19564_;
  assign new_n19566_ = ~new_n19562_ & new_n19565_;
  assign new_n19567_ = new_n9895_ & new_n19518_;
  assign new_n19568_ = new_n9897_ & new_n19518_;
  assign new_n19569_ = new_n9899_ & new_n19518_;
  assign new_n19570_ = ~new_n19568_ & ~new_n19569_;
  assign new_n19571_ = ~new_n19567_ & new_n19570_;
  assign new_n19572_ = new_n19566_ & new_n19571_;
  assign new_n19573_ = new_n19561_ & new_n19572_;
  assign new_n19574_ = new_n9904_ & new_n19518_;
  assign new_n19575_ = new_n9906_ & new_n19518_;
  assign new_n19576_ = new_n9908_ & new_n19518_;
  assign new_n19577_ = ~new_n19575_ & ~new_n19576_;
  assign new_n19578_ = ~new_n19574_ & new_n19577_;
  assign new_n19579_ = new_n9915_ & new_n19518_;
  assign new_n19580_ = new_n9917_ & new_n19518_;
  assign new_n19581_ = new_n9919_ & new_n19518_;
  assign new_n19582_ = ~new_n19580_ & ~new_n19581_;
  assign new_n19583_ = ~new_n19579_ & new_n19582_;
  assign new_n19584_ = new_n19578_ & new_n19583_;
  assign new_n19585_ = new_n6568_ & new_n16978_;
  assign new_n19586_ = new_n9924_ & new_n19585_;
  assign new_n19587_ = new_n9926_ & new_n19585_;
  assign new_n19588_ = new_n9928_ & new_n19585_;
  assign new_n19589_ = ~new_n19587_ & ~new_n19588_;
  assign new_n19590_ = ~new_n19586_ & new_n19589_;
  assign new_n19591_ = new_n9934_ & new_n19585_;
  assign new_n19592_ = new_n9936_ & new_n19585_;
  assign new_n19593_ = new_n9938_ & new_n19585_;
  assign new_n19594_ = ~new_n19592_ & ~new_n19593_;
  assign new_n19595_ = ~new_n19591_ & new_n19594_;
  assign new_n19596_ = new_n19590_ & new_n19595_;
  assign new_n19597_ = new_n19584_ & new_n19596_;
  assign new_n19598_ = new_n19573_ & new_n19597_;
  assign new_n19599_ = new_n9942_ & new_n19585_;
  assign new_n19600_ = new_n9944_ & new_n19585_;
  assign new_n19601_ = new_n9946_ & new_n19585_;
  assign new_n19602_ = ~new_n19600_ & ~new_n19601_;
  assign new_n19603_ = ~new_n19599_ & new_n19602_;
  assign new_n19604_ = new_n9952_ & new_n19585_;
  assign new_n19605_ = new_n9954_ & new_n19585_;
  assign new_n19606_ = new_n9956_ & new_n19585_;
  assign new_n19607_ = ~new_n19605_ & ~new_n19606_;
  assign new_n19608_ = ~new_n19604_ & new_n19607_;
  assign new_n19609_ = new_n19603_ & new_n19608_;
  assign new_n19610_ = new_n9961_ & new_n19585_;
  assign new_n19611_ = new_n9963_ & new_n19585_;
  assign new_n19612_ = new_n9965_ & new_n19585_;
  assign new_n19613_ = ~new_n19611_ & ~new_n19612_;
  assign new_n19614_ = ~new_n19610_ & new_n19613_;
  assign new_n19615_ = new_n9970_ & new_n19585_;
  assign new_n19616_ = new_n9972_ & new_n19585_;
  assign new_n19617_ = new_n9974_ & new_n19585_;
  assign new_n19618_ = ~new_n19616_ & ~new_n19617_;
  assign new_n19619_ = ~new_n19615_ & new_n19618_;
  assign new_n19620_ = new_n19614_ & new_n19619_;
  assign new_n19621_ = new_n19609_ & new_n19620_;
  assign new_n19622_ = new_n9990_ & new_n19585_;
  assign new_n19623_ = new_n9978_ & new_n19585_;
  assign new_n19624_ = new_n9980_ & new_n19585_;
  assign new_n19625_ = ~new_n19623_ & ~new_n19624_;
  assign new_n19626_ = ~new_n19622_ & new_n19625_;
  assign new_n19627_ = new_n9999_ & new_n19585_;
  assign new_n19628_ = new_n9992_ & new_n19585_;
  assign new_n19629_ = new_n9988_ & new_n19585_;
  assign new_n19630_ = ~new_n19628_ & ~new_n19629_;
  assign new_n19631_ = ~new_n19627_ & new_n19630_;
  assign new_n19632_ = new_n19626_ & new_n19631_;
  assign new_n19633_ = new_n10009_ & new_n19585_;
  assign new_n19634_ = new_n10001_ & new_n19585_;
  assign new_n19635_ = new_n9997_ & new_n19585_;
  assign new_n19636_ = ~new_n19634_ & ~new_n19635_;
  assign new_n19637_ = ~new_n19633_ & new_n19636_;
  assign new_n19638_ = new_n10011_ & new_n19585_;
  assign new_n19639_ = new_n10007_ & new_n19585_;
  assign new_n19640_ = ~new_n19638_ & ~new_n19639_;
  assign new_n19641_ = new_n19637_ & new_n19640_;
  assign new_n19642_ = new_n19632_ & new_n19641_;
  assign new_n19643_ = new_n19621_ & new_n19642_;
  assign new_n19644_ = new_n19598_ & new_n19643_;
  assign new_n19645_ = new_n10015_ & new_n19585_;
  assign new_n19646_ = new_n10017_ & new_n19585_;
  assign new_n19647_ = new_n10019_ & new_n19585_;
  assign new_n19648_ = ~new_n19646_ & ~new_n19647_;
  assign new_n19649_ = ~new_n19645_ & new_n19648_;
  assign new_n19650_ = new_n10026_ & new_n19585_;
  assign new_n19651_ = new_n10028_ & new_n19585_;
  assign new_n19652_ = new_n10030_ & new_n19585_;
  assign new_n19653_ = ~new_n19651_ & ~new_n19652_;
  assign new_n19654_ = ~new_n19650_ & new_n19653_;
  assign new_n19655_ = new_n19649_ & new_n19654_;
  assign new_n19656_ = new_n10035_ & new_n19585_;
  assign new_n19657_ = new_n10037_ & new_n19585_;
  assign new_n19658_ = new_n10039_ & new_n19585_;
  assign new_n19659_ = ~new_n19657_ & ~new_n19658_;
  assign new_n19660_ = ~new_n19656_ & new_n19659_;
  assign new_n19661_ = new_n10044_ & new_n19585_;
  assign new_n19662_ = new_n10046_ & new_n19585_;
  assign new_n19663_ = new_n10048_ & new_n19585_;
  assign new_n19664_ = ~new_n19662_ & ~new_n19663_;
  assign new_n19665_ = ~new_n19661_ & new_n19664_;
  assign new_n19666_ = new_n19660_ & new_n19665_;
  assign new_n19667_ = new_n19655_ & new_n19666_;
  assign new_n19668_ = new_n10063_ & new_n19585_;
  assign new_n19669_ = new_n10052_ & new_n19585_;
  assign new_n19670_ = new_n10054_ & new_n19585_;
  assign new_n19671_ = ~new_n19669_ & ~new_n19670_;
  assign new_n19672_ = ~new_n19668_ & new_n19671_;
  assign new_n19673_ = new_n10071_ & new_n19585_;
  assign new_n19674_ = new_n10065_ & new_n19585_;
  assign new_n19675_ = new_n10061_ & new_n19585_;
  assign new_n19676_ = ~new_n19674_ & ~new_n19675_;
  assign new_n19677_ = ~new_n19673_ & new_n19676_;
  assign new_n19678_ = new_n19672_ & new_n19677_;
  assign new_n19679_ = new_n10080_ & new_n19585_;
  assign new_n19680_ = new_n10073_ & new_n19585_;
  assign new_n19681_ = new_n10069_ & new_n19585_;
  assign new_n19682_ = ~new_n19680_ & ~new_n19681_;
  assign new_n19683_ = ~new_n19679_ & new_n19682_;
  assign new_n19684_ = new_n10082_ & new_n19585_;
  assign new_n19685_ = new_n10078_ & new_n19585_;
  assign new_n19686_ = ~new_n19684_ & ~new_n19685_;
  assign new_n19687_ = new_n19683_ & new_n19686_;
  assign new_n19688_ = new_n19678_ & new_n19687_;
  assign new_n19689_ = new_n19667_ & new_n19688_;
  assign new_n19690_ = new_n10087_ & new_n19585_;
  assign new_n19691_ = new_n10089_ & new_n19585_;
  assign new_n19692_ = new_n10091_ & new_n19585_;
  assign new_n19693_ = ~new_n19691_ & ~new_n19692_;
  assign new_n19694_ = ~new_n19690_ & new_n19693_;
  assign new_n19695_ = new_n10098_ & new_n19585_;
  assign new_n19696_ = new_n10100_ & new_n19585_;
  assign new_n19697_ = new_n10102_ & new_n19585_;
  assign new_n19698_ = ~new_n19696_ & ~new_n19697_;
  assign new_n19699_ = ~new_n19695_ & new_n19698_;
  assign new_n19700_ = new_n19694_ & new_n19699_;
  assign new_n19701_ = new_n10107_ & new_n19585_;
  assign new_n19702_ = new_n10109_ & new_n19585_;
  assign new_n19703_ = new_n10111_ & new_n19585_;
  assign new_n19704_ = ~new_n19702_ & ~new_n19703_;
  assign new_n19705_ = ~new_n19701_ & new_n19704_;
  assign new_n19706_ = new_n10116_ & new_n19585_;
  assign new_n19707_ = new_n10118_ & new_n19585_;
  assign new_n19708_ = new_n10120_ & new_n19585_;
  assign new_n19709_ = ~new_n19707_ & ~new_n19708_;
  assign new_n19710_ = ~new_n19706_ & new_n19709_;
  assign new_n19711_ = new_n19705_ & new_n19710_;
  assign new_n19712_ = new_n19700_ & new_n19711_;
  assign new_n19713_ = new_n6655_ & new_n15778_;
  assign new_n19714_ = new_n8630_ & new_n19713_;
  assign new_n19715_ = new_n8617_ & new_n19713_;
  assign new_n19716_ = new_n8628_ & new_n19713_;
  assign new_n19717_ = ~new_n19715_ & ~new_n19716_;
  assign new_n19718_ = ~new_n19714_ & new_n19717_;
  assign new_n19719_ = new_n8639_ & new_n19713_;
  assign new_n19720_ = new_n8625_ & new_n19713_;
  assign new_n19721_ = new_n8637_ & new_n19713_;
  assign new_n19722_ = ~new_n19720_ & ~new_n19721_;
  assign new_n19723_ = ~new_n19719_ & new_n19722_;
  assign new_n19724_ = new_n19718_ & new_n19723_;
  assign new_n19725_ = new_n8650_ & new_n19713_;
  assign new_n19726_ = new_n8635_ & new_n19713_;
  assign new_n19727_ = new_n8648_ & new_n19713_;
  assign new_n19728_ = ~new_n19726_ & ~new_n19727_;
  assign new_n19729_ = ~new_n19725_ & new_n19728_;
  assign new_n19730_ = new_n8646_ & new_n19713_;
  assign new_n19731_ = new_n8657_ & new_n19713_;
  assign new_n19732_ = ~new_n19730_ & ~new_n19731_;
  assign new_n19733_ = new_n19729_ & new_n19732_;
  assign new_n19734_ = new_n19724_ & new_n19733_;
  assign new_n19735_ = new_n19712_ & new_n19734_;
  assign new_n19736_ = new_n19689_ & new_n19735_;
  assign new_n19737_ = new_n19644_ & new_n19736_;
  assign new_n19738_ = new_n8667_ & new_n19713_;
  assign new_n19739_ = new_n8659_ & new_n19713_;
  assign new_n19740_ = new_n8655_ & new_n19713_;
  assign new_n19741_ = ~new_n19739_ & ~new_n19740_;
  assign new_n19742_ = ~new_n19738_ & new_n19741_;
  assign new_n19743_ = new_n8678_ & new_n19713_;
  assign new_n19744_ = new_n8670_ & new_n19713_;
  assign new_n19745_ = new_n8665_ & new_n19713_;
  assign new_n19746_ = ~new_n19744_ & ~new_n19745_;
  assign new_n19747_ = ~new_n19743_ & new_n19746_;
  assign new_n19748_ = new_n19742_ & new_n19747_;
  assign new_n19749_ = new_n8692_ & new_n19713_;
  assign new_n19750_ = new_n8681_ & new_n19713_;
  assign new_n19751_ = new_n8675_ & new_n19713_;
  assign new_n19752_ = ~new_n19750_ & ~new_n19751_;
  assign new_n19753_ = ~new_n19749_ & new_n19752_;
  assign new_n19754_ = new_n8699_ & new_n19713_;
  assign new_n19755_ = new_n8694_ & new_n19713_;
  assign new_n19756_ = new_n8689_ & new_n19713_;
  assign new_n19757_ = ~new_n19755_ & ~new_n19756_;
  assign new_n19758_ = ~new_n19754_ & new_n19757_;
  assign new_n19759_ = new_n19753_ & new_n19758_;
  assign new_n19760_ = new_n19748_ & new_n19759_;
  assign new_n19761_ = new_n6655_ & new_n15830_;
  assign new_n19762_ = new_n8628_ & new_n19761_;
  assign new_n19763_ = new_n8701_ & new_n19713_;
  assign new_n19764_ = new_n8617_ & new_n19761_;
  assign new_n19765_ = ~new_n19763_ & ~new_n19764_;
  assign new_n19766_ = ~new_n19762_ & new_n19765_;
  assign new_n19767_ = new_n8637_ & new_n19761_;
  assign new_n19768_ = new_n8630_ & new_n19761_;
  assign new_n19769_ = new_n8625_ & new_n19761_;
  assign new_n19770_ = ~new_n19768_ & ~new_n19769_;
  assign new_n19771_ = ~new_n19767_ & new_n19770_;
  assign new_n19772_ = new_n19766_ & new_n19771_;
  assign new_n19773_ = new_n8648_ & new_n19761_;
  assign new_n19774_ = new_n8639_ & new_n19761_;
  assign new_n19775_ = new_n8635_ & new_n19761_;
  assign new_n19776_ = ~new_n19774_ & ~new_n19775_;
  assign new_n19777_ = ~new_n19773_ & new_n19776_;
  assign new_n19778_ = new_n8650_ & new_n19761_;
  assign new_n19779_ = new_n8646_ & new_n19761_;
  assign new_n19780_ = ~new_n19778_ & ~new_n19779_;
  assign new_n19781_ = new_n19777_ & new_n19780_;
  assign new_n19782_ = new_n19772_ & new_n19781_;
  assign new_n19783_ = new_n19760_ & new_n19782_;
  assign new_n19784_ = new_n8655_ & new_n19761_;
  assign new_n19785_ = new_n8657_ & new_n19761_;
  assign new_n19786_ = new_n8659_ & new_n19761_;
  assign new_n19787_ = ~new_n19785_ & ~new_n19786_;
  assign new_n19788_ = ~new_n19784_ & new_n19787_;
  assign new_n19789_ = new_n8665_ & new_n19761_;
  assign new_n19790_ = new_n8667_ & new_n19761_;
  assign new_n19791_ = new_n8670_ & new_n19761_;
  assign new_n19792_ = ~new_n19790_ & ~new_n19791_;
  assign new_n19793_ = ~new_n19789_ & new_n19792_;
  assign new_n19794_ = new_n19788_ & new_n19793_;
  assign new_n19795_ = new_n8675_ & new_n19761_;
  assign new_n19796_ = new_n8678_ & new_n19761_;
  assign new_n19797_ = new_n8681_ & new_n19761_;
  assign new_n19798_ = ~new_n19796_ & ~new_n19797_;
  assign new_n19799_ = ~new_n19795_ & new_n19798_;
  assign new_n19800_ = new_n8689_ & new_n19761_;
  assign new_n19801_ = new_n8692_ & new_n19761_;
  assign new_n19802_ = new_n8694_ & new_n19761_;
  assign new_n19803_ = ~new_n19801_ & ~new_n19802_;
  assign new_n19804_ = ~new_n19800_ & new_n19803_;
  assign new_n19805_ = new_n19799_ & new_n19804_;
  assign new_n19806_ = new_n19794_ & new_n19805_;
  assign new_n19807_ = new_n6655_ & new_n15878_;
  assign new_n19808_ = new_n8617_ & new_n19807_;
  assign new_n19809_ = new_n8699_ & new_n19761_;
  assign new_n19810_ = new_n8701_ & new_n19761_;
  assign new_n19811_ = ~new_n19809_ & ~new_n19810_;
  assign new_n19812_ = ~new_n19808_ & new_n19811_;
  assign new_n19813_ = new_n8625_ & new_n19807_;
  assign new_n19814_ = new_n8628_ & new_n19807_;
  assign new_n19815_ = new_n8630_ & new_n19807_;
  assign new_n19816_ = ~new_n19814_ & ~new_n19815_;
  assign new_n19817_ = ~new_n19813_ & new_n19816_;
  assign new_n19818_ = new_n19812_ & new_n19817_;
  assign new_n19819_ = new_n8635_ & new_n19807_;
  assign new_n19820_ = new_n8637_ & new_n19807_;
  assign new_n19821_ = new_n8639_ & new_n19807_;
  assign new_n19822_ = ~new_n19820_ & ~new_n19821_;
  assign new_n19823_ = ~new_n19819_ & new_n19822_;
  assign new_n19824_ = new_n8648_ & new_n19807_;
  assign new_n19825_ = new_n8650_ & new_n19807_;
  assign new_n19826_ = ~new_n19824_ & ~new_n19825_;
  assign new_n19827_ = new_n19823_ & new_n19826_;
  assign new_n19828_ = new_n19818_ & new_n19827_;
  assign new_n19829_ = new_n19806_ & new_n19828_;
  assign new_n19830_ = new_n19783_ & new_n19829_;
  assign new_n19831_ = new_n8659_ & new_n19807_;
  assign new_n19832_ = new_n8646_ & new_n19807_;
  assign new_n19833_ = new_n8657_ & new_n19807_;
  assign new_n19834_ = ~new_n19832_ & ~new_n19833_;
  assign new_n19835_ = ~new_n19831_ & new_n19834_;
  assign new_n19836_ = new_n8670_ & new_n19807_;
  assign new_n19837_ = new_n8655_ & new_n19807_;
  assign new_n19838_ = new_n8667_ & new_n19807_;
  assign new_n19839_ = ~new_n19837_ & ~new_n19838_;
  assign new_n19840_ = ~new_n19836_ & new_n19839_;
  assign new_n19841_ = new_n19835_ & new_n19840_;
  assign new_n19842_ = new_n8681_ & new_n19807_;
  assign new_n19843_ = new_n8665_ & new_n19807_;
  assign new_n19844_ = new_n8678_ & new_n19807_;
  assign new_n19845_ = ~new_n19843_ & ~new_n19844_;
  assign new_n19846_ = ~new_n19842_ & new_n19845_;
  assign new_n19847_ = new_n8694_ & new_n19807_;
  assign new_n19848_ = new_n8675_ & new_n19807_;
  assign new_n19849_ = new_n8692_ & new_n19807_;
  assign new_n19850_ = ~new_n19848_ & ~new_n19849_;
  assign new_n19851_ = ~new_n19847_ & new_n19850_;
  assign new_n19852_ = new_n19846_ & new_n19851_;
  assign new_n19853_ = new_n19841_ & new_n19852_;
  assign new_n19854_ = new_n8701_ & new_n19807_;
  assign new_n19855_ = new_n8689_ & new_n19807_;
  assign new_n19856_ = new_n8699_ & new_n19807_;
  assign new_n19857_ = ~new_n19855_ & ~new_n19856_;
  assign new_n19858_ = ~new_n19854_ & new_n19857_;
  assign new_n19859_ = new_n6655_ & new_n15925_;
  assign new_n19860_ = new_n8630_ & new_n19859_;
  assign new_n19861_ = new_n8617_ & new_n19859_;
  assign new_n19862_ = new_n8628_ & new_n19859_;
  assign new_n19863_ = ~new_n19861_ & ~new_n19862_;
  assign new_n19864_ = ~new_n19860_ & new_n19863_;
  assign new_n19865_ = new_n19858_ & new_n19864_;
  assign new_n19866_ = new_n8639_ & new_n19859_;
  assign new_n19867_ = new_n8625_ & new_n19859_;
  assign new_n19868_ = new_n8637_ & new_n19859_;
  assign new_n19869_ = ~new_n19867_ & ~new_n19868_;
  assign new_n19870_ = ~new_n19866_ & new_n19869_;
  assign new_n19871_ = new_n8635_ & new_n19859_;
  assign new_n19872_ = new_n8648_ & new_n19859_;
  assign new_n19873_ = ~new_n19871_ & ~new_n19872_;
  assign new_n19874_ = new_n19870_ & new_n19873_;
  assign new_n19875_ = new_n19865_ & new_n19874_;
  assign new_n19876_ = new_n19853_ & new_n19875_;
  assign new_n19877_ = new_n8657_ & new_n19859_;
  assign new_n19878_ = new_n8650_ & new_n19859_;
  assign new_n19879_ = new_n8646_ & new_n19859_;
  assign new_n19880_ = ~new_n19878_ & ~new_n19879_;
  assign new_n19881_ = ~new_n19877_ & new_n19880_;
  assign new_n19882_ = new_n8667_ & new_n19859_;
  assign new_n19883_ = new_n8659_ & new_n19859_;
  assign new_n19884_ = new_n8655_ & new_n19859_;
  assign new_n19885_ = ~new_n19883_ & ~new_n19884_;
  assign new_n19886_ = ~new_n19882_ & new_n19885_;
  assign new_n19887_ = new_n19881_ & new_n19886_;
  assign new_n19888_ = new_n8678_ & new_n19859_;
  assign new_n19889_ = new_n8670_ & new_n19859_;
  assign new_n19890_ = new_n8665_ & new_n19859_;
  assign new_n19891_ = ~new_n19889_ & ~new_n19890_;
  assign new_n19892_ = ~new_n19888_ & new_n19891_;
  assign new_n19893_ = new_n8692_ & new_n19859_;
  assign new_n19894_ = new_n8681_ & new_n19859_;
  assign new_n19895_ = new_n8675_ & new_n19859_;
  assign new_n19896_ = ~new_n19894_ & ~new_n19895_;
  assign new_n19897_ = ~new_n19893_ & new_n19896_;
  assign new_n19898_ = new_n19892_ & new_n19897_;
  assign new_n19899_ = new_n19887_ & new_n19898_;
  assign new_n19900_ = new_n8699_ & new_n19859_;
  assign new_n19901_ = new_n8694_ & new_n19859_;
  assign new_n19902_ = new_n8689_ & new_n19859_;
  assign new_n19903_ = ~new_n19901_ & ~new_n19902_;
  assign new_n19904_ = ~new_n19900_ & new_n19903_;
  assign new_n19905_ = new_n6655_ & new_n15981_;
  assign new_n19906_ = new_n8853_ & new_n19905_;
  assign new_n19907_ = new_n8701_ & new_n19859_;
  assign new_n19908_ = new_n8845_ & new_n19905_;
  assign new_n19909_ = ~new_n19907_ & ~new_n19908_;
  assign new_n19910_ = ~new_n19906_ & new_n19909_;
  assign new_n19911_ = new_n19904_ & new_n19910_;
  assign new_n19912_ = new_n8864_ & new_n19905_;
  assign new_n19913_ = new_n8855_ & new_n19905_;
  assign new_n19914_ = new_n8851_ & new_n19905_;
  assign new_n19915_ = ~new_n19913_ & ~new_n19914_;
  assign new_n19916_ = ~new_n19912_ & new_n19915_;
  assign new_n19917_ = new_n8866_ & new_n19905_;
  assign new_n19918_ = new_n8862_ & new_n19905_;
  assign new_n19919_ = ~new_n19917_ & ~new_n19918_;
  assign new_n19920_ = new_n19916_ & new_n19919_;
  assign new_n19921_ = new_n19911_ & new_n19920_;
  assign new_n19922_ = new_n19899_ & new_n19921_;
  assign new_n19923_ = new_n19876_ & new_n19922_;
  assign new_n19924_ = new_n19830_ & new_n19923_;
  assign new_n19925_ = new_n19737_ & new_n19924_;
  assign new_n19926_ = new_n19550_ & new_n19925_;
  assign new_n19927_ = new_n8870_ & new_n19905_;
  assign new_n19928_ = new_n8872_ & new_n19905_;
  assign new_n19929_ = new_n8874_ & new_n19905_;
  assign new_n19930_ = ~new_n19928_ & ~new_n19929_;
  assign new_n19931_ = ~new_n19927_ & new_n19930_;
  assign new_n19932_ = new_n8880_ & new_n19905_;
  assign new_n19933_ = new_n8882_ & new_n19905_;
  assign new_n19934_ = new_n8884_ & new_n19905_;
  assign new_n19935_ = ~new_n19933_ & ~new_n19934_;
  assign new_n19936_ = ~new_n19932_ & new_n19935_;
  assign new_n19937_ = new_n19931_ & new_n19936_;
  assign new_n19938_ = new_n8898_ & new_n19905_;
  assign new_n19939_ = new_n8888_ & new_n19905_;
  assign new_n19940_ = new_n8890_ & new_n19905_;
  assign new_n19941_ = ~new_n19939_ & ~new_n19940_;
  assign new_n19942_ = ~new_n19938_ & new_n19941_;
  assign new_n19943_ = new_n8907_ & new_n19905_;
  assign new_n19944_ = new_n8900_ & new_n19905_;
  assign new_n19945_ = new_n8896_ & new_n19905_;
  assign new_n19946_ = ~new_n19944_ & ~new_n19945_;
  assign new_n19947_ = ~new_n19943_ & new_n19946_;
  assign new_n19948_ = new_n19942_ & new_n19947_;
  assign new_n19949_ = new_n19937_ & new_n19948_;
  assign new_n19950_ = new_n8916_ & new_n19905_;
  assign new_n19951_ = new_n8909_ & new_n19905_;
  assign new_n19952_ = new_n8905_ & new_n19905_;
  assign new_n19953_ = ~new_n19951_ & ~new_n19952_;
  assign new_n19954_ = ~new_n19950_ & new_n19953_;
  assign new_n19955_ = new_n8925_ & new_n19905_;
  assign new_n19956_ = new_n8918_ & new_n19905_;
  assign new_n19957_ = new_n8914_ & new_n19905_;
  assign new_n19958_ = ~new_n19956_ & ~new_n19957_;
  assign new_n19959_ = ~new_n19955_ & new_n19958_;
  assign new_n19960_ = new_n19954_ & new_n19959_;
  assign new_n19961_ = new_n8936_ & new_n19905_;
  assign new_n19962_ = new_n8927_ & new_n19905_;
  assign new_n19963_ = new_n8923_ & new_n19905_;
  assign new_n19964_ = ~new_n19962_ & ~new_n19963_;
  assign new_n19965_ = ~new_n19961_ & new_n19964_;
  assign new_n19966_ = new_n8943_ & new_n19905_;
  assign new_n19967_ = new_n8938_ & new_n19905_;
  assign new_n19968_ = new_n8934_ & new_n19905_;
  assign new_n19969_ = ~new_n19967_ & ~new_n19968_;
  assign new_n19970_ = ~new_n19966_ & new_n19969_;
  assign new_n19971_ = new_n19965_ & new_n19970_;
  assign new_n19972_ = new_n19960_ & new_n19971_;
  assign new_n19973_ = new_n19949_ & new_n19972_;
  assign new_n19974_ = new_n6663_ & new_n16044_;
  assign new_n19975_ = new_n8628_ & new_n19974_;
  assign new_n19976_ = new_n8945_ & new_n19905_;
  assign new_n19977_ = new_n8617_ & new_n19974_;
  assign new_n19978_ = ~new_n19976_ & ~new_n19977_;
  assign new_n19979_ = ~new_n19975_ & new_n19978_;
  assign new_n19980_ = new_n8637_ & new_n19974_;
  assign new_n19981_ = new_n8630_ & new_n19974_;
  assign new_n19982_ = new_n8625_ & new_n19974_;
  assign new_n19983_ = ~new_n19981_ & ~new_n19982_;
  assign new_n19984_ = ~new_n19980_ & new_n19983_;
  assign new_n19985_ = new_n19979_ & new_n19984_;
  assign new_n19986_ = new_n8648_ & new_n19974_;
  assign new_n19987_ = new_n8639_ & new_n19974_;
  assign new_n19988_ = new_n8635_ & new_n19974_;
  assign new_n19989_ = ~new_n19987_ & ~new_n19988_;
  assign new_n19990_ = ~new_n19986_ & new_n19989_;
  assign new_n19991_ = new_n8657_ & new_n19974_;
  assign new_n19992_ = new_n8650_ & new_n19974_;
  assign new_n19993_ = new_n8646_ & new_n19974_;
  assign new_n19994_ = ~new_n19992_ & ~new_n19993_;
  assign new_n19995_ = ~new_n19991_ & new_n19994_;
  assign new_n19996_ = new_n19990_ & new_n19995_;
  assign new_n19997_ = new_n19985_ & new_n19996_;
  assign new_n19998_ = new_n8667_ & new_n19974_;
  assign new_n19999_ = new_n8659_ & new_n19974_;
  assign new_n20000_ = new_n8655_ & new_n19974_;
  assign new_n20001_ = ~new_n19999_ & ~new_n20000_;
  assign new_n20002_ = ~new_n19998_ & new_n20001_;
  assign new_n20003_ = new_n8678_ & new_n19974_;
  assign new_n20004_ = new_n8670_ & new_n19974_;
  assign new_n20005_ = new_n8665_ & new_n19974_;
  assign new_n20006_ = ~new_n20004_ & ~new_n20005_;
  assign new_n20007_ = ~new_n20003_ & new_n20006_;
  assign new_n20008_ = new_n20002_ & new_n20007_;
  assign new_n20009_ = new_n8692_ & new_n19974_;
  assign new_n20010_ = new_n8681_ & new_n19974_;
  assign new_n20011_ = new_n8675_ & new_n19974_;
  assign new_n20012_ = ~new_n20010_ & ~new_n20011_;
  assign new_n20013_ = ~new_n20009_ & new_n20012_;
  assign new_n20014_ = new_n8694_ & new_n19974_;
  assign new_n20015_ = new_n8689_ & new_n19974_;
  assign new_n20016_ = ~new_n20014_ & ~new_n20015_;
  assign new_n20017_ = new_n20013_ & new_n20016_;
  assign new_n20018_ = new_n20008_ & new_n20017_;
  assign new_n20019_ = new_n19997_ & new_n20018_;
  assign new_n20020_ = new_n19973_ & new_n20019_;
  assign new_n20021_ = new_n6663_ & new_n16093_;
  assign new_n20022_ = new_n8617_ & new_n20021_;
  assign new_n20023_ = new_n8699_ & new_n19974_;
  assign new_n20024_ = new_n8701_ & new_n19974_;
  assign new_n20025_ = ~new_n20023_ & ~new_n20024_;
  assign new_n20026_ = ~new_n20022_ & new_n20025_;
  assign new_n20027_ = new_n8625_ & new_n20021_;
  assign new_n20028_ = new_n8628_ & new_n20021_;
  assign new_n20029_ = new_n8630_ & new_n20021_;
  assign new_n20030_ = ~new_n20028_ & ~new_n20029_;
  assign new_n20031_ = ~new_n20027_ & new_n20030_;
  assign new_n20032_ = new_n20026_ & new_n20031_;
  assign new_n20033_ = new_n8635_ & new_n20021_;
  assign new_n20034_ = new_n8637_ & new_n20021_;
  assign new_n20035_ = new_n8639_ & new_n20021_;
  assign new_n20036_ = ~new_n20034_ & ~new_n20035_;
  assign new_n20037_ = ~new_n20033_ & new_n20036_;
  assign new_n20038_ = new_n8646_ & new_n20021_;
  assign new_n20039_ = new_n8648_ & new_n20021_;
  assign new_n20040_ = new_n8650_ & new_n20021_;
  assign new_n20041_ = ~new_n20039_ & ~new_n20040_;
  assign new_n20042_ = ~new_n20038_ & new_n20041_;
  assign new_n20043_ = new_n20037_ & new_n20042_;
  assign new_n20044_ = new_n20032_ & new_n20043_;
  assign new_n20045_ = new_n8655_ & new_n20021_;
  assign new_n20046_ = new_n8657_ & new_n20021_;
  assign new_n20047_ = new_n8659_ & new_n20021_;
  assign new_n20048_ = ~new_n20046_ & ~new_n20047_;
  assign new_n20049_ = ~new_n20045_ & new_n20048_;
  assign new_n20050_ = new_n8665_ & new_n20021_;
  assign new_n20051_ = new_n8667_ & new_n20021_;
  assign new_n20052_ = new_n8670_ & new_n20021_;
  assign new_n20053_ = ~new_n20051_ & ~new_n20052_;
  assign new_n20054_ = ~new_n20050_ & new_n20053_;
  assign new_n20055_ = new_n20049_ & new_n20054_;
  assign new_n20056_ = new_n8675_ & new_n20021_;
  assign new_n20057_ = new_n8678_ & new_n20021_;
  assign new_n20058_ = new_n8681_ & new_n20021_;
  assign new_n20059_ = ~new_n20057_ & ~new_n20058_;
  assign new_n20060_ = ~new_n20056_ & new_n20059_;
  assign new_n20061_ = new_n8692_ & new_n20021_;
  assign new_n20062_ = new_n8694_ & new_n20021_;
  assign new_n20063_ = ~new_n20061_ & ~new_n20062_;
  assign new_n20064_ = new_n20060_ & new_n20063_;
  assign new_n20065_ = new_n20055_ & new_n20064_;
  assign new_n20066_ = new_n20044_ & new_n20065_;
  assign new_n20067_ = new_n8701_ & new_n20021_;
  assign new_n20068_ = new_n8689_ & new_n20021_;
  assign new_n20069_ = new_n8699_ & new_n20021_;
  assign new_n20070_ = ~new_n20068_ & ~new_n20069_;
  assign new_n20071_ = ~new_n20067_ & new_n20070_;
  assign new_n20072_ = new_n6663_ & new_n16151_;
  assign new_n20073_ = new_n8630_ & new_n20072_;
  assign new_n20074_ = new_n8617_ & new_n20072_;
  assign new_n20075_ = new_n8628_ & new_n20072_;
  assign new_n20076_ = ~new_n20074_ & ~new_n20075_;
  assign new_n20077_ = ~new_n20073_ & new_n20076_;
  assign new_n20078_ = new_n20071_ & new_n20077_;
  assign new_n20079_ = new_n8639_ & new_n20072_;
  assign new_n20080_ = new_n8625_ & new_n20072_;
  assign new_n20081_ = new_n8637_ & new_n20072_;
  assign new_n20082_ = ~new_n20080_ & ~new_n20081_;
  assign new_n20083_ = ~new_n20079_ & new_n20082_;
  assign new_n20084_ = new_n8650_ & new_n20072_;
  assign new_n20085_ = new_n8635_ & new_n20072_;
  assign new_n20086_ = new_n8648_ & new_n20072_;
  assign new_n20087_ = ~new_n20085_ & ~new_n20086_;
  assign new_n20088_ = ~new_n20084_ & new_n20087_;
  assign new_n20089_ = new_n20083_ & new_n20088_;
  assign new_n20090_ = new_n20078_ & new_n20089_;
  assign new_n20091_ = new_n8659_ & new_n20072_;
  assign new_n20092_ = new_n8646_ & new_n20072_;
  assign new_n20093_ = new_n8657_ & new_n20072_;
  assign new_n20094_ = ~new_n20092_ & ~new_n20093_;
  assign new_n20095_ = ~new_n20091_ & new_n20094_;
  assign new_n20096_ = new_n8670_ & new_n20072_;
  assign new_n20097_ = new_n8655_ & new_n20072_;
  assign new_n20098_ = new_n8667_ & new_n20072_;
  assign new_n20099_ = ~new_n20097_ & ~new_n20098_;
  assign new_n20100_ = ~new_n20096_ & new_n20099_;
  assign new_n20101_ = new_n20095_ & new_n20100_;
  assign new_n20102_ = new_n8681_ & new_n20072_;
  assign new_n20103_ = new_n8665_ & new_n20072_;
  assign new_n20104_ = new_n8678_ & new_n20072_;
  assign new_n20105_ = ~new_n20103_ & ~new_n20104_;
  assign new_n20106_ = ~new_n20102_ & new_n20105_;
  assign new_n20107_ = new_n8675_ & new_n20072_;
  assign new_n20108_ = new_n8692_ & new_n20072_;
  assign new_n20109_ = ~new_n20107_ & ~new_n20108_;
  assign new_n20110_ = new_n20106_ & new_n20109_;
  assign new_n20111_ = new_n20101_ & new_n20110_;
  assign new_n20112_ = new_n20090_ & new_n20111_;
  assign new_n20113_ = new_n20066_ & new_n20112_;
  assign new_n20114_ = new_n20020_ & new_n20113_;
  assign new_n20115_ = new_n8699_ & new_n20072_;
  assign new_n20116_ = new_n8694_ & new_n20072_;
  assign new_n20117_ = new_n8689_ & new_n20072_;
  assign new_n20118_ = ~new_n20116_ & ~new_n20117_;
  assign new_n20119_ = ~new_n20115_ & new_n20118_;
  assign new_n20120_ = new_n6663_ & new_n16200_;
  assign new_n20121_ = new_n8628_ & new_n20120_;
  assign new_n20122_ = new_n8701_ & new_n20072_;
  assign new_n20123_ = new_n8617_ & new_n20120_;
  assign new_n20124_ = ~new_n20122_ & ~new_n20123_;
  assign new_n20125_ = ~new_n20121_ & new_n20124_;
  assign new_n20126_ = new_n20119_ & new_n20125_;
  assign new_n20127_ = new_n8637_ & new_n20120_;
  assign new_n20128_ = new_n8630_ & new_n20120_;
  assign new_n20129_ = new_n8625_ & new_n20120_;
  assign new_n20130_ = ~new_n20128_ & ~new_n20129_;
  assign new_n20131_ = ~new_n20127_ & new_n20130_;
  assign new_n20132_ = new_n8648_ & new_n20120_;
  assign new_n20133_ = new_n8639_ & new_n20120_;
  assign new_n20134_ = new_n8635_ & new_n20120_;
  assign new_n20135_ = ~new_n20133_ & ~new_n20134_;
  assign new_n20136_ = ~new_n20132_ & new_n20135_;
  assign new_n20137_ = new_n20131_ & new_n20136_;
  assign new_n20138_ = new_n20126_ & new_n20137_;
  assign new_n20139_ = new_n8657_ & new_n20120_;
  assign new_n20140_ = new_n8650_ & new_n20120_;
  assign new_n20141_ = new_n8646_ & new_n20120_;
  assign new_n20142_ = ~new_n20140_ & ~new_n20141_;
  assign new_n20143_ = ~new_n20139_ & new_n20142_;
  assign new_n20144_ = new_n8667_ & new_n20120_;
  assign new_n20145_ = new_n8659_ & new_n20120_;
  assign new_n20146_ = new_n8655_ & new_n20120_;
  assign new_n20147_ = ~new_n20145_ & ~new_n20146_;
  assign new_n20148_ = ~new_n20144_ & new_n20147_;
  assign new_n20149_ = new_n20143_ & new_n20148_;
  assign new_n20150_ = new_n8678_ & new_n20120_;
  assign new_n20151_ = new_n8670_ & new_n20120_;
  assign new_n20152_ = new_n8665_ & new_n20120_;
  assign new_n20153_ = ~new_n20151_ & ~new_n20152_;
  assign new_n20154_ = ~new_n20150_ & new_n20153_;
  assign new_n20155_ = new_n8681_ & new_n20120_;
  assign new_n20156_ = new_n8675_ & new_n20120_;
  assign new_n20157_ = ~new_n20155_ & ~new_n20156_;
  assign new_n20158_ = new_n20154_ & new_n20157_;
  assign new_n20159_ = new_n20149_ & new_n20158_;
  assign new_n20160_ = new_n20138_ & new_n20159_;
  assign new_n20161_ = new_n8689_ & new_n20120_;
  assign new_n20162_ = new_n8692_ & new_n20120_;
  assign new_n20163_ = new_n8694_ & new_n20120_;
  assign new_n20164_ = ~new_n20162_ & ~new_n20163_;
  assign new_n20165_ = ~new_n20161_ & new_n20164_;
  assign new_n20166_ = new_n6663_ & new_n16248_;
  assign new_n20167_ = new_n8845_ & new_n20166_;
  assign new_n20168_ = new_n8699_ & new_n20120_;
  assign new_n20169_ = new_n8701_ & new_n20120_;
  assign new_n20170_ = ~new_n20168_ & ~new_n20169_;
  assign new_n20171_ = ~new_n20167_ & new_n20170_;
  assign new_n20172_ = new_n20165_ & new_n20171_;
  assign new_n20173_ = new_n8851_ & new_n20166_;
  assign new_n20174_ = new_n8853_ & new_n20166_;
  assign new_n20175_ = new_n8855_ & new_n20166_;
  assign new_n20176_ = ~new_n20174_ & ~new_n20175_;
  assign new_n20177_ = ~new_n20173_ & new_n20176_;
  assign new_n20178_ = new_n8862_ & new_n20166_;
  assign new_n20179_ = new_n8864_ & new_n20166_;
  assign new_n20180_ = new_n8866_ & new_n20166_;
  assign new_n20181_ = ~new_n20179_ & ~new_n20180_;
  assign new_n20182_ = ~new_n20178_ & new_n20181_;
  assign new_n20183_ = new_n20177_ & new_n20182_;
  assign new_n20184_ = new_n20172_ & new_n20183_;
  assign new_n20185_ = new_n8870_ & new_n20166_;
  assign new_n20186_ = new_n8872_ & new_n20166_;
  assign new_n20187_ = new_n8874_ & new_n20166_;
  assign new_n20188_ = ~new_n20186_ & ~new_n20187_;
  assign new_n20189_ = ~new_n20185_ & new_n20188_;
  assign new_n20190_ = new_n8880_ & new_n20166_;
  assign new_n20191_ = new_n8882_ & new_n20166_;
  assign new_n20192_ = new_n8884_ & new_n20166_;
  assign new_n20193_ = ~new_n20191_ & ~new_n20192_;
  assign new_n20194_ = ~new_n20190_ & new_n20193_;
  assign new_n20195_ = new_n20189_ & new_n20194_;
  assign new_n20196_ = new_n8898_ & new_n20166_;
  assign new_n20197_ = new_n8888_ & new_n20166_;
  assign new_n20198_ = new_n8890_ & new_n20166_;
  assign new_n20199_ = ~new_n20197_ & ~new_n20198_;
  assign new_n20200_ = ~new_n20196_ & new_n20199_;
  assign new_n20201_ = new_n8900_ & new_n20166_;
  assign new_n20202_ = new_n8896_ & new_n20166_;
  assign new_n20203_ = ~new_n20201_ & ~new_n20202_;
  assign new_n20204_ = new_n20200_ & new_n20203_;
  assign new_n20205_ = new_n20195_ & new_n20204_;
  assign new_n20206_ = new_n20184_ & new_n20205_;
  assign new_n20207_ = new_n20160_ & new_n20206_;
  assign new_n20208_ = new_n8905_ & new_n20166_;
  assign new_n20209_ = new_n8907_ & new_n20166_;
  assign new_n20210_ = new_n8909_ & new_n20166_;
  assign new_n20211_ = ~new_n20209_ & ~new_n20210_;
  assign new_n20212_ = ~new_n20208_ & new_n20211_;
  assign new_n20213_ = new_n8914_ & new_n20166_;
  assign new_n20214_ = new_n8916_ & new_n20166_;
  assign new_n20215_ = new_n8918_ & new_n20166_;
  assign new_n20216_ = ~new_n20214_ & ~new_n20215_;
  assign new_n20217_ = ~new_n20213_ & new_n20216_;
  assign new_n20218_ = new_n20212_ & new_n20217_;
  assign new_n20219_ = new_n8923_ & new_n20166_;
  assign new_n20220_ = new_n8925_ & new_n20166_;
  assign new_n20221_ = new_n8927_ & new_n20166_;
  assign new_n20222_ = ~new_n20220_ & ~new_n20221_;
  assign new_n20223_ = ~new_n20219_ & new_n20222_;
  assign new_n20224_ = new_n8934_ & new_n20166_;
  assign new_n20225_ = new_n8936_ & new_n20166_;
  assign new_n20226_ = new_n8938_ & new_n20166_;
  assign new_n20227_ = ~new_n20225_ & ~new_n20226_;
  assign new_n20228_ = ~new_n20224_ & new_n20227_;
  assign new_n20229_ = new_n20223_ & new_n20228_;
  assign new_n20230_ = new_n20218_ & new_n20229_;
  assign new_n20231_ = new_n6672_ & new_n16311_;
  assign new_n20232_ = new_n8617_ & new_n20231_;
  assign new_n20233_ = new_n8943_ & new_n20166_;
  assign new_n20234_ = new_n8945_ & new_n20166_;
  assign new_n20235_ = ~new_n20233_ & ~new_n20234_;
  assign new_n20236_ = ~new_n20232_ & new_n20235_;
  assign new_n20237_ = new_n8625_ & new_n20231_;
  assign new_n20238_ = new_n8628_ & new_n20231_;
  assign new_n20239_ = new_n8630_ & new_n20231_;
  assign new_n20240_ = ~new_n20238_ & ~new_n20239_;
  assign new_n20241_ = ~new_n20237_ & new_n20240_;
  assign new_n20242_ = new_n20236_ & new_n20241_;
  assign new_n20243_ = new_n8635_ & new_n20231_;
  assign new_n20244_ = new_n8637_ & new_n20231_;
  assign new_n20245_ = new_n8639_ & new_n20231_;
  assign new_n20246_ = ~new_n20244_ & ~new_n20245_;
  assign new_n20247_ = ~new_n20243_ & new_n20246_;
  assign new_n20248_ = new_n8648_ & new_n20231_;
  assign new_n20249_ = new_n8650_ & new_n20231_;
  assign new_n20250_ = ~new_n20248_ & ~new_n20249_;
  assign new_n20251_ = new_n20247_ & new_n20250_;
  assign new_n20252_ = new_n20242_ & new_n20251_;
  assign new_n20253_ = new_n20230_ & new_n20252_;
  assign new_n20254_ = new_n8659_ & new_n20231_;
  assign new_n20255_ = new_n8646_ & new_n20231_;
  assign new_n20256_ = new_n8657_ & new_n20231_;
  assign new_n20257_ = ~new_n20255_ & ~new_n20256_;
  assign new_n20258_ = ~new_n20254_ & new_n20257_;
  assign new_n20259_ = new_n8670_ & new_n20231_;
  assign new_n20260_ = new_n8655_ & new_n20231_;
  assign new_n20261_ = new_n8667_ & new_n20231_;
  assign new_n20262_ = ~new_n20260_ & ~new_n20261_;
  assign new_n20263_ = ~new_n20259_ & new_n20262_;
  assign new_n20264_ = new_n20258_ & new_n20263_;
  assign new_n20265_ = new_n8681_ & new_n20231_;
  assign new_n20266_ = new_n8665_ & new_n20231_;
  assign new_n20267_ = new_n8678_ & new_n20231_;
  assign new_n20268_ = ~new_n20266_ & ~new_n20267_;
  assign new_n20269_ = ~new_n20265_ & new_n20268_;
  assign new_n20270_ = new_n8694_ & new_n20231_;
  assign new_n20271_ = new_n8675_ & new_n20231_;
  assign new_n20272_ = new_n8692_ & new_n20231_;
  assign new_n20273_ = ~new_n20271_ & ~new_n20272_;
  assign new_n20274_ = ~new_n20270_ & new_n20273_;
  assign new_n20275_ = new_n20269_ & new_n20274_;
  assign new_n20276_ = new_n20264_ & new_n20275_;
  assign new_n20277_ = new_n8701_ & new_n20231_;
  assign new_n20278_ = new_n8689_ & new_n20231_;
  assign new_n20279_ = new_n8699_ & new_n20231_;
  assign new_n20280_ = ~new_n20278_ & ~new_n20279_;
  assign new_n20281_ = ~new_n20277_ & new_n20280_;
  assign new_n20282_ = new_n6672_ & new_n16360_;
  assign new_n20283_ = new_n8630_ & new_n20282_;
  assign new_n20284_ = new_n8617_ & new_n20282_;
  assign new_n20285_ = new_n8628_ & new_n20282_;
  assign new_n20286_ = ~new_n20284_ & ~new_n20285_;
  assign new_n20287_ = ~new_n20283_ & new_n20286_;
  assign new_n20288_ = new_n20281_ & new_n20287_;
  assign new_n20289_ = new_n8639_ & new_n20282_;
  assign new_n20290_ = new_n8625_ & new_n20282_;
  assign new_n20291_ = new_n8637_ & new_n20282_;
  assign new_n20292_ = ~new_n20290_ & ~new_n20291_;
  assign new_n20293_ = ~new_n20289_ & new_n20292_;
  assign new_n20294_ = new_n8635_ & new_n20282_;
  assign new_n20295_ = new_n8648_ & new_n20282_;
  assign new_n20296_ = ~new_n20294_ & ~new_n20295_;
  assign new_n20297_ = new_n20293_ & new_n20296_;
  assign new_n20298_ = new_n20288_ & new_n20297_;
  assign new_n20299_ = new_n20276_ & new_n20298_;
  assign new_n20300_ = new_n20253_ & new_n20299_;
  assign new_n20301_ = new_n20207_ & new_n20300_;
  assign new_n20302_ = new_n20114_ & new_n20301_;
  assign new_n20303_ = new_n8657_ & new_n20282_;
  assign new_n20304_ = new_n8650_ & new_n20282_;
  assign new_n20305_ = new_n8646_ & new_n20282_;
  assign new_n20306_ = ~new_n20304_ & ~new_n20305_;
  assign new_n20307_ = ~new_n20303_ & new_n20306_;
  assign new_n20308_ = new_n8667_ & new_n20282_;
  assign new_n20309_ = new_n8659_ & new_n20282_;
  assign new_n20310_ = new_n8655_ & new_n20282_;
  assign new_n20311_ = ~new_n20309_ & ~new_n20310_;
  assign new_n20312_ = ~new_n20308_ & new_n20311_;
  assign new_n20313_ = new_n20307_ & new_n20312_;
  assign new_n20314_ = new_n8678_ & new_n20282_;
  assign new_n20315_ = new_n8670_ & new_n20282_;
  assign new_n20316_ = new_n8665_ & new_n20282_;
  assign new_n20317_ = ~new_n20315_ & ~new_n20316_;
  assign new_n20318_ = ~new_n20314_ & new_n20317_;
  assign new_n20319_ = new_n8692_ & new_n20282_;
  assign new_n20320_ = new_n8681_ & new_n20282_;
  assign new_n20321_ = new_n8675_ & new_n20282_;
  assign new_n20322_ = ~new_n20320_ & ~new_n20321_;
  assign new_n20323_ = ~new_n20319_ & new_n20322_;
  assign new_n20324_ = new_n20318_ & new_n20323_;
  assign new_n20325_ = new_n20313_ & new_n20324_;
  assign new_n20326_ = new_n8699_ & new_n20282_;
  assign new_n20327_ = new_n8694_ & new_n20282_;
  assign new_n20328_ = new_n8689_ & new_n20282_;
  assign new_n20329_ = ~new_n20327_ & ~new_n20328_;
  assign new_n20330_ = ~new_n20326_ & new_n20329_;
  assign new_n20331_ = new_n6672_ & new_n16414_;
  assign new_n20332_ = new_n8628_ & new_n20331_;
  assign new_n20333_ = new_n8701_ & new_n20282_;
  assign new_n20334_ = new_n8617_ & new_n20331_;
  assign new_n20335_ = ~new_n20333_ & ~new_n20334_;
  assign new_n20336_ = ~new_n20332_ & new_n20335_;
  assign new_n20337_ = new_n20330_ & new_n20336_;
  assign new_n20338_ = new_n8637_ & new_n20331_;
  assign new_n20339_ = new_n8630_ & new_n20331_;
  assign new_n20340_ = new_n8625_ & new_n20331_;
  assign new_n20341_ = ~new_n20339_ & ~new_n20340_;
  assign new_n20342_ = ~new_n20338_ & new_n20341_;
  assign new_n20343_ = new_n8639_ & new_n20331_;
  assign new_n20344_ = new_n8635_ & new_n20331_;
  assign new_n20345_ = ~new_n20343_ & ~new_n20344_;
  assign new_n20346_ = new_n20342_ & new_n20345_;
  assign new_n20347_ = new_n20337_ & new_n20346_;
  assign new_n20348_ = new_n20325_ & new_n20347_;
  assign new_n20349_ = new_n8646_ & new_n20331_;
  assign new_n20350_ = new_n8648_ & new_n20331_;
  assign new_n20351_ = new_n8650_ & new_n20331_;
  assign new_n20352_ = ~new_n20350_ & ~new_n20351_;
  assign new_n20353_ = ~new_n20349_ & new_n20352_;
  assign new_n20354_ = new_n8655_ & new_n20331_;
  assign new_n20355_ = new_n8657_ & new_n20331_;
  assign new_n20356_ = new_n8659_ & new_n20331_;
  assign new_n20357_ = ~new_n20355_ & ~new_n20356_;
  assign new_n20358_ = ~new_n20354_ & new_n20357_;
  assign new_n20359_ = new_n20353_ & new_n20358_;
  assign new_n20360_ = new_n8665_ & new_n20331_;
  assign new_n20361_ = new_n8667_ & new_n20331_;
  assign new_n20362_ = new_n8670_ & new_n20331_;
  assign new_n20363_ = ~new_n20361_ & ~new_n20362_;
  assign new_n20364_ = ~new_n20360_ & new_n20363_;
  assign new_n20365_ = new_n8675_ & new_n20331_;
  assign new_n20366_ = new_n8678_ & new_n20331_;
  assign new_n20367_ = new_n8681_ & new_n20331_;
  assign new_n20368_ = ~new_n20366_ & ~new_n20367_;
  assign new_n20369_ = ~new_n20365_ & new_n20368_;
  assign new_n20370_ = new_n20364_ & new_n20369_;
  assign new_n20371_ = new_n20359_ & new_n20370_;
  assign new_n20372_ = new_n8689_ & new_n20331_;
  assign new_n20373_ = new_n8692_ & new_n20331_;
  assign new_n20374_ = new_n8694_ & new_n20331_;
  assign new_n20375_ = ~new_n20373_ & ~new_n20374_;
  assign new_n20376_ = ~new_n20372_ & new_n20375_;
  assign new_n20377_ = new_n6672_ & new_n16462_;
  assign new_n20378_ = new_n8617_ & new_n20377_;
  assign new_n20379_ = new_n8699_ & new_n20331_;
  assign new_n20380_ = new_n8701_ & new_n20331_;
  assign new_n20381_ = ~new_n20379_ & ~new_n20380_;
  assign new_n20382_ = ~new_n20378_ & new_n20381_;
  assign new_n20383_ = new_n20376_ & new_n20382_;
  assign new_n20384_ = new_n8625_ & new_n20377_;
  assign new_n20385_ = new_n8628_ & new_n20377_;
  assign new_n20386_ = new_n8630_ & new_n20377_;
  assign new_n20387_ = ~new_n20385_ & ~new_n20386_;
  assign new_n20388_ = ~new_n20384_ & new_n20387_;
  assign new_n20389_ = new_n8637_ & new_n20377_;
  assign new_n20390_ = new_n8639_ & new_n20377_;
  assign new_n20391_ = ~new_n20389_ & ~new_n20390_;
  assign new_n20392_ = new_n20388_ & new_n20391_;
  assign new_n20393_ = new_n20383_ & new_n20392_;
  assign new_n20394_ = new_n20371_ & new_n20393_;
  assign new_n20395_ = new_n20348_ & new_n20394_;
  assign new_n20396_ = new_n8650_ & new_n20377_;
  assign new_n20397_ = new_n8635_ & new_n20377_;
  assign new_n20398_ = new_n8648_ & new_n20377_;
  assign new_n20399_ = ~new_n20397_ & ~new_n20398_;
  assign new_n20400_ = ~new_n20396_ & new_n20399_;
  assign new_n20401_ = new_n8659_ & new_n20377_;
  assign new_n20402_ = new_n8646_ & new_n20377_;
  assign new_n20403_ = new_n8657_ & new_n20377_;
  assign new_n20404_ = ~new_n20402_ & ~new_n20403_;
  assign new_n20405_ = ~new_n20401_ & new_n20404_;
  assign new_n20406_ = new_n20400_ & new_n20405_;
  assign new_n20407_ = new_n8670_ & new_n20377_;
  assign new_n20408_ = new_n8655_ & new_n20377_;
  assign new_n20409_ = new_n8667_ & new_n20377_;
  assign new_n20410_ = ~new_n20408_ & ~new_n20409_;
  assign new_n20411_ = ~new_n20407_ & new_n20410_;
  assign new_n20412_ = new_n8681_ & new_n20377_;
  assign new_n20413_ = new_n8665_ & new_n20377_;
  assign new_n20414_ = new_n8678_ & new_n20377_;
  assign new_n20415_ = ~new_n20413_ & ~new_n20414_;
  assign new_n20416_ = ~new_n20412_ & new_n20415_;
  assign new_n20417_ = new_n20411_ & new_n20416_;
  assign new_n20418_ = new_n20406_ & new_n20417_;
  assign new_n20419_ = new_n8694_ & new_n20377_;
  assign new_n20420_ = new_n8675_ & new_n20377_;
  assign new_n20421_ = new_n8692_ & new_n20377_;
  assign new_n20422_ = ~new_n20420_ & ~new_n20421_;
  assign new_n20423_ = ~new_n20419_ & new_n20422_;
  assign new_n20424_ = new_n8701_ & new_n20377_;
  assign new_n20425_ = new_n8689_ & new_n20377_;
  assign new_n20426_ = new_n8699_ & new_n20377_;
  assign new_n20427_ = ~new_n20425_ & ~new_n20426_;
  assign new_n20428_ = ~new_n20424_ & new_n20427_;
  assign new_n20429_ = new_n20423_ & new_n20428_;
  assign new_n20430_ = new_n6672_ & new_n16509_;
  assign new_n20431_ = new_n8855_ & new_n20430_;
  assign new_n20432_ = new_n8845_ & new_n20430_;
  assign new_n20433_ = new_n8853_ & new_n20430_;
  assign new_n20434_ = ~new_n20432_ & ~new_n20433_;
  assign new_n20435_ = ~new_n20431_ & new_n20434_;
  assign new_n20436_ = new_n8851_ & new_n20430_;
  assign new_n20437_ = new_n8864_ & new_n20430_;
  assign new_n20438_ = ~new_n20436_ & ~new_n20437_;
  assign new_n20439_ = new_n20435_ & new_n20438_;
  assign new_n20440_ = new_n20429_ & new_n20439_;
  assign new_n20441_ = new_n20418_ & new_n20440_;
  assign new_n20442_ = new_n8872_ & new_n20430_;
  assign new_n20443_ = new_n8866_ & new_n20430_;
  assign new_n20444_ = new_n8862_ & new_n20430_;
  assign new_n20445_ = ~new_n20443_ & ~new_n20444_;
  assign new_n20446_ = ~new_n20442_ & new_n20445_;
  assign new_n20447_ = new_n8882_ & new_n20430_;
  assign new_n20448_ = new_n8874_ & new_n20430_;
  assign new_n20449_ = new_n8870_ & new_n20430_;
  assign new_n20450_ = ~new_n20448_ & ~new_n20449_;
  assign new_n20451_ = ~new_n20447_ & new_n20450_;
  assign new_n20452_ = new_n20446_ & new_n20451_;
  assign new_n20453_ = new_n8888_ & new_n20430_;
  assign new_n20454_ = new_n8884_ & new_n20430_;
  assign new_n20455_ = new_n8880_ & new_n20430_;
  assign new_n20456_ = ~new_n20454_ & ~new_n20455_;
  assign new_n20457_ = ~new_n20453_ & new_n20456_;
  assign new_n20458_ = new_n8900_ & new_n20430_;
  assign new_n20459_ = new_n8890_ & new_n20430_;
  assign new_n20460_ = new_n8898_ & new_n20430_;
  assign new_n20461_ = ~new_n20459_ & ~new_n20460_;
  assign new_n20462_ = ~new_n20458_ & new_n20461_;
  assign new_n20463_ = new_n20457_ & new_n20462_;
  assign new_n20464_ = new_n20452_ & new_n20463_;
  assign new_n20465_ = new_n8909_ & new_n20430_;
  assign new_n20466_ = new_n8896_ & new_n20430_;
  assign new_n20467_ = new_n8907_ & new_n20430_;
  assign new_n20468_ = ~new_n20466_ & ~new_n20467_;
  assign new_n20469_ = ~new_n20465_ & new_n20468_;
  assign new_n20470_ = new_n8918_ & new_n20430_;
  assign new_n20471_ = new_n8905_ & new_n20430_;
  assign new_n20472_ = new_n8916_ & new_n20430_;
  assign new_n20473_ = ~new_n20471_ & ~new_n20472_;
  assign new_n20474_ = ~new_n20470_ & new_n20473_;
  assign new_n20475_ = new_n20469_ & new_n20474_;
  assign new_n20476_ = new_n8927_ & new_n20430_;
  assign new_n20477_ = new_n8914_ & new_n20430_;
  assign new_n20478_ = new_n8925_ & new_n20430_;
  assign new_n20479_ = ~new_n20477_ & ~new_n20478_;
  assign new_n20480_ = ~new_n20476_ & new_n20479_;
  assign new_n20481_ = new_n8923_ & new_n20430_;
  assign new_n20482_ = new_n8936_ & new_n20430_;
  assign new_n20483_ = ~new_n20481_ & ~new_n20482_;
  assign new_n20484_ = new_n20480_ & new_n20483_;
  assign new_n20485_ = new_n20475_ & new_n20484_;
  assign new_n20486_ = new_n20464_ & new_n20485_;
  assign new_n20487_ = new_n20441_ & new_n20486_;
  assign new_n20488_ = new_n20395_ & new_n20487_;
  assign new_n20489_ = new_n8943_ & new_n20430_;
  assign new_n20490_ = new_n8938_ & new_n20430_;
  assign new_n20491_ = new_n8934_ & new_n20430_;
  assign new_n20492_ = ~new_n20490_ & ~new_n20491_;
  assign new_n20493_ = ~new_n20489_ & new_n20492_;
  assign new_n20494_ = new_n6672_ & new_n16575_;
  assign new_n20495_ = new_n8628_ & new_n20494_;
  assign new_n20496_ = new_n8945_ & new_n20430_;
  assign new_n20497_ = new_n8617_ & new_n20494_;
  assign new_n20498_ = ~new_n20496_ & ~new_n20497_;
  assign new_n20499_ = ~new_n20495_ & new_n20498_;
  assign new_n20500_ = new_n20493_ & new_n20499_;
  assign new_n20501_ = new_n8637_ & new_n20494_;
  assign new_n20502_ = new_n8630_ & new_n20494_;
  assign new_n20503_ = new_n8625_ & new_n20494_;
  assign new_n20504_ = ~new_n20502_ & ~new_n20503_;
  assign new_n20505_ = ~new_n20501_ & new_n20504_;
  assign new_n20506_ = new_n8648_ & new_n20494_;
  assign new_n20507_ = new_n8639_ & new_n20494_;
  assign new_n20508_ = new_n8635_ & new_n20494_;
  assign new_n20509_ = ~new_n20507_ & ~new_n20508_;
  assign new_n20510_ = ~new_n20506_ & new_n20509_;
  assign new_n20511_ = new_n20505_ & new_n20510_;
  assign new_n20512_ = new_n20500_ & new_n20511_;
  assign new_n20513_ = new_n8657_ & new_n20494_;
  assign new_n20514_ = new_n8650_ & new_n20494_;
  assign new_n20515_ = new_n8646_ & new_n20494_;
  assign new_n20516_ = ~new_n20514_ & ~new_n20515_;
  assign new_n20517_ = ~new_n20513_ & new_n20516_;
  assign new_n20518_ = new_n8667_ & new_n20494_;
  assign new_n20519_ = new_n8659_ & new_n20494_;
  assign new_n20520_ = new_n8655_ & new_n20494_;
  assign new_n20521_ = ~new_n20519_ & ~new_n20520_;
  assign new_n20522_ = ~new_n20518_ & new_n20521_;
  assign new_n20523_ = new_n20517_ & new_n20522_;
  assign new_n20524_ = new_n8678_ & new_n20494_;
  assign new_n20525_ = new_n8670_ & new_n20494_;
  assign new_n20526_ = new_n8665_ & new_n20494_;
  assign new_n20527_ = ~new_n20525_ & ~new_n20526_;
  assign new_n20528_ = ~new_n20524_ & new_n20527_;
  assign new_n20529_ = new_n8681_ & new_n20494_;
  assign new_n20530_ = new_n8675_ & new_n20494_;
  assign new_n20531_ = ~new_n20529_ & ~new_n20530_;
  assign new_n20532_ = new_n20528_ & new_n20531_;
  assign new_n20533_ = new_n20523_ & new_n20532_;
  assign new_n20534_ = new_n20512_ & new_n20533_;
  assign new_n20535_ = new_n8689_ & new_n20494_;
  assign new_n20536_ = new_n8692_ & new_n20494_;
  assign new_n20537_ = new_n8694_ & new_n20494_;
  assign new_n20538_ = ~new_n20536_ & ~new_n20537_;
  assign new_n20539_ = ~new_n20535_ & new_n20538_;
  assign new_n20540_ = new_n6672_ & new_n16631_;
  assign new_n20541_ = new_n8617_ & new_n20540_;
  assign new_n20542_ = new_n8699_ & new_n20494_;
  assign new_n20543_ = new_n8701_ & new_n20494_;
  assign new_n20544_ = ~new_n20542_ & ~new_n20543_;
  assign new_n20545_ = ~new_n20541_ & new_n20544_;
  assign new_n20546_ = new_n20539_ & new_n20545_;
  assign new_n20547_ = new_n8625_ & new_n20540_;
  assign new_n20548_ = new_n8628_ & new_n20540_;
  assign new_n20549_ = new_n8630_ & new_n20540_;
  assign new_n20550_ = ~new_n20548_ & ~new_n20549_;
  assign new_n20551_ = ~new_n20547_ & new_n20550_;
  assign new_n20552_ = new_n8635_ & new_n20540_;
  assign new_n20553_ = new_n8637_ & new_n20540_;
  assign new_n20554_ = new_n8639_ & new_n20540_;
  assign new_n20555_ = ~new_n20553_ & ~new_n20554_;
  assign new_n20556_ = ~new_n20552_ & new_n20555_;
  assign new_n20557_ = new_n20551_ & new_n20556_;
  assign new_n20558_ = new_n20546_ & new_n20557_;
  assign new_n20559_ = new_n8646_ & new_n20540_;
  assign new_n20560_ = new_n8648_ & new_n20540_;
  assign new_n20561_ = new_n8650_ & new_n20540_;
  assign new_n20562_ = ~new_n20560_ & ~new_n20561_;
  assign new_n20563_ = ~new_n20559_ & new_n20562_;
  assign new_n20564_ = new_n8655_ & new_n20540_;
  assign new_n20565_ = new_n8657_ & new_n20540_;
  assign new_n20566_ = new_n8659_ & new_n20540_;
  assign new_n20567_ = ~new_n20565_ & ~new_n20566_;
  assign new_n20568_ = ~new_n20564_ & new_n20567_;
  assign new_n20569_ = new_n20563_ & new_n20568_;
  assign new_n20570_ = new_n8665_ & new_n20540_;
  assign new_n20571_ = new_n8667_ & new_n20540_;
  assign new_n20572_ = new_n8670_ & new_n20540_;
  assign new_n20573_ = ~new_n20571_ & ~new_n20572_;
  assign new_n20574_ = ~new_n20570_ & new_n20573_;
  assign new_n20575_ = new_n8678_ & new_n20540_;
  assign new_n20576_ = new_n8681_ & new_n20540_;
  assign new_n20577_ = ~new_n20575_ & ~new_n20576_;
  assign new_n20578_ = new_n20574_ & new_n20577_;
  assign new_n20579_ = new_n20569_ & new_n20578_;
  assign new_n20580_ = new_n20558_ & new_n20579_;
  assign new_n20581_ = new_n20534_ & new_n20580_;
  assign new_n20582_ = new_n8694_ & new_n20540_;
  assign new_n20583_ = new_n8675_ & new_n20540_;
  assign new_n20584_ = new_n8692_ & new_n20540_;
  assign new_n20585_ = ~new_n20583_ & ~new_n20584_;
  assign new_n20586_ = ~new_n20582_ & new_n20585_;
  assign new_n20587_ = new_n8701_ & new_n20540_;
  assign new_n20588_ = new_n8689_ & new_n20540_;
  assign new_n20589_ = new_n8699_ & new_n20540_;
  assign new_n20590_ = ~new_n20588_ & ~new_n20589_;
  assign new_n20591_ = ~new_n20587_ & new_n20590_;
  assign new_n20592_ = new_n20586_ & new_n20591_;
  assign new_n20593_ = new_n6672_ & new_n16678_;
  assign new_n20594_ = new_n8630_ & new_n20593_;
  assign new_n20595_ = new_n8617_ & new_n20593_;
  assign new_n20596_ = new_n8628_ & new_n20593_;
  assign new_n20597_ = ~new_n20595_ & ~new_n20596_;
  assign new_n20598_ = ~new_n20594_ & new_n20597_;
  assign new_n20599_ = new_n8639_ & new_n20593_;
  assign new_n20600_ = new_n8625_ & new_n20593_;
  assign new_n20601_ = new_n8637_ & new_n20593_;
  assign new_n20602_ = ~new_n20600_ & ~new_n20601_;
  assign new_n20603_ = ~new_n20599_ & new_n20602_;
  assign new_n20604_ = new_n20598_ & new_n20603_;
  assign new_n20605_ = new_n20592_ & new_n20604_;
  assign new_n20606_ = new_n8650_ & new_n20593_;
  assign new_n20607_ = new_n8635_ & new_n20593_;
  assign new_n20608_ = new_n8648_ & new_n20593_;
  assign new_n20609_ = ~new_n20607_ & ~new_n20608_;
  assign new_n20610_ = ~new_n20606_ & new_n20609_;
  assign new_n20611_ = new_n8659_ & new_n20593_;
  assign new_n20612_ = new_n8646_ & new_n20593_;
  assign new_n20613_ = new_n8657_ & new_n20593_;
  assign new_n20614_ = ~new_n20612_ & ~new_n20613_;
  assign new_n20615_ = ~new_n20611_ & new_n20614_;
  assign new_n20616_ = new_n20610_ & new_n20615_;
  assign new_n20617_ = new_n8670_ & new_n20593_;
  assign new_n20618_ = new_n8655_ & new_n20593_;
  assign new_n20619_ = new_n8667_ & new_n20593_;
  assign new_n20620_ = ~new_n20618_ & ~new_n20619_;
  assign new_n20621_ = ~new_n20617_ & new_n20620_;
  assign new_n20622_ = new_n8665_ & new_n20593_;
  assign new_n20623_ = new_n8678_ & new_n20593_;
  assign new_n20624_ = ~new_n20622_ & ~new_n20623_;
  assign new_n20625_ = new_n20621_ & new_n20624_;
  assign new_n20626_ = new_n20616_ & new_n20625_;
  assign new_n20627_ = new_n20605_ & new_n20626_;
  assign new_n20628_ = new_n8692_ & new_n20593_;
  assign new_n20629_ = new_n8681_ & new_n20593_;
  assign new_n20630_ = new_n8675_ & new_n20593_;
  assign new_n20631_ = ~new_n20629_ & ~new_n20630_;
  assign new_n20632_ = ~new_n20628_ & new_n20631_;
  assign new_n20633_ = new_n8699_ & new_n20593_;
  assign new_n20634_ = new_n8694_ & new_n20593_;
  assign new_n20635_ = new_n8689_ & new_n20593_;
  assign new_n20636_ = ~new_n20634_ & ~new_n20635_;
  assign new_n20637_ = ~new_n20633_ & new_n20636_;
  assign new_n20638_ = new_n20632_ & new_n20637_;
  assign new_n20639_ = new_n6672_ & new_n16727_;
  assign new_n20640_ = new_n8628_ & new_n20639_;
  assign new_n20641_ = new_n8701_ & new_n20593_;
  assign new_n20642_ = new_n8617_ & new_n20639_;
  assign new_n20643_ = ~new_n20641_ & ~new_n20642_;
  assign new_n20644_ = ~new_n20640_ & new_n20643_;
  assign new_n20645_ = new_n8637_ & new_n20639_;
  assign new_n20646_ = new_n8630_ & new_n20639_;
  assign new_n20647_ = new_n8625_ & new_n20639_;
  assign new_n20648_ = ~new_n20646_ & ~new_n20647_;
  assign new_n20649_ = ~new_n20645_ & new_n20648_;
  assign new_n20650_ = new_n20644_ & new_n20649_;
  assign new_n20651_ = new_n20638_ & new_n20650_;
  assign new_n20652_ = new_n8648_ & new_n20639_;
  assign new_n20653_ = new_n8639_ & new_n20639_;
  assign new_n20654_ = new_n8635_ & new_n20639_;
  assign new_n20655_ = ~new_n20653_ & ~new_n20654_;
  assign new_n20656_ = ~new_n20652_ & new_n20655_;
  assign new_n20657_ = new_n8657_ & new_n20639_;
  assign new_n20658_ = new_n8650_ & new_n20639_;
  assign new_n20659_ = new_n8646_ & new_n20639_;
  assign new_n20660_ = ~new_n20658_ & ~new_n20659_;
  assign new_n20661_ = ~new_n20657_ & new_n20660_;
  assign new_n20662_ = new_n20656_ & new_n20661_;
  assign new_n20663_ = new_n8667_ & new_n20639_;
  assign new_n20664_ = new_n8659_ & new_n20639_;
  assign new_n20665_ = new_n8655_ & new_n20639_;
  assign new_n20666_ = ~new_n20664_ & ~new_n20665_;
  assign new_n20667_ = ~new_n20663_ & new_n20666_;
  assign new_n20668_ = new_n8670_ & new_n20639_;
  assign new_n20669_ = new_n8665_ & new_n20639_;
  assign new_n20670_ = ~new_n20668_ & ~new_n20669_;
  assign new_n20671_ = new_n20667_ & new_n20670_;
  assign new_n20672_ = new_n20662_ & new_n20671_;
  assign new_n20673_ = new_n20651_ & new_n20672_;
  assign new_n20674_ = new_n20627_ & new_n20673_;
  assign new_n20675_ = new_n20581_ & new_n20674_;
  assign new_n20676_ = new_n20488_ & new_n20675_;
  assign new_n20677_ = new_n20302_ & new_n20676_;
  assign new_n20678_ = new_n19926_ & new_n20677_;
  assign new_n20679_ = new_n8675_ & new_n20639_;
  assign new_n20680_ = new_n8678_ & new_n20639_;
  assign new_n20681_ = new_n8681_ & new_n20639_;
  assign new_n20682_ = ~new_n20680_ & ~new_n20681_;
  assign new_n20683_ = ~new_n20679_ & new_n20682_;
  assign new_n20684_ = new_n8689_ & new_n20639_;
  assign new_n20685_ = new_n8692_ & new_n20639_;
  assign new_n20686_ = new_n8694_ & new_n20639_;
  assign new_n20687_ = ~new_n20685_ & ~new_n20686_;
  assign new_n20688_ = ~new_n20684_ & new_n20687_;
  assign new_n20689_ = new_n20683_ & new_n20688_;
  assign new_n20690_ = new_n6672_ & new_n16779_;
  assign new_n20691_ = new_n8845_ & new_n20690_;
  assign new_n20692_ = new_n8699_ & new_n20639_;
  assign new_n20693_ = new_n8701_ & new_n20639_;
  assign new_n20694_ = ~new_n20692_ & ~new_n20693_;
  assign new_n20695_ = ~new_n20691_ & new_n20694_;
  assign new_n20696_ = new_n8851_ & new_n20690_;
  assign new_n20697_ = new_n8853_ & new_n20690_;
  assign new_n20698_ = new_n8855_ & new_n20690_;
  assign new_n20699_ = ~new_n20697_ & ~new_n20698_;
  assign new_n20700_ = ~new_n20696_ & new_n20699_;
  assign new_n20701_ = new_n20695_ & new_n20700_;
  assign new_n20702_ = new_n20689_ & new_n20701_;
  assign new_n20703_ = new_n8862_ & new_n20690_;
  assign new_n20704_ = new_n8864_ & new_n20690_;
  assign new_n20705_ = new_n8866_ & new_n20690_;
  assign new_n20706_ = ~new_n20704_ & ~new_n20705_;
  assign new_n20707_ = ~new_n20703_ & new_n20706_;
  assign new_n20708_ = new_n8870_ & new_n20690_;
  assign new_n20709_ = new_n8872_ & new_n20690_;
  assign new_n20710_ = new_n8874_ & new_n20690_;
  assign new_n20711_ = ~new_n20709_ & ~new_n20710_;
  assign new_n20712_ = ~new_n20708_ & new_n20711_;
  assign new_n20713_ = new_n20707_ & new_n20712_;
  assign new_n20714_ = new_n8880_ & new_n20690_;
  assign new_n20715_ = new_n8882_ & new_n20690_;
  assign new_n20716_ = new_n8884_ & new_n20690_;
  assign new_n20717_ = ~new_n20715_ & ~new_n20716_;
  assign new_n20718_ = ~new_n20714_ & new_n20717_;
  assign new_n20719_ = new_n8898_ & new_n20690_;
  assign new_n20720_ = new_n8888_ & new_n20690_;
  assign new_n20721_ = new_n8890_ & new_n20690_;
  assign new_n20722_ = ~new_n20720_ & ~new_n20721_;
  assign new_n20723_ = ~new_n20719_ & new_n20722_;
  assign new_n20724_ = new_n20718_ & new_n20723_;
  assign new_n20725_ = new_n20713_ & new_n20724_;
  assign new_n20726_ = new_n20702_ & new_n20725_;
  assign new_n20727_ = new_n8907_ & new_n20690_;
  assign new_n20728_ = new_n8900_ & new_n20690_;
  assign new_n20729_ = new_n8896_ & new_n20690_;
  assign new_n20730_ = ~new_n20728_ & ~new_n20729_;
  assign new_n20731_ = ~new_n20727_ & new_n20730_;
  assign new_n20732_ = new_n8916_ & new_n20690_;
  assign new_n20733_ = new_n8909_ & new_n20690_;
  assign new_n20734_ = new_n8905_ & new_n20690_;
  assign new_n20735_ = ~new_n20733_ & ~new_n20734_;
  assign new_n20736_ = ~new_n20732_ & new_n20735_;
  assign new_n20737_ = new_n20731_ & new_n20736_;
  assign new_n20738_ = new_n8925_ & new_n20690_;
  assign new_n20739_ = new_n8918_ & new_n20690_;
  assign new_n20740_ = new_n8914_ & new_n20690_;
  assign new_n20741_ = ~new_n20739_ & ~new_n20740_;
  assign new_n20742_ = ~new_n20738_ & new_n20741_;
  assign new_n20743_ = new_n8936_ & new_n20690_;
  assign new_n20744_ = new_n8927_ & new_n20690_;
  assign new_n20745_ = new_n8923_ & new_n20690_;
  assign new_n20746_ = ~new_n20744_ & ~new_n20745_;
  assign new_n20747_ = ~new_n20743_ & new_n20746_;
  assign new_n20748_ = new_n20742_ & new_n20747_;
  assign new_n20749_ = new_n20737_ & new_n20748_;
  assign new_n20750_ = new_n8943_ & new_n20690_;
  assign new_n20751_ = new_n8938_ & new_n20690_;
  assign new_n20752_ = new_n8934_ & new_n20690_;
  assign new_n20753_ = ~new_n20751_ & ~new_n20752_;
  assign new_n20754_ = ~new_n20750_ & new_n20753_;
  assign new_n20755_ = new_n6693_ & new_n16845_;
  assign new_n20756_ = new_n9720_ & new_n20755_;
  assign new_n20757_ = new_n8945_ & new_n20690_;
  assign new_n20758_ = new_n9718_ & new_n20755_;
  assign new_n20759_ = ~new_n20757_ & ~new_n20758_;
  assign new_n20760_ = ~new_n20756_ & new_n20759_;
  assign new_n20761_ = new_n20754_ & new_n20760_;
  assign new_n20762_ = new_n9731_ & new_n20755_;
  assign new_n20763_ = new_n9716_ & new_n20755_;
  assign new_n20764_ = new_n9729_ & new_n20755_;
  assign new_n20765_ = ~new_n20763_ & ~new_n20764_;
  assign new_n20766_ = ~new_n20762_ & new_n20765_;
  assign new_n20767_ = new_n9727_ & new_n20755_;
  assign new_n20768_ = new_n9737_ & new_n20755_;
  assign new_n20769_ = ~new_n20767_ & ~new_n20768_;
  assign new_n20770_ = new_n20766_ & new_n20769_;
  assign new_n20771_ = new_n20761_ & new_n20770_;
  assign new_n20772_ = new_n20749_ & new_n20771_;
  assign new_n20773_ = new_n20726_ & new_n20772_;
  assign new_n20774_ = new_n9746_ & new_n20755_;
  assign new_n20775_ = new_n9739_ & new_n20755_;
  assign new_n20776_ = new_n9735_ & new_n20755_;
  assign new_n20777_ = ~new_n20775_ & ~new_n20776_;
  assign new_n20778_ = ~new_n20774_ & new_n20777_;
  assign new_n20779_ = new_n9753_ & new_n20755_;
  assign new_n20780_ = new_n9748_ & new_n20755_;
  assign new_n20781_ = new_n9744_ & new_n20755_;
  assign new_n20782_ = ~new_n20780_ & ~new_n20781_;
  assign new_n20783_ = ~new_n20779_ & new_n20782_;
  assign new_n20784_ = new_n20778_ & new_n20783_;
  assign new_n20785_ = new_n9765_ & new_n20755_;
  assign new_n20786_ = new_n9755_ & new_n20755_;
  assign new_n20787_ = new_n9763_ & new_n20755_;
  assign new_n20788_ = ~new_n20786_ & ~new_n20787_;
  assign new_n20789_ = ~new_n20785_ & new_n20788_;
  assign new_n20790_ = new_n9773_ & new_n20755_;
  assign new_n20791_ = new_n9761_ & new_n20755_;
  assign new_n20792_ = new_n9771_ & new_n20755_;
  assign new_n20793_ = ~new_n20791_ & ~new_n20792_;
  assign new_n20794_ = ~new_n20790_ & new_n20793_;
  assign new_n20795_ = new_n20789_ & new_n20794_;
  assign new_n20796_ = new_n20784_ & new_n20795_;
  assign new_n20797_ = new_n9783_ & new_n20755_;
  assign new_n20798_ = new_n9769_ & new_n20755_;
  assign new_n20799_ = new_n9781_ & new_n20755_;
  assign new_n20800_ = ~new_n20798_ & ~new_n20799_;
  assign new_n20801_ = ~new_n20797_ & new_n20800_;
  assign new_n20802_ = new_n9792_ & new_n20755_;
  assign new_n20803_ = new_n9779_ & new_n20755_;
  assign new_n20804_ = new_n9790_ & new_n20755_;
  assign new_n20805_ = ~new_n20803_ & ~new_n20804_;
  assign new_n20806_ = ~new_n20802_ & new_n20805_;
  assign new_n20807_ = new_n20801_ & new_n20806_;
  assign new_n20808_ = new_n9803_ & new_n20755_;
  assign new_n20809_ = new_n9788_ & new_n20755_;
  assign new_n20810_ = new_n9801_ & new_n20755_;
  assign new_n20811_ = ~new_n20809_ & ~new_n20810_;
  assign new_n20812_ = ~new_n20808_ & new_n20811_;
  assign new_n20813_ = new_n9799_ & new_n20755_;
  assign new_n20814_ = new_n9809_ & new_n20755_;
  assign new_n20815_ = ~new_n20813_ & ~new_n20814_;
  assign new_n20816_ = new_n20812_ & new_n20815_;
  assign new_n20817_ = new_n20807_ & new_n20816_;
  assign new_n20818_ = new_n20796_ & new_n20817_;
  assign new_n20819_ = new_n6693_ & new_n16908_;
  assign new_n20820_ = new_n9819_ & new_n20819_;
  assign new_n20821_ = new_n9811_ & new_n20755_;
  assign new_n20822_ = new_n9807_ & new_n20755_;
  assign new_n20823_ = ~new_n20821_ & ~new_n20822_;
  assign new_n20824_ = ~new_n20820_ & new_n20823_;
  assign new_n20825_ = new_n9825_ & new_n20819_;
  assign new_n20826_ = new_n9821_ & new_n20819_;
  assign new_n20827_ = new_n9817_ & new_n20819_;
  assign new_n20828_ = ~new_n20826_ & ~new_n20827_;
  assign new_n20829_ = ~new_n20825_ & new_n20828_;
  assign new_n20830_ = new_n20824_ & new_n20829_;
  assign new_n20831_ = new_n9844_ & new_n20819_;
  assign new_n20832_ = new_n9828_ & new_n20819_;
  assign new_n20833_ = new_n9842_ & new_n20819_;
  assign new_n20834_ = ~new_n20832_ & ~new_n20833_;
  assign new_n20835_ = ~new_n20831_ & new_n20834_;
  assign new_n20836_ = new_n9852_ & new_n20819_;
  assign new_n20837_ = new_n9840_ & new_n20819_;
  assign new_n20838_ = new_n9850_ & new_n20819_;
  assign new_n20839_ = ~new_n20837_ & ~new_n20838_;
  assign new_n20840_ = ~new_n20836_ & new_n20839_;
  assign new_n20841_ = new_n20835_ & new_n20840_;
  assign new_n20842_ = new_n20830_ & new_n20841_;
  assign new_n20843_ = new_n9862_ & new_n20819_;
  assign new_n20844_ = new_n9848_ & new_n20819_;
  assign new_n20845_ = new_n9860_ & new_n20819_;
  assign new_n20846_ = ~new_n20844_ & ~new_n20845_;
  assign new_n20847_ = ~new_n20843_ & new_n20846_;
  assign new_n20848_ = new_n9870_ & new_n20819_;
  assign new_n20849_ = new_n9858_ & new_n20819_;
  assign new_n20850_ = new_n9868_ & new_n20819_;
  assign new_n20851_ = ~new_n20849_ & ~new_n20850_;
  assign new_n20852_ = ~new_n20848_ & new_n20851_;
  assign new_n20853_ = new_n20847_ & new_n20852_;
  assign new_n20854_ = new_n9880_ & new_n20819_;
  assign new_n20855_ = new_n9866_ & new_n20819_;
  assign new_n20856_ = new_n9878_ & new_n20819_;
  assign new_n20857_ = ~new_n20855_ & ~new_n20856_;
  assign new_n20858_ = ~new_n20854_ & new_n20857_;
  assign new_n20859_ = new_n9876_ & new_n20819_;
  assign new_n20860_ = new_n9887_ & new_n20819_;
  assign new_n20861_ = ~new_n20859_ & ~new_n20860_;
  assign new_n20862_ = new_n20858_ & new_n20861_;
  assign new_n20863_ = new_n20853_ & new_n20862_;
  assign new_n20864_ = new_n20842_ & new_n20863_;
  assign new_n20865_ = new_n20818_ & new_n20864_;
  assign new_n20866_ = new_n20773_ & new_n20865_;
  assign new_n20867_ = new_n9897_ & new_n20819_;
  assign new_n20868_ = new_n9889_ & new_n20819_;
  assign new_n20869_ = new_n9885_ & new_n20819_;
  assign new_n20870_ = ~new_n20868_ & ~new_n20869_;
  assign new_n20871_ = ~new_n20867_ & new_n20870_;
  assign new_n20872_ = new_n9906_ & new_n20819_;
  assign new_n20873_ = new_n9899_ & new_n20819_;
  assign new_n20874_ = new_n9895_ & new_n20819_;
  assign new_n20875_ = ~new_n20873_ & ~new_n20874_;
  assign new_n20876_ = ~new_n20872_ & new_n20875_;
  assign new_n20877_ = new_n20871_ & new_n20876_;
  assign new_n20878_ = new_n9917_ & new_n20819_;
  assign new_n20879_ = new_n9908_ & new_n20819_;
  assign new_n20880_ = new_n9904_ & new_n20819_;
  assign new_n20881_ = ~new_n20879_ & ~new_n20880_;
  assign new_n20882_ = ~new_n20878_ & new_n20881_;
  assign new_n20883_ = new_n6693_ & new_n16978_;
  assign new_n20884_ = new_n9926_ & new_n20883_;
  assign new_n20885_ = new_n9919_ & new_n20819_;
  assign new_n20886_ = new_n9915_ & new_n20819_;
  assign new_n20887_ = ~new_n20885_ & ~new_n20886_;
  assign new_n20888_ = ~new_n20884_ & new_n20887_;
  assign new_n20889_ = new_n20882_ & new_n20888_;
  assign new_n20890_ = new_n20877_ & new_n20889_;
  assign new_n20891_ = new_n9936_ & new_n20883_;
  assign new_n20892_ = new_n9928_ & new_n20883_;
  assign new_n20893_ = new_n9924_ & new_n20883_;
  assign new_n20894_ = ~new_n20892_ & ~new_n20893_;
  assign new_n20895_ = ~new_n20891_ & new_n20894_;
  assign new_n20896_ = new_n9944_ & new_n20883_;
  assign new_n20897_ = new_n9938_ & new_n20883_;
  assign new_n20898_ = new_n9934_ & new_n20883_;
  assign new_n20899_ = ~new_n20897_ & ~new_n20898_;
  assign new_n20900_ = ~new_n20896_ & new_n20899_;
  assign new_n20901_ = new_n20895_ & new_n20900_;
  assign new_n20902_ = new_n9954_ & new_n20883_;
  assign new_n20903_ = new_n9946_ & new_n20883_;
  assign new_n20904_ = new_n9942_ & new_n20883_;
  assign new_n20905_ = ~new_n20903_ & ~new_n20904_;
  assign new_n20906_ = ~new_n20902_ & new_n20905_;
  assign new_n20907_ = new_n9956_ & new_n20883_;
  assign new_n20908_ = new_n9952_ & new_n20883_;
  assign new_n20909_ = ~new_n20907_ & ~new_n20908_;
  assign new_n20910_ = new_n20906_ & new_n20909_;
  assign new_n20911_ = new_n20901_ & new_n20910_;
  assign new_n20912_ = new_n20890_ & new_n20911_;
  assign new_n20913_ = new_n9961_ & new_n20883_;
  assign new_n20914_ = new_n9963_ & new_n20883_;
  assign new_n20915_ = new_n9965_ & new_n20883_;
  assign new_n20916_ = ~new_n20914_ & ~new_n20915_;
  assign new_n20917_ = ~new_n20913_ & new_n20916_;
  assign new_n20918_ = new_n9970_ & new_n20883_;
  assign new_n20919_ = new_n9972_ & new_n20883_;
  assign new_n20920_ = new_n9974_ & new_n20883_;
  assign new_n20921_ = ~new_n20919_ & ~new_n20920_;
  assign new_n20922_ = ~new_n20918_ & new_n20921_;
  assign new_n20923_ = new_n20917_ & new_n20922_;
  assign new_n20924_ = new_n9990_ & new_n20883_;
  assign new_n20925_ = new_n9978_ & new_n20883_;
  assign new_n20926_ = new_n9980_ & new_n20883_;
  assign new_n20927_ = ~new_n20925_ & ~new_n20926_;
  assign new_n20928_ = ~new_n20924_ & new_n20927_;
  assign new_n20929_ = new_n9999_ & new_n20883_;
  assign new_n20930_ = new_n9992_ & new_n20883_;
  assign new_n20931_ = new_n9988_ & new_n20883_;
  assign new_n20932_ = ~new_n20930_ & ~new_n20931_;
  assign new_n20933_ = ~new_n20929_ & new_n20932_;
  assign new_n20934_ = new_n20928_ & new_n20933_;
  assign new_n20935_ = new_n20923_ & new_n20934_;
  assign new_n20936_ = new_n10009_ & new_n20883_;
  assign new_n20937_ = new_n10001_ & new_n20883_;
  assign new_n20938_ = new_n9997_ & new_n20883_;
  assign new_n20939_ = ~new_n20937_ & ~new_n20938_;
  assign new_n20940_ = ~new_n20936_ & new_n20939_;
  assign new_n20941_ = new_n10017_ & new_n20883_;
  assign new_n20942_ = new_n10011_ & new_n20883_;
  assign new_n20943_ = new_n10007_ & new_n20883_;
  assign new_n20944_ = ~new_n20942_ & ~new_n20943_;
  assign new_n20945_ = ~new_n20941_ & new_n20944_;
  assign new_n20946_ = new_n20940_ & new_n20945_;
  assign new_n20947_ = new_n10028_ & new_n20883_;
  assign new_n20948_ = new_n10019_ & new_n20883_;
  assign new_n20949_ = new_n10015_ & new_n20883_;
  assign new_n20950_ = ~new_n20948_ & ~new_n20949_;
  assign new_n20951_ = ~new_n20947_ & new_n20950_;
  assign new_n20952_ = new_n10030_ & new_n20883_;
  assign new_n20953_ = new_n10026_ & new_n20883_;
  assign new_n20954_ = ~new_n20952_ & ~new_n20953_;
  assign new_n20955_ = new_n20951_ & new_n20954_;
  assign new_n20956_ = new_n20946_ & new_n20955_;
  assign new_n20957_ = new_n20935_ & new_n20956_;
  assign new_n20958_ = new_n20912_ & new_n20957_;
  assign new_n20959_ = new_n10035_ & new_n20883_;
  assign new_n20960_ = new_n10037_ & new_n20883_;
  assign new_n20961_ = new_n10039_ & new_n20883_;
  assign new_n20962_ = ~new_n20960_ & ~new_n20961_;
  assign new_n20963_ = ~new_n20959_ & new_n20962_;
  assign new_n20964_ = new_n10044_ & new_n20883_;
  assign new_n20965_ = new_n10046_ & new_n20883_;
  assign new_n20966_ = new_n10048_ & new_n20883_;
  assign new_n20967_ = ~new_n20965_ & ~new_n20966_;
  assign new_n20968_ = ~new_n20964_ & new_n20967_;
  assign new_n20969_ = new_n20963_ & new_n20968_;
  assign new_n20970_ = new_n10063_ & new_n20883_;
  assign new_n20971_ = new_n10052_ & new_n20883_;
  assign new_n20972_ = new_n10054_ & new_n20883_;
  assign new_n20973_ = ~new_n20971_ & ~new_n20972_;
  assign new_n20974_ = ~new_n20970_ & new_n20973_;
  assign new_n20975_ = new_n10071_ & new_n20883_;
  assign new_n20976_ = new_n10065_ & new_n20883_;
  assign new_n20977_ = new_n10061_ & new_n20883_;
  assign new_n20978_ = ~new_n20976_ & ~new_n20977_;
  assign new_n20979_ = ~new_n20975_ & new_n20978_;
  assign new_n20980_ = new_n20974_ & new_n20979_;
  assign new_n20981_ = new_n20969_ & new_n20980_;
  assign new_n20982_ = new_n10080_ & new_n20883_;
  assign new_n20983_ = new_n10073_ & new_n20883_;
  assign new_n20984_ = new_n10069_ & new_n20883_;
  assign new_n20985_ = ~new_n20983_ & ~new_n20984_;
  assign new_n20986_ = ~new_n20982_ & new_n20985_;
  assign new_n20987_ = new_n10089_ & new_n20883_;
  assign new_n20988_ = new_n10082_ & new_n20883_;
  assign new_n20989_ = new_n10078_ & new_n20883_;
  assign new_n20990_ = ~new_n20988_ & ~new_n20989_;
  assign new_n20991_ = ~new_n20987_ & new_n20990_;
  assign new_n20992_ = new_n20986_ & new_n20991_;
  assign new_n20993_ = new_n10100_ & new_n20883_;
  assign new_n20994_ = new_n10091_ & new_n20883_;
  assign new_n20995_ = new_n10087_ & new_n20883_;
  assign new_n20996_ = ~new_n20994_ & ~new_n20995_;
  assign new_n20997_ = ~new_n20993_ & new_n20996_;
  assign new_n20998_ = new_n10102_ & new_n20883_;
  assign new_n20999_ = new_n10098_ & new_n20883_;
  assign new_n21000_ = ~new_n20998_ & ~new_n20999_;
  assign new_n21001_ = new_n20997_ & new_n21000_;
  assign new_n21002_ = new_n20992_ & new_n21001_;
  assign new_n21003_ = new_n20981_ & new_n21002_;
  assign new_n21004_ = new_n10107_ & new_n20883_;
  assign new_n21005_ = new_n10109_ & new_n20883_;
  assign new_n21006_ = new_n10111_ & new_n20883_;
  assign new_n21007_ = ~new_n21005_ & ~new_n21006_;
  assign new_n21008_ = ~new_n21004_ & new_n21007_;
  assign new_n21009_ = new_n10116_ & new_n20883_;
  assign new_n21010_ = new_n10118_ & new_n20883_;
  assign new_n21011_ = new_n10120_ & new_n20883_;
  assign new_n21012_ = ~new_n21010_ & ~new_n21011_;
  assign new_n21013_ = ~new_n21009_ & new_n21012_;
  assign new_n21014_ = new_n21008_ & new_n21013_;
  assign new_n21015_ = new_n255_ & new_n8627_;
  assign new_n21016_ = new_n15779_ & new_n21015_;
  assign new_n21017_ = new_n229_ & new_n8616_;
  assign new_n21018_ = new_n15779_ & new_n21017_;
  assign new_n21019_ = new_n251_ & new_n8616_;
  assign new_n21020_ = new_n15779_ & new_n21019_;
  assign new_n21021_ = ~new_n21018_ & ~new_n21020_;
  assign new_n21022_ = ~new_n21016_ & new_n21021_;
  assign new_n21023_ = ~A269 & new_n151_;
  assign new_n21024_ = new_n8634_ & new_n21023_;
  assign new_n21025_ = new_n15779_ & new_n21024_;
  assign new_n21026_ = new_n246_ & new_n8627_;
  assign new_n21027_ = new_n15779_ & new_n21026_;
  assign new_n21028_ = ~A269 & new_n161_;
  assign new_n21029_ = new_n8634_ & new_n21028_;
  assign new_n21030_ = new_n15779_ & new_n21029_;
  assign new_n21031_ = ~new_n21027_ & ~new_n21030_;
  assign new_n21032_ = ~new_n21025_ & new_n21031_;
  assign new_n21033_ = new_n21022_ & new_n21032_;
  assign new_n21034_ = new_n21014_ & new_n21033_;
  assign new_n21035_ = A268 & new_n161_;
  assign new_n21036_ = new_n8634_ & new_n21035_;
  assign new_n21037_ = new_n15779_ & new_n21036_;
  assign new_n21038_ = ~A269 & new_n174_;
  assign new_n21039_ = new_n8634_ & new_n21038_;
  assign new_n21040_ = new_n15779_ & new_n21039_;
  assign new_n21041_ = ~A269 & new_n179_;
  assign new_n21042_ = new_n8634_ & new_n21041_;
  assign new_n21043_ = new_n15779_ & new_n21042_;
  assign new_n21044_ = ~new_n21040_ & ~new_n21043_;
  assign new_n21045_ = ~new_n21037_ & new_n21044_;
  assign new_n21046_ = A268 & new_n179_;
  assign new_n21047_ = new_n8634_ & new_n21046_;
  assign new_n21048_ = new_n15779_ & new_n21047_;
  assign new_n21049_ = A268 & new_n151_;
  assign new_n21050_ = new_n8634_ & new_n21049_;
  assign new_n21051_ = new_n15779_ & new_n21050_;
  assign new_n21052_ = A268 & new_n174_;
  assign new_n21053_ = new_n8634_ & new_n21052_;
  assign new_n21054_ = new_n15779_ & new_n21053_;
  assign new_n21055_ = ~new_n21051_ & ~new_n21054_;
  assign new_n21056_ = ~new_n21048_ & new_n21055_;
  assign new_n21057_ = new_n21045_ & new_n21056_;
  assign new_n21058_ = new_n8654_ & new_n21038_;
  assign new_n21059_ = new_n15779_ & new_n21058_;
  assign new_n21060_ = new_n8654_ & new_n21028_;
  assign new_n21061_ = new_n15779_ & new_n21060_;
  assign new_n21062_ = new_n8654_ & new_n21023_;
  assign new_n21063_ = new_n15779_ & new_n21062_;
  assign new_n21064_ = ~new_n21061_ & ~new_n21063_;
  assign new_n21065_ = ~new_n21059_ & new_n21064_;
  assign new_n21066_ = new_n8654_ & new_n21041_;
  assign new_n21067_ = new_n15779_ & new_n21066_;
  assign new_n21068_ = new_n8654_ & new_n21035_;
  assign new_n21069_ = new_n15779_ & new_n21068_;
  assign new_n21070_ = ~new_n21067_ & ~new_n21069_;
  assign new_n21071_ = new_n21065_ & new_n21070_;
  assign new_n21072_ = new_n21057_ & new_n21071_;
  assign new_n21073_ = new_n21034_ & new_n21072_;
  assign new_n21074_ = new_n21003_ & new_n21073_;
  assign new_n21075_ = new_n20958_ & new_n21074_;
  assign new_n21076_ = new_n20866_ & new_n21075_;
  assign new_n21077_ = new_n8654_ & new_n21046_;
  assign new_n21078_ = new_n15779_ & new_n21077_;
  assign new_n21079_ = new_n8654_ & new_n21049_;
  assign new_n21080_ = new_n15779_ & new_n21079_;
  assign new_n21081_ = new_n8654_ & new_n21052_;
  assign new_n21082_ = new_n15779_ & new_n21081_;
  assign new_n21083_ = ~new_n21080_ & ~new_n21082_;
  assign new_n21084_ = ~new_n21078_ & new_n21083_;
  assign new_n21085_ = new_n255_ & new_n8664_;
  assign new_n21086_ = new_n15779_ & new_n21085_;
  assign new_n21087_ = new_n229_ & new_n8669_;
  assign new_n21088_ = new_n15779_ & new_n21087_;
  assign new_n21089_ = new_n251_ & new_n8669_;
  assign new_n21090_ = new_n15779_ & new_n21089_;
  assign new_n21091_ = ~new_n21088_ & ~new_n21090_;
  assign new_n21092_ = ~new_n21086_ & new_n21091_;
  assign new_n21093_ = new_n21084_ & new_n21092_;
  assign new_n21094_ = new_n251_ & new_n8677_;
  assign new_n21095_ = new_n15779_ & new_n21094_;
  assign new_n21096_ = new_n246_ & new_n8664_;
  assign new_n21097_ = new_n15779_ & new_n21096_;
  assign new_n21098_ = new_n229_ & new_n8677_;
  assign new_n21099_ = new_n15779_ & new_n21098_;
  assign new_n21100_ = ~new_n21097_ & ~new_n21099_;
  assign new_n21101_ = ~new_n21095_ & new_n21100_;
  assign new_n21102_ = new_n229_ & new_n8674_;
  assign new_n21103_ = new_n15779_ & new_n21102_;
  assign new_n21104_ = new_n255_ & new_n8680_;
  assign new_n21105_ = new_n15779_ & new_n21104_;
  assign new_n21106_ = new_n246_ & new_n8680_;
  assign new_n21107_ = new_n15779_ & new_n21106_;
  assign new_n21108_ = ~new_n21105_ & ~new_n21107_;
  assign new_n21109_ = ~new_n21103_ & new_n21108_;
  assign new_n21110_ = new_n21101_ & new_n21109_;
  assign new_n21111_ = new_n21093_ & new_n21110_;
  assign new_n21112_ = new_n246_ & new_n8691_;
  assign new_n21113_ = new_n15779_ & new_n21112_;
  assign new_n21114_ = new_n251_ & new_n8674_;
  assign new_n21115_ = new_n15779_ & new_n21114_;
  assign new_n21116_ = new_n255_ & new_n8691_;
  assign new_n21117_ = new_n15779_ & new_n21116_;
  assign new_n21118_ = ~new_n21115_ & ~new_n21117_;
  assign new_n21119_ = ~new_n21113_ & new_n21118_;
  assign new_n21120_ = new_n15831_ & new_n21015_;
  assign new_n21121_ = new_n15831_ & new_n21017_;
  assign new_n21122_ = new_n15831_ & new_n21019_;
  assign new_n21123_ = ~new_n21121_ & ~new_n21122_;
  assign new_n21124_ = ~new_n21120_ & new_n21123_;
  assign new_n21125_ = new_n21119_ & new_n21124_;
  assign new_n21126_ = new_n15831_ & new_n21024_;
  assign new_n21127_ = new_n15831_ & new_n21026_;
  assign new_n21128_ = new_n15831_ & new_n21029_;
  assign new_n21129_ = ~new_n21127_ & ~new_n21128_;
  assign new_n21130_ = ~new_n21126_ & new_n21129_;
  assign new_n21131_ = new_n15831_ & new_n21036_;
  assign new_n21132_ = new_n15831_ & new_n21039_;
  assign new_n21133_ = new_n15831_ & new_n21042_;
  assign new_n21134_ = ~new_n21132_ & ~new_n21133_;
  assign new_n21135_ = ~new_n21131_ & new_n21134_;
  assign new_n21136_ = new_n21130_ & new_n21135_;
  assign new_n21137_ = new_n21125_ & new_n21136_;
  assign new_n21138_ = new_n21111_ & new_n21137_;
  assign new_n21139_ = new_n15831_ & new_n21047_;
  assign new_n21140_ = new_n15831_ & new_n21050_;
  assign new_n21141_ = new_n15831_ & new_n21053_;
  assign new_n21142_ = ~new_n21140_ & ~new_n21141_;
  assign new_n21143_ = ~new_n21139_ & new_n21142_;
  assign new_n21144_ = new_n15831_ & new_n21058_;
  assign new_n21145_ = new_n15831_ & new_n21060_;
  assign new_n21146_ = new_n15831_ & new_n21062_;
  assign new_n21147_ = ~new_n21145_ & ~new_n21146_;
  assign new_n21148_ = ~new_n21144_ & new_n21147_;
  assign new_n21149_ = new_n21143_ & new_n21148_;
  assign new_n21150_ = new_n15831_ & new_n21079_;
  assign new_n21151_ = new_n15831_ & new_n21066_;
  assign new_n21152_ = new_n15831_ & new_n21068_;
  assign new_n21153_ = ~new_n21151_ & ~new_n21152_;
  assign new_n21154_ = ~new_n21150_ & new_n21153_;
  assign new_n21155_ = new_n15831_ & new_n21087_;
  assign new_n21156_ = new_n15831_ & new_n21081_;
  assign new_n21157_ = new_n15831_ & new_n21077_;
  assign new_n21158_ = ~new_n21156_ & ~new_n21157_;
  assign new_n21159_ = ~new_n21155_ & new_n21158_;
  assign new_n21160_ = new_n21154_ & new_n21159_;
  assign new_n21161_ = new_n21149_ & new_n21160_;
  assign new_n21162_ = new_n15831_ & new_n21096_;
  assign new_n21163_ = new_n15831_ & new_n21089_;
  assign new_n21164_ = new_n15831_ & new_n21085_;
  assign new_n21165_ = ~new_n21163_ & ~new_n21164_;
  assign new_n21166_ = ~new_n21162_ & new_n21165_;
  assign new_n21167_ = new_n15831_ & new_n21104_;
  assign new_n21168_ = new_n15831_ & new_n21098_;
  assign new_n21169_ = new_n15831_ & new_n21094_;
  assign new_n21170_ = ~new_n21168_ & ~new_n21169_;
  assign new_n21171_ = ~new_n21167_ & new_n21170_;
  assign new_n21172_ = new_n21166_ & new_n21171_;
  assign new_n21173_ = new_n15831_ & new_n21114_;
  assign new_n21174_ = new_n15831_ & new_n21106_;
  assign new_n21175_ = new_n15831_ & new_n21102_;
  assign new_n21176_ = ~new_n21174_ & ~new_n21175_;
  assign new_n21177_ = ~new_n21173_ & new_n21176_;
  assign new_n21178_ = new_n15831_ & new_n21116_;
  assign new_n21179_ = new_n15831_ & new_n21112_;
  assign new_n21180_ = ~new_n21178_ & ~new_n21179_;
  assign new_n21181_ = new_n21177_ & new_n21180_;
  assign new_n21182_ = new_n21172_ & new_n21181_;
  assign new_n21183_ = new_n21161_ & new_n21182_;
  assign new_n21184_ = new_n21138_ & new_n21183_;
  assign new_n21185_ = new_n15879_ & new_n21015_;
  assign new_n21186_ = new_n15879_ & new_n21017_;
  assign new_n21187_ = new_n15879_ & new_n21019_;
  assign new_n21188_ = ~new_n21186_ & ~new_n21187_;
  assign new_n21189_ = ~new_n21185_ & new_n21188_;
  assign new_n21190_ = new_n15879_ & new_n21024_;
  assign new_n21191_ = new_n15879_ & new_n21026_;
  assign new_n21192_ = new_n15879_ & new_n21029_;
  assign new_n21193_ = ~new_n21191_ & ~new_n21192_;
  assign new_n21194_ = ~new_n21190_ & new_n21193_;
  assign new_n21195_ = new_n21189_ & new_n21194_;
  assign new_n21196_ = new_n15879_ & new_n21036_;
  assign new_n21197_ = new_n15879_ & new_n21039_;
  assign new_n21198_ = new_n15879_ & new_n21042_;
  assign new_n21199_ = ~new_n21197_ & ~new_n21198_;
  assign new_n21200_ = ~new_n21196_ & new_n21199_;
  assign new_n21201_ = new_n15879_ & new_n21047_;
  assign new_n21202_ = new_n15879_ & new_n21050_;
  assign new_n21203_ = new_n15879_ & new_n21053_;
  assign new_n21204_ = ~new_n21202_ & ~new_n21203_;
  assign new_n21205_ = ~new_n21201_ & new_n21204_;
  assign new_n21206_ = new_n21200_ & new_n21205_;
  assign new_n21207_ = new_n21195_ & new_n21206_;
  assign new_n21208_ = new_n15879_ & new_n21058_;
  assign new_n21209_ = new_n15879_ & new_n21060_;
  assign new_n21210_ = new_n15879_ & new_n21062_;
  assign new_n21211_ = ~new_n21209_ & ~new_n21210_;
  assign new_n21212_ = ~new_n21208_ & new_n21211_;
  assign new_n21213_ = new_n15879_ & new_n21079_;
  assign new_n21214_ = new_n15879_ & new_n21066_;
  assign new_n21215_ = new_n15879_ & new_n21068_;
  assign new_n21216_ = ~new_n21214_ & ~new_n21215_;
  assign new_n21217_ = ~new_n21213_ & new_n21216_;
  assign new_n21218_ = new_n21212_ & new_n21217_;
  assign new_n21219_ = new_n15879_ & new_n21087_;
  assign new_n21220_ = new_n15879_ & new_n21081_;
  assign new_n21221_ = new_n15879_ & new_n21077_;
  assign new_n21222_ = ~new_n21220_ & ~new_n21221_;
  assign new_n21223_ = ~new_n21219_ & new_n21222_;
  assign new_n21224_ = new_n15879_ & new_n21089_;
  assign new_n21225_ = new_n15879_ & new_n21085_;
  assign new_n21226_ = ~new_n21224_ & ~new_n21225_;
  assign new_n21227_ = new_n21223_ & new_n21226_;
  assign new_n21228_ = new_n21218_ & new_n21227_;
  assign new_n21229_ = new_n21207_ & new_n21228_;
  assign new_n21230_ = new_n15879_ & new_n21094_;
  assign new_n21231_ = new_n15879_ & new_n21096_;
  assign new_n21232_ = new_n15879_ & new_n21098_;
  assign new_n21233_ = ~new_n21231_ & ~new_n21232_;
  assign new_n21234_ = ~new_n21230_ & new_n21233_;
  assign new_n21235_ = new_n15879_ & new_n21102_;
  assign new_n21236_ = new_n15879_ & new_n21104_;
  assign new_n21237_ = new_n15879_ & new_n21106_;
  assign new_n21238_ = ~new_n21236_ & ~new_n21237_;
  assign new_n21239_ = ~new_n21235_ & new_n21238_;
  assign new_n21240_ = new_n21234_ & new_n21239_;
  assign new_n21241_ = new_n15879_ & new_n21112_;
  assign new_n21242_ = new_n15879_ & new_n21114_;
  assign new_n21243_ = new_n15879_ & new_n21116_;
  assign new_n21244_ = ~new_n21242_ & ~new_n21243_;
  assign new_n21245_ = ~new_n21241_ & new_n21244_;
  assign new_n21246_ = new_n15926_ & new_n21015_;
  assign new_n21247_ = new_n15926_ & new_n21017_;
  assign new_n21248_ = new_n15926_ & new_n21019_;
  assign new_n21249_ = ~new_n21247_ & ~new_n21248_;
  assign new_n21250_ = ~new_n21246_ & new_n21249_;
  assign new_n21251_ = new_n21245_ & new_n21250_;
  assign new_n21252_ = new_n21240_ & new_n21251_;
  assign new_n21253_ = new_n15926_ & new_n21024_;
  assign new_n21254_ = new_n15926_ & new_n21026_;
  assign new_n21255_ = new_n15926_ & new_n21029_;
  assign new_n21256_ = ~new_n21254_ & ~new_n21255_;
  assign new_n21257_ = ~new_n21253_ & new_n21256_;
  assign new_n21258_ = new_n15926_ & new_n21036_;
  assign new_n21259_ = new_n15926_ & new_n21039_;
  assign new_n21260_ = new_n15926_ & new_n21042_;
  assign new_n21261_ = ~new_n21259_ & ~new_n21260_;
  assign new_n21262_ = ~new_n21258_ & new_n21261_;
  assign new_n21263_ = new_n21257_ & new_n21262_;
  assign new_n21264_ = new_n15926_ & new_n21047_;
  assign new_n21265_ = new_n15926_ & new_n21050_;
  assign new_n21266_ = new_n15926_ & new_n21053_;
  assign new_n21267_ = ~new_n21265_ & ~new_n21266_;
  assign new_n21268_ = ~new_n21264_ & new_n21267_;
  assign new_n21269_ = new_n15926_ & new_n21060_;
  assign new_n21270_ = new_n15926_ & new_n21062_;
  assign new_n21271_ = ~new_n21269_ & ~new_n21270_;
  assign new_n21272_ = new_n21268_ & new_n21271_;
  assign new_n21273_ = new_n21263_ & new_n21272_;
  assign new_n21274_ = new_n21252_ & new_n21273_;
  assign new_n21275_ = new_n21229_ & new_n21274_;
  assign new_n21276_ = new_n21184_ & new_n21275_;
  assign new_n21277_ = new_n15926_ & new_n21068_;
  assign new_n21278_ = new_n15926_ & new_n21058_;
  assign new_n21279_ = new_n15926_ & new_n21066_;
  assign new_n21280_ = ~new_n21278_ & ~new_n21279_;
  assign new_n21281_ = ~new_n21277_ & new_n21280_;
  assign new_n21282_ = new_n15926_ & new_n21077_;
  assign new_n21283_ = new_n15926_ & new_n21079_;
  assign new_n21284_ = new_n15926_ & new_n21081_;
  assign new_n21285_ = ~new_n21283_ & ~new_n21284_;
  assign new_n21286_ = ~new_n21282_ & new_n21285_;
  assign new_n21287_ = new_n21281_ & new_n21286_;
  assign new_n21288_ = new_n15926_ & new_n21085_;
  assign new_n21289_ = new_n15926_ & new_n21087_;
  assign new_n21290_ = new_n15926_ & new_n21089_;
  assign new_n21291_ = ~new_n21289_ & ~new_n21290_;
  assign new_n21292_ = ~new_n21288_ & new_n21291_;
  assign new_n21293_ = new_n15926_ & new_n21094_;
  assign new_n21294_ = new_n15926_ & new_n21096_;
  assign new_n21295_ = new_n15926_ & new_n21098_;
  assign new_n21296_ = ~new_n21294_ & ~new_n21295_;
  assign new_n21297_ = ~new_n21293_ & new_n21296_;
  assign new_n21298_ = new_n21292_ & new_n21297_;
  assign new_n21299_ = new_n21287_ & new_n21298_;
  assign new_n21300_ = new_n15926_ & new_n21102_;
  assign new_n21301_ = new_n15926_ & new_n21104_;
  assign new_n21302_ = new_n15926_ & new_n21106_;
  assign new_n21303_ = ~new_n21301_ & ~new_n21302_;
  assign new_n21304_ = ~new_n21300_ & new_n21303_;
  assign new_n21305_ = new_n15926_ & new_n21112_;
  assign new_n21306_ = new_n15926_ & new_n21114_;
  assign new_n21307_ = new_n15926_ & new_n21116_;
  assign new_n21308_ = ~new_n21306_ & ~new_n21307_;
  assign new_n21309_ = ~new_n21305_ & new_n21308_;
  assign new_n21310_ = new_n21304_ & new_n21309_;
  assign new_n21311_ = new_n16045_ & new_n21015_;
  assign new_n21312_ = new_n16045_ & new_n21017_;
  assign new_n21313_ = new_n16045_ & new_n21019_;
  assign new_n21314_ = ~new_n21312_ & ~new_n21313_;
  assign new_n21315_ = ~new_n21311_ & new_n21314_;
  assign new_n21316_ = new_n16045_ & new_n21026_;
  assign new_n21317_ = new_n16045_ & new_n21029_;
  assign new_n21318_ = ~new_n21316_ & ~new_n21317_;
  assign new_n21319_ = new_n21315_ & new_n21318_;
  assign new_n21320_ = new_n21310_ & new_n21319_;
  assign new_n21321_ = new_n21299_ & new_n21320_;
  assign new_n21322_ = new_n16045_ & new_n21042_;
  assign new_n21323_ = new_n16045_ & new_n21024_;
  assign new_n21324_ = new_n16045_ & new_n21039_;
  assign new_n21325_ = ~new_n21323_ & ~new_n21324_;
  assign new_n21326_ = ~new_n21322_ & new_n21325_;
  assign new_n21327_ = new_n16045_ & new_n21053_;
  assign new_n21328_ = new_n16045_ & new_n21036_;
  assign new_n21329_ = new_n16045_ & new_n21050_;
  assign new_n21330_ = ~new_n21328_ & ~new_n21329_;
  assign new_n21331_ = ~new_n21327_ & new_n21330_;
  assign new_n21332_ = new_n21326_ & new_n21331_;
  assign new_n21333_ = new_n16045_ & new_n21062_;
  assign new_n21334_ = new_n16045_ & new_n21047_;
  assign new_n21335_ = new_n16045_ & new_n21060_;
  assign new_n21336_ = ~new_n21334_ & ~new_n21335_;
  assign new_n21337_ = ~new_n21333_ & new_n21336_;
  assign new_n21338_ = new_n16045_ & new_n21068_;
  assign new_n21339_ = new_n16045_ & new_n21058_;
  assign new_n21340_ = new_n16045_ & new_n21066_;
  assign new_n21341_ = ~new_n21339_ & ~new_n21340_;
  assign new_n21342_ = ~new_n21338_ & new_n21341_;
  assign new_n21343_ = new_n21337_ & new_n21342_;
  assign new_n21344_ = new_n21332_ & new_n21343_;
  assign new_n21345_ = new_n16045_ & new_n21077_;
  assign new_n21346_ = new_n16045_ & new_n21079_;
  assign new_n21347_ = new_n16045_ & new_n21081_;
  assign new_n21348_ = ~new_n21346_ & ~new_n21347_;
  assign new_n21349_ = ~new_n21345_ & new_n21348_;
  assign new_n21350_ = new_n16045_ & new_n21085_;
  assign new_n21351_ = new_n16045_ & new_n21087_;
  assign new_n21352_ = new_n16045_ & new_n21089_;
  assign new_n21353_ = ~new_n21351_ & ~new_n21352_;
  assign new_n21354_ = ~new_n21350_ & new_n21353_;
  assign new_n21355_ = new_n21349_ & new_n21354_;
  assign new_n21356_ = new_n16045_ & new_n21094_;
  assign new_n21357_ = new_n16045_ & new_n21096_;
  assign new_n21358_ = new_n16045_ & new_n21098_;
  assign new_n21359_ = ~new_n21357_ & ~new_n21358_;
  assign new_n21360_ = ~new_n21356_ & new_n21359_;
  assign new_n21361_ = new_n16045_ & new_n21104_;
  assign new_n21362_ = new_n16045_ & new_n21106_;
  assign new_n21363_ = ~new_n21361_ & ~new_n21362_;
  assign new_n21364_ = new_n21360_ & new_n21363_;
  assign new_n21365_ = new_n21355_ & new_n21364_;
  assign new_n21366_ = new_n21344_ & new_n21365_;
  assign new_n21367_ = new_n21321_ & new_n21366_;
  assign new_n21368_ = new_n16045_ & new_n21116_;
  assign new_n21369_ = new_n16045_ & new_n21102_;
  assign new_n21370_ = new_n16045_ & new_n21114_;
  assign new_n21371_ = ~new_n21369_ & ~new_n21370_;
  assign new_n21372_ = ~new_n21368_ & new_n21371_;
  assign new_n21373_ = new_n16094_ & new_n21019_;
  assign new_n21374_ = new_n16045_ & new_n21112_;
  assign new_n21375_ = new_n16094_ & new_n21017_;
  assign new_n21376_ = ~new_n21374_ & ~new_n21375_;
  assign new_n21377_ = ~new_n21373_ & new_n21376_;
  assign new_n21378_ = new_n21372_ & new_n21377_;
  assign new_n21379_ = new_n16094_ & new_n21029_;
  assign new_n21380_ = new_n16094_ & new_n21015_;
  assign new_n21381_ = new_n16094_ & new_n21026_;
  assign new_n21382_ = ~new_n21380_ & ~new_n21381_;
  assign new_n21383_ = ~new_n21379_ & new_n21382_;
  assign new_n21384_ = new_n16094_ & new_n21042_;
  assign new_n21385_ = new_n16094_ & new_n21024_;
  assign new_n21386_ = new_n16094_ & new_n21039_;
  assign new_n21387_ = ~new_n21385_ & ~new_n21386_;
  assign new_n21388_ = ~new_n21384_ & new_n21387_;
  assign new_n21389_ = new_n21383_ & new_n21388_;
  assign new_n21390_ = new_n21378_ & new_n21389_;
  assign new_n21391_ = new_n16094_ & new_n21053_;
  assign new_n21392_ = new_n16094_ & new_n21036_;
  assign new_n21393_ = new_n16094_ & new_n21050_;
  assign new_n21394_ = ~new_n21392_ & ~new_n21393_;
  assign new_n21395_ = ~new_n21391_ & new_n21394_;
  assign new_n21396_ = new_n16094_ & new_n21062_;
  assign new_n21397_ = new_n16094_ & new_n21047_;
  assign new_n21398_ = new_n16094_ & new_n21060_;
  assign new_n21399_ = ~new_n21397_ & ~new_n21398_;
  assign new_n21400_ = ~new_n21396_ & new_n21399_;
  assign new_n21401_ = new_n21395_ & new_n21400_;
  assign new_n21402_ = new_n16094_ & new_n21068_;
  assign new_n21403_ = new_n16094_ & new_n21058_;
  assign new_n21404_ = new_n16094_ & new_n21066_;
  assign new_n21405_ = ~new_n21403_ & ~new_n21404_;
  assign new_n21406_ = ~new_n21402_ & new_n21405_;
  assign new_n21407_ = new_n16094_ & new_n21079_;
  assign new_n21408_ = new_n16094_ & new_n21081_;
  assign new_n21409_ = ~new_n21407_ & ~new_n21408_;
  assign new_n21410_ = new_n21406_ & new_n21409_;
  assign new_n21411_ = new_n21401_ & new_n21410_;
  assign new_n21412_ = new_n21390_ & new_n21411_;
  assign new_n21413_ = new_n16094_ & new_n21089_;
  assign new_n21414_ = new_n16094_ & new_n21077_;
  assign new_n21415_ = new_n16094_ & new_n21087_;
  assign new_n21416_ = ~new_n21414_ & ~new_n21415_;
  assign new_n21417_ = ~new_n21413_ & new_n21416_;
  assign new_n21418_ = new_n16094_ & new_n21098_;
  assign new_n21419_ = new_n16094_ & new_n21085_;
  assign new_n21420_ = new_n16094_ & new_n21096_;
  assign new_n21421_ = ~new_n21419_ & ~new_n21420_;
  assign new_n21422_ = ~new_n21418_ & new_n21421_;
  assign new_n21423_ = new_n21417_ & new_n21422_;
  assign new_n21424_ = new_n16094_ & new_n21106_;
  assign new_n21425_ = new_n16094_ & new_n21094_;
  assign new_n21426_ = new_n16094_ & new_n21104_;
  assign new_n21427_ = ~new_n21425_ & ~new_n21426_;
  assign new_n21428_ = ~new_n21424_ & new_n21427_;
  assign new_n21429_ = new_n16094_ & new_n21116_;
  assign new_n21430_ = new_n16094_ & new_n21102_;
  assign new_n21431_ = new_n16094_ & new_n21114_;
  assign new_n21432_ = ~new_n21430_ & ~new_n21431_;
  assign new_n21433_ = ~new_n21429_ & new_n21432_;
  assign new_n21434_ = new_n21428_ & new_n21433_;
  assign new_n21435_ = new_n21423_ & new_n21434_;
  assign new_n21436_ = new_n16152_ & new_n21019_;
  assign new_n21437_ = new_n16094_ & new_n21112_;
  assign new_n21438_ = new_n16152_ & new_n21017_;
  assign new_n21439_ = ~new_n21437_ & ~new_n21438_;
  assign new_n21440_ = ~new_n21436_ & new_n21439_;
  assign new_n21441_ = new_n16152_ & new_n21029_;
  assign new_n21442_ = new_n16152_ & new_n21015_;
  assign new_n21443_ = new_n16152_ & new_n21026_;
  assign new_n21444_ = ~new_n21442_ & ~new_n21443_;
  assign new_n21445_ = ~new_n21441_ & new_n21444_;
  assign new_n21446_ = new_n21440_ & new_n21445_;
  assign new_n21447_ = new_n16152_ & new_n21042_;
  assign new_n21448_ = new_n16152_ & new_n21024_;
  assign new_n21449_ = new_n16152_ & new_n21039_;
  assign new_n21450_ = ~new_n21448_ & ~new_n21449_;
  assign new_n21451_ = ~new_n21447_ & new_n21450_;
  assign new_n21452_ = new_n16152_ & new_n21036_;
  assign new_n21453_ = new_n16152_ & new_n21050_;
  assign new_n21454_ = ~new_n21452_ & ~new_n21453_;
  assign new_n21455_ = new_n21451_ & new_n21454_;
  assign new_n21456_ = new_n21446_ & new_n21455_;
  assign new_n21457_ = new_n21435_ & new_n21456_;
  assign new_n21458_ = new_n21412_ & new_n21457_;
  assign new_n21459_ = new_n21367_ & new_n21458_;
  assign new_n21460_ = new_n21276_ & new_n21459_;
  assign new_n21461_ = new_n21076_ & new_n21460_;
  assign new_n21462_ = new_n16152_ & new_n21060_;
  assign new_n21463_ = new_n16152_ & new_n21053_;
  assign new_n21464_ = new_n16152_ & new_n21047_;
  assign new_n21465_ = ~new_n21463_ & ~new_n21464_;
  assign new_n21466_ = ~new_n21462_ & new_n21465_;
  assign new_n21467_ = new_n16152_ & new_n21066_;
  assign new_n21468_ = new_n16152_ & new_n21062_;
  assign new_n21469_ = new_n16152_ & new_n21058_;
  assign new_n21470_ = ~new_n21468_ & ~new_n21469_;
  assign new_n21471_ = ~new_n21467_ & new_n21470_;
  assign new_n21472_ = new_n21466_ & new_n21471_;
  assign new_n21473_ = new_n16152_ & new_n21081_;
  assign new_n21474_ = new_n16152_ & new_n21068_;
  assign new_n21475_ = new_n16152_ & new_n21079_;
  assign new_n21476_ = ~new_n21474_ & ~new_n21475_;
  assign new_n21477_ = ~new_n21473_ & new_n21476_;
  assign new_n21478_ = new_n16152_ & new_n21089_;
  assign new_n21479_ = new_n16152_ & new_n21077_;
  assign new_n21480_ = new_n16152_ & new_n21087_;
  assign new_n21481_ = ~new_n21479_ & ~new_n21480_;
  assign new_n21482_ = ~new_n21478_ & new_n21481_;
  assign new_n21483_ = new_n21477_ & new_n21482_;
  assign new_n21484_ = new_n21472_ & new_n21483_;
  assign new_n21485_ = new_n16152_ & new_n21098_;
  assign new_n21486_ = new_n16152_ & new_n21085_;
  assign new_n21487_ = new_n16152_ & new_n21096_;
  assign new_n21488_ = ~new_n21486_ & ~new_n21487_;
  assign new_n21489_ = ~new_n21485_ & new_n21488_;
  assign new_n21490_ = new_n16152_ & new_n21106_;
  assign new_n21491_ = new_n16152_ & new_n21094_;
  assign new_n21492_ = new_n16152_ & new_n21104_;
  assign new_n21493_ = ~new_n21491_ & ~new_n21492_;
  assign new_n21494_ = ~new_n21490_ & new_n21493_;
  assign new_n21495_ = new_n21489_ & new_n21494_;
  assign new_n21496_ = new_n16152_ & new_n21116_;
  assign new_n21497_ = new_n16152_ & new_n21102_;
  assign new_n21498_ = new_n16152_ & new_n21114_;
  assign new_n21499_ = ~new_n21497_ & ~new_n21498_;
  assign new_n21500_ = ~new_n21496_ & new_n21499_;
  assign new_n21501_ = new_n16201_ & new_n21019_;
  assign new_n21502_ = new_n16152_ & new_n21112_;
  assign new_n21503_ = new_n16201_ & new_n21017_;
  assign new_n21504_ = ~new_n21502_ & ~new_n21503_;
  assign new_n21505_ = ~new_n21501_ & new_n21504_;
  assign new_n21506_ = new_n21500_ & new_n21505_;
  assign new_n21507_ = new_n21495_ & new_n21506_;
  assign new_n21508_ = new_n21484_ & new_n21507_;
  assign new_n21509_ = new_n16201_ & new_n21029_;
  assign new_n21510_ = new_n16201_ & new_n21015_;
  assign new_n21511_ = new_n16201_ & new_n21026_;
  assign new_n21512_ = ~new_n21510_ & ~new_n21511_;
  assign new_n21513_ = ~new_n21509_ & new_n21512_;
  assign new_n21514_ = new_n16201_ & new_n21042_;
  assign new_n21515_ = new_n16201_ & new_n21024_;
  assign new_n21516_ = new_n16201_ & new_n21039_;
  assign new_n21517_ = ~new_n21515_ & ~new_n21516_;
  assign new_n21518_ = ~new_n21514_ & new_n21517_;
  assign new_n21519_ = new_n21513_ & new_n21518_;
  assign new_n21520_ = new_n16201_ & new_n21053_;
  assign new_n21521_ = new_n16201_ & new_n21036_;
  assign new_n21522_ = new_n16201_ & new_n21050_;
  assign new_n21523_ = ~new_n21521_ & ~new_n21522_;
  assign new_n21524_ = ~new_n21520_ & new_n21523_;
  assign new_n21525_ = new_n16201_ & new_n21062_;
  assign new_n21526_ = new_n16201_ & new_n21047_;
  assign new_n21527_ = new_n16201_ & new_n21060_;
  assign new_n21528_ = ~new_n21526_ & ~new_n21527_;
  assign new_n21529_ = ~new_n21525_ & new_n21528_;
  assign new_n21530_ = new_n21524_ & new_n21529_;
  assign new_n21531_ = new_n21519_ & new_n21530_;
  assign new_n21532_ = new_n16201_ & new_n21068_;
  assign new_n21533_ = new_n16201_ & new_n21058_;
  assign new_n21534_ = new_n16201_ & new_n21066_;
  assign new_n21535_ = ~new_n21533_ & ~new_n21534_;
  assign new_n21536_ = ~new_n21532_ & new_n21535_;
  assign new_n21537_ = new_n16201_ & new_n21077_;
  assign new_n21538_ = new_n16201_ & new_n21079_;
  assign new_n21539_ = new_n16201_ & new_n21081_;
  assign new_n21540_ = ~new_n21538_ & ~new_n21539_;
  assign new_n21541_ = ~new_n21537_ & new_n21540_;
  assign new_n21542_ = new_n21536_ & new_n21541_;
  assign new_n21543_ = new_n16201_ & new_n21085_;
  assign new_n21544_ = new_n16201_ & new_n21087_;
  assign new_n21545_ = new_n16201_ & new_n21089_;
  assign new_n21546_ = ~new_n21544_ & ~new_n21545_;
  assign new_n21547_ = ~new_n21543_ & new_n21546_;
  assign new_n21548_ = new_n16201_ & new_n21096_;
  assign new_n21549_ = new_n16201_ & new_n21098_;
  assign new_n21550_ = ~new_n21548_ & ~new_n21549_;
  assign new_n21551_ = new_n21547_ & new_n21550_;
  assign new_n21552_ = new_n21542_ & new_n21551_;
  assign new_n21553_ = new_n21531_ & new_n21552_;
  assign new_n21554_ = new_n21508_ & new_n21553_;
  assign new_n21555_ = new_n16201_ & new_n21106_;
  assign new_n21556_ = new_n16201_ & new_n21094_;
  assign new_n21557_ = new_n16201_ & new_n21104_;
  assign new_n21558_ = ~new_n21556_ & ~new_n21557_;
  assign new_n21559_ = ~new_n21555_ & new_n21558_;
  assign new_n21560_ = new_n16201_ & new_n21116_;
  assign new_n21561_ = new_n16201_ & new_n21102_;
  assign new_n21562_ = new_n16201_ & new_n21114_;
  assign new_n21563_ = ~new_n21561_ & ~new_n21562_;
  assign new_n21564_ = ~new_n21560_ & new_n21563_;
  assign new_n21565_ = new_n21559_ & new_n21564_;
  assign new_n21566_ = new_n16312_ & new_n21019_;
  assign new_n21567_ = new_n16201_ & new_n21112_;
  assign new_n21568_ = new_n16312_ & new_n21017_;
  assign new_n21569_ = ~new_n21567_ & ~new_n21568_;
  assign new_n21570_ = ~new_n21566_ & new_n21569_;
  assign new_n21571_ = new_n16312_ & new_n21029_;
  assign new_n21572_ = new_n16312_ & new_n21015_;
  assign new_n21573_ = new_n16312_ & new_n21026_;
  assign new_n21574_ = ~new_n21572_ & ~new_n21573_;
  assign new_n21575_ = ~new_n21571_ & new_n21574_;
  assign new_n21576_ = new_n21570_ & new_n21575_;
  assign new_n21577_ = new_n21565_ & new_n21576_;
  assign new_n21578_ = new_n16312_ & new_n21042_;
  assign new_n21579_ = new_n16312_ & new_n21024_;
  assign new_n21580_ = new_n16312_ & new_n21039_;
  assign new_n21581_ = ~new_n21579_ & ~new_n21580_;
  assign new_n21582_ = ~new_n21578_ & new_n21581_;
  assign new_n21583_ = new_n16312_ & new_n21053_;
  assign new_n21584_ = new_n16312_ & new_n21036_;
  assign new_n21585_ = new_n16312_ & new_n21050_;
  assign new_n21586_ = ~new_n21584_ & ~new_n21585_;
  assign new_n21587_ = ~new_n21583_ & new_n21586_;
  assign new_n21588_ = new_n21582_ & new_n21587_;
  assign new_n21589_ = new_n16312_ & new_n21062_;
  assign new_n21590_ = new_n16312_ & new_n21047_;
  assign new_n21591_ = new_n16312_ & new_n21060_;
  assign new_n21592_ = ~new_n21590_ & ~new_n21591_;
  assign new_n21593_ = ~new_n21589_ & new_n21592_;
  assign new_n21594_ = new_n16312_ & new_n21058_;
  assign new_n21595_ = new_n16312_ & new_n21066_;
  assign new_n21596_ = ~new_n21594_ & ~new_n21595_;
  assign new_n21597_ = new_n21593_ & new_n21596_;
  assign new_n21598_ = new_n21588_ & new_n21597_;
  assign new_n21599_ = new_n21577_ & new_n21598_;
  assign new_n21600_ = new_n16312_ & new_n21081_;
  assign new_n21601_ = new_n16312_ & new_n21068_;
  assign new_n21602_ = new_n16312_ & new_n21079_;
  assign new_n21603_ = ~new_n21601_ & ~new_n21602_;
  assign new_n21604_ = ~new_n21600_ & new_n21603_;
  assign new_n21605_ = new_n16312_ & new_n21089_;
  assign new_n21606_ = new_n16312_ & new_n21077_;
  assign new_n21607_ = new_n16312_ & new_n21087_;
  assign new_n21608_ = ~new_n21606_ & ~new_n21607_;
  assign new_n21609_ = ~new_n21605_ & new_n21608_;
  assign new_n21610_ = new_n21604_ & new_n21609_;
  assign new_n21611_ = new_n16312_ & new_n21098_;
  assign new_n21612_ = new_n16312_ & new_n21085_;
  assign new_n21613_ = new_n16312_ & new_n21096_;
  assign new_n21614_ = ~new_n21612_ & ~new_n21613_;
  assign new_n21615_ = ~new_n21611_ & new_n21614_;
  assign new_n21616_ = new_n16312_ & new_n21106_;
  assign new_n21617_ = new_n16312_ & new_n21094_;
  assign new_n21618_ = new_n16312_ & new_n21104_;
  assign new_n21619_ = ~new_n21617_ & ~new_n21618_;
  assign new_n21620_ = ~new_n21616_ & new_n21619_;
  assign new_n21621_ = new_n21615_ & new_n21620_;
  assign new_n21622_ = new_n21610_ & new_n21621_;
  assign new_n21623_ = new_n16312_ & new_n21116_;
  assign new_n21624_ = new_n16312_ & new_n21102_;
  assign new_n21625_ = new_n16312_ & new_n21114_;
  assign new_n21626_ = ~new_n21624_ & ~new_n21625_;
  assign new_n21627_ = ~new_n21623_ & new_n21626_;
  assign new_n21628_ = new_n16361_ & new_n21019_;
  assign new_n21629_ = new_n16312_ & new_n21112_;
  assign new_n21630_ = new_n16361_ & new_n21017_;
  assign new_n21631_ = ~new_n21629_ & ~new_n21630_;
  assign new_n21632_ = ~new_n21628_ & new_n21631_;
  assign new_n21633_ = new_n21627_ & new_n21632_;
  assign new_n21634_ = new_n16361_ & new_n21029_;
  assign new_n21635_ = new_n16361_ & new_n21015_;
  assign new_n21636_ = new_n16361_ & new_n21026_;
  assign new_n21637_ = ~new_n21635_ & ~new_n21636_;
  assign new_n21638_ = ~new_n21634_ & new_n21637_;
  assign new_n21639_ = new_n16361_ & new_n21024_;
  assign new_n21640_ = new_n16361_ & new_n21039_;
  assign new_n21641_ = ~new_n21639_ & ~new_n21640_;
  assign new_n21642_ = new_n21638_ & new_n21641_;
  assign new_n21643_ = new_n21633_ & new_n21642_;
  assign new_n21644_ = new_n21622_ & new_n21643_;
  assign new_n21645_ = new_n21599_ & new_n21644_;
  assign new_n21646_ = new_n21554_ & new_n21645_;
  assign new_n21647_ = new_n16361_ & new_n21050_;
  assign new_n21648_ = new_n16361_ & new_n21042_;
  assign new_n21649_ = new_n16361_ & new_n21036_;
  assign new_n21650_ = ~new_n21648_ & ~new_n21649_;
  assign new_n21651_ = ~new_n21647_ & new_n21650_;
  assign new_n21652_ = new_n16361_ & new_n21060_;
  assign new_n21653_ = new_n16361_ & new_n21053_;
  assign new_n21654_ = new_n16361_ & new_n21047_;
  assign new_n21655_ = ~new_n21653_ & ~new_n21654_;
  assign new_n21656_ = ~new_n21652_ & new_n21655_;
  assign new_n21657_ = new_n21651_ & new_n21656_;
  assign new_n21658_ = new_n16361_ & new_n21066_;
  assign new_n21659_ = new_n16361_ & new_n21062_;
  assign new_n21660_ = new_n16361_ & new_n21058_;
  assign new_n21661_ = ~new_n21659_ & ~new_n21660_;
  assign new_n21662_ = ~new_n21658_ & new_n21661_;
  assign new_n21663_ = new_n16361_ & new_n21081_;
  assign new_n21664_ = new_n16361_ & new_n21068_;
  assign new_n21665_ = new_n16361_ & new_n21079_;
  assign new_n21666_ = ~new_n21664_ & ~new_n21665_;
  assign new_n21667_ = ~new_n21663_ & new_n21666_;
  assign new_n21668_ = new_n21662_ & new_n21667_;
  assign new_n21669_ = new_n21657_ & new_n21668_;
  assign new_n21670_ = new_n16361_ & new_n21089_;
  assign new_n21671_ = new_n16361_ & new_n21077_;
  assign new_n21672_ = new_n16361_ & new_n21087_;
  assign new_n21673_ = ~new_n21671_ & ~new_n21672_;
  assign new_n21674_ = ~new_n21670_ & new_n21673_;
  assign new_n21675_ = new_n16361_ & new_n21098_;
  assign new_n21676_ = new_n16361_ & new_n21085_;
  assign new_n21677_ = new_n16361_ & new_n21096_;
  assign new_n21678_ = ~new_n21676_ & ~new_n21677_;
  assign new_n21679_ = ~new_n21675_ & new_n21678_;
  assign new_n21680_ = new_n21674_ & new_n21679_;
  assign new_n21681_ = new_n16361_ & new_n21106_;
  assign new_n21682_ = new_n16361_ & new_n21094_;
  assign new_n21683_ = new_n16361_ & new_n21104_;
  assign new_n21684_ = ~new_n21682_ & ~new_n21683_;
  assign new_n21685_ = ~new_n21681_ & new_n21684_;
  assign new_n21686_ = new_n16361_ & new_n21102_;
  assign new_n21687_ = new_n16361_ & new_n21114_;
  assign new_n21688_ = ~new_n21686_ & ~new_n21687_;
  assign new_n21689_ = new_n21685_ & new_n21688_;
  assign new_n21690_ = new_n21680_ & new_n21689_;
  assign new_n21691_ = new_n21669_ & new_n21690_;
  assign new_n21692_ = new_n16415_ & new_n21017_;
  assign new_n21693_ = new_n16361_ & new_n21116_;
  assign new_n21694_ = new_n16361_ & new_n21112_;
  assign new_n21695_ = ~new_n21693_ & ~new_n21694_;
  assign new_n21696_ = ~new_n21692_ & new_n21695_;
  assign new_n21697_ = new_n16415_ & new_n21026_;
  assign new_n21698_ = new_n16415_ & new_n21019_;
  assign new_n21699_ = new_n16415_ & new_n21015_;
  assign new_n21700_ = ~new_n21698_ & ~new_n21699_;
  assign new_n21701_ = ~new_n21697_ & new_n21700_;
  assign new_n21702_ = new_n21696_ & new_n21701_;
  assign new_n21703_ = new_n16415_ & new_n21039_;
  assign new_n21704_ = new_n16415_ & new_n21029_;
  assign new_n21705_ = new_n16415_ & new_n21024_;
  assign new_n21706_ = ~new_n21704_ & ~new_n21705_;
  assign new_n21707_ = ~new_n21703_ & new_n21706_;
  assign new_n21708_ = new_n16415_ & new_n21050_;
  assign new_n21709_ = new_n16415_ & new_n21042_;
  assign new_n21710_ = new_n16415_ & new_n21036_;
  assign new_n21711_ = ~new_n21709_ & ~new_n21710_;
  assign new_n21712_ = ~new_n21708_ & new_n21711_;
  assign new_n21713_ = new_n21707_ & new_n21712_;
  assign new_n21714_ = new_n21702_ & new_n21713_;
  assign new_n21715_ = new_n16415_ & new_n21060_;
  assign new_n21716_ = new_n16415_ & new_n21053_;
  assign new_n21717_ = new_n16415_ & new_n21047_;
  assign new_n21718_ = ~new_n21716_ & ~new_n21717_;
  assign new_n21719_ = ~new_n21715_ & new_n21718_;
  assign new_n21720_ = new_n16415_ & new_n21066_;
  assign new_n21721_ = new_n16415_ & new_n21062_;
  assign new_n21722_ = new_n16415_ & new_n21058_;
  assign new_n21723_ = ~new_n21721_ & ~new_n21722_;
  assign new_n21724_ = ~new_n21720_ & new_n21723_;
  assign new_n21725_ = new_n21719_ & new_n21724_;
  assign new_n21726_ = new_n16415_ & new_n21081_;
  assign new_n21727_ = new_n16415_ & new_n21068_;
  assign new_n21728_ = new_n16415_ & new_n21079_;
  assign new_n21729_ = ~new_n21727_ & ~new_n21728_;
  assign new_n21730_ = ~new_n21726_ & new_n21729_;
  assign new_n21731_ = new_n16415_ & new_n21077_;
  assign new_n21732_ = new_n16415_ & new_n21087_;
  assign new_n21733_ = ~new_n21731_ & ~new_n21732_;
  assign new_n21734_ = new_n21730_ & new_n21733_;
  assign new_n21735_ = new_n21725_ & new_n21734_;
  assign new_n21736_ = new_n21714_ & new_n21735_;
  assign new_n21737_ = new_n21691_ & new_n21736_;
  assign new_n21738_ = new_n16415_ & new_n21096_;
  assign new_n21739_ = new_n16415_ & new_n21089_;
  assign new_n21740_ = new_n16415_ & new_n21085_;
  assign new_n21741_ = ~new_n21739_ & ~new_n21740_;
  assign new_n21742_ = ~new_n21738_ & new_n21741_;
  assign new_n21743_ = new_n16415_ & new_n21104_;
  assign new_n21744_ = new_n16415_ & new_n21098_;
  assign new_n21745_ = new_n16415_ & new_n21094_;
  assign new_n21746_ = ~new_n21744_ & ~new_n21745_;
  assign new_n21747_ = ~new_n21743_ & new_n21746_;
  assign new_n21748_ = new_n21742_ & new_n21747_;
  assign new_n21749_ = new_n16415_ & new_n21114_;
  assign new_n21750_ = new_n16415_ & new_n21106_;
  assign new_n21751_ = new_n16415_ & new_n21102_;
  assign new_n21752_ = ~new_n21750_ & ~new_n21751_;
  assign new_n21753_ = ~new_n21749_ & new_n21752_;
  assign new_n21754_ = new_n16463_ & new_n21017_;
  assign new_n21755_ = new_n16415_ & new_n21116_;
  assign new_n21756_ = new_n16415_ & new_n21112_;
  assign new_n21757_ = ~new_n21755_ & ~new_n21756_;
  assign new_n21758_ = ~new_n21754_ & new_n21757_;
  assign new_n21759_ = new_n21753_ & new_n21758_;
  assign new_n21760_ = new_n21748_ & new_n21759_;
  assign new_n21761_ = new_n16463_ & new_n21026_;
  assign new_n21762_ = new_n16463_ & new_n21019_;
  assign new_n21763_ = new_n16463_ & new_n21015_;
  assign new_n21764_ = ~new_n21762_ & ~new_n21763_;
  assign new_n21765_ = ~new_n21761_ & new_n21764_;
  assign new_n21766_ = new_n16463_ & new_n21039_;
  assign new_n21767_ = new_n16463_ & new_n21029_;
  assign new_n21768_ = new_n16463_ & new_n21024_;
  assign new_n21769_ = ~new_n21767_ & ~new_n21768_;
  assign new_n21770_ = ~new_n21766_ & new_n21769_;
  assign new_n21771_ = new_n21765_ & new_n21770_;
  assign new_n21772_ = new_n16463_ & new_n21050_;
  assign new_n21773_ = new_n16463_ & new_n21042_;
  assign new_n21774_ = new_n16463_ & new_n21036_;
  assign new_n21775_ = ~new_n21773_ & ~new_n21774_;
  assign new_n21776_ = ~new_n21772_ & new_n21775_;
  assign new_n21777_ = new_n16463_ & new_n21053_;
  assign new_n21778_ = new_n16463_ & new_n21047_;
  assign new_n21779_ = ~new_n21777_ & ~new_n21778_;
  assign new_n21780_ = new_n21776_ & new_n21779_;
  assign new_n21781_ = new_n21771_ & new_n21780_;
  assign new_n21782_ = new_n21760_ & new_n21781_;
  assign new_n21783_ = new_n16463_ & new_n21058_;
  assign new_n21784_ = new_n16463_ & new_n21060_;
  assign new_n21785_ = new_n16463_ & new_n21062_;
  assign new_n21786_ = ~new_n21784_ & ~new_n21785_;
  assign new_n21787_ = ~new_n21783_ & new_n21786_;
  assign new_n21788_ = new_n16463_ & new_n21079_;
  assign new_n21789_ = new_n16463_ & new_n21066_;
  assign new_n21790_ = new_n16463_ & new_n21068_;
  assign new_n21791_ = ~new_n21789_ & ~new_n21790_;
  assign new_n21792_ = ~new_n21788_ & new_n21791_;
  assign new_n21793_ = new_n21787_ & new_n21792_;
  assign new_n21794_ = new_n16463_ & new_n21087_;
  assign new_n21795_ = new_n16463_ & new_n21081_;
  assign new_n21796_ = new_n16463_ & new_n21077_;
  assign new_n21797_ = ~new_n21795_ & ~new_n21796_;
  assign new_n21798_ = ~new_n21794_ & new_n21797_;
  assign new_n21799_ = new_n16463_ & new_n21096_;
  assign new_n21800_ = new_n16463_ & new_n21089_;
  assign new_n21801_ = new_n16463_ & new_n21085_;
  assign new_n21802_ = ~new_n21800_ & ~new_n21801_;
  assign new_n21803_ = ~new_n21799_ & new_n21802_;
  assign new_n21804_ = new_n21798_ & new_n21803_;
  assign new_n21805_ = new_n21793_ & new_n21804_;
  assign new_n21806_ = new_n16463_ & new_n21104_;
  assign new_n21807_ = new_n16463_ & new_n21098_;
  assign new_n21808_ = new_n16463_ & new_n21094_;
  assign new_n21809_ = ~new_n21807_ & ~new_n21808_;
  assign new_n21810_ = ~new_n21806_ & new_n21809_;
  assign new_n21811_ = new_n16463_ & new_n21114_;
  assign new_n21812_ = new_n16463_ & new_n21106_;
  assign new_n21813_ = new_n16463_ & new_n21102_;
  assign new_n21814_ = ~new_n21812_ & ~new_n21813_;
  assign new_n21815_ = ~new_n21811_ & new_n21814_;
  assign new_n21816_ = new_n21810_ & new_n21815_;
  assign new_n21817_ = new_n16576_ & new_n21017_;
  assign new_n21818_ = new_n16463_ & new_n21116_;
  assign new_n21819_ = new_n16463_ & new_n21112_;
  assign new_n21820_ = ~new_n21818_ & ~new_n21819_;
  assign new_n21821_ = ~new_n21817_ & new_n21820_;
  assign new_n21822_ = new_n16576_ & new_n21019_;
  assign new_n21823_ = new_n16576_ & new_n21015_;
  assign new_n21824_ = ~new_n21822_ & ~new_n21823_;
  assign new_n21825_ = new_n21821_ & new_n21824_;
  assign new_n21826_ = new_n21816_ & new_n21825_;
  assign new_n21827_ = new_n21805_ & new_n21826_;
  assign new_n21828_ = new_n21782_ & new_n21827_;
  assign new_n21829_ = new_n21737_ & new_n21828_;
  assign new_n21830_ = new_n21646_ & new_n21829_;
  assign new_n21831_ = new_n16576_ & new_n21024_;
  assign new_n21832_ = new_n16576_ & new_n21026_;
  assign new_n21833_ = new_n16576_ & new_n21029_;
  assign new_n21834_ = ~new_n21832_ & ~new_n21833_;
  assign new_n21835_ = ~new_n21831_ & new_n21834_;
  assign new_n21836_ = new_n16576_ & new_n21036_;
  assign new_n21837_ = new_n16576_ & new_n21039_;
  assign new_n21838_ = new_n16576_ & new_n21042_;
  assign new_n21839_ = ~new_n21837_ & ~new_n21838_;
  assign new_n21840_ = ~new_n21836_ & new_n21839_;
  assign new_n21841_ = new_n21835_ & new_n21840_;
  assign new_n21842_ = new_n16576_ & new_n21047_;
  assign new_n21843_ = new_n16576_ & new_n21050_;
  assign new_n21844_ = new_n16576_ & new_n21053_;
  assign new_n21845_ = ~new_n21843_ & ~new_n21844_;
  assign new_n21846_ = ~new_n21842_ & new_n21845_;
  assign new_n21847_ = new_n16576_ & new_n21058_;
  assign new_n21848_ = new_n16576_ & new_n21060_;
  assign new_n21849_ = new_n16576_ & new_n21062_;
  assign new_n21850_ = ~new_n21848_ & ~new_n21849_;
  assign new_n21851_ = ~new_n21847_ & new_n21850_;
  assign new_n21852_ = new_n21846_ & new_n21851_;
  assign new_n21853_ = new_n21841_ & new_n21852_;
  assign new_n21854_ = new_n16576_ & new_n21079_;
  assign new_n21855_ = new_n16576_ & new_n21066_;
  assign new_n21856_ = new_n16576_ & new_n21068_;
  assign new_n21857_ = ~new_n21855_ & ~new_n21856_;
  assign new_n21858_ = ~new_n21854_ & new_n21857_;
  assign new_n21859_ = new_n16576_ & new_n21087_;
  assign new_n21860_ = new_n16576_ & new_n21081_;
  assign new_n21861_ = new_n16576_ & new_n21077_;
  assign new_n21862_ = ~new_n21860_ & ~new_n21861_;
  assign new_n21863_ = ~new_n21859_ & new_n21862_;
  assign new_n21864_ = new_n21858_ & new_n21863_;
  assign new_n21865_ = new_n16576_ & new_n21096_;
  assign new_n21866_ = new_n16576_ & new_n21089_;
  assign new_n21867_ = new_n16576_ & new_n21085_;
  assign new_n21868_ = ~new_n21866_ & ~new_n21867_;
  assign new_n21869_ = ~new_n21865_ & new_n21868_;
  assign new_n21870_ = new_n16576_ & new_n21098_;
  assign new_n21871_ = new_n16576_ & new_n21094_;
  assign new_n21872_ = ~new_n21870_ & ~new_n21871_;
  assign new_n21873_ = new_n21869_ & new_n21872_;
  assign new_n21874_ = new_n21864_ & new_n21873_;
  assign new_n21875_ = new_n21853_ & new_n21874_;
  assign new_n21876_ = new_n16576_ & new_n21102_;
  assign new_n21877_ = new_n16576_ & new_n21104_;
  assign new_n21878_ = new_n16576_ & new_n21106_;
  assign new_n21879_ = ~new_n21877_ & ~new_n21878_;
  assign new_n21880_ = ~new_n21876_ & new_n21879_;
  assign new_n21881_ = new_n16576_ & new_n21112_;
  assign new_n21882_ = new_n16576_ & new_n21114_;
  assign new_n21883_ = new_n16576_ & new_n21116_;
  assign new_n21884_ = ~new_n21882_ & ~new_n21883_;
  assign new_n21885_ = ~new_n21881_ & new_n21884_;
  assign new_n21886_ = new_n21880_ & new_n21885_;
  assign new_n21887_ = new_n16632_ & new_n21015_;
  assign new_n21888_ = new_n16632_ & new_n21017_;
  assign new_n21889_ = new_n16632_ & new_n21019_;
  assign new_n21890_ = ~new_n21888_ & ~new_n21889_;
  assign new_n21891_ = ~new_n21887_ & new_n21890_;
  assign new_n21892_ = new_n16632_ & new_n21024_;
  assign new_n21893_ = new_n16632_ & new_n21026_;
  assign new_n21894_ = new_n16632_ & new_n21029_;
  assign new_n21895_ = ~new_n21893_ & ~new_n21894_;
  assign new_n21896_ = ~new_n21892_ & new_n21895_;
  assign new_n21897_ = new_n21891_ & new_n21896_;
  assign new_n21898_ = new_n21886_ & new_n21897_;
  assign new_n21899_ = new_n16632_ & new_n21036_;
  assign new_n21900_ = new_n16632_ & new_n21039_;
  assign new_n21901_ = new_n16632_ & new_n21042_;
  assign new_n21902_ = ~new_n21900_ & ~new_n21901_;
  assign new_n21903_ = ~new_n21899_ & new_n21902_;
  assign new_n21904_ = new_n16632_ & new_n21047_;
  assign new_n21905_ = new_n16632_ & new_n21050_;
  assign new_n21906_ = new_n16632_ & new_n21053_;
  assign new_n21907_ = ~new_n21905_ & ~new_n21906_;
  assign new_n21908_ = ~new_n21904_ & new_n21907_;
  assign new_n21909_ = new_n21903_ & new_n21908_;
  assign new_n21910_ = new_n16632_ & new_n21058_;
  assign new_n21911_ = new_n16632_ & new_n21060_;
  assign new_n21912_ = new_n16632_ & new_n21062_;
  assign new_n21913_ = ~new_n21911_ & ~new_n21912_;
  assign new_n21914_ = ~new_n21910_ & new_n21913_;
  assign new_n21915_ = new_n16632_ & new_n21066_;
  assign new_n21916_ = new_n16632_ & new_n21068_;
  assign new_n21917_ = ~new_n21915_ & ~new_n21916_;
  assign new_n21918_ = new_n21914_ & new_n21917_;
  assign new_n21919_ = new_n21909_ & new_n21918_;
  assign new_n21920_ = new_n21898_ & new_n21919_;
  assign new_n21921_ = new_n21875_ & new_n21920_;
  assign new_n21922_ = new_n16632_ & new_n21077_;
  assign new_n21923_ = new_n16632_ & new_n21079_;
  assign new_n21924_ = new_n16632_ & new_n21081_;
  assign new_n21925_ = ~new_n21923_ & ~new_n21924_;
  assign new_n21926_ = ~new_n21922_ & new_n21925_;
  assign new_n21927_ = new_n16632_ & new_n21085_;
  assign new_n21928_ = new_n16632_ & new_n21087_;
  assign new_n21929_ = new_n16632_ & new_n21089_;
  assign new_n21930_ = ~new_n21928_ & ~new_n21929_;
  assign new_n21931_ = ~new_n21927_ & new_n21930_;
  assign new_n21932_ = new_n21926_ & new_n21931_;
  assign new_n21933_ = new_n16632_ & new_n21094_;
  assign new_n21934_ = new_n16632_ & new_n21096_;
  assign new_n21935_ = new_n16632_ & new_n21098_;
  assign new_n21936_ = ~new_n21934_ & ~new_n21935_;
  assign new_n21937_ = ~new_n21933_ & new_n21936_;
  assign new_n21938_ = new_n16632_ & new_n21102_;
  assign new_n21939_ = new_n16632_ & new_n21104_;
  assign new_n21940_ = new_n16632_ & new_n21106_;
  assign new_n21941_ = ~new_n21939_ & ~new_n21940_;
  assign new_n21942_ = ~new_n21938_ & new_n21941_;
  assign new_n21943_ = new_n21937_ & new_n21942_;
  assign new_n21944_ = new_n21932_ & new_n21943_;
  assign new_n21945_ = new_n16632_ & new_n21112_;
  assign new_n21946_ = new_n16632_ & new_n21114_;
  assign new_n21947_ = new_n16632_ & new_n21116_;
  assign new_n21948_ = ~new_n21946_ & ~new_n21947_;
  assign new_n21949_ = ~new_n21945_ & new_n21948_;
  assign new_n21950_ = new_n16679_ & new_n21015_;
  assign new_n21951_ = new_n16679_ & new_n21017_;
  assign new_n21952_ = new_n16679_ & new_n21019_;
  assign new_n21953_ = ~new_n21951_ & ~new_n21952_;
  assign new_n21954_ = ~new_n21950_ & new_n21953_;
  assign new_n21955_ = new_n21949_ & new_n21954_;
  assign new_n21956_ = new_n16679_ & new_n21024_;
  assign new_n21957_ = new_n16679_ & new_n21026_;
  assign new_n21958_ = new_n16679_ & new_n21029_;
  assign new_n21959_ = ~new_n21957_ & ~new_n21958_;
  assign new_n21960_ = ~new_n21956_ & new_n21959_;
  assign new_n21961_ = new_n16679_ & new_n21039_;
  assign new_n21962_ = new_n16679_ & new_n21042_;
  assign new_n21963_ = ~new_n21961_ & ~new_n21962_;
  assign new_n21964_ = new_n21960_ & new_n21963_;
  assign new_n21965_ = new_n21955_ & new_n21964_;
  assign new_n21966_ = new_n21944_ & new_n21965_;
  assign new_n21967_ = new_n16679_ & new_n21053_;
  assign new_n21968_ = new_n16679_ & new_n21036_;
  assign new_n21969_ = new_n16679_ & new_n21050_;
  assign new_n21970_ = ~new_n21968_ & ~new_n21969_;
  assign new_n21971_ = ~new_n21967_ & new_n21970_;
  assign new_n21972_ = new_n16679_ & new_n21062_;
  assign new_n21973_ = new_n16679_ & new_n21047_;
  assign new_n21974_ = new_n16679_ & new_n21060_;
  assign new_n21975_ = ~new_n21973_ & ~new_n21974_;
  assign new_n21976_ = ~new_n21972_ & new_n21975_;
  assign new_n21977_ = new_n21971_ & new_n21976_;
  assign new_n21978_ = new_n16679_ & new_n21068_;
  assign new_n21979_ = new_n16679_ & new_n21058_;
  assign new_n21980_ = new_n16679_ & new_n21066_;
  assign new_n21981_ = ~new_n21979_ & ~new_n21980_;
  assign new_n21982_ = ~new_n21978_ & new_n21981_;
  assign new_n21983_ = new_n16679_ & new_n21077_;
  assign new_n21984_ = new_n16679_ & new_n21079_;
  assign new_n21985_ = new_n16679_ & new_n21081_;
  assign new_n21986_ = ~new_n21984_ & ~new_n21985_;
  assign new_n21987_ = ~new_n21983_ & new_n21986_;
  assign new_n21988_ = new_n21982_ & new_n21987_;
  assign new_n21989_ = new_n21977_ & new_n21988_;
  assign new_n21990_ = new_n16679_ & new_n21085_;
  assign new_n21991_ = new_n16679_ & new_n21087_;
  assign new_n21992_ = new_n16679_ & new_n21089_;
  assign new_n21993_ = ~new_n21991_ & ~new_n21992_;
  assign new_n21994_ = ~new_n21990_ & new_n21993_;
  assign new_n21995_ = new_n16679_ & new_n21094_;
  assign new_n21996_ = new_n16679_ & new_n21096_;
  assign new_n21997_ = new_n16679_ & new_n21098_;
  assign new_n21998_ = ~new_n21996_ & ~new_n21997_;
  assign new_n21999_ = ~new_n21995_ & new_n21998_;
  assign new_n22000_ = new_n21994_ & new_n21999_;
  assign new_n22001_ = new_n16679_ & new_n21102_;
  assign new_n22002_ = new_n16679_ & new_n21104_;
  assign new_n22003_ = new_n16679_ & new_n21106_;
  assign new_n22004_ = ~new_n22002_ & ~new_n22003_;
  assign new_n22005_ = ~new_n22001_ & new_n22004_;
  assign new_n22006_ = new_n16679_ & new_n21114_;
  assign new_n22007_ = new_n16679_ & new_n21116_;
  assign new_n22008_ = ~new_n22006_ & ~new_n22007_;
  assign new_n22009_ = new_n22005_ & new_n22008_;
  assign new_n22010_ = new_n22000_ & new_n22009_;
  assign new_n22011_ = new_n21989_ & new_n22010_;
  assign new_n22012_ = new_n21966_ & new_n22011_;
  assign new_n22013_ = new_n21921_ & new_n22012_;
  assign new_n22014_ = new_n16728_ & new_n21019_;
  assign new_n22015_ = new_n16679_ & new_n21112_;
  assign new_n22016_ = new_n16728_ & new_n21017_;
  assign new_n22017_ = ~new_n22015_ & ~new_n22016_;
  assign new_n22018_ = ~new_n22014_ & new_n22017_;
  assign new_n22019_ = new_n16728_ & new_n21029_;
  assign new_n22020_ = new_n16728_ & new_n21015_;
  assign new_n22021_ = new_n16728_ & new_n21026_;
  assign new_n22022_ = ~new_n22020_ & ~new_n22021_;
  assign new_n22023_ = ~new_n22019_ & new_n22022_;
  assign new_n22024_ = new_n22018_ & new_n22023_;
  assign new_n22025_ = new_n16728_ & new_n21042_;
  assign new_n22026_ = new_n16728_ & new_n21024_;
  assign new_n22027_ = new_n16728_ & new_n21039_;
  assign new_n22028_ = ~new_n22026_ & ~new_n22027_;
  assign new_n22029_ = ~new_n22025_ & new_n22028_;
  assign new_n22030_ = new_n16728_ & new_n21053_;
  assign new_n22031_ = new_n16728_ & new_n21036_;
  assign new_n22032_ = new_n16728_ & new_n21050_;
  assign new_n22033_ = ~new_n22031_ & ~new_n22032_;
  assign new_n22034_ = ~new_n22030_ & new_n22033_;
  assign new_n22035_ = new_n22029_ & new_n22034_;
  assign new_n22036_ = new_n22024_ & new_n22035_;
  assign new_n22037_ = new_n16728_ & new_n21062_;
  assign new_n22038_ = new_n16728_ & new_n21047_;
  assign new_n22039_ = new_n16728_ & new_n21060_;
  assign new_n22040_ = ~new_n22038_ & ~new_n22039_;
  assign new_n22041_ = ~new_n22037_ & new_n22040_;
  assign new_n22042_ = new_n16728_ & new_n21068_;
  assign new_n22043_ = new_n16728_ & new_n21058_;
  assign new_n22044_ = new_n16728_ & new_n21066_;
  assign new_n22045_ = ~new_n22043_ & ~new_n22044_;
  assign new_n22046_ = ~new_n22042_ & new_n22045_;
  assign new_n22047_ = new_n22041_ & new_n22046_;
  assign new_n22048_ = new_n16728_ & new_n21077_;
  assign new_n22049_ = new_n16728_ & new_n21079_;
  assign new_n22050_ = new_n16728_ & new_n21081_;
  assign new_n22051_ = ~new_n22049_ & ~new_n22050_;
  assign new_n22052_ = ~new_n22048_ & new_n22051_;
  assign new_n22053_ = new_n16728_ & new_n21087_;
  assign new_n22054_ = new_n16728_ & new_n21089_;
  assign new_n22055_ = ~new_n22053_ & ~new_n22054_;
  assign new_n22056_ = new_n22052_ & new_n22055_;
  assign new_n22057_ = new_n22047_ & new_n22056_;
  assign new_n22058_ = new_n22036_ & new_n22057_;
  assign new_n22059_ = new_n16728_ & new_n21098_;
  assign new_n22060_ = new_n16728_ & new_n21085_;
  assign new_n22061_ = new_n16728_ & new_n21096_;
  assign new_n22062_ = ~new_n22060_ & ~new_n22061_;
  assign new_n22063_ = ~new_n22059_ & new_n22062_;
  assign new_n22064_ = new_n16728_ & new_n21106_;
  assign new_n22065_ = new_n16728_ & new_n21094_;
  assign new_n22066_ = new_n16728_ & new_n21104_;
  assign new_n22067_ = ~new_n22065_ & ~new_n22066_;
  assign new_n22068_ = ~new_n22064_ & new_n22067_;
  assign new_n22069_ = new_n22063_ & new_n22068_;
  assign new_n22070_ = new_n16728_ & new_n21116_;
  assign new_n22071_ = new_n16728_ & new_n21102_;
  assign new_n22072_ = new_n16728_ & new_n21114_;
  assign new_n22073_ = ~new_n22071_ & ~new_n22072_;
  assign new_n22074_ = ~new_n22070_ & new_n22073_;
  assign new_n22075_ = new_n17107_ & new_n21019_;
  assign new_n22076_ = new_n16728_ & new_n21112_;
  assign new_n22077_ = new_n17107_ & new_n21017_;
  assign new_n22078_ = ~new_n22076_ & ~new_n22077_;
  assign new_n22079_ = ~new_n22075_ & new_n22078_;
  assign new_n22080_ = new_n22074_ & new_n22079_;
  assign new_n22081_ = new_n22069_ & new_n22080_;
  assign new_n22082_ = new_n17107_ & new_n21029_;
  assign new_n22083_ = new_n17107_ & new_n21015_;
  assign new_n22084_ = new_n17107_ & new_n21026_;
  assign new_n22085_ = ~new_n22083_ & ~new_n22084_;
  assign new_n22086_ = ~new_n22082_ & new_n22085_;
  assign new_n22087_ = new_n17107_ & new_n21042_;
  assign new_n22088_ = new_n17107_ & new_n21024_;
  assign new_n22089_ = new_n17107_ & new_n21039_;
  assign new_n22090_ = ~new_n22088_ & ~new_n22089_;
  assign new_n22091_ = ~new_n22087_ & new_n22090_;
  assign new_n22092_ = new_n22086_ & new_n22091_;
  assign new_n22093_ = new_n17107_ & new_n21053_;
  assign new_n22094_ = new_n17107_ & new_n21036_;
  assign new_n22095_ = new_n17107_ & new_n21050_;
  assign new_n22096_ = ~new_n22094_ & ~new_n22095_;
  assign new_n22097_ = ~new_n22093_ & new_n22096_;
  assign new_n22098_ = new_n17107_ & new_n21047_;
  assign new_n22099_ = new_n17107_ & new_n21060_;
  assign new_n22100_ = ~new_n22098_ & ~new_n22099_;
  assign new_n22101_ = new_n22097_ & new_n22100_;
  assign new_n22102_ = new_n22092_ & new_n22101_;
  assign new_n22103_ = new_n22081_ & new_n22102_;
  assign new_n22104_ = new_n22058_ & new_n22103_;
  assign new_n22105_ = new_n17107_ & new_n21066_;
  assign new_n22106_ = new_n17107_ & new_n21062_;
  assign new_n22107_ = new_n17107_ & new_n21058_;
  assign new_n22108_ = ~new_n22106_ & ~new_n22107_;
  assign new_n22109_ = ~new_n22105_ & new_n22108_;
  assign new_n22110_ = new_n17107_ & new_n21081_;
  assign new_n22111_ = new_n17107_ & new_n21068_;
  assign new_n22112_ = new_n17107_ & new_n21079_;
  assign new_n22113_ = ~new_n22111_ & ~new_n22112_;
  assign new_n22114_ = ~new_n22110_ & new_n22113_;
  assign new_n22115_ = new_n22109_ & new_n22114_;
  assign new_n22116_ = new_n17107_ & new_n21089_;
  assign new_n22117_ = new_n17107_ & new_n21077_;
  assign new_n22118_ = new_n17107_ & new_n21087_;
  assign new_n22119_ = ~new_n22117_ & ~new_n22118_;
  assign new_n22120_ = ~new_n22116_ & new_n22119_;
  assign new_n22121_ = new_n17107_ & new_n21098_;
  assign new_n22122_ = new_n17107_ & new_n21085_;
  assign new_n22123_ = new_n17107_ & new_n21096_;
  assign new_n22124_ = ~new_n22122_ & ~new_n22123_;
  assign new_n22125_ = ~new_n22121_ & new_n22124_;
  assign new_n22126_ = new_n22120_ & new_n22125_;
  assign new_n22127_ = new_n22115_ & new_n22126_;
  assign new_n22128_ = new_n17107_ & new_n21106_;
  assign new_n22129_ = new_n17107_ & new_n21094_;
  assign new_n22130_ = new_n17107_ & new_n21104_;
  assign new_n22131_ = ~new_n22129_ & ~new_n22130_;
  assign new_n22132_ = ~new_n22128_ & new_n22131_;
  assign new_n22133_ = new_n17107_ & new_n21116_;
  assign new_n22134_ = new_n17107_ & new_n21102_;
  assign new_n22135_ = new_n17107_ & new_n21114_;
  assign new_n22136_ = ~new_n22134_ & ~new_n22135_;
  assign new_n22137_ = ~new_n22133_ & new_n22136_;
  assign new_n22138_ = new_n22132_ & new_n22137_;
  assign new_n22139_ = new_n17153_ & new_n21019_;
  assign new_n22140_ = new_n17107_ & new_n21112_;
  assign new_n22141_ = new_n17153_ & new_n21017_;
  assign new_n22142_ = ~new_n22140_ & ~new_n22141_;
  assign new_n22143_ = ~new_n22139_ & new_n22142_;
  assign new_n22144_ = new_n17153_ & new_n21015_;
  assign new_n22145_ = new_n17153_ & new_n21026_;
  assign new_n22146_ = ~new_n22144_ & ~new_n22145_;
  assign new_n22147_ = new_n22143_ & new_n22146_;
  assign new_n22148_ = new_n22138_ & new_n22147_;
  assign new_n22149_ = new_n22127_ & new_n22148_;
  assign new_n22150_ = new_n17153_ & new_n21039_;
  assign new_n22151_ = new_n17153_ & new_n21029_;
  assign new_n22152_ = new_n17153_ & new_n21024_;
  assign new_n22153_ = ~new_n22151_ & ~new_n22152_;
  assign new_n22154_ = ~new_n22150_ & new_n22153_;
  assign new_n22155_ = new_n17153_ & new_n21050_;
  assign new_n22156_ = new_n17153_ & new_n21042_;
  assign new_n22157_ = new_n17153_ & new_n21036_;
  assign new_n22158_ = ~new_n22156_ & ~new_n22157_;
  assign new_n22159_ = ~new_n22155_ & new_n22158_;
  assign new_n22160_ = new_n22154_ & new_n22159_;
  assign new_n22161_ = new_n17153_ & new_n21060_;
  assign new_n22162_ = new_n17153_ & new_n21053_;
  assign new_n22163_ = new_n17153_ & new_n21047_;
  assign new_n22164_ = ~new_n22162_ & ~new_n22163_;
  assign new_n22165_ = ~new_n22161_ & new_n22164_;
  assign new_n22166_ = new_n17153_ & new_n21066_;
  assign new_n22167_ = new_n17153_ & new_n21062_;
  assign new_n22168_ = new_n17153_ & new_n21058_;
  assign new_n22169_ = ~new_n22167_ & ~new_n22168_;
  assign new_n22170_ = ~new_n22166_ & new_n22169_;
  assign new_n22171_ = new_n22165_ & new_n22170_;
  assign new_n22172_ = new_n22160_ & new_n22171_;
  assign new_n22173_ = new_n17153_ & new_n21081_;
  assign new_n22174_ = new_n17153_ & new_n21068_;
  assign new_n22175_ = new_n17153_ & new_n21079_;
  assign new_n22176_ = ~new_n22174_ & ~new_n22175_;
  assign new_n22177_ = ~new_n22173_ & new_n22176_;
  assign new_n22178_ = new_n17153_ & new_n21089_;
  assign new_n22179_ = new_n17153_ & new_n21077_;
  assign new_n22180_ = new_n17153_ & new_n21087_;
  assign new_n22181_ = ~new_n22179_ & ~new_n22180_;
  assign new_n22182_ = ~new_n22178_ & new_n22181_;
  assign new_n22183_ = new_n22177_ & new_n22182_;
  assign new_n22184_ = new_n17153_ & new_n21098_;
  assign new_n22185_ = new_n17153_ & new_n21085_;
  assign new_n22186_ = new_n17153_ & new_n21096_;
  assign new_n22187_ = ~new_n22185_ & ~new_n22186_;
  assign new_n22188_ = ~new_n22184_ & new_n22187_;
  assign new_n22189_ = new_n17153_ & new_n21094_;
  assign new_n22190_ = new_n17153_ & new_n21104_;
  assign new_n22191_ = ~new_n22189_ & ~new_n22190_;
  assign new_n22192_ = new_n22188_ & new_n22191_;
  assign new_n22193_ = new_n22183_ & new_n22192_;
  assign new_n22194_ = new_n22172_ & new_n22193_;
  assign new_n22195_ = new_n22149_ & new_n22194_;
  assign new_n22196_ = new_n22104_ & new_n22195_;
  assign new_n22197_ = new_n22013_ & new_n22196_;
  assign new_n22198_ = new_n21830_ & new_n22197_;
  assign new_n22199_ = new_n21461_ & new_n22198_;
  assign new_n22200_ = new_n20678_ & new_n22199_;
  assign new_n22201_ = new_n17153_ & new_n21114_;
  assign new_n22202_ = new_n17153_ & new_n21106_;
  assign new_n22203_ = new_n17153_ & new_n21102_;
  assign new_n22204_ = ~new_n22202_ & ~new_n22203_;
  assign new_n22205_ = ~new_n22201_ & new_n22204_;
  assign new_n22206_ = new_n17205_ & new_n21017_;
  assign new_n22207_ = new_n17153_ & new_n21116_;
  assign new_n22208_ = new_n17153_ & new_n21112_;
  assign new_n22209_ = ~new_n22207_ & ~new_n22208_;
  assign new_n22210_ = ~new_n22206_ & new_n22209_;
  assign new_n22211_ = new_n22205_ & new_n22210_;
  assign new_n22212_ = new_n17205_ & new_n21026_;
  assign new_n22213_ = new_n17205_ & new_n21019_;
  assign new_n22214_ = new_n17205_ & new_n21015_;
  assign new_n22215_ = ~new_n22213_ & ~new_n22214_;
  assign new_n22216_ = ~new_n22212_ & new_n22215_;
  assign new_n22217_ = new_n17205_ & new_n21039_;
  assign new_n22218_ = new_n17205_ & new_n21029_;
  assign new_n22219_ = new_n17205_ & new_n21024_;
  assign new_n22220_ = ~new_n22218_ & ~new_n22219_;
  assign new_n22221_ = ~new_n22217_ & new_n22220_;
  assign new_n22222_ = new_n22216_ & new_n22221_;
  assign new_n22223_ = new_n22211_ & new_n22222_;
  assign new_n22224_ = new_n17205_ & new_n21050_;
  assign new_n22225_ = new_n17205_ & new_n21042_;
  assign new_n22226_ = new_n17205_ & new_n21036_;
  assign new_n22227_ = ~new_n22225_ & ~new_n22226_;
  assign new_n22228_ = ~new_n22224_ & new_n22227_;
  assign new_n22229_ = new_n17205_ & new_n21060_;
  assign new_n22230_ = new_n17205_ & new_n21053_;
  assign new_n22231_ = new_n17205_ & new_n21047_;
  assign new_n22232_ = ~new_n22230_ & ~new_n22231_;
  assign new_n22233_ = ~new_n22229_ & new_n22232_;
  assign new_n22234_ = new_n22228_ & new_n22233_;
  assign new_n22235_ = new_n17205_ & new_n21066_;
  assign new_n22236_ = new_n17205_ & new_n21062_;
  assign new_n22237_ = new_n17205_ & new_n21058_;
  assign new_n22238_ = ~new_n22236_ & ~new_n22237_;
  assign new_n22239_ = ~new_n22235_ & new_n22238_;
  assign new_n22240_ = new_n17205_ & new_n21081_;
  assign new_n22241_ = new_n17205_ & new_n21068_;
  assign new_n22242_ = new_n17205_ & new_n21079_;
  assign new_n22243_ = ~new_n22241_ & ~new_n22242_;
  assign new_n22244_ = ~new_n22240_ & new_n22243_;
  assign new_n22245_ = new_n22239_ & new_n22244_;
  assign new_n22246_ = new_n22234_ & new_n22245_;
  assign new_n22247_ = new_n22223_ & new_n22246_;
  assign new_n22248_ = new_n17205_ & new_n21089_;
  assign new_n22249_ = new_n17205_ & new_n21077_;
  assign new_n22250_ = new_n17205_ & new_n21087_;
  assign new_n22251_ = ~new_n22249_ & ~new_n22250_;
  assign new_n22252_ = ~new_n22248_ & new_n22251_;
  assign new_n22253_ = new_n17205_ & new_n21098_;
  assign new_n22254_ = new_n17205_ & new_n21085_;
  assign new_n22255_ = new_n17205_ & new_n21096_;
  assign new_n22256_ = ~new_n22254_ & ~new_n22255_;
  assign new_n22257_ = ~new_n22253_ & new_n22256_;
  assign new_n22258_ = new_n22252_ & new_n22257_;
  assign new_n22259_ = new_n17205_ & new_n21106_;
  assign new_n22260_ = new_n17205_ & new_n21094_;
  assign new_n22261_ = new_n17205_ & new_n21104_;
  assign new_n22262_ = ~new_n22260_ & ~new_n22261_;
  assign new_n22263_ = ~new_n22259_ & new_n22262_;
  assign new_n22264_ = new_n17205_ & new_n21116_;
  assign new_n22265_ = new_n17205_ & new_n21102_;
  assign new_n22266_ = new_n17205_ & new_n21114_;
  assign new_n22267_ = ~new_n22265_ & ~new_n22266_;
  assign new_n22268_ = ~new_n22264_ & new_n22267_;
  assign new_n22269_ = new_n22263_ & new_n22268_;
  assign new_n22270_ = new_n22258_ & new_n22269_;
  assign new_n22271_ = new_n17251_ & new_n21019_;
  assign new_n22272_ = new_n17205_ & new_n21112_;
  assign new_n22273_ = new_n17251_ & new_n21017_;
  assign new_n22274_ = ~new_n22272_ & ~new_n22273_;
  assign new_n22275_ = ~new_n22271_ & new_n22274_;
  assign new_n22276_ = new_n17251_ & new_n21029_;
  assign new_n22277_ = new_n17251_ & new_n21015_;
  assign new_n22278_ = new_n17251_ & new_n21026_;
  assign new_n22279_ = ~new_n22277_ & ~new_n22278_;
  assign new_n22280_ = ~new_n22276_ & new_n22279_;
  assign new_n22281_ = new_n22275_ & new_n22280_;
  assign new_n22282_ = new_n17251_ & new_n21042_;
  assign new_n22283_ = new_n17251_ & new_n21024_;
  assign new_n22284_ = new_n17251_ & new_n21039_;
  assign new_n22285_ = ~new_n22283_ & ~new_n22284_;
  assign new_n22286_ = ~new_n22282_ & new_n22285_;
  assign new_n22287_ = new_n17251_ & new_n21036_;
  assign new_n22288_ = new_n17251_ & new_n21050_;
  assign new_n22289_ = ~new_n22287_ & ~new_n22288_;
  assign new_n22290_ = new_n22286_ & new_n22289_;
  assign new_n22291_ = new_n22281_ & new_n22290_;
  assign new_n22292_ = new_n22270_ & new_n22291_;
  assign new_n22293_ = new_n22247_ & new_n22292_;
  assign new_n22294_ = new_n17251_ & new_n21060_;
  assign new_n22295_ = new_n17251_ & new_n21053_;
  assign new_n22296_ = new_n17251_ & new_n21047_;
  assign new_n22297_ = ~new_n22295_ & ~new_n22296_;
  assign new_n22298_ = ~new_n22294_ & new_n22297_;
  assign new_n22299_ = new_n17251_ & new_n21066_;
  assign new_n22300_ = new_n17251_ & new_n21062_;
  assign new_n22301_ = new_n17251_ & new_n21058_;
  assign new_n22302_ = ~new_n22300_ & ~new_n22301_;
  assign new_n22303_ = ~new_n22299_ & new_n22302_;
  assign new_n22304_ = new_n22298_ & new_n22303_;
  assign new_n22305_ = new_n17251_ & new_n21081_;
  assign new_n22306_ = new_n17251_ & new_n21068_;
  assign new_n22307_ = new_n17251_ & new_n21079_;
  assign new_n22308_ = ~new_n22306_ & ~new_n22307_;
  assign new_n22309_ = ~new_n22305_ & new_n22308_;
  assign new_n22310_ = new_n17251_ & new_n21089_;
  assign new_n22311_ = new_n17251_ & new_n21077_;
  assign new_n22312_ = new_n17251_ & new_n21087_;
  assign new_n22313_ = ~new_n22311_ & ~new_n22312_;
  assign new_n22314_ = ~new_n22310_ & new_n22313_;
  assign new_n22315_ = new_n22309_ & new_n22314_;
  assign new_n22316_ = new_n22304_ & new_n22315_;
  assign new_n22317_ = new_n17251_ & new_n21098_;
  assign new_n22318_ = new_n17251_ & new_n21085_;
  assign new_n22319_ = new_n17251_ & new_n21096_;
  assign new_n22320_ = ~new_n22318_ & ~new_n22319_;
  assign new_n22321_ = ~new_n22317_ & new_n22320_;
  assign new_n22322_ = new_n17251_ & new_n21106_;
  assign new_n22323_ = new_n17251_ & new_n21094_;
  assign new_n22324_ = new_n17251_ & new_n21104_;
  assign new_n22325_ = ~new_n22323_ & ~new_n22324_;
  assign new_n22326_ = ~new_n22322_ & new_n22325_;
  assign new_n22327_ = new_n22321_ & new_n22326_;
  assign new_n22328_ = new_n17251_ & new_n21116_;
  assign new_n22329_ = new_n17251_ & new_n21102_;
  assign new_n22330_ = new_n17251_ & new_n21114_;
  assign new_n22331_ = ~new_n22329_ & ~new_n22330_;
  assign new_n22332_ = ~new_n22328_ & new_n22331_;
  assign new_n22333_ = new_n17251_ & new_n21112_;
  assign new_n22334_ = new_n17364_ & new_n21017_;
  assign new_n22335_ = ~new_n22333_ & ~new_n22334_;
  assign new_n22336_ = new_n22332_ & new_n22335_;
  assign new_n22337_ = new_n22327_ & new_n22336_;
  assign new_n22338_ = new_n22316_ & new_n22337_;
  assign new_n22339_ = new_n17364_ & new_n21026_;
  assign new_n22340_ = new_n17364_ & new_n21019_;
  assign new_n22341_ = new_n17364_ & new_n21015_;
  assign new_n22342_ = ~new_n22340_ & ~new_n22341_;
  assign new_n22343_ = ~new_n22339_ & new_n22342_;
  assign new_n22344_ = new_n17364_ & new_n21039_;
  assign new_n22345_ = new_n17364_ & new_n21029_;
  assign new_n22346_ = new_n17364_ & new_n21024_;
  assign new_n22347_ = ~new_n22345_ & ~new_n22346_;
  assign new_n22348_ = ~new_n22344_ & new_n22347_;
  assign new_n22349_ = new_n22343_ & new_n22348_;
  assign new_n22350_ = new_n17364_ & new_n21050_;
  assign new_n22351_ = new_n17364_ & new_n21042_;
  assign new_n22352_ = new_n17364_ & new_n21036_;
  assign new_n22353_ = ~new_n22351_ & ~new_n22352_;
  assign new_n22354_ = ~new_n22350_ & new_n22353_;
  assign new_n22355_ = new_n17364_ & new_n21060_;
  assign new_n22356_ = new_n17364_ & new_n21053_;
  assign new_n22357_ = new_n17364_ & new_n21047_;
  assign new_n22358_ = ~new_n22356_ & ~new_n22357_;
  assign new_n22359_ = ~new_n22355_ & new_n22358_;
  assign new_n22360_ = new_n22354_ & new_n22359_;
  assign new_n22361_ = new_n22349_ & new_n22360_;
  assign new_n22362_ = new_n17364_ & new_n21066_;
  assign new_n22363_ = new_n17364_ & new_n21062_;
  assign new_n22364_ = new_n17364_ & new_n21058_;
  assign new_n22365_ = ~new_n22363_ & ~new_n22364_;
  assign new_n22366_ = ~new_n22362_ & new_n22365_;
  assign new_n22367_ = new_n17364_ & new_n21081_;
  assign new_n22368_ = new_n17364_ & new_n21068_;
  assign new_n22369_ = new_n17364_ & new_n21079_;
  assign new_n22370_ = ~new_n22368_ & ~new_n22369_;
  assign new_n22371_ = ~new_n22367_ & new_n22370_;
  assign new_n22372_ = new_n22366_ & new_n22371_;
  assign new_n22373_ = new_n17364_ & new_n21089_;
  assign new_n22374_ = new_n17364_ & new_n21077_;
  assign new_n22375_ = new_n17364_ & new_n21087_;
  assign new_n22376_ = ~new_n22374_ & ~new_n22375_;
  assign new_n22377_ = ~new_n22373_ & new_n22376_;
  assign new_n22378_ = new_n17364_ & new_n21085_;
  assign new_n22379_ = new_n17364_ & new_n21096_;
  assign new_n22380_ = ~new_n22378_ & ~new_n22379_;
  assign new_n22381_ = new_n22377_ & new_n22380_;
  assign new_n22382_ = new_n22372_ & new_n22381_;
  assign new_n22383_ = new_n22361_ & new_n22382_;
  assign new_n22384_ = new_n22338_ & new_n22383_;
  assign new_n22385_ = new_n22293_ & new_n22384_;
  assign new_n22386_ = new_n17364_ & new_n21104_;
  assign new_n22387_ = new_n17364_ & new_n21098_;
  assign new_n22388_ = new_n17364_ & new_n21094_;
  assign new_n22389_ = ~new_n22387_ & ~new_n22388_;
  assign new_n22390_ = ~new_n22386_ & new_n22389_;
  assign new_n22391_ = new_n17364_ & new_n21114_;
  assign new_n22392_ = new_n17364_ & new_n21106_;
  assign new_n22393_ = new_n17364_ & new_n21102_;
  assign new_n22394_ = ~new_n22392_ & ~new_n22393_;
  assign new_n22395_ = ~new_n22391_ & new_n22394_;
  assign new_n22396_ = new_n22390_ & new_n22395_;
  assign new_n22397_ = new_n17416_ & new_n21017_;
  assign new_n22398_ = new_n17364_ & new_n21116_;
  assign new_n22399_ = new_n17364_ & new_n21112_;
  assign new_n22400_ = ~new_n22398_ & ~new_n22399_;
  assign new_n22401_ = ~new_n22397_ & new_n22400_;
  assign new_n22402_ = new_n17416_ & new_n21026_;
  assign new_n22403_ = new_n17416_ & new_n21019_;
  assign new_n22404_ = new_n17416_ & new_n21015_;
  assign new_n22405_ = ~new_n22403_ & ~new_n22404_;
  assign new_n22406_ = ~new_n22402_ & new_n22405_;
  assign new_n22407_ = new_n22401_ & new_n22406_;
  assign new_n22408_ = new_n22396_ & new_n22407_;
  assign new_n22409_ = new_n17416_ & new_n21039_;
  assign new_n22410_ = new_n17416_ & new_n21029_;
  assign new_n22411_ = new_n17416_ & new_n21024_;
  assign new_n22412_ = ~new_n22410_ & ~new_n22411_;
  assign new_n22413_ = ~new_n22409_ & new_n22412_;
  assign new_n22414_ = new_n17416_ & new_n21050_;
  assign new_n22415_ = new_n17416_ & new_n21042_;
  assign new_n22416_ = new_n17416_ & new_n21036_;
  assign new_n22417_ = ~new_n22415_ & ~new_n22416_;
  assign new_n22418_ = ~new_n22414_ & new_n22417_;
  assign new_n22419_ = new_n22413_ & new_n22418_;
  assign new_n22420_ = new_n17416_ & new_n21060_;
  assign new_n22421_ = new_n17416_ & new_n21053_;
  assign new_n22422_ = new_n17416_ & new_n21047_;
  assign new_n22423_ = ~new_n22421_ & ~new_n22422_;
  assign new_n22424_ = ~new_n22420_ & new_n22423_;
  assign new_n22425_ = new_n17416_ & new_n21062_;
  assign new_n22426_ = new_n17416_ & new_n21058_;
  assign new_n22427_ = ~new_n22425_ & ~new_n22426_;
  assign new_n22428_ = new_n22424_ & new_n22427_;
  assign new_n22429_ = new_n22419_ & new_n22428_;
  assign new_n22430_ = new_n22408_ & new_n22429_;
  assign new_n22431_ = new_n17416_ & new_n21079_;
  assign new_n22432_ = new_n17416_ & new_n21066_;
  assign new_n22433_ = new_n17416_ & new_n21068_;
  assign new_n22434_ = ~new_n22432_ & ~new_n22433_;
  assign new_n22435_ = ~new_n22431_ & new_n22434_;
  assign new_n22436_ = new_n17416_ & new_n21087_;
  assign new_n22437_ = new_n17416_ & new_n21081_;
  assign new_n22438_ = new_n17416_ & new_n21077_;
  assign new_n22439_ = ~new_n22437_ & ~new_n22438_;
  assign new_n22440_ = ~new_n22436_ & new_n22439_;
  assign new_n22441_ = new_n22435_ & new_n22440_;
  assign new_n22442_ = new_n17416_ & new_n21096_;
  assign new_n22443_ = new_n17416_ & new_n21089_;
  assign new_n22444_ = new_n17416_ & new_n21085_;
  assign new_n22445_ = ~new_n22443_ & ~new_n22444_;
  assign new_n22446_ = ~new_n22442_ & new_n22445_;
  assign new_n22447_ = new_n17416_ & new_n21104_;
  assign new_n22448_ = new_n17416_ & new_n21098_;
  assign new_n22449_ = new_n17416_ & new_n21094_;
  assign new_n22450_ = ~new_n22448_ & ~new_n22449_;
  assign new_n22451_ = ~new_n22447_ & new_n22450_;
  assign new_n22452_ = new_n22446_ & new_n22451_;
  assign new_n22453_ = new_n22441_ & new_n22452_;
  assign new_n22454_ = new_n17416_ & new_n21114_;
  assign new_n22455_ = new_n17416_ & new_n21106_;
  assign new_n22456_ = new_n17416_ & new_n21102_;
  assign new_n22457_ = ~new_n22455_ & ~new_n22456_;
  assign new_n22458_ = ~new_n22454_ & new_n22457_;
  assign new_n22459_ = new_n17462_ & new_n21017_;
  assign new_n22460_ = new_n17416_ & new_n21116_;
  assign new_n22461_ = new_n17416_ & new_n21112_;
  assign new_n22462_ = ~new_n22460_ & ~new_n22461_;
  assign new_n22463_ = ~new_n22459_ & new_n22462_;
  assign new_n22464_ = new_n22458_ & new_n22463_;
  assign new_n22465_ = new_n17462_ & new_n21026_;
  assign new_n22466_ = new_n17462_ & new_n21019_;
  assign new_n22467_ = new_n17462_ & new_n21015_;
  assign new_n22468_ = ~new_n22466_ & ~new_n22467_;
  assign new_n22469_ = ~new_n22465_ & new_n22468_;
  assign new_n22470_ = new_n17462_ & new_n21029_;
  assign new_n22471_ = new_n17462_ & new_n21024_;
  assign new_n22472_ = ~new_n22470_ & ~new_n22471_;
  assign new_n22473_ = new_n22469_ & new_n22472_;
  assign new_n22474_ = new_n22464_ & new_n22473_;
  assign new_n22475_ = new_n22453_ & new_n22474_;
  assign new_n22476_ = new_n22430_ & new_n22475_;
  assign new_n22477_ = new_n17462_ & new_n21036_;
  assign new_n22478_ = new_n17462_ & new_n21039_;
  assign new_n22479_ = new_n17462_ & new_n21042_;
  assign new_n22480_ = ~new_n22478_ & ~new_n22479_;
  assign new_n22481_ = ~new_n22477_ & new_n22480_;
  assign new_n22482_ = new_n17462_ & new_n21047_;
  assign new_n22483_ = new_n17462_ & new_n21050_;
  assign new_n22484_ = new_n17462_ & new_n21053_;
  assign new_n22485_ = ~new_n22483_ & ~new_n22484_;
  assign new_n22486_ = ~new_n22482_ & new_n22485_;
  assign new_n22487_ = new_n22481_ & new_n22486_;
  assign new_n22488_ = new_n17462_ & new_n21058_;
  assign new_n22489_ = new_n17462_ & new_n21060_;
  assign new_n22490_ = new_n17462_ & new_n21062_;
  assign new_n22491_ = ~new_n22489_ & ~new_n22490_;
  assign new_n22492_ = ~new_n22488_ & new_n22491_;
  assign new_n22493_ = new_n17462_ & new_n21079_;
  assign new_n22494_ = new_n17462_ & new_n21066_;
  assign new_n22495_ = new_n17462_ & new_n21068_;
  assign new_n22496_ = ~new_n22494_ & ~new_n22495_;
  assign new_n22497_ = ~new_n22493_ & new_n22496_;
  assign new_n22498_ = new_n22492_ & new_n22497_;
  assign new_n22499_ = new_n22487_ & new_n22498_;
  assign new_n22500_ = new_n17462_ & new_n21087_;
  assign new_n22501_ = new_n17462_ & new_n21081_;
  assign new_n22502_ = new_n17462_ & new_n21077_;
  assign new_n22503_ = ~new_n22501_ & ~new_n22502_;
  assign new_n22504_ = ~new_n22500_ & new_n22503_;
  assign new_n22505_ = new_n17462_ & new_n21096_;
  assign new_n22506_ = new_n17462_ & new_n21089_;
  assign new_n22507_ = new_n17462_ & new_n21085_;
  assign new_n22508_ = ~new_n22506_ & ~new_n22507_;
  assign new_n22509_ = ~new_n22505_ & new_n22508_;
  assign new_n22510_ = new_n22504_ & new_n22509_;
  assign new_n22511_ = new_n17462_ & new_n21104_;
  assign new_n22512_ = new_n17462_ & new_n21098_;
  assign new_n22513_ = new_n17462_ & new_n21094_;
  assign new_n22514_ = ~new_n22512_ & ~new_n22513_;
  assign new_n22515_ = ~new_n22511_ & new_n22514_;
  assign new_n22516_ = new_n17462_ & new_n21106_;
  assign new_n22517_ = new_n17462_ & new_n21102_;
  assign new_n22518_ = ~new_n22516_ & ~new_n22517_;
  assign new_n22519_ = new_n22515_ & new_n22518_;
  assign new_n22520_ = new_n22510_ & new_n22519_;
  assign new_n22521_ = new_n22499_ & new_n22520_;
  assign new_n22522_ = new_n17462_ & new_n21112_;
  assign new_n22523_ = new_n17462_ & new_n21114_;
  assign new_n22524_ = new_n17462_ & new_n21116_;
  assign new_n22525_ = ~new_n22523_ & ~new_n22524_;
  assign new_n22526_ = ~new_n22522_ & new_n22525_;
  assign new_n22527_ = new_n17510_ & new_n21015_;
  assign new_n22528_ = new_n17510_ & new_n21017_;
  assign new_n22529_ = new_n17510_ & new_n21019_;
  assign new_n22530_ = ~new_n22528_ & ~new_n22529_;
  assign new_n22531_ = ~new_n22527_ & new_n22530_;
  assign new_n22532_ = new_n22526_ & new_n22531_;
  assign new_n22533_ = new_n17510_ & new_n21024_;
  assign new_n22534_ = new_n17510_ & new_n21026_;
  assign new_n22535_ = new_n17510_ & new_n21029_;
  assign new_n22536_ = ~new_n22534_ & ~new_n22535_;
  assign new_n22537_ = ~new_n22533_ & new_n22536_;
  assign new_n22538_ = new_n17510_ & new_n21036_;
  assign new_n22539_ = new_n17510_ & new_n21039_;
  assign new_n22540_ = new_n17510_ & new_n21042_;
  assign new_n22541_ = ~new_n22539_ & ~new_n22540_;
  assign new_n22542_ = ~new_n22538_ & new_n22541_;
  assign new_n22543_ = new_n22537_ & new_n22542_;
  assign new_n22544_ = new_n22532_ & new_n22543_;
  assign new_n22545_ = new_n17510_ & new_n21047_;
  assign new_n22546_ = new_n17510_ & new_n21050_;
  assign new_n22547_ = new_n17510_ & new_n21053_;
  assign new_n22548_ = ~new_n22546_ & ~new_n22547_;
  assign new_n22549_ = ~new_n22545_ & new_n22548_;
  assign new_n22550_ = new_n17510_ & new_n21058_;
  assign new_n22551_ = new_n17510_ & new_n21060_;
  assign new_n22552_ = new_n17510_ & new_n21062_;
  assign new_n22553_ = ~new_n22551_ & ~new_n22552_;
  assign new_n22554_ = ~new_n22550_ & new_n22553_;
  assign new_n22555_ = new_n22549_ & new_n22554_;
  assign new_n22556_ = new_n17510_ & new_n21079_;
  assign new_n22557_ = new_n17510_ & new_n21066_;
  assign new_n22558_ = new_n17510_ & new_n21068_;
  assign new_n22559_ = ~new_n22557_ & ~new_n22558_;
  assign new_n22560_ = ~new_n22556_ & new_n22559_;
  assign new_n22561_ = new_n17510_ & new_n21081_;
  assign new_n22562_ = new_n17510_ & new_n21077_;
  assign new_n22563_ = ~new_n22561_ & ~new_n22562_;
  assign new_n22564_ = new_n22560_ & new_n22563_;
  assign new_n22565_ = new_n22555_ & new_n22564_;
  assign new_n22566_ = new_n22544_ & new_n22565_;
  assign new_n22567_ = new_n22521_ & new_n22566_;
  assign new_n22568_ = new_n22476_ & new_n22567_;
  assign new_n22569_ = new_n22385_ & new_n22568_;
  assign new_n22570_ = new_n17510_ & new_n21085_;
  assign new_n22571_ = new_n17510_ & new_n21087_;
  assign new_n22572_ = new_n17510_ & new_n21089_;
  assign new_n22573_ = ~new_n22571_ & ~new_n22572_;
  assign new_n22574_ = ~new_n22570_ & new_n22573_;
  assign new_n22575_ = new_n17510_ & new_n21094_;
  assign new_n22576_ = new_n17510_ & new_n21096_;
  assign new_n22577_ = new_n17510_ & new_n21098_;
  assign new_n22578_ = ~new_n22576_ & ~new_n22577_;
  assign new_n22579_ = ~new_n22575_ & new_n22578_;
  assign new_n22580_ = new_n22574_ & new_n22579_;
  assign new_n22581_ = new_n17510_ & new_n21102_;
  assign new_n22582_ = new_n17510_ & new_n21104_;
  assign new_n22583_ = new_n17510_ & new_n21106_;
  assign new_n22584_ = ~new_n22582_ & ~new_n22583_;
  assign new_n22585_ = ~new_n22581_ & new_n22584_;
  assign new_n22586_ = new_n17510_ & new_n21112_;
  assign new_n22587_ = new_n17510_ & new_n21114_;
  assign new_n22588_ = new_n17510_ & new_n21116_;
  assign new_n22589_ = ~new_n22587_ & ~new_n22588_;
  assign new_n22590_ = ~new_n22586_ & new_n22589_;
  assign new_n22591_ = new_n22585_ & new_n22590_;
  assign new_n22592_ = new_n22580_ & new_n22591_;
  assign new_n22593_ = new_n17625_ & new_n21015_;
  assign new_n22594_ = new_n17625_ & new_n21017_;
  assign new_n22595_ = new_n17625_ & new_n21019_;
  assign new_n22596_ = ~new_n22594_ & ~new_n22595_;
  assign new_n22597_ = ~new_n22593_ & new_n22596_;
  assign new_n22598_ = new_n17625_ & new_n21024_;
  assign new_n22599_ = new_n17625_ & new_n21026_;
  assign new_n22600_ = new_n17625_ & new_n21029_;
  assign new_n22601_ = ~new_n22599_ & ~new_n22600_;
  assign new_n22602_ = ~new_n22598_ & new_n22601_;
  assign new_n22603_ = new_n22597_ & new_n22602_;
  assign new_n22604_ = new_n17625_ & new_n21036_;
  assign new_n22605_ = new_n17625_ & new_n21039_;
  assign new_n22606_ = new_n17625_ & new_n21042_;
  assign new_n22607_ = ~new_n22605_ & ~new_n22606_;
  assign new_n22608_ = ~new_n22604_ & new_n22607_;
  assign new_n22609_ = new_n17625_ & new_n21047_;
  assign new_n22610_ = new_n17625_ & new_n21050_;
  assign new_n22611_ = new_n17625_ & new_n21053_;
  assign new_n22612_ = ~new_n22610_ & ~new_n22611_;
  assign new_n22613_ = ~new_n22609_ & new_n22612_;
  assign new_n22614_ = new_n22608_ & new_n22613_;
  assign new_n22615_ = new_n22603_ & new_n22614_;
  assign new_n22616_ = new_n22592_ & new_n22615_;
  assign new_n22617_ = new_n17625_ & new_n21058_;
  assign new_n22618_ = new_n17625_ & new_n21060_;
  assign new_n22619_ = new_n17625_ & new_n21062_;
  assign new_n22620_ = ~new_n22618_ & ~new_n22619_;
  assign new_n22621_ = ~new_n22617_ & new_n22620_;
  assign new_n22622_ = new_n17625_ & new_n21079_;
  assign new_n22623_ = new_n17625_ & new_n21066_;
  assign new_n22624_ = new_n17625_ & new_n21068_;
  assign new_n22625_ = ~new_n22623_ & ~new_n22624_;
  assign new_n22626_ = ~new_n22622_ & new_n22625_;
  assign new_n22627_ = new_n22621_ & new_n22626_;
  assign new_n22628_ = new_n17625_ & new_n21087_;
  assign new_n22629_ = new_n17625_ & new_n21081_;
  assign new_n22630_ = new_n17625_ & new_n21077_;
  assign new_n22631_ = ~new_n22629_ & ~new_n22630_;
  assign new_n22632_ = ~new_n22628_ & new_n22631_;
  assign new_n22633_ = new_n17625_ & new_n21096_;
  assign new_n22634_ = new_n17625_ & new_n21089_;
  assign new_n22635_ = new_n17625_ & new_n21085_;
  assign new_n22636_ = ~new_n22634_ & ~new_n22635_;
  assign new_n22637_ = ~new_n22633_ & new_n22636_;
  assign new_n22638_ = new_n22632_ & new_n22637_;
  assign new_n22639_ = new_n22627_ & new_n22638_;
  assign new_n22640_ = new_n17625_ & new_n21104_;
  assign new_n22641_ = new_n17625_ & new_n21098_;
  assign new_n22642_ = new_n17625_ & new_n21094_;
  assign new_n22643_ = ~new_n22641_ & ~new_n22642_;
  assign new_n22644_ = ~new_n22640_ & new_n22643_;
  assign new_n22645_ = new_n17625_ & new_n21114_;
  assign new_n22646_ = new_n17625_ & new_n21106_;
  assign new_n22647_ = new_n17625_ & new_n21102_;
  assign new_n22648_ = ~new_n22646_ & ~new_n22647_;
  assign new_n22649_ = ~new_n22645_ & new_n22648_;
  assign new_n22650_ = new_n22644_ & new_n22649_;
  assign new_n22651_ = new_n17676_ & new_n21017_;
  assign new_n22652_ = new_n17625_ & new_n21116_;
  assign new_n22653_ = new_n17625_ & new_n21112_;
  assign new_n22654_ = ~new_n22652_ & ~new_n22653_;
  assign new_n22655_ = ~new_n22651_ & new_n22654_;
  assign new_n22656_ = new_n17676_ & new_n21019_;
  assign new_n22657_ = new_n17676_ & new_n21015_;
  assign new_n22658_ = ~new_n22656_ & ~new_n22657_;
  assign new_n22659_ = new_n22655_ & new_n22658_;
  assign new_n22660_ = new_n22650_ & new_n22659_;
  assign new_n22661_ = new_n22639_ & new_n22660_;
  assign new_n22662_ = new_n22616_ & new_n22661_;
  assign new_n22663_ = new_n17676_ & new_n21024_;
  assign new_n22664_ = new_n17676_ & new_n21026_;
  assign new_n22665_ = new_n17676_ & new_n21029_;
  assign new_n22666_ = ~new_n22664_ & ~new_n22665_;
  assign new_n22667_ = ~new_n22663_ & new_n22666_;
  assign new_n22668_ = new_n17676_ & new_n21036_;
  assign new_n22669_ = new_n17676_ & new_n21039_;
  assign new_n22670_ = new_n17676_ & new_n21042_;
  assign new_n22671_ = ~new_n22669_ & ~new_n22670_;
  assign new_n22672_ = ~new_n22668_ & new_n22671_;
  assign new_n22673_ = new_n22667_ & new_n22672_;
  assign new_n22674_ = new_n17676_ & new_n21047_;
  assign new_n22675_ = new_n17676_ & new_n21050_;
  assign new_n22676_ = new_n17676_ & new_n21053_;
  assign new_n22677_ = ~new_n22675_ & ~new_n22676_;
  assign new_n22678_ = ~new_n22674_ & new_n22677_;
  assign new_n22679_ = new_n17676_ & new_n21058_;
  assign new_n22680_ = new_n17676_ & new_n21060_;
  assign new_n22681_ = new_n17676_ & new_n21062_;
  assign new_n22682_ = ~new_n22680_ & ~new_n22681_;
  assign new_n22683_ = ~new_n22679_ & new_n22682_;
  assign new_n22684_ = new_n22678_ & new_n22683_;
  assign new_n22685_ = new_n22673_ & new_n22684_;
  assign new_n22686_ = new_n17676_ & new_n21079_;
  assign new_n22687_ = new_n17676_ & new_n21066_;
  assign new_n22688_ = new_n17676_ & new_n21068_;
  assign new_n22689_ = ~new_n22687_ & ~new_n22688_;
  assign new_n22690_ = ~new_n22686_ & new_n22689_;
  assign new_n22691_ = new_n17676_ & new_n21087_;
  assign new_n22692_ = new_n17676_ & new_n21081_;
  assign new_n22693_ = new_n17676_ & new_n21077_;
  assign new_n22694_ = ~new_n22692_ & ~new_n22693_;
  assign new_n22695_ = ~new_n22691_ & new_n22694_;
  assign new_n22696_ = new_n22690_ & new_n22695_;
  assign new_n22697_ = new_n17676_ & new_n21096_;
  assign new_n22698_ = new_n17676_ & new_n21089_;
  assign new_n22699_ = new_n17676_ & new_n21085_;
  assign new_n22700_ = ~new_n22698_ & ~new_n22699_;
  assign new_n22701_ = ~new_n22697_ & new_n22700_;
  assign new_n22702_ = new_n17676_ & new_n21098_;
  assign new_n22703_ = new_n17676_ & new_n21094_;
  assign new_n22704_ = ~new_n22702_ & ~new_n22703_;
  assign new_n22705_ = new_n22701_ & new_n22704_;
  assign new_n22706_ = new_n22696_ & new_n22705_;
  assign new_n22707_ = new_n22685_ & new_n22706_;
  assign new_n22708_ = new_n17676_ & new_n21102_;
  assign new_n22709_ = new_n17676_ & new_n21104_;
  assign new_n22710_ = new_n17676_ & new_n21106_;
  assign new_n22711_ = ~new_n22709_ & ~new_n22710_;
  assign new_n22712_ = ~new_n22708_ & new_n22711_;
  assign new_n22713_ = new_n17676_ & new_n21112_;
  assign new_n22714_ = new_n17676_ & new_n21114_;
  assign new_n22715_ = new_n17676_ & new_n21116_;
  assign new_n22716_ = ~new_n22714_ & ~new_n22715_;
  assign new_n22717_ = ~new_n22713_ & new_n22716_;
  assign new_n22718_ = new_n22712_ & new_n22717_;
  assign new_n22719_ = new_n17724_ & new_n21015_;
  assign new_n22720_ = new_n17724_ & new_n21017_;
  assign new_n22721_ = new_n17724_ & new_n21019_;
  assign new_n22722_ = ~new_n22720_ & ~new_n22721_;
  assign new_n22723_ = ~new_n22719_ & new_n22722_;
  assign new_n22724_ = new_n17724_ & new_n21024_;
  assign new_n22725_ = new_n17724_ & new_n21026_;
  assign new_n22726_ = new_n17724_ & new_n21029_;
  assign new_n22727_ = ~new_n22725_ & ~new_n22726_;
  assign new_n22728_ = ~new_n22724_ & new_n22727_;
  assign new_n22729_ = new_n22723_ & new_n22728_;
  assign new_n22730_ = new_n22718_ & new_n22729_;
  assign new_n22731_ = new_n17724_ & new_n21036_;
  assign new_n22732_ = new_n17724_ & new_n21039_;
  assign new_n22733_ = new_n17724_ & new_n21042_;
  assign new_n22734_ = ~new_n22732_ & ~new_n22733_;
  assign new_n22735_ = ~new_n22731_ & new_n22734_;
  assign new_n22736_ = new_n17724_ & new_n21047_;
  assign new_n22737_ = new_n17724_ & new_n21050_;
  assign new_n22738_ = new_n17724_ & new_n21053_;
  assign new_n22739_ = ~new_n22737_ & ~new_n22738_;
  assign new_n22740_ = ~new_n22736_ & new_n22739_;
  assign new_n22741_ = new_n22735_ & new_n22740_;
  assign new_n22742_ = new_n17724_ & new_n21058_;
  assign new_n22743_ = new_n17724_ & new_n21060_;
  assign new_n22744_ = new_n17724_ & new_n21062_;
  assign new_n22745_ = ~new_n22743_ & ~new_n22744_;
  assign new_n22746_ = ~new_n22742_ & new_n22745_;
  assign new_n22747_ = new_n17724_ & new_n21066_;
  assign new_n22748_ = new_n17724_ & new_n21068_;
  assign new_n22749_ = ~new_n22747_ & ~new_n22748_;
  assign new_n22750_ = new_n22746_ & new_n22749_;
  assign new_n22751_ = new_n22741_ & new_n22750_;
  assign new_n22752_ = new_n22730_ & new_n22751_;
  assign new_n22753_ = new_n22707_ & new_n22752_;
  assign new_n22754_ = new_n22662_ & new_n22753_;
  assign new_n22755_ = new_n17724_ & new_n21077_;
  assign new_n22756_ = new_n17724_ & new_n21079_;
  assign new_n22757_ = new_n17724_ & new_n21081_;
  assign new_n22758_ = ~new_n22756_ & ~new_n22757_;
  assign new_n22759_ = ~new_n22755_ & new_n22758_;
  assign new_n22760_ = new_n17724_ & new_n21085_;
  assign new_n22761_ = new_n17724_ & new_n21087_;
  assign new_n22762_ = new_n17724_ & new_n21089_;
  assign new_n22763_ = ~new_n22761_ & ~new_n22762_;
  assign new_n22764_ = ~new_n22760_ & new_n22763_;
  assign new_n22765_ = new_n22759_ & new_n22764_;
  assign new_n22766_ = new_n17724_ & new_n21094_;
  assign new_n22767_ = new_n17724_ & new_n21096_;
  assign new_n22768_ = new_n17724_ & new_n21098_;
  assign new_n22769_ = ~new_n22767_ & ~new_n22768_;
  assign new_n22770_ = ~new_n22766_ & new_n22769_;
  assign new_n22771_ = new_n17724_ & new_n21102_;
  assign new_n22772_ = new_n17724_ & new_n21104_;
  assign new_n22773_ = new_n17724_ & new_n21106_;
  assign new_n22774_ = ~new_n22772_ & ~new_n22773_;
  assign new_n22775_ = ~new_n22771_ & new_n22774_;
  assign new_n22776_ = new_n22770_ & new_n22775_;
  assign new_n22777_ = new_n22765_ & new_n22776_;
  assign new_n22778_ = new_n17724_ & new_n21112_;
  assign new_n22779_ = new_n17724_ & new_n21114_;
  assign new_n22780_ = new_n17724_ & new_n21116_;
  assign new_n22781_ = ~new_n22779_ & ~new_n22780_;
  assign new_n22782_ = ~new_n22778_ & new_n22781_;
  assign new_n22783_ = new_n17777_ & new_n21015_;
  assign new_n22784_ = new_n17777_ & new_n21017_;
  assign new_n22785_ = new_n17777_ & new_n21019_;
  assign new_n22786_ = ~new_n22784_ & ~new_n22785_;
  assign new_n22787_ = ~new_n22783_ & new_n22786_;
  assign new_n22788_ = new_n22782_ & new_n22787_;
  assign new_n22789_ = new_n17777_ & new_n21024_;
  assign new_n22790_ = new_n17777_ & new_n21026_;
  assign new_n22791_ = new_n17777_ & new_n21029_;
  assign new_n22792_ = ~new_n22790_ & ~new_n22791_;
  assign new_n22793_ = ~new_n22789_ & new_n22792_;
  assign new_n22794_ = new_n17777_ & new_n21039_;
  assign new_n22795_ = new_n17777_ & new_n21042_;
  assign new_n22796_ = ~new_n22794_ & ~new_n22795_;
  assign new_n22797_ = new_n22793_ & new_n22796_;
  assign new_n22798_ = new_n22788_ & new_n22797_;
  assign new_n22799_ = new_n22777_ & new_n22798_;
  assign new_n22800_ = new_n17777_ & new_n21053_;
  assign new_n22801_ = new_n17777_ & new_n21036_;
  assign new_n22802_ = new_n17777_ & new_n21050_;
  assign new_n22803_ = ~new_n22801_ & ~new_n22802_;
  assign new_n22804_ = ~new_n22800_ & new_n22803_;
  assign new_n22805_ = new_n17777_ & new_n21062_;
  assign new_n22806_ = new_n17777_ & new_n21047_;
  assign new_n22807_ = new_n17777_ & new_n21060_;
  assign new_n22808_ = ~new_n22806_ & ~new_n22807_;
  assign new_n22809_ = ~new_n22805_ & new_n22808_;
  assign new_n22810_ = new_n22804_ & new_n22809_;
  assign new_n22811_ = new_n17777_ & new_n21068_;
  assign new_n22812_ = new_n17777_ & new_n21058_;
  assign new_n22813_ = new_n17777_ & new_n21066_;
  assign new_n22814_ = ~new_n22812_ & ~new_n22813_;
  assign new_n22815_ = ~new_n22811_ & new_n22814_;
  assign new_n22816_ = new_n17777_ & new_n21077_;
  assign new_n22817_ = new_n17777_ & new_n21079_;
  assign new_n22818_ = new_n17777_ & new_n21081_;
  assign new_n22819_ = ~new_n22817_ & ~new_n22818_;
  assign new_n22820_ = ~new_n22816_ & new_n22819_;
  assign new_n22821_ = new_n22815_ & new_n22820_;
  assign new_n22822_ = new_n22810_ & new_n22821_;
  assign new_n22823_ = new_n17777_ & new_n21085_;
  assign new_n22824_ = new_n17777_ & new_n21087_;
  assign new_n22825_ = new_n17777_ & new_n21089_;
  assign new_n22826_ = ~new_n22824_ & ~new_n22825_;
  assign new_n22827_ = ~new_n22823_ & new_n22826_;
  assign new_n22828_ = new_n17777_ & new_n21094_;
  assign new_n22829_ = new_n17777_ & new_n21096_;
  assign new_n22830_ = new_n17777_ & new_n21098_;
  assign new_n22831_ = ~new_n22829_ & ~new_n22830_;
  assign new_n22832_ = ~new_n22828_ & new_n22831_;
  assign new_n22833_ = new_n22827_ & new_n22832_;
  assign new_n22834_ = new_n17777_ & new_n21102_;
  assign new_n22835_ = new_n17777_ & new_n21104_;
  assign new_n22836_ = new_n17777_ & new_n21106_;
  assign new_n22837_ = ~new_n22835_ & ~new_n22836_;
  assign new_n22838_ = ~new_n22834_ & new_n22837_;
  assign new_n22839_ = new_n17777_ & new_n21114_;
  assign new_n22840_ = new_n17777_ & new_n21116_;
  assign new_n22841_ = ~new_n22839_ & ~new_n22840_;
  assign new_n22842_ = new_n22838_ & new_n22841_;
  assign new_n22843_ = new_n22833_ & new_n22842_;
  assign new_n22844_ = new_n22822_ & new_n22843_;
  assign new_n22845_ = new_n22799_ & new_n22844_;
  assign new_n22846_ = new_n17888_ & new_n21019_;
  assign new_n22847_ = new_n17777_ & new_n21112_;
  assign new_n22848_ = new_n17888_ & new_n21017_;
  assign new_n22849_ = ~new_n22847_ & ~new_n22848_;
  assign new_n22850_ = ~new_n22846_ & new_n22849_;
  assign new_n22851_ = new_n17888_ & new_n21029_;
  assign new_n22852_ = new_n17888_ & new_n21015_;
  assign new_n22853_ = new_n17888_ & new_n21026_;
  assign new_n22854_ = ~new_n22852_ & ~new_n22853_;
  assign new_n22855_ = ~new_n22851_ & new_n22854_;
  assign new_n22856_ = new_n22850_ & new_n22855_;
  assign new_n22857_ = new_n17888_ & new_n21042_;
  assign new_n22858_ = new_n17888_ & new_n21024_;
  assign new_n22859_ = new_n17888_ & new_n21039_;
  assign new_n22860_ = ~new_n22858_ & ~new_n22859_;
  assign new_n22861_ = ~new_n22857_ & new_n22860_;
  assign new_n22862_ = new_n17888_ & new_n21053_;
  assign new_n22863_ = new_n17888_ & new_n21036_;
  assign new_n22864_ = new_n17888_ & new_n21050_;
  assign new_n22865_ = ~new_n22863_ & ~new_n22864_;
  assign new_n22866_ = ~new_n22862_ & new_n22865_;
  assign new_n22867_ = new_n22861_ & new_n22866_;
  assign new_n22868_ = new_n22856_ & new_n22867_;
  assign new_n22869_ = new_n17888_ & new_n21062_;
  assign new_n22870_ = new_n17888_ & new_n21047_;
  assign new_n22871_ = new_n17888_ & new_n21060_;
  assign new_n22872_ = ~new_n22870_ & ~new_n22871_;
  assign new_n22873_ = ~new_n22869_ & new_n22872_;
  assign new_n22874_ = new_n17888_ & new_n21068_;
  assign new_n22875_ = new_n17888_ & new_n21058_;
  assign new_n22876_ = new_n17888_ & new_n21066_;
  assign new_n22877_ = ~new_n22875_ & ~new_n22876_;
  assign new_n22878_ = ~new_n22874_ & new_n22877_;
  assign new_n22879_ = new_n22873_ & new_n22878_;
  assign new_n22880_ = new_n17888_ & new_n21077_;
  assign new_n22881_ = new_n17888_ & new_n21079_;
  assign new_n22882_ = new_n17888_ & new_n21081_;
  assign new_n22883_ = ~new_n22881_ & ~new_n22882_;
  assign new_n22884_ = ~new_n22880_ & new_n22883_;
  assign new_n22885_ = new_n17888_ & new_n21087_;
  assign new_n22886_ = new_n17888_ & new_n21089_;
  assign new_n22887_ = ~new_n22885_ & ~new_n22886_;
  assign new_n22888_ = new_n22884_ & new_n22887_;
  assign new_n22889_ = new_n22879_ & new_n22888_;
  assign new_n22890_ = new_n22868_ & new_n22889_;
  assign new_n22891_ = new_n17888_ & new_n21098_;
  assign new_n22892_ = new_n17888_ & new_n21085_;
  assign new_n22893_ = new_n17888_ & new_n21096_;
  assign new_n22894_ = ~new_n22892_ & ~new_n22893_;
  assign new_n22895_ = ~new_n22891_ & new_n22894_;
  assign new_n22896_ = new_n17888_ & new_n21106_;
  assign new_n22897_ = new_n17888_ & new_n21094_;
  assign new_n22898_ = new_n17888_ & new_n21104_;
  assign new_n22899_ = ~new_n22897_ & ~new_n22898_;
  assign new_n22900_ = ~new_n22896_ & new_n22899_;
  assign new_n22901_ = new_n22895_ & new_n22900_;
  assign new_n22902_ = new_n17888_ & new_n21116_;
  assign new_n22903_ = new_n17888_ & new_n21102_;
  assign new_n22904_ = new_n17888_ & new_n21114_;
  assign new_n22905_ = ~new_n22903_ & ~new_n22904_;
  assign new_n22906_ = ~new_n22902_ & new_n22905_;
  assign new_n22907_ = new_n17934_ & new_n21019_;
  assign new_n22908_ = new_n17888_ & new_n21112_;
  assign new_n22909_ = new_n17934_ & new_n21017_;
  assign new_n22910_ = ~new_n22908_ & ~new_n22909_;
  assign new_n22911_ = ~new_n22907_ & new_n22910_;
  assign new_n22912_ = new_n22906_ & new_n22911_;
  assign new_n22913_ = new_n22901_ & new_n22912_;
  assign new_n22914_ = new_n17934_ & new_n21029_;
  assign new_n22915_ = new_n17934_ & new_n21015_;
  assign new_n22916_ = new_n17934_ & new_n21026_;
  assign new_n22917_ = ~new_n22915_ & ~new_n22916_;
  assign new_n22918_ = ~new_n22914_ & new_n22917_;
  assign new_n22919_ = new_n17934_ & new_n21042_;
  assign new_n22920_ = new_n17934_ & new_n21024_;
  assign new_n22921_ = new_n17934_ & new_n21039_;
  assign new_n22922_ = ~new_n22920_ & ~new_n22921_;
  assign new_n22923_ = ~new_n22919_ & new_n22922_;
  assign new_n22924_ = new_n22918_ & new_n22923_;
  assign new_n22925_ = new_n17934_ & new_n21053_;
  assign new_n22926_ = new_n17934_ & new_n21036_;
  assign new_n22927_ = new_n17934_ & new_n21050_;
  assign new_n22928_ = ~new_n22926_ & ~new_n22927_;
  assign new_n22929_ = ~new_n22925_ & new_n22928_;
  assign new_n22930_ = new_n17934_ & new_n21047_;
  assign new_n22931_ = new_n17934_ & new_n21060_;
  assign new_n22932_ = ~new_n22930_ & ~new_n22931_;
  assign new_n22933_ = new_n22929_ & new_n22932_;
  assign new_n22934_ = new_n22924_ & new_n22933_;
  assign new_n22935_ = new_n22913_ & new_n22934_;
  assign new_n22936_ = new_n22890_ & new_n22935_;
  assign new_n22937_ = new_n22845_ & new_n22936_;
  assign new_n22938_ = new_n22754_ & new_n22937_;
  assign new_n22939_ = new_n22569_ & new_n22938_;
  assign new_n22940_ = new_n17934_ & new_n21066_;
  assign new_n22941_ = new_n17934_ & new_n21062_;
  assign new_n22942_ = new_n17934_ & new_n21058_;
  assign new_n22943_ = ~new_n22941_ & ~new_n22942_;
  assign new_n22944_ = ~new_n22940_ & new_n22943_;
  assign new_n22945_ = new_n17934_ & new_n21081_;
  assign new_n22946_ = new_n17934_ & new_n21068_;
  assign new_n22947_ = new_n17934_ & new_n21079_;
  assign new_n22948_ = ~new_n22946_ & ~new_n22947_;
  assign new_n22949_ = ~new_n22945_ & new_n22948_;
  assign new_n22950_ = new_n22944_ & new_n22949_;
  assign new_n22951_ = new_n17934_ & new_n21089_;
  assign new_n22952_ = new_n17934_ & new_n21077_;
  assign new_n22953_ = new_n17934_ & new_n21087_;
  assign new_n22954_ = ~new_n22952_ & ~new_n22953_;
  assign new_n22955_ = ~new_n22951_ & new_n22954_;
  assign new_n22956_ = new_n17934_ & new_n21098_;
  assign new_n22957_ = new_n17934_ & new_n21085_;
  assign new_n22958_ = new_n17934_ & new_n21096_;
  assign new_n22959_ = ~new_n22957_ & ~new_n22958_;
  assign new_n22960_ = ~new_n22956_ & new_n22959_;
  assign new_n22961_ = new_n22955_ & new_n22960_;
  assign new_n22962_ = new_n22950_ & new_n22961_;
  assign new_n22963_ = new_n17934_ & new_n21106_;
  assign new_n22964_ = new_n17934_ & new_n21094_;
  assign new_n22965_ = new_n17934_ & new_n21104_;
  assign new_n22966_ = ~new_n22964_ & ~new_n22965_;
  assign new_n22967_ = ~new_n22963_ & new_n22966_;
  assign new_n22968_ = new_n17934_ & new_n21116_;
  assign new_n22969_ = new_n17934_ & new_n21102_;
  assign new_n22970_ = new_n17934_ & new_n21114_;
  assign new_n22971_ = ~new_n22969_ & ~new_n22970_;
  assign new_n22972_ = ~new_n22968_ & new_n22971_;
  assign new_n22973_ = new_n22967_ & new_n22972_;
  assign new_n22974_ = new_n17987_ & new_n21019_;
  assign new_n22975_ = new_n17934_ & new_n21112_;
  assign new_n22976_ = new_n17987_ & new_n21017_;
  assign new_n22977_ = ~new_n22975_ & ~new_n22976_;
  assign new_n22978_ = ~new_n22974_ & new_n22977_;
  assign new_n22979_ = new_n17987_ & new_n21029_;
  assign new_n22980_ = new_n17987_ & new_n21015_;
  assign new_n22981_ = new_n17987_ & new_n21026_;
  assign new_n22982_ = ~new_n22980_ & ~new_n22981_;
  assign new_n22983_ = ~new_n22979_ & new_n22982_;
  assign new_n22984_ = new_n22978_ & new_n22983_;
  assign new_n22985_ = new_n22973_ & new_n22984_;
  assign new_n22986_ = new_n22962_ & new_n22985_;
  assign new_n22987_ = new_n17987_ & new_n21042_;
  assign new_n22988_ = new_n17987_ & new_n21024_;
  assign new_n22989_ = new_n17987_ & new_n21039_;
  assign new_n22990_ = ~new_n22988_ & ~new_n22989_;
  assign new_n22991_ = ~new_n22987_ & new_n22990_;
  assign new_n22992_ = new_n17987_ & new_n21053_;
  assign new_n22993_ = new_n17987_ & new_n21036_;
  assign new_n22994_ = new_n17987_ & new_n21050_;
  assign new_n22995_ = ~new_n22993_ & ~new_n22994_;
  assign new_n22996_ = ~new_n22992_ & new_n22995_;
  assign new_n22997_ = new_n22991_ & new_n22996_;
  assign new_n22998_ = new_n17987_ & new_n21062_;
  assign new_n22999_ = new_n17987_ & new_n21047_;
  assign new_n23000_ = new_n17987_ & new_n21060_;
  assign new_n23001_ = ~new_n22999_ & ~new_n23000_;
  assign new_n23002_ = ~new_n22998_ & new_n23001_;
  assign new_n23003_ = new_n17987_ & new_n21068_;
  assign new_n23004_ = new_n17987_ & new_n21058_;
  assign new_n23005_ = new_n17987_ & new_n21066_;
  assign new_n23006_ = ~new_n23004_ & ~new_n23005_;
  assign new_n23007_ = ~new_n23003_ & new_n23006_;
  assign new_n23008_ = new_n23002_ & new_n23007_;
  assign new_n23009_ = new_n22997_ & new_n23008_;
  assign new_n23010_ = new_n17987_ & new_n21077_;
  assign new_n23011_ = new_n17987_ & new_n21079_;
  assign new_n23012_ = new_n17987_ & new_n21081_;
  assign new_n23013_ = ~new_n23011_ & ~new_n23012_;
  assign new_n23014_ = ~new_n23010_ & new_n23013_;
  assign new_n23015_ = new_n17987_ & new_n21085_;
  assign new_n23016_ = new_n17987_ & new_n21087_;
  assign new_n23017_ = new_n17987_ & new_n21089_;
  assign new_n23018_ = ~new_n23016_ & ~new_n23017_;
  assign new_n23019_ = ~new_n23015_ & new_n23018_;
  assign new_n23020_ = new_n23014_ & new_n23019_;
  assign new_n23021_ = new_n17987_ & new_n21094_;
  assign new_n23022_ = new_n17987_ & new_n21096_;
  assign new_n23023_ = new_n17987_ & new_n21098_;
  assign new_n23024_ = ~new_n23022_ & ~new_n23023_;
  assign new_n23025_ = ~new_n23021_ & new_n23024_;
  assign new_n23026_ = new_n17987_ & new_n21104_;
  assign new_n23027_ = new_n17987_ & new_n21106_;
  assign new_n23028_ = ~new_n23026_ & ~new_n23027_;
  assign new_n23029_ = new_n23025_ & new_n23028_;
  assign new_n23030_ = new_n23020_ & new_n23029_;
  assign new_n23031_ = new_n23009_ & new_n23030_;
  assign new_n23032_ = new_n22986_ & new_n23031_;
  assign new_n23033_ = new_n17987_ & new_n21116_;
  assign new_n23034_ = new_n17987_ & new_n21102_;
  assign new_n23035_ = new_n17987_ & new_n21114_;
  assign new_n23036_ = ~new_n23034_ & ~new_n23035_;
  assign new_n23037_ = ~new_n23033_ & new_n23036_;
  assign new_n23038_ = new_n18033_ & new_n21019_;
  assign new_n23039_ = new_n17987_ & new_n21112_;
  assign new_n23040_ = new_n18033_ & new_n21017_;
  assign new_n23041_ = ~new_n23039_ & ~new_n23040_;
  assign new_n23042_ = ~new_n23038_ & new_n23041_;
  assign new_n23043_ = new_n23037_ & new_n23042_;
  assign new_n23044_ = new_n18033_ & new_n21029_;
  assign new_n23045_ = new_n18033_ & new_n21015_;
  assign new_n23046_ = new_n18033_ & new_n21026_;
  assign new_n23047_ = ~new_n23045_ & ~new_n23046_;
  assign new_n23048_ = ~new_n23044_ & new_n23047_;
  assign new_n23049_ = new_n18033_ & new_n21042_;
  assign new_n23050_ = new_n18033_ & new_n21024_;
  assign new_n23051_ = new_n18033_ & new_n21039_;
  assign new_n23052_ = ~new_n23050_ & ~new_n23051_;
  assign new_n23053_ = ~new_n23049_ & new_n23052_;
  assign new_n23054_ = new_n23048_ & new_n23053_;
  assign new_n23055_ = new_n23043_ & new_n23054_;
  assign new_n23056_ = new_n18033_ & new_n21053_;
  assign new_n23057_ = new_n18033_ & new_n21036_;
  assign new_n23058_ = new_n18033_ & new_n21050_;
  assign new_n23059_ = ~new_n23057_ & ~new_n23058_;
  assign new_n23060_ = ~new_n23056_ & new_n23059_;
  assign new_n23061_ = new_n18033_ & new_n21062_;
  assign new_n23062_ = new_n18033_ & new_n21047_;
  assign new_n23063_ = new_n18033_ & new_n21060_;
  assign new_n23064_ = ~new_n23062_ & ~new_n23063_;
  assign new_n23065_ = ~new_n23061_ & new_n23064_;
  assign new_n23066_ = new_n23060_ & new_n23065_;
  assign new_n23067_ = new_n18033_ & new_n21068_;
  assign new_n23068_ = new_n18033_ & new_n21058_;
  assign new_n23069_ = new_n18033_ & new_n21066_;
  assign new_n23070_ = ~new_n23068_ & ~new_n23069_;
  assign new_n23071_ = ~new_n23067_ & new_n23070_;
  assign new_n23072_ = new_n18033_ & new_n21079_;
  assign new_n23073_ = new_n18033_ & new_n21081_;
  assign new_n23074_ = ~new_n23072_ & ~new_n23073_;
  assign new_n23075_ = new_n23071_ & new_n23074_;
  assign new_n23076_ = new_n23066_ & new_n23075_;
  assign new_n23077_ = new_n23055_ & new_n23076_;
  assign new_n23078_ = new_n18033_ & new_n21089_;
  assign new_n23079_ = new_n18033_ & new_n21077_;
  assign new_n23080_ = new_n18033_ & new_n21087_;
  assign new_n23081_ = ~new_n23079_ & ~new_n23080_;
  assign new_n23082_ = ~new_n23078_ & new_n23081_;
  assign new_n23083_ = new_n18033_ & new_n21098_;
  assign new_n23084_ = new_n18033_ & new_n21085_;
  assign new_n23085_ = new_n18033_ & new_n21096_;
  assign new_n23086_ = ~new_n23084_ & ~new_n23085_;
  assign new_n23087_ = ~new_n23083_ & new_n23086_;
  assign new_n23088_ = new_n23082_ & new_n23087_;
  assign new_n23089_ = new_n18033_ & new_n21106_;
  assign new_n23090_ = new_n18033_ & new_n21094_;
  assign new_n23091_ = new_n18033_ & new_n21104_;
  assign new_n23092_ = ~new_n23090_ & ~new_n23091_;
  assign new_n23093_ = ~new_n23089_ & new_n23092_;
  assign new_n23094_ = new_n18033_ & new_n21116_;
  assign new_n23095_ = new_n18033_ & new_n21102_;
  assign new_n23096_ = new_n18033_ & new_n21114_;
  assign new_n23097_ = ~new_n23095_ & ~new_n23096_;
  assign new_n23098_ = ~new_n23094_ & new_n23097_;
  assign new_n23099_ = new_n23093_ & new_n23098_;
  assign new_n23100_ = new_n23088_ & new_n23099_;
  assign new_n23101_ = new_n18405_ & new_n21019_;
  assign new_n23102_ = new_n18033_ & new_n21112_;
  assign new_n23103_ = new_n18405_ & new_n21017_;
  assign new_n23104_ = ~new_n23102_ & ~new_n23103_;
  assign new_n23105_ = ~new_n23101_ & new_n23104_;
  assign new_n23106_ = new_n18405_ & new_n21029_;
  assign new_n23107_ = new_n18405_ & new_n21015_;
  assign new_n23108_ = new_n18405_ & new_n21026_;
  assign new_n23109_ = ~new_n23107_ & ~new_n23108_;
  assign new_n23110_ = ~new_n23106_ & new_n23109_;
  assign new_n23111_ = new_n23105_ & new_n23110_;
  assign new_n23112_ = new_n18405_ & new_n21042_;
  assign new_n23113_ = new_n18405_ & new_n21024_;
  assign new_n23114_ = new_n18405_ & new_n21039_;
  assign new_n23115_ = ~new_n23113_ & ~new_n23114_;
  assign new_n23116_ = ~new_n23112_ & new_n23115_;
  assign new_n23117_ = new_n18405_ & new_n21036_;
  assign new_n23118_ = new_n18405_ & new_n21050_;
  assign new_n23119_ = ~new_n23117_ & ~new_n23118_;
  assign new_n23120_ = new_n23116_ & new_n23119_;
  assign new_n23121_ = new_n23111_ & new_n23120_;
  assign new_n23122_ = new_n23100_ & new_n23121_;
  assign new_n23123_ = new_n23077_ & new_n23122_;
  assign new_n23124_ = new_n23032_ & new_n23123_;
  assign new_n23125_ = new_n18405_ & new_n21060_;
  assign new_n23126_ = new_n18405_ & new_n21053_;
  assign new_n23127_ = new_n18405_ & new_n21047_;
  assign new_n23128_ = ~new_n23126_ & ~new_n23127_;
  assign new_n23129_ = ~new_n23125_ & new_n23128_;
  assign new_n23130_ = new_n18405_ & new_n21066_;
  assign new_n23131_ = new_n18405_ & new_n21062_;
  assign new_n23132_ = new_n18405_ & new_n21058_;
  assign new_n23133_ = ~new_n23131_ & ~new_n23132_;
  assign new_n23134_ = ~new_n23130_ & new_n23133_;
  assign new_n23135_ = new_n23129_ & new_n23134_;
  assign new_n23136_ = new_n18405_ & new_n21081_;
  assign new_n23137_ = new_n18405_ & new_n21068_;
  assign new_n23138_ = new_n18405_ & new_n21079_;
  assign new_n23139_ = ~new_n23137_ & ~new_n23138_;
  assign new_n23140_ = ~new_n23136_ & new_n23139_;
  assign new_n23141_ = new_n18405_ & new_n21089_;
  assign new_n23142_ = new_n18405_ & new_n21077_;
  assign new_n23143_ = new_n18405_ & new_n21087_;
  assign new_n23144_ = ~new_n23142_ & ~new_n23143_;
  assign new_n23145_ = ~new_n23141_ & new_n23144_;
  assign new_n23146_ = new_n23140_ & new_n23145_;
  assign new_n23147_ = new_n23135_ & new_n23146_;
  assign new_n23148_ = new_n18405_ & new_n21098_;
  assign new_n23149_ = new_n18405_ & new_n21085_;
  assign new_n23150_ = new_n18405_ & new_n21096_;
  assign new_n23151_ = ~new_n23149_ & ~new_n23150_;
  assign new_n23152_ = ~new_n23148_ & new_n23151_;
  assign new_n23153_ = new_n18405_ & new_n21106_;
  assign new_n23154_ = new_n18405_ & new_n21094_;
  assign new_n23155_ = new_n18405_ & new_n21104_;
  assign new_n23156_ = ~new_n23154_ & ~new_n23155_;
  assign new_n23157_ = ~new_n23153_ & new_n23156_;
  assign new_n23158_ = new_n23152_ & new_n23157_;
  assign new_n23159_ = new_n18405_ & new_n21116_;
  assign new_n23160_ = new_n18405_ & new_n21102_;
  assign new_n23161_ = new_n18405_ & new_n21114_;
  assign new_n23162_ = ~new_n23160_ & ~new_n23161_;
  assign new_n23163_ = ~new_n23159_ & new_n23162_;
  assign new_n23164_ = new_n18405_ & new_n21112_;
  assign new_n23165_ = new_n18455_ & new_n21017_;
  assign new_n23166_ = ~new_n23164_ & ~new_n23165_;
  assign new_n23167_ = new_n23163_ & new_n23166_;
  assign new_n23168_ = new_n23158_ & new_n23167_;
  assign new_n23169_ = new_n23147_ & new_n23168_;
  assign new_n23170_ = new_n18455_ & new_n21026_;
  assign new_n23171_ = new_n18455_ & new_n21019_;
  assign new_n23172_ = new_n18455_ & new_n21015_;
  assign new_n23173_ = ~new_n23171_ & ~new_n23172_;
  assign new_n23174_ = ~new_n23170_ & new_n23173_;
  assign new_n23175_ = new_n18455_ & new_n21039_;
  assign new_n23176_ = new_n18455_ & new_n21029_;
  assign new_n23177_ = new_n18455_ & new_n21024_;
  assign new_n23178_ = ~new_n23176_ & ~new_n23177_;
  assign new_n23179_ = ~new_n23175_ & new_n23178_;
  assign new_n23180_ = new_n23174_ & new_n23179_;
  assign new_n23181_ = new_n18455_ & new_n21050_;
  assign new_n23182_ = new_n18455_ & new_n21042_;
  assign new_n23183_ = new_n18455_ & new_n21036_;
  assign new_n23184_ = ~new_n23182_ & ~new_n23183_;
  assign new_n23185_ = ~new_n23181_ & new_n23184_;
  assign new_n23186_ = new_n18455_ & new_n21060_;
  assign new_n23187_ = new_n18455_ & new_n21053_;
  assign new_n23188_ = new_n18455_ & new_n21047_;
  assign new_n23189_ = ~new_n23187_ & ~new_n23188_;
  assign new_n23190_ = ~new_n23186_ & new_n23189_;
  assign new_n23191_ = new_n23185_ & new_n23190_;
  assign new_n23192_ = new_n23180_ & new_n23191_;
  assign new_n23193_ = new_n18455_ & new_n21066_;
  assign new_n23194_ = new_n18455_ & new_n21062_;
  assign new_n23195_ = new_n18455_ & new_n21058_;
  assign new_n23196_ = ~new_n23194_ & ~new_n23195_;
  assign new_n23197_ = ~new_n23193_ & new_n23196_;
  assign new_n23198_ = new_n18455_ & new_n21081_;
  assign new_n23199_ = new_n18455_ & new_n21068_;
  assign new_n23200_ = new_n18455_ & new_n21079_;
  assign new_n23201_ = ~new_n23199_ & ~new_n23200_;
  assign new_n23202_ = ~new_n23198_ & new_n23201_;
  assign new_n23203_ = new_n23197_ & new_n23202_;
  assign new_n23204_ = new_n18455_ & new_n21089_;
  assign new_n23205_ = new_n18455_ & new_n21077_;
  assign new_n23206_ = new_n18455_ & new_n21087_;
  assign new_n23207_ = ~new_n23205_ & ~new_n23206_;
  assign new_n23208_ = ~new_n23204_ & new_n23207_;
  assign new_n23209_ = new_n18455_ & new_n21085_;
  assign new_n23210_ = new_n18455_ & new_n21096_;
  assign new_n23211_ = ~new_n23209_ & ~new_n23210_;
  assign new_n23212_ = new_n23208_ & new_n23211_;
  assign new_n23213_ = new_n23203_ & new_n23212_;
  assign new_n23214_ = new_n23192_ & new_n23213_;
  assign new_n23215_ = new_n23169_ & new_n23214_;
  assign new_n23216_ = new_n18455_ & new_n21104_;
  assign new_n23217_ = new_n18455_ & new_n21098_;
  assign new_n23218_ = new_n18455_ & new_n21094_;
  assign new_n23219_ = ~new_n23217_ & ~new_n23218_;
  assign new_n23220_ = ~new_n23216_ & new_n23219_;
  assign new_n23221_ = new_n18455_ & new_n21114_;
  assign new_n23222_ = new_n18455_ & new_n21106_;
  assign new_n23223_ = new_n18455_ & new_n21102_;
  assign new_n23224_ = ~new_n23222_ & ~new_n23223_;
  assign new_n23225_ = ~new_n23221_ & new_n23224_;
  assign new_n23226_ = new_n23220_ & new_n23225_;
  assign new_n23227_ = new_n18503_ & new_n21017_;
  assign new_n23228_ = new_n18455_ & new_n21116_;
  assign new_n23229_ = new_n18455_ & new_n21112_;
  assign new_n23230_ = ~new_n23228_ & ~new_n23229_;
  assign new_n23231_ = ~new_n23227_ & new_n23230_;
  assign new_n23232_ = new_n18503_ & new_n21026_;
  assign new_n23233_ = new_n18503_ & new_n21019_;
  assign new_n23234_ = new_n18503_ & new_n21015_;
  assign new_n23235_ = ~new_n23233_ & ~new_n23234_;
  assign new_n23236_ = ~new_n23232_ & new_n23235_;
  assign new_n23237_ = new_n23231_ & new_n23236_;
  assign new_n23238_ = new_n23226_ & new_n23237_;
  assign new_n23239_ = new_n18503_ & new_n21039_;
  assign new_n23240_ = new_n18503_ & new_n21029_;
  assign new_n23241_ = new_n18503_ & new_n21024_;
  assign new_n23242_ = ~new_n23240_ & ~new_n23241_;
  assign new_n23243_ = ~new_n23239_ & new_n23242_;
  assign new_n23244_ = new_n18503_ & new_n21050_;
  assign new_n23245_ = new_n18503_ & new_n21042_;
  assign new_n23246_ = new_n18503_ & new_n21036_;
  assign new_n23247_ = ~new_n23245_ & ~new_n23246_;
  assign new_n23248_ = ~new_n23244_ & new_n23247_;
  assign new_n23249_ = new_n23243_ & new_n23248_;
  assign new_n23250_ = new_n18503_ & new_n21060_;
  assign new_n23251_ = new_n18503_ & new_n21053_;
  assign new_n23252_ = new_n18503_ & new_n21047_;
  assign new_n23253_ = ~new_n23251_ & ~new_n23252_;
  assign new_n23254_ = ~new_n23250_ & new_n23253_;
  assign new_n23255_ = new_n18503_ & new_n21062_;
  assign new_n23256_ = new_n18503_ & new_n21058_;
  assign new_n23257_ = ~new_n23255_ & ~new_n23256_;
  assign new_n23258_ = new_n23254_ & new_n23257_;
  assign new_n23259_ = new_n23249_ & new_n23258_;
  assign new_n23260_ = new_n23238_ & new_n23259_;
  assign new_n23261_ = new_n18503_ & new_n21079_;
  assign new_n23262_ = new_n18503_ & new_n21066_;
  assign new_n23263_ = new_n18503_ & new_n21068_;
  assign new_n23264_ = ~new_n23262_ & ~new_n23263_;
  assign new_n23265_ = ~new_n23261_ & new_n23264_;
  assign new_n23266_ = new_n18503_ & new_n21087_;
  assign new_n23267_ = new_n18503_ & new_n21081_;
  assign new_n23268_ = new_n18503_ & new_n21077_;
  assign new_n23269_ = ~new_n23267_ & ~new_n23268_;
  assign new_n23270_ = ~new_n23266_ & new_n23269_;
  assign new_n23271_ = new_n23265_ & new_n23270_;
  assign new_n23272_ = new_n18503_ & new_n21096_;
  assign new_n23273_ = new_n18503_ & new_n21089_;
  assign new_n23274_ = new_n18503_ & new_n21085_;
  assign new_n23275_ = ~new_n23273_ & ~new_n23274_;
  assign new_n23276_ = ~new_n23272_ & new_n23275_;
  assign new_n23277_ = new_n18503_ & new_n21104_;
  assign new_n23278_ = new_n18503_ & new_n21098_;
  assign new_n23279_ = new_n18503_ & new_n21094_;
  assign new_n23280_ = ~new_n23278_ & ~new_n23279_;
  assign new_n23281_ = ~new_n23277_ & new_n23280_;
  assign new_n23282_ = new_n23276_ & new_n23281_;
  assign new_n23283_ = new_n23271_ & new_n23282_;
  assign new_n23284_ = new_n18503_ & new_n21114_;
  assign new_n23285_ = new_n18503_ & new_n21106_;
  assign new_n23286_ = new_n18503_ & new_n21102_;
  assign new_n23287_ = ~new_n23285_ & ~new_n23286_;
  assign new_n23288_ = ~new_n23284_ & new_n23287_;
  assign new_n23289_ = new_n18555_ & new_n21017_;
  assign new_n23290_ = new_n18503_ & new_n21116_;
  assign new_n23291_ = new_n18503_ & new_n21112_;
  assign new_n23292_ = ~new_n23290_ & ~new_n23291_;
  assign new_n23293_ = ~new_n23289_ & new_n23292_;
  assign new_n23294_ = new_n23288_ & new_n23293_;
  assign new_n23295_ = new_n18555_ & new_n21026_;
  assign new_n23296_ = new_n18555_ & new_n21019_;
  assign new_n23297_ = new_n18555_ & new_n21015_;
  assign new_n23298_ = ~new_n23296_ & ~new_n23297_;
  assign new_n23299_ = ~new_n23295_ & new_n23298_;
  assign new_n23300_ = new_n18555_ & new_n21029_;
  assign new_n23301_ = new_n18555_ & new_n21024_;
  assign new_n23302_ = ~new_n23300_ & ~new_n23301_;
  assign new_n23303_ = new_n23299_ & new_n23302_;
  assign new_n23304_ = new_n23294_ & new_n23303_;
  assign new_n23305_ = new_n23283_ & new_n23304_;
  assign new_n23306_ = new_n23260_ & new_n23305_;
  assign new_n23307_ = new_n23215_ & new_n23306_;
  assign new_n23308_ = new_n23124_ & new_n23307_;
  assign new_n23309_ = new_n18555_ & new_n21036_;
  assign new_n23310_ = new_n18555_ & new_n21039_;
  assign new_n23311_ = new_n18555_ & new_n21042_;
  assign new_n23312_ = ~new_n23310_ & ~new_n23311_;
  assign new_n23313_ = ~new_n23309_ & new_n23312_;
  assign new_n23314_ = new_n18555_ & new_n21047_;
  assign new_n23315_ = new_n18555_ & new_n21050_;
  assign new_n23316_ = new_n18555_ & new_n21053_;
  assign new_n23317_ = ~new_n23315_ & ~new_n23316_;
  assign new_n23318_ = ~new_n23314_ & new_n23317_;
  assign new_n23319_ = new_n23313_ & new_n23318_;
  assign new_n23320_ = new_n18555_ & new_n21058_;
  assign new_n23321_ = new_n18555_ & new_n21060_;
  assign new_n23322_ = new_n18555_ & new_n21062_;
  assign new_n23323_ = ~new_n23321_ & ~new_n23322_;
  assign new_n23324_ = ~new_n23320_ & new_n23323_;
  assign new_n23325_ = new_n18555_ & new_n21079_;
  assign new_n23326_ = new_n18555_ & new_n21066_;
  assign new_n23327_ = new_n18555_ & new_n21068_;
  assign new_n23328_ = ~new_n23326_ & ~new_n23327_;
  assign new_n23329_ = ~new_n23325_ & new_n23328_;
  assign new_n23330_ = new_n23324_ & new_n23329_;
  assign new_n23331_ = new_n23319_ & new_n23330_;
  assign new_n23332_ = new_n18555_ & new_n21087_;
  assign new_n23333_ = new_n18555_ & new_n21081_;
  assign new_n23334_ = new_n18555_ & new_n21077_;
  assign new_n23335_ = ~new_n23333_ & ~new_n23334_;
  assign new_n23336_ = ~new_n23332_ & new_n23335_;
  assign new_n23337_ = new_n18555_ & new_n21096_;
  assign new_n23338_ = new_n18555_ & new_n21089_;
  assign new_n23339_ = new_n18555_ & new_n21085_;
  assign new_n23340_ = ~new_n23338_ & ~new_n23339_;
  assign new_n23341_ = ~new_n23337_ & new_n23340_;
  assign new_n23342_ = new_n23336_ & new_n23341_;
  assign new_n23343_ = new_n18555_ & new_n21104_;
  assign new_n23344_ = new_n18555_ & new_n21098_;
  assign new_n23345_ = new_n18555_ & new_n21094_;
  assign new_n23346_ = ~new_n23344_ & ~new_n23345_;
  assign new_n23347_ = ~new_n23343_ & new_n23346_;
  assign new_n23348_ = new_n18555_ & new_n21106_;
  assign new_n23349_ = new_n18555_ & new_n21102_;
  assign new_n23350_ = ~new_n23348_ & ~new_n23349_;
  assign new_n23351_ = new_n23347_ & new_n23350_;
  assign new_n23352_ = new_n23342_ & new_n23351_;
  assign new_n23353_ = new_n23331_ & new_n23352_;
  assign new_n23354_ = new_n18555_ & new_n21112_;
  assign new_n23355_ = new_n18555_ & new_n21114_;
  assign new_n23356_ = new_n18555_ & new_n21116_;
  assign new_n23357_ = ~new_n23355_ & ~new_n23356_;
  assign new_n23358_ = ~new_n23354_ & new_n23357_;
  assign new_n23359_ = new_n18666_ & new_n21015_;
  assign new_n23360_ = new_n18666_ & new_n21017_;
  assign new_n23361_ = new_n18666_ & new_n21019_;
  assign new_n23362_ = ~new_n23360_ & ~new_n23361_;
  assign new_n23363_ = ~new_n23359_ & new_n23362_;
  assign new_n23364_ = new_n23358_ & new_n23363_;
  assign new_n23365_ = new_n18666_ & new_n21024_;
  assign new_n23366_ = new_n18666_ & new_n21026_;
  assign new_n23367_ = new_n18666_ & new_n21029_;
  assign new_n23368_ = ~new_n23366_ & ~new_n23367_;
  assign new_n23369_ = ~new_n23365_ & new_n23368_;
  assign new_n23370_ = new_n18666_ & new_n21036_;
  assign new_n23371_ = new_n18666_ & new_n21039_;
  assign new_n23372_ = new_n18666_ & new_n21042_;
  assign new_n23373_ = ~new_n23371_ & ~new_n23372_;
  assign new_n23374_ = ~new_n23370_ & new_n23373_;
  assign new_n23375_ = new_n23369_ & new_n23374_;
  assign new_n23376_ = new_n23364_ & new_n23375_;
  assign new_n23377_ = new_n18666_ & new_n21047_;
  assign new_n23378_ = new_n18666_ & new_n21050_;
  assign new_n23379_ = new_n18666_ & new_n21053_;
  assign new_n23380_ = ~new_n23378_ & ~new_n23379_;
  assign new_n23381_ = ~new_n23377_ & new_n23380_;
  assign new_n23382_ = new_n18666_ & new_n21058_;
  assign new_n23383_ = new_n18666_ & new_n21060_;
  assign new_n23384_ = new_n18666_ & new_n21062_;
  assign new_n23385_ = ~new_n23383_ & ~new_n23384_;
  assign new_n23386_ = ~new_n23382_ & new_n23385_;
  assign new_n23387_ = new_n23381_ & new_n23386_;
  assign new_n23388_ = new_n18666_ & new_n21079_;
  assign new_n23389_ = new_n18666_ & new_n21066_;
  assign new_n23390_ = new_n18666_ & new_n21068_;
  assign new_n23391_ = ~new_n23389_ & ~new_n23390_;
  assign new_n23392_ = ~new_n23388_ & new_n23391_;
  assign new_n23393_ = new_n18666_ & new_n21081_;
  assign new_n23394_ = new_n18666_ & new_n21077_;
  assign new_n23395_ = ~new_n23393_ & ~new_n23394_;
  assign new_n23396_ = new_n23392_ & new_n23395_;
  assign new_n23397_ = new_n23387_ & new_n23396_;
  assign new_n23398_ = new_n23376_ & new_n23397_;
  assign new_n23399_ = new_n23353_ & new_n23398_;
  assign new_n23400_ = new_n18666_ & new_n21085_;
  assign new_n23401_ = new_n18666_ & new_n21087_;
  assign new_n23402_ = new_n18666_ & new_n21089_;
  assign new_n23403_ = ~new_n23401_ & ~new_n23402_;
  assign new_n23404_ = ~new_n23400_ & new_n23403_;
  assign new_n23405_ = new_n18666_ & new_n21094_;
  assign new_n23406_ = new_n18666_ & new_n21096_;
  assign new_n23407_ = new_n18666_ & new_n21098_;
  assign new_n23408_ = ~new_n23406_ & ~new_n23407_;
  assign new_n23409_ = ~new_n23405_ & new_n23408_;
  assign new_n23410_ = new_n23404_ & new_n23409_;
  assign new_n23411_ = new_n18666_ & new_n21102_;
  assign new_n23412_ = new_n18666_ & new_n21104_;
  assign new_n23413_ = new_n18666_ & new_n21106_;
  assign new_n23414_ = ~new_n23412_ & ~new_n23413_;
  assign new_n23415_ = ~new_n23411_ & new_n23414_;
  assign new_n23416_ = new_n18666_ & new_n21112_;
  assign new_n23417_ = new_n18666_ & new_n21114_;
  assign new_n23418_ = new_n18666_ & new_n21116_;
  assign new_n23419_ = ~new_n23417_ & ~new_n23418_;
  assign new_n23420_ = ~new_n23416_ & new_n23419_;
  assign new_n23421_ = new_n23415_ & new_n23420_;
  assign new_n23422_ = new_n23410_ & new_n23421_;
  assign new_n23423_ = new_n18718_ & new_n21015_;
  assign new_n23424_ = new_n18718_ & new_n21017_;
  assign new_n23425_ = new_n18718_ & new_n21019_;
  assign new_n23426_ = ~new_n23424_ & ~new_n23425_;
  assign new_n23427_ = ~new_n23423_ & new_n23426_;
  assign new_n23428_ = new_n18718_ & new_n21024_;
  assign new_n23429_ = new_n18718_ & new_n21026_;
  assign new_n23430_ = new_n18718_ & new_n21029_;
  assign new_n23431_ = ~new_n23429_ & ~new_n23430_;
  assign new_n23432_ = ~new_n23428_ & new_n23431_;
  assign new_n23433_ = new_n23427_ & new_n23432_;
  assign new_n23434_ = new_n18718_ & new_n21036_;
  assign new_n23435_ = new_n18718_ & new_n21039_;
  assign new_n23436_ = new_n18718_ & new_n21042_;
  assign new_n23437_ = ~new_n23435_ & ~new_n23436_;
  assign new_n23438_ = ~new_n23434_ & new_n23437_;
  assign new_n23439_ = new_n18718_ & new_n21050_;
  assign new_n23440_ = new_n18718_ & new_n21053_;
  assign new_n23441_ = ~new_n23439_ & ~new_n23440_;
  assign new_n23442_ = new_n23438_ & new_n23441_;
  assign new_n23443_ = new_n23433_ & new_n23442_;
  assign new_n23444_ = new_n23422_ & new_n23443_;
  assign new_n23445_ = new_n18718_ & new_n21062_;
  assign new_n23446_ = new_n18718_ & new_n21047_;
  assign new_n23447_ = new_n18718_ & new_n21060_;
  assign new_n23448_ = ~new_n23446_ & ~new_n23447_;
  assign new_n23449_ = ~new_n23445_ & new_n23448_;
  assign new_n23450_ = new_n18718_ & new_n21068_;
  assign new_n23451_ = new_n18718_ & new_n21058_;
  assign new_n23452_ = new_n18718_ & new_n21066_;
  assign new_n23453_ = ~new_n23451_ & ~new_n23452_;
  assign new_n23454_ = ~new_n23450_ & new_n23453_;
  assign new_n23455_ = new_n23449_ & new_n23454_;
  assign new_n23456_ = new_n18718_ & new_n21077_;
  assign new_n23457_ = new_n18718_ & new_n21079_;
  assign new_n23458_ = new_n18718_ & new_n21081_;
  assign new_n23459_ = ~new_n23457_ & ~new_n23458_;
  assign new_n23460_ = ~new_n23456_ & new_n23459_;
  assign new_n23461_ = new_n18718_ & new_n21085_;
  assign new_n23462_ = new_n18718_ & new_n21087_;
  assign new_n23463_ = new_n18718_ & new_n21089_;
  assign new_n23464_ = ~new_n23462_ & ~new_n23463_;
  assign new_n23465_ = ~new_n23461_ & new_n23464_;
  assign new_n23466_ = new_n23460_ & new_n23465_;
  assign new_n23467_ = new_n23455_ & new_n23466_;
  assign new_n23468_ = new_n18718_ & new_n21094_;
  assign new_n23469_ = new_n18718_ & new_n21096_;
  assign new_n23470_ = new_n18718_ & new_n21098_;
  assign new_n23471_ = ~new_n23469_ & ~new_n23470_;
  assign new_n23472_ = ~new_n23468_ & new_n23471_;
  assign new_n23473_ = new_n18718_ & new_n21102_;
  assign new_n23474_ = new_n18718_ & new_n21104_;
  assign new_n23475_ = new_n18718_ & new_n21106_;
  assign new_n23476_ = ~new_n23474_ & ~new_n23475_;
  assign new_n23477_ = ~new_n23473_ & new_n23476_;
  assign new_n23478_ = new_n23472_ & new_n23477_;
  assign new_n23479_ = new_n18718_ & new_n21112_;
  assign new_n23480_ = new_n18718_ & new_n21114_;
  assign new_n23481_ = new_n18718_ & new_n21116_;
  assign new_n23482_ = ~new_n23480_ & ~new_n23481_;
  assign new_n23483_ = ~new_n23479_ & new_n23482_;
  assign new_n23484_ = new_n18764_ & new_n21017_;
  assign new_n23485_ = new_n18764_ & new_n21019_;
  assign new_n23486_ = ~new_n23484_ & ~new_n23485_;
  assign new_n23487_ = new_n23483_ & new_n23486_;
  assign new_n23488_ = new_n23478_ & new_n23487_;
  assign new_n23489_ = new_n23467_ & new_n23488_;
  assign new_n23490_ = new_n23444_ & new_n23489_;
  assign new_n23491_ = new_n23399_ & new_n23490_;
  assign new_n23492_ = new_n18764_ & new_n21029_;
  assign new_n23493_ = new_n18764_ & new_n21015_;
  assign new_n23494_ = new_n18764_ & new_n21026_;
  assign new_n23495_ = ~new_n23493_ & ~new_n23494_;
  assign new_n23496_ = ~new_n23492_ & new_n23495_;
  assign new_n23497_ = new_n18764_ & new_n21042_;
  assign new_n23498_ = new_n18764_ & new_n21024_;
  assign new_n23499_ = new_n18764_ & new_n21039_;
  assign new_n23500_ = ~new_n23498_ & ~new_n23499_;
  assign new_n23501_ = ~new_n23497_ & new_n23500_;
  assign new_n23502_ = new_n23496_ & new_n23501_;
  assign new_n23503_ = new_n18764_ & new_n21053_;
  assign new_n23504_ = new_n18764_ & new_n21036_;
  assign new_n23505_ = new_n18764_ & new_n21050_;
  assign new_n23506_ = ~new_n23504_ & ~new_n23505_;
  assign new_n23507_ = ~new_n23503_ & new_n23506_;
  assign new_n23508_ = new_n18764_ & new_n21062_;
  assign new_n23509_ = new_n18764_ & new_n21047_;
  assign new_n23510_ = new_n18764_ & new_n21060_;
  assign new_n23511_ = ~new_n23509_ & ~new_n23510_;
  assign new_n23512_ = ~new_n23508_ & new_n23511_;
  assign new_n23513_ = new_n23507_ & new_n23512_;
  assign new_n23514_ = new_n23502_ & new_n23513_;
  assign new_n23515_ = new_n18764_ & new_n21068_;
  assign new_n23516_ = new_n18764_ & new_n21058_;
  assign new_n23517_ = new_n18764_ & new_n21066_;
  assign new_n23518_ = ~new_n23516_ & ~new_n23517_;
  assign new_n23519_ = ~new_n23515_ & new_n23518_;
  assign new_n23520_ = new_n18764_ & new_n21077_;
  assign new_n23521_ = new_n18764_ & new_n21079_;
  assign new_n23522_ = new_n18764_ & new_n21081_;
  assign new_n23523_ = ~new_n23521_ & ~new_n23522_;
  assign new_n23524_ = ~new_n23520_ & new_n23523_;
  assign new_n23525_ = new_n23519_ & new_n23524_;
  assign new_n23526_ = new_n18764_ & new_n21085_;
  assign new_n23527_ = new_n18764_ & new_n21087_;
  assign new_n23528_ = new_n18764_ & new_n21089_;
  assign new_n23529_ = ~new_n23527_ & ~new_n23528_;
  assign new_n23530_ = ~new_n23526_ & new_n23529_;
  assign new_n23531_ = new_n18764_ & new_n21096_;
  assign new_n23532_ = new_n18764_ & new_n21098_;
  assign new_n23533_ = ~new_n23531_ & ~new_n23532_;
  assign new_n23534_ = new_n23530_ & new_n23533_;
  assign new_n23535_ = new_n23525_ & new_n23534_;
  assign new_n23536_ = new_n23514_ & new_n23535_;
  assign new_n23537_ = new_n18764_ & new_n21106_;
  assign new_n23538_ = new_n18764_ & new_n21094_;
  assign new_n23539_ = new_n18764_ & new_n21104_;
  assign new_n23540_ = ~new_n23538_ & ~new_n23539_;
  assign new_n23541_ = ~new_n23537_ & new_n23540_;
  assign new_n23542_ = new_n18764_ & new_n21116_;
  assign new_n23543_ = new_n18764_ & new_n21102_;
  assign new_n23544_ = new_n18764_ & new_n21114_;
  assign new_n23545_ = ~new_n23543_ & ~new_n23544_;
  assign new_n23546_ = ~new_n23542_ & new_n23545_;
  assign new_n23547_ = new_n23541_ & new_n23546_;
  assign new_n23548_ = new_n18813_ & new_n21019_;
  assign new_n23549_ = new_n18764_ & new_n21112_;
  assign new_n23550_ = new_n18813_ & new_n21017_;
  assign new_n23551_ = ~new_n23549_ & ~new_n23550_;
  assign new_n23552_ = ~new_n23548_ & new_n23551_;
  assign new_n23553_ = new_n18813_ & new_n21029_;
  assign new_n23554_ = new_n18813_ & new_n21015_;
  assign new_n23555_ = new_n18813_ & new_n21026_;
  assign new_n23556_ = ~new_n23554_ & ~new_n23555_;
  assign new_n23557_ = ~new_n23553_ & new_n23556_;
  assign new_n23558_ = new_n23552_ & new_n23557_;
  assign new_n23559_ = new_n23547_ & new_n23558_;
  assign new_n23560_ = new_n18813_ & new_n21042_;
  assign new_n23561_ = new_n18813_ & new_n21024_;
  assign new_n23562_ = new_n18813_ & new_n21039_;
  assign new_n23563_ = ~new_n23561_ & ~new_n23562_;
  assign new_n23564_ = ~new_n23560_ & new_n23563_;
  assign new_n23565_ = new_n18813_ & new_n21053_;
  assign new_n23566_ = new_n18813_ & new_n21036_;
  assign new_n23567_ = new_n18813_ & new_n21050_;
  assign new_n23568_ = ~new_n23566_ & ~new_n23567_;
  assign new_n23569_ = ~new_n23565_ & new_n23568_;
  assign new_n23570_ = new_n23564_ & new_n23569_;
  assign new_n23571_ = new_n18813_ & new_n21062_;
  assign new_n23572_ = new_n18813_ & new_n21047_;
  assign new_n23573_ = new_n18813_ & new_n21060_;
  assign new_n23574_ = ~new_n23572_ & ~new_n23573_;
  assign new_n23575_ = ~new_n23571_ & new_n23574_;
  assign new_n23576_ = new_n18813_ & new_n21058_;
  assign new_n23577_ = new_n18813_ & new_n21066_;
  assign new_n23578_ = ~new_n23576_ & ~new_n23577_;
  assign new_n23579_ = new_n23575_ & new_n23578_;
  assign new_n23580_ = new_n23570_ & new_n23579_;
  assign new_n23581_ = new_n23559_ & new_n23580_;
  assign new_n23582_ = new_n23536_ & new_n23581_;
  assign new_n23583_ = new_n18813_ & new_n21081_;
  assign new_n23584_ = new_n18813_ & new_n21068_;
  assign new_n23585_ = new_n18813_ & new_n21079_;
  assign new_n23586_ = ~new_n23584_ & ~new_n23585_;
  assign new_n23587_ = ~new_n23583_ & new_n23586_;
  assign new_n23588_ = new_n18813_ & new_n21089_;
  assign new_n23589_ = new_n18813_ & new_n21077_;
  assign new_n23590_ = new_n18813_ & new_n21087_;
  assign new_n23591_ = ~new_n23589_ & ~new_n23590_;
  assign new_n23592_ = ~new_n23588_ & new_n23591_;
  assign new_n23593_ = new_n23587_ & new_n23592_;
  assign new_n23594_ = new_n18813_ & new_n21098_;
  assign new_n23595_ = new_n18813_ & new_n21085_;
  assign new_n23596_ = new_n18813_ & new_n21096_;
  assign new_n23597_ = ~new_n23595_ & ~new_n23596_;
  assign new_n23598_ = ~new_n23594_ & new_n23597_;
  assign new_n23599_ = new_n18813_ & new_n21106_;
  assign new_n23600_ = new_n18813_ & new_n21094_;
  assign new_n23601_ = new_n18813_ & new_n21104_;
  assign new_n23602_ = ~new_n23600_ & ~new_n23601_;
  assign new_n23603_ = ~new_n23599_ & new_n23602_;
  assign new_n23604_ = new_n23598_ & new_n23603_;
  assign new_n23605_ = new_n23593_ & new_n23604_;
  assign new_n23606_ = new_n18813_ & new_n21116_;
  assign new_n23607_ = new_n18813_ & new_n21102_;
  assign new_n23608_ = new_n18813_ & new_n21114_;
  assign new_n23609_ = ~new_n23607_ & ~new_n23608_;
  assign new_n23610_ = ~new_n23606_ & new_n23609_;
  assign new_n23611_ = new_n18929_ & new_n21019_;
  assign new_n23612_ = new_n18813_ & new_n21112_;
  assign new_n23613_ = new_n18929_ & new_n21017_;
  assign new_n23614_ = ~new_n23612_ & ~new_n23613_;
  assign new_n23615_ = ~new_n23611_ & new_n23614_;
  assign new_n23616_ = new_n23610_ & new_n23615_;
  assign new_n23617_ = new_n18929_ & new_n21029_;
  assign new_n23618_ = new_n18929_ & new_n21015_;
  assign new_n23619_ = new_n18929_ & new_n21026_;
  assign new_n23620_ = ~new_n23618_ & ~new_n23619_;
  assign new_n23621_ = ~new_n23617_ & new_n23620_;
  assign new_n23622_ = new_n18929_ & new_n21024_;
  assign new_n23623_ = new_n18929_ & new_n21039_;
  assign new_n23624_ = ~new_n23622_ & ~new_n23623_;
  assign new_n23625_ = new_n23621_ & new_n23624_;
  assign new_n23626_ = new_n23616_ & new_n23625_;
  assign new_n23627_ = new_n23605_ & new_n23626_;
  assign new_n23628_ = new_n18929_ & new_n21050_;
  assign new_n23629_ = new_n18929_ & new_n21042_;
  assign new_n23630_ = new_n18929_ & new_n21036_;
  assign new_n23631_ = ~new_n23629_ & ~new_n23630_;
  assign new_n23632_ = ~new_n23628_ & new_n23631_;
  assign new_n23633_ = new_n18929_ & new_n21060_;
  assign new_n23634_ = new_n18929_ & new_n21053_;
  assign new_n23635_ = new_n18929_ & new_n21047_;
  assign new_n23636_ = ~new_n23634_ & ~new_n23635_;
  assign new_n23637_ = ~new_n23633_ & new_n23636_;
  assign new_n23638_ = new_n23632_ & new_n23637_;
  assign new_n23639_ = new_n18929_ & new_n21066_;
  assign new_n23640_ = new_n18929_ & new_n21062_;
  assign new_n23641_ = new_n18929_ & new_n21058_;
  assign new_n23642_ = ~new_n23640_ & ~new_n23641_;
  assign new_n23643_ = ~new_n23639_ & new_n23642_;
  assign new_n23644_ = new_n18929_ & new_n21081_;
  assign new_n23645_ = new_n18929_ & new_n21068_;
  assign new_n23646_ = new_n18929_ & new_n21079_;
  assign new_n23647_ = ~new_n23645_ & ~new_n23646_;
  assign new_n23648_ = ~new_n23644_ & new_n23647_;
  assign new_n23649_ = new_n23643_ & new_n23648_;
  assign new_n23650_ = new_n23638_ & new_n23649_;
  assign new_n23651_ = new_n18929_ & new_n21089_;
  assign new_n23652_ = new_n18929_ & new_n21077_;
  assign new_n23653_ = new_n18929_ & new_n21087_;
  assign new_n23654_ = ~new_n23652_ & ~new_n23653_;
  assign new_n23655_ = ~new_n23651_ & new_n23654_;
  assign new_n23656_ = new_n18929_ & new_n21098_;
  assign new_n23657_ = new_n18929_ & new_n21085_;
  assign new_n23658_ = new_n18929_ & new_n21096_;
  assign new_n23659_ = ~new_n23657_ & ~new_n23658_;
  assign new_n23660_ = ~new_n23656_ & new_n23659_;
  assign new_n23661_ = new_n23655_ & new_n23660_;
  assign new_n23662_ = new_n18929_ & new_n21106_;
  assign new_n23663_ = new_n18929_ & new_n21094_;
  assign new_n23664_ = new_n18929_ & new_n21104_;
  assign new_n23665_ = ~new_n23663_ & ~new_n23664_;
  assign new_n23666_ = ~new_n23662_ & new_n23665_;
  assign new_n23667_ = new_n18929_ & new_n21102_;
  assign new_n23668_ = new_n18929_ & new_n21114_;
  assign new_n23669_ = ~new_n23667_ & ~new_n23668_;
  assign new_n23670_ = new_n23666_ & new_n23669_;
  assign new_n23671_ = new_n23661_ & new_n23670_;
  assign new_n23672_ = new_n23650_ & new_n23671_;
  assign new_n23673_ = new_n23627_ & new_n23672_;
  assign new_n23674_ = new_n23582_ & new_n23673_;
  assign new_n23675_ = new_n23491_ & new_n23674_;
  assign new_n23676_ = new_n23308_ & new_n23675_;
  assign new_n23677_ = new_n22939_ & new_n23676_;
  assign new_n23678_ = new_n18976_ & new_n21017_;
  assign new_n23679_ = new_n18929_ & new_n21116_;
  assign new_n23680_ = new_n18929_ & new_n21112_;
  assign new_n23681_ = ~new_n23679_ & ~new_n23680_;
  assign new_n23682_ = ~new_n23678_ & new_n23681_;
  assign new_n23683_ = new_n18976_ & new_n21026_;
  assign new_n23684_ = new_n18976_ & new_n21019_;
  assign new_n23685_ = new_n18976_ & new_n21015_;
  assign new_n23686_ = ~new_n23684_ & ~new_n23685_;
  assign new_n23687_ = ~new_n23683_ & new_n23686_;
  assign new_n23688_ = new_n23682_ & new_n23687_;
  assign new_n23689_ = new_n18976_ & new_n21039_;
  assign new_n23690_ = new_n18976_ & new_n21029_;
  assign new_n23691_ = new_n18976_ & new_n21024_;
  assign new_n23692_ = ~new_n23690_ & ~new_n23691_;
  assign new_n23693_ = ~new_n23689_ & new_n23692_;
  assign new_n23694_ = new_n18976_ & new_n21050_;
  assign new_n23695_ = new_n18976_ & new_n21042_;
  assign new_n23696_ = new_n18976_ & new_n21036_;
  assign new_n23697_ = ~new_n23695_ & ~new_n23696_;
  assign new_n23698_ = ~new_n23694_ & new_n23697_;
  assign new_n23699_ = new_n23693_ & new_n23698_;
  assign new_n23700_ = new_n23688_ & new_n23699_;
  assign new_n23701_ = new_n18976_ & new_n21060_;
  assign new_n23702_ = new_n18976_ & new_n21053_;
  assign new_n23703_ = new_n18976_ & new_n21047_;
  assign new_n23704_ = ~new_n23702_ & ~new_n23703_;
  assign new_n23705_ = ~new_n23701_ & new_n23704_;
  assign new_n23706_ = new_n18976_ & new_n21066_;
  assign new_n23707_ = new_n18976_ & new_n21062_;
  assign new_n23708_ = new_n18976_ & new_n21058_;
  assign new_n23709_ = ~new_n23707_ & ~new_n23708_;
  assign new_n23710_ = ~new_n23706_ & new_n23709_;
  assign new_n23711_ = new_n23705_ & new_n23710_;
  assign new_n23712_ = new_n18976_ & new_n21081_;
  assign new_n23713_ = new_n18976_ & new_n21068_;
  assign new_n23714_ = new_n18976_ & new_n21079_;
  assign new_n23715_ = ~new_n23713_ & ~new_n23714_;
  assign new_n23716_ = ~new_n23712_ & new_n23715_;
  assign new_n23717_ = new_n18976_ & new_n21089_;
  assign new_n23718_ = new_n18976_ & new_n21077_;
  assign new_n23719_ = new_n18976_ & new_n21087_;
  assign new_n23720_ = ~new_n23718_ & ~new_n23719_;
  assign new_n23721_ = ~new_n23717_ & new_n23720_;
  assign new_n23722_ = new_n23716_ & new_n23721_;
  assign new_n23723_ = new_n23711_ & new_n23722_;
  assign new_n23724_ = new_n23700_ & new_n23723_;
  assign new_n23725_ = new_n18976_ & new_n21098_;
  assign new_n23726_ = new_n18976_ & new_n21085_;
  assign new_n23727_ = new_n18976_ & new_n21096_;
  assign new_n23728_ = ~new_n23726_ & ~new_n23727_;
  assign new_n23729_ = ~new_n23725_ & new_n23728_;
  assign new_n23730_ = new_n18976_ & new_n21106_;
  assign new_n23731_ = new_n18976_ & new_n21094_;
  assign new_n23732_ = new_n18976_ & new_n21104_;
  assign new_n23733_ = ~new_n23731_ & ~new_n23732_;
  assign new_n23734_ = ~new_n23730_ & new_n23733_;
  assign new_n23735_ = new_n23729_ & new_n23734_;
  assign new_n23736_ = new_n18976_ & new_n21116_;
  assign new_n23737_ = new_n18976_ & new_n21102_;
  assign new_n23738_ = new_n18976_ & new_n21114_;
  assign new_n23739_ = ~new_n23737_ & ~new_n23738_;
  assign new_n23740_ = ~new_n23736_ & new_n23739_;
  assign new_n23741_ = new_n19029_ & new_n21019_;
  assign new_n23742_ = new_n18976_ & new_n21112_;
  assign new_n23743_ = new_n19029_ & new_n21017_;
  assign new_n23744_ = ~new_n23742_ & ~new_n23743_;
  assign new_n23745_ = ~new_n23741_ & new_n23744_;
  assign new_n23746_ = new_n23740_ & new_n23745_;
  assign new_n23747_ = new_n23735_ & new_n23746_;
  assign new_n23748_ = new_n19029_ & new_n21029_;
  assign new_n23749_ = new_n19029_ & new_n21015_;
  assign new_n23750_ = new_n19029_ & new_n21026_;
  assign new_n23751_ = ~new_n23749_ & ~new_n23750_;
  assign new_n23752_ = ~new_n23748_ & new_n23751_;
  assign new_n23753_ = new_n19029_ & new_n21042_;
  assign new_n23754_ = new_n19029_ & new_n21024_;
  assign new_n23755_ = new_n19029_ & new_n21039_;
  assign new_n23756_ = ~new_n23754_ & ~new_n23755_;
  assign new_n23757_ = ~new_n23753_ & new_n23756_;
  assign new_n23758_ = new_n23752_ & new_n23757_;
  assign new_n23759_ = new_n19029_ & new_n21053_;
  assign new_n23760_ = new_n19029_ & new_n21036_;
  assign new_n23761_ = new_n19029_ & new_n21050_;
  assign new_n23762_ = ~new_n23760_ & ~new_n23761_;
  assign new_n23763_ = ~new_n23759_ & new_n23762_;
  assign new_n23764_ = new_n19029_ & new_n21047_;
  assign new_n23765_ = new_n19029_ & new_n21060_;
  assign new_n23766_ = ~new_n23764_ & ~new_n23765_;
  assign new_n23767_ = new_n23763_ & new_n23766_;
  assign new_n23768_ = new_n23758_ & new_n23767_;
  assign new_n23769_ = new_n23747_ & new_n23768_;
  assign new_n23770_ = new_n23724_ & new_n23769_;
  assign new_n23771_ = new_n19029_ & new_n21066_;
  assign new_n23772_ = new_n19029_ & new_n21062_;
  assign new_n23773_ = new_n19029_ & new_n21058_;
  assign new_n23774_ = ~new_n23772_ & ~new_n23773_;
  assign new_n23775_ = ~new_n23771_ & new_n23774_;
  assign new_n23776_ = new_n19029_ & new_n21081_;
  assign new_n23777_ = new_n19029_ & new_n21068_;
  assign new_n23778_ = new_n19029_ & new_n21079_;
  assign new_n23779_ = ~new_n23777_ & ~new_n23778_;
  assign new_n23780_ = ~new_n23776_ & new_n23779_;
  assign new_n23781_ = new_n23775_ & new_n23780_;
  assign new_n23782_ = new_n19029_ & new_n21089_;
  assign new_n23783_ = new_n19029_ & new_n21077_;
  assign new_n23784_ = new_n19029_ & new_n21087_;
  assign new_n23785_ = ~new_n23783_ & ~new_n23784_;
  assign new_n23786_ = ~new_n23782_ & new_n23785_;
  assign new_n23787_ = new_n19029_ & new_n21098_;
  assign new_n23788_ = new_n19029_ & new_n21085_;
  assign new_n23789_ = new_n19029_ & new_n21096_;
  assign new_n23790_ = ~new_n23788_ & ~new_n23789_;
  assign new_n23791_ = ~new_n23787_ & new_n23790_;
  assign new_n23792_ = new_n23786_ & new_n23791_;
  assign new_n23793_ = new_n23781_ & new_n23792_;
  assign new_n23794_ = new_n19029_ & new_n21106_;
  assign new_n23795_ = new_n19029_ & new_n21094_;
  assign new_n23796_ = new_n19029_ & new_n21104_;
  assign new_n23797_ = ~new_n23795_ & ~new_n23796_;
  assign new_n23798_ = ~new_n23794_ & new_n23797_;
  assign new_n23799_ = new_n19029_ & new_n21116_;
  assign new_n23800_ = new_n19029_ & new_n21102_;
  assign new_n23801_ = new_n19029_ & new_n21114_;
  assign new_n23802_ = ~new_n23800_ & ~new_n23801_;
  assign new_n23803_ = ~new_n23799_ & new_n23802_;
  assign new_n23804_ = new_n23798_ & new_n23803_;
  assign new_n23805_ = new_n19076_ & new_n21019_;
  assign new_n23806_ = new_n19029_ & new_n21112_;
  assign new_n23807_ = new_n19076_ & new_n21017_;
  assign new_n23808_ = ~new_n23806_ & ~new_n23807_;
  assign new_n23809_ = ~new_n23805_ & new_n23808_;
  assign new_n23810_ = new_n19076_ & new_n21015_;
  assign new_n23811_ = new_n19076_ & new_n21026_;
  assign new_n23812_ = ~new_n23810_ & ~new_n23811_;
  assign new_n23813_ = new_n23809_ & new_n23812_;
  assign new_n23814_ = new_n23804_ & new_n23813_;
  assign new_n23815_ = new_n23793_ & new_n23814_;
  assign new_n23816_ = new_n19076_ & new_n21039_;
  assign new_n23817_ = new_n19076_ & new_n21029_;
  assign new_n23818_ = new_n19076_ & new_n21024_;
  assign new_n23819_ = ~new_n23817_ & ~new_n23818_;
  assign new_n23820_ = ~new_n23816_ & new_n23819_;
  assign new_n23821_ = new_n19076_ & new_n21050_;
  assign new_n23822_ = new_n19076_ & new_n21042_;
  assign new_n23823_ = new_n19076_ & new_n21036_;
  assign new_n23824_ = ~new_n23822_ & ~new_n23823_;
  assign new_n23825_ = ~new_n23821_ & new_n23824_;
  assign new_n23826_ = new_n23820_ & new_n23825_;
  assign new_n23827_ = new_n19076_ & new_n21060_;
  assign new_n23828_ = new_n19076_ & new_n21053_;
  assign new_n23829_ = new_n19076_ & new_n21047_;
  assign new_n23830_ = ~new_n23828_ & ~new_n23829_;
  assign new_n23831_ = ~new_n23827_ & new_n23830_;
  assign new_n23832_ = new_n19076_ & new_n21066_;
  assign new_n23833_ = new_n19076_ & new_n21062_;
  assign new_n23834_ = new_n19076_ & new_n21058_;
  assign new_n23835_ = ~new_n23833_ & ~new_n23834_;
  assign new_n23836_ = ~new_n23832_ & new_n23835_;
  assign new_n23837_ = new_n23831_ & new_n23836_;
  assign new_n23838_ = new_n23826_ & new_n23837_;
  assign new_n23839_ = new_n19076_ & new_n21081_;
  assign new_n23840_ = new_n19076_ & new_n21068_;
  assign new_n23841_ = new_n19076_ & new_n21079_;
  assign new_n23842_ = ~new_n23840_ & ~new_n23841_;
  assign new_n23843_ = ~new_n23839_ & new_n23842_;
  assign new_n23844_ = new_n19076_ & new_n21089_;
  assign new_n23845_ = new_n19076_ & new_n21077_;
  assign new_n23846_ = new_n19076_ & new_n21087_;
  assign new_n23847_ = ~new_n23845_ & ~new_n23846_;
  assign new_n23848_ = ~new_n23844_ & new_n23847_;
  assign new_n23849_ = new_n23843_ & new_n23848_;
  assign new_n23850_ = new_n19076_ & new_n21098_;
  assign new_n23851_ = new_n19076_ & new_n21085_;
  assign new_n23852_ = new_n19076_ & new_n21096_;
  assign new_n23853_ = ~new_n23851_ & ~new_n23852_;
  assign new_n23854_ = ~new_n23850_ & new_n23853_;
  assign new_n23855_ = new_n19076_ & new_n21094_;
  assign new_n23856_ = new_n19076_ & new_n21104_;
  assign new_n23857_ = ~new_n23855_ & ~new_n23856_;
  assign new_n23858_ = new_n23854_ & new_n23857_;
  assign new_n23859_ = new_n23849_ & new_n23858_;
  assign new_n23860_ = new_n23838_ & new_n23859_;
  assign new_n23861_ = new_n23815_ & new_n23860_;
  assign new_n23862_ = new_n23770_ & new_n23861_;
  assign new_n23863_ = new_n19076_ & new_n21114_;
  assign new_n23864_ = new_n19076_ & new_n21106_;
  assign new_n23865_ = new_n19076_ & new_n21102_;
  assign new_n23866_ = ~new_n23864_ & ~new_n23865_;
  assign new_n23867_ = ~new_n23863_ & new_n23866_;
  assign new_n23868_ = new_n19191_ & new_n21017_;
  assign new_n23869_ = new_n19076_ & new_n21116_;
  assign new_n23870_ = new_n19076_ & new_n21112_;
  assign new_n23871_ = ~new_n23869_ & ~new_n23870_;
  assign new_n23872_ = ~new_n23868_ & new_n23871_;
  assign new_n23873_ = new_n23867_ & new_n23872_;
  assign new_n23874_ = new_n19191_ & new_n21026_;
  assign new_n23875_ = new_n19191_ & new_n21019_;
  assign new_n23876_ = new_n19191_ & new_n21015_;
  assign new_n23877_ = ~new_n23875_ & ~new_n23876_;
  assign new_n23878_ = ~new_n23874_ & new_n23877_;
  assign new_n23879_ = new_n19191_ & new_n21039_;
  assign new_n23880_ = new_n19191_ & new_n21029_;
  assign new_n23881_ = new_n19191_ & new_n21024_;
  assign new_n23882_ = ~new_n23880_ & ~new_n23881_;
  assign new_n23883_ = ~new_n23879_ & new_n23882_;
  assign new_n23884_ = new_n23878_ & new_n23883_;
  assign new_n23885_ = new_n23873_ & new_n23884_;
  assign new_n23886_ = new_n19191_ & new_n21050_;
  assign new_n23887_ = new_n19191_ & new_n21042_;
  assign new_n23888_ = new_n19191_ & new_n21036_;
  assign new_n23889_ = ~new_n23887_ & ~new_n23888_;
  assign new_n23890_ = ~new_n23886_ & new_n23889_;
  assign new_n23891_ = new_n19191_ & new_n21060_;
  assign new_n23892_ = new_n19191_ & new_n21053_;
  assign new_n23893_ = new_n19191_ & new_n21047_;
  assign new_n23894_ = ~new_n23892_ & ~new_n23893_;
  assign new_n23895_ = ~new_n23891_ & new_n23894_;
  assign new_n23896_ = new_n23890_ & new_n23895_;
  assign new_n23897_ = new_n19191_ & new_n21066_;
  assign new_n23898_ = new_n19191_ & new_n21062_;
  assign new_n23899_ = new_n19191_ & new_n21058_;
  assign new_n23900_ = ~new_n23898_ & ~new_n23899_;
  assign new_n23901_ = ~new_n23897_ & new_n23900_;
  assign new_n23902_ = new_n19191_ & new_n21068_;
  assign new_n23903_ = new_n19191_ & new_n21079_;
  assign new_n23904_ = ~new_n23902_ & ~new_n23903_;
  assign new_n23905_ = new_n23901_ & new_n23904_;
  assign new_n23906_ = new_n23896_ & new_n23905_;
  assign new_n23907_ = new_n23885_ & new_n23906_;
  assign new_n23908_ = new_n19191_ & new_n21087_;
  assign new_n23909_ = new_n19191_ & new_n21081_;
  assign new_n23910_ = new_n19191_ & new_n21077_;
  assign new_n23911_ = ~new_n23909_ & ~new_n23910_;
  assign new_n23912_ = ~new_n23908_ & new_n23911_;
  assign new_n23913_ = new_n19191_ & new_n21096_;
  assign new_n23914_ = new_n19191_ & new_n21089_;
  assign new_n23915_ = new_n19191_ & new_n21085_;
  assign new_n23916_ = ~new_n23914_ & ~new_n23915_;
  assign new_n23917_ = ~new_n23913_ & new_n23916_;
  assign new_n23918_ = new_n23912_ & new_n23917_;
  assign new_n23919_ = new_n19191_ & new_n21104_;
  assign new_n23920_ = new_n19191_ & new_n21098_;
  assign new_n23921_ = new_n19191_ & new_n21094_;
  assign new_n23922_ = ~new_n23920_ & ~new_n23921_;
  assign new_n23923_ = ~new_n23919_ & new_n23922_;
  assign new_n23924_ = new_n19191_ & new_n21114_;
  assign new_n23925_ = new_n19191_ & new_n21106_;
  assign new_n23926_ = new_n19191_ & new_n21102_;
  assign new_n23927_ = ~new_n23925_ & ~new_n23926_;
  assign new_n23928_ = ~new_n23924_ & new_n23927_;
  assign new_n23929_ = new_n23923_ & new_n23928_;
  assign new_n23930_ = new_n23918_ & new_n23929_;
  assign new_n23931_ = new_n19239_ & new_n21017_;
  assign new_n23932_ = new_n19191_ & new_n21116_;
  assign new_n23933_ = new_n19191_ & new_n21112_;
  assign new_n23934_ = ~new_n23932_ & ~new_n23933_;
  assign new_n23935_ = ~new_n23931_ & new_n23934_;
  assign new_n23936_ = new_n19239_ & new_n21026_;
  assign new_n23937_ = new_n19239_ & new_n21019_;
  assign new_n23938_ = new_n19239_ & new_n21015_;
  assign new_n23939_ = ~new_n23937_ & ~new_n23938_;
  assign new_n23940_ = ~new_n23936_ & new_n23939_;
  assign new_n23941_ = new_n23935_ & new_n23940_;
  assign new_n23942_ = new_n19239_ & new_n21039_;
  assign new_n23943_ = new_n19239_ & new_n21029_;
  assign new_n23944_ = new_n19239_ & new_n21024_;
  assign new_n23945_ = ~new_n23943_ & ~new_n23944_;
  assign new_n23946_ = ~new_n23942_ & new_n23945_;
  assign new_n23947_ = new_n19239_ & new_n21042_;
  assign new_n23948_ = new_n19239_ & new_n21036_;
  assign new_n23949_ = ~new_n23947_ & ~new_n23948_;
  assign new_n23950_ = new_n23946_ & new_n23949_;
  assign new_n23951_ = new_n23941_ & new_n23950_;
  assign new_n23952_ = new_n23930_ & new_n23951_;
  assign new_n23953_ = new_n23907_ & new_n23952_;
  assign new_n23954_ = new_n19239_ & new_n21047_;
  assign new_n23955_ = new_n19239_ & new_n21050_;
  assign new_n23956_ = new_n19239_ & new_n21053_;
  assign new_n23957_ = ~new_n23955_ & ~new_n23956_;
  assign new_n23958_ = ~new_n23954_ & new_n23957_;
  assign new_n23959_ = new_n19239_ & new_n21058_;
  assign new_n23960_ = new_n19239_ & new_n21060_;
  assign new_n23961_ = new_n19239_ & new_n21062_;
  assign new_n23962_ = ~new_n23960_ & ~new_n23961_;
  assign new_n23963_ = ~new_n23959_ & new_n23962_;
  assign new_n23964_ = new_n23958_ & new_n23963_;
  assign new_n23965_ = new_n19239_ & new_n21079_;
  assign new_n23966_ = new_n19239_ & new_n21066_;
  assign new_n23967_ = new_n19239_ & new_n21068_;
  assign new_n23968_ = ~new_n23966_ & ~new_n23967_;
  assign new_n23969_ = ~new_n23965_ & new_n23968_;
  assign new_n23970_ = new_n19239_ & new_n21087_;
  assign new_n23971_ = new_n19239_ & new_n21081_;
  assign new_n23972_ = new_n19239_ & new_n21077_;
  assign new_n23973_ = ~new_n23971_ & ~new_n23972_;
  assign new_n23974_ = ~new_n23970_ & new_n23973_;
  assign new_n23975_ = new_n23969_ & new_n23974_;
  assign new_n23976_ = new_n23964_ & new_n23975_;
  assign new_n23977_ = new_n19239_ & new_n21096_;
  assign new_n23978_ = new_n19239_ & new_n21089_;
  assign new_n23979_ = new_n19239_ & new_n21085_;
  assign new_n23980_ = ~new_n23978_ & ~new_n23979_;
  assign new_n23981_ = ~new_n23977_ & new_n23980_;
  assign new_n23982_ = new_n19239_ & new_n21104_;
  assign new_n23983_ = new_n19239_ & new_n21098_;
  assign new_n23984_ = new_n19239_ & new_n21094_;
  assign new_n23985_ = ~new_n23983_ & ~new_n23984_;
  assign new_n23986_ = ~new_n23982_ & new_n23985_;
  assign new_n23987_ = new_n23981_ & new_n23986_;
  assign new_n23988_ = new_n19239_ & new_n21114_;
  assign new_n23989_ = new_n19239_ & new_n21106_;
  assign new_n23990_ = new_n19239_ & new_n21102_;
  assign new_n23991_ = ~new_n23989_ & ~new_n23990_;
  assign new_n23992_ = ~new_n23988_ & new_n23991_;
  assign new_n23993_ = new_n19239_ & new_n21116_;
  assign new_n23994_ = new_n19239_ & new_n21112_;
  assign new_n23995_ = ~new_n23993_ & ~new_n23994_;
  assign new_n23996_ = new_n23992_ & new_n23995_;
  assign new_n23997_ = new_n23987_ & new_n23996_;
  assign new_n23998_ = new_n23976_ & new_n23997_;
  assign new_n23999_ = new_n19293_ & new_n21015_;
  assign new_n24000_ = new_n19293_ & new_n21017_;
  assign new_n24001_ = new_n19293_ & new_n21019_;
  assign new_n24002_ = ~new_n24000_ & ~new_n24001_;
  assign new_n24003_ = ~new_n23999_ & new_n24002_;
  assign new_n24004_ = new_n19293_ & new_n21024_;
  assign new_n24005_ = new_n19293_ & new_n21026_;
  assign new_n24006_ = new_n19293_ & new_n21029_;
  assign new_n24007_ = ~new_n24005_ & ~new_n24006_;
  assign new_n24008_ = ~new_n24004_ & new_n24007_;
  assign new_n24009_ = new_n24003_ & new_n24008_;
  assign new_n24010_ = new_n19293_ & new_n21036_;
  assign new_n24011_ = new_n19293_ & new_n21039_;
  assign new_n24012_ = new_n19293_ & new_n21042_;
  assign new_n24013_ = ~new_n24011_ & ~new_n24012_;
  assign new_n24014_ = ~new_n24010_ & new_n24013_;
  assign new_n24015_ = new_n19293_ & new_n21047_;
  assign new_n24016_ = new_n19293_ & new_n21050_;
  assign new_n24017_ = new_n19293_ & new_n21053_;
  assign new_n24018_ = ~new_n24016_ & ~new_n24017_;
  assign new_n24019_ = ~new_n24015_ & new_n24018_;
  assign new_n24020_ = new_n24014_ & new_n24019_;
  assign new_n24021_ = new_n24009_ & new_n24020_;
  assign new_n24022_ = new_n19293_ & new_n21058_;
  assign new_n24023_ = new_n19293_ & new_n21060_;
  assign new_n24024_ = new_n19293_ & new_n21062_;
  assign new_n24025_ = ~new_n24023_ & ~new_n24024_;
  assign new_n24026_ = ~new_n24022_ & new_n24025_;
  assign new_n24027_ = new_n19293_ & new_n21079_;
  assign new_n24028_ = new_n19293_ & new_n21066_;
  assign new_n24029_ = new_n19293_ & new_n21068_;
  assign new_n24030_ = ~new_n24028_ & ~new_n24029_;
  assign new_n24031_ = ~new_n24027_ & new_n24030_;
  assign new_n24032_ = new_n24026_ & new_n24031_;
  assign new_n24033_ = new_n19293_ & new_n21087_;
  assign new_n24034_ = new_n19293_ & new_n21081_;
  assign new_n24035_ = new_n19293_ & new_n21077_;
  assign new_n24036_ = ~new_n24034_ & ~new_n24035_;
  assign new_n24037_ = ~new_n24033_ & new_n24036_;
  assign new_n24038_ = new_n19293_ & new_n21089_;
  assign new_n24039_ = new_n19293_ & new_n21085_;
  assign new_n24040_ = ~new_n24038_ & ~new_n24039_;
  assign new_n24041_ = new_n24037_ & new_n24040_;
  assign new_n24042_ = new_n24032_ & new_n24041_;
  assign new_n24043_ = new_n24021_ & new_n24042_;
  assign new_n24044_ = new_n23998_ & new_n24043_;
  assign new_n24045_ = new_n23953_ & new_n24044_;
  assign new_n24046_ = new_n23862_ & new_n24045_;
  assign new_n24047_ = new_n19293_ & new_n21094_;
  assign new_n24048_ = new_n19293_ & new_n21096_;
  assign new_n24049_ = new_n19293_ & new_n21098_;
  assign new_n24050_ = ~new_n24048_ & ~new_n24049_;
  assign new_n24051_ = ~new_n24047_ & new_n24050_;
  assign new_n24052_ = new_n19293_ & new_n21102_;
  assign new_n24053_ = new_n19293_ & new_n21104_;
  assign new_n24054_ = new_n19293_ & new_n21106_;
  assign new_n24055_ = ~new_n24053_ & ~new_n24054_;
  assign new_n24056_ = ~new_n24052_ & new_n24055_;
  assign new_n24057_ = new_n24051_ & new_n24056_;
  assign new_n24058_ = new_n19293_ & new_n21112_;
  assign new_n24059_ = new_n19293_ & new_n21114_;
  assign new_n24060_ = new_n19293_ & new_n21116_;
  assign new_n24061_ = ~new_n24059_ & ~new_n24060_;
  assign new_n24062_ = ~new_n24058_ & new_n24061_;
  assign new_n24063_ = new_n19339_ & new_n21015_;
  assign new_n24064_ = new_n19339_ & new_n21017_;
  assign new_n24065_ = new_n19339_ & new_n21019_;
  assign new_n24066_ = ~new_n24064_ & ~new_n24065_;
  assign new_n24067_ = ~new_n24063_ & new_n24066_;
  assign new_n24068_ = new_n24062_ & new_n24067_;
  assign new_n24069_ = new_n24057_ & new_n24068_;
  assign new_n24070_ = new_n19339_ & new_n21024_;
  assign new_n24071_ = new_n19339_ & new_n21026_;
  assign new_n24072_ = new_n19339_ & new_n21029_;
  assign new_n24073_ = ~new_n24071_ & ~new_n24072_;
  assign new_n24074_ = ~new_n24070_ & new_n24073_;
  assign new_n24075_ = new_n19339_ & new_n21036_;
  assign new_n24076_ = new_n19339_ & new_n21039_;
  assign new_n24077_ = new_n19339_ & new_n21042_;
  assign new_n24078_ = ~new_n24076_ & ~new_n24077_;
  assign new_n24079_ = ~new_n24075_ & new_n24078_;
  assign new_n24080_ = new_n24074_ & new_n24079_;
  assign new_n24081_ = new_n19339_ & new_n21047_;
  assign new_n24082_ = new_n19339_ & new_n21050_;
  assign new_n24083_ = new_n19339_ & new_n21053_;
  assign new_n24084_ = ~new_n24082_ & ~new_n24083_;
  assign new_n24085_ = ~new_n24081_ & new_n24084_;
  assign new_n24086_ = new_n19339_ & new_n21060_;
  assign new_n24087_ = new_n19339_ & new_n21062_;
  assign new_n24088_ = ~new_n24086_ & ~new_n24087_;
  assign new_n24089_ = new_n24085_ & new_n24088_;
  assign new_n24090_ = new_n24080_ & new_n24089_;
  assign new_n24091_ = new_n24069_ & new_n24090_;
  assign new_n24092_ = new_n19339_ & new_n21068_;
  assign new_n24093_ = new_n19339_ & new_n21058_;
  assign new_n24094_ = new_n19339_ & new_n21066_;
  assign new_n24095_ = ~new_n24093_ & ~new_n24094_;
  assign new_n24096_ = ~new_n24092_ & new_n24095_;
  assign new_n24097_ = new_n19339_ & new_n21077_;
  assign new_n24098_ = new_n19339_ & new_n21079_;
  assign new_n24099_ = new_n19339_ & new_n21081_;
  assign new_n24100_ = ~new_n24098_ & ~new_n24099_;
  assign new_n24101_ = ~new_n24097_ & new_n24100_;
  assign new_n24102_ = new_n24096_ & new_n24101_;
  assign new_n24103_ = new_n19339_ & new_n21085_;
  assign new_n24104_ = new_n19339_ & new_n21087_;
  assign new_n24105_ = new_n19339_ & new_n21089_;
  assign new_n24106_ = ~new_n24104_ & ~new_n24105_;
  assign new_n24107_ = ~new_n24103_ & new_n24106_;
  assign new_n24108_ = new_n19339_ & new_n21094_;
  assign new_n24109_ = new_n19339_ & new_n21096_;
  assign new_n24110_ = new_n19339_ & new_n21098_;
  assign new_n24111_ = ~new_n24109_ & ~new_n24110_;
  assign new_n24112_ = ~new_n24108_ & new_n24111_;
  assign new_n24113_ = new_n24107_ & new_n24112_;
  assign new_n24114_ = new_n24102_ & new_n24113_;
  assign new_n24115_ = new_n19339_ & new_n21102_;
  assign new_n24116_ = new_n19339_ & new_n21104_;
  assign new_n24117_ = new_n19339_ & new_n21106_;
  assign new_n24118_ = ~new_n24116_ & ~new_n24117_;
  assign new_n24119_ = ~new_n24115_ & new_n24118_;
  assign new_n24120_ = new_n19339_ & new_n21112_;
  assign new_n24121_ = new_n19339_ & new_n21114_;
  assign new_n24122_ = new_n19339_ & new_n21116_;
  assign new_n24123_ = ~new_n24121_ & ~new_n24122_;
  assign new_n24124_ = ~new_n24120_ & new_n24123_;
  assign new_n24125_ = new_n24119_ & new_n24124_;
  assign new_n24126_ = new_n19713_ & new_n21015_;
  assign new_n24127_ = new_n19713_ & new_n21017_;
  assign new_n24128_ = new_n19713_ & new_n21019_;
  assign new_n24129_ = ~new_n24127_ & ~new_n24128_;
  assign new_n24130_ = ~new_n24126_ & new_n24129_;
  assign new_n24131_ = new_n19713_ & new_n21026_;
  assign new_n24132_ = new_n19713_ & new_n21029_;
  assign new_n24133_ = ~new_n24131_ & ~new_n24132_;
  assign new_n24134_ = new_n24130_ & new_n24133_;
  assign new_n24135_ = new_n24125_ & new_n24134_;
  assign new_n24136_ = new_n24114_ & new_n24135_;
  assign new_n24137_ = new_n24091_ & new_n24136_;
  assign new_n24138_ = new_n19713_ & new_n21042_;
  assign new_n24139_ = new_n19713_ & new_n21024_;
  assign new_n24140_ = new_n19713_ & new_n21039_;
  assign new_n24141_ = ~new_n24139_ & ~new_n24140_;
  assign new_n24142_ = ~new_n24138_ & new_n24141_;
  assign new_n24143_ = new_n19713_ & new_n21053_;
  assign new_n24144_ = new_n19713_ & new_n21036_;
  assign new_n24145_ = new_n19713_ & new_n21050_;
  assign new_n24146_ = ~new_n24144_ & ~new_n24145_;
  assign new_n24147_ = ~new_n24143_ & new_n24146_;
  assign new_n24148_ = new_n24142_ & new_n24147_;
  assign new_n24149_ = new_n19713_ & new_n21062_;
  assign new_n24150_ = new_n19713_ & new_n21047_;
  assign new_n24151_ = new_n19713_ & new_n21060_;
  assign new_n24152_ = ~new_n24150_ & ~new_n24151_;
  assign new_n24153_ = ~new_n24149_ & new_n24152_;
  assign new_n24154_ = new_n19713_ & new_n21068_;
  assign new_n24155_ = new_n19713_ & new_n21058_;
  assign new_n24156_ = new_n19713_ & new_n21066_;
  assign new_n24157_ = ~new_n24155_ & ~new_n24156_;
  assign new_n24158_ = ~new_n24154_ & new_n24157_;
  assign new_n24159_ = new_n24153_ & new_n24158_;
  assign new_n24160_ = new_n24148_ & new_n24159_;
  assign new_n24161_ = new_n19713_ & new_n21077_;
  assign new_n24162_ = new_n19713_ & new_n21079_;
  assign new_n24163_ = new_n19713_ & new_n21081_;
  assign new_n24164_ = ~new_n24162_ & ~new_n24163_;
  assign new_n24165_ = ~new_n24161_ & new_n24164_;
  assign new_n24166_ = new_n19713_ & new_n21085_;
  assign new_n24167_ = new_n19713_ & new_n21087_;
  assign new_n24168_ = new_n19713_ & new_n21089_;
  assign new_n24169_ = ~new_n24167_ & ~new_n24168_;
  assign new_n24170_ = ~new_n24166_ & new_n24169_;
  assign new_n24171_ = new_n24165_ & new_n24170_;
  assign new_n24172_ = new_n19713_ & new_n21094_;
  assign new_n24173_ = new_n19713_ & new_n21096_;
  assign new_n24174_ = new_n19713_ & new_n21098_;
  assign new_n24175_ = ~new_n24173_ & ~new_n24174_;
  assign new_n24176_ = ~new_n24172_ & new_n24175_;
  assign new_n24177_ = new_n19713_ & new_n21104_;
  assign new_n24178_ = new_n19713_ & new_n21106_;
  assign new_n24179_ = ~new_n24177_ & ~new_n24178_;
  assign new_n24180_ = new_n24176_ & new_n24179_;
  assign new_n24181_ = new_n24171_ & new_n24180_;
  assign new_n24182_ = new_n24160_ & new_n24181_;
  assign new_n24183_ = new_n19713_ & new_n21116_;
  assign new_n24184_ = new_n19713_ & new_n21102_;
  assign new_n24185_ = new_n19713_ & new_n21114_;
  assign new_n24186_ = ~new_n24184_ & ~new_n24185_;
  assign new_n24187_ = ~new_n24183_ & new_n24186_;
  assign new_n24188_ = new_n19761_ & new_n21019_;
  assign new_n24189_ = new_n19713_ & new_n21112_;
  assign new_n24190_ = new_n19761_ & new_n21017_;
  assign new_n24191_ = ~new_n24189_ & ~new_n24190_;
  assign new_n24192_ = ~new_n24188_ & new_n24191_;
  assign new_n24193_ = new_n24187_ & new_n24192_;
  assign new_n24194_ = new_n19761_ & new_n21029_;
  assign new_n24195_ = new_n19761_ & new_n21015_;
  assign new_n24196_ = new_n19761_ & new_n21026_;
  assign new_n24197_ = ~new_n24195_ & ~new_n24196_;
  assign new_n24198_ = ~new_n24194_ & new_n24197_;
  assign new_n24199_ = new_n19761_ & new_n21042_;
  assign new_n24200_ = new_n19761_ & new_n21024_;
  assign new_n24201_ = new_n19761_ & new_n21039_;
  assign new_n24202_ = ~new_n24200_ & ~new_n24201_;
  assign new_n24203_ = ~new_n24199_ & new_n24202_;
  assign new_n24204_ = new_n24198_ & new_n24203_;
  assign new_n24205_ = new_n24193_ & new_n24204_;
  assign new_n24206_ = new_n19761_ & new_n21053_;
  assign new_n24207_ = new_n19761_ & new_n21036_;
  assign new_n24208_ = new_n19761_ & new_n21050_;
  assign new_n24209_ = ~new_n24207_ & ~new_n24208_;
  assign new_n24210_ = ~new_n24206_ & new_n24209_;
  assign new_n24211_ = new_n19761_ & new_n21062_;
  assign new_n24212_ = new_n19761_ & new_n21047_;
  assign new_n24213_ = new_n19761_ & new_n21060_;
  assign new_n24214_ = ~new_n24212_ & ~new_n24213_;
  assign new_n24215_ = ~new_n24211_ & new_n24214_;
  assign new_n24216_ = new_n24210_ & new_n24215_;
  assign new_n24217_ = new_n19761_ & new_n21068_;
  assign new_n24218_ = new_n19761_ & new_n21058_;
  assign new_n24219_ = new_n19761_ & new_n21066_;
  assign new_n24220_ = ~new_n24218_ & ~new_n24219_;
  assign new_n24221_ = ~new_n24217_ & new_n24220_;
  assign new_n24222_ = new_n19761_ & new_n21079_;
  assign new_n24223_ = new_n19761_ & new_n21081_;
  assign new_n24224_ = ~new_n24222_ & ~new_n24223_;
  assign new_n24225_ = new_n24221_ & new_n24224_;
  assign new_n24226_ = new_n24216_ & new_n24225_;
  assign new_n24227_ = new_n24205_ & new_n24226_;
  assign new_n24228_ = new_n24182_ & new_n24227_;
  assign new_n24229_ = new_n24137_ & new_n24228_;
  assign new_n24230_ = new_n19761_ & new_n21089_;
  assign new_n24231_ = new_n19761_ & new_n21077_;
  assign new_n24232_ = new_n19761_ & new_n21087_;
  assign new_n24233_ = ~new_n24231_ & ~new_n24232_;
  assign new_n24234_ = ~new_n24230_ & new_n24233_;
  assign new_n24235_ = new_n19761_ & new_n21098_;
  assign new_n24236_ = new_n19761_ & new_n21085_;
  assign new_n24237_ = new_n19761_ & new_n21096_;
  assign new_n24238_ = ~new_n24236_ & ~new_n24237_;
  assign new_n24239_ = ~new_n24235_ & new_n24238_;
  assign new_n24240_ = new_n24234_ & new_n24239_;
  assign new_n24241_ = new_n19761_ & new_n21106_;
  assign new_n24242_ = new_n19761_ & new_n21094_;
  assign new_n24243_ = new_n19761_ & new_n21104_;
  assign new_n24244_ = ~new_n24242_ & ~new_n24243_;
  assign new_n24245_ = ~new_n24241_ & new_n24244_;
  assign new_n24246_ = new_n19761_ & new_n21116_;
  assign new_n24247_ = new_n19761_ & new_n21102_;
  assign new_n24248_ = new_n19761_ & new_n21114_;
  assign new_n24249_ = ~new_n24247_ & ~new_n24248_;
  assign new_n24250_ = ~new_n24246_ & new_n24249_;
  assign new_n24251_ = new_n24245_ & new_n24250_;
  assign new_n24252_ = new_n24240_ & new_n24251_;
  assign new_n24253_ = new_n19807_ & new_n21019_;
  assign new_n24254_ = new_n19761_ & new_n21112_;
  assign new_n24255_ = new_n19807_ & new_n21017_;
  assign new_n24256_ = ~new_n24254_ & ~new_n24255_;
  assign new_n24257_ = ~new_n24253_ & new_n24256_;
  assign new_n24258_ = new_n19807_ & new_n21029_;
  assign new_n24259_ = new_n19807_ & new_n21015_;
  assign new_n24260_ = new_n19807_ & new_n21026_;
  assign new_n24261_ = ~new_n24259_ & ~new_n24260_;
  assign new_n24262_ = ~new_n24258_ & new_n24261_;
  assign new_n24263_ = new_n24257_ & new_n24262_;
  assign new_n24264_ = new_n19807_ & new_n21042_;
  assign new_n24265_ = new_n19807_ & new_n21024_;
  assign new_n24266_ = new_n19807_ & new_n21039_;
  assign new_n24267_ = ~new_n24265_ & ~new_n24266_;
  assign new_n24268_ = ~new_n24264_ & new_n24267_;
  assign new_n24269_ = new_n19807_ & new_n21036_;
  assign new_n24270_ = new_n19807_ & new_n21050_;
  assign new_n24271_ = ~new_n24269_ & ~new_n24270_;
  assign new_n24272_ = new_n24268_ & new_n24271_;
  assign new_n24273_ = new_n24263_ & new_n24272_;
  assign new_n24274_ = new_n24252_ & new_n24273_;
  assign new_n24275_ = new_n19807_ & new_n21060_;
  assign new_n24276_ = new_n19807_ & new_n21053_;
  assign new_n24277_ = new_n19807_ & new_n21047_;
  assign new_n24278_ = ~new_n24276_ & ~new_n24277_;
  assign new_n24279_ = ~new_n24275_ & new_n24278_;
  assign new_n24280_ = new_n19807_ & new_n21066_;
  assign new_n24281_ = new_n19807_ & new_n21062_;
  assign new_n24282_ = new_n19807_ & new_n21058_;
  assign new_n24283_ = ~new_n24281_ & ~new_n24282_;
  assign new_n24284_ = ~new_n24280_ & new_n24283_;
  assign new_n24285_ = new_n24279_ & new_n24284_;
  assign new_n24286_ = new_n19807_ & new_n21081_;
  assign new_n24287_ = new_n19807_ & new_n21068_;
  assign new_n24288_ = new_n19807_ & new_n21079_;
  assign new_n24289_ = ~new_n24287_ & ~new_n24288_;
  assign new_n24290_ = ~new_n24286_ & new_n24289_;
  assign new_n24291_ = new_n19807_ & new_n21089_;
  assign new_n24292_ = new_n19807_ & new_n21077_;
  assign new_n24293_ = new_n19807_ & new_n21087_;
  assign new_n24294_ = ~new_n24292_ & ~new_n24293_;
  assign new_n24295_ = ~new_n24291_ & new_n24294_;
  assign new_n24296_ = new_n24290_ & new_n24295_;
  assign new_n24297_ = new_n24285_ & new_n24296_;
  assign new_n24298_ = new_n19807_ & new_n21098_;
  assign new_n24299_ = new_n19807_ & new_n21085_;
  assign new_n24300_ = new_n19807_ & new_n21096_;
  assign new_n24301_ = ~new_n24299_ & ~new_n24300_;
  assign new_n24302_ = ~new_n24298_ & new_n24301_;
  assign new_n24303_ = new_n19807_ & new_n21106_;
  assign new_n24304_ = new_n19807_ & new_n21094_;
  assign new_n24305_ = new_n19807_ & new_n21104_;
  assign new_n24306_ = ~new_n24304_ & ~new_n24305_;
  assign new_n24307_ = ~new_n24303_ & new_n24306_;
  assign new_n24308_ = new_n24302_ & new_n24307_;
  assign new_n24309_ = new_n19807_ & new_n21116_;
  assign new_n24310_ = new_n19807_ & new_n21102_;
  assign new_n24311_ = new_n19807_ & new_n21114_;
  assign new_n24312_ = ~new_n24310_ & ~new_n24311_;
  assign new_n24313_ = ~new_n24309_ & new_n24312_;
  assign new_n24314_ = new_n19807_ & new_n21112_;
  assign new_n24315_ = new_n19859_ & new_n21017_;
  assign new_n24316_ = ~new_n24314_ & ~new_n24315_;
  assign new_n24317_ = new_n24313_ & new_n24316_;
  assign new_n24318_ = new_n24308_ & new_n24317_;
  assign new_n24319_ = new_n24297_ & new_n24318_;
  assign new_n24320_ = new_n24274_ & new_n24319_;
  assign new_n24321_ = new_n19859_ & new_n21026_;
  assign new_n24322_ = new_n19859_ & new_n21019_;
  assign new_n24323_ = new_n19859_ & new_n21015_;
  assign new_n24324_ = ~new_n24322_ & ~new_n24323_;
  assign new_n24325_ = ~new_n24321_ & new_n24324_;
  assign new_n24326_ = new_n19859_ & new_n21039_;
  assign new_n24327_ = new_n19859_ & new_n21029_;
  assign new_n24328_ = new_n19859_ & new_n21024_;
  assign new_n24329_ = ~new_n24327_ & ~new_n24328_;
  assign new_n24330_ = ~new_n24326_ & new_n24329_;
  assign new_n24331_ = new_n24325_ & new_n24330_;
  assign new_n24332_ = new_n19859_ & new_n21050_;
  assign new_n24333_ = new_n19859_ & new_n21042_;
  assign new_n24334_ = new_n19859_ & new_n21036_;
  assign new_n24335_ = ~new_n24333_ & ~new_n24334_;
  assign new_n24336_ = ~new_n24332_ & new_n24335_;
  assign new_n24337_ = new_n19859_ & new_n21060_;
  assign new_n24338_ = new_n19859_ & new_n21053_;
  assign new_n24339_ = new_n19859_ & new_n21047_;
  assign new_n24340_ = ~new_n24338_ & ~new_n24339_;
  assign new_n24341_ = ~new_n24337_ & new_n24340_;
  assign new_n24342_ = new_n24336_ & new_n24341_;
  assign new_n24343_ = new_n24331_ & new_n24342_;
  assign new_n24344_ = new_n19859_ & new_n21066_;
  assign new_n24345_ = new_n19859_ & new_n21062_;
  assign new_n24346_ = new_n19859_ & new_n21058_;
  assign new_n24347_ = ~new_n24345_ & ~new_n24346_;
  assign new_n24348_ = ~new_n24344_ & new_n24347_;
  assign new_n24349_ = new_n19859_ & new_n21081_;
  assign new_n24350_ = new_n19859_ & new_n21068_;
  assign new_n24351_ = new_n19859_ & new_n21079_;
  assign new_n24352_ = ~new_n24350_ & ~new_n24351_;
  assign new_n24353_ = ~new_n24349_ & new_n24352_;
  assign new_n24354_ = new_n24348_ & new_n24353_;
  assign new_n24355_ = new_n19859_ & new_n21089_;
  assign new_n24356_ = new_n19859_ & new_n21077_;
  assign new_n24357_ = new_n19859_ & new_n21087_;
  assign new_n24358_ = ~new_n24356_ & ~new_n24357_;
  assign new_n24359_ = ~new_n24355_ & new_n24358_;
  assign new_n24360_ = new_n19859_ & new_n21085_;
  assign new_n24361_ = new_n19859_ & new_n21096_;
  assign new_n24362_ = ~new_n24360_ & ~new_n24361_;
  assign new_n24363_ = new_n24359_ & new_n24362_;
  assign new_n24364_ = new_n24354_ & new_n24363_;
  assign new_n24365_ = new_n24343_ & new_n24364_;
  assign new_n24366_ = new_n19859_ & new_n21104_;
  assign new_n24367_ = new_n19859_ & new_n21098_;
  assign new_n24368_ = new_n19859_ & new_n21094_;
  assign new_n24369_ = ~new_n24367_ & ~new_n24368_;
  assign new_n24370_ = ~new_n24366_ & new_n24369_;
  assign new_n24371_ = new_n19859_ & new_n21114_;
  assign new_n24372_ = new_n19859_ & new_n21106_;
  assign new_n24373_ = new_n19859_ & new_n21102_;
  assign new_n24374_ = ~new_n24372_ & ~new_n24373_;
  assign new_n24375_ = ~new_n24371_ & new_n24374_;
  assign new_n24376_ = new_n24370_ & new_n24375_;
  assign new_n24377_ = new_n19974_ & new_n21017_;
  assign new_n24378_ = new_n19859_ & new_n21116_;
  assign new_n24379_ = new_n19859_ & new_n21112_;
  assign new_n24380_ = ~new_n24378_ & ~new_n24379_;
  assign new_n24381_ = ~new_n24377_ & new_n24380_;
  assign new_n24382_ = new_n19974_ & new_n21026_;
  assign new_n24383_ = new_n19974_ & new_n21019_;
  assign new_n24384_ = new_n19974_ & new_n21015_;
  assign new_n24385_ = ~new_n24383_ & ~new_n24384_;
  assign new_n24386_ = ~new_n24382_ & new_n24385_;
  assign new_n24387_ = new_n24381_ & new_n24386_;
  assign new_n24388_ = new_n24376_ & new_n24387_;
  assign new_n24389_ = new_n19974_ & new_n21039_;
  assign new_n24390_ = new_n19974_ & new_n21029_;
  assign new_n24391_ = new_n19974_ & new_n21024_;
  assign new_n24392_ = ~new_n24390_ & ~new_n24391_;
  assign new_n24393_ = ~new_n24389_ & new_n24392_;
  assign new_n24394_ = new_n19974_ & new_n21050_;
  assign new_n24395_ = new_n19974_ & new_n21042_;
  assign new_n24396_ = new_n19974_ & new_n21036_;
  assign new_n24397_ = ~new_n24395_ & ~new_n24396_;
  assign new_n24398_ = ~new_n24394_ & new_n24397_;
  assign new_n24399_ = new_n24393_ & new_n24398_;
  assign new_n24400_ = new_n19974_ & new_n21060_;
  assign new_n24401_ = new_n19974_ & new_n21053_;
  assign new_n24402_ = new_n19974_ & new_n21047_;
  assign new_n24403_ = ~new_n24401_ & ~new_n24402_;
  assign new_n24404_ = ~new_n24400_ & new_n24403_;
  assign new_n24405_ = new_n19974_ & new_n21062_;
  assign new_n24406_ = new_n19974_ & new_n21058_;
  assign new_n24407_ = ~new_n24405_ & ~new_n24406_;
  assign new_n24408_ = new_n24404_ & new_n24407_;
  assign new_n24409_ = new_n24399_ & new_n24408_;
  assign new_n24410_ = new_n24388_ & new_n24409_;
  assign new_n24411_ = new_n24365_ & new_n24410_;
  assign new_n24412_ = new_n24320_ & new_n24411_;
  assign new_n24413_ = new_n24229_ & new_n24412_;
  assign new_n24414_ = new_n24046_ & new_n24413_;
  assign new_n24415_ = new_n19974_ & new_n21079_;
  assign new_n24416_ = new_n19974_ & new_n21066_;
  assign new_n24417_ = new_n19974_ & new_n21068_;
  assign new_n24418_ = ~new_n24416_ & ~new_n24417_;
  assign new_n24419_ = ~new_n24415_ & new_n24418_;
  assign new_n24420_ = new_n19974_ & new_n21087_;
  assign new_n24421_ = new_n19974_ & new_n21081_;
  assign new_n24422_ = new_n19974_ & new_n21077_;
  assign new_n24423_ = ~new_n24421_ & ~new_n24422_;
  assign new_n24424_ = ~new_n24420_ & new_n24423_;
  assign new_n24425_ = new_n24419_ & new_n24424_;
  assign new_n24426_ = new_n19974_ & new_n21096_;
  assign new_n24427_ = new_n19974_ & new_n21089_;
  assign new_n24428_ = new_n19974_ & new_n21085_;
  assign new_n24429_ = ~new_n24427_ & ~new_n24428_;
  assign new_n24430_ = ~new_n24426_ & new_n24429_;
  assign new_n24431_ = new_n19974_ & new_n21104_;
  assign new_n24432_ = new_n19974_ & new_n21098_;
  assign new_n24433_ = new_n19974_ & new_n21094_;
  assign new_n24434_ = ~new_n24432_ & ~new_n24433_;
  assign new_n24435_ = ~new_n24431_ & new_n24434_;
  assign new_n24436_ = new_n24430_ & new_n24435_;
  assign new_n24437_ = new_n24425_ & new_n24436_;
  assign new_n24438_ = new_n19974_ & new_n21114_;
  assign new_n24439_ = new_n19974_ & new_n21106_;
  assign new_n24440_ = new_n19974_ & new_n21102_;
  assign new_n24441_ = ~new_n24439_ & ~new_n24440_;
  assign new_n24442_ = ~new_n24438_ & new_n24441_;
  assign new_n24443_ = new_n20021_ & new_n21017_;
  assign new_n24444_ = new_n19974_ & new_n21116_;
  assign new_n24445_ = new_n19974_ & new_n21112_;
  assign new_n24446_ = ~new_n24444_ & ~new_n24445_;
  assign new_n24447_ = ~new_n24443_ & new_n24446_;
  assign new_n24448_ = new_n24442_ & new_n24447_;
  assign new_n24449_ = new_n20021_ & new_n21026_;
  assign new_n24450_ = new_n20021_ & new_n21019_;
  assign new_n24451_ = new_n20021_ & new_n21015_;
  assign new_n24452_ = ~new_n24450_ & ~new_n24451_;
  assign new_n24453_ = ~new_n24449_ & new_n24452_;
  assign new_n24454_ = new_n20021_ & new_n21039_;
  assign new_n24455_ = new_n20021_ & new_n21029_;
  assign new_n24456_ = new_n20021_ & new_n21024_;
  assign new_n24457_ = ~new_n24455_ & ~new_n24456_;
  assign new_n24458_ = ~new_n24454_ & new_n24457_;
  assign new_n24459_ = new_n24453_ & new_n24458_;
  assign new_n24460_ = new_n24448_ & new_n24459_;
  assign new_n24461_ = new_n24437_ & new_n24460_;
  assign new_n24462_ = new_n20021_ & new_n21050_;
  assign new_n24463_ = new_n20021_ & new_n21042_;
  assign new_n24464_ = new_n20021_ & new_n21036_;
  assign new_n24465_ = ~new_n24463_ & ~new_n24464_;
  assign new_n24466_ = ~new_n24462_ & new_n24465_;
  assign new_n24467_ = new_n20021_ & new_n21060_;
  assign new_n24468_ = new_n20021_ & new_n21053_;
  assign new_n24469_ = new_n20021_ & new_n21047_;
  assign new_n24470_ = ~new_n24468_ & ~new_n24469_;
  assign new_n24471_ = ~new_n24467_ & new_n24470_;
  assign new_n24472_ = new_n24466_ & new_n24471_;
  assign new_n24473_ = new_n20021_ & new_n21066_;
  assign new_n24474_ = new_n20021_ & new_n21062_;
  assign new_n24475_ = new_n20021_ & new_n21058_;
  assign new_n24476_ = ~new_n24474_ & ~new_n24475_;
  assign new_n24477_ = ~new_n24473_ & new_n24476_;
  assign new_n24478_ = new_n20021_ & new_n21081_;
  assign new_n24479_ = new_n20021_ & new_n21068_;
  assign new_n24480_ = new_n20021_ & new_n21079_;
  assign new_n24481_ = ~new_n24479_ & ~new_n24480_;
  assign new_n24482_ = ~new_n24478_ & new_n24481_;
  assign new_n24483_ = new_n24477_ & new_n24482_;
  assign new_n24484_ = new_n24472_ & new_n24483_;
  assign new_n24485_ = new_n20021_ & new_n21089_;
  assign new_n24486_ = new_n20021_ & new_n21077_;
  assign new_n24487_ = new_n20021_ & new_n21087_;
  assign new_n24488_ = ~new_n24486_ & ~new_n24487_;
  assign new_n24489_ = ~new_n24485_ & new_n24488_;
  assign new_n24490_ = new_n20021_ & new_n21098_;
  assign new_n24491_ = new_n20021_ & new_n21085_;
  assign new_n24492_ = new_n20021_ & new_n21096_;
  assign new_n24493_ = ~new_n24491_ & ~new_n24492_;
  assign new_n24494_ = ~new_n24490_ & new_n24493_;
  assign new_n24495_ = new_n24489_ & new_n24494_;
  assign new_n24496_ = new_n20021_ & new_n21106_;
  assign new_n24497_ = new_n20021_ & new_n21094_;
  assign new_n24498_ = new_n20021_ & new_n21104_;
  assign new_n24499_ = ~new_n24497_ & ~new_n24498_;
  assign new_n24500_ = ~new_n24496_ & new_n24499_;
  assign new_n24501_ = new_n20021_ & new_n21102_;
  assign new_n24502_ = new_n20021_ & new_n21114_;
  assign new_n24503_ = ~new_n24501_ & ~new_n24502_;
  assign new_n24504_ = new_n24500_ & new_n24503_;
  assign new_n24505_ = new_n24495_ & new_n24504_;
  assign new_n24506_ = new_n24484_ & new_n24505_;
  assign new_n24507_ = new_n24461_ & new_n24506_;
  assign new_n24508_ = new_n20072_ & new_n21017_;
  assign new_n24509_ = new_n20021_ & new_n21116_;
  assign new_n24510_ = new_n20021_ & new_n21112_;
  assign new_n24511_ = ~new_n24509_ & ~new_n24510_;
  assign new_n24512_ = ~new_n24508_ & new_n24511_;
  assign new_n24513_ = new_n20072_ & new_n21026_;
  assign new_n24514_ = new_n20072_ & new_n21019_;
  assign new_n24515_ = new_n20072_ & new_n21015_;
  assign new_n24516_ = ~new_n24514_ & ~new_n24515_;
  assign new_n24517_ = ~new_n24513_ & new_n24516_;
  assign new_n24518_ = new_n24512_ & new_n24517_;
  assign new_n24519_ = new_n20072_ & new_n21039_;
  assign new_n24520_ = new_n20072_ & new_n21029_;
  assign new_n24521_ = new_n20072_ & new_n21024_;
  assign new_n24522_ = ~new_n24520_ & ~new_n24521_;
  assign new_n24523_ = ~new_n24519_ & new_n24522_;
  assign new_n24524_ = new_n20072_ & new_n21050_;
  assign new_n24525_ = new_n20072_ & new_n21042_;
  assign new_n24526_ = new_n20072_ & new_n21036_;
  assign new_n24527_ = ~new_n24525_ & ~new_n24526_;
  assign new_n24528_ = ~new_n24524_ & new_n24527_;
  assign new_n24529_ = new_n24523_ & new_n24528_;
  assign new_n24530_ = new_n24518_ & new_n24529_;
  assign new_n24531_ = new_n20072_ & new_n21060_;
  assign new_n24532_ = new_n20072_ & new_n21053_;
  assign new_n24533_ = new_n20072_ & new_n21047_;
  assign new_n24534_ = ~new_n24532_ & ~new_n24533_;
  assign new_n24535_ = ~new_n24531_ & new_n24534_;
  assign new_n24536_ = new_n20072_ & new_n21066_;
  assign new_n24537_ = new_n20072_ & new_n21062_;
  assign new_n24538_ = new_n20072_ & new_n21058_;
  assign new_n24539_ = ~new_n24537_ & ~new_n24538_;
  assign new_n24540_ = ~new_n24536_ & new_n24539_;
  assign new_n24541_ = new_n24535_ & new_n24540_;
  assign new_n24542_ = new_n20072_ & new_n21081_;
  assign new_n24543_ = new_n20072_ & new_n21068_;
  assign new_n24544_ = new_n20072_ & new_n21079_;
  assign new_n24545_ = ~new_n24543_ & ~new_n24544_;
  assign new_n24546_ = ~new_n24542_ & new_n24545_;
  assign new_n24547_ = new_n20072_ & new_n21077_;
  assign new_n24548_ = new_n20072_ & new_n21087_;
  assign new_n24549_ = ~new_n24547_ & ~new_n24548_;
  assign new_n24550_ = new_n24546_ & new_n24549_;
  assign new_n24551_ = new_n24541_ & new_n24550_;
  assign new_n24552_ = new_n24530_ & new_n24551_;
  assign new_n24553_ = new_n20072_ & new_n21096_;
  assign new_n24554_ = new_n20072_ & new_n21089_;
  assign new_n24555_ = new_n20072_ & new_n21085_;
  assign new_n24556_ = ~new_n24554_ & ~new_n24555_;
  assign new_n24557_ = ~new_n24553_ & new_n24556_;
  assign new_n24558_ = new_n20072_ & new_n21104_;
  assign new_n24559_ = new_n20072_ & new_n21098_;
  assign new_n24560_ = new_n20072_ & new_n21094_;
  assign new_n24561_ = ~new_n24559_ & ~new_n24560_;
  assign new_n24562_ = ~new_n24558_ & new_n24561_;
  assign new_n24563_ = new_n24557_ & new_n24562_;
  assign new_n24564_ = new_n20072_ & new_n21114_;
  assign new_n24565_ = new_n20072_ & new_n21106_;
  assign new_n24566_ = new_n20072_ & new_n21102_;
  assign new_n24567_ = ~new_n24565_ & ~new_n24566_;
  assign new_n24568_ = ~new_n24564_ & new_n24567_;
  assign new_n24569_ = new_n20120_ & new_n21017_;
  assign new_n24570_ = new_n20072_ & new_n21116_;
  assign new_n24571_ = new_n20072_ & new_n21112_;
  assign new_n24572_ = ~new_n24570_ & ~new_n24571_;
  assign new_n24573_ = ~new_n24569_ & new_n24572_;
  assign new_n24574_ = new_n24568_ & new_n24573_;
  assign new_n24575_ = new_n24563_ & new_n24574_;
  assign new_n24576_ = new_n20120_ & new_n21026_;
  assign new_n24577_ = new_n20120_ & new_n21019_;
  assign new_n24578_ = new_n20120_ & new_n21015_;
  assign new_n24579_ = ~new_n24577_ & ~new_n24578_;
  assign new_n24580_ = ~new_n24576_ & new_n24579_;
  assign new_n24581_ = new_n20120_ & new_n21039_;
  assign new_n24582_ = new_n20120_ & new_n21029_;
  assign new_n24583_ = new_n20120_ & new_n21024_;
  assign new_n24584_ = ~new_n24582_ & ~new_n24583_;
  assign new_n24585_ = ~new_n24581_ & new_n24584_;
  assign new_n24586_ = new_n24580_ & new_n24585_;
  assign new_n24587_ = new_n20120_ & new_n21050_;
  assign new_n24588_ = new_n20120_ & new_n21042_;
  assign new_n24589_ = new_n20120_ & new_n21036_;
  assign new_n24590_ = ~new_n24588_ & ~new_n24589_;
  assign new_n24591_ = ~new_n24587_ & new_n24590_;
  assign new_n24592_ = new_n20120_ & new_n21053_;
  assign new_n24593_ = new_n20120_ & new_n21047_;
  assign new_n24594_ = ~new_n24592_ & ~new_n24593_;
  assign new_n24595_ = new_n24591_ & new_n24594_;
  assign new_n24596_ = new_n24586_ & new_n24595_;
  assign new_n24597_ = new_n24575_ & new_n24596_;
  assign new_n24598_ = new_n24552_ & new_n24597_;
  assign new_n24599_ = new_n24507_ & new_n24598_;
  assign new_n24600_ = new_n20120_ & new_n21058_;
  assign new_n24601_ = new_n20120_ & new_n21060_;
  assign new_n24602_ = new_n20120_ & new_n21062_;
  assign new_n24603_ = ~new_n24601_ & ~new_n24602_;
  assign new_n24604_ = ~new_n24600_ & new_n24603_;
  assign new_n24605_ = new_n20120_ & new_n21079_;
  assign new_n24606_ = new_n20120_ & new_n21066_;
  assign new_n24607_ = new_n20120_ & new_n21068_;
  assign new_n24608_ = ~new_n24606_ & ~new_n24607_;
  assign new_n24609_ = ~new_n24605_ & new_n24608_;
  assign new_n24610_ = new_n24604_ & new_n24609_;
  assign new_n24611_ = new_n20120_ & new_n21087_;
  assign new_n24612_ = new_n20120_ & new_n21081_;
  assign new_n24613_ = new_n20120_ & new_n21077_;
  assign new_n24614_ = ~new_n24612_ & ~new_n24613_;
  assign new_n24615_ = ~new_n24611_ & new_n24614_;
  assign new_n24616_ = new_n20120_ & new_n21096_;
  assign new_n24617_ = new_n20120_ & new_n21089_;
  assign new_n24618_ = new_n20120_ & new_n21085_;
  assign new_n24619_ = ~new_n24617_ & ~new_n24618_;
  assign new_n24620_ = ~new_n24616_ & new_n24619_;
  assign new_n24621_ = new_n24615_ & new_n24620_;
  assign new_n24622_ = new_n24610_ & new_n24621_;
  assign new_n24623_ = new_n20120_ & new_n21104_;
  assign new_n24624_ = new_n20120_ & new_n21098_;
  assign new_n24625_ = new_n20120_ & new_n21094_;
  assign new_n24626_ = ~new_n24624_ & ~new_n24625_;
  assign new_n24627_ = ~new_n24623_ & new_n24626_;
  assign new_n24628_ = new_n20120_ & new_n21114_;
  assign new_n24629_ = new_n20120_ & new_n21106_;
  assign new_n24630_ = new_n20120_ & new_n21102_;
  assign new_n24631_ = ~new_n24629_ & ~new_n24630_;
  assign new_n24632_ = ~new_n24628_ & new_n24631_;
  assign new_n24633_ = new_n24627_ & new_n24632_;
  assign new_n24634_ = new_n20231_ & new_n21017_;
  assign new_n24635_ = new_n20120_ & new_n21116_;
  assign new_n24636_ = new_n20120_ & new_n21112_;
  assign new_n24637_ = ~new_n24635_ & ~new_n24636_;
  assign new_n24638_ = ~new_n24634_ & new_n24637_;
  assign new_n24639_ = new_n20231_ & new_n21019_;
  assign new_n24640_ = new_n20231_ & new_n21015_;
  assign new_n24641_ = ~new_n24639_ & ~new_n24640_;
  assign new_n24642_ = new_n24638_ & new_n24641_;
  assign new_n24643_ = new_n24633_ & new_n24642_;
  assign new_n24644_ = new_n24622_ & new_n24643_;
  assign new_n24645_ = new_n20231_ & new_n21024_;
  assign new_n24646_ = new_n20231_ & new_n21026_;
  assign new_n24647_ = new_n20231_ & new_n21029_;
  assign new_n24648_ = ~new_n24646_ & ~new_n24647_;
  assign new_n24649_ = ~new_n24645_ & new_n24648_;
  assign new_n24650_ = new_n20231_ & new_n21036_;
  assign new_n24651_ = new_n20231_ & new_n21039_;
  assign new_n24652_ = new_n20231_ & new_n21042_;
  assign new_n24653_ = ~new_n24651_ & ~new_n24652_;
  assign new_n24654_ = ~new_n24650_ & new_n24653_;
  assign new_n24655_ = new_n24649_ & new_n24654_;
  assign new_n24656_ = new_n20231_ & new_n21047_;
  assign new_n24657_ = new_n20231_ & new_n21050_;
  assign new_n24658_ = new_n20231_ & new_n21053_;
  assign new_n24659_ = ~new_n24657_ & ~new_n24658_;
  assign new_n24660_ = ~new_n24656_ & new_n24659_;
  assign new_n24661_ = new_n20231_ & new_n21058_;
  assign new_n24662_ = new_n20231_ & new_n21060_;
  assign new_n24663_ = new_n20231_ & new_n21062_;
  assign new_n24664_ = ~new_n24662_ & ~new_n24663_;
  assign new_n24665_ = ~new_n24661_ & new_n24664_;
  assign new_n24666_ = new_n24660_ & new_n24665_;
  assign new_n24667_ = new_n24655_ & new_n24666_;
  assign new_n24668_ = new_n20231_ & new_n21079_;
  assign new_n24669_ = new_n20231_ & new_n21066_;
  assign new_n24670_ = new_n20231_ & new_n21068_;
  assign new_n24671_ = ~new_n24669_ & ~new_n24670_;
  assign new_n24672_ = ~new_n24668_ & new_n24671_;
  assign new_n24673_ = new_n20231_ & new_n21087_;
  assign new_n24674_ = new_n20231_ & new_n21081_;
  assign new_n24675_ = new_n20231_ & new_n21077_;
  assign new_n24676_ = ~new_n24674_ & ~new_n24675_;
  assign new_n24677_ = ~new_n24673_ & new_n24676_;
  assign new_n24678_ = new_n24672_ & new_n24677_;
  assign new_n24679_ = new_n20231_ & new_n21096_;
  assign new_n24680_ = new_n20231_ & new_n21089_;
  assign new_n24681_ = new_n20231_ & new_n21085_;
  assign new_n24682_ = ~new_n24680_ & ~new_n24681_;
  assign new_n24683_ = ~new_n24679_ & new_n24682_;
  assign new_n24684_ = new_n20231_ & new_n21098_;
  assign new_n24685_ = new_n20231_ & new_n21094_;
  assign new_n24686_ = ~new_n24684_ & ~new_n24685_;
  assign new_n24687_ = new_n24683_ & new_n24686_;
  assign new_n24688_ = new_n24678_ & new_n24687_;
  assign new_n24689_ = new_n24667_ & new_n24688_;
  assign new_n24690_ = new_n24644_ & new_n24689_;
  assign new_n24691_ = new_n20231_ & new_n21102_;
  assign new_n24692_ = new_n20231_ & new_n21104_;
  assign new_n24693_ = new_n20231_ & new_n21106_;
  assign new_n24694_ = ~new_n24692_ & ~new_n24693_;
  assign new_n24695_ = ~new_n24691_ & new_n24694_;
  assign new_n24696_ = new_n20231_ & new_n21112_;
  assign new_n24697_ = new_n20231_ & new_n21114_;
  assign new_n24698_ = new_n20231_ & new_n21116_;
  assign new_n24699_ = ~new_n24697_ & ~new_n24698_;
  assign new_n24700_ = ~new_n24696_ & new_n24699_;
  assign new_n24701_ = new_n24695_ & new_n24700_;
  assign new_n24702_ = new_n20282_ & new_n21015_;
  assign new_n24703_ = new_n20282_ & new_n21017_;
  assign new_n24704_ = new_n20282_ & new_n21019_;
  assign new_n24705_ = ~new_n24703_ & ~new_n24704_;
  assign new_n24706_ = ~new_n24702_ & new_n24705_;
  assign new_n24707_ = new_n20282_ & new_n21024_;
  assign new_n24708_ = new_n20282_ & new_n21026_;
  assign new_n24709_ = new_n20282_ & new_n21029_;
  assign new_n24710_ = ~new_n24708_ & ~new_n24709_;
  assign new_n24711_ = ~new_n24707_ & new_n24710_;
  assign new_n24712_ = new_n24706_ & new_n24711_;
  assign new_n24713_ = new_n24701_ & new_n24712_;
  assign new_n24714_ = new_n20282_ & new_n21036_;
  assign new_n24715_ = new_n20282_ & new_n21039_;
  assign new_n24716_ = new_n20282_ & new_n21042_;
  assign new_n24717_ = ~new_n24715_ & ~new_n24716_;
  assign new_n24718_ = ~new_n24714_ & new_n24717_;
  assign new_n24719_ = new_n20282_ & new_n21047_;
  assign new_n24720_ = new_n20282_ & new_n21050_;
  assign new_n24721_ = new_n20282_ & new_n21053_;
  assign new_n24722_ = ~new_n24720_ & ~new_n24721_;
  assign new_n24723_ = ~new_n24719_ & new_n24722_;
  assign new_n24724_ = new_n24718_ & new_n24723_;
  assign new_n24725_ = new_n20282_ & new_n21058_;
  assign new_n24726_ = new_n20282_ & new_n21060_;
  assign new_n24727_ = new_n20282_ & new_n21062_;
  assign new_n24728_ = ~new_n24726_ & ~new_n24727_;
  assign new_n24729_ = ~new_n24725_ & new_n24728_;
  assign new_n24730_ = new_n20282_ & new_n21066_;
  assign new_n24731_ = new_n20282_ & new_n21068_;
  assign new_n24732_ = ~new_n24730_ & ~new_n24731_;
  assign new_n24733_ = new_n24729_ & new_n24732_;
  assign new_n24734_ = new_n24724_ & new_n24733_;
  assign new_n24735_ = new_n24713_ & new_n24734_;
  assign new_n24736_ = new_n20282_ & new_n21077_;
  assign new_n24737_ = new_n20282_ & new_n21079_;
  assign new_n24738_ = new_n20282_ & new_n21081_;
  assign new_n24739_ = ~new_n24737_ & ~new_n24738_;
  assign new_n24740_ = ~new_n24736_ & new_n24739_;
  assign new_n24741_ = new_n20282_ & new_n21085_;
  assign new_n24742_ = new_n20282_ & new_n21087_;
  assign new_n24743_ = new_n20282_ & new_n21089_;
  assign new_n24744_ = ~new_n24742_ & ~new_n24743_;
  assign new_n24745_ = ~new_n24741_ & new_n24744_;
  assign new_n24746_ = new_n24740_ & new_n24745_;
  assign new_n24747_ = new_n20282_ & new_n21094_;
  assign new_n24748_ = new_n20282_ & new_n21096_;
  assign new_n24749_ = new_n20282_ & new_n21098_;
  assign new_n24750_ = ~new_n24748_ & ~new_n24749_;
  assign new_n24751_ = ~new_n24747_ & new_n24750_;
  assign new_n24752_ = new_n20282_ & new_n21102_;
  assign new_n24753_ = new_n20282_ & new_n21104_;
  assign new_n24754_ = new_n20282_ & new_n21106_;
  assign new_n24755_ = ~new_n24753_ & ~new_n24754_;
  assign new_n24756_ = ~new_n24752_ & new_n24755_;
  assign new_n24757_ = new_n24751_ & new_n24756_;
  assign new_n24758_ = new_n24746_ & new_n24757_;
  assign new_n24759_ = new_n20282_ & new_n21112_;
  assign new_n24760_ = new_n20282_ & new_n21114_;
  assign new_n24761_ = new_n20282_ & new_n21116_;
  assign new_n24762_ = ~new_n24760_ & ~new_n24761_;
  assign new_n24763_ = ~new_n24759_ & new_n24762_;
  assign new_n24764_ = new_n20331_ & new_n21015_;
  assign new_n24765_ = new_n20331_ & new_n21017_;
  assign new_n24766_ = new_n20331_ & new_n21019_;
  assign new_n24767_ = ~new_n24765_ & ~new_n24766_;
  assign new_n24768_ = ~new_n24764_ & new_n24767_;
  assign new_n24769_ = new_n24763_ & new_n24768_;
  assign new_n24770_ = new_n20331_ & new_n21024_;
  assign new_n24771_ = new_n20331_ & new_n21026_;
  assign new_n24772_ = new_n20331_ & new_n21029_;
  assign new_n24773_ = ~new_n24771_ & ~new_n24772_;
  assign new_n24774_ = ~new_n24770_ & new_n24773_;
  assign new_n24775_ = new_n20331_ & new_n21039_;
  assign new_n24776_ = new_n20331_ & new_n21042_;
  assign new_n24777_ = ~new_n24775_ & ~new_n24776_;
  assign new_n24778_ = new_n24774_ & new_n24777_;
  assign new_n24779_ = new_n24769_ & new_n24778_;
  assign new_n24780_ = new_n24758_ & new_n24779_;
  assign new_n24781_ = new_n24735_ & new_n24780_;
  assign new_n24782_ = new_n24690_ & new_n24781_;
  assign new_n24783_ = new_n24599_ & new_n24782_;
  assign new_n24784_ = new_n20331_ & new_n21053_;
  assign new_n24785_ = new_n20331_ & new_n21036_;
  assign new_n24786_ = new_n20331_ & new_n21050_;
  assign new_n24787_ = ~new_n24785_ & ~new_n24786_;
  assign new_n24788_ = ~new_n24784_ & new_n24787_;
  assign new_n24789_ = new_n20331_ & new_n21062_;
  assign new_n24790_ = new_n20331_ & new_n21047_;
  assign new_n24791_ = new_n20331_ & new_n21060_;
  assign new_n24792_ = ~new_n24790_ & ~new_n24791_;
  assign new_n24793_ = ~new_n24789_ & new_n24792_;
  assign new_n24794_ = new_n24788_ & new_n24793_;
  assign new_n24795_ = new_n20331_ & new_n21068_;
  assign new_n24796_ = new_n20331_ & new_n21058_;
  assign new_n24797_ = new_n20331_ & new_n21066_;
  assign new_n24798_ = ~new_n24796_ & ~new_n24797_;
  assign new_n24799_ = ~new_n24795_ & new_n24798_;
  assign new_n24800_ = new_n20331_ & new_n21077_;
  assign new_n24801_ = new_n20331_ & new_n21079_;
  assign new_n24802_ = new_n20331_ & new_n21081_;
  assign new_n24803_ = ~new_n24801_ & ~new_n24802_;
  assign new_n24804_ = ~new_n24800_ & new_n24803_;
  assign new_n24805_ = new_n24799_ & new_n24804_;
  assign new_n24806_ = new_n24794_ & new_n24805_;
  assign new_n24807_ = new_n20331_ & new_n21085_;
  assign new_n24808_ = new_n20331_ & new_n21087_;
  assign new_n24809_ = new_n20331_ & new_n21089_;
  assign new_n24810_ = ~new_n24808_ & ~new_n24809_;
  assign new_n24811_ = ~new_n24807_ & new_n24810_;
  assign new_n24812_ = new_n20331_ & new_n21094_;
  assign new_n24813_ = new_n20331_ & new_n21096_;
  assign new_n24814_ = new_n20331_ & new_n21098_;
  assign new_n24815_ = ~new_n24813_ & ~new_n24814_;
  assign new_n24816_ = ~new_n24812_ & new_n24815_;
  assign new_n24817_ = new_n24811_ & new_n24816_;
  assign new_n24818_ = new_n20331_ & new_n21102_;
  assign new_n24819_ = new_n20331_ & new_n21104_;
  assign new_n24820_ = new_n20331_ & new_n21106_;
  assign new_n24821_ = ~new_n24819_ & ~new_n24820_;
  assign new_n24822_ = ~new_n24818_ & new_n24821_;
  assign new_n24823_ = new_n20331_ & new_n21114_;
  assign new_n24824_ = new_n20331_ & new_n21116_;
  assign new_n24825_ = ~new_n24823_ & ~new_n24824_;
  assign new_n24826_ = new_n24822_ & new_n24825_;
  assign new_n24827_ = new_n24817_ & new_n24826_;
  assign new_n24828_ = new_n24806_ & new_n24827_;
  assign new_n24829_ = new_n20377_ & new_n21019_;
  assign new_n24830_ = new_n20331_ & new_n21112_;
  assign new_n24831_ = new_n20377_ & new_n21017_;
  assign new_n24832_ = ~new_n24830_ & ~new_n24831_;
  assign new_n24833_ = ~new_n24829_ & new_n24832_;
  assign new_n24834_ = new_n20377_ & new_n21029_;
  assign new_n24835_ = new_n20377_ & new_n21015_;
  assign new_n24836_ = new_n20377_ & new_n21026_;
  assign new_n24837_ = ~new_n24835_ & ~new_n24836_;
  assign new_n24838_ = ~new_n24834_ & new_n24837_;
  assign new_n24839_ = new_n24833_ & new_n24838_;
  assign new_n24840_ = new_n20377_ & new_n21042_;
  assign new_n24841_ = new_n20377_ & new_n21024_;
  assign new_n24842_ = new_n20377_ & new_n21039_;
  assign new_n24843_ = ~new_n24841_ & ~new_n24842_;
  assign new_n24844_ = ~new_n24840_ & new_n24843_;
  assign new_n24845_ = new_n20377_ & new_n21053_;
  assign new_n24846_ = new_n20377_ & new_n21036_;
  assign new_n24847_ = new_n20377_ & new_n21050_;
  assign new_n24848_ = ~new_n24846_ & ~new_n24847_;
  assign new_n24849_ = ~new_n24845_ & new_n24848_;
  assign new_n24850_ = new_n24844_ & new_n24849_;
  assign new_n24851_ = new_n24839_ & new_n24850_;
  assign new_n24852_ = new_n20377_ & new_n21062_;
  assign new_n24853_ = new_n20377_ & new_n21047_;
  assign new_n24854_ = new_n20377_ & new_n21060_;
  assign new_n24855_ = ~new_n24853_ & ~new_n24854_;
  assign new_n24856_ = ~new_n24852_ & new_n24855_;
  assign new_n24857_ = new_n20377_ & new_n21068_;
  assign new_n24858_ = new_n20377_ & new_n21058_;
  assign new_n24859_ = new_n20377_ & new_n21066_;
  assign new_n24860_ = ~new_n24858_ & ~new_n24859_;
  assign new_n24861_ = ~new_n24857_ & new_n24860_;
  assign new_n24862_ = new_n24856_ & new_n24861_;
  assign new_n24863_ = new_n20377_ & new_n21077_;
  assign new_n24864_ = new_n20377_ & new_n21079_;
  assign new_n24865_ = new_n20377_ & new_n21081_;
  assign new_n24866_ = ~new_n24864_ & ~new_n24865_;
  assign new_n24867_ = ~new_n24863_ & new_n24866_;
  assign new_n24868_ = new_n20377_ & new_n21087_;
  assign new_n24869_ = new_n20377_ & new_n21089_;
  assign new_n24870_ = ~new_n24868_ & ~new_n24869_;
  assign new_n24871_ = new_n24867_ & new_n24870_;
  assign new_n24872_ = new_n24862_ & new_n24871_;
  assign new_n24873_ = new_n24851_ & new_n24872_;
  assign new_n24874_ = new_n24828_ & new_n24873_;
  assign new_n24875_ = new_n20377_ & new_n21098_;
  assign new_n24876_ = new_n20377_ & new_n21085_;
  assign new_n24877_ = new_n20377_ & new_n21096_;
  assign new_n24878_ = ~new_n24876_ & ~new_n24877_;
  assign new_n24879_ = ~new_n24875_ & new_n24878_;
  assign new_n24880_ = new_n20377_ & new_n21106_;
  assign new_n24881_ = new_n20377_ & new_n21094_;
  assign new_n24882_ = new_n20377_ & new_n21104_;
  assign new_n24883_ = ~new_n24881_ & ~new_n24882_;
  assign new_n24884_ = ~new_n24880_ & new_n24883_;
  assign new_n24885_ = new_n24879_ & new_n24884_;
  assign new_n24886_ = new_n20377_ & new_n21116_;
  assign new_n24887_ = new_n20377_ & new_n21102_;
  assign new_n24888_ = new_n20377_ & new_n21114_;
  assign new_n24889_ = ~new_n24887_ & ~new_n24888_;
  assign new_n24890_ = ~new_n24886_ & new_n24889_;
  assign new_n24891_ = new_n20494_ & new_n21019_;
  assign new_n24892_ = new_n20377_ & new_n21112_;
  assign new_n24893_ = new_n20494_ & new_n21017_;
  assign new_n24894_ = ~new_n24892_ & ~new_n24893_;
  assign new_n24895_ = ~new_n24891_ & new_n24894_;
  assign new_n24896_ = new_n24890_ & new_n24895_;
  assign new_n24897_ = new_n24885_ & new_n24896_;
  assign new_n24898_ = new_n20494_ & new_n21029_;
  assign new_n24899_ = new_n20494_ & new_n21015_;
  assign new_n24900_ = new_n20494_ & new_n21026_;
  assign new_n24901_ = ~new_n24899_ & ~new_n24900_;
  assign new_n24902_ = ~new_n24898_ & new_n24901_;
  assign new_n24903_ = new_n20494_ & new_n21042_;
  assign new_n24904_ = new_n20494_ & new_n21024_;
  assign new_n24905_ = new_n20494_ & new_n21039_;
  assign new_n24906_ = ~new_n24904_ & ~new_n24905_;
  assign new_n24907_ = ~new_n24903_ & new_n24906_;
  assign new_n24908_ = new_n24902_ & new_n24907_;
  assign new_n24909_ = new_n20494_ & new_n21053_;
  assign new_n24910_ = new_n20494_ & new_n21036_;
  assign new_n24911_ = new_n20494_ & new_n21050_;
  assign new_n24912_ = ~new_n24910_ & ~new_n24911_;
  assign new_n24913_ = ~new_n24909_ & new_n24912_;
  assign new_n24914_ = new_n20494_ & new_n21047_;
  assign new_n24915_ = new_n20494_ & new_n21060_;
  assign new_n24916_ = ~new_n24914_ & ~new_n24915_;
  assign new_n24917_ = new_n24913_ & new_n24916_;
  assign new_n24918_ = new_n24908_ & new_n24917_;
  assign new_n24919_ = new_n24897_ & new_n24918_;
  assign new_n24920_ = new_n20494_ & new_n21066_;
  assign new_n24921_ = new_n20494_ & new_n21062_;
  assign new_n24922_ = new_n20494_ & new_n21058_;
  assign new_n24923_ = ~new_n24921_ & ~new_n24922_;
  assign new_n24924_ = ~new_n24920_ & new_n24923_;
  assign new_n24925_ = new_n20494_ & new_n21081_;
  assign new_n24926_ = new_n20494_ & new_n21068_;
  assign new_n24927_ = new_n20494_ & new_n21079_;
  assign new_n24928_ = ~new_n24926_ & ~new_n24927_;
  assign new_n24929_ = ~new_n24925_ & new_n24928_;
  assign new_n24930_ = new_n24924_ & new_n24929_;
  assign new_n24931_ = new_n20494_ & new_n21089_;
  assign new_n24932_ = new_n20494_ & new_n21077_;
  assign new_n24933_ = new_n20494_ & new_n21087_;
  assign new_n24934_ = ~new_n24932_ & ~new_n24933_;
  assign new_n24935_ = ~new_n24931_ & new_n24934_;
  assign new_n24936_ = new_n20494_ & new_n21098_;
  assign new_n24937_ = new_n20494_ & new_n21085_;
  assign new_n24938_ = new_n20494_ & new_n21096_;
  assign new_n24939_ = ~new_n24937_ & ~new_n24938_;
  assign new_n24940_ = ~new_n24936_ & new_n24939_;
  assign new_n24941_ = new_n24935_ & new_n24940_;
  assign new_n24942_ = new_n24930_ & new_n24941_;
  assign new_n24943_ = new_n20494_ & new_n21106_;
  assign new_n24944_ = new_n20494_ & new_n21094_;
  assign new_n24945_ = new_n20494_ & new_n21104_;
  assign new_n24946_ = ~new_n24944_ & ~new_n24945_;
  assign new_n24947_ = ~new_n24943_ & new_n24946_;
  assign new_n24948_ = new_n20494_ & new_n21116_;
  assign new_n24949_ = new_n20494_ & new_n21102_;
  assign new_n24950_ = new_n20494_ & new_n21114_;
  assign new_n24951_ = ~new_n24949_ & ~new_n24950_;
  assign new_n24952_ = ~new_n24948_ & new_n24951_;
  assign new_n24953_ = new_n24947_ & new_n24952_;
  assign new_n24954_ = new_n20540_ & new_n21019_;
  assign new_n24955_ = new_n20494_ & new_n21112_;
  assign new_n24956_ = new_n20540_ & new_n21017_;
  assign new_n24957_ = ~new_n24955_ & ~new_n24956_;
  assign new_n24958_ = ~new_n24954_ & new_n24957_;
  assign new_n24959_ = new_n20540_ & new_n21015_;
  assign new_n24960_ = new_n20540_ & new_n21026_;
  assign new_n24961_ = ~new_n24959_ & ~new_n24960_;
  assign new_n24962_ = new_n24958_ & new_n24961_;
  assign new_n24963_ = new_n24953_ & new_n24962_;
  assign new_n24964_ = new_n24942_ & new_n24963_;
  assign new_n24965_ = new_n24919_ & new_n24964_;
  assign new_n24966_ = new_n24874_ & new_n24965_;
  assign new_n24967_ = new_n20540_ & new_n21039_;
  assign new_n24968_ = new_n20540_ & new_n21029_;
  assign new_n24969_ = new_n20540_ & new_n21024_;
  assign new_n24970_ = ~new_n24968_ & ~new_n24969_;
  assign new_n24971_ = ~new_n24967_ & new_n24970_;
  assign new_n24972_ = new_n20540_ & new_n21050_;
  assign new_n24973_ = new_n20540_ & new_n21042_;
  assign new_n24974_ = new_n20540_ & new_n21036_;
  assign new_n24975_ = ~new_n24973_ & ~new_n24974_;
  assign new_n24976_ = ~new_n24972_ & new_n24975_;
  assign new_n24977_ = new_n24971_ & new_n24976_;
  assign new_n24978_ = new_n20540_ & new_n21060_;
  assign new_n24979_ = new_n20540_ & new_n21053_;
  assign new_n24980_ = new_n20540_ & new_n21047_;
  assign new_n24981_ = ~new_n24979_ & ~new_n24980_;
  assign new_n24982_ = ~new_n24978_ & new_n24981_;
  assign new_n24983_ = new_n20540_ & new_n21066_;
  assign new_n24984_ = new_n20540_ & new_n21062_;
  assign new_n24985_ = new_n20540_ & new_n21058_;
  assign new_n24986_ = ~new_n24984_ & ~new_n24985_;
  assign new_n24987_ = ~new_n24983_ & new_n24986_;
  assign new_n24988_ = new_n24982_ & new_n24987_;
  assign new_n24989_ = new_n24977_ & new_n24988_;
  assign new_n24990_ = new_n20540_ & new_n21081_;
  assign new_n24991_ = new_n20540_ & new_n21068_;
  assign new_n24992_ = new_n20540_ & new_n21079_;
  assign new_n24993_ = ~new_n24991_ & ~new_n24992_;
  assign new_n24994_ = ~new_n24990_ & new_n24993_;
  assign new_n24995_ = new_n20540_ & new_n21089_;
  assign new_n24996_ = new_n20540_ & new_n21077_;
  assign new_n24997_ = new_n20540_ & new_n21087_;
  assign new_n24998_ = ~new_n24996_ & ~new_n24997_;
  assign new_n24999_ = ~new_n24995_ & new_n24998_;
  assign new_n25000_ = new_n24994_ & new_n24999_;
  assign new_n25001_ = new_n20540_ & new_n21098_;
  assign new_n25002_ = new_n20540_ & new_n21085_;
  assign new_n25003_ = new_n20540_ & new_n21096_;
  assign new_n25004_ = ~new_n25002_ & ~new_n25003_;
  assign new_n25005_ = ~new_n25001_ & new_n25004_;
  assign new_n25006_ = new_n20540_ & new_n21094_;
  assign new_n25007_ = new_n20540_ & new_n21104_;
  assign new_n25008_ = ~new_n25006_ & ~new_n25007_;
  assign new_n25009_ = new_n25005_ & new_n25008_;
  assign new_n25010_ = new_n25000_ & new_n25009_;
  assign new_n25011_ = new_n24989_ & new_n25010_;
  assign new_n25012_ = new_n20540_ & new_n21114_;
  assign new_n25013_ = new_n20540_ & new_n21106_;
  assign new_n25014_ = new_n20540_ & new_n21102_;
  assign new_n25015_ = ~new_n25013_ & ~new_n25014_;
  assign new_n25016_ = ~new_n25012_ & new_n25015_;
  assign new_n25017_ = new_n20593_ & new_n21017_;
  assign new_n25018_ = new_n20540_ & new_n21116_;
  assign new_n25019_ = new_n20540_ & new_n21112_;
  assign new_n25020_ = ~new_n25018_ & ~new_n25019_;
  assign new_n25021_ = ~new_n25017_ & new_n25020_;
  assign new_n25022_ = new_n25016_ & new_n25021_;
  assign new_n25023_ = new_n20593_ & new_n21026_;
  assign new_n25024_ = new_n20593_ & new_n21019_;
  assign new_n25025_ = new_n20593_ & new_n21015_;
  assign new_n25026_ = ~new_n25024_ & ~new_n25025_;
  assign new_n25027_ = ~new_n25023_ & new_n25026_;
  assign new_n25028_ = new_n20593_ & new_n21039_;
  assign new_n25029_ = new_n20593_ & new_n21029_;
  assign new_n25030_ = new_n20593_ & new_n21024_;
  assign new_n25031_ = ~new_n25029_ & ~new_n25030_;
  assign new_n25032_ = ~new_n25028_ & new_n25031_;
  assign new_n25033_ = new_n25027_ & new_n25032_;
  assign new_n25034_ = new_n25022_ & new_n25033_;
  assign new_n25035_ = new_n20593_ & new_n21050_;
  assign new_n25036_ = new_n20593_ & new_n21042_;
  assign new_n25037_ = new_n20593_ & new_n21036_;
  assign new_n25038_ = ~new_n25036_ & ~new_n25037_;
  assign new_n25039_ = ~new_n25035_ & new_n25038_;
  assign new_n25040_ = new_n20593_ & new_n21060_;
  assign new_n25041_ = new_n20593_ & new_n21053_;
  assign new_n25042_ = new_n20593_ & new_n21047_;
  assign new_n25043_ = ~new_n25041_ & ~new_n25042_;
  assign new_n25044_ = ~new_n25040_ & new_n25043_;
  assign new_n25045_ = new_n25039_ & new_n25044_;
  assign new_n25046_ = new_n20593_ & new_n21066_;
  assign new_n25047_ = new_n20593_ & new_n21062_;
  assign new_n25048_ = new_n20593_ & new_n21058_;
  assign new_n25049_ = ~new_n25047_ & ~new_n25048_;
  assign new_n25050_ = ~new_n25046_ & new_n25049_;
  assign new_n25051_ = new_n20593_ & new_n21068_;
  assign new_n25052_ = new_n20593_ & new_n21079_;
  assign new_n25053_ = ~new_n25051_ & ~new_n25052_;
  assign new_n25054_ = new_n25050_ & new_n25053_;
  assign new_n25055_ = new_n25045_ & new_n25054_;
  assign new_n25056_ = new_n25034_ & new_n25055_;
  assign new_n25057_ = new_n25011_ & new_n25056_;
  assign new_n25058_ = new_n20593_ & new_n21087_;
  assign new_n25059_ = new_n20593_ & new_n21081_;
  assign new_n25060_ = new_n20593_ & new_n21077_;
  assign new_n25061_ = ~new_n25059_ & ~new_n25060_;
  assign new_n25062_ = ~new_n25058_ & new_n25061_;
  assign new_n25063_ = new_n20593_ & new_n21096_;
  assign new_n25064_ = new_n20593_ & new_n21089_;
  assign new_n25065_ = new_n20593_ & new_n21085_;
  assign new_n25066_ = ~new_n25064_ & ~new_n25065_;
  assign new_n25067_ = ~new_n25063_ & new_n25066_;
  assign new_n25068_ = new_n25062_ & new_n25067_;
  assign new_n25069_ = new_n20593_ & new_n21104_;
  assign new_n25070_ = new_n20593_ & new_n21098_;
  assign new_n25071_ = new_n20593_ & new_n21094_;
  assign new_n25072_ = ~new_n25070_ & ~new_n25071_;
  assign new_n25073_ = ~new_n25069_ & new_n25072_;
  assign new_n25074_ = new_n20593_ & new_n21114_;
  assign new_n25075_ = new_n20593_ & new_n21106_;
  assign new_n25076_ = new_n20593_ & new_n21102_;
  assign new_n25077_ = ~new_n25075_ & ~new_n25076_;
  assign new_n25078_ = ~new_n25074_ & new_n25077_;
  assign new_n25079_ = new_n25073_ & new_n25078_;
  assign new_n25080_ = new_n25068_ & new_n25079_;
  assign new_n25081_ = new_n20639_ & new_n21017_;
  assign new_n25082_ = new_n20593_ & new_n21116_;
  assign new_n25083_ = new_n20593_ & new_n21112_;
  assign new_n25084_ = ~new_n25082_ & ~new_n25083_;
  assign new_n25085_ = ~new_n25081_ & new_n25084_;
  assign new_n25086_ = new_n20639_ & new_n21026_;
  assign new_n25087_ = new_n20639_ & new_n21019_;
  assign new_n25088_ = new_n20639_ & new_n21015_;
  assign new_n25089_ = ~new_n25087_ & ~new_n25088_;
  assign new_n25090_ = ~new_n25086_ & new_n25089_;
  assign new_n25091_ = new_n25085_ & new_n25090_;
  assign new_n25092_ = new_n20639_ & new_n21039_;
  assign new_n25093_ = new_n20639_ & new_n21029_;
  assign new_n25094_ = new_n20639_ & new_n21024_;
  assign new_n25095_ = ~new_n25093_ & ~new_n25094_;
  assign new_n25096_ = ~new_n25092_ & new_n25095_;
  assign new_n25097_ = new_n20639_ & new_n21042_;
  assign new_n25098_ = new_n20639_ & new_n21036_;
  assign new_n25099_ = ~new_n25097_ & ~new_n25098_;
  assign new_n25100_ = new_n25096_ & new_n25099_;
  assign new_n25101_ = new_n25091_ & new_n25100_;
  assign new_n25102_ = new_n25080_ & new_n25101_;
  assign new_n25103_ = new_n20639_ & new_n21047_;
  assign new_n25104_ = new_n20639_ & new_n21050_;
  assign new_n25105_ = new_n20639_ & new_n21053_;
  assign new_n25106_ = ~new_n25104_ & ~new_n25105_;
  assign new_n25107_ = ~new_n25103_ & new_n25106_;
  assign new_n25108_ = new_n20639_ & new_n21058_;
  assign new_n25109_ = new_n20639_ & new_n21060_;
  assign new_n25110_ = new_n20639_ & new_n21062_;
  assign new_n25111_ = ~new_n25109_ & ~new_n25110_;
  assign new_n25112_ = ~new_n25108_ & new_n25111_;
  assign new_n25113_ = new_n25107_ & new_n25112_;
  assign new_n25114_ = new_n20639_ & new_n21079_;
  assign new_n25115_ = new_n20639_ & new_n21066_;
  assign new_n25116_ = new_n20639_ & new_n21068_;
  assign new_n25117_ = ~new_n25115_ & ~new_n25116_;
  assign new_n25118_ = ~new_n25114_ & new_n25117_;
  assign new_n25119_ = new_n20639_ & new_n21087_;
  assign new_n25120_ = new_n20639_ & new_n21081_;
  assign new_n25121_ = new_n20639_ & new_n21077_;
  assign new_n25122_ = ~new_n25120_ & ~new_n25121_;
  assign new_n25123_ = ~new_n25119_ & new_n25122_;
  assign new_n25124_ = new_n25118_ & new_n25123_;
  assign new_n25125_ = new_n25113_ & new_n25124_;
  assign new_n25126_ = new_n20639_ & new_n21096_;
  assign new_n25127_ = new_n20639_ & new_n21089_;
  assign new_n25128_ = new_n20639_ & new_n21085_;
  assign new_n25129_ = ~new_n25127_ & ~new_n25128_;
  assign new_n25130_ = ~new_n25126_ & new_n25129_;
  assign new_n25131_ = new_n20639_ & new_n21104_;
  assign new_n25132_ = new_n20639_ & new_n21098_;
  assign new_n25133_ = new_n20639_ & new_n21094_;
  assign new_n25134_ = ~new_n25132_ & ~new_n25133_;
  assign new_n25135_ = ~new_n25131_ & new_n25134_;
  assign new_n25136_ = new_n25130_ & new_n25135_;
  assign new_n25137_ = new_n20639_ & new_n21114_;
  assign new_n25138_ = new_n20639_ & new_n21106_;
  assign new_n25139_ = new_n20639_ & new_n21102_;
  assign new_n25140_ = ~new_n25138_ & ~new_n25139_;
  assign new_n25141_ = ~new_n25137_ & new_n25140_;
  assign new_n25142_ = new_n20639_ & new_n21116_;
  assign new_n25143_ = new_n20639_ & new_n21112_;
  assign new_n25144_ = ~new_n25142_ & ~new_n25143_;
  assign new_n25145_ = new_n25141_ & new_n25144_;
  assign new_n25146_ = new_n25136_ & new_n25145_;
  assign new_n25147_ = new_n25125_ & new_n25146_;
  assign new_n25148_ = new_n25102_ & new_n25147_;
  assign new_n25149_ = new_n25057_ & new_n25148_;
  assign new_n25150_ = new_n24966_ & new_n25149_;
  assign new_n25151_ = new_n24783_ & new_n25150_;
  assign new_n25152_ = new_n24414_ & new_n25151_;
  assign new_n25153_ = new_n23677_ & new_n25152_;
  assign new_n25154_ = new_n22200_ & new_n25153_;
  assign new_n25155_ = new_n19174_ & new_n25154_;
  assign A10 = ~new_n13117_ | ~new_n25155_;
endmodule


