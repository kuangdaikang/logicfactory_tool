// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:34 2022

module amd  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13,
    \v14.0 , \v14.1 , \v14.2 , \v14.3 , \v14.4 , \v14.5 , \v14.6 , \v14.7 ,
    \v14.8 , \v14.9 , \v14.10 , \v14.11 , \v14.12 , \v14.13 , \v14.14 ,
    \v14.15 , \v14.16 , \v14.17 , \v14.18 , \v14.19 , \v14.20 , \v14.21 ,
    \v14.22 , \v14.23   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13;
  output \v14.0 , \v14.1 , \v14.2 , \v14.3 , \v14.4 , \v14.5 , \v14.6 ,
    \v14.7 , \v14.8 , \v14.9 , \v14.10 , \v14.11 , \v14.12 , \v14.13 ,
    \v14.14 , \v14.15 , \v14.16 , \v14.17 , \v14.18 , \v14.19 , \v14.20 ,
    \v14.21 , \v14.22 , \v14.23 ;
  wire new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_,
    new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n337_, new_n338_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n414_, new_n415_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n579_, new_n580_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_;
  assign new_n39_ = v0 & ~v4;
  assign new_n40_ = v0 & ~new_n39_;
  assign new_n41_ = ~v12 & ~new_n40_;
  assign new_n42_ = ~v0 & v12;
  assign new_n43_ = ~new_n41_ & ~new_n42_;
  assign new_n44_ = ~v5 & ~new_n43_;
  assign new_n45_ = ~v3 & v5;
  assign new_n46_ = ~new_n44_ & ~new_n45_;
  assign new_n47_ = v13 & ~new_n46_;
  assign new_n48_ = v12 & ~v13;
  assign new_n49_ = new_n45_ & new_n48_;
  assign new_n50_ = ~new_n47_ & ~new_n49_;
  assign new_n51_ = ~v4 & ~v11;
  assign new_n52_ = v12 & v13;
  assign new_n53_ = new_n51_ & new_n52_;
  assign new_n54_ = ~v12 & ~v13;
  assign new_n55_ = v11 & new_n54_;
  assign new_n56_ = ~new_n53_ & ~new_n55_;
  assign new_n57_ = ~v5 & ~new_n56_;
  assign new_n58_ = v0 & new_n57_;
  assign new_n59_ = new_n45_ & new_n55_;
  assign new_n60_ = ~new_n58_ & ~new_n59_;
  assign new_n61_ = new_n50_ & new_n60_;
  assign new_n62_ = ~v10 & ~new_n61_;
  assign new_n63_ = ~v12 & v13;
  assign new_n64_ = ~v0 & new_n63_;
  assign new_n65_ = v0 & new_n48_;
  assign new_n66_ = ~new_n64_ & ~new_n65_;
  assign new_n67_ = ~v5 & ~new_n66_;
  assign new_n68_ = v12 & ~new_n48_;
  assign new_n69_ = v5 & ~new_n68_;
  assign new_n70_ = ~v3 & new_n69_;
  assign new_n71_ = ~new_n67_ & ~new_n70_;
  assign new_n72_ = ~v11 & ~new_n71_;
  assign new_n73_ = ~v1 & ~v3;
  assign new_n74_ = ~v1 & ~new_n73_;
  assign new_n75_ = v13 & ~new_n74_;
  assign new_n76_ = v12 & new_n75_;
  assign new_n77_ = v11 & new_n76_;
  assign new_n78_ = ~new_n72_ & ~new_n77_;
  assign new_n79_ = v10 & ~new_n78_;
  assign new_n80_ = ~new_n62_ & ~new_n79_;
  assign new_n81_ = ~v9 & ~new_n80_;
  assign new_n82_ = v4 & v12;
  assign new_n83_ = ~v0 & new_n82_;
  assign new_n84_ = ~new_n39_ & ~new_n83_;
  assign new_n85_ = ~v5 & ~new_n84_;
  assign new_n86_ = ~new_n45_ & ~new_n85_;
  assign new_n87_ = ~v13 & ~new_n86_;
  assign new_n88_ = ~v11 & new_n87_;
  assign new_n89_ = ~v10 & new_n88_;
  assign new_n90_ = v9 & new_n89_;
  assign new_n91_ = ~new_n81_ & ~new_n90_;
  assign new_n92_ = ~v5 & v12;
  assign new_n93_ = v4 & new_n92_;
  assign new_n94_ = ~new_n45_ & ~new_n93_;
  assign new_n95_ = ~v10 & ~new_n94_;
  assign new_n96_ = v9 & new_n95_;
  assign new_n97_ = v10 & v12;
  assign new_n98_ = ~v9 & new_n97_;
  assign new_n99_ = ~new_n96_ & ~new_n98_;
  assign new_n100_ = ~v11 & ~new_n99_;
  assign new_n101_ = ~v9 & v10;
  assign new_n102_ = v11 & ~v12;
  assign new_n103_ = new_n101_ & new_n102_;
  assign new_n104_ = ~new_n100_ & ~new_n103_;
  assign new_n105_ = v13 & ~new_n104_;
  assign new_n106_ = new_n91_ & ~new_n105_;
  assign new_n107_ = v6 & ~new_n106_;
  assign new_n108_ = v10 & v11;
  assign new_n109_ = ~v6 & new_n108_;
  assign new_n110_ = ~v10 & ~v11;
  assign new_n111_ = v3 & new_n110_;
  assign new_n112_ = ~new_n109_ & ~new_n111_;
  assign new_n113_ = ~v9 & ~new_n112_;
  assign new_n114_ = v8 & new_n113_;
  assign new_n115_ = ~v10 & v11;
  assign new_n116_ = v9 & new_n115_;
  assign new_n117_ = ~new_n114_ & ~new_n116_;
  assign new_n118_ = ~v13 & ~new_n117_;
  assign new_n119_ = ~v6 & v9;
  assign new_n120_ = ~v11 & v13;
  assign new_n121_ = ~v10 & new_n120_;
  assign new_n122_ = new_n119_ & new_n121_;
  assign new_n123_ = ~new_n118_ & ~new_n122_;
  assign new_n124_ = ~v12 & ~new_n123_;
  assign new_n125_ = v9 & ~v10;
  assign new_n126_ = ~v6 & new_n125_;
  assign new_n127_ = ~v11 & new_n52_;
  assign new_n128_ = new_n126_ & new_n127_;
  assign new_n129_ = ~new_n124_ & ~new_n128_;
  assign new_n130_ = ~v5 & ~new_n129_;
  assign \v14.0  = new_n107_ | new_n130_;
  assign new_n132_ = ~v9 & new_n63_;
  assign new_n133_ = v9 & new_n48_;
  assign new_n134_ = ~new_n132_ & ~new_n133_;
  assign new_n135_ = v4 & ~v5;
  assign new_n136_ = v0 & new_n135_;
  assign new_n137_ = ~v5 & ~new_n136_;
  assign new_n138_ = ~new_n134_ & ~new_n137_;
  assign new_n139_ = v0 & ~v12;
  assign new_n140_ = ~new_n42_ & ~new_n139_;
  assign new_n141_ = ~v5 & ~new_n140_;
  assign new_n142_ = v5 & ~v12;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = v9 & ~new_n143_;
  assign new_n145_ = ~v0 & ~v5;
  assign new_n146_ = ~v5 & ~new_n145_;
  assign new_n147_ = v12 & ~new_n146_;
  assign new_n148_ = ~v9 & new_n147_;
  assign new_n149_ = ~new_n144_ & ~new_n148_;
  assign new_n150_ = ~v13 & ~new_n149_;
  assign new_n151_ = v0 & v4;
  assign new_n152_ = v0 & ~new_n151_;
  assign new_n153_ = ~v5 & ~new_n152_;
  assign new_n154_ = ~v5 & ~new_n153_;
  assign new_n155_ = v13 & ~new_n154_;
  assign new_n156_ = v12 & new_n155_;
  assign new_n157_ = ~v9 & new_n156_;
  assign new_n158_ = ~new_n150_ & ~new_n157_;
  assign new_n159_ = ~new_n138_ & new_n158_;
  assign new_n160_ = ~v10 & ~new_n159_;
  assign new_n161_ = v0 & ~v5;
  assign new_n162_ = ~v5 & ~new_n161_;
  assign new_n163_ = ~v0 & new_n92_;
  assign new_n164_ = new_n162_ & ~new_n163_;
  assign new_n165_ = ~v13 & ~new_n164_;
  assign new_n166_ = v5 & new_n63_;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = v10 & ~new_n167_;
  assign new_n169_ = ~v9 & new_n168_;
  assign new_n170_ = ~new_n160_ & ~new_n169_;
  assign new_n171_ = ~v11 & ~new_n170_;
  assign new_n172_ = ~v12 & ~new_n137_;
  assign new_n173_ = ~new_n147_ & ~new_n172_;
  assign new_n174_ = v13 & ~new_n173_;
  assign new_n175_ = ~v5 & ~new_n163_;
  assign new_n176_ = ~v13 & ~new_n175_;
  assign new_n177_ = ~new_n174_ & ~new_n176_;
  assign new_n178_ = ~v10 & ~new_n177_;
  assign new_n179_ = ~v1 & new_n97_;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = v11 & ~new_n180_;
  assign new_n182_ = ~v9 & new_n181_;
  assign new_n183_ = ~new_n171_ & ~new_n182_;
  assign new_n184_ = ~v5 & ~new_n92_;
  assign new_n185_ = ~v10 & ~new_n184_;
  assign new_n186_ = v9 & new_n185_;
  assign new_n187_ = ~new_n98_ & ~new_n186_;
  assign new_n188_ = v13 & ~new_n187_;
  assign new_n189_ = ~v11 & new_n188_;
  assign new_n190_ = new_n183_ & ~new_n189_;
  assign new_n191_ = v6 & ~new_n190_;
  assign new_n192_ = ~v6 & ~v11;
  assign new_n193_ = new_n52_ & new_n192_;
  assign new_n194_ = ~new_n55_ & ~new_n193_;
  assign new_n195_ = ~v10 & ~new_n194_;
  assign new_n196_ = v9 & new_n195_;
  assign new_n197_ = ~v5 & new_n196_;
  assign \v14.1  = new_n191_ | new_n197_;
  assign new_n199_ = ~v13 & ~new_n112_;
  assign new_n200_ = ~v8 & new_n199_;
  assign new_n201_ = ~v10 & v13;
  assign new_n202_ = v6 & new_n201_;
  assign new_n203_ = v0 & new_n202_;
  assign new_n204_ = ~new_n200_ & ~new_n203_;
  assign new_n205_ = ~v4 & ~new_n204_;
  assign new_n206_ = v13 & ~new_n152_;
  assign new_n207_ = ~v0 & ~v13;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = v11 & ~new_n208_;
  assign new_n210_ = v4 & new_n120_;
  assign new_n211_ = v0 & new_n210_;
  assign new_n212_ = ~new_n209_ & ~new_n211_;
  assign new_n213_ = ~v10 & ~new_n212_;
  assign new_n214_ = v6 & new_n213_;
  assign new_n215_ = ~new_n205_ & ~new_n214_;
  assign new_n216_ = ~v5 & ~new_n215_;
  assign new_n217_ = v10 & ~v11;
  assign new_n218_ = ~new_n115_ & ~new_n217_;
  assign new_n219_ = ~new_n121_ & new_n218_;
  assign new_n220_ = v5 & ~new_n219_;
  assign new_n221_ = ~new_n108_ & ~new_n220_;
  assign new_n222_ = v6 & ~new_n221_;
  assign new_n223_ = ~new_n216_ & ~new_n222_;
  assign new_n224_ = ~v12 & ~new_n223_;
  assign new_n225_ = v5 & ~v11;
  assign new_n226_ = ~v11 & ~new_n225_;
  assign new_n227_ = ~v10 & ~new_n226_;
  assign new_n228_ = v1 & new_n108_;
  assign new_n229_ = ~new_n227_ & ~new_n228_;
  assign new_n230_ = v4 & v13;
  assign new_n231_ = v13 & ~new_n230_;
  assign new_n232_ = ~v10 & ~new_n231_;
  assign new_n233_ = ~v5 & new_n232_;
  assign new_n234_ = v0 & new_n233_;
  assign new_n235_ = v10 & ~v13;
  assign new_n236_ = v5 & new_n235_;
  assign new_n237_ = ~new_n234_ & ~new_n236_;
  assign new_n238_ = ~v11 & ~new_n237_;
  assign new_n239_ = ~v1 & new_n108_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = new_n229_ & new_n240_;
  assign new_n242_ = v12 & ~new_n241_;
  assign new_n243_ = v6 & new_n242_;
  assign new_n244_ = ~new_n224_ & ~new_n243_;
  assign new_n245_ = ~v9 & ~new_n244_;
  assign new_n246_ = ~v0 & v4;
  assign new_n247_ = ~v0 & ~new_n246_;
  assign new_n248_ = ~v5 & ~new_n247_;
  assign new_n249_ = ~v5 & ~new_n248_;
  assign new_n250_ = v12 & ~new_n249_;
  assign new_n251_ = ~new_n142_ & ~new_n250_;
  assign new_n252_ = ~v13 & ~new_n251_;
  assign new_n253_ = ~v5 & ~new_n93_;
  assign new_n254_ = v13 & ~new_n253_;
  assign new_n255_ = ~new_n252_ & ~new_n254_;
  assign new_n256_ = ~v11 & ~new_n255_;
  assign new_n257_ = ~v10 & new_n256_;
  assign new_n258_ = v9 & new_n257_;
  assign new_n259_ = v6 & new_n258_;
  assign \v14.2  = new_n245_ | new_n259_;
  assign new_n261_ = ~v10 & v12;
  assign new_n262_ = v10 & ~v12;
  assign new_n263_ = ~new_n261_ & ~new_n262_;
  assign new_n264_ = v5 & ~new_n263_;
  assign new_n265_ = ~v5 & new_n262_;
  assign new_n266_ = ~new_n264_ & ~new_n265_;
  assign new_n267_ = ~v11 & ~new_n266_;
  assign new_n268_ = v5 & ~v10;
  assign new_n269_ = v1 & new_n97_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = v11 & ~new_n270_;
  assign new_n272_ = ~new_n267_ & ~new_n271_;
  assign new_n273_ = v10 & new_n102_;
  assign new_n274_ = new_n272_ & ~new_n273_;
  assign new_n275_ = ~v11 & v12;
  assign new_n276_ = v10 & new_n275_;
  assign new_n277_ = ~v10 & new_n102_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = v0 & ~new_n278_;
  assign new_n280_ = ~v0 & v10;
  assign new_n281_ = new_n275_ & new_n280_;
  assign new_n282_ = ~new_n279_ & ~new_n281_;
  assign new_n283_ = ~v5 & ~new_n282_;
  assign new_n284_ = ~v1 & v11;
  assign new_n285_ = ~new_n225_ & ~new_n284_;
  assign new_n286_ = v12 & ~new_n285_;
  assign new_n287_ = v10 & new_n286_;
  assign new_n288_ = ~new_n283_ & ~new_n287_;
  assign new_n289_ = ~v13 & ~new_n288_;
  assign new_n290_ = ~v1 & v10;
  assign new_n291_ = v11 & v12;
  assign new_n292_ = new_n290_ & new_n291_;
  assign new_n293_ = ~v11 & ~v12;
  assign new_n294_ = new_n268_ & new_n293_;
  assign new_n295_ = ~new_n292_ & ~new_n294_;
  assign new_n296_ = v13 & ~new_n295_;
  assign new_n297_ = ~new_n289_ & ~new_n296_;
  assign new_n298_ = new_n52_ & new_n217_;
  assign new_n299_ = new_n297_ & ~new_n298_;
  assign new_n300_ = new_n274_ & new_n299_;
  assign new_n301_ = ~v9 & ~new_n300_;
  assign new_n302_ = v9 & new_n110_;
  assign new_n303_ = v5 & new_n302_;
  assign new_n304_ = ~new_n301_ & ~new_n303_;
  assign \v14.3  = v6 & ~new_n304_;
  assign new_n306_ = v9 & v11;
  assign new_n307_ = v6 & v9;
  assign new_n308_ = ~v0 & new_n307_;
  assign new_n309_ = v4 & v8;
  assign new_n310_ = v4 & ~new_n309_;
  assign new_n311_ = ~v9 & ~new_n310_;
  assign new_n312_ = v3 & new_n311_;
  assign new_n313_ = ~new_n308_ & ~new_n312_;
  assign new_n314_ = ~v11 & ~new_n313_;
  assign new_n315_ = ~new_n306_ & ~new_n314_;
  assign new_n316_ = ~v10 & ~new_n315_;
  assign new_n317_ = v11 & ~new_n310_;
  assign new_n318_ = v10 & new_n317_;
  assign new_n319_ = ~v9 & new_n318_;
  assign new_n320_ = ~v6 & new_n319_;
  assign new_n321_ = ~new_n316_ & ~new_n320_;
  assign new_n322_ = ~v13 & ~new_n321_;
  assign new_n323_ = v9 & new_n121_;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign new_n325_ = ~v12 & ~new_n324_;
  assign new_n326_ = ~v13 & ~new_n207_;
  assign new_n327_ = v6 & ~new_n326_;
  assign new_n328_ = ~v4 & new_n327_;
  assign new_n329_ = ~v6 & v13;
  assign new_n330_ = ~new_n328_ & ~new_n329_;
  assign new_n331_ = v12 & ~new_n330_;
  assign new_n332_ = ~v11 & new_n331_;
  assign new_n333_ = ~v10 & new_n332_;
  assign new_n334_ = v9 & new_n333_;
  assign new_n335_ = ~new_n325_ & ~new_n334_;
  assign \v14.4  = ~v5 & ~new_n335_;
  assign new_n337_ = ~v12 & new_n199_;
  assign new_n338_ = ~v9 & new_n337_;
  assign \v14.5  = ~v5 & new_n338_;
  assign new_n340_ = v9 & ~v11;
  assign new_n341_ = new_n48_ & new_n340_;
  assign new_n342_ = ~new_n132_ & ~new_n341_;
  assign new_n343_ = ~v9 & new_n291_;
  assign new_n344_ = new_n342_ & ~new_n343_;
  assign new_n345_ = ~v10 & ~new_n344_;
  assign new_n346_ = v6 & new_n345_;
  assign new_n347_ = ~v5 & new_n346_;
  assign new_n348_ = v2 & new_n347_;
  assign \v14.6  = v0 & new_n348_;
  assign new_n350_ = ~v12 & ~new_n146_;
  assign new_n351_ = ~v12 & ~new_n350_;
  assign new_n352_ = v11 & ~new_n351_;
  assign new_n353_ = ~v11 & new_n147_;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = ~v10 & ~new_n354_;
  assign new_n356_ = v1 & new_n291_;
  assign new_n357_ = ~new_n293_ & ~new_n356_;
  assign new_n358_ = v10 & ~new_n357_;
  assign new_n359_ = ~new_n355_ & ~new_n358_;
  assign new_n360_ = v6 & ~new_n359_;
  assign new_n361_ = ~new_n291_ & ~new_n293_;
  assign new_n362_ = v10 & ~new_n361_;
  assign new_n363_ = ~v11 & ~new_n275_;
  assign new_n364_ = ~v10 & ~new_n363_;
  assign new_n365_ = ~new_n362_ & ~new_n364_;
  assign new_n366_ = ~v6 & ~new_n365_;
  assign new_n367_ = ~new_n360_ & ~new_n366_;
  assign new_n368_ = ~v10 & new_n63_;
  assign new_n369_ = v10 & new_n48_;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = v6 & ~new_n146_;
  assign new_n372_ = v6 & ~new_n371_;
  assign new_n373_ = ~new_n370_ & ~new_n372_;
  assign new_n374_ = ~v13 & ~new_n48_;
  assign new_n375_ = ~v10 & ~new_n374_;
  assign new_n376_ = ~new_n369_ & ~new_n375_;
  assign new_n377_ = v6 & ~new_n376_;
  assign new_n378_ = ~v5 & new_n377_;
  assign new_n379_ = v0 & new_n378_;
  assign new_n380_ = ~new_n373_ & ~new_n379_;
  assign new_n381_ = ~v11 & ~new_n380_;
  assign new_n382_ = ~v10 & ~v12;
  assign new_n383_ = ~v5 & new_n382_;
  assign new_n384_ = v0 & new_n383_;
  assign new_n385_ = ~new_n179_ & ~new_n384_;
  assign new_n386_ = v13 & ~new_n385_;
  assign new_n387_ = new_n161_ & new_n382_;
  assign new_n388_ = ~new_n179_ & ~new_n387_;
  assign new_n389_ = ~v13 & ~new_n388_;
  assign new_n390_ = ~new_n386_ & ~new_n389_;
  assign new_n391_ = v11 & ~new_n390_;
  assign new_n392_ = v6 & new_n391_;
  assign new_n393_ = ~new_n381_ & ~new_n392_;
  assign new_n394_ = new_n367_ & new_n393_;
  assign new_n395_ = ~v9 & ~new_n394_;
  assign new_n396_ = ~v0 & ~v12;
  assign new_n397_ = ~v0 & ~new_n42_;
  assign new_n398_ = ~new_n396_ & new_n397_;
  assign new_n399_ = ~v5 & ~new_n398_;
  assign new_n400_ = ~v5 & ~new_n399_;
  assign new_n401_ = v6 & ~new_n400_;
  assign new_n402_ = v6 & ~new_n401_;
  assign new_n403_ = ~v13 & ~new_n402_;
  assign new_n404_ = ~v11 & new_n403_;
  assign new_n405_ = ~v10 & new_n404_;
  assign new_n406_ = v9 & new_n405_;
  assign new_n407_ = ~new_n395_ & ~new_n406_;
  assign \v14.7  = v7 & ~new_n407_;
  assign new_n409_ = ~v6 & ~v9;
  assign new_n410_ = v10 & new_n409_;
  assign new_n411_ = v11 & new_n410_;
  assign new_n412_ = ~v12 & new_n411_;
  assign \v14.8  = v13 & new_n412_;
  assign new_n414_ = ~v11 & new_n410_;
  assign new_n415_ = v12 & new_n414_;
  assign \v14.9  = v13 & new_n415_;
  assign new_n417_ = ~v9 & ~v11;
  assign new_n418_ = new_n52_ & new_n417_;
  assign new_n419_ = new_n342_ & ~new_n418_;
  assign new_n420_ = v6 & ~new_n419_;
  assign new_n421_ = v0 & new_n420_;
  assign new_n422_ = new_n54_ & new_n306_;
  assign new_n423_ = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~v10 & ~new_n423_;
  assign \v14.10  = ~v5 & new_n424_;
  assign new_n426_ = ~v11 & ~v13;
  assign new_n427_ = v9 & new_n426_;
  assign new_n428_ = v11 & v13;
  assign new_n429_ = ~v9 & new_n428_;
  assign new_n430_ = ~new_n427_ & ~new_n429_;
  assign new_n431_ = v12 & ~new_n430_;
  assign new_n432_ = ~v11 & new_n54_;
  assign new_n433_ = v9 & new_n432_;
  assign new_n434_ = ~new_n431_ & ~new_n433_;
  assign new_n435_ = ~v10 & ~new_n434_;
  assign new_n436_ = v6 & new_n435_;
  assign new_n437_ = ~v5 & new_n436_;
  assign \v14.11  = v0 & new_n437_;
  assign new_n439_ = v8 & ~new_n112_;
  assign new_n440_ = ~v5 & new_n439_;
  assign new_n441_ = v6 & ~new_n218_;
  assign new_n442_ = v5 & new_n441_;
  assign new_n443_ = ~new_n440_ & ~new_n442_;
  assign new_n444_ = ~v13 & ~new_n443_;
  assign new_n445_ = v10 & ~new_n217_;
  assign new_n446_ = v13 & ~new_n445_;
  assign new_n447_ = v6 & new_n446_;
  assign new_n448_ = v5 & new_n447_;
  assign new_n449_ = ~new_n444_ & ~new_n448_;
  assign new_n450_ = ~v12 & ~new_n449_;
  assign new_n451_ = v10 & new_n426_;
  assign new_n452_ = v10 & ~new_n451_;
  assign new_n453_ = v12 & ~new_n452_;
  assign new_n454_ = v6 & new_n453_;
  assign new_n455_ = v5 & new_n454_;
  assign new_n456_ = ~new_n450_ & ~new_n455_;
  assign new_n457_ = ~v9 & ~new_n456_;
  assign new_n458_ = v5 & v6;
  assign new_n459_ = ~v5 & new_n329_;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~v11 & ~new_n460_;
  assign new_n462_ = ~v5 & v11;
  assign new_n463_ = new_n54_ & new_n462_;
  assign new_n464_ = ~new_n461_ & ~new_n463_;
  assign new_n465_ = ~v10 & ~new_n464_;
  assign new_n466_ = v9 & new_n465_;
  assign \v14.12  = new_n457_ | new_n466_;
  assign new_n468_ = ~v11 & ~new_n120_;
  assign new_n469_ = ~v10 & ~new_n468_;
  assign new_n470_ = ~new_n451_ & ~new_n469_;
  assign new_n471_ = ~v9 & ~new_n470_;
  assign new_n472_ = new_n125_ & new_n426_;
  assign new_n473_ = ~new_n471_ & ~new_n472_;
  assign new_n474_ = ~new_n323_ & new_n473_;
  assign new_n475_ = v10 & new_n63_;
  assign new_n476_ = ~v10 & new_n48_;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign new_n478_ = ~v11 & ~new_n477_;
  assign new_n479_ = ~v9 & new_n478_;
  assign new_n480_ = new_n474_ & ~new_n479_;
  assign new_n481_ = v6 & ~new_n480_;
  assign \v14.13  = v5 & new_n481_;
  assign new_n483_ = v6 & ~v11;
  assign new_n484_ = v0 & new_n483_;
  assign new_n485_ = v8 & v11;
  assign new_n486_ = ~v6 & new_n485_;
  assign new_n487_ = ~new_n484_ & ~new_n486_;
  assign new_n488_ = v10 & ~new_n487_;
  assign new_n489_ = v8 & new_n110_;
  assign new_n490_ = v3 & new_n489_;
  assign new_n491_ = ~new_n488_ & ~new_n490_;
  assign new_n492_ = ~v9 & ~new_n491_;
  assign new_n493_ = ~new_n116_ & ~new_n492_;
  assign new_n494_ = ~v13 & ~new_n493_;
  assign new_n495_ = ~new_n122_ & ~new_n494_;
  assign new_n496_ = ~v12 & ~new_n495_;
  assign new_n497_ = ~new_n128_ & ~new_n496_;
  assign \v14.14  = ~v5 & ~new_n497_;
  assign new_n499_ = ~v10 & new_n275_;
  assign new_n500_ = ~v9 & new_n499_;
  assign new_n501_ = v6 & new_n500_;
  assign new_n502_ = ~v5 & new_n501_;
  assign \v14.15  = v0 & new_n502_;
  assign new_n504_ = ~v10 & new_n432_;
  assign new_n505_ = v9 & new_n504_;
  assign new_n506_ = v6 & new_n505_;
  assign new_n507_ = ~v5 & new_n506_;
  assign \v14.16  = v0 & new_n507_;
  assign \v14.17  = v0 & new_n347_;
  assign new_n510_ = v8 & new_n199_;
  assign new_n511_ = ~new_n203_ & ~new_n510_;
  assign new_n512_ = ~v12 & ~new_n511_;
  assign new_n513_ = ~v10 & new_n127_;
  assign new_n514_ = v6 & new_n513_;
  assign new_n515_ = v0 & new_n514_;
  assign new_n516_ = ~new_n512_ & ~new_n515_;
  assign new_n517_ = ~v9 & ~new_n516_;
  assign new_n518_ = ~v10 & new_n426_;
  assign new_n519_ = v9 & new_n518_;
  assign new_n520_ = v6 & new_n519_;
  assign new_n521_ = v0 & new_n520_;
  assign new_n522_ = ~new_n517_ & ~new_n521_;
  assign new_n523_ = ~v9 & v11;
  assign new_n524_ = v6 & new_n523_;
  assign new_n525_ = v0 & new_n524_;
  assign new_n526_ = ~v6 & new_n340_;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_ = v12 & ~new_n527_;
  assign new_n529_ = new_n119_ & new_n293_;
  assign new_n530_ = ~new_n528_ & ~new_n529_;
  assign new_n531_ = v13 & ~new_n530_;
  assign new_n532_ = ~v9 & v12;
  assign new_n533_ = v6 & new_n532_;
  assign new_n534_ = v0 & new_n533_;
  assign new_n535_ = v9 & new_n102_;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = ~v13 & ~new_n536_;
  assign new_n538_ = ~new_n531_ & ~new_n537_;
  assign new_n539_ = ~v10 & ~new_n538_;
  assign new_n540_ = v10 & new_n432_;
  assign new_n541_ = ~v9 & new_n540_;
  assign new_n542_ = v6 & new_n541_;
  assign new_n543_ = v0 & new_n542_;
  assign new_n544_ = ~new_n539_ & ~new_n543_;
  assign new_n545_ = new_n522_ & new_n544_;
  assign new_n546_ = ~v5 & ~new_n545_;
  assign \v14.18  = \v14.13  | new_n546_;
  assign new_n548_ = new_n125_ & new_n127_;
  assign new_n549_ = ~v8 & ~v9;
  assign new_n550_ = ~v4 & new_n549_;
  assign new_n551_ = new_n54_ & new_n108_;
  assign new_n552_ = new_n550_ & new_n551_;
  assign new_n553_ = ~new_n548_ & ~new_n552_;
  assign new_n554_ = ~v6 & ~new_n553_;
  assign new_n555_ = v12 & ~new_n40_;
  assign new_n556_ = ~v11 & new_n555_;
  assign new_n557_ = ~new_n41_ & ~new_n556_;
  assign new_n558_ = v13 & ~new_n557_;
  assign new_n559_ = ~v9 & new_n558_;
  assign new_n560_ = ~v13 & ~new_n397_;
  assign new_n561_ = ~v11 & new_n560_;
  assign new_n562_ = v9 & new_n561_;
  assign new_n563_ = ~v4 & new_n562_;
  assign new_n564_ = ~new_n559_ & ~new_n563_;
  assign new_n565_ = ~v4 & v9;
  assign new_n566_ = new_n127_ & new_n565_;
  assign new_n567_ = new_n564_ & ~new_n566_;
  assign new_n568_ = v6 & ~new_n567_;
  assign new_n569_ = v3 & ~v4;
  assign new_n570_ = ~v8 & new_n417_;
  assign new_n571_ = new_n569_ & new_n570_;
  assign new_n572_ = ~new_n306_ & ~new_n571_;
  assign new_n573_ = ~v13 & ~new_n572_;
  assign new_n574_ = ~v12 & new_n573_;
  assign new_n575_ = ~new_n568_ & ~new_n574_;
  assign new_n576_ = ~v10 & ~new_n575_;
  assign new_n577_ = ~new_n554_ & ~new_n576_;
  assign \v14.19  = ~v5 & ~new_n577_;
  assign new_n579_ = ~v8 & new_n338_;
  assign new_n580_ = ~v5 & new_n579_;
  assign \v14.20  = ~v4 & new_n580_;
  assign new_n582_ = v0 & v12;
  assign new_n583_ = ~new_n396_ & ~new_n582_;
  assign new_n584_ = v11 & ~new_n583_;
  assign new_n585_ = ~v0 & new_n275_;
  assign new_n586_ = ~new_n584_ & ~new_n585_;
  assign new_n587_ = ~v10 & ~new_n586_;
  assign new_n588_ = new_n280_ & new_n293_;
  assign new_n589_ = ~new_n587_ & ~new_n588_;
  assign new_n590_ = ~v11 & new_n63_;
  assign new_n591_ = v11 & new_n48_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = ~v0 & ~new_n592_;
  assign new_n594_ = ~new_n102_ & ~new_n275_;
  assign new_n595_ = ~v13 & ~new_n594_;
  assign new_n596_ = v12 & ~new_n275_;
  assign new_n597_ = v13 & ~new_n596_;
  assign new_n598_ = ~new_n595_ & ~new_n597_;
  assign new_n599_ = v0 & ~new_n598_;
  assign new_n600_ = ~new_n593_ & ~new_n599_;
  assign new_n601_ = ~v10 & ~new_n600_;
  assign new_n602_ = v0 & v10;
  assign new_n603_ = new_n590_ & new_n602_;
  assign new_n604_ = ~new_n601_ & ~new_n603_;
  assign new_n605_ = new_n589_ & new_n604_;
  assign new_n606_ = ~v9 & ~new_n605_;
  assign new_n607_ = v0 & new_n519_;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = v6 & ~new_n608_;
  assign \v14.21  = ~v5 & new_n609_;
  assign new_n611_ = v10 & new_n120_;
  assign new_n612_ = v11 & ~v13;
  assign new_n613_ = ~v10 & new_n612_;
  assign new_n614_ = ~new_n611_ & ~new_n613_;
  assign new_n615_ = v0 & ~new_n614_;
  assign new_n616_ = ~v0 & new_n217_;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = ~v12 & ~new_n617_;
  assign new_n619_ = ~v9 & new_n618_;
  assign new_n620_ = v6 & new_n619_;
  assign \v14.22  = ~v5 & new_n620_;
  assign new_n622_ = ~v9 & new_n52_;
  assign new_n623_ = v9 & new_n54_;
  assign new_n624_ = ~new_n622_ & ~new_n623_;
  assign new_n625_ = ~v11 & ~new_n624_;
  assign new_n626_ = new_n342_ & ~new_n625_;
  assign new_n627_ = v0 & ~new_n626_;
  assign new_n628_ = ~v0 & v9;
  assign new_n629_ = ~v11 & new_n48_;
  assign new_n630_ = new_n628_ & new_n629_;
  assign new_n631_ = ~new_n627_ & ~new_n630_;
  assign new_n632_ = new_n52_ & new_n340_;
  assign new_n633_ = new_n631_ & ~new_n632_;
  assign new_n634_ = v6 & ~new_n633_;
  assign new_n635_ = v8 & ~v9;
  assign new_n636_ = v3 & new_n635_;
  assign new_n637_ = new_n432_ & new_n636_;
  assign new_n638_ = ~new_n634_ & ~new_n637_;
  assign new_n639_ = ~v10 & ~new_n638_;
  assign new_n640_ = ~v6 & new_n635_;
  assign new_n641_ = new_n551_ & new_n640_;
  assign new_n642_ = ~new_n639_ & ~new_n641_;
  assign new_n643_ = v6 & new_n471_;
  assign new_n644_ = ~v0 & new_n643_;
  assign new_n645_ = ~new_n122_ & ~new_n644_;
  assign new_n646_ = new_n54_ & new_n602_;
  assign new_n647_ = new_n477_ & ~new_n646_;
  assign new_n648_ = ~v11 & ~new_n647_;
  assign new_n649_ = ~v12 & ~new_n54_;
  assign new_n650_ = v11 & ~new_n649_;
  assign new_n651_ = ~v10 & new_n650_;
  assign new_n652_ = v0 & new_n651_;
  assign new_n653_ = ~new_n648_ & ~new_n652_;
  assign new_n654_ = ~v9 & ~new_n653_;
  assign new_n655_ = ~v0 & new_n125_;
  assign new_n656_ = new_n432_ & new_n655_;
  assign new_n657_ = ~new_n654_ & ~new_n656_;
  assign new_n658_ = new_n125_ & new_n590_;
  assign new_n659_ = new_n657_ & ~new_n658_;
  assign new_n660_ = v6 & ~new_n659_;
  assign new_n661_ = new_n55_ & new_n125_;
  assign new_n662_ = ~new_n660_ & ~new_n661_;
  assign new_n663_ = new_n645_ & new_n662_;
  assign new_n664_ = new_n642_ & new_n663_;
  assign new_n665_ = ~v5 & ~new_n664_;
  assign new_n666_ = new_n473_ & ~new_n479_;
  assign new_n667_ = v5 & ~new_n666_;
  assign new_n668_ = ~v1 & new_n101_;
  assign new_n669_ = v11 & new_n52_;
  assign new_n670_ = new_n668_ & new_n669_;
  assign new_n671_ = ~new_n667_ & ~new_n670_;
  assign new_n672_ = new_n591_ & new_n668_;
  assign new_n673_ = new_n671_ & ~new_n672_;
  assign new_n674_ = v5 & new_n323_;
  assign new_n675_ = new_n673_ & ~new_n674_;
  assign new_n676_ = v6 & ~new_n675_;
  assign \v14.23  = new_n665_ | new_n676_;
endmodule


