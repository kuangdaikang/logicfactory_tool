// Benchmark "arbiter" written by ABC on Fri Sep 15 11:24:47 2023

module arbiter ( 
    \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ,
    \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] ,
    \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] ,
    \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] ,
    \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] ,
    \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] ,
    \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] ,
    \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] ,
    \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] ,
    \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] ,
    \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] ,
    \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] ,
    \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] ,
    \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] ,
    \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] ,
    \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] ,
    \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] ,
    \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] ,
    \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] ,
    \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] ,
    \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] ,
    \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] ,
    \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] ,
    \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
    \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] ,
    \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] ,
    \grant[126] , \grant[127] , anyGrant  );
  input  \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
    \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
    \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
    \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
    \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
    \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
    \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
    \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
    \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
    \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
    \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
    \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
    \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
    \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
    \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
    \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
    \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
    \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
    \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
    \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
    \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] ,
    \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] ,
    \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] ,
    \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
    \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] ,
    \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_,
    new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_,
    new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_,
    new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_,
    new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_,
    new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3782_, new_n3783_, new_n3784_,
    new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_,
    new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_,
    new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_,
    new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_,
    new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4046_, new_n4047_, new_n4048_,
    new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_,
    new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_,
    new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_,
    new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_,
    new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_,
    new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_,
    new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_,
    new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_,
    new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_,
    new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_,
    new_n4263_, new_n4264_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_,
    new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_,
    new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_,
    new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_,
    new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_,
    new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_,
    new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4662_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_,
    new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_,
    new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4926_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_,
    new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_,
    new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_,
    new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_,
    new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_,
    new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_,
    new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_,
    new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_,
    new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_,
    new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_,
    new_n5055_, new_n5056_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_,
    new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_,
    new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_,
    new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_,
    new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_,
    new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_,
    new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_,
    new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_,
    new_n5319_, new_n5320_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_,
    new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_,
    new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5894_, new_n5895_, new_n5896_,
    new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_,
    new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_,
    new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_,
    new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_,
    new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6158_, new_n6159_, new_n6160_,
    new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_,
    new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_,
    new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_,
    new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_,
    new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_,
    new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_,
    new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_,
    new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_,
    new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_,
    new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_,
    new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_,
    new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_,
    new_n6375_, new_n6376_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_,
    new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_,
    new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6422_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_,
    new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_,
    new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_,
    new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_,
    new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_,
    new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_,
    new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_,
    new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_,
    new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_,
    new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_,
    new_n6639_, new_n6640_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6686_, new_n6687_, new_n6688_,
    new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_,
    new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_,
    new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_,
    new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_,
    new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_,
    new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_,
    new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6906_, new_n6907_, new_n6908_, new_n6909_,
    new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_,
    new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_,
    new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_,
    new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_,
    new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_,
    new_n6946_, new_n6947_, new_n6948_, new_n6950_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_,
    new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6994_, new_n6995_,
    new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_,
    new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_,
    new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_,
    new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7170_, new_n7171_, new_n7172_, new_n7173_,
    new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_,
    new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_, new_n7189_;
  INV_X1     g0000(.I(\priority[122] ), .ZN(new_n386_));
  INV_X1     g0001(.I(\req[120] ), .ZN(new_n387_));
  AOI21_X1   g0002(.A1(new_n387_), .A2(\priority[120] ), .B(\priority[121] ), .ZN(new_n388_));
  NAND2_X1   g0003(.A1(new_n388_), .A2(new_n386_), .ZN(new_n389_));
  INV_X1     g0004(.I(new_n389_), .ZN(new_n390_));
  INV_X1     g0005(.I(\priority[119] ), .ZN(new_n391_));
  INV_X1     g0006(.I(\req[117] ), .ZN(new_n392_));
  AOI21_X1   g0007(.A1(new_n392_), .A2(\priority[117] ), .B(\priority[118] ), .ZN(new_n393_));
  NAND2_X1   g0008(.A1(new_n393_), .A2(new_n391_), .ZN(new_n394_));
  INV_X1     g0009(.I(\priority[113] ), .ZN(new_n395_));
  INV_X1     g0010(.I(\req[111] ), .ZN(new_n396_));
  AOI21_X1   g0011(.A1(new_n396_), .A2(\priority[111] ), .B(\priority[112] ), .ZN(new_n397_));
  NAND2_X1   g0012(.A1(new_n397_), .A2(new_n395_), .ZN(new_n398_));
  INV_X1     g0013(.I(\priority[110] ), .ZN(new_n399_));
  INV_X1     g0014(.I(\req[108] ), .ZN(new_n400_));
  AOI21_X1   g0015(.A1(new_n400_), .A2(\priority[108] ), .B(\priority[109] ), .ZN(new_n401_));
  NAND2_X1   g0016(.A1(new_n401_), .A2(new_n399_), .ZN(new_n402_));
  INV_X1     g0017(.I(new_n402_), .ZN(new_n403_));
  INV_X1     g0018(.I(\priority[104] ), .ZN(new_n404_));
  INV_X1     g0019(.I(\req[102] ), .ZN(new_n405_));
  AOI21_X1   g0020(.A1(new_n405_), .A2(\priority[102] ), .B(\priority[103] ), .ZN(new_n406_));
  NAND2_X1   g0021(.A1(new_n406_), .A2(new_n404_), .ZN(new_n407_));
  INV_X1     g0022(.I(new_n407_), .ZN(new_n408_));
  INV_X1     g0023(.I(\priority[101] ), .ZN(new_n409_));
  INV_X1     g0024(.I(\req[99] ), .ZN(new_n410_));
  AOI21_X1   g0025(.A1(new_n410_), .A2(\priority[99] ), .B(\priority[100] ), .ZN(new_n411_));
  NAND2_X1   g0026(.A1(new_n411_), .A2(new_n409_), .ZN(new_n412_));
  INV_X1     g0027(.I(\priority[95] ), .ZN(new_n413_));
  INV_X1     g0028(.I(\req[93] ), .ZN(new_n414_));
  AOI21_X1   g0029(.A1(new_n414_), .A2(\priority[93] ), .B(\priority[94] ), .ZN(new_n415_));
  NAND2_X1   g0030(.A1(new_n415_), .A2(new_n413_), .ZN(new_n416_));
  INV_X1     g0031(.I(\priority[92] ), .ZN(new_n417_));
  INV_X1     g0032(.I(\req[90] ), .ZN(new_n418_));
  AOI21_X1   g0033(.A1(new_n418_), .A2(\priority[90] ), .B(\priority[91] ), .ZN(new_n419_));
  NAND2_X1   g0034(.A1(new_n419_), .A2(new_n417_), .ZN(new_n420_));
  INV_X1     g0035(.I(new_n420_), .ZN(new_n421_));
  INV_X1     g0036(.I(\priority[86] ), .ZN(new_n422_));
  INV_X1     g0037(.I(\req[84] ), .ZN(new_n423_));
  AOI21_X1   g0038(.A1(new_n423_), .A2(\priority[84] ), .B(\priority[85] ), .ZN(new_n424_));
  NAND2_X1   g0039(.A1(new_n424_), .A2(new_n422_), .ZN(new_n425_));
  INV_X1     g0040(.I(new_n425_), .ZN(new_n426_));
  INV_X1     g0041(.I(\priority[83] ), .ZN(new_n427_));
  INV_X1     g0042(.I(\req[81] ), .ZN(new_n428_));
  AOI21_X1   g0043(.A1(new_n428_), .A2(\priority[81] ), .B(\priority[82] ), .ZN(new_n429_));
  NAND2_X1   g0044(.A1(new_n429_), .A2(new_n427_), .ZN(new_n430_));
  INV_X1     g0045(.I(\priority[77] ), .ZN(new_n431_));
  INV_X1     g0046(.I(\req[75] ), .ZN(new_n432_));
  AOI21_X1   g0047(.A1(new_n432_), .A2(\priority[75] ), .B(\priority[76] ), .ZN(new_n433_));
  NAND2_X1   g0048(.A1(new_n433_), .A2(new_n431_), .ZN(new_n434_));
  INV_X1     g0049(.I(\priority[74] ), .ZN(new_n435_));
  INV_X1     g0050(.I(\req[72] ), .ZN(new_n436_));
  AOI21_X1   g0051(.A1(new_n436_), .A2(\priority[72] ), .B(\priority[73] ), .ZN(new_n437_));
  NAND2_X1   g0052(.A1(new_n437_), .A2(new_n435_), .ZN(new_n438_));
  INV_X1     g0053(.I(new_n438_), .ZN(new_n439_));
  INV_X1     g0054(.I(\priority[68] ), .ZN(new_n440_));
  INV_X1     g0055(.I(\req[66] ), .ZN(new_n441_));
  AOI21_X1   g0056(.A1(new_n441_), .A2(\priority[66] ), .B(\priority[67] ), .ZN(new_n442_));
  NAND2_X1   g0057(.A1(new_n442_), .A2(new_n440_), .ZN(new_n443_));
  INV_X1     g0058(.I(new_n443_), .ZN(new_n444_));
  INV_X1     g0059(.I(\priority[65] ), .ZN(new_n445_));
  INV_X1     g0060(.I(\req[63] ), .ZN(new_n446_));
  AOI21_X1   g0061(.A1(new_n446_), .A2(\priority[63] ), .B(\priority[64] ), .ZN(new_n447_));
  NAND2_X1   g0062(.A1(new_n447_), .A2(new_n445_), .ZN(new_n448_));
  INV_X1     g0063(.I(\priority[59] ), .ZN(new_n449_));
  INV_X1     g0064(.I(\req[57] ), .ZN(new_n450_));
  AOI21_X1   g0065(.A1(new_n450_), .A2(\priority[57] ), .B(\priority[58] ), .ZN(new_n451_));
  NAND2_X1   g0066(.A1(new_n451_), .A2(new_n449_), .ZN(new_n452_));
  INV_X1     g0067(.I(\priority[56] ), .ZN(new_n453_));
  INV_X1     g0068(.I(\req[54] ), .ZN(new_n454_));
  AOI21_X1   g0069(.A1(new_n454_), .A2(\priority[54] ), .B(\priority[55] ), .ZN(new_n455_));
  NAND2_X1   g0070(.A1(new_n455_), .A2(new_n453_), .ZN(new_n456_));
  INV_X1     g0071(.I(new_n456_), .ZN(new_n457_));
  INV_X1     g0072(.I(\priority[50] ), .ZN(new_n458_));
  INV_X1     g0073(.I(\req[48] ), .ZN(new_n459_));
  AOI21_X1   g0074(.A1(new_n459_), .A2(\priority[48] ), .B(\priority[49] ), .ZN(new_n460_));
  NAND2_X1   g0075(.A1(new_n460_), .A2(new_n458_), .ZN(new_n461_));
  INV_X1     g0076(.I(new_n461_), .ZN(new_n462_));
  INV_X1     g0077(.I(\priority[47] ), .ZN(new_n463_));
  INV_X1     g0078(.I(\req[45] ), .ZN(new_n464_));
  AOI21_X1   g0079(.A1(new_n464_), .A2(\priority[45] ), .B(\priority[46] ), .ZN(new_n465_));
  NAND2_X1   g0080(.A1(new_n465_), .A2(new_n463_), .ZN(new_n466_));
  INV_X1     g0081(.I(\priority[41] ), .ZN(new_n467_));
  INV_X1     g0082(.I(\req[39] ), .ZN(new_n468_));
  AOI21_X1   g0083(.A1(new_n468_), .A2(\priority[39] ), .B(\priority[40] ), .ZN(new_n469_));
  NAND2_X1   g0084(.A1(new_n469_), .A2(new_n467_), .ZN(new_n470_));
  INV_X1     g0085(.I(\priority[38] ), .ZN(new_n471_));
  INV_X1     g0086(.I(\req[36] ), .ZN(new_n472_));
  AOI21_X1   g0087(.A1(new_n472_), .A2(\priority[36] ), .B(\priority[37] ), .ZN(new_n473_));
  NAND2_X1   g0088(.A1(new_n473_), .A2(new_n471_), .ZN(new_n474_));
  INV_X1     g0089(.I(new_n474_), .ZN(new_n475_));
  INV_X1     g0090(.I(\priority[32] ), .ZN(new_n476_));
  INV_X1     g0091(.I(\req[30] ), .ZN(new_n477_));
  AOI21_X1   g0092(.A1(new_n477_), .A2(\priority[30] ), .B(\priority[31] ), .ZN(new_n478_));
  NAND2_X1   g0093(.A1(new_n478_), .A2(new_n476_), .ZN(new_n479_));
  INV_X1     g0094(.I(new_n479_), .ZN(new_n480_));
  INV_X1     g0095(.I(\priority[29] ), .ZN(new_n481_));
  INV_X1     g0096(.I(\req[27] ), .ZN(new_n482_));
  AOI21_X1   g0097(.A1(new_n482_), .A2(\priority[27] ), .B(\priority[28] ), .ZN(new_n483_));
  NAND2_X1   g0098(.A1(new_n483_), .A2(new_n481_), .ZN(new_n484_));
  INV_X1     g0099(.I(\priority[23] ), .ZN(new_n485_));
  INV_X1     g0100(.I(\req[21] ), .ZN(new_n486_));
  AOI21_X1   g0101(.A1(new_n486_), .A2(\priority[21] ), .B(\priority[22] ), .ZN(new_n487_));
  NAND2_X1   g0102(.A1(new_n487_), .A2(new_n485_), .ZN(new_n488_));
  INV_X1     g0103(.I(\priority[20] ), .ZN(new_n489_));
  INV_X1     g0104(.I(\req[18] ), .ZN(new_n490_));
  AOI21_X1   g0105(.A1(new_n490_), .A2(\priority[18] ), .B(\priority[19] ), .ZN(new_n491_));
  NAND2_X1   g0106(.A1(new_n491_), .A2(new_n489_), .ZN(new_n492_));
  INV_X1     g0107(.I(new_n492_), .ZN(new_n493_));
  INV_X1     g0108(.I(\priority[14] ), .ZN(new_n494_));
  INV_X1     g0109(.I(\req[12] ), .ZN(new_n495_));
  AOI21_X1   g0110(.A1(new_n495_), .A2(\priority[12] ), .B(\priority[13] ), .ZN(new_n496_));
  NAND2_X1   g0111(.A1(new_n496_), .A2(new_n494_), .ZN(new_n497_));
  INV_X1     g0112(.I(new_n497_), .ZN(new_n498_));
  INV_X1     g0113(.I(\priority[11] ), .ZN(new_n499_));
  INV_X1     g0114(.I(\req[9] ), .ZN(new_n500_));
  AOI21_X1   g0115(.A1(new_n500_), .A2(\priority[9] ), .B(\priority[10] ), .ZN(new_n501_));
  NAND2_X1   g0116(.A1(new_n501_), .A2(new_n499_), .ZN(new_n502_));
  INV_X1     g0117(.I(\priority[5] ), .ZN(new_n503_));
  INV_X1     g0118(.I(\req[3] ), .ZN(new_n504_));
  AOI21_X1   g0119(.A1(new_n504_), .A2(\priority[3] ), .B(\priority[4] ), .ZN(new_n505_));
  NAND2_X1   g0120(.A1(new_n505_), .A2(new_n503_), .ZN(new_n506_));
  INV_X1     g0121(.I(\req[1] ), .ZN(new_n507_));
  AOI21_X1   g0122(.A1(new_n507_), .A2(\priority[1] ), .B(\priority[2] ), .ZN(new_n508_));
  OR2_X2     g0123(.A1(\req[2] ), .A2(\req[3] ), .Z(new_n509_));
  NOR2_X1    g0124(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1     g0125(.I(\req[4] ), .ZN(new_n511_));
  NOR2_X1    g0126(.A1(new_n511_), .A2(\priority[5] ), .ZN(new_n512_));
  OR2_X2     g0127(.A1(\req[5] ), .A2(\req[6] ), .Z(new_n513_));
  NOR2_X1    g0128(.A1(new_n513_), .A2(new_n512_), .ZN(new_n514_));
  OAI21_X1   g0129(.A1(new_n506_), .A2(new_n510_), .B(new_n514_), .ZN(new_n515_));
  INV_X1     g0130(.I(\priority[8] ), .ZN(new_n516_));
  INV_X1     g0131(.I(\req[6] ), .ZN(new_n517_));
  AOI21_X1   g0132(.A1(new_n517_), .A2(\priority[6] ), .B(\priority[7] ), .ZN(new_n518_));
  NAND2_X1   g0133(.A1(new_n518_), .A2(new_n516_), .ZN(new_n519_));
  INV_X1     g0134(.I(new_n519_), .ZN(new_n520_));
  INV_X1     g0135(.I(\req[7] ), .ZN(new_n521_));
  NOR2_X1    g0136(.A1(new_n521_), .A2(\priority[8] ), .ZN(new_n522_));
  OR2_X2     g0137(.A1(\req[8] ), .A2(\req[9] ), .Z(new_n523_));
  NOR2_X1    g0138(.A1(new_n523_), .A2(new_n522_), .ZN(new_n524_));
  INV_X1     g0139(.I(new_n524_), .ZN(new_n525_));
  AOI21_X1   g0140(.A1(new_n515_), .A2(new_n520_), .B(new_n525_), .ZN(new_n526_));
  INV_X1     g0141(.I(\req[10] ), .ZN(new_n527_));
  NOR2_X1    g0142(.A1(new_n527_), .A2(\priority[11] ), .ZN(new_n528_));
  OR2_X2     g0143(.A1(\req[11] ), .A2(\req[12] ), .Z(new_n529_));
  NOR2_X1    g0144(.A1(new_n529_), .A2(new_n528_), .ZN(new_n530_));
  OAI21_X1   g0145(.A1(new_n526_), .A2(new_n502_), .B(new_n530_), .ZN(new_n531_));
  INV_X1     g0146(.I(\req[13] ), .ZN(new_n532_));
  NOR2_X1    g0147(.A1(new_n532_), .A2(\priority[14] ), .ZN(new_n533_));
  OR2_X2     g0148(.A1(\req[14] ), .A2(\req[15] ), .Z(new_n534_));
  NOR2_X1    g0149(.A1(new_n534_), .A2(new_n533_), .ZN(new_n535_));
  INV_X1     g0150(.I(new_n535_), .ZN(new_n536_));
  AOI21_X1   g0151(.A1(new_n531_), .A2(new_n498_), .B(new_n536_), .ZN(new_n537_));
  INV_X1     g0152(.I(\priority[17] ), .ZN(new_n538_));
  INV_X1     g0153(.I(\req[15] ), .ZN(new_n539_));
  AOI21_X1   g0154(.A1(new_n539_), .A2(\priority[15] ), .B(\priority[16] ), .ZN(new_n540_));
  NAND2_X1   g0155(.A1(new_n540_), .A2(new_n538_), .ZN(new_n541_));
  INV_X1     g0156(.I(\req[16] ), .ZN(new_n542_));
  NOR2_X1    g0157(.A1(new_n542_), .A2(\priority[17] ), .ZN(new_n543_));
  OR2_X2     g0158(.A1(\req[17] ), .A2(\req[18] ), .Z(new_n544_));
  NOR2_X1    g0159(.A1(new_n544_), .A2(new_n543_), .ZN(new_n545_));
  OAI21_X1   g0160(.A1(new_n537_), .A2(new_n541_), .B(new_n545_), .ZN(new_n546_));
  INV_X1     g0161(.I(\req[19] ), .ZN(new_n547_));
  NOR2_X1    g0162(.A1(new_n547_), .A2(\priority[20] ), .ZN(new_n548_));
  OR2_X2     g0163(.A1(\req[20] ), .A2(\req[21] ), .Z(new_n549_));
  NOR2_X1    g0164(.A1(new_n549_), .A2(new_n548_), .ZN(new_n550_));
  INV_X1     g0165(.I(new_n550_), .ZN(new_n551_));
  AOI21_X1   g0166(.A1(new_n546_), .A2(new_n493_), .B(new_n551_), .ZN(new_n552_));
  INV_X1     g0167(.I(\req[22] ), .ZN(new_n553_));
  NOR2_X1    g0168(.A1(new_n553_), .A2(\priority[23] ), .ZN(new_n554_));
  OR2_X2     g0169(.A1(\req[23] ), .A2(\req[24] ), .Z(new_n555_));
  NOR2_X1    g0170(.A1(new_n555_), .A2(new_n554_), .ZN(new_n556_));
  OAI21_X1   g0171(.A1(new_n552_), .A2(new_n488_), .B(new_n556_), .ZN(new_n557_));
  INV_X1     g0172(.I(\priority[26] ), .ZN(new_n558_));
  INV_X1     g0173(.I(\req[24] ), .ZN(new_n559_));
  AOI21_X1   g0174(.A1(new_n559_), .A2(\priority[24] ), .B(\priority[25] ), .ZN(new_n560_));
  NAND2_X1   g0175(.A1(new_n560_), .A2(new_n558_), .ZN(new_n561_));
  INV_X1     g0176(.I(new_n561_), .ZN(new_n562_));
  INV_X1     g0177(.I(\req[25] ), .ZN(new_n563_));
  NOR2_X1    g0178(.A1(new_n563_), .A2(\priority[26] ), .ZN(new_n564_));
  OR2_X2     g0179(.A1(\req[26] ), .A2(\req[27] ), .Z(new_n565_));
  NOR2_X1    g0180(.A1(new_n565_), .A2(new_n564_), .ZN(new_n566_));
  INV_X1     g0181(.I(new_n566_), .ZN(new_n567_));
  AOI21_X1   g0182(.A1(new_n557_), .A2(new_n562_), .B(new_n567_), .ZN(new_n568_));
  INV_X1     g0183(.I(\req[28] ), .ZN(new_n569_));
  NOR2_X1    g0184(.A1(new_n569_), .A2(\priority[29] ), .ZN(new_n570_));
  OR2_X2     g0185(.A1(\req[29] ), .A2(\req[30] ), .Z(new_n571_));
  NOR2_X1    g0186(.A1(new_n571_), .A2(new_n570_), .ZN(new_n572_));
  OAI21_X1   g0187(.A1(new_n568_), .A2(new_n484_), .B(new_n572_), .ZN(new_n573_));
  INV_X1     g0188(.I(\req[31] ), .ZN(new_n574_));
  NOR2_X1    g0189(.A1(new_n574_), .A2(\priority[32] ), .ZN(new_n575_));
  OR2_X2     g0190(.A1(\req[32] ), .A2(\req[33] ), .Z(new_n576_));
  NOR2_X1    g0191(.A1(new_n576_), .A2(new_n575_), .ZN(new_n577_));
  INV_X1     g0192(.I(new_n577_), .ZN(new_n578_));
  AOI21_X1   g0193(.A1(new_n573_), .A2(new_n480_), .B(new_n578_), .ZN(new_n579_));
  INV_X1     g0194(.I(\priority[35] ), .ZN(new_n580_));
  INV_X1     g0195(.I(\req[33] ), .ZN(new_n581_));
  AOI21_X1   g0196(.A1(new_n581_), .A2(\priority[33] ), .B(\priority[34] ), .ZN(new_n582_));
  NAND2_X1   g0197(.A1(new_n582_), .A2(new_n580_), .ZN(new_n583_));
  INV_X1     g0198(.I(\req[34] ), .ZN(new_n584_));
  NOR2_X1    g0199(.A1(new_n584_), .A2(\priority[35] ), .ZN(new_n585_));
  OR2_X2     g0200(.A1(\req[35] ), .A2(\req[36] ), .Z(new_n586_));
  NOR2_X1    g0201(.A1(new_n586_), .A2(new_n585_), .ZN(new_n587_));
  OAI21_X1   g0202(.A1(new_n579_), .A2(new_n583_), .B(new_n587_), .ZN(new_n588_));
  INV_X1     g0203(.I(\req[37] ), .ZN(new_n589_));
  NOR2_X1    g0204(.A1(new_n589_), .A2(\priority[38] ), .ZN(new_n590_));
  OR2_X2     g0205(.A1(\req[38] ), .A2(\req[39] ), .Z(new_n591_));
  NOR2_X1    g0206(.A1(new_n591_), .A2(new_n590_), .ZN(new_n592_));
  INV_X1     g0207(.I(new_n592_), .ZN(new_n593_));
  AOI21_X1   g0208(.A1(new_n588_), .A2(new_n475_), .B(new_n593_), .ZN(new_n594_));
  INV_X1     g0209(.I(\req[40] ), .ZN(new_n595_));
  NOR2_X1    g0210(.A1(new_n595_), .A2(\priority[41] ), .ZN(new_n596_));
  OR2_X2     g0211(.A1(\req[41] ), .A2(\req[42] ), .Z(new_n597_));
  NOR2_X1    g0212(.A1(new_n597_), .A2(new_n596_), .ZN(new_n598_));
  OAI21_X1   g0213(.A1(new_n594_), .A2(new_n470_), .B(new_n598_), .ZN(new_n599_));
  INV_X1     g0214(.I(\priority[44] ), .ZN(new_n600_));
  INV_X1     g0215(.I(\req[42] ), .ZN(new_n601_));
  AOI21_X1   g0216(.A1(new_n601_), .A2(\priority[42] ), .B(\priority[43] ), .ZN(new_n602_));
  NAND2_X1   g0217(.A1(new_n602_), .A2(new_n600_), .ZN(new_n603_));
  INV_X1     g0218(.I(new_n603_), .ZN(new_n604_));
  INV_X1     g0219(.I(\req[43] ), .ZN(new_n605_));
  NOR2_X1    g0220(.A1(new_n605_), .A2(\priority[44] ), .ZN(new_n606_));
  OR2_X2     g0221(.A1(\req[44] ), .A2(\req[45] ), .Z(new_n607_));
  NOR2_X1    g0222(.A1(new_n607_), .A2(new_n606_), .ZN(new_n608_));
  INV_X1     g0223(.I(new_n608_), .ZN(new_n609_));
  AOI21_X1   g0224(.A1(new_n599_), .A2(new_n604_), .B(new_n609_), .ZN(new_n610_));
  INV_X1     g0225(.I(\req[46] ), .ZN(new_n611_));
  NOR2_X1    g0226(.A1(new_n611_), .A2(\priority[47] ), .ZN(new_n612_));
  OR2_X2     g0227(.A1(\req[47] ), .A2(\req[48] ), .Z(new_n613_));
  NOR2_X1    g0228(.A1(new_n613_), .A2(new_n612_), .ZN(new_n614_));
  OAI21_X1   g0229(.A1(new_n610_), .A2(new_n466_), .B(new_n614_), .ZN(new_n615_));
  INV_X1     g0230(.I(\req[49] ), .ZN(new_n616_));
  NOR2_X1    g0231(.A1(new_n616_), .A2(\priority[50] ), .ZN(new_n617_));
  OR2_X2     g0232(.A1(\req[50] ), .A2(\req[51] ), .Z(new_n618_));
  NOR2_X1    g0233(.A1(new_n618_), .A2(new_n617_), .ZN(new_n619_));
  INV_X1     g0234(.I(new_n619_), .ZN(new_n620_));
  AOI21_X1   g0235(.A1(new_n615_), .A2(new_n462_), .B(new_n620_), .ZN(new_n621_));
  INV_X1     g0236(.I(\priority[53] ), .ZN(new_n622_));
  INV_X1     g0237(.I(\req[51] ), .ZN(new_n623_));
  AOI21_X1   g0238(.A1(new_n623_), .A2(\priority[51] ), .B(\priority[52] ), .ZN(new_n624_));
  NAND2_X1   g0239(.A1(new_n624_), .A2(new_n622_), .ZN(new_n625_));
  INV_X1     g0240(.I(\req[52] ), .ZN(new_n626_));
  NOR2_X1    g0241(.A1(new_n626_), .A2(\priority[53] ), .ZN(new_n627_));
  OR2_X2     g0242(.A1(\req[53] ), .A2(\req[54] ), .Z(new_n628_));
  NOR2_X1    g0243(.A1(new_n628_), .A2(new_n627_), .ZN(new_n629_));
  OAI21_X1   g0244(.A1(new_n621_), .A2(new_n625_), .B(new_n629_), .ZN(new_n630_));
  INV_X1     g0245(.I(\req[55] ), .ZN(new_n631_));
  NOR2_X1    g0246(.A1(new_n631_), .A2(\priority[56] ), .ZN(new_n632_));
  OR2_X2     g0247(.A1(\req[56] ), .A2(\req[57] ), .Z(new_n633_));
  NOR2_X1    g0248(.A1(new_n633_), .A2(new_n632_), .ZN(new_n634_));
  INV_X1     g0249(.I(new_n634_), .ZN(new_n635_));
  AOI21_X1   g0250(.A1(new_n630_), .A2(new_n457_), .B(new_n635_), .ZN(new_n636_));
  INV_X1     g0251(.I(\req[58] ), .ZN(new_n637_));
  NOR2_X1    g0252(.A1(new_n637_), .A2(\priority[59] ), .ZN(new_n638_));
  OR2_X2     g0253(.A1(\req[59] ), .A2(\req[60] ), .Z(new_n639_));
  NOR2_X1    g0254(.A1(new_n639_), .A2(new_n638_), .ZN(new_n640_));
  OAI21_X1   g0255(.A1(new_n636_), .A2(new_n452_), .B(new_n640_), .ZN(new_n641_));
  INV_X1     g0256(.I(\priority[62] ), .ZN(new_n642_));
  INV_X1     g0257(.I(\req[60] ), .ZN(new_n643_));
  AOI21_X1   g0258(.A1(new_n643_), .A2(\priority[60] ), .B(\priority[61] ), .ZN(new_n644_));
  NAND2_X1   g0259(.A1(new_n644_), .A2(new_n642_), .ZN(new_n645_));
  INV_X1     g0260(.I(new_n645_), .ZN(new_n646_));
  INV_X1     g0261(.I(\req[61] ), .ZN(new_n647_));
  NOR2_X1    g0262(.A1(new_n647_), .A2(\priority[62] ), .ZN(new_n648_));
  OR2_X2     g0263(.A1(\req[62] ), .A2(\req[63] ), .Z(new_n649_));
  NOR2_X1    g0264(.A1(new_n649_), .A2(new_n648_), .ZN(new_n650_));
  INV_X1     g0265(.I(new_n650_), .ZN(new_n651_));
  AOI21_X1   g0266(.A1(new_n641_), .A2(new_n646_), .B(new_n651_), .ZN(new_n652_));
  INV_X1     g0267(.I(\req[64] ), .ZN(new_n653_));
  NOR2_X1    g0268(.A1(new_n653_), .A2(\priority[65] ), .ZN(new_n654_));
  OR2_X2     g0269(.A1(\req[65] ), .A2(\req[66] ), .Z(new_n655_));
  NOR2_X1    g0270(.A1(new_n655_), .A2(new_n654_), .ZN(new_n656_));
  OAI21_X1   g0271(.A1(new_n652_), .A2(new_n448_), .B(new_n656_), .ZN(new_n657_));
  INV_X1     g0272(.I(\req[67] ), .ZN(new_n658_));
  NOR2_X1    g0273(.A1(new_n658_), .A2(\priority[68] ), .ZN(new_n659_));
  OR2_X2     g0274(.A1(\req[68] ), .A2(\req[69] ), .Z(new_n660_));
  NOR2_X1    g0275(.A1(new_n660_), .A2(new_n659_), .ZN(new_n661_));
  INV_X1     g0276(.I(new_n661_), .ZN(new_n662_));
  AOI21_X1   g0277(.A1(new_n657_), .A2(new_n444_), .B(new_n662_), .ZN(new_n663_));
  INV_X1     g0278(.I(\priority[71] ), .ZN(new_n664_));
  INV_X1     g0279(.I(\req[69] ), .ZN(new_n665_));
  AOI21_X1   g0280(.A1(new_n665_), .A2(\priority[69] ), .B(\priority[70] ), .ZN(new_n666_));
  NAND2_X1   g0281(.A1(new_n666_), .A2(new_n664_), .ZN(new_n667_));
  INV_X1     g0282(.I(\req[70] ), .ZN(new_n668_));
  NOR2_X1    g0283(.A1(new_n668_), .A2(\priority[71] ), .ZN(new_n669_));
  OR2_X2     g0284(.A1(\req[71] ), .A2(\req[72] ), .Z(new_n670_));
  NOR2_X1    g0285(.A1(new_n670_), .A2(new_n669_), .ZN(new_n671_));
  OAI21_X1   g0286(.A1(new_n663_), .A2(new_n667_), .B(new_n671_), .ZN(new_n672_));
  INV_X1     g0287(.I(\req[73] ), .ZN(new_n673_));
  NOR2_X1    g0288(.A1(new_n673_), .A2(\priority[74] ), .ZN(new_n674_));
  OR2_X2     g0289(.A1(\req[74] ), .A2(\req[75] ), .Z(new_n675_));
  NOR2_X1    g0290(.A1(new_n675_), .A2(new_n674_), .ZN(new_n676_));
  INV_X1     g0291(.I(new_n676_), .ZN(new_n677_));
  AOI21_X1   g0292(.A1(new_n672_), .A2(new_n439_), .B(new_n677_), .ZN(new_n678_));
  INV_X1     g0293(.I(\req[76] ), .ZN(new_n679_));
  NOR2_X1    g0294(.A1(new_n679_), .A2(\priority[77] ), .ZN(new_n680_));
  OR2_X2     g0295(.A1(\req[77] ), .A2(\req[78] ), .Z(new_n681_));
  NOR2_X1    g0296(.A1(new_n681_), .A2(new_n680_), .ZN(new_n682_));
  OAI21_X1   g0297(.A1(new_n678_), .A2(new_n434_), .B(new_n682_), .ZN(new_n683_));
  INV_X1     g0298(.I(\priority[80] ), .ZN(new_n684_));
  INV_X1     g0299(.I(\req[78] ), .ZN(new_n685_));
  AOI21_X1   g0300(.A1(new_n685_), .A2(\priority[78] ), .B(\priority[79] ), .ZN(new_n686_));
  NAND2_X1   g0301(.A1(new_n686_), .A2(new_n684_), .ZN(new_n687_));
  INV_X1     g0302(.I(new_n687_), .ZN(new_n688_));
  INV_X1     g0303(.I(\req[79] ), .ZN(new_n689_));
  NOR2_X1    g0304(.A1(new_n689_), .A2(\priority[80] ), .ZN(new_n690_));
  OR2_X2     g0305(.A1(\req[80] ), .A2(\req[81] ), .Z(new_n691_));
  NOR2_X1    g0306(.A1(new_n691_), .A2(new_n690_), .ZN(new_n692_));
  INV_X1     g0307(.I(new_n692_), .ZN(new_n693_));
  AOI21_X1   g0308(.A1(new_n683_), .A2(new_n688_), .B(new_n693_), .ZN(new_n694_));
  INV_X1     g0309(.I(\req[82] ), .ZN(new_n695_));
  NOR2_X1    g0310(.A1(new_n695_), .A2(\priority[83] ), .ZN(new_n696_));
  OR2_X2     g0311(.A1(\req[83] ), .A2(\req[84] ), .Z(new_n697_));
  NOR2_X1    g0312(.A1(new_n697_), .A2(new_n696_), .ZN(new_n698_));
  OAI21_X1   g0313(.A1(new_n694_), .A2(new_n430_), .B(new_n698_), .ZN(new_n699_));
  INV_X1     g0314(.I(\req[85] ), .ZN(new_n700_));
  NOR2_X1    g0315(.A1(new_n700_), .A2(\priority[86] ), .ZN(new_n701_));
  OR2_X2     g0316(.A1(\req[86] ), .A2(\req[87] ), .Z(new_n702_));
  NOR2_X1    g0317(.A1(new_n702_), .A2(new_n701_), .ZN(new_n703_));
  INV_X1     g0318(.I(new_n703_), .ZN(new_n704_));
  AOI21_X1   g0319(.A1(new_n699_), .A2(new_n426_), .B(new_n704_), .ZN(new_n705_));
  INV_X1     g0320(.I(\priority[89] ), .ZN(new_n706_));
  INV_X1     g0321(.I(\req[87] ), .ZN(new_n707_));
  AOI21_X1   g0322(.A1(new_n707_), .A2(\priority[87] ), .B(\priority[88] ), .ZN(new_n708_));
  NAND2_X1   g0323(.A1(new_n708_), .A2(new_n706_), .ZN(new_n709_));
  INV_X1     g0324(.I(\req[88] ), .ZN(new_n710_));
  NOR2_X1    g0325(.A1(new_n710_), .A2(\priority[89] ), .ZN(new_n711_));
  OR2_X2     g0326(.A1(\req[89] ), .A2(\req[90] ), .Z(new_n712_));
  NOR2_X1    g0327(.A1(new_n712_), .A2(new_n711_), .ZN(new_n713_));
  OAI21_X1   g0328(.A1(new_n705_), .A2(new_n709_), .B(new_n713_), .ZN(new_n714_));
  INV_X1     g0329(.I(\req[91] ), .ZN(new_n715_));
  NOR2_X1    g0330(.A1(new_n715_), .A2(\priority[92] ), .ZN(new_n716_));
  OR2_X2     g0331(.A1(\req[92] ), .A2(\req[93] ), .Z(new_n717_));
  NOR2_X1    g0332(.A1(new_n717_), .A2(new_n716_), .ZN(new_n718_));
  INV_X1     g0333(.I(new_n718_), .ZN(new_n719_));
  AOI21_X1   g0334(.A1(new_n714_), .A2(new_n421_), .B(new_n719_), .ZN(new_n720_));
  INV_X1     g0335(.I(\req[94] ), .ZN(new_n721_));
  NOR2_X1    g0336(.A1(new_n721_), .A2(\priority[95] ), .ZN(new_n722_));
  OR2_X2     g0337(.A1(\req[95] ), .A2(\req[96] ), .Z(new_n723_));
  NOR2_X1    g0338(.A1(new_n723_), .A2(new_n722_), .ZN(new_n724_));
  OAI21_X1   g0339(.A1(new_n720_), .A2(new_n416_), .B(new_n724_), .ZN(new_n725_));
  INV_X1     g0340(.I(\priority[98] ), .ZN(new_n726_));
  INV_X1     g0341(.I(\req[96] ), .ZN(new_n727_));
  AOI21_X1   g0342(.A1(new_n727_), .A2(\priority[96] ), .B(\priority[97] ), .ZN(new_n728_));
  NAND2_X1   g0343(.A1(new_n728_), .A2(new_n726_), .ZN(new_n729_));
  INV_X1     g0344(.I(new_n729_), .ZN(new_n730_));
  INV_X1     g0345(.I(\req[97] ), .ZN(new_n731_));
  NOR2_X1    g0346(.A1(new_n731_), .A2(\priority[98] ), .ZN(new_n732_));
  OR2_X2     g0347(.A1(\req[98] ), .A2(\req[99] ), .Z(new_n733_));
  NOR2_X1    g0348(.A1(new_n733_), .A2(new_n732_), .ZN(new_n734_));
  INV_X1     g0349(.I(new_n734_), .ZN(new_n735_));
  AOI21_X1   g0350(.A1(new_n725_), .A2(new_n730_), .B(new_n735_), .ZN(new_n736_));
  INV_X1     g0351(.I(\req[100] ), .ZN(new_n737_));
  NOR2_X1    g0352(.A1(new_n737_), .A2(\priority[101] ), .ZN(new_n738_));
  OR2_X2     g0353(.A1(\req[101] ), .A2(\req[102] ), .Z(new_n739_));
  NOR2_X1    g0354(.A1(new_n739_), .A2(new_n738_), .ZN(new_n740_));
  OAI21_X1   g0355(.A1(new_n736_), .A2(new_n412_), .B(new_n740_), .ZN(new_n741_));
  INV_X1     g0356(.I(\req[103] ), .ZN(new_n742_));
  NOR2_X1    g0357(.A1(new_n742_), .A2(\priority[104] ), .ZN(new_n743_));
  OR2_X2     g0358(.A1(\req[104] ), .A2(\req[105] ), .Z(new_n744_));
  NOR2_X1    g0359(.A1(new_n744_), .A2(new_n743_), .ZN(new_n745_));
  INV_X1     g0360(.I(new_n745_), .ZN(new_n746_));
  AOI21_X1   g0361(.A1(new_n741_), .A2(new_n408_), .B(new_n746_), .ZN(new_n747_));
  INV_X1     g0362(.I(\priority[107] ), .ZN(new_n748_));
  INV_X1     g0363(.I(\req[105] ), .ZN(new_n749_));
  AOI21_X1   g0364(.A1(new_n749_), .A2(\priority[105] ), .B(\priority[106] ), .ZN(new_n750_));
  NAND2_X1   g0365(.A1(new_n750_), .A2(new_n748_), .ZN(new_n751_));
  INV_X1     g0366(.I(\req[106] ), .ZN(new_n752_));
  NOR2_X1    g0367(.A1(new_n752_), .A2(\priority[107] ), .ZN(new_n753_));
  OR2_X2     g0368(.A1(\req[107] ), .A2(\req[108] ), .Z(new_n754_));
  NOR2_X1    g0369(.A1(new_n754_), .A2(new_n753_), .ZN(new_n755_));
  OAI21_X1   g0370(.A1(new_n747_), .A2(new_n751_), .B(new_n755_), .ZN(new_n756_));
  INV_X1     g0371(.I(\req[109] ), .ZN(new_n757_));
  NOR2_X1    g0372(.A1(new_n757_), .A2(\priority[110] ), .ZN(new_n758_));
  OR2_X2     g0373(.A1(\req[110] ), .A2(\req[111] ), .Z(new_n759_));
  NOR2_X1    g0374(.A1(new_n759_), .A2(new_n758_), .ZN(new_n760_));
  INV_X1     g0375(.I(new_n760_), .ZN(new_n761_));
  AOI21_X1   g0376(.A1(new_n756_), .A2(new_n403_), .B(new_n761_), .ZN(new_n762_));
  INV_X1     g0377(.I(\req[112] ), .ZN(new_n763_));
  NOR2_X1    g0378(.A1(new_n763_), .A2(\priority[113] ), .ZN(new_n764_));
  OR2_X2     g0379(.A1(\req[113] ), .A2(\req[114] ), .Z(new_n765_));
  NOR2_X1    g0380(.A1(new_n765_), .A2(new_n764_), .ZN(new_n766_));
  OAI21_X1   g0381(.A1(new_n762_), .A2(new_n398_), .B(new_n766_), .ZN(new_n767_));
  INV_X1     g0382(.I(\priority[116] ), .ZN(new_n768_));
  INV_X1     g0383(.I(\req[114] ), .ZN(new_n769_));
  AOI21_X1   g0384(.A1(new_n769_), .A2(\priority[114] ), .B(\priority[115] ), .ZN(new_n770_));
  NAND2_X1   g0385(.A1(new_n770_), .A2(new_n768_), .ZN(new_n771_));
  INV_X1     g0386(.I(new_n771_), .ZN(new_n772_));
  INV_X1     g0387(.I(\req[115] ), .ZN(new_n773_));
  NOR2_X1    g0388(.A1(new_n773_), .A2(\priority[116] ), .ZN(new_n774_));
  OR2_X2     g0389(.A1(\req[116] ), .A2(\req[117] ), .Z(new_n775_));
  NOR2_X1    g0390(.A1(new_n775_), .A2(new_n774_), .ZN(new_n776_));
  INV_X1     g0391(.I(new_n776_), .ZN(new_n777_));
  AOI21_X1   g0392(.A1(new_n767_), .A2(new_n772_), .B(new_n777_), .ZN(new_n778_));
  INV_X1     g0393(.I(\req[118] ), .ZN(new_n779_));
  NOR2_X1    g0394(.A1(new_n779_), .A2(\priority[119] ), .ZN(new_n780_));
  OR2_X2     g0395(.A1(\req[119] ), .A2(\req[120] ), .Z(new_n781_));
  NOR2_X1    g0396(.A1(new_n781_), .A2(new_n780_), .ZN(new_n782_));
  OAI21_X1   g0397(.A1(new_n778_), .A2(new_n394_), .B(new_n782_), .ZN(new_n783_));
  INV_X1     g0398(.I(\req[121] ), .ZN(new_n784_));
  NOR2_X1    g0399(.A1(new_n784_), .A2(\priority[122] ), .ZN(new_n785_));
  OR2_X2     g0400(.A1(\req[122] ), .A2(\req[123] ), .Z(new_n786_));
  NOR2_X1    g0401(.A1(new_n786_), .A2(new_n785_), .ZN(new_n787_));
  INV_X1     g0402(.I(new_n787_), .ZN(new_n788_));
  AOI21_X1   g0403(.A1(new_n783_), .A2(new_n390_), .B(new_n788_), .ZN(new_n789_));
  INV_X1     g0404(.I(\priority[125] ), .ZN(new_n790_));
  INV_X1     g0405(.I(\req[123] ), .ZN(new_n791_));
  AOI21_X1   g0406(.A1(new_n791_), .A2(\priority[123] ), .B(\priority[124] ), .ZN(new_n792_));
  NAND2_X1   g0407(.A1(new_n792_), .A2(new_n790_), .ZN(new_n793_));
  INV_X1     g0408(.I(\req[124] ), .ZN(new_n794_));
  NOR2_X1    g0409(.A1(new_n794_), .A2(\priority[125] ), .ZN(new_n795_));
  OR2_X2     g0410(.A1(\req[125] ), .A2(\req[126] ), .Z(new_n796_));
  NOR2_X1    g0411(.A1(new_n796_), .A2(new_n795_), .ZN(new_n797_));
  OAI21_X1   g0412(.A1(new_n789_), .A2(new_n793_), .B(new_n797_), .ZN(new_n798_));
  INV_X1     g0413(.I(\priority[0] ), .ZN(new_n799_));
  INV_X1     g0414(.I(\req[126] ), .ZN(new_n800_));
  AOI21_X1   g0415(.A1(new_n800_), .A2(\priority[126] ), .B(\priority[127] ), .ZN(new_n801_));
  NAND2_X1   g0416(.A1(new_n801_), .A2(new_n799_), .ZN(new_n802_));
  INV_X1     g0417(.I(new_n802_), .ZN(new_n803_));
  INV_X1     g0418(.I(\req[127] ), .ZN(new_n804_));
  OAI21_X1   g0419(.A1(new_n804_), .A2(\priority[0] ), .B(\req[0] ), .ZN(new_n805_));
  AOI21_X1   g0420(.A1(new_n798_), .A2(new_n803_), .B(new_n805_), .ZN(\grant[0] ));
  INV_X1     g0421(.I(\priority[123] ), .ZN(new_n807_));
  AOI21_X1   g0422(.A1(new_n784_), .A2(\priority[121] ), .B(\priority[122] ), .ZN(new_n808_));
  NAND2_X1   g0423(.A1(new_n808_), .A2(new_n807_), .ZN(new_n809_));
  INV_X1     g0424(.I(new_n809_), .ZN(new_n810_));
  INV_X1     g0425(.I(\priority[120] ), .ZN(new_n811_));
  AOI21_X1   g0426(.A1(new_n779_), .A2(\priority[118] ), .B(\priority[119] ), .ZN(new_n812_));
  NAND2_X1   g0427(.A1(new_n812_), .A2(new_n811_), .ZN(new_n813_));
  INV_X1     g0428(.I(\priority[114] ), .ZN(new_n814_));
  AOI21_X1   g0429(.A1(new_n763_), .A2(\priority[112] ), .B(\priority[113] ), .ZN(new_n815_));
  NAND2_X1   g0430(.A1(new_n815_), .A2(new_n814_), .ZN(new_n816_));
  INV_X1     g0431(.I(\priority[111] ), .ZN(new_n817_));
  AOI21_X1   g0432(.A1(new_n757_), .A2(\priority[109] ), .B(\priority[110] ), .ZN(new_n818_));
  NAND2_X1   g0433(.A1(new_n818_), .A2(new_n817_), .ZN(new_n819_));
  INV_X1     g0434(.I(new_n819_), .ZN(new_n820_));
  INV_X1     g0435(.I(\priority[105] ), .ZN(new_n821_));
  AOI21_X1   g0436(.A1(new_n742_), .A2(\priority[103] ), .B(\priority[104] ), .ZN(new_n822_));
  NAND2_X1   g0437(.A1(new_n822_), .A2(new_n821_), .ZN(new_n823_));
  INV_X1     g0438(.I(new_n823_), .ZN(new_n824_));
  INV_X1     g0439(.I(\priority[102] ), .ZN(new_n825_));
  AOI21_X1   g0440(.A1(new_n737_), .A2(\priority[100] ), .B(\priority[101] ), .ZN(new_n826_));
  NAND2_X1   g0441(.A1(new_n826_), .A2(new_n825_), .ZN(new_n827_));
  INV_X1     g0442(.I(\priority[96] ), .ZN(new_n828_));
  AOI21_X1   g0443(.A1(new_n721_), .A2(\priority[94] ), .B(\priority[95] ), .ZN(new_n829_));
  NAND2_X1   g0444(.A1(new_n829_), .A2(new_n828_), .ZN(new_n830_));
  INV_X1     g0445(.I(\priority[93] ), .ZN(new_n831_));
  AOI21_X1   g0446(.A1(new_n715_), .A2(\priority[91] ), .B(\priority[92] ), .ZN(new_n832_));
  NAND2_X1   g0447(.A1(new_n832_), .A2(new_n831_), .ZN(new_n833_));
  INV_X1     g0448(.I(new_n833_), .ZN(new_n834_));
  INV_X1     g0449(.I(\priority[87] ), .ZN(new_n835_));
  AOI21_X1   g0450(.A1(new_n700_), .A2(\priority[85] ), .B(\priority[86] ), .ZN(new_n836_));
  NAND2_X1   g0451(.A1(new_n836_), .A2(new_n835_), .ZN(new_n837_));
  INV_X1     g0452(.I(new_n837_), .ZN(new_n838_));
  INV_X1     g0453(.I(\priority[84] ), .ZN(new_n839_));
  AOI21_X1   g0454(.A1(new_n695_), .A2(\priority[82] ), .B(\priority[83] ), .ZN(new_n840_));
  NAND2_X1   g0455(.A1(new_n840_), .A2(new_n839_), .ZN(new_n841_));
  INV_X1     g0456(.I(\priority[78] ), .ZN(new_n842_));
  AOI21_X1   g0457(.A1(new_n679_), .A2(\priority[76] ), .B(\priority[77] ), .ZN(new_n843_));
  NAND2_X1   g0458(.A1(new_n843_), .A2(new_n842_), .ZN(new_n844_));
  INV_X1     g0459(.I(\priority[75] ), .ZN(new_n845_));
  AOI21_X1   g0460(.A1(new_n673_), .A2(\priority[73] ), .B(\priority[74] ), .ZN(new_n846_));
  NAND2_X1   g0461(.A1(new_n846_), .A2(new_n845_), .ZN(new_n847_));
  INV_X1     g0462(.I(new_n847_), .ZN(new_n848_));
  INV_X1     g0463(.I(\priority[69] ), .ZN(new_n849_));
  AOI21_X1   g0464(.A1(new_n658_), .A2(\priority[67] ), .B(\priority[68] ), .ZN(new_n850_));
  NAND2_X1   g0465(.A1(new_n850_), .A2(new_n849_), .ZN(new_n851_));
  INV_X1     g0466(.I(new_n851_), .ZN(new_n852_));
  INV_X1     g0467(.I(\priority[66] ), .ZN(new_n853_));
  AOI21_X1   g0468(.A1(new_n653_), .A2(\priority[64] ), .B(\priority[65] ), .ZN(new_n854_));
  NAND2_X1   g0469(.A1(new_n854_), .A2(new_n853_), .ZN(new_n855_));
  INV_X1     g0470(.I(\priority[60] ), .ZN(new_n856_));
  AOI21_X1   g0471(.A1(new_n637_), .A2(\priority[58] ), .B(\priority[59] ), .ZN(new_n857_));
  NAND2_X1   g0472(.A1(new_n857_), .A2(new_n856_), .ZN(new_n858_));
  INV_X1     g0473(.I(\priority[57] ), .ZN(new_n859_));
  AOI21_X1   g0474(.A1(new_n631_), .A2(\priority[55] ), .B(\priority[56] ), .ZN(new_n860_));
  NAND2_X1   g0475(.A1(new_n860_), .A2(new_n859_), .ZN(new_n861_));
  INV_X1     g0476(.I(new_n861_), .ZN(new_n862_));
  INV_X1     g0477(.I(\priority[51] ), .ZN(new_n863_));
  AOI21_X1   g0478(.A1(new_n616_), .A2(\priority[49] ), .B(\priority[50] ), .ZN(new_n864_));
  NAND2_X1   g0479(.A1(new_n864_), .A2(new_n863_), .ZN(new_n865_));
  INV_X1     g0480(.I(new_n865_), .ZN(new_n866_));
  INV_X1     g0481(.I(\priority[48] ), .ZN(new_n867_));
  AOI21_X1   g0482(.A1(new_n611_), .A2(\priority[46] ), .B(\priority[47] ), .ZN(new_n868_));
  NAND2_X1   g0483(.A1(new_n868_), .A2(new_n867_), .ZN(new_n869_));
  INV_X1     g0484(.I(\priority[42] ), .ZN(new_n870_));
  AOI21_X1   g0485(.A1(new_n595_), .A2(\priority[40] ), .B(\priority[41] ), .ZN(new_n871_));
  NAND2_X1   g0486(.A1(new_n871_), .A2(new_n870_), .ZN(new_n872_));
  INV_X1     g0487(.I(\priority[39] ), .ZN(new_n873_));
  AOI21_X1   g0488(.A1(new_n589_), .A2(\priority[37] ), .B(\priority[38] ), .ZN(new_n874_));
  NAND2_X1   g0489(.A1(new_n874_), .A2(new_n873_), .ZN(new_n875_));
  INV_X1     g0490(.I(new_n875_), .ZN(new_n876_));
  INV_X1     g0491(.I(\priority[33] ), .ZN(new_n877_));
  AOI21_X1   g0492(.A1(new_n574_), .A2(\priority[31] ), .B(\priority[32] ), .ZN(new_n878_));
  NAND2_X1   g0493(.A1(new_n878_), .A2(new_n877_), .ZN(new_n879_));
  INV_X1     g0494(.I(new_n879_), .ZN(new_n880_));
  INV_X1     g0495(.I(\priority[30] ), .ZN(new_n881_));
  AOI21_X1   g0496(.A1(new_n569_), .A2(\priority[28] ), .B(\priority[29] ), .ZN(new_n882_));
  NAND2_X1   g0497(.A1(new_n882_), .A2(new_n881_), .ZN(new_n883_));
  INV_X1     g0498(.I(\priority[24] ), .ZN(new_n884_));
  AOI21_X1   g0499(.A1(new_n553_), .A2(\priority[22] ), .B(\priority[23] ), .ZN(new_n885_));
  NAND2_X1   g0500(.A1(new_n885_), .A2(new_n884_), .ZN(new_n886_));
  INV_X1     g0501(.I(\priority[21] ), .ZN(new_n887_));
  AOI21_X1   g0502(.A1(new_n547_), .A2(\priority[19] ), .B(\priority[20] ), .ZN(new_n888_));
  NAND2_X1   g0503(.A1(new_n888_), .A2(new_n887_), .ZN(new_n889_));
  INV_X1     g0504(.I(new_n889_), .ZN(new_n890_));
  INV_X1     g0505(.I(\priority[15] ), .ZN(new_n891_));
  AOI21_X1   g0506(.A1(new_n532_), .A2(\priority[13] ), .B(\priority[14] ), .ZN(new_n892_));
  NAND2_X1   g0507(.A1(new_n892_), .A2(new_n891_), .ZN(new_n893_));
  INV_X1     g0508(.I(new_n893_), .ZN(new_n894_));
  INV_X1     g0509(.I(\priority[12] ), .ZN(new_n895_));
  AOI21_X1   g0510(.A1(new_n527_), .A2(\priority[10] ), .B(\priority[11] ), .ZN(new_n896_));
  NAND2_X1   g0511(.A1(new_n896_), .A2(new_n895_), .ZN(new_n897_));
  INV_X1     g0512(.I(\priority[6] ), .ZN(new_n898_));
  AOI21_X1   g0513(.A1(new_n511_), .A2(\priority[4] ), .B(\priority[5] ), .ZN(new_n899_));
  NAND2_X1   g0514(.A1(new_n899_), .A2(new_n898_), .ZN(new_n900_));
  INV_X1     g0515(.I(\req[2] ), .ZN(new_n901_));
  AOI21_X1   g0516(.A1(new_n901_), .A2(\priority[2] ), .B(\priority[3] ), .ZN(new_n902_));
  OR2_X2     g0517(.A1(\req[3] ), .A2(\req[4] ), .Z(new_n903_));
  NOR2_X1    g0518(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1     g0519(.I(\req[5] ), .ZN(new_n905_));
  NOR2_X1    g0520(.A1(new_n905_), .A2(\priority[6] ), .ZN(new_n906_));
  OR2_X2     g0521(.A1(\req[6] ), .A2(\req[7] ), .Z(new_n907_));
  NOR2_X1    g0522(.A1(new_n907_), .A2(new_n906_), .ZN(new_n908_));
  OAI21_X1   g0523(.A1(new_n900_), .A2(new_n904_), .B(new_n908_), .ZN(new_n909_));
  INV_X1     g0524(.I(\priority[9] ), .ZN(new_n910_));
  AOI21_X1   g0525(.A1(new_n521_), .A2(\priority[7] ), .B(\priority[8] ), .ZN(new_n911_));
  NAND2_X1   g0526(.A1(new_n911_), .A2(new_n910_), .ZN(new_n912_));
  INV_X1     g0527(.I(new_n912_), .ZN(new_n913_));
  INV_X1     g0528(.I(\req[8] ), .ZN(new_n914_));
  NOR2_X1    g0529(.A1(new_n914_), .A2(\priority[9] ), .ZN(new_n915_));
  OR2_X2     g0530(.A1(\req[9] ), .A2(\req[10] ), .Z(new_n916_));
  NOR2_X1    g0531(.A1(new_n916_), .A2(new_n915_), .ZN(new_n917_));
  INV_X1     g0532(.I(new_n917_), .ZN(new_n918_));
  AOI21_X1   g0533(.A1(new_n909_), .A2(new_n913_), .B(new_n918_), .ZN(new_n919_));
  INV_X1     g0534(.I(\req[11] ), .ZN(new_n920_));
  NOR2_X1    g0535(.A1(new_n920_), .A2(\priority[12] ), .ZN(new_n921_));
  OR2_X2     g0536(.A1(\req[12] ), .A2(\req[13] ), .Z(new_n922_));
  NOR2_X1    g0537(.A1(new_n922_), .A2(new_n921_), .ZN(new_n923_));
  OAI21_X1   g0538(.A1(new_n919_), .A2(new_n897_), .B(new_n923_), .ZN(new_n924_));
  INV_X1     g0539(.I(\req[14] ), .ZN(new_n925_));
  NOR2_X1    g0540(.A1(new_n925_), .A2(\priority[15] ), .ZN(new_n926_));
  OR2_X2     g0541(.A1(\req[15] ), .A2(\req[16] ), .Z(new_n927_));
  NOR2_X1    g0542(.A1(new_n927_), .A2(new_n926_), .ZN(new_n928_));
  INV_X1     g0543(.I(new_n928_), .ZN(new_n929_));
  AOI21_X1   g0544(.A1(new_n924_), .A2(new_n894_), .B(new_n929_), .ZN(new_n930_));
  INV_X1     g0545(.I(\priority[18] ), .ZN(new_n931_));
  AOI21_X1   g0546(.A1(new_n542_), .A2(\priority[16] ), .B(\priority[17] ), .ZN(new_n932_));
  NAND2_X1   g0547(.A1(new_n932_), .A2(new_n931_), .ZN(new_n933_));
  INV_X1     g0548(.I(\req[17] ), .ZN(new_n934_));
  NOR2_X1    g0549(.A1(new_n934_), .A2(\priority[18] ), .ZN(new_n935_));
  OR2_X2     g0550(.A1(\req[18] ), .A2(\req[19] ), .Z(new_n936_));
  NOR2_X1    g0551(.A1(new_n936_), .A2(new_n935_), .ZN(new_n937_));
  OAI21_X1   g0552(.A1(new_n930_), .A2(new_n933_), .B(new_n937_), .ZN(new_n938_));
  INV_X1     g0553(.I(\req[20] ), .ZN(new_n939_));
  NOR2_X1    g0554(.A1(new_n939_), .A2(\priority[21] ), .ZN(new_n940_));
  OR2_X2     g0555(.A1(\req[21] ), .A2(\req[22] ), .Z(new_n941_));
  NOR2_X1    g0556(.A1(new_n941_), .A2(new_n940_), .ZN(new_n942_));
  INV_X1     g0557(.I(new_n942_), .ZN(new_n943_));
  AOI21_X1   g0558(.A1(new_n938_), .A2(new_n890_), .B(new_n943_), .ZN(new_n944_));
  INV_X1     g0559(.I(\req[23] ), .ZN(new_n945_));
  NOR2_X1    g0560(.A1(new_n945_), .A2(\priority[24] ), .ZN(new_n946_));
  OR2_X2     g0561(.A1(\req[24] ), .A2(\req[25] ), .Z(new_n947_));
  NOR2_X1    g0562(.A1(new_n947_), .A2(new_n946_), .ZN(new_n948_));
  OAI21_X1   g0563(.A1(new_n944_), .A2(new_n886_), .B(new_n948_), .ZN(new_n949_));
  INV_X1     g0564(.I(\priority[27] ), .ZN(new_n950_));
  AOI21_X1   g0565(.A1(new_n563_), .A2(\priority[25] ), .B(\priority[26] ), .ZN(new_n951_));
  NAND2_X1   g0566(.A1(new_n951_), .A2(new_n950_), .ZN(new_n952_));
  INV_X1     g0567(.I(new_n952_), .ZN(new_n953_));
  INV_X1     g0568(.I(\req[26] ), .ZN(new_n954_));
  NOR2_X1    g0569(.A1(new_n954_), .A2(\priority[27] ), .ZN(new_n955_));
  OR2_X2     g0570(.A1(\req[27] ), .A2(\req[28] ), .Z(new_n956_));
  NOR2_X1    g0571(.A1(new_n956_), .A2(new_n955_), .ZN(new_n957_));
  INV_X1     g0572(.I(new_n957_), .ZN(new_n958_));
  AOI21_X1   g0573(.A1(new_n949_), .A2(new_n953_), .B(new_n958_), .ZN(new_n959_));
  INV_X1     g0574(.I(\req[29] ), .ZN(new_n960_));
  NOR2_X1    g0575(.A1(new_n960_), .A2(\priority[30] ), .ZN(new_n961_));
  OR2_X2     g0576(.A1(\req[30] ), .A2(\req[31] ), .Z(new_n962_));
  NOR2_X1    g0577(.A1(new_n962_), .A2(new_n961_), .ZN(new_n963_));
  OAI21_X1   g0578(.A1(new_n959_), .A2(new_n883_), .B(new_n963_), .ZN(new_n964_));
  INV_X1     g0579(.I(\req[32] ), .ZN(new_n965_));
  NOR2_X1    g0580(.A1(new_n965_), .A2(\priority[33] ), .ZN(new_n966_));
  OR2_X2     g0581(.A1(\req[33] ), .A2(\req[34] ), .Z(new_n967_));
  NOR2_X1    g0582(.A1(new_n967_), .A2(new_n966_), .ZN(new_n968_));
  INV_X1     g0583(.I(new_n968_), .ZN(new_n969_));
  AOI21_X1   g0584(.A1(new_n964_), .A2(new_n880_), .B(new_n969_), .ZN(new_n970_));
  INV_X1     g0585(.I(\priority[36] ), .ZN(new_n971_));
  AOI21_X1   g0586(.A1(new_n584_), .A2(\priority[34] ), .B(\priority[35] ), .ZN(new_n972_));
  NAND2_X1   g0587(.A1(new_n972_), .A2(new_n971_), .ZN(new_n973_));
  INV_X1     g0588(.I(\req[35] ), .ZN(new_n974_));
  NOR2_X1    g0589(.A1(new_n974_), .A2(\priority[36] ), .ZN(new_n975_));
  OR2_X2     g0590(.A1(\req[36] ), .A2(\req[37] ), .Z(new_n976_));
  NOR2_X1    g0591(.A1(new_n976_), .A2(new_n975_), .ZN(new_n977_));
  OAI21_X1   g0592(.A1(new_n970_), .A2(new_n973_), .B(new_n977_), .ZN(new_n978_));
  INV_X1     g0593(.I(\req[38] ), .ZN(new_n979_));
  NOR2_X1    g0594(.A1(new_n979_), .A2(\priority[39] ), .ZN(new_n980_));
  OR2_X2     g0595(.A1(\req[39] ), .A2(\req[40] ), .Z(new_n981_));
  NOR2_X1    g0596(.A1(new_n981_), .A2(new_n980_), .ZN(new_n982_));
  INV_X1     g0597(.I(new_n982_), .ZN(new_n983_));
  AOI21_X1   g0598(.A1(new_n978_), .A2(new_n876_), .B(new_n983_), .ZN(new_n984_));
  INV_X1     g0599(.I(\req[41] ), .ZN(new_n985_));
  NOR2_X1    g0600(.A1(new_n985_), .A2(\priority[42] ), .ZN(new_n986_));
  OR2_X2     g0601(.A1(\req[42] ), .A2(\req[43] ), .Z(new_n987_));
  NOR2_X1    g0602(.A1(new_n987_), .A2(new_n986_), .ZN(new_n988_));
  OAI21_X1   g0603(.A1(new_n984_), .A2(new_n872_), .B(new_n988_), .ZN(new_n989_));
  INV_X1     g0604(.I(\priority[45] ), .ZN(new_n990_));
  AOI21_X1   g0605(.A1(new_n605_), .A2(\priority[43] ), .B(\priority[44] ), .ZN(new_n991_));
  NAND2_X1   g0606(.A1(new_n991_), .A2(new_n990_), .ZN(new_n992_));
  INV_X1     g0607(.I(new_n992_), .ZN(new_n993_));
  INV_X1     g0608(.I(\req[44] ), .ZN(new_n994_));
  NOR2_X1    g0609(.A1(new_n994_), .A2(\priority[45] ), .ZN(new_n995_));
  OR2_X2     g0610(.A1(\req[45] ), .A2(\req[46] ), .Z(new_n996_));
  NOR2_X1    g0611(.A1(new_n996_), .A2(new_n995_), .ZN(new_n997_));
  INV_X1     g0612(.I(new_n997_), .ZN(new_n998_));
  AOI21_X1   g0613(.A1(new_n989_), .A2(new_n993_), .B(new_n998_), .ZN(new_n999_));
  INV_X1     g0614(.I(\req[47] ), .ZN(new_n1000_));
  NOR2_X1    g0615(.A1(new_n1000_), .A2(\priority[48] ), .ZN(new_n1001_));
  OR2_X2     g0616(.A1(\req[48] ), .A2(\req[49] ), .Z(new_n1002_));
  NOR2_X1    g0617(.A1(new_n1002_), .A2(new_n1001_), .ZN(new_n1003_));
  OAI21_X1   g0618(.A1(new_n999_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n1004_));
  INV_X1     g0619(.I(\req[50] ), .ZN(new_n1005_));
  NOR2_X1    g0620(.A1(new_n1005_), .A2(\priority[51] ), .ZN(new_n1006_));
  OR2_X2     g0621(.A1(\req[51] ), .A2(\req[52] ), .Z(new_n1007_));
  NOR2_X1    g0622(.A1(new_n1007_), .A2(new_n1006_), .ZN(new_n1008_));
  INV_X1     g0623(.I(new_n1008_), .ZN(new_n1009_));
  AOI21_X1   g0624(.A1(new_n1004_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n1010_));
  INV_X1     g0625(.I(\priority[54] ), .ZN(new_n1011_));
  AOI21_X1   g0626(.A1(new_n626_), .A2(\priority[52] ), .B(\priority[53] ), .ZN(new_n1012_));
  NAND2_X1   g0627(.A1(new_n1012_), .A2(new_n1011_), .ZN(new_n1013_));
  INV_X1     g0628(.I(\req[53] ), .ZN(new_n1014_));
  NOR2_X1    g0629(.A1(new_n1014_), .A2(\priority[54] ), .ZN(new_n1015_));
  OR2_X2     g0630(.A1(\req[54] ), .A2(\req[55] ), .Z(new_n1016_));
  NOR2_X1    g0631(.A1(new_n1016_), .A2(new_n1015_), .ZN(new_n1017_));
  OAI21_X1   g0632(.A1(new_n1010_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n1018_));
  INV_X1     g0633(.I(\req[56] ), .ZN(new_n1019_));
  NOR2_X1    g0634(.A1(new_n1019_), .A2(\priority[57] ), .ZN(new_n1020_));
  OR2_X2     g0635(.A1(\req[57] ), .A2(\req[58] ), .Z(new_n1021_));
  NOR2_X1    g0636(.A1(new_n1021_), .A2(new_n1020_), .ZN(new_n1022_));
  INV_X1     g0637(.I(new_n1022_), .ZN(new_n1023_));
  AOI21_X1   g0638(.A1(new_n1018_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n1024_));
  INV_X1     g0639(.I(\req[59] ), .ZN(new_n1025_));
  NOR2_X1    g0640(.A1(new_n1025_), .A2(\priority[60] ), .ZN(new_n1026_));
  OR2_X2     g0641(.A1(\req[60] ), .A2(\req[61] ), .Z(new_n1027_));
  NOR2_X1    g0642(.A1(new_n1027_), .A2(new_n1026_), .ZN(new_n1028_));
  OAI21_X1   g0643(.A1(new_n1024_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n1029_));
  INV_X1     g0644(.I(\priority[63] ), .ZN(new_n1030_));
  AOI21_X1   g0645(.A1(new_n647_), .A2(\priority[61] ), .B(\priority[62] ), .ZN(new_n1031_));
  NAND2_X1   g0646(.A1(new_n1031_), .A2(new_n1030_), .ZN(new_n1032_));
  INV_X1     g0647(.I(new_n1032_), .ZN(new_n1033_));
  INV_X1     g0648(.I(\req[62] ), .ZN(new_n1034_));
  NOR2_X1    g0649(.A1(new_n1034_), .A2(\priority[63] ), .ZN(new_n1035_));
  OR2_X2     g0650(.A1(\req[63] ), .A2(\req[64] ), .Z(new_n1036_));
  NOR2_X1    g0651(.A1(new_n1036_), .A2(new_n1035_), .ZN(new_n1037_));
  INV_X1     g0652(.I(new_n1037_), .ZN(new_n1038_));
  AOI21_X1   g0653(.A1(new_n1029_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n1039_));
  INV_X1     g0654(.I(\req[65] ), .ZN(new_n1040_));
  NOR2_X1    g0655(.A1(new_n1040_), .A2(\priority[66] ), .ZN(new_n1041_));
  OR2_X2     g0656(.A1(\req[66] ), .A2(\req[67] ), .Z(new_n1042_));
  NOR2_X1    g0657(.A1(new_n1042_), .A2(new_n1041_), .ZN(new_n1043_));
  OAI21_X1   g0658(.A1(new_n1039_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n1044_));
  INV_X1     g0659(.I(\req[68] ), .ZN(new_n1045_));
  NOR2_X1    g0660(.A1(new_n1045_), .A2(\priority[69] ), .ZN(new_n1046_));
  OR2_X2     g0661(.A1(\req[69] ), .A2(\req[70] ), .Z(new_n1047_));
  NOR2_X1    g0662(.A1(new_n1047_), .A2(new_n1046_), .ZN(new_n1048_));
  INV_X1     g0663(.I(new_n1048_), .ZN(new_n1049_));
  AOI21_X1   g0664(.A1(new_n1044_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n1050_));
  INV_X1     g0665(.I(\priority[72] ), .ZN(new_n1051_));
  AOI21_X1   g0666(.A1(new_n668_), .A2(\priority[70] ), .B(\priority[71] ), .ZN(new_n1052_));
  NAND2_X1   g0667(.A1(new_n1052_), .A2(new_n1051_), .ZN(new_n1053_));
  INV_X1     g0668(.I(\req[71] ), .ZN(new_n1054_));
  NOR2_X1    g0669(.A1(new_n1054_), .A2(\priority[72] ), .ZN(new_n1055_));
  OR2_X2     g0670(.A1(\req[72] ), .A2(\req[73] ), .Z(new_n1056_));
  NOR2_X1    g0671(.A1(new_n1056_), .A2(new_n1055_), .ZN(new_n1057_));
  OAI21_X1   g0672(.A1(new_n1050_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n1058_));
  INV_X1     g0673(.I(\req[74] ), .ZN(new_n1059_));
  NOR2_X1    g0674(.A1(new_n1059_), .A2(\priority[75] ), .ZN(new_n1060_));
  OR2_X2     g0675(.A1(\req[75] ), .A2(\req[76] ), .Z(new_n1061_));
  NOR2_X1    g0676(.A1(new_n1061_), .A2(new_n1060_), .ZN(new_n1062_));
  INV_X1     g0677(.I(new_n1062_), .ZN(new_n1063_));
  AOI21_X1   g0678(.A1(new_n1058_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n1064_));
  INV_X1     g0679(.I(\req[77] ), .ZN(new_n1065_));
  NOR2_X1    g0680(.A1(new_n1065_), .A2(\priority[78] ), .ZN(new_n1066_));
  OR2_X2     g0681(.A1(\req[78] ), .A2(\req[79] ), .Z(new_n1067_));
  NOR2_X1    g0682(.A1(new_n1067_), .A2(new_n1066_), .ZN(new_n1068_));
  OAI21_X1   g0683(.A1(new_n1064_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n1069_));
  INV_X1     g0684(.I(\priority[81] ), .ZN(new_n1070_));
  AOI21_X1   g0685(.A1(new_n689_), .A2(\priority[79] ), .B(\priority[80] ), .ZN(new_n1071_));
  NAND2_X1   g0686(.A1(new_n1071_), .A2(new_n1070_), .ZN(new_n1072_));
  INV_X1     g0687(.I(new_n1072_), .ZN(new_n1073_));
  INV_X1     g0688(.I(\req[80] ), .ZN(new_n1074_));
  NOR2_X1    g0689(.A1(new_n1074_), .A2(\priority[81] ), .ZN(new_n1075_));
  OR2_X2     g0690(.A1(\req[81] ), .A2(\req[82] ), .Z(new_n1076_));
  NOR2_X1    g0691(.A1(new_n1076_), .A2(new_n1075_), .ZN(new_n1077_));
  INV_X1     g0692(.I(new_n1077_), .ZN(new_n1078_));
  AOI21_X1   g0693(.A1(new_n1069_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n1079_));
  INV_X1     g0694(.I(\req[83] ), .ZN(new_n1080_));
  NOR2_X1    g0695(.A1(new_n1080_), .A2(\priority[84] ), .ZN(new_n1081_));
  OR2_X2     g0696(.A1(\req[84] ), .A2(\req[85] ), .Z(new_n1082_));
  NOR2_X1    g0697(.A1(new_n1082_), .A2(new_n1081_), .ZN(new_n1083_));
  OAI21_X1   g0698(.A1(new_n1079_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n1084_));
  INV_X1     g0699(.I(\req[86] ), .ZN(new_n1085_));
  NOR2_X1    g0700(.A1(new_n1085_), .A2(\priority[87] ), .ZN(new_n1086_));
  OR2_X2     g0701(.A1(\req[87] ), .A2(\req[88] ), .Z(new_n1087_));
  NOR2_X1    g0702(.A1(new_n1087_), .A2(new_n1086_), .ZN(new_n1088_));
  INV_X1     g0703(.I(new_n1088_), .ZN(new_n1089_));
  AOI21_X1   g0704(.A1(new_n1084_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n1090_));
  INV_X1     g0705(.I(\priority[90] ), .ZN(new_n1091_));
  AOI21_X1   g0706(.A1(new_n710_), .A2(\priority[88] ), .B(\priority[89] ), .ZN(new_n1092_));
  NAND2_X1   g0707(.A1(new_n1092_), .A2(new_n1091_), .ZN(new_n1093_));
  INV_X1     g0708(.I(\req[89] ), .ZN(new_n1094_));
  NOR2_X1    g0709(.A1(new_n1094_), .A2(\priority[90] ), .ZN(new_n1095_));
  OR2_X2     g0710(.A1(\req[90] ), .A2(\req[91] ), .Z(new_n1096_));
  NOR2_X1    g0711(.A1(new_n1096_), .A2(new_n1095_), .ZN(new_n1097_));
  OAI21_X1   g0712(.A1(new_n1090_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n1098_));
  INV_X1     g0713(.I(\req[92] ), .ZN(new_n1099_));
  NOR2_X1    g0714(.A1(new_n1099_), .A2(\priority[93] ), .ZN(new_n1100_));
  OR2_X2     g0715(.A1(\req[93] ), .A2(\req[94] ), .Z(new_n1101_));
  NOR2_X1    g0716(.A1(new_n1101_), .A2(new_n1100_), .ZN(new_n1102_));
  INV_X1     g0717(.I(new_n1102_), .ZN(new_n1103_));
  AOI21_X1   g0718(.A1(new_n1098_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n1104_));
  INV_X1     g0719(.I(\req[95] ), .ZN(new_n1105_));
  NOR2_X1    g0720(.A1(new_n1105_), .A2(\priority[96] ), .ZN(new_n1106_));
  OR2_X2     g0721(.A1(\req[96] ), .A2(\req[97] ), .Z(new_n1107_));
  NOR2_X1    g0722(.A1(new_n1107_), .A2(new_n1106_), .ZN(new_n1108_));
  OAI21_X1   g0723(.A1(new_n1104_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n1109_));
  INV_X1     g0724(.I(\priority[99] ), .ZN(new_n1110_));
  AOI21_X1   g0725(.A1(new_n731_), .A2(\priority[97] ), .B(\priority[98] ), .ZN(new_n1111_));
  NAND2_X1   g0726(.A1(new_n1111_), .A2(new_n1110_), .ZN(new_n1112_));
  INV_X1     g0727(.I(new_n1112_), .ZN(new_n1113_));
  INV_X1     g0728(.I(\req[98] ), .ZN(new_n1114_));
  NOR2_X1    g0729(.A1(new_n1114_), .A2(\priority[99] ), .ZN(new_n1115_));
  OR2_X2     g0730(.A1(\req[99] ), .A2(\req[100] ), .Z(new_n1116_));
  NOR2_X1    g0731(.A1(new_n1116_), .A2(new_n1115_), .ZN(new_n1117_));
  INV_X1     g0732(.I(new_n1117_), .ZN(new_n1118_));
  AOI21_X1   g0733(.A1(new_n1109_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n1119_));
  INV_X1     g0734(.I(\req[101] ), .ZN(new_n1120_));
  NOR2_X1    g0735(.A1(new_n1120_), .A2(\priority[102] ), .ZN(new_n1121_));
  OR2_X2     g0736(.A1(\req[102] ), .A2(\req[103] ), .Z(new_n1122_));
  NOR2_X1    g0737(.A1(new_n1122_), .A2(new_n1121_), .ZN(new_n1123_));
  OAI21_X1   g0738(.A1(new_n1119_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n1124_));
  INV_X1     g0739(.I(\req[104] ), .ZN(new_n1125_));
  NOR2_X1    g0740(.A1(new_n1125_), .A2(\priority[105] ), .ZN(new_n1126_));
  OR2_X2     g0741(.A1(\req[105] ), .A2(\req[106] ), .Z(new_n1127_));
  NOR2_X1    g0742(.A1(new_n1127_), .A2(new_n1126_), .ZN(new_n1128_));
  INV_X1     g0743(.I(new_n1128_), .ZN(new_n1129_));
  AOI21_X1   g0744(.A1(new_n1124_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n1130_));
  INV_X1     g0745(.I(\priority[108] ), .ZN(new_n1131_));
  AOI21_X1   g0746(.A1(new_n752_), .A2(\priority[106] ), .B(\priority[107] ), .ZN(new_n1132_));
  NAND2_X1   g0747(.A1(new_n1132_), .A2(new_n1131_), .ZN(new_n1133_));
  INV_X1     g0748(.I(\req[107] ), .ZN(new_n1134_));
  NOR2_X1    g0749(.A1(new_n1134_), .A2(\priority[108] ), .ZN(new_n1135_));
  OR2_X2     g0750(.A1(\req[108] ), .A2(\req[109] ), .Z(new_n1136_));
  NOR2_X1    g0751(.A1(new_n1136_), .A2(new_n1135_), .ZN(new_n1137_));
  OAI21_X1   g0752(.A1(new_n1130_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n1138_));
  INV_X1     g0753(.I(\req[110] ), .ZN(new_n1139_));
  NOR2_X1    g0754(.A1(new_n1139_), .A2(\priority[111] ), .ZN(new_n1140_));
  OR2_X2     g0755(.A1(\req[111] ), .A2(\req[112] ), .Z(new_n1141_));
  NOR2_X1    g0756(.A1(new_n1141_), .A2(new_n1140_), .ZN(new_n1142_));
  INV_X1     g0757(.I(new_n1142_), .ZN(new_n1143_));
  AOI21_X1   g0758(.A1(new_n1138_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n1144_));
  INV_X1     g0759(.I(\req[113] ), .ZN(new_n1145_));
  NOR2_X1    g0760(.A1(new_n1145_), .A2(\priority[114] ), .ZN(new_n1146_));
  OR2_X2     g0761(.A1(\req[114] ), .A2(\req[115] ), .Z(new_n1147_));
  NOR2_X1    g0762(.A1(new_n1147_), .A2(new_n1146_), .ZN(new_n1148_));
  OAI21_X1   g0763(.A1(new_n1144_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n1149_));
  INV_X1     g0764(.I(\priority[117] ), .ZN(new_n1150_));
  AOI21_X1   g0765(.A1(new_n773_), .A2(\priority[115] ), .B(\priority[116] ), .ZN(new_n1151_));
  NAND2_X1   g0766(.A1(new_n1151_), .A2(new_n1150_), .ZN(new_n1152_));
  INV_X1     g0767(.I(new_n1152_), .ZN(new_n1153_));
  INV_X1     g0768(.I(\req[116] ), .ZN(new_n1154_));
  NOR2_X1    g0769(.A1(new_n1154_), .A2(\priority[117] ), .ZN(new_n1155_));
  OR2_X2     g0770(.A1(\req[117] ), .A2(\req[118] ), .Z(new_n1156_));
  NOR2_X1    g0771(.A1(new_n1156_), .A2(new_n1155_), .ZN(new_n1157_));
  INV_X1     g0772(.I(new_n1157_), .ZN(new_n1158_));
  AOI21_X1   g0773(.A1(new_n1149_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n1159_));
  INV_X1     g0774(.I(\req[119] ), .ZN(new_n1160_));
  NOR2_X1    g0775(.A1(new_n1160_), .A2(\priority[120] ), .ZN(new_n1161_));
  OR2_X2     g0776(.A1(\req[120] ), .A2(\req[121] ), .Z(new_n1162_));
  NOR2_X1    g0777(.A1(new_n1162_), .A2(new_n1161_), .ZN(new_n1163_));
  OAI21_X1   g0778(.A1(new_n1159_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n1164_));
  INV_X1     g0779(.I(\req[122] ), .ZN(new_n1165_));
  NOR2_X1    g0780(.A1(new_n1165_), .A2(\priority[123] ), .ZN(new_n1166_));
  OR2_X2     g0781(.A1(\req[123] ), .A2(\req[124] ), .Z(new_n1167_));
  NOR2_X1    g0782(.A1(new_n1167_), .A2(new_n1166_), .ZN(new_n1168_));
  INV_X1     g0783(.I(new_n1168_), .ZN(new_n1169_));
  AOI21_X1   g0784(.A1(new_n1164_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n1170_));
  INV_X1     g0785(.I(\priority[126] ), .ZN(new_n1171_));
  AOI21_X1   g0786(.A1(new_n794_), .A2(\priority[124] ), .B(\priority[125] ), .ZN(new_n1172_));
  NAND2_X1   g0787(.A1(new_n1172_), .A2(new_n1171_), .ZN(new_n1173_));
  INV_X1     g0788(.I(\req[125] ), .ZN(new_n1174_));
  NOR2_X1    g0789(.A1(new_n1174_), .A2(\priority[126] ), .ZN(new_n1175_));
  OR2_X2     g0790(.A1(\req[126] ), .A2(\req[127] ), .Z(new_n1176_));
  NOR2_X1    g0791(.A1(new_n1176_), .A2(new_n1175_), .ZN(new_n1177_));
  OAI21_X1   g0792(.A1(new_n1170_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n1178_));
  INV_X1     g0793(.I(\priority[1] ), .ZN(new_n1179_));
  AOI21_X1   g0794(.A1(new_n804_), .A2(\priority[127] ), .B(\priority[0] ), .ZN(new_n1180_));
  NAND2_X1   g0795(.A1(new_n1180_), .A2(new_n1179_), .ZN(new_n1181_));
  INV_X1     g0796(.I(new_n1181_), .ZN(new_n1182_));
  INV_X1     g0797(.I(\req[0] ), .ZN(new_n1183_));
  OAI21_X1   g0798(.A1(new_n1183_), .A2(\priority[1] ), .B(\req[1] ), .ZN(new_n1184_));
  AOI21_X1   g0799(.A1(new_n1178_), .A2(new_n1182_), .B(new_n1184_), .ZN(\grant[1] ));
  INV_X1     g0800(.I(\priority[2] ), .ZN(new_n1186_));
  AOI21_X1   g0801(.A1(new_n1183_), .A2(\priority[0] ), .B(\priority[1] ), .ZN(new_n1187_));
  NAND2_X1   g0802(.A1(new_n1187_), .A2(new_n1186_), .ZN(new_n1188_));
  INV_X1     g0803(.I(new_n1188_), .ZN(new_n1189_));
  INV_X1     g0804(.I(\priority[124] ), .ZN(new_n1190_));
  AOI21_X1   g0805(.A1(new_n1165_), .A2(\priority[122] ), .B(\priority[123] ), .ZN(new_n1191_));
  NAND2_X1   g0806(.A1(new_n1191_), .A2(new_n1190_), .ZN(new_n1192_));
  INV_X1     g0807(.I(new_n1192_), .ZN(new_n1193_));
  INV_X1     g0808(.I(\priority[121] ), .ZN(new_n1194_));
  AOI21_X1   g0809(.A1(new_n1160_), .A2(\priority[119] ), .B(\priority[120] ), .ZN(new_n1195_));
  NAND2_X1   g0810(.A1(new_n1195_), .A2(new_n1194_), .ZN(new_n1196_));
  INV_X1     g0811(.I(\priority[115] ), .ZN(new_n1197_));
  AOI21_X1   g0812(.A1(new_n1145_), .A2(\priority[113] ), .B(\priority[114] ), .ZN(new_n1198_));
  NAND2_X1   g0813(.A1(new_n1198_), .A2(new_n1197_), .ZN(new_n1199_));
  INV_X1     g0814(.I(\priority[112] ), .ZN(new_n1200_));
  AOI21_X1   g0815(.A1(new_n1139_), .A2(\priority[110] ), .B(\priority[111] ), .ZN(new_n1201_));
  NAND2_X1   g0816(.A1(new_n1201_), .A2(new_n1200_), .ZN(new_n1202_));
  INV_X1     g0817(.I(new_n1202_), .ZN(new_n1203_));
  INV_X1     g0818(.I(\priority[106] ), .ZN(new_n1204_));
  AOI21_X1   g0819(.A1(new_n1125_), .A2(\priority[104] ), .B(\priority[105] ), .ZN(new_n1205_));
  NAND2_X1   g0820(.A1(new_n1205_), .A2(new_n1204_), .ZN(new_n1206_));
  INV_X1     g0821(.I(new_n1206_), .ZN(new_n1207_));
  INV_X1     g0822(.I(\priority[103] ), .ZN(new_n1208_));
  AOI21_X1   g0823(.A1(new_n1120_), .A2(\priority[101] ), .B(\priority[102] ), .ZN(new_n1209_));
  NAND2_X1   g0824(.A1(new_n1209_), .A2(new_n1208_), .ZN(new_n1210_));
  INV_X1     g0825(.I(\priority[97] ), .ZN(new_n1211_));
  AOI21_X1   g0826(.A1(new_n1105_), .A2(\priority[95] ), .B(\priority[96] ), .ZN(new_n1212_));
  NAND2_X1   g0827(.A1(new_n1212_), .A2(new_n1211_), .ZN(new_n1213_));
  INV_X1     g0828(.I(\priority[94] ), .ZN(new_n1214_));
  AOI21_X1   g0829(.A1(new_n1099_), .A2(\priority[92] ), .B(\priority[93] ), .ZN(new_n1215_));
  NAND2_X1   g0830(.A1(new_n1215_), .A2(new_n1214_), .ZN(new_n1216_));
  INV_X1     g0831(.I(new_n1216_), .ZN(new_n1217_));
  INV_X1     g0832(.I(\priority[88] ), .ZN(new_n1218_));
  AOI21_X1   g0833(.A1(new_n1085_), .A2(\priority[86] ), .B(\priority[87] ), .ZN(new_n1219_));
  NAND2_X1   g0834(.A1(new_n1219_), .A2(new_n1218_), .ZN(new_n1220_));
  INV_X1     g0835(.I(new_n1220_), .ZN(new_n1221_));
  INV_X1     g0836(.I(\priority[85] ), .ZN(new_n1222_));
  AOI21_X1   g0837(.A1(new_n1080_), .A2(\priority[83] ), .B(\priority[84] ), .ZN(new_n1223_));
  NAND2_X1   g0838(.A1(new_n1223_), .A2(new_n1222_), .ZN(new_n1224_));
  INV_X1     g0839(.I(\priority[79] ), .ZN(new_n1225_));
  AOI21_X1   g0840(.A1(new_n1065_), .A2(\priority[77] ), .B(\priority[78] ), .ZN(new_n1226_));
  NAND2_X1   g0841(.A1(new_n1226_), .A2(new_n1225_), .ZN(new_n1227_));
  INV_X1     g0842(.I(\priority[76] ), .ZN(new_n1228_));
  AOI21_X1   g0843(.A1(new_n1059_), .A2(\priority[74] ), .B(\priority[75] ), .ZN(new_n1229_));
  NAND2_X1   g0844(.A1(new_n1229_), .A2(new_n1228_), .ZN(new_n1230_));
  INV_X1     g0845(.I(new_n1230_), .ZN(new_n1231_));
  INV_X1     g0846(.I(\priority[70] ), .ZN(new_n1232_));
  AOI21_X1   g0847(.A1(new_n1045_), .A2(\priority[68] ), .B(\priority[69] ), .ZN(new_n1233_));
  NAND2_X1   g0848(.A1(new_n1233_), .A2(new_n1232_), .ZN(new_n1234_));
  INV_X1     g0849(.I(new_n1234_), .ZN(new_n1235_));
  INV_X1     g0850(.I(\priority[67] ), .ZN(new_n1236_));
  AOI21_X1   g0851(.A1(new_n1040_), .A2(\priority[65] ), .B(\priority[66] ), .ZN(new_n1237_));
  NAND2_X1   g0852(.A1(new_n1237_), .A2(new_n1236_), .ZN(new_n1238_));
  INV_X1     g0853(.I(\priority[61] ), .ZN(new_n1239_));
  AOI21_X1   g0854(.A1(new_n1025_), .A2(\priority[59] ), .B(\priority[60] ), .ZN(new_n1240_));
  NAND2_X1   g0855(.A1(new_n1240_), .A2(new_n1239_), .ZN(new_n1241_));
  INV_X1     g0856(.I(\priority[58] ), .ZN(new_n1242_));
  AOI21_X1   g0857(.A1(new_n1019_), .A2(\priority[56] ), .B(\priority[57] ), .ZN(new_n1243_));
  NAND2_X1   g0858(.A1(new_n1243_), .A2(new_n1242_), .ZN(new_n1244_));
  INV_X1     g0859(.I(new_n1244_), .ZN(new_n1245_));
  INV_X1     g0860(.I(\priority[52] ), .ZN(new_n1246_));
  AOI21_X1   g0861(.A1(new_n1005_), .A2(\priority[50] ), .B(\priority[51] ), .ZN(new_n1247_));
  NAND2_X1   g0862(.A1(new_n1247_), .A2(new_n1246_), .ZN(new_n1248_));
  INV_X1     g0863(.I(new_n1248_), .ZN(new_n1249_));
  INV_X1     g0864(.I(\priority[49] ), .ZN(new_n1250_));
  AOI21_X1   g0865(.A1(new_n1000_), .A2(\priority[47] ), .B(\priority[48] ), .ZN(new_n1251_));
  NAND2_X1   g0866(.A1(new_n1251_), .A2(new_n1250_), .ZN(new_n1252_));
  INV_X1     g0867(.I(\priority[43] ), .ZN(new_n1253_));
  AOI21_X1   g0868(.A1(new_n985_), .A2(\priority[41] ), .B(\priority[42] ), .ZN(new_n1254_));
  NAND2_X1   g0869(.A1(new_n1254_), .A2(new_n1253_), .ZN(new_n1255_));
  INV_X1     g0870(.I(\priority[40] ), .ZN(new_n1256_));
  AOI21_X1   g0871(.A1(new_n979_), .A2(\priority[38] ), .B(\priority[39] ), .ZN(new_n1257_));
  NAND2_X1   g0872(.A1(new_n1257_), .A2(new_n1256_), .ZN(new_n1258_));
  INV_X1     g0873(.I(new_n1258_), .ZN(new_n1259_));
  INV_X1     g0874(.I(\priority[34] ), .ZN(new_n1260_));
  AOI21_X1   g0875(.A1(new_n965_), .A2(\priority[32] ), .B(\priority[33] ), .ZN(new_n1261_));
  NAND2_X1   g0876(.A1(new_n1261_), .A2(new_n1260_), .ZN(new_n1262_));
  INV_X1     g0877(.I(new_n1262_), .ZN(new_n1263_));
  INV_X1     g0878(.I(\priority[31] ), .ZN(new_n1264_));
  AOI21_X1   g0879(.A1(new_n960_), .A2(\priority[29] ), .B(\priority[30] ), .ZN(new_n1265_));
  NAND2_X1   g0880(.A1(new_n1265_), .A2(new_n1264_), .ZN(new_n1266_));
  INV_X1     g0881(.I(\priority[25] ), .ZN(new_n1267_));
  AOI21_X1   g0882(.A1(new_n945_), .A2(\priority[23] ), .B(\priority[24] ), .ZN(new_n1268_));
  NAND2_X1   g0883(.A1(new_n1268_), .A2(new_n1267_), .ZN(new_n1269_));
  INV_X1     g0884(.I(\priority[22] ), .ZN(new_n1270_));
  AOI21_X1   g0885(.A1(new_n939_), .A2(\priority[20] ), .B(\priority[21] ), .ZN(new_n1271_));
  NAND2_X1   g0886(.A1(new_n1271_), .A2(new_n1270_), .ZN(new_n1272_));
  INV_X1     g0887(.I(new_n1272_), .ZN(new_n1273_));
  INV_X1     g0888(.I(\priority[16] ), .ZN(new_n1274_));
  AOI21_X1   g0889(.A1(new_n925_), .A2(\priority[14] ), .B(\priority[15] ), .ZN(new_n1275_));
  NAND2_X1   g0890(.A1(new_n1275_), .A2(new_n1274_), .ZN(new_n1276_));
  INV_X1     g0891(.I(new_n1276_), .ZN(new_n1277_));
  INV_X1     g0892(.I(\priority[13] ), .ZN(new_n1278_));
  AOI21_X1   g0893(.A1(new_n920_), .A2(\priority[11] ), .B(\priority[12] ), .ZN(new_n1279_));
  NAND2_X1   g0894(.A1(new_n1279_), .A2(new_n1278_), .ZN(new_n1280_));
  INV_X1     g0895(.I(\priority[7] ), .ZN(new_n1281_));
  AOI21_X1   g0896(.A1(new_n905_), .A2(\priority[5] ), .B(\priority[6] ), .ZN(new_n1282_));
  NAND2_X1   g0897(.A1(new_n1282_), .A2(new_n1281_), .ZN(new_n1283_));
  OR2_X2     g0898(.A1(\req[4] ), .A2(\req[5] ), .Z(new_n1284_));
  NOR2_X1    g0899(.A1(new_n505_), .A2(new_n1284_), .ZN(new_n1285_));
  NOR2_X1    g0900(.A1(new_n517_), .A2(\priority[7] ), .ZN(new_n1286_));
  OR2_X2     g0901(.A1(\req[7] ), .A2(\req[8] ), .Z(new_n1287_));
  NOR2_X1    g0902(.A1(new_n1287_), .A2(new_n1286_), .ZN(new_n1288_));
  OAI21_X1   g0903(.A1(new_n1283_), .A2(new_n1285_), .B(new_n1288_), .ZN(new_n1289_));
  INV_X1     g0904(.I(\priority[10] ), .ZN(new_n1290_));
  AOI21_X1   g0905(.A1(new_n914_), .A2(\priority[8] ), .B(\priority[9] ), .ZN(new_n1291_));
  NAND2_X1   g0906(.A1(new_n1291_), .A2(new_n1290_), .ZN(new_n1292_));
  INV_X1     g0907(.I(new_n1292_), .ZN(new_n1293_));
  NOR2_X1    g0908(.A1(new_n500_), .A2(\priority[10] ), .ZN(new_n1294_));
  OR2_X2     g0909(.A1(\req[10] ), .A2(\req[11] ), .Z(new_n1295_));
  NOR2_X1    g0910(.A1(new_n1295_), .A2(new_n1294_), .ZN(new_n1296_));
  INV_X1     g0911(.I(new_n1296_), .ZN(new_n1297_));
  AOI21_X1   g0912(.A1(new_n1289_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n1298_));
  NOR2_X1    g0913(.A1(new_n495_), .A2(\priority[13] ), .ZN(new_n1299_));
  OR2_X2     g0914(.A1(\req[13] ), .A2(\req[14] ), .Z(new_n1300_));
  NOR2_X1    g0915(.A1(new_n1300_), .A2(new_n1299_), .ZN(new_n1301_));
  OAI21_X1   g0916(.A1(new_n1298_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n1302_));
  NOR2_X1    g0917(.A1(new_n539_), .A2(\priority[16] ), .ZN(new_n1303_));
  OR2_X2     g0918(.A1(\req[16] ), .A2(\req[17] ), .Z(new_n1304_));
  NOR2_X1    g0919(.A1(new_n1304_), .A2(new_n1303_), .ZN(new_n1305_));
  INV_X1     g0920(.I(new_n1305_), .ZN(new_n1306_));
  AOI21_X1   g0921(.A1(new_n1302_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n1307_));
  INV_X1     g0922(.I(\priority[19] ), .ZN(new_n1308_));
  AOI21_X1   g0923(.A1(new_n934_), .A2(\priority[17] ), .B(\priority[18] ), .ZN(new_n1309_));
  NAND2_X1   g0924(.A1(new_n1309_), .A2(new_n1308_), .ZN(new_n1310_));
  NOR2_X1    g0925(.A1(new_n490_), .A2(\priority[19] ), .ZN(new_n1311_));
  OR2_X2     g0926(.A1(\req[19] ), .A2(\req[20] ), .Z(new_n1312_));
  NOR2_X1    g0927(.A1(new_n1312_), .A2(new_n1311_), .ZN(new_n1313_));
  OAI21_X1   g0928(.A1(new_n1307_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n1314_));
  NOR2_X1    g0929(.A1(new_n486_), .A2(\priority[22] ), .ZN(new_n1315_));
  OR2_X2     g0930(.A1(\req[22] ), .A2(\req[23] ), .Z(new_n1316_));
  NOR2_X1    g0931(.A1(new_n1316_), .A2(new_n1315_), .ZN(new_n1317_));
  INV_X1     g0932(.I(new_n1317_), .ZN(new_n1318_));
  AOI21_X1   g0933(.A1(new_n1314_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n1319_));
  NOR2_X1    g0934(.A1(new_n559_), .A2(\priority[25] ), .ZN(new_n1320_));
  OR2_X2     g0935(.A1(\req[25] ), .A2(\req[26] ), .Z(new_n1321_));
  NOR2_X1    g0936(.A1(new_n1321_), .A2(new_n1320_), .ZN(new_n1322_));
  OAI21_X1   g0937(.A1(new_n1319_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n1323_));
  INV_X1     g0938(.I(\priority[28] ), .ZN(new_n1324_));
  AOI21_X1   g0939(.A1(new_n954_), .A2(\priority[26] ), .B(\priority[27] ), .ZN(new_n1325_));
  NAND2_X1   g0940(.A1(new_n1325_), .A2(new_n1324_), .ZN(new_n1326_));
  INV_X1     g0941(.I(new_n1326_), .ZN(new_n1327_));
  NOR2_X1    g0942(.A1(new_n482_), .A2(\priority[28] ), .ZN(new_n1328_));
  OR2_X2     g0943(.A1(\req[28] ), .A2(\req[29] ), .Z(new_n1329_));
  NOR2_X1    g0944(.A1(new_n1329_), .A2(new_n1328_), .ZN(new_n1330_));
  INV_X1     g0945(.I(new_n1330_), .ZN(new_n1331_));
  AOI21_X1   g0946(.A1(new_n1323_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n1332_));
  NOR2_X1    g0947(.A1(new_n477_), .A2(\priority[31] ), .ZN(new_n1333_));
  OR2_X2     g0948(.A1(\req[31] ), .A2(\req[32] ), .Z(new_n1334_));
  NOR2_X1    g0949(.A1(new_n1334_), .A2(new_n1333_), .ZN(new_n1335_));
  OAI21_X1   g0950(.A1(new_n1332_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n1336_));
  NOR2_X1    g0951(.A1(new_n581_), .A2(\priority[34] ), .ZN(new_n1337_));
  OR2_X2     g0952(.A1(\req[34] ), .A2(\req[35] ), .Z(new_n1338_));
  NOR2_X1    g0953(.A1(new_n1338_), .A2(new_n1337_), .ZN(new_n1339_));
  INV_X1     g0954(.I(new_n1339_), .ZN(new_n1340_));
  AOI21_X1   g0955(.A1(new_n1336_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n1341_));
  INV_X1     g0956(.I(\priority[37] ), .ZN(new_n1342_));
  AOI21_X1   g0957(.A1(new_n974_), .A2(\priority[35] ), .B(\priority[36] ), .ZN(new_n1343_));
  NAND2_X1   g0958(.A1(new_n1343_), .A2(new_n1342_), .ZN(new_n1344_));
  NOR2_X1    g0959(.A1(new_n472_), .A2(\priority[37] ), .ZN(new_n1345_));
  OR2_X2     g0960(.A1(\req[37] ), .A2(\req[38] ), .Z(new_n1346_));
  NOR2_X1    g0961(.A1(new_n1346_), .A2(new_n1345_), .ZN(new_n1347_));
  OAI21_X1   g0962(.A1(new_n1341_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n1348_));
  NOR2_X1    g0963(.A1(new_n468_), .A2(\priority[40] ), .ZN(new_n1349_));
  OR2_X2     g0964(.A1(\req[40] ), .A2(\req[41] ), .Z(new_n1350_));
  NOR2_X1    g0965(.A1(new_n1350_), .A2(new_n1349_), .ZN(new_n1351_));
  INV_X1     g0966(.I(new_n1351_), .ZN(new_n1352_));
  AOI21_X1   g0967(.A1(new_n1348_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n1353_));
  NOR2_X1    g0968(.A1(new_n601_), .A2(\priority[43] ), .ZN(new_n1354_));
  OR2_X2     g0969(.A1(\req[43] ), .A2(\req[44] ), .Z(new_n1355_));
  NOR2_X1    g0970(.A1(new_n1355_), .A2(new_n1354_), .ZN(new_n1356_));
  OAI21_X1   g0971(.A1(new_n1353_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n1357_));
  INV_X1     g0972(.I(\priority[46] ), .ZN(new_n1358_));
  AOI21_X1   g0973(.A1(new_n994_), .A2(\priority[44] ), .B(\priority[45] ), .ZN(new_n1359_));
  NAND2_X1   g0974(.A1(new_n1359_), .A2(new_n1358_), .ZN(new_n1360_));
  INV_X1     g0975(.I(new_n1360_), .ZN(new_n1361_));
  NOR2_X1    g0976(.A1(new_n464_), .A2(\priority[46] ), .ZN(new_n1362_));
  OR2_X2     g0977(.A1(\req[46] ), .A2(\req[47] ), .Z(new_n1363_));
  NOR2_X1    g0978(.A1(new_n1363_), .A2(new_n1362_), .ZN(new_n1364_));
  INV_X1     g0979(.I(new_n1364_), .ZN(new_n1365_));
  AOI21_X1   g0980(.A1(new_n1357_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n1366_));
  NOR2_X1    g0981(.A1(new_n459_), .A2(\priority[49] ), .ZN(new_n1367_));
  OR2_X2     g0982(.A1(\req[49] ), .A2(\req[50] ), .Z(new_n1368_));
  NOR2_X1    g0983(.A1(new_n1368_), .A2(new_n1367_), .ZN(new_n1369_));
  OAI21_X1   g0984(.A1(new_n1366_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n1370_));
  NOR2_X1    g0985(.A1(new_n623_), .A2(\priority[52] ), .ZN(new_n1371_));
  OR2_X2     g0986(.A1(\req[52] ), .A2(\req[53] ), .Z(new_n1372_));
  NOR2_X1    g0987(.A1(new_n1372_), .A2(new_n1371_), .ZN(new_n1373_));
  INV_X1     g0988(.I(new_n1373_), .ZN(new_n1374_));
  AOI21_X1   g0989(.A1(new_n1370_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n1375_));
  INV_X1     g0990(.I(\priority[55] ), .ZN(new_n1376_));
  AOI21_X1   g0991(.A1(new_n1014_), .A2(\priority[53] ), .B(\priority[54] ), .ZN(new_n1377_));
  NAND2_X1   g0992(.A1(new_n1377_), .A2(new_n1376_), .ZN(new_n1378_));
  NOR2_X1    g0993(.A1(new_n454_), .A2(\priority[55] ), .ZN(new_n1379_));
  OR2_X2     g0994(.A1(\req[55] ), .A2(\req[56] ), .Z(new_n1380_));
  NOR2_X1    g0995(.A1(new_n1380_), .A2(new_n1379_), .ZN(new_n1381_));
  OAI21_X1   g0996(.A1(new_n1375_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n1382_));
  NOR2_X1    g0997(.A1(new_n450_), .A2(\priority[58] ), .ZN(new_n1383_));
  OR2_X2     g0998(.A1(\req[58] ), .A2(\req[59] ), .Z(new_n1384_));
  NOR2_X1    g0999(.A1(new_n1384_), .A2(new_n1383_), .ZN(new_n1385_));
  INV_X1     g1000(.I(new_n1385_), .ZN(new_n1386_));
  AOI21_X1   g1001(.A1(new_n1382_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n1387_));
  NOR2_X1    g1002(.A1(new_n643_), .A2(\priority[61] ), .ZN(new_n1388_));
  OR2_X2     g1003(.A1(\req[61] ), .A2(\req[62] ), .Z(new_n1389_));
  NOR2_X1    g1004(.A1(new_n1389_), .A2(new_n1388_), .ZN(new_n1390_));
  OAI21_X1   g1005(.A1(new_n1387_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n1391_));
  INV_X1     g1006(.I(\priority[64] ), .ZN(new_n1392_));
  AOI21_X1   g1007(.A1(new_n1034_), .A2(\priority[62] ), .B(\priority[63] ), .ZN(new_n1393_));
  NAND2_X1   g1008(.A1(new_n1393_), .A2(new_n1392_), .ZN(new_n1394_));
  INV_X1     g1009(.I(new_n1394_), .ZN(new_n1395_));
  NOR2_X1    g1010(.A1(new_n446_), .A2(\priority[64] ), .ZN(new_n1396_));
  OR2_X2     g1011(.A1(\req[64] ), .A2(\req[65] ), .Z(new_n1397_));
  NOR2_X1    g1012(.A1(new_n1397_), .A2(new_n1396_), .ZN(new_n1398_));
  INV_X1     g1013(.I(new_n1398_), .ZN(new_n1399_));
  AOI21_X1   g1014(.A1(new_n1391_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n1400_));
  NOR2_X1    g1015(.A1(new_n441_), .A2(\priority[67] ), .ZN(new_n1401_));
  OR2_X2     g1016(.A1(\req[67] ), .A2(\req[68] ), .Z(new_n1402_));
  NOR2_X1    g1017(.A1(new_n1402_), .A2(new_n1401_), .ZN(new_n1403_));
  OAI21_X1   g1018(.A1(new_n1400_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n1404_));
  NOR2_X1    g1019(.A1(new_n665_), .A2(\priority[70] ), .ZN(new_n1405_));
  OR2_X2     g1020(.A1(\req[70] ), .A2(\req[71] ), .Z(new_n1406_));
  NOR2_X1    g1021(.A1(new_n1406_), .A2(new_n1405_), .ZN(new_n1407_));
  INV_X1     g1022(.I(new_n1407_), .ZN(new_n1408_));
  AOI21_X1   g1023(.A1(new_n1404_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n1409_));
  INV_X1     g1024(.I(\priority[73] ), .ZN(new_n1410_));
  AOI21_X1   g1025(.A1(new_n1054_), .A2(\priority[71] ), .B(\priority[72] ), .ZN(new_n1411_));
  NAND2_X1   g1026(.A1(new_n1411_), .A2(new_n1410_), .ZN(new_n1412_));
  NOR2_X1    g1027(.A1(new_n436_), .A2(\priority[73] ), .ZN(new_n1413_));
  OR2_X2     g1028(.A1(\req[73] ), .A2(\req[74] ), .Z(new_n1414_));
  NOR2_X1    g1029(.A1(new_n1414_), .A2(new_n1413_), .ZN(new_n1415_));
  OAI21_X1   g1030(.A1(new_n1409_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n1416_));
  NOR2_X1    g1031(.A1(new_n432_), .A2(\priority[76] ), .ZN(new_n1417_));
  OR2_X2     g1032(.A1(\req[76] ), .A2(\req[77] ), .Z(new_n1418_));
  NOR2_X1    g1033(.A1(new_n1418_), .A2(new_n1417_), .ZN(new_n1419_));
  INV_X1     g1034(.I(new_n1419_), .ZN(new_n1420_));
  AOI21_X1   g1035(.A1(new_n1416_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n1421_));
  NOR2_X1    g1036(.A1(new_n685_), .A2(\priority[79] ), .ZN(new_n1422_));
  OR2_X2     g1037(.A1(\req[79] ), .A2(\req[80] ), .Z(new_n1423_));
  NOR2_X1    g1038(.A1(new_n1423_), .A2(new_n1422_), .ZN(new_n1424_));
  OAI21_X1   g1039(.A1(new_n1421_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n1425_));
  INV_X1     g1040(.I(\priority[82] ), .ZN(new_n1426_));
  AOI21_X1   g1041(.A1(new_n1074_), .A2(\priority[80] ), .B(\priority[81] ), .ZN(new_n1427_));
  NAND2_X1   g1042(.A1(new_n1427_), .A2(new_n1426_), .ZN(new_n1428_));
  INV_X1     g1043(.I(new_n1428_), .ZN(new_n1429_));
  NOR2_X1    g1044(.A1(new_n428_), .A2(\priority[82] ), .ZN(new_n1430_));
  OR2_X2     g1045(.A1(\req[82] ), .A2(\req[83] ), .Z(new_n1431_));
  NOR2_X1    g1046(.A1(new_n1431_), .A2(new_n1430_), .ZN(new_n1432_));
  INV_X1     g1047(.I(new_n1432_), .ZN(new_n1433_));
  AOI21_X1   g1048(.A1(new_n1425_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n1434_));
  NOR2_X1    g1049(.A1(new_n423_), .A2(\priority[85] ), .ZN(new_n1435_));
  OR2_X2     g1050(.A1(\req[85] ), .A2(\req[86] ), .Z(new_n1436_));
  NOR2_X1    g1051(.A1(new_n1436_), .A2(new_n1435_), .ZN(new_n1437_));
  OAI21_X1   g1052(.A1(new_n1434_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n1438_));
  NOR2_X1    g1053(.A1(new_n707_), .A2(\priority[88] ), .ZN(new_n1439_));
  OR2_X2     g1054(.A1(\req[88] ), .A2(\req[89] ), .Z(new_n1440_));
  NOR2_X1    g1055(.A1(new_n1440_), .A2(new_n1439_), .ZN(new_n1441_));
  INV_X1     g1056(.I(new_n1441_), .ZN(new_n1442_));
  AOI21_X1   g1057(.A1(new_n1438_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n1443_));
  INV_X1     g1058(.I(\priority[91] ), .ZN(new_n1444_));
  AOI21_X1   g1059(.A1(new_n1094_), .A2(\priority[89] ), .B(\priority[90] ), .ZN(new_n1445_));
  NAND2_X1   g1060(.A1(new_n1445_), .A2(new_n1444_), .ZN(new_n1446_));
  NOR2_X1    g1061(.A1(new_n418_), .A2(\priority[91] ), .ZN(new_n1447_));
  OR2_X2     g1062(.A1(\req[91] ), .A2(\req[92] ), .Z(new_n1448_));
  NOR2_X1    g1063(.A1(new_n1448_), .A2(new_n1447_), .ZN(new_n1449_));
  OAI21_X1   g1064(.A1(new_n1443_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n1450_));
  NOR2_X1    g1065(.A1(new_n414_), .A2(\priority[94] ), .ZN(new_n1451_));
  OR2_X2     g1066(.A1(\req[94] ), .A2(\req[95] ), .Z(new_n1452_));
  NOR2_X1    g1067(.A1(new_n1452_), .A2(new_n1451_), .ZN(new_n1453_));
  INV_X1     g1068(.I(new_n1453_), .ZN(new_n1454_));
  AOI21_X1   g1069(.A1(new_n1450_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n1455_));
  NOR2_X1    g1070(.A1(new_n727_), .A2(\priority[97] ), .ZN(new_n1456_));
  OR2_X2     g1071(.A1(\req[97] ), .A2(\req[98] ), .Z(new_n1457_));
  NOR2_X1    g1072(.A1(new_n1457_), .A2(new_n1456_), .ZN(new_n1458_));
  OAI21_X1   g1073(.A1(new_n1455_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n1459_));
  INV_X1     g1074(.I(\priority[100] ), .ZN(new_n1460_));
  AOI21_X1   g1075(.A1(new_n1114_), .A2(\priority[98] ), .B(\priority[99] ), .ZN(new_n1461_));
  NAND2_X1   g1076(.A1(new_n1461_), .A2(new_n1460_), .ZN(new_n1462_));
  INV_X1     g1077(.I(new_n1462_), .ZN(new_n1463_));
  NOR2_X1    g1078(.A1(new_n410_), .A2(\priority[100] ), .ZN(new_n1464_));
  OR2_X2     g1079(.A1(\req[100] ), .A2(\req[101] ), .Z(new_n1465_));
  NOR2_X1    g1080(.A1(new_n1465_), .A2(new_n1464_), .ZN(new_n1466_));
  INV_X1     g1081(.I(new_n1466_), .ZN(new_n1467_));
  AOI21_X1   g1082(.A1(new_n1459_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n1468_));
  NOR2_X1    g1083(.A1(new_n405_), .A2(\priority[103] ), .ZN(new_n1469_));
  OR2_X2     g1084(.A1(\req[103] ), .A2(\req[104] ), .Z(new_n1470_));
  NOR2_X1    g1085(.A1(new_n1470_), .A2(new_n1469_), .ZN(new_n1471_));
  OAI21_X1   g1086(.A1(new_n1468_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n1472_));
  NOR2_X1    g1087(.A1(new_n749_), .A2(\priority[106] ), .ZN(new_n1473_));
  OR2_X2     g1088(.A1(\req[106] ), .A2(\req[107] ), .Z(new_n1474_));
  NOR2_X1    g1089(.A1(new_n1474_), .A2(new_n1473_), .ZN(new_n1475_));
  INV_X1     g1090(.I(new_n1475_), .ZN(new_n1476_));
  AOI21_X1   g1091(.A1(new_n1472_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n1477_));
  INV_X1     g1092(.I(\priority[109] ), .ZN(new_n1478_));
  AOI21_X1   g1093(.A1(new_n1134_), .A2(\priority[107] ), .B(\priority[108] ), .ZN(new_n1479_));
  NAND2_X1   g1094(.A1(new_n1479_), .A2(new_n1478_), .ZN(new_n1480_));
  NOR2_X1    g1095(.A1(new_n400_), .A2(\priority[109] ), .ZN(new_n1481_));
  OR2_X2     g1096(.A1(\req[109] ), .A2(\req[110] ), .Z(new_n1482_));
  NOR2_X1    g1097(.A1(new_n1482_), .A2(new_n1481_), .ZN(new_n1483_));
  OAI21_X1   g1098(.A1(new_n1477_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n1484_));
  NOR2_X1    g1099(.A1(new_n396_), .A2(\priority[112] ), .ZN(new_n1485_));
  OR2_X2     g1100(.A1(\req[112] ), .A2(\req[113] ), .Z(new_n1486_));
  NOR2_X1    g1101(.A1(new_n1486_), .A2(new_n1485_), .ZN(new_n1487_));
  INV_X1     g1102(.I(new_n1487_), .ZN(new_n1488_));
  AOI21_X1   g1103(.A1(new_n1484_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n1489_));
  NOR2_X1    g1104(.A1(new_n769_), .A2(\priority[115] ), .ZN(new_n1490_));
  OR2_X2     g1105(.A1(\req[115] ), .A2(\req[116] ), .Z(new_n1491_));
  NOR2_X1    g1106(.A1(new_n1491_), .A2(new_n1490_), .ZN(new_n1492_));
  OAI21_X1   g1107(.A1(new_n1489_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n1493_));
  INV_X1     g1108(.I(\priority[118] ), .ZN(new_n1494_));
  AOI21_X1   g1109(.A1(new_n1154_), .A2(\priority[116] ), .B(\priority[117] ), .ZN(new_n1495_));
  NAND2_X1   g1110(.A1(new_n1495_), .A2(new_n1494_), .ZN(new_n1496_));
  INV_X1     g1111(.I(new_n1496_), .ZN(new_n1497_));
  NOR2_X1    g1112(.A1(new_n392_), .A2(\priority[118] ), .ZN(new_n1498_));
  OR2_X2     g1113(.A1(\req[118] ), .A2(\req[119] ), .Z(new_n1499_));
  NOR2_X1    g1114(.A1(new_n1499_), .A2(new_n1498_), .ZN(new_n1500_));
  INV_X1     g1115(.I(new_n1500_), .ZN(new_n1501_));
  AOI21_X1   g1116(.A1(new_n1493_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n1502_));
  NOR2_X1    g1117(.A1(new_n387_), .A2(\priority[121] ), .ZN(new_n1503_));
  OR2_X2     g1118(.A1(\req[121] ), .A2(\req[122] ), .Z(new_n1504_));
  NOR2_X1    g1119(.A1(new_n1504_), .A2(new_n1503_), .ZN(new_n1505_));
  OAI21_X1   g1120(.A1(new_n1502_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n1506_));
  NOR2_X1    g1121(.A1(new_n791_), .A2(\priority[124] ), .ZN(new_n1507_));
  OR2_X2     g1122(.A1(\req[124] ), .A2(\req[125] ), .Z(new_n1508_));
  NOR2_X1    g1123(.A1(new_n1508_), .A2(new_n1507_), .ZN(new_n1509_));
  INV_X1     g1124(.I(new_n1509_), .ZN(new_n1510_));
  AOI21_X1   g1125(.A1(new_n1506_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n1511_));
  INV_X1     g1126(.I(\priority[127] ), .ZN(new_n1512_));
  AOI21_X1   g1127(.A1(new_n1174_), .A2(\priority[125] ), .B(\priority[126] ), .ZN(new_n1513_));
  NAND2_X1   g1128(.A1(new_n1513_), .A2(new_n1512_), .ZN(new_n1514_));
  NOR2_X1    g1129(.A1(new_n800_), .A2(\priority[127] ), .ZN(new_n1515_));
  OR2_X2     g1130(.A1(\req[0] ), .A2(\req[127] ), .Z(new_n1516_));
  NOR2_X1    g1131(.A1(new_n1516_), .A2(new_n1515_), .ZN(new_n1517_));
  OAI21_X1   g1132(.A1(new_n1511_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n1518_));
  OAI21_X1   g1133(.A1(new_n507_), .A2(\priority[2] ), .B(\req[2] ), .ZN(new_n1519_));
  AOI21_X1   g1134(.A1(new_n1518_), .A2(new_n1189_), .B(new_n1519_), .ZN(\grant[2] ));
  INV_X1     g1135(.I(\priority[3] ), .ZN(new_n1521_));
  NAND2_X1   g1136(.A1(new_n508_), .A2(new_n1521_), .ZN(new_n1522_));
  INV_X1     g1137(.I(new_n1522_), .ZN(new_n1523_));
  INV_X1     g1138(.I(new_n793_), .ZN(new_n1524_));
  INV_X1     g1139(.I(new_n797_), .ZN(new_n1525_));
  INV_X1     g1140(.I(new_n394_), .ZN(new_n1526_));
  INV_X1     g1141(.I(new_n782_), .ZN(new_n1527_));
  INV_X1     g1142(.I(new_n398_), .ZN(new_n1528_));
  INV_X1     g1143(.I(new_n766_), .ZN(new_n1529_));
  INV_X1     g1144(.I(new_n751_), .ZN(new_n1530_));
  INV_X1     g1145(.I(new_n755_), .ZN(new_n1531_));
  INV_X1     g1146(.I(new_n412_), .ZN(new_n1532_));
  INV_X1     g1147(.I(new_n740_), .ZN(new_n1533_));
  INV_X1     g1148(.I(new_n416_), .ZN(new_n1534_));
  INV_X1     g1149(.I(new_n724_), .ZN(new_n1535_));
  INV_X1     g1150(.I(new_n709_), .ZN(new_n1536_));
  INV_X1     g1151(.I(new_n713_), .ZN(new_n1537_));
  INV_X1     g1152(.I(new_n430_), .ZN(new_n1538_));
  INV_X1     g1153(.I(new_n698_), .ZN(new_n1539_));
  INV_X1     g1154(.I(new_n434_), .ZN(new_n1540_));
  INV_X1     g1155(.I(new_n682_), .ZN(new_n1541_));
  INV_X1     g1156(.I(new_n667_), .ZN(new_n1542_));
  INV_X1     g1157(.I(new_n671_), .ZN(new_n1543_));
  INV_X1     g1158(.I(new_n448_), .ZN(new_n1544_));
  INV_X1     g1159(.I(new_n656_), .ZN(new_n1545_));
  INV_X1     g1160(.I(new_n452_), .ZN(new_n1546_));
  INV_X1     g1161(.I(new_n640_), .ZN(new_n1547_));
  INV_X1     g1162(.I(new_n625_), .ZN(new_n1548_));
  INV_X1     g1163(.I(new_n629_), .ZN(new_n1549_));
  INV_X1     g1164(.I(new_n466_), .ZN(new_n1550_));
  INV_X1     g1165(.I(new_n614_), .ZN(new_n1551_));
  INV_X1     g1166(.I(new_n470_), .ZN(new_n1552_));
  INV_X1     g1167(.I(new_n598_), .ZN(new_n1553_));
  INV_X1     g1168(.I(new_n583_), .ZN(new_n1554_));
  INV_X1     g1169(.I(new_n587_), .ZN(new_n1555_));
  INV_X1     g1170(.I(new_n484_), .ZN(new_n1556_));
  INV_X1     g1171(.I(new_n572_), .ZN(new_n1557_));
  INV_X1     g1172(.I(new_n488_), .ZN(new_n1558_));
  INV_X1     g1173(.I(new_n556_), .ZN(new_n1559_));
  INV_X1     g1174(.I(new_n541_), .ZN(new_n1560_));
  INV_X1     g1175(.I(new_n545_), .ZN(new_n1561_));
  INV_X1     g1176(.I(new_n502_), .ZN(new_n1562_));
  INV_X1     g1177(.I(new_n530_), .ZN(new_n1563_));
  NOR2_X1    g1178(.A1(new_n899_), .A2(new_n513_), .ZN(new_n1564_));
  OAI21_X1   g1179(.A1(new_n519_), .A2(new_n1564_), .B(new_n524_), .ZN(new_n1565_));
  AOI21_X1   g1180(.A1(new_n1565_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n1566_));
  OAI21_X1   g1181(.A1(new_n1566_), .A2(new_n497_), .B(new_n535_), .ZN(new_n1567_));
  AOI21_X1   g1182(.A1(new_n1567_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n1568_));
  OAI21_X1   g1183(.A1(new_n1568_), .A2(new_n492_), .B(new_n550_), .ZN(new_n1569_));
  AOI21_X1   g1184(.A1(new_n1569_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n1570_));
  OAI21_X1   g1185(.A1(new_n1570_), .A2(new_n561_), .B(new_n566_), .ZN(new_n1571_));
  AOI21_X1   g1186(.A1(new_n1571_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n1572_));
  OAI21_X1   g1187(.A1(new_n1572_), .A2(new_n479_), .B(new_n577_), .ZN(new_n1573_));
  AOI21_X1   g1188(.A1(new_n1573_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n1574_));
  OAI21_X1   g1189(.A1(new_n1574_), .A2(new_n474_), .B(new_n592_), .ZN(new_n1575_));
  AOI21_X1   g1190(.A1(new_n1575_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n1576_));
  OAI21_X1   g1191(.A1(new_n1576_), .A2(new_n603_), .B(new_n608_), .ZN(new_n1577_));
  AOI21_X1   g1192(.A1(new_n1577_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n1578_));
  OAI21_X1   g1193(.A1(new_n1578_), .A2(new_n461_), .B(new_n619_), .ZN(new_n1579_));
  AOI21_X1   g1194(.A1(new_n1579_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n1580_));
  OAI21_X1   g1195(.A1(new_n1580_), .A2(new_n456_), .B(new_n634_), .ZN(new_n1581_));
  AOI21_X1   g1196(.A1(new_n1581_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n1582_));
  OAI21_X1   g1197(.A1(new_n1582_), .A2(new_n645_), .B(new_n650_), .ZN(new_n1583_));
  AOI21_X1   g1198(.A1(new_n1583_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n1584_));
  OAI21_X1   g1199(.A1(new_n1584_), .A2(new_n443_), .B(new_n661_), .ZN(new_n1585_));
  AOI21_X1   g1200(.A1(new_n1585_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n1586_));
  OAI21_X1   g1201(.A1(new_n1586_), .A2(new_n438_), .B(new_n676_), .ZN(new_n1587_));
  AOI21_X1   g1202(.A1(new_n1587_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n1588_));
  OAI21_X1   g1203(.A1(new_n1588_), .A2(new_n687_), .B(new_n692_), .ZN(new_n1589_));
  AOI21_X1   g1204(.A1(new_n1589_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n1590_));
  OAI21_X1   g1205(.A1(new_n1590_), .A2(new_n425_), .B(new_n703_), .ZN(new_n1591_));
  AOI21_X1   g1206(.A1(new_n1591_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n1592_));
  OAI21_X1   g1207(.A1(new_n1592_), .A2(new_n420_), .B(new_n718_), .ZN(new_n1593_));
  AOI21_X1   g1208(.A1(new_n1593_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n1594_));
  OAI21_X1   g1209(.A1(new_n1594_), .A2(new_n729_), .B(new_n734_), .ZN(new_n1595_));
  AOI21_X1   g1210(.A1(new_n1595_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n1596_));
  OAI21_X1   g1211(.A1(new_n1596_), .A2(new_n407_), .B(new_n745_), .ZN(new_n1597_));
  AOI21_X1   g1212(.A1(new_n1597_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n1598_));
  OAI21_X1   g1213(.A1(new_n1598_), .A2(new_n402_), .B(new_n760_), .ZN(new_n1599_));
  AOI21_X1   g1214(.A1(new_n1599_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n1600_));
  OAI21_X1   g1215(.A1(new_n1600_), .A2(new_n771_), .B(new_n776_), .ZN(new_n1601_));
  AOI21_X1   g1216(.A1(new_n1601_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n1602_));
  OAI21_X1   g1217(.A1(new_n1602_), .A2(new_n389_), .B(new_n787_), .ZN(new_n1603_));
  AOI21_X1   g1218(.A1(new_n1603_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n1604_));
  NOR2_X1    g1219(.A1(new_n804_), .A2(\priority[0] ), .ZN(new_n1605_));
  OR2_X2     g1220(.A1(\req[0] ), .A2(\req[1] ), .Z(new_n1606_));
  NOR2_X1    g1221(.A1(new_n1606_), .A2(new_n1605_), .ZN(new_n1607_));
  OAI21_X1   g1222(.A1(new_n1604_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n1608_));
  OAI21_X1   g1223(.A1(new_n901_), .A2(\priority[3] ), .B(\req[3] ), .ZN(new_n1609_));
  AOI21_X1   g1224(.A1(new_n1608_), .A2(new_n1523_), .B(new_n1609_), .ZN(\grant[3] ));
  INV_X1     g1225(.I(\priority[4] ), .ZN(new_n1611_));
  NAND2_X1   g1226(.A1(new_n902_), .A2(new_n1611_), .ZN(new_n1612_));
  INV_X1     g1227(.I(new_n1612_), .ZN(new_n1613_));
  INV_X1     g1228(.I(new_n1173_), .ZN(new_n1614_));
  INV_X1     g1229(.I(new_n1177_), .ZN(new_n1615_));
  INV_X1     g1230(.I(new_n813_), .ZN(new_n1616_));
  INV_X1     g1231(.I(new_n1163_), .ZN(new_n1617_));
  INV_X1     g1232(.I(new_n816_), .ZN(new_n1618_));
  INV_X1     g1233(.I(new_n1148_), .ZN(new_n1619_));
  INV_X1     g1234(.I(new_n1133_), .ZN(new_n1620_));
  INV_X1     g1235(.I(new_n1137_), .ZN(new_n1621_));
  INV_X1     g1236(.I(new_n827_), .ZN(new_n1622_));
  INV_X1     g1237(.I(new_n1123_), .ZN(new_n1623_));
  INV_X1     g1238(.I(new_n830_), .ZN(new_n1624_));
  INV_X1     g1239(.I(new_n1108_), .ZN(new_n1625_));
  INV_X1     g1240(.I(new_n1093_), .ZN(new_n1626_));
  INV_X1     g1241(.I(new_n1097_), .ZN(new_n1627_));
  INV_X1     g1242(.I(new_n841_), .ZN(new_n1628_));
  INV_X1     g1243(.I(new_n1083_), .ZN(new_n1629_));
  INV_X1     g1244(.I(new_n844_), .ZN(new_n1630_));
  INV_X1     g1245(.I(new_n1068_), .ZN(new_n1631_));
  INV_X1     g1246(.I(new_n1053_), .ZN(new_n1632_));
  INV_X1     g1247(.I(new_n1057_), .ZN(new_n1633_));
  INV_X1     g1248(.I(new_n855_), .ZN(new_n1634_));
  INV_X1     g1249(.I(new_n1043_), .ZN(new_n1635_));
  INV_X1     g1250(.I(new_n858_), .ZN(new_n1636_));
  INV_X1     g1251(.I(new_n1028_), .ZN(new_n1637_));
  INV_X1     g1252(.I(new_n1013_), .ZN(new_n1638_));
  INV_X1     g1253(.I(new_n1017_), .ZN(new_n1639_));
  INV_X1     g1254(.I(new_n869_), .ZN(new_n1640_));
  INV_X1     g1255(.I(new_n1003_), .ZN(new_n1641_));
  INV_X1     g1256(.I(new_n872_), .ZN(new_n1642_));
  INV_X1     g1257(.I(new_n988_), .ZN(new_n1643_));
  INV_X1     g1258(.I(new_n973_), .ZN(new_n1644_));
  INV_X1     g1259(.I(new_n977_), .ZN(new_n1645_));
  INV_X1     g1260(.I(new_n883_), .ZN(new_n1646_));
  INV_X1     g1261(.I(new_n963_), .ZN(new_n1647_));
  INV_X1     g1262(.I(new_n886_), .ZN(new_n1648_));
  INV_X1     g1263(.I(new_n948_), .ZN(new_n1649_));
  INV_X1     g1264(.I(new_n933_), .ZN(new_n1650_));
  INV_X1     g1265(.I(new_n937_), .ZN(new_n1651_));
  INV_X1     g1266(.I(new_n897_), .ZN(new_n1652_));
  INV_X1     g1267(.I(new_n923_), .ZN(new_n1653_));
  NOR2_X1    g1268(.A1(new_n1282_), .A2(new_n907_), .ZN(new_n1654_));
  OAI21_X1   g1269(.A1(new_n912_), .A2(new_n1654_), .B(new_n917_), .ZN(new_n1655_));
  AOI21_X1   g1270(.A1(new_n1655_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n1656_));
  OAI21_X1   g1271(.A1(new_n1656_), .A2(new_n893_), .B(new_n928_), .ZN(new_n1657_));
  AOI21_X1   g1272(.A1(new_n1657_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n1658_));
  OAI21_X1   g1273(.A1(new_n1658_), .A2(new_n889_), .B(new_n942_), .ZN(new_n1659_));
  AOI21_X1   g1274(.A1(new_n1659_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n1660_));
  OAI21_X1   g1275(.A1(new_n1660_), .A2(new_n952_), .B(new_n957_), .ZN(new_n1661_));
  AOI21_X1   g1276(.A1(new_n1661_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n1662_));
  OAI21_X1   g1277(.A1(new_n1662_), .A2(new_n879_), .B(new_n968_), .ZN(new_n1663_));
  AOI21_X1   g1278(.A1(new_n1663_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n1664_));
  OAI21_X1   g1279(.A1(new_n1664_), .A2(new_n875_), .B(new_n982_), .ZN(new_n1665_));
  AOI21_X1   g1280(.A1(new_n1665_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n1666_));
  OAI21_X1   g1281(.A1(new_n1666_), .A2(new_n992_), .B(new_n997_), .ZN(new_n1667_));
  AOI21_X1   g1282(.A1(new_n1667_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n1668_));
  OAI21_X1   g1283(.A1(new_n1668_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n1669_));
  AOI21_X1   g1284(.A1(new_n1669_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n1670_));
  OAI21_X1   g1285(.A1(new_n1670_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n1671_));
  AOI21_X1   g1286(.A1(new_n1671_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n1672_));
  OAI21_X1   g1287(.A1(new_n1672_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n1673_));
  AOI21_X1   g1288(.A1(new_n1673_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n1674_));
  OAI21_X1   g1289(.A1(new_n1674_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n1675_));
  AOI21_X1   g1290(.A1(new_n1675_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n1676_));
  OAI21_X1   g1291(.A1(new_n1676_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n1677_));
  AOI21_X1   g1292(.A1(new_n1677_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n1678_));
  OAI21_X1   g1293(.A1(new_n1678_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n1679_));
  AOI21_X1   g1294(.A1(new_n1679_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n1680_));
  OAI21_X1   g1295(.A1(new_n1680_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n1681_));
  AOI21_X1   g1296(.A1(new_n1681_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n1682_));
  OAI21_X1   g1297(.A1(new_n1682_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n1683_));
  AOI21_X1   g1298(.A1(new_n1683_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n1684_));
  OAI21_X1   g1299(.A1(new_n1684_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n1685_));
  AOI21_X1   g1300(.A1(new_n1685_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n1686_));
  OAI21_X1   g1301(.A1(new_n1686_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n1687_));
  AOI21_X1   g1302(.A1(new_n1687_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n1688_));
  OAI21_X1   g1303(.A1(new_n1688_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n1689_));
  AOI21_X1   g1304(.A1(new_n1689_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n1690_));
  OAI21_X1   g1305(.A1(new_n1690_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n1691_));
  AOI21_X1   g1306(.A1(new_n1691_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n1692_));
  OAI21_X1   g1307(.A1(new_n1692_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n1693_));
  AOI21_X1   g1308(.A1(new_n1693_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n1694_));
  NOR2_X1    g1309(.A1(new_n1183_), .A2(\priority[1] ), .ZN(new_n1695_));
  OR2_X2     g1310(.A1(\req[1] ), .A2(\req[2] ), .Z(new_n1696_));
  NOR2_X1    g1311(.A1(new_n1696_), .A2(new_n1695_), .ZN(new_n1697_));
  OAI21_X1   g1312(.A1(new_n1694_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n1698_));
  OAI21_X1   g1313(.A1(new_n504_), .A2(\priority[4] ), .B(\req[4] ), .ZN(new_n1699_));
  AOI21_X1   g1314(.A1(new_n1698_), .A2(new_n1613_), .B(new_n1699_), .ZN(\grant[4] ));
  INV_X1     g1315(.I(new_n506_), .ZN(new_n1701_));
  INV_X1     g1316(.I(new_n1514_), .ZN(new_n1702_));
  INV_X1     g1317(.I(new_n1517_), .ZN(new_n1703_));
  INV_X1     g1318(.I(new_n1196_), .ZN(new_n1704_));
  INV_X1     g1319(.I(new_n1505_), .ZN(new_n1705_));
  INV_X1     g1320(.I(new_n1199_), .ZN(new_n1706_));
  INV_X1     g1321(.I(new_n1492_), .ZN(new_n1707_));
  INV_X1     g1322(.I(new_n1480_), .ZN(new_n1708_));
  INV_X1     g1323(.I(new_n1483_), .ZN(new_n1709_));
  INV_X1     g1324(.I(new_n1210_), .ZN(new_n1710_));
  INV_X1     g1325(.I(new_n1471_), .ZN(new_n1711_));
  INV_X1     g1326(.I(new_n1213_), .ZN(new_n1712_));
  INV_X1     g1327(.I(new_n1458_), .ZN(new_n1713_));
  INV_X1     g1328(.I(new_n1446_), .ZN(new_n1714_));
  INV_X1     g1329(.I(new_n1449_), .ZN(new_n1715_));
  INV_X1     g1330(.I(new_n1224_), .ZN(new_n1716_));
  INV_X1     g1331(.I(new_n1437_), .ZN(new_n1717_));
  INV_X1     g1332(.I(new_n1227_), .ZN(new_n1718_));
  INV_X1     g1333(.I(new_n1424_), .ZN(new_n1719_));
  INV_X1     g1334(.I(new_n1412_), .ZN(new_n1720_));
  INV_X1     g1335(.I(new_n1415_), .ZN(new_n1721_));
  INV_X1     g1336(.I(new_n1238_), .ZN(new_n1722_));
  INV_X1     g1337(.I(new_n1403_), .ZN(new_n1723_));
  INV_X1     g1338(.I(new_n1241_), .ZN(new_n1724_));
  INV_X1     g1339(.I(new_n1390_), .ZN(new_n1725_));
  INV_X1     g1340(.I(new_n1378_), .ZN(new_n1726_));
  INV_X1     g1341(.I(new_n1381_), .ZN(new_n1727_));
  INV_X1     g1342(.I(new_n1252_), .ZN(new_n1728_));
  INV_X1     g1343(.I(new_n1369_), .ZN(new_n1729_));
  INV_X1     g1344(.I(new_n1255_), .ZN(new_n1730_));
  INV_X1     g1345(.I(new_n1356_), .ZN(new_n1731_));
  INV_X1     g1346(.I(new_n1344_), .ZN(new_n1732_));
  INV_X1     g1347(.I(new_n1347_), .ZN(new_n1733_));
  INV_X1     g1348(.I(new_n1266_), .ZN(new_n1734_));
  INV_X1     g1349(.I(new_n1335_), .ZN(new_n1735_));
  INV_X1     g1350(.I(new_n1269_), .ZN(new_n1736_));
  INV_X1     g1351(.I(new_n1322_), .ZN(new_n1737_));
  INV_X1     g1352(.I(new_n1310_), .ZN(new_n1738_));
  INV_X1     g1353(.I(new_n1313_), .ZN(new_n1739_));
  INV_X1     g1354(.I(new_n1280_), .ZN(new_n1740_));
  INV_X1     g1355(.I(new_n1301_), .ZN(new_n1741_));
  NOR2_X1    g1356(.A1(new_n518_), .A2(new_n1287_), .ZN(new_n1742_));
  OAI21_X1   g1357(.A1(new_n1292_), .A2(new_n1742_), .B(new_n1296_), .ZN(new_n1743_));
  AOI21_X1   g1358(.A1(new_n1743_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n1744_));
  OAI21_X1   g1359(.A1(new_n1744_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n1745_));
  AOI21_X1   g1360(.A1(new_n1745_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n1746_));
  OAI21_X1   g1361(.A1(new_n1746_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n1747_));
  AOI21_X1   g1362(.A1(new_n1747_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n1748_));
  OAI21_X1   g1363(.A1(new_n1748_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n1749_));
  AOI21_X1   g1364(.A1(new_n1749_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n1750_));
  OAI21_X1   g1365(.A1(new_n1750_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n1751_));
  AOI21_X1   g1366(.A1(new_n1751_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n1752_));
  OAI21_X1   g1367(.A1(new_n1752_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n1753_));
  AOI21_X1   g1368(.A1(new_n1753_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n1754_));
  OAI21_X1   g1369(.A1(new_n1754_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n1755_));
  AOI21_X1   g1370(.A1(new_n1755_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n1756_));
  OAI21_X1   g1371(.A1(new_n1756_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n1757_));
  AOI21_X1   g1372(.A1(new_n1757_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n1758_));
  OAI21_X1   g1373(.A1(new_n1758_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n1759_));
  AOI21_X1   g1374(.A1(new_n1759_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n1760_));
  OAI21_X1   g1375(.A1(new_n1760_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n1761_));
  AOI21_X1   g1376(.A1(new_n1761_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n1762_));
  OAI21_X1   g1377(.A1(new_n1762_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n1763_));
  AOI21_X1   g1378(.A1(new_n1763_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n1764_));
  OAI21_X1   g1379(.A1(new_n1764_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n1765_));
  AOI21_X1   g1380(.A1(new_n1765_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n1766_));
  OAI21_X1   g1381(.A1(new_n1766_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n1767_));
  AOI21_X1   g1382(.A1(new_n1767_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n1768_));
  OAI21_X1   g1383(.A1(new_n1768_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n1769_));
  AOI21_X1   g1384(.A1(new_n1769_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n1770_));
  OAI21_X1   g1385(.A1(new_n1770_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n1771_));
  AOI21_X1   g1386(.A1(new_n1771_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n1772_));
  OAI21_X1   g1387(.A1(new_n1772_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n1773_));
  AOI21_X1   g1388(.A1(new_n1773_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n1774_));
  OAI21_X1   g1389(.A1(new_n1774_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n1775_));
  AOI21_X1   g1390(.A1(new_n1775_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n1776_));
  OAI21_X1   g1391(.A1(new_n1776_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n1777_));
  AOI21_X1   g1392(.A1(new_n1777_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n1778_));
  OAI21_X1   g1393(.A1(new_n1778_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n1779_));
  AOI21_X1   g1394(.A1(new_n1779_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n1780_));
  OAI21_X1   g1395(.A1(new_n1780_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n1781_));
  AOI21_X1   g1396(.A1(new_n1781_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n1782_));
  NOR2_X1    g1397(.A1(new_n507_), .A2(\priority[2] ), .ZN(new_n1783_));
  NOR2_X1    g1398(.A1(new_n509_), .A2(new_n1783_), .ZN(new_n1784_));
  OAI21_X1   g1399(.A1(new_n1782_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n1785_));
  OAI21_X1   g1400(.A1(new_n511_), .A2(\priority[5] ), .B(\req[5] ), .ZN(new_n1786_));
  AOI21_X1   g1401(.A1(new_n1785_), .A2(new_n1701_), .B(new_n1786_), .ZN(\grant[5] ));
  INV_X1     g1402(.I(new_n900_), .ZN(new_n1788_));
  INV_X1     g1403(.I(new_n1607_), .ZN(new_n1789_));
  NOR2_X1    g1404(.A1(new_n911_), .A2(new_n523_), .ZN(new_n1790_));
  OAI21_X1   g1405(.A1(new_n502_), .A2(new_n1790_), .B(new_n530_), .ZN(new_n1791_));
  AOI21_X1   g1406(.A1(new_n1791_), .A2(new_n498_), .B(new_n536_), .ZN(new_n1792_));
  OAI21_X1   g1407(.A1(new_n1792_), .A2(new_n541_), .B(new_n545_), .ZN(new_n1793_));
  AOI21_X1   g1408(.A1(new_n1793_), .A2(new_n493_), .B(new_n551_), .ZN(new_n1794_));
  OAI21_X1   g1409(.A1(new_n1794_), .A2(new_n488_), .B(new_n556_), .ZN(new_n1795_));
  AOI21_X1   g1410(.A1(new_n1795_), .A2(new_n562_), .B(new_n567_), .ZN(new_n1796_));
  OAI21_X1   g1411(.A1(new_n1796_), .A2(new_n484_), .B(new_n572_), .ZN(new_n1797_));
  AOI21_X1   g1412(.A1(new_n1797_), .A2(new_n480_), .B(new_n578_), .ZN(new_n1798_));
  OAI21_X1   g1413(.A1(new_n1798_), .A2(new_n583_), .B(new_n587_), .ZN(new_n1799_));
  AOI21_X1   g1414(.A1(new_n1799_), .A2(new_n475_), .B(new_n593_), .ZN(new_n1800_));
  OAI21_X1   g1415(.A1(new_n1800_), .A2(new_n470_), .B(new_n598_), .ZN(new_n1801_));
  AOI21_X1   g1416(.A1(new_n1801_), .A2(new_n604_), .B(new_n609_), .ZN(new_n1802_));
  OAI21_X1   g1417(.A1(new_n1802_), .A2(new_n466_), .B(new_n614_), .ZN(new_n1803_));
  AOI21_X1   g1418(.A1(new_n1803_), .A2(new_n462_), .B(new_n620_), .ZN(new_n1804_));
  OAI21_X1   g1419(.A1(new_n1804_), .A2(new_n625_), .B(new_n629_), .ZN(new_n1805_));
  AOI21_X1   g1420(.A1(new_n1805_), .A2(new_n457_), .B(new_n635_), .ZN(new_n1806_));
  OAI21_X1   g1421(.A1(new_n1806_), .A2(new_n452_), .B(new_n640_), .ZN(new_n1807_));
  AOI21_X1   g1422(.A1(new_n1807_), .A2(new_n646_), .B(new_n651_), .ZN(new_n1808_));
  OAI21_X1   g1423(.A1(new_n1808_), .A2(new_n448_), .B(new_n656_), .ZN(new_n1809_));
  AOI21_X1   g1424(.A1(new_n1809_), .A2(new_n444_), .B(new_n662_), .ZN(new_n1810_));
  OAI21_X1   g1425(.A1(new_n1810_), .A2(new_n667_), .B(new_n671_), .ZN(new_n1811_));
  AOI21_X1   g1426(.A1(new_n1811_), .A2(new_n439_), .B(new_n677_), .ZN(new_n1812_));
  OAI21_X1   g1427(.A1(new_n1812_), .A2(new_n434_), .B(new_n682_), .ZN(new_n1813_));
  AOI21_X1   g1428(.A1(new_n1813_), .A2(new_n688_), .B(new_n693_), .ZN(new_n1814_));
  OAI21_X1   g1429(.A1(new_n1814_), .A2(new_n430_), .B(new_n698_), .ZN(new_n1815_));
  AOI21_X1   g1430(.A1(new_n1815_), .A2(new_n426_), .B(new_n704_), .ZN(new_n1816_));
  OAI21_X1   g1431(.A1(new_n1816_), .A2(new_n709_), .B(new_n713_), .ZN(new_n1817_));
  AOI21_X1   g1432(.A1(new_n1817_), .A2(new_n421_), .B(new_n719_), .ZN(new_n1818_));
  OAI21_X1   g1433(.A1(new_n1818_), .A2(new_n416_), .B(new_n724_), .ZN(new_n1819_));
  AOI21_X1   g1434(.A1(new_n1819_), .A2(new_n730_), .B(new_n735_), .ZN(new_n1820_));
  OAI21_X1   g1435(.A1(new_n1820_), .A2(new_n412_), .B(new_n740_), .ZN(new_n1821_));
  AOI21_X1   g1436(.A1(new_n1821_), .A2(new_n408_), .B(new_n746_), .ZN(new_n1822_));
  OAI21_X1   g1437(.A1(new_n1822_), .A2(new_n751_), .B(new_n755_), .ZN(new_n1823_));
  AOI21_X1   g1438(.A1(new_n1823_), .A2(new_n403_), .B(new_n761_), .ZN(new_n1824_));
  OAI21_X1   g1439(.A1(new_n1824_), .A2(new_n398_), .B(new_n766_), .ZN(new_n1825_));
  AOI21_X1   g1440(.A1(new_n1825_), .A2(new_n772_), .B(new_n777_), .ZN(new_n1826_));
  OAI21_X1   g1441(.A1(new_n1826_), .A2(new_n394_), .B(new_n782_), .ZN(new_n1827_));
  AOI21_X1   g1442(.A1(new_n1827_), .A2(new_n390_), .B(new_n788_), .ZN(new_n1828_));
  OAI21_X1   g1443(.A1(new_n1828_), .A2(new_n793_), .B(new_n797_), .ZN(new_n1829_));
  AOI21_X1   g1444(.A1(new_n1829_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n1830_));
  NOR2_X1    g1445(.A1(new_n901_), .A2(\priority[3] ), .ZN(new_n1831_));
  NOR2_X1    g1446(.A1(new_n903_), .A2(new_n1831_), .ZN(new_n1832_));
  OAI21_X1   g1447(.A1(new_n1830_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n1833_));
  OAI21_X1   g1448(.A1(new_n905_), .A2(\priority[6] ), .B(\req[6] ), .ZN(new_n1834_));
  AOI21_X1   g1449(.A1(new_n1833_), .A2(new_n1788_), .B(new_n1834_), .ZN(\grant[6] ));
  INV_X1     g1450(.I(new_n1283_), .ZN(new_n1836_));
  INV_X1     g1451(.I(new_n1697_), .ZN(new_n1837_));
  NOR2_X1    g1452(.A1(new_n1291_), .A2(new_n916_), .ZN(new_n1838_));
  OAI21_X1   g1453(.A1(new_n897_), .A2(new_n1838_), .B(new_n923_), .ZN(new_n1839_));
  AOI21_X1   g1454(.A1(new_n1839_), .A2(new_n894_), .B(new_n929_), .ZN(new_n1840_));
  OAI21_X1   g1455(.A1(new_n1840_), .A2(new_n933_), .B(new_n937_), .ZN(new_n1841_));
  AOI21_X1   g1456(.A1(new_n1841_), .A2(new_n890_), .B(new_n943_), .ZN(new_n1842_));
  OAI21_X1   g1457(.A1(new_n1842_), .A2(new_n886_), .B(new_n948_), .ZN(new_n1843_));
  AOI21_X1   g1458(.A1(new_n1843_), .A2(new_n953_), .B(new_n958_), .ZN(new_n1844_));
  OAI21_X1   g1459(.A1(new_n1844_), .A2(new_n883_), .B(new_n963_), .ZN(new_n1845_));
  AOI21_X1   g1460(.A1(new_n1845_), .A2(new_n880_), .B(new_n969_), .ZN(new_n1846_));
  OAI21_X1   g1461(.A1(new_n1846_), .A2(new_n973_), .B(new_n977_), .ZN(new_n1847_));
  AOI21_X1   g1462(.A1(new_n1847_), .A2(new_n876_), .B(new_n983_), .ZN(new_n1848_));
  OAI21_X1   g1463(.A1(new_n1848_), .A2(new_n872_), .B(new_n988_), .ZN(new_n1849_));
  AOI21_X1   g1464(.A1(new_n1849_), .A2(new_n993_), .B(new_n998_), .ZN(new_n1850_));
  OAI21_X1   g1465(.A1(new_n1850_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n1851_));
  AOI21_X1   g1466(.A1(new_n1851_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n1852_));
  OAI21_X1   g1467(.A1(new_n1852_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n1853_));
  AOI21_X1   g1468(.A1(new_n1853_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n1854_));
  OAI21_X1   g1469(.A1(new_n1854_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n1855_));
  AOI21_X1   g1470(.A1(new_n1855_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n1856_));
  OAI21_X1   g1471(.A1(new_n1856_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n1857_));
  AOI21_X1   g1472(.A1(new_n1857_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n1858_));
  OAI21_X1   g1473(.A1(new_n1858_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n1859_));
  AOI21_X1   g1474(.A1(new_n1859_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n1860_));
  OAI21_X1   g1475(.A1(new_n1860_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n1861_));
  AOI21_X1   g1476(.A1(new_n1861_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n1862_));
  OAI21_X1   g1477(.A1(new_n1862_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n1863_));
  AOI21_X1   g1478(.A1(new_n1863_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n1864_));
  OAI21_X1   g1479(.A1(new_n1864_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n1865_));
  AOI21_X1   g1480(.A1(new_n1865_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n1866_));
  OAI21_X1   g1481(.A1(new_n1866_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n1867_));
  AOI21_X1   g1482(.A1(new_n1867_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n1868_));
  OAI21_X1   g1483(.A1(new_n1868_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n1869_));
  AOI21_X1   g1484(.A1(new_n1869_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n1870_));
  OAI21_X1   g1485(.A1(new_n1870_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n1871_));
  AOI21_X1   g1486(.A1(new_n1871_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n1872_));
  OAI21_X1   g1487(.A1(new_n1872_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n1873_));
  AOI21_X1   g1488(.A1(new_n1873_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n1874_));
  OAI21_X1   g1489(.A1(new_n1874_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n1875_));
  AOI21_X1   g1490(.A1(new_n1875_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n1876_));
  OAI21_X1   g1491(.A1(new_n1876_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n1877_));
  AOI21_X1   g1492(.A1(new_n1877_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n1878_));
  NOR2_X1    g1493(.A1(new_n504_), .A2(\priority[4] ), .ZN(new_n1879_));
  NOR2_X1    g1494(.A1(new_n1284_), .A2(new_n1879_), .ZN(new_n1880_));
  OAI21_X1   g1495(.A1(new_n1878_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n1881_));
  OAI21_X1   g1496(.A1(new_n517_), .A2(\priority[7] ), .B(\req[7] ), .ZN(new_n1882_));
  AOI21_X1   g1497(.A1(new_n1881_), .A2(new_n1836_), .B(new_n1882_), .ZN(\grant[7] ));
  INV_X1     g1498(.I(new_n1784_), .ZN(new_n1884_));
  NOR2_X1    g1499(.A1(new_n501_), .A2(new_n1295_), .ZN(new_n1885_));
  OAI21_X1   g1500(.A1(new_n1280_), .A2(new_n1885_), .B(new_n1301_), .ZN(new_n1886_));
  AOI21_X1   g1501(.A1(new_n1886_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n1887_));
  OAI21_X1   g1502(.A1(new_n1887_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n1888_));
  AOI21_X1   g1503(.A1(new_n1888_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n1889_));
  OAI21_X1   g1504(.A1(new_n1889_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n1890_));
  AOI21_X1   g1505(.A1(new_n1890_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n1891_));
  OAI21_X1   g1506(.A1(new_n1891_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n1892_));
  AOI21_X1   g1507(.A1(new_n1892_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n1893_));
  OAI21_X1   g1508(.A1(new_n1893_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n1894_));
  AOI21_X1   g1509(.A1(new_n1894_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n1895_));
  OAI21_X1   g1510(.A1(new_n1895_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n1896_));
  AOI21_X1   g1511(.A1(new_n1896_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n1897_));
  OAI21_X1   g1512(.A1(new_n1897_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n1898_));
  AOI21_X1   g1513(.A1(new_n1898_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n1899_));
  OAI21_X1   g1514(.A1(new_n1899_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n1900_));
  AOI21_X1   g1515(.A1(new_n1900_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n1901_));
  OAI21_X1   g1516(.A1(new_n1901_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n1902_));
  AOI21_X1   g1517(.A1(new_n1902_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n1903_));
  OAI21_X1   g1518(.A1(new_n1903_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n1904_));
  AOI21_X1   g1519(.A1(new_n1904_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n1905_));
  OAI21_X1   g1520(.A1(new_n1905_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n1906_));
  AOI21_X1   g1521(.A1(new_n1906_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n1907_));
  OAI21_X1   g1522(.A1(new_n1907_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n1908_));
  AOI21_X1   g1523(.A1(new_n1908_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n1909_));
  OAI21_X1   g1524(.A1(new_n1909_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n1910_));
  AOI21_X1   g1525(.A1(new_n1910_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n1911_));
  OAI21_X1   g1526(.A1(new_n1911_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n1912_));
  AOI21_X1   g1527(.A1(new_n1912_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n1913_));
  OAI21_X1   g1528(.A1(new_n1913_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n1914_));
  AOI21_X1   g1529(.A1(new_n1914_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n1915_));
  OAI21_X1   g1530(.A1(new_n1915_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n1916_));
  AOI21_X1   g1531(.A1(new_n1916_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n1917_));
  OAI21_X1   g1532(.A1(new_n1917_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n1918_));
  AOI21_X1   g1533(.A1(new_n1918_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n1919_));
  OAI21_X1   g1534(.A1(new_n1919_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n1920_));
  AOI21_X1   g1535(.A1(new_n1920_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n1921_));
  OAI21_X1   g1536(.A1(new_n1921_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n1922_));
  AOI21_X1   g1537(.A1(new_n1922_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n1923_));
  OAI21_X1   g1538(.A1(new_n1923_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n1924_));
  AOI21_X1   g1539(.A1(new_n1924_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n1925_));
  OAI21_X1   g1540(.A1(new_n1925_), .A2(new_n506_), .B(new_n514_), .ZN(new_n1926_));
  OAI21_X1   g1541(.A1(new_n521_), .A2(\priority[8] ), .B(\req[8] ), .ZN(new_n1927_));
  AOI21_X1   g1542(.A1(new_n1926_), .A2(new_n520_), .B(new_n1927_), .ZN(\grant[8] ));
  INV_X1     g1543(.I(new_n1832_), .ZN(new_n1929_));
  NOR2_X1    g1544(.A1(new_n896_), .A2(new_n529_), .ZN(new_n1930_));
  OAI21_X1   g1545(.A1(new_n497_), .A2(new_n1930_), .B(new_n535_), .ZN(new_n1931_));
  AOI21_X1   g1546(.A1(new_n1931_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n1932_));
  OAI21_X1   g1547(.A1(new_n1932_), .A2(new_n492_), .B(new_n550_), .ZN(new_n1933_));
  AOI21_X1   g1548(.A1(new_n1933_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n1934_));
  OAI21_X1   g1549(.A1(new_n1934_), .A2(new_n561_), .B(new_n566_), .ZN(new_n1935_));
  AOI21_X1   g1550(.A1(new_n1935_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n1936_));
  OAI21_X1   g1551(.A1(new_n1936_), .A2(new_n479_), .B(new_n577_), .ZN(new_n1937_));
  AOI21_X1   g1552(.A1(new_n1937_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n1938_));
  OAI21_X1   g1553(.A1(new_n1938_), .A2(new_n474_), .B(new_n592_), .ZN(new_n1939_));
  AOI21_X1   g1554(.A1(new_n1939_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n1940_));
  OAI21_X1   g1555(.A1(new_n1940_), .A2(new_n603_), .B(new_n608_), .ZN(new_n1941_));
  AOI21_X1   g1556(.A1(new_n1941_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n1942_));
  OAI21_X1   g1557(.A1(new_n1942_), .A2(new_n461_), .B(new_n619_), .ZN(new_n1943_));
  AOI21_X1   g1558(.A1(new_n1943_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n1944_));
  OAI21_X1   g1559(.A1(new_n1944_), .A2(new_n456_), .B(new_n634_), .ZN(new_n1945_));
  AOI21_X1   g1560(.A1(new_n1945_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n1946_));
  OAI21_X1   g1561(.A1(new_n1946_), .A2(new_n645_), .B(new_n650_), .ZN(new_n1947_));
  AOI21_X1   g1562(.A1(new_n1947_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n1948_));
  OAI21_X1   g1563(.A1(new_n1948_), .A2(new_n443_), .B(new_n661_), .ZN(new_n1949_));
  AOI21_X1   g1564(.A1(new_n1949_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n1950_));
  OAI21_X1   g1565(.A1(new_n1950_), .A2(new_n438_), .B(new_n676_), .ZN(new_n1951_));
  AOI21_X1   g1566(.A1(new_n1951_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n1952_));
  OAI21_X1   g1567(.A1(new_n1952_), .A2(new_n687_), .B(new_n692_), .ZN(new_n1953_));
  AOI21_X1   g1568(.A1(new_n1953_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n1954_));
  OAI21_X1   g1569(.A1(new_n1954_), .A2(new_n425_), .B(new_n703_), .ZN(new_n1955_));
  AOI21_X1   g1570(.A1(new_n1955_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n1956_));
  OAI21_X1   g1571(.A1(new_n1956_), .A2(new_n420_), .B(new_n718_), .ZN(new_n1957_));
  AOI21_X1   g1572(.A1(new_n1957_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n1958_));
  OAI21_X1   g1573(.A1(new_n1958_), .A2(new_n729_), .B(new_n734_), .ZN(new_n1959_));
  AOI21_X1   g1574(.A1(new_n1959_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n1960_));
  OAI21_X1   g1575(.A1(new_n1960_), .A2(new_n407_), .B(new_n745_), .ZN(new_n1961_));
  AOI21_X1   g1576(.A1(new_n1961_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n1962_));
  OAI21_X1   g1577(.A1(new_n1962_), .A2(new_n402_), .B(new_n760_), .ZN(new_n1963_));
  AOI21_X1   g1578(.A1(new_n1963_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n1964_));
  OAI21_X1   g1579(.A1(new_n1964_), .A2(new_n771_), .B(new_n776_), .ZN(new_n1965_));
  AOI21_X1   g1580(.A1(new_n1965_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n1966_));
  OAI21_X1   g1581(.A1(new_n1966_), .A2(new_n389_), .B(new_n787_), .ZN(new_n1967_));
  AOI21_X1   g1582(.A1(new_n1967_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n1968_));
  OAI21_X1   g1583(.A1(new_n1968_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n1969_));
  AOI21_X1   g1584(.A1(new_n1969_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n1970_));
  OAI21_X1   g1585(.A1(new_n1970_), .A2(new_n900_), .B(new_n908_), .ZN(new_n1971_));
  OAI21_X1   g1586(.A1(new_n914_), .A2(\priority[9] ), .B(\req[9] ), .ZN(new_n1972_));
  AOI21_X1   g1587(.A1(new_n1971_), .A2(new_n913_), .B(new_n1972_), .ZN(\grant[9] ));
  INV_X1     g1588(.I(new_n1880_), .ZN(new_n1974_));
  NOR2_X1    g1589(.A1(new_n1279_), .A2(new_n922_), .ZN(new_n1975_));
  OAI21_X1   g1590(.A1(new_n893_), .A2(new_n1975_), .B(new_n928_), .ZN(new_n1976_));
  AOI21_X1   g1591(.A1(new_n1976_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n1977_));
  OAI21_X1   g1592(.A1(new_n1977_), .A2(new_n889_), .B(new_n942_), .ZN(new_n1978_));
  AOI21_X1   g1593(.A1(new_n1978_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n1979_));
  OAI21_X1   g1594(.A1(new_n1979_), .A2(new_n952_), .B(new_n957_), .ZN(new_n1980_));
  AOI21_X1   g1595(.A1(new_n1980_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n1981_));
  OAI21_X1   g1596(.A1(new_n1981_), .A2(new_n879_), .B(new_n968_), .ZN(new_n1982_));
  AOI21_X1   g1597(.A1(new_n1982_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n1983_));
  OAI21_X1   g1598(.A1(new_n1983_), .A2(new_n875_), .B(new_n982_), .ZN(new_n1984_));
  AOI21_X1   g1599(.A1(new_n1984_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n1985_));
  OAI21_X1   g1600(.A1(new_n1985_), .A2(new_n992_), .B(new_n997_), .ZN(new_n1986_));
  AOI21_X1   g1601(.A1(new_n1986_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n1987_));
  OAI21_X1   g1602(.A1(new_n1987_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n1988_));
  AOI21_X1   g1603(.A1(new_n1988_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n1989_));
  OAI21_X1   g1604(.A1(new_n1989_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n1990_));
  AOI21_X1   g1605(.A1(new_n1990_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n1991_));
  OAI21_X1   g1606(.A1(new_n1991_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n1992_));
  AOI21_X1   g1607(.A1(new_n1992_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n1993_));
  OAI21_X1   g1608(.A1(new_n1993_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n1994_));
  AOI21_X1   g1609(.A1(new_n1994_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n1995_));
  OAI21_X1   g1610(.A1(new_n1995_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n1996_));
  AOI21_X1   g1611(.A1(new_n1996_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n1997_));
  OAI21_X1   g1612(.A1(new_n1997_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n1998_));
  AOI21_X1   g1613(.A1(new_n1998_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n1999_));
  OAI21_X1   g1614(.A1(new_n1999_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n2000_));
  AOI21_X1   g1615(.A1(new_n2000_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n2001_));
  OAI21_X1   g1616(.A1(new_n2001_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n2002_));
  AOI21_X1   g1617(.A1(new_n2002_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n2003_));
  OAI21_X1   g1618(.A1(new_n2003_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n2004_));
  AOI21_X1   g1619(.A1(new_n2004_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n2005_));
  OAI21_X1   g1620(.A1(new_n2005_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n2006_));
  AOI21_X1   g1621(.A1(new_n2006_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n2007_));
  OAI21_X1   g1622(.A1(new_n2007_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n2008_));
  AOI21_X1   g1623(.A1(new_n2008_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n2009_));
  OAI21_X1   g1624(.A1(new_n2009_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n2010_));
  AOI21_X1   g1625(.A1(new_n2010_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n2011_));
  OAI21_X1   g1626(.A1(new_n2011_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n2012_));
  AOI21_X1   g1627(.A1(new_n2012_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n2013_));
  OAI21_X1   g1628(.A1(new_n2013_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n2014_));
  AOI21_X1   g1629(.A1(new_n2014_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n2015_));
  OAI21_X1   g1630(.A1(new_n2015_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n2016_));
  OAI21_X1   g1631(.A1(new_n500_), .A2(\priority[10] ), .B(\req[10] ), .ZN(new_n2017_));
  AOI21_X1   g1632(.A1(new_n2016_), .A2(new_n1293_), .B(new_n2017_), .ZN(\grant[10] ));
  INV_X1     g1633(.I(new_n514_), .ZN(new_n2019_));
  NOR2_X1    g1634(.A1(new_n496_), .A2(new_n1300_), .ZN(new_n2020_));
  OAI21_X1   g1635(.A1(new_n1276_), .A2(new_n2020_), .B(new_n1305_), .ZN(new_n2021_));
  AOI21_X1   g1636(.A1(new_n2021_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n2022_));
  OAI21_X1   g1637(.A1(new_n2022_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n2023_));
  AOI21_X1   g1638(.A1(new_n2023_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n2024_));
  OAI21_X1   g1639(.A1(new_n2024_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n2025_));
  AOI21_X1   g1640(.A1(new_n2025_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n2026_));
  OAI21_X1   g1641(.A1(new_n2026_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n2027_));
  AOI21_X1   g1642(.A1(new_n2027_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n2028_));
  OAI21_X1   g1643(.A1(new_n2028_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n2029_));
  AOI21_X1   g1644(.A1(new_n2029_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n2030_));
  OAI21_X1   g1645(.A1(new_n2030_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n2031_));
  AOI21_X1   g1646(.A1(new_n2031_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n2032_));
  OAI21_X1   g1647(.A1(new_n2032_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n2033_));
  AOI21_X1   g1648(.A1(new_n2033_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n2034_));
  OAI21_X1   g1649(.A1(new_n2034_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n2035_));
  AOI21_X1   g1650(.A1(new_n2035_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n2036_));
  OAI21_X1   g1651(.A1(new_n2036_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n2037_));
  AOI21_X1   g1652(.A1(new_n2037_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n2038_));
  OAI21_X1   g1653(.A1(new_n2038_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n2039_));
  AOI21_X1   g1654(.A1(new_n2039_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n2040_));
  OAI21_X1   g1655(.A1(new_n2040_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n2041_));
  AOI21_X1   g1656(.A1(new_n2041_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n2042_));
  OAI21_X1   g1657(.A1(new_n2042_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n2043_));
  AOI21_X1   g1658(.A1(new_n2043_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n2044_));
  OAI21_X1   g1659(.A1(new_n2044_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n2045_));
  AOI21_X1   g1660(.A1(new_n2045_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n2046_));
  OAI21_X1   g1661(.A1(new_n2046_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n2047_));
  AOI21_X1   g1662(.A1(new_n2047_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n2048_));
  OAI21_X1   g1663(.A1(new_n2048_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n2049_));
  AOI21_X1   g1664(.A1(new_n2049_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n2050_));
  OAI21_X1   g1665(.A1(new_n2050_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n2051_));
  AOI21_X1   g1666(.A1(new_n2051_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n2052_));
  OAI21_X1   g1667(.A1(new_n2052_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n2053_));
  AOI21_X1   g1668(.A1(new_n2053_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n2054_));
  OAI21_X1   g1669(.A1(new_n2054_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n2055_));
  AOI21_X1   g1670(.A1(new_n2055_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n2056_));
  OAI21_X1   g1671(.A1(new_n2056_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n2057_));
  AOI21_X1   g1672(.A1(new_n2057_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n2058_));
  OAI21_X1   g1673(.A1(new_n2058_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n2059_));
  AOI21_X1   g1674(.A1(new_n2059_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n2060_));
  OAI21_X1   g1675(.A1(new_n2060_), .A2(new_n519_), .B(new_n524_), .ZN(new_n2061_));
  OAI21_X1   g1676(.A1(new_n527_), .A2(\priority[11] ), .B(\req[11] ), .ZN(new_n2062_));
  AOI21_X1   g1677(.A1(new_n2061_), .A2(new_n1562_), .B(new_n2062_), .ZN(\grant[11] ));
  INV_X1     g1678(.I(new_n908_), .ZN(new_n2064_));
  NOR2_X1    g1679(.A1(new_n892_), .A2(new_n534_), .ZN(new_n2065_));
  OAI21_X1   g1680(.A1(new_n541_), .A2(new_n2065_), .B(new_n545_), .ZN(new_n2066_));
  AOI21_X1   g1681(.A1(new_n2066_), .A2(new_n493_), .B(new_n551_), .ZN(new_n2067_));
  OAI21_X1   g1682(.A1(new_n2067_), .A2(new_n488_), .B(new_n556_), .ZN(new_n2068_));
  AOI21_X1   g1683(.A1(new_n2068_), .A2(new_n562_), .B(new_n567_), .ZN(new_n2069_));
  OAI21_X1   g1684(.A1(new_n2069_), .A2(new_n484_), .B(new_n572_), .ZN(new_n2070_));
  AOI21_X1   g1685(.A1(new_n2070_), .A2(new_n480_), .B(new_n578_), .ZN(new_n2071_));
  OAI21_X1   g1686(.A1(new_n2071_), .A2(new_n583_), .B(new_n587_), .ZN(new_n2072_));
  AOI21_X1   g1687(.A1(new_n2072_), .A2(new_n475_), .B(new_n593_), .ZN(new_n2073_));
  OAI21_X1   g1688(.A1(new_n2073_), .A2(new_n470_), .B(new_n598_), .ZN(new_n2074_));
  AOI21_X1   g1689(.A1(new_n2074_), .A2(new_n604_), .B(new_n609_), .ZN(new_n2075_));
  OAI21_X1   g1690(.A1(new_n2075_), .A2(new_n466_), .B(new_n614_), .ZN(new_n2076_));
  AOI21_X1   g1691(.A1(new_n2076_), .A2(new_n462_), .B(new_n620_), .ZN(new_n2077_));
  OAI21_X1   g1692(.A1(new_n2077_), .A2(new_n625_), .B(new_n629_), .ZN(new_n2078_));
  AOI21_X1   g1693(.A1(new_n2078_), .A2(new_n457_), .B(new_n635_), .ZN(new_n2079_));
  OAI21_X1   g1694(.A1(new_n2079_), .A2(new_n452_), .B(new_n640_), .ZN(new_n2080_));
  AOI21_X1   g1695(.A1(new_n2080_), .A2(new_n646_), .B(new_n651_), .ZN(new_n2081_));
  OAI21_X1   g1696(.A1(new_n2081_), .A2(new_n448_), .B(new_n656_), .ZN(new_n2082_));
  AOI21_X1   g1697(.A1(new_n2082_), .A2(new_n444_), .B(new_n662_), .ZN(new_n2083_));
  OAI21_X1   g1698(.A1(new_n2083_), .A2(new_n667_), .B(new_n671_), .ZN(new_n2084_));
  AOI21_X1   g1699(.A1(new_n2084_), .A2(new_n439_), .B(new_n677_), .ZN(new_n2085_));
  OAI21_X1   g1700(.A1(new_n2085_), .A2(new_n434_), .B(new_n682_), .ZN(new_n2086_));
  AOI21_X1   g1701(.A1(new_n2086_), .A2(new_n688_), .B(new_n693_), .ZN(new_n2087_));
  OAI21_X1   g1702(.A1(new_n2087_), .A2(new_n430_), .B(new_n698_), .ZN(new_n2088_));
  AOI21_X1   g1703(.A1(new_n2088_), .A2(new_n426_), .B(new_n704_), .ZN(new_n2089_));
  OAI21_X1   g1704(.A1(new_n2089_), .A2(new_n709_), .B(new_n713_), .ZN(new_n2090_));
  AOI21_X1   g1705(.A1(new_n2090_), .A2(new_n421_), .B(new_n719_), .ZN(new_n2091_));
  OAI21_X1   g1706(.A1(new_n2091_), .A2(new_n416_), .B(new_n724_), .ZN(new_n2092_));
  AOI21_X1   g1707(.A1(new_n2092_), .A2(new_n730_), .B(new_n735_), .ZN(new_n2093_));
  OAI21_X1   g1708(.A1(new_n2093_), .A2(new_n412_), .B(new_n740_), .ZN(new_n2094_));
  AOI21_X1   g1709(.A1(new_n2094_), .A2(new_n408_), .B(new_n746_), .ZN(new_n2095_));
  OAI21_X1   g1710(.A1(new_n2095_), .A2(new_n751_), .B(new_n755_), .ZN(new_n2096_));
  AOI21_X1   g1711(.A1(new_n2096_), .A2(new_n403_), .B(new_n761_), .ZN(new_n2097_));
  OAI21_X1   g1712(.A1(new_n2097_), .A2(new_n398_), .B(new_n766_), .ZN(new_n2098_));
  AOI21_X1   g1713(.A1(new_n2098_), .A2(new_n772_), .B(new_n777_), .ZN(new_n2099_));
  OAI21_X1   g1714(.A1(new_n2099_), .A2(new_n394_), .B(new_n782_), .ZN(new_n2100_));
  AOI21_X1   g1715(.A1(new_n2100_), .A2(new_n390_), .B(new_n788_), .ZN(new_n2101_));
  OAI21_X1   g1716(.A1(new_n2101_), .A2(new_n793_), .B(new_n797_), .ZN(new_n2102_));
  AOI21_X1   g1717(.A1(new_n2102_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n2103_));
  OAI21_X1   g1718(.A1(new_n2103_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n2104_));
  AOI21_X1   g1719(.A1(new_n2104_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n2105_));
  OAI21_X1   g1720(.A1(new_n2105_), .A2(new_n912_), .B(new_n917_), .ZN(new_n2106_));
  OAI21_X1   g1721(.A1(new_n920_), .A2(\priority[12] ), .B(\req[12] ), .ZN(new_n2107_));
  AOI21_X1   g1722(.A1(new_n2106_), .A2(new_n1652_), .B(new_n2107_), .ZN(\grant[12] ));
  INV_X1     g1723(.I(new_n1288_), .ZN(new_n2109_));
  NOR2_X1    g1724(.A1(new_n1275_), .A2(new_n927_), .ZN(new_n2110_));
  OAI21_X1   g1725(.A1(new_n933_), .A2(new_n2110_), .B(new_n937_), .ZN(new_n2111_));
  AOI21_X1   g1726(.A1(new_n2111_), .A2(new_n890_), .B(new_n943_), .ZN(new_n2112_));
  OAI21_X1   g1727(.A1(new_n2112_), .A2(new_n886_), .B(new_n948_), .ZN(new_n2113_));
  AOI21_X1   g1728(.A1(new_n2113_), .A2(new_n953_), .B(new_n958_), .ZN(new_n2114_));
  OAI21_X1   g1729(.A1(new_n2114_), .A2(new_n883_), .B(new_n963_), .ZN(new_n2115_));
  AOI21_X1   g1730(.A1(new_n2115_), .A2(new_n880_), .B(new_n969_), .ZN(new_n2116_));
  OAI21_X1   g1731(.A1(new_n2116_), .A2(new_n973_), .B(new_n977_), .ZN(new_n2117_));
  AOI21_X1   g1732(.A1(new_n2117_), .A2(new_n876_), .B(new_n983_), .ZN(new_n2118_));
  OAI21_X1   g1733(.A1(new_n2118_), .A2(new_n872_), .B(new_n988_), .ZN(new_n2119_));
  AOI21_X1   g1734(.A1(new_n2119_), .A2(new_n993_), .B(new_n998_), .ZN(new_n2120_));
  OAI21_X1   g1735(.A1(new_n2120_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n2121_));
  AOI21_X1   g1736(.A1(new_n2121_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n2122_));
  OAI21_X1   g1737(.A1(new_n2122_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n2123_));
  AOI21_X1   g1738(.A1(new_n2123_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n2124_));
  OAI21_X1   g1739(.A1(new_n2124_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n2125_));
  AOI21_X1   g1740(.A1(new_n2125_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n2126_));
  OAI21_X1   g1741(.A1(new_n2126_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n2127_));
  AOI21_X1   g1742(.A1(new_n2127_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n2128_));
  OAI21_X1   g1743(.A1(new_n2128_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n2129_));
  AOI21_X1   g1744(.A1(new_n2129_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n2130_));
  OAI21_X1   g1745(.A1(new_n2130_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n2131_));
  AOI21_X1   g1746(.A1(new_n2131_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n2132_));
  OAI21_X1   g1747(.A1(new_n2132_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n2133_));
  AOI21_X1   g1748(.A1(new_n2133_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n2134_));
  OAI21_X1   g1749(.A1(new_n2134_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n2135_));
  AOI21_X1   g1750(.A1(new_n2135_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n2136_));
  OAI21_X1   g1751(.A1(new_n2136_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n2137_));
  AOI21_X1   g1752(.A1(new_n2137_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n2138_));
  OAI21_X1   g1753(.A1(new_n2138_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n2139_));
  AOI21_X1   g1754(.A1(new_n2139_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n2140_));
  OAI21_X1   g1755(.A1(new_n2140_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n2141_));
  AOI21_X1   g1756(.A1(new_n2141_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n2142_));
  OAI21_X1   g1757(.A1(new_n2142_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n2143_));
  AOI21_X1   g1758(.A1(new_n2143_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n2144_));
  OAI21_X1   g1759(.A1(new_n2144_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n2145_));
  AOI21_X1   g1760(.A1(new_n2145_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n2146_));
  OAI21_X1   g1761(.A1(new_n2146_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n2147_));
  AOI21_X1   g1762(.A1(new_n2147_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n2148_));
  OAI21_X1   g1763(.A1(new_n2148_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n2149_));
  AOI21_X1   g1764(.A1(new_n2149_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n2150_));
  OAI21_X1   g1765(.A1(new_n2150_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n2151_));
  OAI21_X1   g1766(.A1(new_n495_), .A2(\priority[13] ), .B(\req[13] ), .ZN(new_n2152_));
  AOI21_X1   g1767(.A1(new_n2151_), .A2(new_n1740_), .B(new_n2152_), .ZN(\grant[13] ));
  NOR2_X1    g1768(.A1(new_n540_), .A2(new_n1304_), .ZN(new_n2154_));
  OAI21_X1   g1769(.A1(new_n1310_), .A2(new_n2154_), .B(new_n1313_), .ZN(new_n2155_));
  AOI21_X1   g1770(.A1(new_n2155_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n2156_));
  OAI21_X1   g1771(.A1(new_n2156_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n2157_));
  AOI21_X1   g1772(.A1(new_n2157_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n2158_));
  OAI21_X1   g1773(.A1(new_n2158_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n2159_));
  AOI21_X1   g1774(.A1(new_n2159_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n2160_));
  OAI21_X1   g1775(.A1(new_n2160_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n2161_));
  AOI21_X1   g1776(.A1(new_n2161_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n2162_));
  OAI21_X1   g1777(.A1(new_n2162_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n2163_));
  AOI21_X1   g1778(.A1(new_n2163_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n2164_));
  OAI21_X1   g1779(.A1(new_n2164_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n2165_));
  AOI21_X1   g1780(.A1(new_n2165_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n2166_));
  OAI21_X1   g1781(.A1(new_n2166_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n2167_));
  AOI21_X1   g1782(.A1(new_n2167_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n2168_));
  OAI21_X1   g1783(.A1(new_n2168_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n2169_));
  AOI21_X1   g1784(.A1(new_n2169_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n2170_));
  OAI21_X1   g1785(.A1(new_n2170_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n2171_));
  AOI21_X1   g1786(.A1(new_n2171_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n2172_));
  OAI21_X1   g1787(.A1(new_n2172_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n2173_));
  AOI21_X1   g1788(.A1(new_n2173_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n2174_));
  OAI21_X1   g1789(.A1(new_n2174_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n2175_));
  AOI21_X1   g1790(.A1(new_n2175_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n2176_));
  OAI21_X1   g1791(.A1(new_n2176_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n2177_));
  AOI21_X1   g1792(.A1(new_n2177_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n2178_));
  OAI21_X1   g1793(.A1(new_n2178_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n2179_));
  AOI21_X1   g1794(.A1(new_n2179_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n2180_));
  OAI21_X1   g1795(.A1(new_n2180_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n2181_));
  AOI21_X1   g1796(.A1(new_n2181_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n2182_));
  OAI21_X1   g1797(.A1(new_n2182_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n2183_));
  AOI21_X1   g1798(.A1(new_n2183_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n2184_));
  OAI21_X1   g1799(.A1(new_n2184_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n2185_));
  AOI21_X1   g1800(.A1(new_n2185_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n2186_));
  OAI21_X1   g1801(.A1(new_n2186_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n2187_));
  AOI21_X1   g1802(.A1(new_n2187_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n2188_));
  OAI21_X1   g1803(.A1(new_n2188_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n2189_));
  AOI21_X1   g1804(.A1(new_n2189_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n2190_));
  OAI21_X1   g1805(.A1(new_n2190_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n2191_));
  AOI21_X1   g1806(.A1(new_n2191_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n2192_));
  OAI21_X1   g1807(.A1(new_n2192_), .A2(new_n506_), .B(new_n514_), .ZN(new_n2193_));
  AOI21_X1   g1808(.A1(new_n2193_), .A2(new_n520_), .B(new_n525_), .ZN(new_n2194_));
  OAI21_X1   g1809(.A1(new_n2194_), .A2(new_n502_), .B(new_n530_), .ZN(new_n2195_));
  OAI21_X1   g1810(.A1(new_n532_), .A2(\priority[14] ), .B(\req[14] ), .ZN(new_n2196_));
  AOI21_X1   g1811(.A1(new_n2195_), .A2(new_n498_), .B(new_n2196_), .ZN(\grant[14] ));
  NOR2_X1    g1812(.A1(new_n932_), .A2(new_n544_), .ZN(new_n2198_));
  OAI21_X1   g1813(.A1(new_n492_), .A2(new_n2198_), .B(new_n550_), .ZN(new_n2199_));
  AOI21_X1   g1814(.A1(new_n2199_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n2200_));
  OAI21_X1   g1815(.A1(new_n2200_), .A2(new_n561_), .B(new_n566_), .ZN(new_n2201_));
  AOI21_X1   g1816(.A1(new_n2201_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n2202_));
  OAI21_X1   g1817(.A1(new_n2202_), .A2(new_n479_), .B(new_n577_), .ZN(new_n2203_));
  AOI21_X1   g1818(.A1(new_n2203_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n2204_));
  OAI21_X1   g1819(.A1(new_n2204_), .A2(new_n474_), .B(new_n592_), .ZN(new_n2205_));
  AOI21_X1   g1820(.A1(new_n2205_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n2206_));
  OAI21_X1   g1821(.A1(new_n2206_), .A2(new_n603_), .B(new_n608_), .ZN(new_n2207_));
  AOI21_X1   g1822(.A1(new_n2207_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n2208_));
  OAI21_X1   g1823(.A1(new_n2208_), .A2(new_n461_), .B(new_n619_), .ZN(new_n2209_));
  AOI21_X1   g1824(.A1(new_n2209_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n2210_));
  OAI21_X1   g1825(.A1(new_n2210_), .A2(new_n456_), .B(new_n634_), .ZN(new_n2211_));
  AOI21_X1   g1826(.A1(new_n2211_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n2212_));
  OAI21_X1   g1827(.A1(new_n2212_), .A2(new_n645_), .B(new_n650_), .ZN(new_n2213_));
  AOI21_X1   g1828(.A1(new_n2213_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n2214_));
  OAI21_X1   g1829(.A1(new_n2214_), .A2(new_n443_), .B(new_n661_), .ZN(new_n2215_));
  AOI21_X1   g1830(.A1(new_n2215_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n2216_));
  OAI21_X1   g1831(.A1(new_n2216_), .A2(new_n438_), .B(new_n676_), .ZN(new_n2217_));
  AOI21_X1   g1832(.A1(new_n2217_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n2218_));
  OAI21_X1   g1833(.A1(new_n2218_), .A2(new_n687_), .B(new_n692_), .ZN(new_n2219_));
  AOI21_X1   g1834(.A1(new_n2219_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n2220_));
  OAI21_X1   g1835(.A1(new_n2220_), .A2(new_n425_), .B(new_n703_), .ZN(new_n2221_));
  AOI21_X1   g1836(.A1(new_n2221_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n2222_));
  OAI21_X1   g1837(.A1(new_n2222_), .A2(new_n420_), .B(new_n718_), .ZN(new_n2223_));
  AOI21_X1   g1838(.A1(new_n2223_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n2224_));
  OAI21_X1   g1839(.A1(new_n2224_), .A2(new_n729_), .B(new_n734_), .ZN(new_n2225_));
  AOI21_X1   g1840(.A1(new_n2225_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n2226_));
  OAI21_X1   g1841(.A1(new_n2226_), .A2(new_n407_), .B(new_n745_), .ZN(new_n2227_));
  AOI21_X1   g1842(.A1(new_n2227_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n2228_));
  OAI21_X1   g1843(.A1(new_n2228_), .A2(new_n402_), .B(new_n760_), .ZN(new_n2229_));
  AOI21_X1   g1844(.A1(new_n2229_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n2230_));
  OAI21_X1   g1845(.A1(new_n2230_), .A2(new_n771_), .B(new_n776_), .ZN(new_n2231_));
  AOI21_X1   g1846(.A1(new_n2231_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n2232_));
  OAI21_X1   g1847(.A1(new_n2232_), .A2(new_n389_), .B(new_n787_), .ZN(new_n2233_));
  AOI21_X1   g1848(.A1(new_n2233_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n2234_));
  OAI21_X1   g1849(.A1(new_n2234_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n2235_));
  AOI21_X1   g1850(.A1(new_n2235_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n2236_));
  OAI21_X1   g1851(.A1(new_n2236_), .A2(new_n900_), .B(new_n908_), .ZN(new_n2237_));
  AOI21_X1   g1852(.A1(new_n2237_), .A2(new_n913_), .B(new_n918_), .ZN(new_n2238_));
  OAI21_X1   g1853(.A1(new_n2238_), .A2(new_n897_), .B(new_n923_), .ZN(new_n2239_));
  OAI21_X1   g1854(.A1(new_n925_), .A2(\priority[15] ), .B(\req[15] ), .ZN(new_n2240_));
  AOI21_X1   g1855(.A1(new_n2239_), .A2(new_n894_), .B(new_n2240_), .ZN(\grant[15] ));
  NOR2_X1    g1856(.A1(new_n1309_), .A2(new_n936_), .ZN(new_n2242_));
  OAI21_X1   g1857(.A1(new_n889_), .A2(new_n2242_), .B(new_n942_), .ZN(new_n2243_));
  AOI21_X1   g1858(.A1(new_n2243_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n2244_));
  OAI21_X1   g1859(.A1(new_n2244_), .A2(new_n952_), .B(new_n957_), .ZN(new_n2245_));
  AOI21_X1   g1860(.A1(new_n2245_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n2246_));
  OAI21_X1   g1861(.A1(new_n2246_), .A2(new_n879_), .B(new_n968_), .ZN(new_n2247_));
  AOI21_X1   g1862(.A1(new_n2247_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n2248_));
  OAI21_X1   g1863(.A1(new_n2248_), .A2(new_n875_), .B(new_n982_), .ZN(new_n2249_));
  AOI21_X1   g1864(.A1(new_n2249_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n2250_));
  OAI21_X1   g1865(.A1(new_n2250_), .A2(new_n992_), .B(new_n997_), .ZN(new_n2251_));
  AOI21_X1   g1866(.A1(new_n2251_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n2252_));
  OAI21_X1   g1867(.A1(new_n2252_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n2253_));
  AOI21_X1   g1868(.A1(new_n2253_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n2254_));
  OAI21_X1   g1869(.A1(new_n2254_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n2255_));
  AOI21_X1   g1870(.A1(new_n2255_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n2256_));
  OAI21_X1   g1871(.A1(new_n2256_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n2257_));
  AOI21_X1   g1872(.A1(new_n2257_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n2258_));
  OAI21_X1   g1873(.A1(new_n2258_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n2259_));
  AOI21_X1   g1874(.A1(new_n2259_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n2260_));
  OAI21_X1   g1875(.A1(new_n2260_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n2261_));
  AOI21_X1   g1876(.A1(new_n2261_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n2262_));
  OAI21_X1   g1877(.A1(new_n2262_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n2263_));
  AOI21_X1   g1878(.A1(new_n2263_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n2264_));
  OAI21_X1   g1879(.A1(new_n2264_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n2265_));
  AOI21_X1   g1880(.A1(new_n2265_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n2266_));
  OAI21_X1   g1881(.A1(new_n2266_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n2267_));
  AOI21_X1   g1882(.A1(new_n2267_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n2268_));
  OAI21_X1   g1883(.A1(new_n2268_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n2269_));
  AOI21_X1   g1884(.A1(new_n2269_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n2270_));
  OAI21_X1   g1885(.A1(new_n2270_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n2271_));
  AOI21_X1   g1886(.A1(new_n2271_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n2272_));
  OAI21_X1   g1887(.A1(new_n2272_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n2273_));
  AOI21_X1   g1888(.A1(new_n2273_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n2274_));
  OAI21_X1   g1889(.A1(new_n2274_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n2275_));
  AOI21_X1   g1890(.A1(new_n2275_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n2276_));
  OAI21_X1   g1891(.A1(new_n2276_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n2277_));
  AOI21_X1   g1892(.A1(new_n2277_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n2278_));
  OAI21_X1   g1893(.A1(new_n2278_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n2279_));
  AOI21_X1   g1894(.A1(new_n2279_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n2280_));
  OAI21_X1   g1895(.A1(new_n2280_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n2281_));
  AOI21_X1   g1896(.A1(new_n2281_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n2282_));
  OAI21_X1   g1897(.A1(new_n2282_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n2283_));
  OAI21_X1   g1898(.A1(new_n539_), .A2(\priority[16] ), .B(\req[16] ), .ZN(new_n2284_));
  AOI21_X1   g1899(.A1(new_n2283_), .A2(new_n1277_), .B(new_n2284_), .ZN(\grant[16] ));
  NOR2_X1    g1900(.A1(new_n491_), .A2(new_n1312_), .ZN(new_n2286_));
  OAI21_X1   g1901(.A1(new_n1272_), .A2(new_n2286_), .B(new_n1317_), .ZN(new_n2287_));
  AOI21_X1   g1902(.A1(new_n2287_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n2288_));
  OAI21_X1   g1903(.A1(new_n2288_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n2289_));
  AOI21_X1   g1904(.A1(new_n2289_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n2290_));
  OAI21_X1   g1905(.A1(new_n2290_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n2291_));
  AOI21_X1   g1906(.A1(new_n2291_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n2292_));
  OAI21_X1   g1907(.A1(new_n2292_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n2293_));
  AOI21_X1   g1908(.A1(new_n2293_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n2294_));
  OAI21_X1   g1909(.A1(new_n2294_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n2295_));
  AOI21_X1   g1910(.A1(new_n2295_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n2296_));
  OAI21_X1   g1911(.A1(new_n2296_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n2297_));
  AOI21_X1   g1912(.A1(new_n2297_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n2298_));
  OAI21_X1   g1913(.A1(new_n2298_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n2299_));
  AOI21_X1   g1914(.A1(new_n2299_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n2300_));
  OAI21_X1   g1915(.A1(new_n2300_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n2301_));
  AOI21_X1   g1916(.A1(new_n2301_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n2302_));
  OAI21_X1   g1917(.A1(new_n2302_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n2303_));
  AOI21_X1   g1918(.A1(new_n2303_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n2304_));
  OAI21_X1   g1919(.A1(new_n2304_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n2305_));
  AOI21_X1   g1920(.A1(new_n2305_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n2306_));
  OAI21_X1   g1921(.A1(new_n2306_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n2307_));
  AOI21_X1   g1922(.A1(new_n2307_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n2308_));
  OAI21_X1   g1923(.A1(new_n2308_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n2309_));
  AOI21_X1   g1924(.A1(new_n2309_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n2310_));
  OAI21_X1   g1925(.A1(new_n2310_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n2311_));
  AOI21_X1   g1926(.A1(new_n2311_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n2312_));
  OAI21_X1   g1927(.A1(new_n2312_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n2313_));
  AOI21_X1   g1928(.A1(new_n2313_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n2314_));
  OAI21_X1   g1929(.A1(new_n2314_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n2315_));
  AOI21_X1   g1930(.A1(new_n2315_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n2316_));
  OAI21_X1   g1931(.A1(new_n2316_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n2317_));
  AOI21_X1   g1932(.A1(new_n2317_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n2318_));
  OAI21_X1   g1933(.A1(new_n2318_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n2319_));
  AOI21_X1   g1934(.A1(new_n2319_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n2320_));
  OAI21_X1   g1935(.A1(new_n2320_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n2321_));
  AOI21_X1   g1936(.A1(new_n2321_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n2322_));
  OAI21_X1   g1937(.A1(new_n2322_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n2323_));
  AOI21_X1   g1938(.A1(new_n2323_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n2324_));
  OAI21_X1   g1939(.A1(new_n2324_), .A2(new_n519_), .B(new_n524_), .ZN(new_n2325_));
  AOI21_X1   g1940(.A1(new_n2325_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n2326_));
  OAI21_X1   g1941(.A1(new_n2326_), .A2(new_n497_), .B(new_n535_), .ZN(new_n2327_));
  OAI21_X1   g1942(.A1(new_n542_), .A2(\priority[17] ), .B(\req[17] ), .ZN(new_n2328_));
  AOI21_X1   g1943(.A1(new_n2327_), .A2(new_n1560_), .B(new_n2328_), .ZN(\grant[17] ));
  NOR2_X1    g1944(.A1(new_n888_), .A2(new_n549_), .ZN(new_n2330_));
  OAI21_X1   g1945(.A1(new_n488_), .A2(new_n2330_), .B(new_n556_), .ZN(new_n2331_));
  AOI21_X1   g1946(.A1(new_n2331_), .A2(new_n562_), .B(new_n567_), .ZN(new_n2332_));
  OAI21_X1   g1947(.A1(new_n2332_), .A2(new_n484_), .B(new_n572_), .ZN(new_n2333_));
  AOI21_X1   g1948(.A1(new_n2333_), .A2(new_n480_), .B(new_n578_), .ZN(new_n2334_));
  OAI21_X1   g1949(.A1(new_n2334_), .A2(new_n583_), .B(new_n587_), .ZN(new_n2335_));
  AOI21_X1   g1950(.A1(new_n2335_), .A2(new_n475_), .B(new_n593_), .ZN(new_n2336_));
  OAI21_X1   g1951(.A1(new_n2336_), .A2(new_n470_), .B(new_n598_), .ZN(new_n2337_));
  AOI21_X1   g1952(.A1(new_n2337_), .A2(new_n604_), .B(new_n609_), .ZN(new_n2338_));
  OAI21_X1   g1953(.A1(new_n2338_), .A2(new_n466_), .B(new_n614_), .ZN(new_n2339_));
  AOI21_X1   g1954(.A1(new_n2339_), .A2(new_n462_), .B(new_n620_), .ZN(new_n2340_));
  OAI21_X1   g1955(.A1(new_n2340_), .A2(new_n625_), .B(new_n629_), .ZN(new_n2341_));
  AOI21_X1   g1956(.A1(new_n2341_), .A2(new_n457_), .B(new_n635_), .ZN(new_n2342_));
  OAI21_X1   g1957(.A1(new_n2342_), .A2(new_n452_), .B(new_n640_), .ZN(new_n2343_));
  AOI21_X1   g1958(.A1(new_n2343_), .A2(new_n646_), .B(new_n651_), .ZN(new_n2344_));
  OAI21_X1   g1959(.A1(new_n2344_), .A2(new_n448_), .B(new_n656_), .ZN(new_n2345_));
  AOI21_X1   g1960(.A1(new_n2345_), .A2(new_n444_), .B(new_n662_), .ZN(new_n2346_));
  OAI21_X1   g1961(.A1(new_n2346_), .A2(new_n667_), .B(new_n671_), .ZN(new_n2347_));
  AOI21_X1   g1962(.A1(new_n2347_), .A2(new_n439_), .B(new_n677_), .ZN(new_n2348_));
  OAI21_X1   g1963(.A1(new_n2348_), .A2(new_n434_), .B(new_n682_), .ZN(new_n2349_));
  AOI21_X1   g1964(.A1(new_n2349_), .A2(new_n688_), .B(new_n693_), .ZN(new_n2350_));
  OAI21_X1   g1965(.A1(new_n2350_), .A2(new_n430_), .B(new_n698_), .ZN(new_n2351_));
  AOI21_X1   g1966(.A1(new_n2351_), .A2(new_n426_), .B(new_n704_), .ZN(new_n2352_));
  OAI21_X1   g1967(.A1(new_n2352_), .A2(new_n709_), .B(new_n713_), .ZN(new_n2353_));
  AOI21_X1   g1968(.A1(new_n2353_), .A2(new_n421_), .B(new_n719_), .ZN(new_n2354_));
  OAI21_X1   g1969(.A1(new_n2354_), .A2(new_n416_), .B(new_n724_), .ZN(new_n2355_));
  AOI21_X1   g1970(.A1(new_n2355_), .A2(new_n730_), .B(new_n735_), .ZN(new_n2356_));
  OAI21_X1   g1971(.A1(new_n2356_), .A2(new_n412_), .B(new_n740_), .ZN(new_n2357_));
  AOI21_X1   g1972(.A1(new_n2357_), .A2(new_n408_), .B(new_n746_), .ZN(new_n2358_));
  OAI21_X1   g1973(.A1(new_n2358_), .A2(new_n751_), .B(new_n755_), .ZN(new_n2359_));
  AOI21_X1   g1974(.A1(new_n2359_), .A2(new_n403_), .B(new_n761_), .ZN(new_n2360_));
  OAI21_X1   g1975(.A1(new_n2360_), .A2(new_n398_), .B(new_n766_), .ZN(new_n2361_));
  AOI21_X1   g1976(.A1(new_n2361_), .A2(new_n772_), .B(new_n777_), .ZN(new_n2362_));
  OAI21_X1   g1977(.A1(new_n2362_), .A2(new_n394_), .B(new_n782_), .ZN(new_n2363_));
  AOI21_X1   g1978(.A1(new_n2363_), .A2(new_n390_), .B(new_n788_), .ZN(new_n2364_));
  OAI21_X1   g1979(.A1(new_n2364_), .A2(new_n793_), .B(new_n797_), .ZN(new_n2365_));
  AOI21_X1   g1980(.A1(new_n2365_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n2366_));
  OAI21_X1   g1981(.A1(new_n2366_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n2367_));
  AOI21_X1   g1982(.A1(new_n2367_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n2368_));
  OAI21_X1   g1983(.A1(new_n2368_), .A2(new_n912_), .B(new_n917_), .ZN(new_n2369_));
  AOI21_X1   g1984(.A1(new_n2369_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n2370_));
  OAI21_X1   g1985(.A1(new_n2370_), .A2(new_n893_), .B(new_n928_), .ZN(new_n2371_));
  OAI21_X1   g1986(.A1(new_n934_), .A2(\priority[18] ), .B(\req[18] ), .ZN(new_n2372_));
  AOI21_X1   g1987(.A1(new_n2371_), .A2(new_n1650_), .B(new_n2372_), .ZN(\grant[18] ));
  NOR2_X1    g1988(.A1(new_n1271_), .A2(new_n941_), .ZN(new_n2374_));
  OAI21_X1   g1989(.A1(new_n886_), .A2(new_n2374_), .B(new_n948_), .ZN(new_n2375_));
  AOI21_X1   g1990(.A1(new_n2375_), .A2(new_n953_), .B(new_n958_), .ZN(new_n2376_));
  OAI21_X1   g1991(.A1(new_n2376_), .A2(new_n883_), .B(new_n963_), .ZN(new_n2377_));
  AOI21_X1   g1992(.A1(new_n2377_), .A2(new_n880_), .B(new_n969_), .ZN(new_n2378_));
  OAI21_X1   g1993(.A1(new_n2378_), .A2(new_n973_), .B(new_n977_), .ZN(new_n2379_));
  AOI21_X1   g1994(.A1(new_n2379_), .A2(new_n876_), .B(new_n983_), .ZN(new_n2380_));
  OAI21_X1   g1995(.A1(new_n2380_), .A2(new_n872_), .B(new_n988_), .ZN(new_n2381_));
  AOI21_X1   g1996(.A1(new_n2381_), .A2(new_n993_), .B(new_n998_), .ZN(new_n2382_));
  OAI21_X1   g1997(.A1(new_n2382_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n2383_));
  AOI21_X1   g1998(.A1(new_n2383_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n2384_));
  OAI21_X1   g1999(.A1(new_n2384_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n2385_));
  AOI21_X1   g2000(.A1(new_n2385_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n2386_));
  OAI21_X1   g2001(.A1(new_n2386_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n2387_));
  AOI21_X1   g2002(.A1(new_n2387_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n2388_));
  OAI21_X1   g2003(.A1(new_n2388_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n2389_));
  AOI21_X1   g2004(.A1(new_n2389_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n2390_));
  OAI21_X1   g2005(.A1(new_n2390_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n2391_));
  AOI21_X1   g2006(.A1(new_n2391_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n2392_));
  OAI21_X1   g2007(.A1(new_n2392_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n2393_));
  AOI21_X1   g2008(.A1(new_n2393_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n2394_));
  OAI21_X1   g2009(.A1(new_n2394_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n2395_));
  AOI21_X1   g2010(.A1(new_n2395_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n2396_));
  OAI21_X1   g2011(.A1(new_n2396_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n2397_));
  AOI21_X1   g2012(.A1(new_n2397_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n2398_));
  OAI21_X1   g2013(.A1(new_n2398_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n2399_));
  AOI21_X1   g2014(.A1(new_n2399_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n2400_));
  OAI21_X1   g2015(.A1(new_n2400_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n2401_));
  AOI21_X1   g2016(.A1(new_n2401_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n2402_));
  OAI21_X1   g2017(.A1(new_n2402_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n2403_));
  AOI21_X1   g2018(.A1(new_n2403_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n2404_));
  OAI21_X1   g2019(.A1(new_n2404_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n2405_));
  AOI21_X1   g2020(.A1(new_n2405_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n2406_));
  OAI21_X1   g2021(.A1(new_n2406_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n2407_));
  AOI21_X1   g2022(.A1(new_n2407_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n2408_));
  OAI21_X1   g2023(.A1(new_n2408_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n2409_));
  AOI21_X1   g2024(.A1(new_n2409_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n2410_));
  OAI21_X1   g2025(.A1(new_n2410_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n2411_));
  AOI21_X1   g2026(.A1(new_n2411_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n2412_));
  OAI21_X1   g2027(.A1(new_n2412_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n2413_));
  AOI21_X1   g2028(.A1(new_n2413_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n2414_));
  OAI21_X1   g2029(.A1(new_n2414_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n2415_));
  OAI21_X1   g2030(.A1(new_n490_), .A2(\priority[19] ), .B(\req[19] ), .ZN(new_n2416_));
  AOI21_X1   g2031(.A1(new_n2415_), .A2(new_n1738_), .B(new_n2416_), .ZN(\grant[19] ));
  NOR2_X1    g2032(.A1(new_n487_), .A2(new_n1316_), .ZN(new_n2418_));
  OAI21_X1   g2033(.A1(new_n1269_), .A2(new_n2418_), .B(new_n1322_), .ZN(new_n2419_));
  AOI21_X1   g2034(.A1(new_n2419_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n2420_));
  OAI21_X1   g2035(.A1(new_n2420_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n2421_));
  AOI21_X1   g2036(.A1(new_n2421_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n2422_));
  OAI21_X1   g2037(.A1(new_n2422_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n2423_));
  AOI21_X1   g2038(.A1(new_n2423_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n2424_));
  OAI21_X1   g2039(.A1(new_n2424_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n2425_));
  AOI21_X1   g2040(.A1(new_n2425_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n2426_));
  OAI21_X1   g2041(.A1(new_n2426_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n2427_));
  AOI21_X1   g2042(.A1(new_n2427_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n2428_));
  OAI21_X1   g2043(.A1(new_n2428_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n2429_));
  AOI21_X1   g2044(.A1(new_n2429_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n2430_));
  OAI21_X1   g2045(.A1(new_n2430_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n2431_));
  AOI21_X1   g2046(.A1(new_n2431_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n2432_));
  OAI21_X1   g2047(.A1(new_n2432_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n2433_));
  AOI21_X1   g2048(.A1(new_n2433_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n2434_));
  OAI21_X1   g2049(.A1(new_n2434_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n2435_));
  AOI21_X1   g2050(.A1(new_n2435_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n2436_));
  OAI21_X1   g2051(.A1(new_n2436_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n2437_));
  AOI21_X1   g2052(.A1(new_n2437_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n2438_));
  OAI21_X1   g2053(.A1(new_n2438_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n2439_));
  AOI21_X1   g2054(.A1(new_n2439_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n2440_));
  OAI21_X1   g2055(.A1(new_n2440_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n2441_));
  AOI21_X1   g2056(.A1(new_n2441_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n2442_));
  OAI21_X1   g2057(.A1(new_n2442_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n2443_));
  AOI21_X1   g2058(.A1(new_n2443_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n2444_));
  OAI21_X1   g2059(.A1(new_n2444_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n2445_));
  AOI21_X1   g2060(.A1(new_n2445_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n2446_));
  OAI21_X1   g2061(.A1(new_n2446_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n2447_));
  AOI21_X1   g2062(.A1(new_n2447_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n2448_));
  OAI21_X1   g2063(.A1(new_n2448_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n2449_));
  AOI21_X1   g2064(.A1(new_n2449_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n2450_));
  OAI21_X1   g2065(.A1(new_n2450_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n2451_));
  AOI21_X1   g2066(.A1(new_n2451_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n2452_));
  OAI21_X1   g2067(.A1(new_n2452_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n2453_));
  AOI21_X1   g2068(.A1(new_n2453_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n2454_));
  OAI21_X1   g2069(.A1(new_n2454_), .A2(new_n506_), .B(new_n514_), .ZN(new_n2455_));
  AOI21_X1   g2070(.A1(new_n2455_), .A2(new_n520_), .B(new_n525_), .ZN(new_n2456_));
  OAI21_X1   g2071(.A1(new_n2456_), .A2(new_n502_), .B(new_n530_), .ZN(new_n2457_));
  AOI21_X1   g2072(.A1(new_n2457_), .A2(new_n498_), .B(new_n536_), .ZN(new_n2458_));
  OAI21_X1   g2073(.A1(new_n2458_), .A2(new_n541_), .B(new_n545_), .ZN(new_n2459_));
  OAI21_X1   g2074(.A1(new_n547_), .A2(\priority[20] ), .B(\req[20] ), .ZN(new_n2460_));
  AOI21_X1   g2075(.A1(new_n2459_), .A2(new_n493_), .B(new_n2460_), .ZN(\grant[20] ));
  NOR2_X1    g2076(.A1(new_n885_), .A2(new_n555_), .ZN(new_n2462_));
  OAI21_X1   g2077(.A1(new_n561_), .A2(new_n2462_), .B(new_n566_), .ZN(new_n2463_));
  AOI21_X1   g2078(.A1(new_n2463_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n2464_));
  OAI21_X1   g2079(.A1(new_n2464_), .A2(new_n479_), .B(new_n577_), .ZN(new_n2465_));
  AOI21_X1   g2080(.A1(new_n2465_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n2466_));
  OAI21_X1   g2081(.A1(new_n2466_), .A2(new_n474_), .B(new_n592_), .ZN(new_n2467_));
  AOI21_X1   g2082(.A1(new_n2467_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n2468_));
  OAI21_X1   g2083(.A1(new_n2468_), .A2(new_n603_), .B(new_n608_), .ZN(new_n2469_));
  AOI21_X1   g2084(.A1(new_n2469_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n2470_));
  OAI21_X1   g2085(.A1(new_n2470_), .A2(new_n461_), .B(new_n619_), .ZN(new_n2471_));
  AOI21_X1   g2086(.A1(new_n2471_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n2472_));
  OAI21_X1   g2087(.A1(new_n2472_), .A2(new_n456_), .B(new_n634_), .ZN(new_n2473_));
  AOI21_X1   g2088(.A1(new_n2473_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n2474_));
  OAI21_X1   g2089(.A1(new_n2474_), .A2(new_n645_), .B(new_n650_), .ZN(new_n2475_));
  AOI21_X1   g2090(.A1(new_n2475_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n2476_));
  OAI21_X1   g2091(.A1(new_n2476_), .A2(new_n443_), .B(new_n661_), .ZN(new_n2477_));
  AOI21_X1   g2092(.A1(new_n2477_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n2478_));
  OAI21_X1   g2093(.A1(new_n2478_), .A2(new_n438_), .B(new_n676_), .ZN(new_n2479_));
  AOI21_X1   g2094(.A1(new_n2479_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n2480_));
  OAI21_X1   g2095(.A1(new_n2480_), .A2(new_n687_), .B(new_n692_), .ZN(new_n2481_));
  AOI21_X1   g2096(.A1(new_n2481_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n2482_));
  OAI21_X1   g2097(.A1(new_n2482_), .A2(new_n425_), .B(new_n703_), .ZN(new_n2483_));
  AOI21_X1   g2098(.A1(new_n2483_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n2484_));
  OAI21_X1   g2099(.A1(new_n2484_), .A2(new_n420_), .B(new_n718_), .ZN(new_n2485_));
  AOI21_X1   g2100(.A1(new_n2485_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n2486_));
  OAI21_X1   g2101(.A1(new_n2486_), .A2(new_n729_), .B(new_n734_), .ZN(new_n2487_));
  AOI21_X1   g2102(.A1(new_n2487_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n2488_));
  OAI21_X1   g2103(.A1(new_n2488_), .A2(new_n407_), .B(new_n745_), .ZN(new_n2489_));
  AOI21_X1   g2104(.A1(new_n2489_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n2490_));
  OAI21_X1   g2105(.A1(new_n2490_), .A2(new_n402_), .B(new_n760_), .ZN(new_n2491_));
  AOI21_X1   g2106(.A1(new_n2491_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n2492_));
  OAI21_X1   g2107(.A1(new_n2492_), .A2(new_n771_), .B(new_n776_), .ZN(new_n2493_));
  AOI21_X1   g2108(.A1(new_n2493_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n2494_));
  OAI21_X1   g2109(.A1(new_n2494_), .A2(new_n389_), .B(new_n787_), .ZN(new_n2495_));
  AOI21_X1   g2110(.A1(new_n2495_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n2496_));
  OAI21_X1   g2111(.A1(new_n2496_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n2497_));
  AOI21_X1   g2112(.A1(new_n2497_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n2498_));
  OAI21_X1   g2113(.A1(new_n2498_), .A2(new_n900_), .B(new_n908_), .ZN(new_n2499_));
  AOI21_X1   g2114(.A1(new_n2499_), .A2(new_n913_), .B(new_n918_), .ZN(new_n2500_));
  OAI21_X1   g2115(.A1(new_n2500_), .A2(new_n897_), .B(new_n923_), .ZN(new_n2501_));
  AOI21_X1   g2116(.A1(new_n2501_), .A2(new_n894_), .B(new_n929_), .ZN(new_n2502_));
  OAI21_X1   g2117(.A1(new_n2502_), .A2(new_n933_), .B(new_n937_), .ZN(new_n2503_));
  OAI21_X1   g2118(.A1(new_n939_), .A2(\priority[21] ), .B(\req[21] ), .ZN(new_n2504_));
  AOI21_X1   g2119(.A1(new_n2503_), .A2(new_n890_), .B(new_n2504_), .ZN(\grant[21] ));
  NOR2_X1    g2120(.A1(new_n1268_), .A2(new_n947_), .ZN(new_n2506_));
  OAI21_X1   g2121(.A1(new_n952_), .A2(new_n2506_), .B(new_n957_), .ZN(new_n2507_));
  AOI21_X1   g2122(.A1(new_n2507_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n2508_));
  OAI21_X1   g2123(.A1(new_n2508_), .A2(new_n879_), .B(new_n968_), .ZN(new_n2509_));
  AOI21_X1   g2124(.A1(new_n2509_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n2510_));
  OAI21_X1   g2125(.A1(new_n2510_), .A2(new_n875_), .B(new_n982_), .ZN(new_n2511_));
  AOI21_X1   g2126(.A1(new_n2511_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n2512_));
  OAI21_X1   g2127(.A1(new_n2512_), .A2(new_n992_), .B(new_n997_), .ZN(new_n2513_));
  AOI21_X1   g2128(.A1(new_n2513_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n2514_));
  OAI21_X1   g2129(.A1(new_n2514_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n2515_));
  AOI21_X1   g2130(.A1(new_n2515_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n2516_));
  OAI21_X1   g2131(.A1(new_n2516_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n2517_));
  AOI21_X1   g2132(.A1(new_n2517_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n2518_));
  OAI21_X1   g2133(.A1(new_n2518_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n2519_));
  AOI21_X1   g2134(.A1(new_n2519_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n2520_));
  OAI21_X1   g2135(.A1(new_n2520_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n2521_));
  AOI21_X1   g2136(.A1(new_n2521_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n2522_));
  OAI21_X1   g2137(.A1(new_n2522_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n2523_));
  AOI21_X1   g2138(.A1(new_n2523_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n2524_));
  OAI21_X1   g2139(.A1(new_n2524_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n2525_));
  AOI21_X1   g2140(.A1(new_n2525_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n2526_));
  OAI21_X1   g2141(.A1(new_n2526_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n2527_));
  AOI21_X1   g2142(.A1(new_n2527_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n2528_));
  OAI21_X1   g2143(.A1(new_n2528_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n2529_));
  AOI21_X1   g2144(.A1(new_n2529_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n2530_));
  OAI21_X1   g2145(.A1(new_n2530_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n2531_));
  AOI21_X1   g2146(.A1(new_n2531_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n2532_));
  OAI21_X1   g2147(.A1(new_n2532_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n2533_));
  AOI21_X1   g2148(.A1(new_n2533_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n2534_));
  OAI21_X1   g2149(.A1(new_n2534_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n2535_));
  AOI21_X1   g2150(.A1(new_n2535_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n2536_));
  OAI21_X1   g2151(.A1(new_n2536_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n2537_));
  AOI21_X1   g2152(.A1(new_n2537_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n2538_));
  OAI21_X1   g2153(.A1(new_n2538_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n2539_));
  AOI21_X1   g2154(.A1(new_n2539_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n2540_));
  OAI21_X1   g2155(.A1(new_n2540_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n2541_));
  AOI21_X1   g2156(.A1(new_n2541_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n2542_));
  OAI21_X1   g2157(.A1(new_n2542_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n2543_));
  AOI21_X1   g2158(.A1(new_n2543_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n2544_));
  OAI21_X1   g2159(.A1(new_n2544_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n2545_));
  AOI21_X1   g2160(.A1(new_n2545_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n2546_));
  OAI21_X1   g2161(.A1(new_n2546_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n2547_));
  OAI21_X1   g2162(.A1(new_n486_), .A2(\priority[22] ), .B(\req[22] ), .ZN(new_n2548_));
  AOI21_X1   g2163(.A1(new_n2547_), .A2(new_n1273_), .B(new_n2548_), .ZN(\grant[22] ));
  NOR2_X1    g2164(.A1(new_n560_), .A2(new_n1321_), .ZN(new_n2550_));
  OAI21_X1   g2165(.A1(new_n1326_), .A2(new_n2550_), .B(new_n1330_), .ZN(new_n2551_));
  AOI21_X1   g2166(.A1(new_n2551_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n2552_));
  OAI21_X1   g2167(.A1(new_n2552_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n2553_));
  AOI21_X1   g2168(.A1(new_n2553_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n2554_));
  OAI21_X1   g2169(.A1(new_n2554_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n2555_));
  AOI21_X1   g2170(.A1(new_n2555_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n2556_));
  OAI21_X1   g2171(.A1(new_n2556_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n2557_));
  AOI21_X1   g2172(.A1(new_n2557_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n2558_));
  OAI21_X1   g2173(.A1(new_n2558_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n2559_));
  AOI21_X1   g2174(.A1(new_n2559_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n2560_));
  OAI21_X1   g2175(.A1(new_n2560_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n2561_));
  AOI21_X1   g2176(.A1(new_n2561_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n2562_));
  OAI21_X1   g2177(.A1(new_n2562_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n2563_));
  AOI21_X1   g2178(.A1(new_n2563_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n2564_));
  OAI21_X1   g2179(.A1(new_n2564_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n2565_));
  AOI21_X1   g2180(.A1(new_n2565_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n2566_));
  OAI21_X1   g2181(.A1(new_n2566_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n2567_));
  AOI21_X1   g2182(.A1(new_n2567_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n2568_));
  OAI21_X1   g2183(.A1(new_n2568_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n2569_));
  AOI21_X1   g2184(.A1(new_n2569_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n2570_));
  OAI21_X1   g2185(.A1(new_n2570_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n2571_));
  AOI21_X1   g2186(.A1(new_n2571_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n2572_));
  OAI21_X1   g2187(.A1(new_n2572_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n2573_));
  AOI21_X1   g2188(.A1(new_n2573_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n2574_));
  OAI21_X1   g2189(.A1(new_n2574_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n2575_));
  AOI21_X1   g2190(.A1(new_n2575_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n2576_));
  OAI21_X1   g2191(.A1(new_n2576_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n2577_));
  AOI21_X1   g2192(.A1(new_n2577_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n2578_));
  OAI21_X1   g2193(.A1(new_n2578_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n2579_));
  AOI21_X1   g2194(.A1(new_n2579_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n2580_));
  OAI21_X1   g2195(.A1(new_n2580_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n2581_));
  AOI21_X1   g2196(.A1(new_n2581_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n2582_));
  OAI21_X1   g2197(.A1(new_n2582_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n2583_));
  AOI21_X1   g2198(.A1(new_n2583_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n2584_));
  OAI21_X1   g2199(.A1(new_n2584_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n2585_));
  AOI21_X1   g2200(.A1(new_n2585_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n2586_));
  OAI21_X1   g2201(.A1(new_n2586_), .A2(new_n519_), .B(new_n524_), .ZN(new_n2587_));
  AOI21_X1   g2202(.A1(new_n2587_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n2588_));
  OAI21_X1   g2203(.A1(new_n2588_), .A2(new_n497_), .B(new_n535_), .ZN(new_n2589_));
  AOI21_X1   g2204(.A1(new_n2589_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n2590_));
  OAI21_X1   g2205(.A1(new_n2590_), .A2(new_n492_), .B(new_n550_), .ZN(new_n2591_));
  OAI21_X1   g2206(.A1(new_n553_), .A2(\priority[23] ), .B(\req[23] ), .ZN(new_n2592_));
  AOI21_X1   g2207(.A1(new_n2591_), .A2(new_n1558_), .B(new_n2592_), .ZN(\grant[23] ));
  NOR2_X1    g2208(.A1(new_n951_), .A2(new_n565_), .ZN(new_n2594_));
  OAI21_X1   g2209(.A1(new_n484_), .A2(new_n2594_), .B(new_n572_), .ZN(new_n2595_));
  AOI21_X1   g2210(.A1(new_n2595_), .A2(new_n480_), .B(new_n578_), .ZN(new_n2596_));
  OAI21_X1   g2211(.A1(new_n2596_), .A2(new_n583_), .B(new_n587_), .ZN(new_n2597_));
  AOI21_X1   g2212(.A1(new_n2597_), .A2(new_n475_), .B(new_n593_), .ZN(new_n2598_));
  OAI21_X1   g2213(.A1(new_n2598_), .A2(new_n470_), .B(new_n598_), .ZN(new_n2599_));
  AOI21_X1   g2214(.A1(new_n2599_), .A2(new_n604_), .B(new_n609_), .ZN(new_n2600_));
  OAI21_X1   g2215(.A1(new_n2600_), .A2(new_n466_), .B(new_n614_), .ZN(new_n2601_));
  AOI21_X1   g2216(.A1(new_n2601_), .A2(new_n462_), .B(new_n620_), .ZN(new_n2602_));
  OAI21_X1   g2217(.A1(new_n2602_), .A2(new_n625_), .B(new_n629_), .ZN(new_n2603_));
  AOI21_X1   g2218(.A1(new_n2603_), .A2(new_n457_), .B(new_n635_), .ZN(new_n2604_));
  OAI21_X1   g2219(.A1(new_n2604_), .A2(new_n452_), .B(new_n640_), .ZN(new_n2605_));
  AOI21_X1   g2220(.A1(new_n2605_), .A2(new_n646_), .B(new_n651_), .ZN(new_n2606_));
  OAI21_X1   g2221(.A1(new_n2606_), .A2(new_n448_), .B(new_n656_), .ZN(new_n2607_));
  AOI21_X1   g2222(.A1(new_n2607_), .A2(new_n444_), .B(new_n662_), .ZN(new_n2608_));
  OAI21_X1   g2223(.A1(new_n2608_), .A2(new_n667_), .B(new_n671_), .ZN(new_n2609_));
  AOI21_X1   g2224(.A1(new_n2609_), .A2(new_n439_), .B(new_n677_), .ZN(new_n2610_));
  OAI21_X1   g2225(.A1(new_n2610_), .A2(new_n434_), .B(new_n682_), .ZN(new_n2611_));
  AOI21_X1   g2226(.A1(new_n2611_), .A2(new_n688_), .B(new_n693_), .ZN(new_n2612_));
  OAI21_X1   g2227(.A1(new_n2612_), .A2(new_n430_), .B(new_n698_), .ZN(new_n2613_));
  AOI21_X1   g2228(.A1(new_n2613_), .A2(new_n426_), .B(new_n704_), .ZN(new_n2614_));
  OAI21_X1   g2229(.A1(new_n2614_), .A2(new_n709_), .B(new_n713_), .ZN(new_n2615_));
  AOI21_X1   g2230(.A1(new_n2615_), .A2(new_n421_), .B(new_n719_), .ZN(new_n2616_));
  OAI21_X1   g2231(.A1(new_n2616_), .A2(new_n416_), .B(new_n724_), .ZN(new_n2617_));
  AOI21_X1   g2232(.A1(new_n2617_), .A2(new_n730_), .B(new_n735_), .ZN(new_n2618_));
  OAI21_X1   g2233(.A1(new_n2618_), .A2(new_n412_), .B(new_n740_), .ZN(new_n2619_));
  AOI21_X1   g2234(.A1(new_n2619_), .A2(new_n408_), .B(new_n746_), .ZN(new_n2620_));
  OAI21_X1   g2235(.A1(new_n2620_), .A2(new_n751_), .B(new_n755_), .ZN(new_n2621_));
  AOI21_X1   g2236(.A1(new_n2621_), .A2(new_n403_), .B(new_n761_), .ZN(new_n2622_));
  OAI21_X1   g2237(.A1(new_n2622_), .A2(new_n398_), .B(new_n766_), .ZN(new_n2623_));
  AOI21_X1   g2238(.A1(new_n2623_), .A2(new_n772_), .B(new_n777_), .ZN(new_n2624_));
  OAI21_X1   g2239(.A1(new_n2624_), .A2(new_n394_), .B(new_n782_), .ZN(new_n2625_));
  AOI21_X1   g2240(.A1(new_n2625_), .A2(new_n390_), .B(new_n788_), .ZN(new_n2626_));
  OAI21_X1   g2241(.A1(new_n2626_), .A2(new_n793_), .B(new_n797_), .ZN(new_n2627_));
  AOI21_X1   g2242(.A1(new_n2627_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n2628_));
  OAI21_X1   g2243(.A1(new_n2628_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n2629_));
  AOI21_X1   g2244(.A1(new_n2629_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n2630_));
  OAI21_X1   g2245(.A1(new_n2630_), .A2(new_n912_), .B(new_n917_), .ZN(new_n2631_));
  AOI21_X1   g2246(.A1(new_n2631_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n2632_));
  OAI21_X1   g2247(.A1(new_n2632_), .A2(new_n893_), .B(new_n928_), .ZN(new_n2633_));
  AOI21_X1   g2248(.A1(new_n2633_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n2634_));
  OAI21_X1   g2249(.A1(new_n2634_), .A2(new_n889_), .B(new_n942_), .ZN(new_n2635_));
  OAI21_X1   g2250(.A1(new_n945_), .A2(\priority[24] ), .B(\req[24] ), .ZN(new_n2636_));
  AOI21_X1   g2251(.A1(new_n2635_), .A2(new_n1648_), .B(new_n2636_), .ZN(\grant[24] ));
  NOR2_X1    g2252(.A1(new_n1325_), .A2(new_n956_), .ZN(new_n2638_));
  OAI21_X1   g2253(.A1(new_n883_), .A2(new_n2638_), .B(new_n963_), .ZN(new_n2639_));
  AOI21_X1   g2254(.A1(new_n2639_), .A2(new_n880_), .B(new_n969_), .ZN(new_n2640_));
  OAI21_X1   g2255(.A1(new_n2640_), .A2(new_n973_), .B(new_n977_), .ZN(new_n2641_));
  AOI21_X1   g2256(.A1(new_n2641_), .A2(new_n876_), .B(new_n983_), .ZN(new_n2642_));
  OAI21_X1   g2257(.A1(new_n2642_), .A2(new_n872_), .B(new_n988_), .ZN(new_n2643_));
  AOI21_X1   g2258(.A1(new_n2643_), .A2(new_n993_), .B(new_n998_), .ZN(new_n2644_));
  OAI21_X1   g2259(.A1(new_n2644_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n2645_));
  AOI21_X1   g2260(.A1(new_n2645_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n2646_));
  OAI21_X1   g2261(.A1(new_n2646_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n2647_));
  AOI21_X1   g2262(.A1(new_n2647_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n2648_));
  OAI21_X1   g2263(.A1(new_n2648_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n2649_));
  AOI21_X1   g2264(.A1(new_n2649_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n2650_));
  OAI21_X1   g2265(.A1(new_n2650_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n2651_));
  AOI21_X1   g2266(.A1(new_n2651_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n2652_));
  OAI21_X1   g2267(.A1(new_n2652_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n2653_));
  AOI21_X1   g2268(.A1(new_n2653_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n2654_));
  OAI21_X1   g2269(.A1(new_n2654_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n2655_));
  AOI21_X1   g2270(.A1(new_n2655_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n2656_));
  OAI21_X1   g2271(.A1(new_n2656_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n2657_));
  AOI21_X1   g2272(.A1(new_n2657_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n2658_));
  OAI21_X1   g2273(.A1(new_n2658_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n2659_));
  AOI21_X1   g2274(.A1(new_n2659_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n2660_));
  OAI21_X1   g2275(.A1(new_n2660_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n2661_));
  AOI21_X1   g2276(.A1(new_n2661_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n2662_));
  OAI21_X1   g2277(.A1(new_n2662_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n2663_));
  AOI21_X1   g2278(.A1(new_n2663_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n2664_));
  OAI21_X1   g2279(.A1(new_n2664_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n2665_));
  AOI21_X1   g2280(.A1(new_n2665_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n2666_));
  OAI21_X1   g2281(.A1(new_n2666_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n2667_));
  AOI21_X1   g2282(.A1(new_n2667_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n2668_));
  OAI21_X1   g2283(.A1(new_n2668_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n2669_));
  AOI21_X1   g2284(.A1(new_n2669_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n2670_));
  OAI21_X1   g2285(.A1(new_n2670_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n2671_));
  AOI21_X1   g2286(.A1(new_n2671_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n2672_));
  OAI21_X1   g2287(.A1(new_n2672_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n2673_));
  AOI21_X1   g2288(.A1(new_n2673_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n2674_));
  OAI21_X1   g2289(.A1(new_n2674_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n2675_));
  AOI21_X1   g2290(.A1(new_n2675_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n2676_));
  OAI21_X1   g2291(.A1(new_n2676_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n2677_));
  AOI21_X1   g2292(.A1(new_n2677_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n2678_));
  OAI21_X1   g2293(.A1(new_n2678_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n2679_));
  OAI21_X1   g2294(.A1(new_n559_), .A2(\priority[25] ), .B(\req[25] ), .ZN(new_n2680_));
  AOI21_X1   g2295(.A1(new_n2679_), .A2(new_n1736_), .B(new_n2680_), .ZN(\grant[25] ));
  NOR2_X1    g2296(.A1(new_n483_), .A2(new_n1329_), .ZN(new_n2682_));
  OAI21_X1   g2297(.A1(new_n1266_), .A2(new_n2682_), .B(new_n1335_), .ZN(new_n2683_));
  AOI21_X1   g2298(.A1(new_n2683_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n2684_));
  OAI21_X1   g2299(.A1(new_n2684_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n2685_));
  AOI21_X1   g2300(.A1(new_n2685_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n2686_));
  OAI21_X1   g2301(.A1(new_n2686_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n2687_));
  AOI21_X1   g2302(.A1(new_n2687_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n2688_));
  OAI21_X1   g2303(.A1(new_n2688_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n2689_));
  AOI21_X1   g2304(.A1(new_n2689_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n2690_));
  OAI21_X1   g2305(.A1(new_n2690_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n2691_));
  AOI21_X1   g2306(.A1(new_n2691_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n2692_));
  OAI21_X1   g2307(.A1(new_n2692_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n2693_));
  AOI21_X1   g2308(.A1(new_n2693_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n2694_));
  OAI21_X1   g2309(.A1(new_n2694_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n2695_));
  AOI21_X1   g2310(.A1(new_n2695_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n2696_));
  OAI21_X1   g2311(.A1(new_n2696_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n2697_));
  AOI21_X1   g2312(.A1(new_n2697_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n2698_));
  OAI21_X1   g2313(.A1(new_n2698_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n2699_));
  AOI21_X1   g2314(.A1(new_n2699_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n2700_));
  OAI21_X1   g2315(.A1(new_n2700_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n2701_));
  AOI21_X1   g2316(.A1(new_n2701_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n2702_));
  OAI21_X1   g2317(.A1(new_n2702_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n2703_));
  AOI21_X1   g2318(.A1(new_n2703_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n2704_));
  OAI21_X1   g2319(.A1(new_n2704_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n2705_));
  AOI21_X1   g2320(.A1(new_n2705_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n2706_));
  OAI21_X1   g2321(.A1(new_n2706_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n2707_));
  AOI21_X1   g2322(.A1(new_n2707_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n2708_));
  OAI21_X1   g2323(.A1(new_n2708_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n2709_));
  AOI21_X1   g2324(.A1(new_n2709_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n2710_));
  OAI21_X1   g2325(.A1(new_n2710_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n2711_));
  AOI21_X1   g2326(.A1(new_n2711_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n2712_));
  OAI21_X1   g2327(.A1(new_n2712_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n2713_));
  AOI21_X1   g2328(.A1(new_n2713_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n2714_));
  OAI21_X1   g2329(.A1(new_n2714_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n2715_));
  AOI21_X1   g2330(.A1(new_n2715_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n2716_));
  OAI21_X1   g2331(.A1(new_n2716_), .A2(new_n506_), .B(new_n514_), .ZN(new_n2717_));
  AOI21_X1   g2332(.A1(new_n2717_), .A2(new_n520_), .B(new_n525_), .ZN(new_n2718_));
  OAI21_X1   g2333(.A1(new_n2718_), .A2(new_n502_), .B(new_n530_), .ZN(new_n2719_));
  AOI21_X1   g2334(.A1(new_n2719_), .A2(new_n498_), .B(new_n536_), .ZN(new_n2720_));
  OAI21_X1   g2335(.A1(new_n2720_), .A2(new_n541_), .B(new_n545_), .ZN(new_n2721_));
  AOI21_X1   g2336(.A1(new_n2721_), .A2(new_n493_), .B(new_n551_), .ZN(new_n2722_));
  OAI21_X1   g2337(.A1(new_n2722_), .A2(new_n488_), .B(new_n556_), .ZN(new_n2723_));
  OAI21_X1   g2338(.A1(new_n563_), .A2(\priority[26] ), .B(\req[26] ), .ZN(new_n2724_));
  AOI21_X1   g2339(.A1(new_n2723_), .A2(new_n562_), .B(new_n2724_), .ZN(\grant[26] ));
  NOR2_X1    g2340(.A1(new_n882_), .A2(new_n571_), .ZN(new_n2726_));
  OAI21_X1   g2341(.A1(new_n479_), .A2(new_n2726_), .B(new_n577_), .ZN(new_n2727_));
  AOI21_X1   g2342(.A1(new_n2727_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n2728_));
  OAI21_X1   g2343(.A1(new_n2728_), .A2(new_n474_), .B(new_n592_), .ZN(new_n2729_));
  AOI21_X1   g2344(.A1(new_n2729_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n2730_));
  OAI21_X1   g2345(.A1(new_n2730_), .A2(new_n603_), .B(new_n608_), .ZN(new_n2731_));
  AOI21_X1   g2346(.A1(new_n2731_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n2732_));
  OAI21_X1   g2347(.A1(new_n2732_), .A2(new_n461_), .B(new_n619_), .ZN(new_n2733_));
  AOI21_X1   g2348(.A1(new_n2733_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n2734_));
  OAI21_X1   g2349(.A1(new_n2734_), .A2(new_n456_), .B(new_n634_), .ZN(new_n2735_));
  AOI21_X1   g2350(.A1(new_n2735_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n2736_));
  OAI21_X1   g2351(.A1(new_n2736_), .A2(new_n645_), .B(new_n650_), .ZN(new_n2737_));
  AOI21_X1   g2352(.A1(new_n2737_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n2738_));
  OAI21_X1   g2353(.A1(new_n2738_), .A2(new_n443_), .B(new_n661_), .ZN(new_n2739_));
  AOI21_X1   g2354(.A1(new_n2739_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n2740_));
  OAI21_X1   g2355(.A1(new_n2740_), .A2(new_n438_), .B(new_n676_), .ZN(new_n2741_));
  AOI21_X1   g2356(.A1(new_n2741_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n2742_));
  OAI21_X1   g2357(.A1(new_n2742_), .A2(new_n687_), .B(new_n692_), .ZN(new_n2743_));
  AOI21_X1   g2358(.A1(new_n2743_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n2744_));
  OAI21_X1   g2359(.A1(new_n2744_), .A2(new_n425_), .B(new_n703_), .ZN(new_n2745_));
  AOI21_X1   g2360(.A1(new_n2745_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n2746_));
  OAI21_X1   g2361(.A1(new_n2746_), .A2(new_n420_), .B(new_n718_), .ZN(new_n2747_));
  AOI21_X1   g2362(.A1(new_n2747_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n2748_));
  OAI21_X1   g2363(.A1(new_n2748_), .A2(new_n729_), .B(new_n734_), .ZN(new_n2749_));
  AOI21_X1   g2364(.A1(new_n2749_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n2750_));
  OAI21_X1   g2365(.A1(new_n2750_), .A2(new_n407_), .B(new_n745_), .ZN(new_n2751_));
  AOI21_X1   g2366(.A1(new_n2751_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n2752_));
  OAI21_X1   g2367(.A1(new_n2752_), .A2(new_n402_), .B(new_n760_), .ZN(new_n2753_));
  AOI21_X1   g2368(.A1(new_n2753_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n2754_));
  OAI21_X1   g2369(.A1(new_n2754_), .A2(new_n771_), .B(new_n776_), .ZN(new_n2755_));
  AOI21_X1   g2370(.A1(new_n2755_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n2756_));
  OAI21_X1   g2371(.A1(new_n2756_), .A2(new_n389_), .B(new_n787_), .ZN(new_n2757_));
  AOI21_X1   g2372(.A1(new_n2757_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n2758_));
  OAI21_X1   g2373(.A1(new_n2758_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n2759_));
  AOI21_X1   g2374(.A1(new_n2759_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n2760_));
  OAI21_X1   g2375(.A1(new_n2760_), .A2(new_n900_), .B(new_n908_), .ZN(new_n2761_));
  AOI21_X1   g2376(.A1(new_n2761_), .A2(new_n913_), .B(new_n918_), .ZN(new_n2762_));
  OAI21_X1   g2377(.A1(new_n2762_), .A2(new_n897_), .B(new_n923_), .ZN(new_n2763_));
  AOI21_X1   g2378(.A1(new_n2763_), .A2(new_n894_), .B(new_n929_), .ZN(new_n2764_));
  OAI21_X1   g2379(.A1(new_n2764_), .A2(new_n933_), .B(new_n937_), .ZN(new_n2765_));
  AOI21_X1   g2380(.A1(new_n2765_), .A2(new_n890_), .B(new_n943_), .ZN(new_n2766_));
  OAI21_X1   g2381(.A1(new_n2766_), .A2(new_n886_), .B(new_n948_), .ZN(new_n2767_));
  OAI21_X1   g2382(.A1(new_n954_), .A2(\priority[27] ), .B(\req[27] ), .ZN(new_n2768_));
  AOI21_X1   g2383(.A1(new_n2767_), .A2(new_n953_), .B(new_n2768_), .ZN(\grant[27] ));
  NOR2_X1    g2384(.A1(new_n1265_), .A2(new_n962_), .ZN(new_n2770_));
  OAI21_X1   g2385(.A1(new_n879_), .A2(new_n2770_), .B(new_n968_), .ZN(new_n2771_));
  AOI21_X1   g2386(.A1(new_n2771_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n2772_));
  OAI21_X1   g2387(.A1(new_n2772_), .A2(new_n875_), .B(new_n982_), .ZN(new_n2773_));
  AOI21_X1   g2388(.A1(new_n2773_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n2774_));
  OAI21_X1   g2389(.A1(new_n2774_), .A2(new_n992_), .B(new_n997_), .ZN(new_n2775_));
  AOI21_X1   g2390(.A1(new_n2775_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n2776_));
  OAI21_X1   g2391(.A1(new_n2776_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n2777_));
  AOI21_X1   g2392(.A1(new_n2777_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n2778_));
  OAI21_X1   g2393(.A1(new_n2778_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n2779_));
  AOI21_X1   g2394(.A1(new_n2779_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n2780_));
  OAI21_X1   g2395(.A1(new_n2780_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n2781_));
  AOI21_X1   g2396(.A1(new_n2781_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n2782_));
  OAI21_X1   g2397(.A1(new_n2782_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n2783_));
  AOI21_X1   g2398(.A1(new_n2783_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n2784_));
  OAI21_X1   g2399(.A1(new_n2784_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n2785_));
  AOI21_X1   g2400(.A1(new_n2785_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n2786_));
  OAI21_X1   g2401(.A1(new_n2786_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n2787_));
  AOI21_X1   g2402(.A1(new_n2787_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n2788_));
  OAI21_X1   g2403(.A1(new_n2788_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n2789_));
  AOI21_X1   g2404(.A1(new_n2789_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n2790_));
  OAI21_X1   g2405(.A1(new_n2790_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n2791_));
  AOI21_X1   g2406(.A1(new_n2791_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n2792_));
  OAI21_X1   g2407(.A1(new_n2792_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n2793_));
  AOI21_X1   g2408(.A1(new_n2793_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n2794_));
  OAI21_X1   g2409(.A1(new_n2794_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n2795_));
  AOI21_X1   g2410(.A1(new_n2795_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n2796_));
  OAI21_X1   g2411(.A1(new_n2796_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n2797_));
  AOI21_X1   g2412(.A1(new_n2797_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n2798_));
  OAI21_X1   g2413(.A1(new_n2798_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n2799_));
  AOI21_X1   g2414(.A1(new_n2799_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n2800_));
  OAI21_X1   g2415(.A1(new_n2800_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n2801_));
  AOI21_X1   g2416(.A1(new_n2801_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n2802_));
  OAI21_X1   g2417(.A1(new_n2802_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n2803_));
  AOI21_X1   g2418(.A1(new_n2803_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n2804_));
  OAI21_X1   g2419(.A1(new_n2804_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n2805_));
  AOI21_X1   g2420(.A1(new_n2805_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n2806_));
  OAI21_X1   g2421(.A1(new_n2806_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n2807_));
  AOI21_X1   g2422(.A1(new_n2807_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n2808_));
  OAI21_X1   g2423(.A1(new_n2808_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n2809_));
  AOI21_X1   g2424(.A1(new_n2809_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n2810_));
  OAI21_X1   g2425(.A1(new_n2810_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n2811_));
  OAI21_X1   g2426(.A1(new_n482_), .A2(\priority[28] ), .B(\req[28] ), .ZN(new_n2812_));
  AOI21_X1   g2427(.A1(new_n2811_), .A2(new_n1327_), .B(new_n2812_), .ZN(\grant[28] ));
  NOR2_X1    g2428(.A1(new_n478_), .A2(new_n1334_), .ZN(new_n2814_));
  OAI21_X1   g2429(.A1(new_n1262_), .A2(new_n2814_), .B(new_n1339_), .ZN(new_n2815_));
  AOI21_X1   g2430(.A1(new_n2815_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n2816_));
  OAI21_X1   g2431(.A1(new_n2816_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n2817_));
  AOI21_X1   g2432(.A1(new_n2817_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n2818_));
  OAI21_X1   g2433(.A1(new_n2818_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n2819_));
  AOI21_X1   g2434(.A1(new_n2819_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n2820_));
  OAI21_X1   g2435(.A1(new_n2820_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n2821_));
  AOI21_X1   g2436(.A1(new_n2821_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n2822_));
  OAI21_X1   g2437(.A1(new_n2822_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n2823_));
  AOI21_X1   g2438(.A1(new_n2823_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n2824_));
  OAI21_X1   g2439(.A1(new_n2824_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n2825_));
  AOI21_X1   g2440(.A1(new_n2825_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n2826_));
  OAI21_X1   g2441(.A1(new_n2826_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n2827_));
  AOI21_X1   g2442(.A1(new_n2827_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n2828_));
  OAI21_X1   g2443(.A1(new_n2828_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n2829_));
  AOI21_X1   g2444(.A1(new_n2829_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n2830_));
  OAI21_X1   g2445(.A1(new_n2830_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n2831_));
  AOI21_X1   g2446(.A1(new_n2831_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n2832_));
  OAI21_X1   g2447(.A1(new_n2832_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n2833_));
  AOI21_X1   g2448(.A1(new_n2833_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n2834_));
  OAI21_X1   g2449(.A1(new_n2834_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n2835_));
  AOI21_X1   g2450(.A1(new_n2835_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n2836_));
  OAI21_X1   g2451(.A1(new_n2836_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n2837_));
  AOI21_X1   g2452(.A1(new_n2837_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n2838_));
  OAI21_X1   g2453(.A1(new_n2838_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n2839_));
  AOI21_X1   g2454(.A1(new_n2839_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n2840_));
  OAI21_X1   g2455(.A1(new_n2840_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n2841_));
  AOI21_X1   g2456(.A1(new_n2841_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n2842_));
  OAI21_X1   g2457(.A1(new_n2842_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n2843_));
  AOI21_X1   g2458(.A1(new_n2843_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n2844_));
  OAI21_X1   g2459(.A1(new_n2844_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n2845_));
  AOI21_X1   g2460(.A1(new_n2845_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n2846_));
  OAI21_X1   g2461(.A1(new_n2846_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n2847_));
  AOI21_X1   g2462(.A1(new_n2847_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n2848_));
  OAI21_X1   g2463(.A1(new_n2848_), .A2(new_n519_), .B(new_n524_), .ZN(new_n2849_));
  AOI21_X1   g2464(.A1(new_n2849_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n2850_));
  OAI21_X1   g2465(.A1(new_n2850_), .A2(new_n497_), .B(new_n535_), .ZN(new_n2851_));
  AOI21_X1   g2466(.A1(new_n2851_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n2852_));
  OAI21_X1   g2467(.A1(new_n2852_), .A2(new_n492_), .B(new_n550_), .ZN(new_n2853_));
  AOI21_X1   g2468(.A1(new_n2853_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n2854_));
  OAI21_X1   g2469(.A1(new_n2854_), .A2(new_n561_), .B(new_n566_), .ZN(new_n2855_));
  OAI21_X1   g2470(.A1(new_n569_), .A2(\priority[29] ), .B(\req[29] ), .ZN(new_n2856_));
  AOI21_X1   g2471(.A1(new_n2855_), .A2(new_n1556_), .B(new_n2856_), .ZN(\grant[29] ));
  NOR2_X1    g2472(.A1(new_n878_), .A2(new_n576_), .ZN(new_n2858_));
  OAI21_X1   g2473(.A1(new_n583_), .A2(new_n2858_), .B(new_n587_), .ZN(new_n2859_));
  AOI21_X1   g2474(.A1(new_n2859_), .A2(new_n475_), .B(new_n593_), .ZN(new_n2860_));
  OAI21_X1   g2475(.A1(new_n2860_), .A2(new_n470_), .B(new_n598_), .ZN(new_n2861_));
  AOI21_X1   g2476(.A1(new_n2861_), .A2(new_n604_), .B(new_n609_), .ZN(new_n2862_));
  OAI21_X1   g2477(.A1(new_n2862_), .A2(new_n466_), .B(new_n614_), .ZN(new_n2863_));
  AOI21_X1   g2478(.A1(new_n2863_), .A2(new_n462_), .B(new_n620_), .ZN(new_n2864_));
  OAI21_X1   g2479(.A1(new_n2864_), .A2(new_n625_), .B(new_n629_), .ZN(new_n2865_));
  AOI21_X1   g2480(.A1(new_n2865_), .A2(new_n457_), .B(new_n635_), .ZN(new_n2866_));
  OAI21_X1   g2481(.A1(new_n2866_), .A2(new_n452_), .B(new_n640_), .ZN(new_n2867_));
  AOI21_X1   g2482(.A1(new_n2867_), .A2(new_n646_), .B(new_n651_), .ZN(new_n2868_));
  OAI21_X1   g2483(.A1(new_n2868_), .A2(new_n448_), .B(new_n656_), .ZN(new_n2869_));
  AOI21_X1   g2484(.A1(new_n2869_), .A2(new_n444_), .B(new_n662_), .ZN(new_n2870_));
  OAI21_X1   g2485(.A1(new_n2870_), .A2(new_n667_), .B(new_n671_), .ZN(new_n2871_));
  AOI21_X1   g2486(.A1(new_n2871_), .A2(new_n439_), .B(new_n677_), .ZN(new_n2872_));
  OAI21_X1   g2487(.A1(new_n2872_), .A2(new_n434_), .B(new_n682_), .ZN(new_n2873_));
  AOI21_X1   g2488(.A1(new_n2873_), .A2(new_n688_), .B(new_n693_), .ZN(new_n2874_));
  OAI21_X1   g2489(.A1(new_n2874_), .A2(new_n430_), .B(new_n698_), .ZN(new_n2875_));
  AOI21_X1   g2490(.A1(new_n2875_), .A2(new_n426_), .B(new_n704_), .ZN(new_n2876_));
  OAI21_X1   g2491(.A1(new_n2876_), .A2(new_n709_), .B(new_n713_), .ZN(new_n2877_));
  AOI21_X1   g2492(.A1(new_n2877_), .A2(new_n421_), .B(new_n719_), .ZN(new_n2878_));
  OAI21_X1   g2493(.A1(new_n2878_), .A2(new_n416_), .B(new_n724_), .ZN(new_n2879_));
  AOI21_X1   g2494(.A1(new_n2879_), .A2(new_n730_), .B(new_n735_), .ZN(new_n2880_));
  OAI21_X1   g2495(.A1(new_n2880_), .A2(new_n412_), .B(new_n740_), .ZN(new_n2881_));
  AOI21_X1   g2496(.A1(new_n2881_), .A2(new_n408_), .B(new_n746_), .ZN(new_n2882_));
  OAI21_X1   g2497(.A1(new_n2882_), .A2(new_n751_), .B(new_n755_), .ZN(new_n2883_));
  AOI21_X1   g2498(.A1(new_n2883_), .A2(new_n403_), .B(new_n761_), .ZN(new_n2884_));
  OAI21_X1   g2499(.A1(new_n2884_), .A2(new_n398_), .B(new_n766_), .ZN(new_n2885_));
  AOI21_X1   g2500(.A1(new_n2885_), .A2(new_n772_), .B(new_n777_), .ZN(new_n2886_));
  OAI21_X1   g2501(.A1(new_n2886_), .A2(new_n394_), .B(new_n782_), .ZN(new_n2887_));
  AOI21_X1   g2502(.A1(new_n2887_), .A2(new_n390_), .B(new_n788_), .ZN(new_n2888_));
  OAI21_X1   g2503(.A1(new_n2888_), .A2(new_n793_), .B(new_n797_), .ZN(new_n2889_));
  AOI21_X1   g2504(.A1(new_n2889_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n2890_));
  OAI21_X1   g2505(.A1(new_n2890_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n2891_));
  AOI21_X1   g2506(.A1(new_n2891_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n2892_));
  OAI21_X1   g2507(.A1(new_n2892_), .A2(new_n912_), .B(new_n917_), .ZN(new_n2893_));
  AOI21_X1   g2508(.A1(new_n2893_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n2894_));
  OAI21_X1   g2509(.A1(new_n2894_), .A2(new_n893_), .B(new_n928_), .ZN(new_n2895_));
  AOI21_X1   g2510(.A1(new_n2895_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n2896_));
  OAI21_X1   g2511(.A1(new_n2896_), .A2(new_n889_), .B(new_n942_), .ZN(new_n2897_));
  AOI21_X1   g2512(.A1(new_n2897_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n2898_));
  OAI21_X1   g2513(.A1(new_n2898_), .A2(new_n952_), .B(new_n957_), .ZN(new_n2899_));
  OAI21_X1   g2514(.A1(new_n960_), .A2(\priority[30] ), .B(\req[30] ), .ZN(new_n2900_));
  AOI21_X1   g2515(.A1(new_n2899_), .A2(new_n1646_), .B(new_n2900_), .ZN(\grant[30] ));
  NOR2_X1    g2516(.A1(new_n1261_), .A2(new_n967_), .ZN(new_n2902_));
  OAI21_X1   g2517(.A1(new_n973_), .A2(new_n2902_), .B(new_n977_), .ZN(new_n2903_));
  AOI21_X1   g2518(.A1(new_n2903_), .A2(new_n876_), .B(new_n983_), .ZN(new_n2904_));
  OAI21_X1   g2519(.A1(new_n2904_), .A2(new_n872_), .B(new_n988_), .ZN(new_n2905_));
  AOI21_X1   g2520(.A1(new_n2905_), .A2(new_n993_), .B(new_n998_), .ZN(new_n2906_));
  OAI21_X1   g2521(.A1(new_n2906_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n2907_));
  AOI21_X1   g2522(.A1(new_n2907_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n2908_));
  OAI21_X1   g2523(.A1(new_n2908_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n2909_));
  AOI21_X1   g2524(.A1(new_n2909_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n2910_));
  OAI21_X1   g2525(.A1(new_n2910_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n2911_));
  AOI21_X1   g2526(.A1(new_n2911_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n2912_));
  OAI21_X1   g2527(.A1(new_n2912_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n2913_));
  AOI21_X1   g2528(.A1(new_n2913_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n2914_));
  OAI21_X1   g2529(.A1(new_n2914_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n2915_));
  AOI21_X1   g2530(.A1(new_n2915_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n2916_));
  OAI21_X1   g2531(.A1(new_n2916_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n2917_));
  AOI21_X1   g2532(.A1(new_n2917_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n2918_));
  OAI21_X1   g2533(.A1(new_n2918_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n2919_));
  AOI21_X1   g2534(.A1(new_n2919_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n2920_));
  OAI21_X1   g2535(.A1(new_n2920_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n2921_));
  AOI21_X1   g2536(.A1(new_n2921_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n2922_));
  OAI21_X1   g2537(.A1(new_n2922_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n2923_));
  AOI21_X1   g2538(.A1(new_n2923_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n2924_));
  OAI21_X1   g2539(.A1(new_n2924_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n2925_));
  AOI21_X1   g2540(.A1(new_n2925_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n2926_));
  OAI21_X1   g2541(.A1(new_n2926_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n2927_));
  AOI21_X1   g2542(.A1(new_n2927_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n2928_));
  OAI21_X1   g2543(.A1(new_n2928_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n2929_));
  AOI21_X1   g2544(.A1(new_n2929_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n2930_));
  OAI21_X1   g2545(.A1(new_n2930_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n2931_));
  AOI21_X1   g2546(.A1(new_n2931_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n2932_));
  OAI21_X1   g2547(.A1(new_n2932_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n2933_));
  AOI21_X1   g2548(.A1(new_n2933_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n2934_));
  OAI21_X1   g2549(.A1(new_n2934_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n2935_));
  AOI21_X1   g2550(.A1(new_n2935_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n2936_));
  OAI21_X1   g2551(.A1(new_n2936_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n2937_));
  AOI21_X1   g2552(.A1(new_n2937_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n2938_));
  OAI21_X1   g2553(.A1(new_n2938_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n2939_));
  AOI21_X1   g2554(.A1(new_n2939_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n2940_));
  OAI21_X1   g2555(.A1(new_n2940_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n2941_));
  AOI21_X1   g2556(.A1(new_n2941_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n2942_));
  OAI21_X1   g2557(.A1(new_n2942_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n2943_));
  OAI21_X1   g2558(.A1(new_n477_), .A2(\priority[31] ), .B(\req[31] ), .ZN(new_n2944_));
  AOI21_X1   g2559(.A1(new_n2943_), .A2(new_n1734_), .B(new_n2944_), .ZN(\grant[31] ));
  NOR2_X1    g2560(.A1(new_n582_), .A2(new_n1338_), .ZN(new_n2946_));
  OAI21_X1   g2561(.A1(new_n1344_), .A2(new_n2946_), .B(new_n1347_), .ZN(new_n2947_));
  AOI21_X1   g2562(.A1(new_n2947_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n2948_));
  OAI21_X1   g2563(.A1(new_n2948_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n2949_));
  AOI21_X1   g2564(.A1(new_n2949_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n2950_));
  OAI21_X1   g2565(.A1(new_n2950_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n2951_));
  AOI21_X1   g2566(.A1(new_n2951_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n2952_));
  OAI21_X1   g2567(.A1(new_n2952_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n2953_));
  AOI21_X1   g2568(.A1(new_n2953_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n2954_));
  OAI21_X1   g2569(.A1(new_n2954_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n2955_));
  AOI21_X1   g2570(.A1(new_n2955_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n2956_));
  OAI21_X1   g2571(.A1(new_n2956_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n2957_));
  AOI21_X1   g2572(.A1(new_n2957_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n2958_));
  OAI21_X1   g2573(.A1(new_n2958_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n2959_));
  AOI21_X1   g2574(.A1(new_n2959_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n2960_));
  OAI21_X1   g2575(.A1(new_n2960_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n2961_));
  AOI21_X1   g2576(.A1(new_n2961_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n2962_));
  OAI21_X1   g2577(.A1(new_n2962_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n2963_));
  AOI21_X1   g2578(.A1(new_n2963_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n2964_));
  OAI21_X1   g2579(.A1(new_n2964_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n2965_));
  AOI21_X1   g2580(.A1(new_n2965_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n2966_));
  OAI21_X1   g2581(.A1(new_n2966_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n2967_));
  AOI21_X1   g2582(.A1(new_n2967_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n2968_));
  OAI21_X1   g2583(.A1(new_n2968_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n2969_));
  AOI21_X1   g2584(.A1(new_n2969_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n2970_));
  OAI21_X1   g2585(.A1(new_n2970_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n2971_));
  AOI21_X1   g2586(.A1(new_n2971_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n2972_));
  OAI21_X1   g2587(.A1(new_n2972_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n2973_));
  AOI21_X1   g2588(.A1(new_n2973_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n2974_));
  OAI21_X1   g2589(.A1(new_n2974_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n2975_));
  AOI21_X1   g2590(.A1(new_n2975_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n2976_));
  OAI21_X1   g2591(.A1(new_n2976_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n2977_));
  AOI21_X1   g2592(.A1(new_n2977_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n2978_));
  OAI21_X1   g2593(.A1(new_n2978_), .A2(new_n506_), .B(new_n514_), .ZN(new_n2979_));
  AOI21_X1   g2594(.A1(new_n2979_), .A2(new_n520_), .B(new_n525_), .ZN(new_n2980_));
  OAI21_X1   g2595(.A1(new_n2980_), .A2(new_n502_), .B(new_n530_), .ZN(new_n2981_));
  AOI21_X1   g2596(.A1(new_n2981_), .A2(new_n498_), .B(new_n536_), .ZN(new_n2982_));
  OAI21_X1   g2597(.A1(new_n2982_), .A2(new_n541_), .B(new_n545_), .ZN(new_n2983_));
  AOI21_X1   g2598(.A1(new_n2983_), .A2(new_n493_), .B(new_n551_), .ZN(new_n2984_));
  OAI21_X1   g2599(.A1(new_n2984_), .A2(new_n488_), .B(new_n556_), .ZN(new_n2985_));
  AOI21_X1   g2600(.A1(new_n2985_), .A2(new_n562_), .B(new_n567_), .ZN(new_n2986_));
  OAI21_X1   g2601(.A1(new_n2986_), .A2(new_n484_), .B(new_n572_), .ZN(new_n2987_));
  OAI21_X1   g2602(.A1(new_n574_), .A2(\priority[32] ), .B(\req[32] ), .ZN(new_n2988_));
  AOI21_X1   g2603(.A1(new_n2987_), .A2(new_n480_), .B(new_n2988_), .ZN(\grant[32] ));
  NOR2_X1    g2604(.A1(new_n972_), .A2(new_n586_), .ZN(new_n2990_));
  OAI21_X1   g2605(.A1(new_n474_), .A2(new_n2990_), .B(new_n592_), .ZN(new_n2991_));
  AOI21_X1   g2606(.A1(new_n2991_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n2992_));
  OAI21_X1   g2607(.A1(new_n2992_), .A2(new_n603_), .B(new_n608_), .ZN(new_n2993_));
  AOI21_X1   g2608(.A1(new_n2993_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n2994_));
  OAI21_X1   g2609(.A1(new_n2994_), .A2(new_n461_), .B(new_n619_), .ZN(new_n2995_));
  AOI21_X1   g2610(.A1(new_n2995_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n2996_));
  OAI21_X1   g2611(.A1(new_n2996_), .A2(new_n456_), .B(new_n634_), .ZN(new_n2997_));
  AOI21_X1   g2612(.A1(new_n2997_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n2998_));
  OAI21_X1   g2613(.A1(new_n2998_), .A2(new_n645_), .B(new_n650_), .ZN(new_n2999_));
  AOI21_X1   g2614(.A1(new_n2999_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n3000_));
  OAI21_X1   g2615(.A1(new_n3000_), .A2(new_n443_), .B(new_n661_), .ZN(new_n3001_));
  AOI21_X1   g2616(.A1(new_n3001_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n3002_));
  OAI21_X1   g2617(.A1(new_n3002_), .A2(new_n438_), .B(new_n676_), .ZN(new_n3003_));
  AOI21_X1   g2618(.A1(new_n3003_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n3004_));
  OAI21_X1   g2619(.A1(new_n3004_), .A2(new_n687_), .B(new_n692_), .ZN(new_n3005_));
  AOI21_X1   g2620(.A1(new_n3005_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n3006_));
  OAI21_X1   g2621(.A1(new_n3006_), .A2(new_n425_), .B(new_n703_), .ZN(new_n3007_));
  AOI21_X1   g2622(.A1(new_n3007_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n3008_));
  OAI21_X1   g2623(.A1(new_n3008_), .A2(new_n420_), .B(new_n718_), .ZN(new_n3009_));
  AOI21_X1   g2624(.A1(new_n3009_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n3010_));
  OAI21_X1   g2625(.A1(new_n3010_), .A2(new_n729_), .B(new_n734_), .ZN(new_n3011_));
  AOI21_X1   g2626(.A1(new_n3011_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n3012_));
  OAI21_X1   g2627(.A1(new_n3012_), .A2(new_n407_), .B(new_n745_), .ZN(new_n3013_));
  AOI21_X1   g2628(.A1(new_n3013_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n3014_));
  OAI21_X1   g2629(.A1(new_n3014_), .A2(new_n402_), .B(new_n760_), .ZN(new_n3015_));
  AOI21_X1   g2630(.A1(new_n3015_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n3016_));
  OAI21_X1   g2631(.A1(new_n3016_), .A2(new_n771_), .B(new_n776_), .ZN(new_n3017_));
  AOI21_X1   g2632(.A1(new_n3017_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n3018_));
  OAI21_X1   g2633(.A1(new_n3018_), .A2(new_n389_), .B(new_n787_), .ZN(new_n3019_));
  AOI21_X1   g2634(.A1(new_n3019_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n3020_));
  OAI21_X1   g2635(.A1(new_n3020_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n3021_));
  AOI21_X1   g2636(.A1(new_n3021_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n3022_));
  OAI21_X1   g2637(.A1(new_n3022_), .A2(new_n900_), .B(new_n908_), .ZN(new_n3023_));
  AOI21_X1   g2638(.A1(new_n3023_), .A2(new_n913_), .B(new_n918_), .ZN(new_n3024_));
  OAI21_X1   g2639(.A1(new_n3024_), .A2(new_n897_), .B(new_n923_), .ZN(new_n3025_));
  AOI21_X1   g2640(.A1(new_n3025_), .A2(new_n894_), .B(new_n929_), .ZN(new_n3026_));
  OAI21_X1   g2641(.A1(new_n3026_), .A2(new_n933_), .B(new_n937_), .ZN(new_n3027_));
  AOI21_X1   g2642(.A1(new_n3027_), .A2(new_n890_), .B(new_n943_), .ZN(new_n3028_));
  OAI21_X1   g2643(.A1(new_n3028_), .A2(new_n886_), .B(new_n948_), .ZN(new_n3029_));
  AOI21_X1   g2644(.A1(new_n3029_), .A2(new_n953_), .B(new_n958_), .ZN(new_n3030_));
  OAI21_X1   g2645(.A1(new_n3030_), .A2(new_n883_), .B(new_n963_), .ZN(new_n3031_));
  OAI21_X1   g2646(.A1(new_n965_), .A2(\priority[33] ), .B(\req[33] ), .ZN(new_n3032_));
  AOI21_X1   g2647(.A1(new_n3031_), .A2(new_n880_), .B(new_n3032_), .ZN(\grant[33] ));
  NOR2_X1    g2648(.A1(new_n1343_), .A2(new_n976_), .ZN(new_n3034_));
  OAI21_X1   g2649(.A1(new_n875_), .A2(new_n3034_), .B(new_n982_), .ZN(new_n3035_));
  AOI21_X1   g2650(.A1(new_n3035_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n3036_));
  OAI21_X1   g2651(.A1(new_n3036_), .A2(new_n992_), .B(new_n997_), .ZN(new_n3037_));
  AOI21_X1   g2652(.A1(new_n3037_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n3038_));
  OAI21_X1   g2653(.A1(new_n3038_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n3039_));
  AOI21_X1   g2654(.A1(new_n3039_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n3040_));
  OAI21_X1   g2655(.A1(new_n3040_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n3041_));
  AOI21_X1   g2656(.A1(new_n3041_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n3042_));
  OAI21_X1   g2657(.A1(new_n3042_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n3043_));
  AOI21_X1   g2658(.A1(new_n3043_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n3044_));
  OAI21_X1   g2659(.A1(new_n3044_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n3045_));
  AOI21_X1   g2660(.A1(new_n3045_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n3046_));
  OAI21_X1   g2661(.A1(new_n3046_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n3047_));
  AOI21_X1   g2662(.A1(new_n3047_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n3048_));
  OAI21_X1   g2663(.A1(new_n3048_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n3049_));
  AOI21_X1   g2664(.A1(new_n3049_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n3050_));
  OAI21_X1   g2665(.A1(new_n3050_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n3051_));
  AOI21_X1   g2666(.A1(new_n3051_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n3052_));
  OAI21_X1   g2667(.A1(new_n3052_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n3053_));
  AOI21_X1   g2668(.A1(new_n3053_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n3054_));
  OAI21_X1   g2669(.A1(new_n3054_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n3055_));
  AOI21_X1   g2670(.A1(new_n3055_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n3056_));
  OAI21_X1   g2671(.A1(new_n3056_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n3057_));
  AOI21_X1   g2672(.A1(new_n3057_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n3058_));
  OAI21_X1   g2673(.A1(new_n3058_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n3059_));
  AOI21_X1   g2674(.A1(new_n3059_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n3060_));
  OAI21_X1   g2675(.A1(new_n3060_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n3061_));
  AOI21_X1   g2676(.A1(new_n3061_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n3062_));
  OAI21_X1   g2677(.A1(new_n3062_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n3063_));
  AOI21_X1   g2678(.A1(new_n3063_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n3064_));
  OAI21_X1   g2679(.A1(new_n3064_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n3065_));
  AOI21_X1   g2680(.A1(new_n3065_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n3066_));
  OAI21_X1   g2681(.A1(new_n3066_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n3067_));
  AOI21_X1   g2682(.A1(new_n3067_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n3068_));
  OAI21_X1   g2683(.A1(new_n3068_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n3069_));
  AOI21_X1   g2684(.A1(new_n3069_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n3070_));
  OAI21_X1   g2685(.A1(new_n3070_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n3071_));
  AOI21_X1   g2686(.A1(new_n3071_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n3072_));
  OAI21_X1   g2687(.A1(new_n3072_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n3073_));
  AOI21_X1   g2688(.A1(new_n3073_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n3074_));
  OAI21_X1   g2689(.A1(new_n3074_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n3075_));
  OAI21_X1   g2690(.A1(new_n581_), .A2(\priority[34] ), .B(\req[34] ), .ZN(new_n3076_));
  AOI21_X1   g2691(.A1(new_n3075_), .A2(new_n1263_), .B(new_n3076_), .ZN(\grant[34] ));
  NOR2_X1    g2692(.A1(new_n473_), .A2(new_n1346_), .ZN(new_n3078_));
  OAI21_X1   g2693(.A1(new_n1258_), .A2(new_n3078_), .B(new_n1351_), .ZN(new_n3079_));
  AOI21_X1   g2694(.A1(new_n3079_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n3080_));
  OAI21_X1   g2695(.A1(new_n3080_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n3081_));
  AOI21_X1   g2696(.A1(new_n3081_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n3082_));
  OAI21_X1   g2697(.A1(new_n3082_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n3083_));
  AOI21_X1   g2698(.A1(new_n3083_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n3084_));
  OAI21_X1   g2699(.A1(new_n3084_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n3085_));
  AOI21_X1   g2700(.A1(new_n3085_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n3086_));
  OAI21_X1   g2701(.A1(new_n3086_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n3087_));
  AOI21_X1   g2702(.A1(new_n3087_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n3088_));
  OAI21_X1   g2703(.A1(new_n3088_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n3089_));
  AOI21_X1   g2704(.A1(new_n3089_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n3090_));
  OAI21_X1   g2705(.A1(new_n3090_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n3091_));
  AOI21_X1   g2706(.A1(new_n3091_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n3092_));
  OAI21_X1   g2707(.A1(new_n3092_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n3093_));
  AOI21_X1   g2708(.A1(new_n3093_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n3094_));
  OAI21_X1   g2709(.A1(new_n3094_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n3095_));
  AOI21_X1   g2710(.A1(new_n3095_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n3096_));
  OAI21_X1   g2711(.A1(new_n3096_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n3097_));
  AOI21_X1   g2712(.A1(new_n3097_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n3098_));
  OAI21_X1   g2713(.A1(new_n3098_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n3099_));
  AOI21_X1   g2714(.A1(new_n3099_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n3100_));
  OAI21_X1   g2715(.A1(new_n3100_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n3101_));
  AOI21_X1   g2716(.A1(new_n3101_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n3102_));
  OAI21_X1   g2717(.A1(new_n3102_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n3103_));
  AOI21_X1   g2718(.A1(new_n3103_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n3104_));
  OAI21_X1   g2719(.A1(new_n3104_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n3105_));
  AOI21_X1   g2720(.A1(new_n3105_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n3106_));
  OAI21_X1   g2721(.A1(new_n3106_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n3107_));
  AOI21_X1   g2722(.A1(new_n3107_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n3108_));
  OAI21_X1   g2723(.A1(new_n3108_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n3109_));
  AOI21_X1   g2724(.A1(new_n3109_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n3110_));
  OAI21_X1   g2725(.A1(new_n3110_), .A2(new_n519_), .B(new_n524_), .ZN(new_n3111_));
  AOI21_X1   g2726(.A1(new_n3111_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n3112_));
  OAI21_X1   g2727(.A1(new_n3112_), .A2(new_n497_), .B(new_n535_), .ZN(new_n3113_));
  AOI21_X1   g2728(.A1(new_n3113_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n3114_));
  OAI21_X1   g2729(.A1(new_n3114_), .A2(new_n492_), .B(new_n550_), .ZN(new_n3115_));
  AOI21_X1   g2730(.A1(new_n3115_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n3116_));
  OAI21_X1   g2731(.A1(new_n3116_), .A2(new_n561_), .B(new_n566_), .ZN(new_n3117_));
  AOI21_X1   g2732(.A1(new_n3117_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n3118_));
  OAI21_X1   g2733(.A1(new_n3118_), .A2(new_n479_), .B(new_n577_), .ZN(new_n3119_));
  OAI21_X1   g2734(.A1(new_n584_), .A2(\priority[35] ), .B(\req[35] ), .ZN(new_n3120_));
  AOI21_X1   g2735(.A1(new_n3119_), .A2(new_n1554_), .B(new_n3120_), .ZN(\grant[35] ));
  NOR2_X1    g2736(.A1(new_n874_), .A2(new_n591_), .ZN(new_n3122_));
  OAI21_X1   g2737(.A1(new_n470_), .A2(new_n3122_), .B(new_n598_), .ZN(new_n3123_));
  AOI21_X1   g2738(.A1(new_n3123_), .A2(new_n604_), .B(new_n609_), .ZN(new_n3124_));
  OAI21_X1   g2739(.A1(new_n3124_), .A2(new_n466_), .B(new_n614_), .ZN(new_n3125_));
  AOI21_X1   g2740(.A1(new_n3125_), .A2(new_n462_), .B(new_n620_), .ZN(new_n3126_));
  OAI21_X1   g2741(.A1(new_n3126_), .A2(new_n625_), .B(new_n629_), .ZN(new_n3127_));
  AOI21_X1   g2742(.A1(new_n3127_), .A2(new_n457_), .B(new_n635_), .ZN(new_n3128_));
  OAI21_X1   g2743(.A1(new_n3128_), .A2(new_n452_), .B(new_n640_), .ZN(new_n3129_));
  AOI21_X1   g2744(.A1(new_n3129_), .A2(new_n646_), .B(new_n651_), .ZN(new_n3130_));
  OAI21_X1   g2745(.A1(new_n3130_), .A2(new_n448_), .B(new_n656_), .ZN(new_n3131_));
  AOI21_X1   g2746(.A1(new_n3131_), .A2(new_n444_), .B(new_n662_), .ZN(new_n3132_));
  OAI21_X1   g2747(.A1(new_n3132_), .A2(new_n667_), .B(new_n671_), .ZN(new_n3133_));
  AOI21_X1   g2748(.A1(new_n3133_), .A2(new_n439_), .B(new_n677_), .ZN(new_n3134_));
  OAI21_X1   g2749(.A1(new_n3134_), .A2(new_n434_), .B(new_n682_), .ZN(new_n3135_));
  AOI21_X1   g2750(.A1(new_n3135_), .A2(new_n688_), .B(new_n693_), .ZN(new_n3136_));
  OAI21_X1   g2751(.A1(new_n3136_), .A2(new_n430_), .B(new_n698_), .ZN(new_n3137_));
  AOI21_X1   g2752(.A1(new_n3137_), .A2(new_n426_), .B(new_n704_), .ZN(new_n3138_));
  OAI21_X1   g2753(.A1(new_n3138_), .A2(new_n709_), .B(new_n713_), .ZN(new_n3139_));
  AOI21_X1   g2754(.A1(new_n3139_), .A2(new_n421_), .B(new_n719_), .ZN(new_n3140_));
  OAI21_X1   g2755(.A1(new_n3140_), .A2(new_n416_), .B(new_n724_), .ZN(new_n3141_));
  AOI21_X1   g2756(.A1(new_n3141_), .A2(new_n730_), .B(new_n735_), .ZN(new_n3142_));
  OAI21_X1   g2757(.A1(new_n3142_), .A2(new_n412_), .B(new_n740_), .ZN(new_n3143_));
  AOI21_X1   g2758(.A1(new_n3143_), .A2(new_n408_), .B(new_n746_), .ZN(new_n3144_));
  OAI21_X1   g2759(.A1(new_n3144_), .A2(new_n751_), .B(new_n755_), .ZN(new_n3145_));
  AOI21_X1   g2760(.A1(new_n3145_), .A2(new_n403_), .B(new_n761_), .ZN(new_n3146_));
  OAI21_X1   g2761(.A1(new_n3146_), .A2(new_n398_), .B(new_n766_), .ZN(new_n3147_));
  AOI21_X1   g2762(.A1(new_n3147_), .A2(new_n772_), .B(new_n777_), .ZN(new_n3148_));
  OAI21_X1   g2763(.A1(new_n3148_), .A2(new_n394_), .B(new_n782_), .ZN(new_n3149_));
  AOI21_X1   g2764(.A1(new_n3149_), .A2(new_n390_), .B(new_n788_), .ZN(new_n3150_));
  OAI21_X1   g2765(.A1(new_n3150_), .A2(new_n793_), .B(new_n797_), .ZN(new_n3151_));
  AOI21_X1   g2766(.A1(new_n3151_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n3152_));
  OAI21_X1   g2767(.A1(new_n3152_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n3153_));
  AOI21_X1   g2768(.A1(new_n3153_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n3154_));
  OAI21_X1   g2769(.A1(new_n3154_), .A2(new_n912_), .B(new_n917_), .ZN(new_n3155_));
  AOI21_X1   g2770(.A1(new_n3155_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n3156_));
  OAI21_X1   g2771(.A1(new_n3156_), .A2(new_n893_), .B(new_n928_), .ZN(new_n3157_));
  AOI21_X1   g2772(.A1(new_n3157_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n3158_));
  OAI21_X1   g2773(.A1(new_n3158_), .A2(new_n889_), .B(new_n942_), .ZN(new_n3159_));
  AOI21_X1   g2774(.A1(new_n3159_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n3160_));
  OAI21_X1   g2775(.A1(new_n3160_), .A2(new_n952_), .B(new_n957_), .ZN(new_n3161_));
  AOI21_X1   g2776(.A1(new_n3161_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n3162_));
  OAI21_X1   g2777(.A1(new_n3162_), .A2(new_n879_), .B(new_n968_), .ZN(new_n3163_));
  OAI21_X1   g2778(.A1(new_n974_), .A2(\priority[36] ), .B(\req[36] ), .ZN(new_n3164_));
  AOI21_X1   g2779(.A1(new_n3163_), .A2(new_n1644_), .B(new_n3164_), .ZN(\grant[36] ));
  NOR2_X1    g2780(.A1(new_n1257_), .A2(new_n981_), .ZN(new_n3166_));
  OAI21_X1   g2781(.A1(new_n872_), .A2(new_n3166_), .B(new_n988_), .ZN(new_n3167_));
  AOI21_X1   g2782(.A1(new_n3167_), .A2(new_n993_), .B(new_n998_), .ZN(new_n3168_));
  OAI21_X1   g2783(.A1(new_n3168_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n3169_));
  AOI21_X1   g2784(.A1(new_n3169_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n3170_));
  OAI21_X1   g2785(.A1(new_n3170_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n3171_));
  AOI21_X1   g2786(.A1(new_n3171_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n3172_));
  OAI21_X1   g2787(.A1(new_n3172_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n3173_));
  AOI21_X1   g2788(.A1(new_n3173_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n3174_));
  OAI21_X1   g2789(.A1(new_n3174_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n3175_));
  AOI21_X1   g2790(.A1(new_n3175_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n3176_));
  OAI21_X1   g2791(.A1(new_n3176_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n3177_));
  AOI21_X1   g2792(.A1(new_n3177_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n3178_));
  OAI21_X1   g2793(.A1(new_n3178_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n3179_));
  AOI21_X1   g2794(.A1(new_n3179_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n3180_));
  OAI21_X1   g2795(.A1(new_n3180_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n3181_));
  AOI21_X1   g2796(.A1(new_n3181_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n3182_));
  OAI21_X1   g2797(.A1(new_n3182_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n3183_));
  AOI21_X1   g2798(.A1(new_n3183_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n3184_));
  OAI21_X1   g2799(.A1(new_n3184_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n3185_));
  AOI21_X1   g2800(.A1(new_n3185_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n3186_));
  OAI21_X1   g2801(.A1(new_n3186_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n3187_));
  AOI21_X1   g2802(.A1(new_n3187_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n3188_));
  OAI21_X1   g2803(.A1(new_n3188_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n3189_));
  AOI21_X1   g2804(.A1(new_n3189_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n3190_));
  OAI21_X1   g2805(.A1(new_n3190_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n3191_));
  AOI21_X1   g2806(.A1(new_n3191_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n3192_));
  OAI21_X1   g2807(.A1(new_n3192_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n3193_));
  AOI21_X1   g2808(.A1(new_n3193_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n3194_));
  OAI21_X1   g2809(.A1(new_n3194_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n3195_));
  AOI21_X1   g2810(.A1(new_n3195_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n3196_));
  OAI21_X1   g2811(.A1(new_n3196_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n3197_));
  AOI21_X1   g2812(.A1(new_n3197_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n3198_));
  OAI21_X1   g2813(.A1(new_n3198_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n3199_));
  AOI21_X1   g2814(.A1(new_n3199_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n3200_));
  OAI21_X1   g2815(.A1(new_n3200_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n3201_));
  AOI21_X1   g2816(.A1(new_n3201_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n3202_));
  OAI21_X1   g2817(.A1(new_n3202_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n3203_));
  AOI21_X1   g2818(.A1(new_n3203_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n3204_));
  OAI21_X1   g2819(.A1(new_n3204_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n3205_));
  AOI21_X1   g2820(.A1(new_n3205_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n3206_));
  OAI21_X1   g2821(.A1(new_n3206_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n3207_));
  OAI21_X1   g2822(.A1(new_n472_), .A2(\priority[37] ), .B(\req[37] ), .ZN(new_n3208_));
  AOI21_X1   g2823(.A1(new_n3207_), .A2(new_n1732_), .B(new_n3208_), .ZN(\grant[37] ));
  NOR2_X1    g2824(.A1(new_n469_), .A2(new_n1350_), .ZN(new_n3210_));
  OAI21_X1   g2825(.A1(new_n1255_), .A2(new_n3210_), .B(new_n1356_), .ZN(new_n3211_));
  AOI21_X1   g2826(.A1(new_n3211_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n3212_));
  OAI21_X1   g2827(.A1(new_n3212_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n3213_));
  AOI21_X1   g2828(.A1(new_n3213_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n3214_));
  OAI21_X1   g2829(.A1(new_n3214_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n3215_));
  AOI21_X1   g2830(.A1(new_n3215_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n3216_));
  OAI21_X1   g2831(.A1(new_n3216_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n3217_));
  AOI21_X1   g2832(.A1(new_n3217_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n3218_));
  OAI21_X1   g2833(.A1(new_n3218_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n3219_));
  AOI21_X1   g2834(.A1(new_n3219_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n3220_));
  OAI21_X1   g2835(.A1(new_n3220_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n3221_));
  AOI21_X1   g2836(.A1(new_n3221_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n3222_));
  OAI21_X1   g2837(.A1(new_n3222_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n3223_));
  AOI21_X1   g2838(.A1(new_n3223_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n3224_));
  OAI21_X1   g2839(.A1(new_n3224_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n3225_));
  AOI21_X1   g2840(.A1(new_n3225_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n3226_));
  OAI21_X1   g2841(.A1(new_n3226_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n3227_));
  AOI21_X1   g2842(.A1(new_n3227_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n3228_));
  OAI21_X1   g2843(.A1(new_n3228_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n3229_));
  AOI21_X1   g2844(.A1(new_n3229_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n3230_));
  OAI21_X1   g2845(.A1(new_n3230_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n3231_));
  AOI21_X1   g2846(.A1(new_n3231_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n3232_));
  OAI21_X1   g2847(.A1(new_n3232_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n3233_));
  AOI21_X1   g2848(.A1(new_n3233_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n3234_));
  OAI21_X1   g2849(.A1(new_n3234_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n3235_));
  AOI21_X1   g2850(.A1(new_n3235_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n3236_));
  OAI21_X1   g2851(.A1(new_n3236_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n3237_));
  AOI21_X1   g2852(.A1(new_n3237_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n3238_));
  OAI21_X1   g2853(.A1(new_n3238_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n3239_));
  AOI21_X1   g2854(.A1(new_n3239_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n3240_));
  OAI21_X1   g2855(.A1(new_n3240_), .A2(new_n506_), .B(new_n514_), .ZN(new_n3241_));
  AOI21_X1   g2856(.A1(new_n3241_), .A2(new_n520_), .B(new_n525_), .ZN(new_n3242_));
  OAI21_X1   g2857(.A1(new_n3242_), .A2(new_n502_), .B(new_n530_), .ZN(new_n3243_));
  AOI21_X1   g2858(.A1(new_n3243_), .A2(new_n498_), .B(new_n536_), .ZN(new_n3244_));
  OAI21_X1   g2859(.A1(new_n3244_), .A2(new_n541_), .B(new_n545_), .ZN(new_n3245_));
  AOI21_X1   g2860(.A1(new_n3245_), .A2(new_n493_), .B(new_n551_), .ZN(new_n3246_));
  OAI21_X1   g2861(.A1(new_n3246_), .A2(new_n488_), .B(new_n556_), .ZN(new_n3247_));
  AOI21_X1   g2862(.A1(new_n3247_), .A2(new_n562_), .B(new_n567_), .ZN(new_n3248_));
  OAI21_X1   g2863(.A1(new_n3248_), .A2(new_n484_), .B(new_n572_), .ZN(new_n3249_));
  AOI21_X1   g2864(.A1(new_n3249_), .A2(new_n480_), .B(new_n578_), .ZN(new_n3250_));
  OAI21_X1   g2865(.A1(new_n3250_), .A2(new_n583_), .B(new_n587_), .ZN(new_n3251_));
  OAI21_X1   g2866(.A1(new_n589_), .A2(\priority[38] ), .B(\req[38] ), .ZN(new_n3252_));
  AOI21_X1   g2867(.A1(new_n3251_), .A2(new_n475_), .B(new_n3252_), .ZN(\grant[38] ));
  NOR2_X1    g2868(.A1(new_n871_), .A2(new_n597_), .ZN(new_n3254_));
  OAI21_X1   g2869(.A1(new_n603_), .A2(new_n3254_), .B(new_n608_), .ZN(new_n3255_));
  AOI21_X1   g2870(.A1(new_n3255_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n3256_));
  OAI21_X1   g2871(.A1(new_n3256_), .A2(new_n461_), .B(new_n619_), .ZN(new_n3257_));
  AOI21_X1   g2872(.A1(new_n3257_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n3258_));
  OAI21_X1   g2873(.A1(new_n3258_), .A2(new_n456_), .B(new_n634_), .ZN(new_n3259_));
  AOI21_X1   g2874(.A1(new_n3259_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n3260_));
  OAI21_X1   g2875(.A1(new_n3260_), .A2(new_n645_), .B(new_n650_), .ZN(new_n3261_));
  AOI21_X1   g2876(.A1(new_n3261_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n3262_));
  OAI21_X1   g2877(.A1(new_n3262_), .A2(new_n443_), .B(new_n661_), .ZN(new_n3263_));
  AOI21_X1   g2878(.A1(new_n3263_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n3264_));
  OAI21_X1   g2879(.A1(new_n3264_), .A2(new_n438_), .B(new_n676_), .ZN(new_n3265_));
  AOI21_X1   g2880(.A1(new_n3265_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n3266_));
  OAI21_X1   g2881(.A1(new_n3266_), .A2(new_n687_), .B(new_n692_), .ZN(new_n3267_));
  AOI21_X1   g2882(.A1(new_n3267_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n3268_));
  OAI21_X1   g2883(.A1(new_n3268_), .A2(new_n425_), .B(new_n703_), .ZN(new_n3269_));
  AOI21_X1   g2884(.A1(new_n3269_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n3270_));
  OAI21_X1   g2885(.A1(new_n3270_), .A2(new_n420_), .B(new_n718_), .ZN(new_n3271_));
  AOI21_X1   g2886(.A1(new_n3271_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n3272_));
  OAI21_X1   g2887(.A1(new_n3272_), .A2(new_n729_), .B(new_n734_), .ZN(new_n3273_));
  AOI21_X1   g2888(.A1(new_n3273_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n3274_));
  OAI21_X1   g2889(.A1(new_n3274_), .A2(new_n407_), .B(new_n745_), .ZN(new_n3275_));
  AOI21_X1   g2890(.A1(new_n3275_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n3276_));
  OAI21_X1   g2891(.A1(new_n3276_), .A2(new_n402_), .B(new_n760_), .ZN(new_n3277_));
  AOI21_X1   g2892(.A1(new_n3277_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n3278_));
  OAI21_X1   g2893(.A1(new_n3278_), .A2(new_n771_), .B(new_n776_), .ZN(new_n3279_));
  AOI21_X1   g2894(.A1(new_n3279_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n3280_));
  OAI21_X1   g2895(.A1(new_n3280_), .A2(new_n389_), .B(new_n787_), .ZN(new_n3281_));
  AOI21_X1   g2896(.A1(new_n3281_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n3282_));
  OAI21_X1   g2897(.A1(new_n3282_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n3283_));
  AOI21_X1   g2898(.A1(new_n3283_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n3284_));
  OAI21_X1   g2899(.A1(new_n3284_), .A2(new_n900_), .B(new_n908_), .ZN(new_n3285_));
  AOI21_X1   g2900(.A1(new_n3285_), .A2(new_n913_), .B(new_n918_), .ZN(new_n3286_));
  OAI21_X1   g2901(.A1(new_n3286_), .A2(new_n897_), .B(new_n923_), .ZN(new_n3287_));
  AOI21_X1   g2902(.A1(new_n3287_), .A2(new_n894_), .B(new_n929_), .ZN(new_n3288_));
  OAI21_X1   g2903(.A1(new_n3288_), .A2(new_n933_), .B(new_n937_), .ZN(new_n3289_));
  AOI21_X1   g2904(.A1(new_n3289_), .A2(new_n890_), .B(new_n943_), .ZN(new_n3290_));
  OAI21_X1   g2905(.A1(new_n3290_), .A2(new_n886_), .B(new_n948_), .ZN(new_n3291_));
  AOI21_X1   g2906(.A1(new_n3291_), .A2(new_n953_), .B(new_n958_), .ZN(new_n3292_));
  OAI21_X1   g2907(.A1(new_n3292_), .A2(new_n883_), .B(new_n963_), .ZN(new_n3293_));
  AOI21_X1   g2908(.A1(new_n3293_), .A2(new_n880_), .B(new_n969_), .ZN(new_n3294_));
  OAI21_X1   g2909(.A1(new_n3294_), .A2(new_n973_), .B(new_n977_), .ZN(new_n3295_));
  OAI21_X1   g2910(.A1(new_n979_), .A2(\priority[39] ), .B(\req[39] ), .ZN(new_n3296_));
  AOI21_X1   g2911(.A1(new_n3295_), .A2(new_n876_), .B(new_n3296_), .ZN(\grant[39] ));
  NOR2_X1    g2912(.A1(new_n1254_), .A2(new_n987_), .ZN(new_n3298_));
  OAI21_X1   g2913(.A1(new_n992_), .A2(new_n3298_), .B(new_n997_), .ZN(new_n3299_));
  AOI21_X1   g2914(.A1(new_n3299_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n3300_));
  OAI21_X1   g2915(.A1(new_n3300_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n3301_));
  AOI21_X1   g2916(.A1(new_n3301_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n3302_));
  OAI21_X1   g2917(.A1(new_n3302_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n3303_));
  AOI21_X1   g2918(.A1(new_n3303_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n3304_));
  OAI21_X1   g2919(.A1(new_n3304_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n3305_));
  AOI21_X1   g2920(.A1(new_n3305_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n3306_));
  OAI21_X1   g2921(.A1(new_n3306_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n3307_));
  AOI21_X1   g2922(.A1(new_n3307_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n3308_));
  OAI21_X1   g2923(.A1(new_n3308_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n3309_));
  AOI21_X1   g2924(.A1(new_n3309_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n3310_));
  OAI21_X1   g2925(.A1(new_n3310_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n3311_));
  AOI21_X1   g2926(.A1(new_n3311_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n3312_));
  OAI21_X1   g2927(.A1(new_n3312_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n3313_));
  AOI21_X1   g2928(.A1(new_n3313_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n3314_));
  OAI21_X1   g2929(.A1(new_n3314_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n3315_));
  AOI21_X1   g2930(.A1(new_n3315_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n3316_));
  OAI21_X1   g2931(.A1(new_n3316_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n3317_));
  AOI21_X1   g2932(.A1(new_n3317_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n3318_));
  OAI21_X1   g2933(.A1(new_n3318_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n3319_));
  AOI21_X1   g2934(.A1(new_n3319_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n3320_));
  OAI21_X1   g2935(.A1(new_n3320_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n3321_));
  AOI21_X1   g2936(.A1(new_n3321_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n3322_));
  OAI21_X1   g2937(.A1(new_n3322_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n3323_));
  AOI21_X1   g2938(.A1(new_n3323_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n3324_));
  OAI21_X1   g2939(.A1(new_n3324_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n3325_));
  AOI21_X1   g2940(.A1(new_n3325_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n3326_));
  OAI21_X1   g2941(.A1(new_n3326_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n3327_));
  AOI21_X1   g2942(.A1(new_n3327_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n3328_));
  OAI21_X1   g2943(.A1(new_n3328_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n3329_));
  AOI21_X1   g2944(.A1(new_n3329_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n3330_));
  OAI21_X1   g2945(.A1(new_n3330_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n3331_));
  AOI21_X1   g2946(.A1(new_n3331_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n3332_));
  OAI21_X1   g2947(.A1(new_n3332_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n3333_));
  AOI21_X1   g2948(.A1(new_n3333_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n3334_));
  OAI21_X1   g2949(.A1(new_n3334_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n3335_));
  AOI21_X1   g2950(.A1(new_n3335_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n3336_));
  OAI21_X1   g2951(.A1(new_n3336_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n3337_));
  AOI21_X1   g2952(.A1(new_n3337_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n3338_));
  OAI21_X1   g2953(.A1(new_n3338_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n3339_));
  OAI21_X1   g2954(.A1(new_n468_), .A2(\priority[40] ), .B(\req[40] ), .ZN(new_n3340_));
  AOI21_X1   g2955(.A1(new_n3339_), .A2(new_n1259_), .B(new_n3340_), .ZN(\grant[40] ));
  NOR2_X1    g2956(.A1(new_n602_), .A2(new_n1355_), .ZN(new_n3342_));
  OAI21_X1   g2957(.A1(new_n1360_), .A2(new_n3342_), .B(new_n1364_), .ZN(new_n3343_));
  AOI21_X1   g2958(.A1(new_n3343_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n3344_));
  OAI21_X1   g2959(.A1(new_n3344_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n3345_));
  AOI21_X1   g2960(.A1(new_n3345_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n3346_));
  OAI21_X1   g2961(.A1(new_n3346_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n3347_));
  AOI21_X1   g2962(.A1(new_n3347_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n3348_));
  OAI21_X1   g2963(.A1(new_n3348_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n3349_));
  AOI21_X1   g2964(.A1(new_n3349_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n3350_));
  OAI21_X1   g2965(.A1(new_n3350_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n3351_));
  AOI21_X1   g2966(.A1(new_n3351_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n3352_));
  OAI21_X1   g2967(.A1(new_n3352_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n3353_));
  AOI21_X1   g2968(.A1(new_n3353_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n3354_));
  OAI21_X1   g2969(.A1(new_n3354_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n3355_));
  AOI21_X1   g2970(.A1(new_n3355_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n3356_));
  OAI21_X1   g2971(.A1(new_n3356_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n3357_));
  AOI21_X1   g2972(.A1(new_n3357_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n3358_));
  OAI21_X1   g2973(.A1(new_n3358_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n3359_));
  AOI21_X1   g2974(.A1(new_n3359_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n3360_));
  OAI21_X1   g2975(.A1(new_n3360_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n3361_));
  AOI21_X1   g2976(.A1(new_n3361_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n3362_));
  OAI21_X1   g2977(.A1(new_n3362_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n3363_));
  AOI21_X1   g2978(.A1(new_n3363_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n3364_));
  OAI21_X1   g2979(.A1(new_n3364_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n3365_));
  AOI21_X1   g2980(.A1(new_n3365_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n3366_));
  OAI21_X1   g2981(.A1(new_n3366_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n3367_));
  AOI21_X1   g2982(.A1(new_n3367_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n3368_));
  OAI21_X1   g2983(.A1(new_n3368_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n3369_));
  AOI21_X1   g2984(.A1(new_n3369_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n3370_));
  OAI21_X1   g2985(.A1(new_n3370_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n3371_));
  AOI21_X1   g2986(.A1(new_n3371_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n3372_));
  OAI21_X1   g2987(.A1(new_n3372_), .A2(new_n519_), .B(new_n524_), .ZN(new_n3373_));
  AOI21_X1   g2988(.A1(new_n3373_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n3374_));
  OAI21_X1   g2989(.A1(new_n3374_), .A2(new_n497_), .B(new_n535_), .ZN(new_n3375_));
  AOI21_X1   g2990(.A1(new_n3375_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n3376_));
  OAI21_X1   g2991(.A1(new_n3376_), .A2(new_n492_), .B(new_n550_), .ZN(new_n3377_));
  AOI21_X1   g2992(.A1(new_n3377_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n3378_));
  OAI21_X1   g2993(.A1(new_n3378_), .A2(new_n561_), .B(new_n566_), .ZN(new_n3379_));
  AOI21_X1   g2994(.A1(new_n3379_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n3380_));
  OAI21_X1   g2995(.A1(new_n3380_), .A2(new_n479_), .B(new_n577_), .ZN(new_n3381_));
  AOI21_X1   g2996(.A1(new_n3381_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n3382_));
  OAI21_X1   g2997(.A1(new_n3382_), .A2(new_n474_), .B(new_n592_), .ZN(new_n3383_));
  OAI21_X1   g2998(.A1(new_n595_), .A2(\priority[41] ), .B(\req[41] ), .ZN(new_n3384_));
  AOI21_X1   g2999(.A1(new_n3383_), .A2(new_n1552_), .B(new_n3384_), .ZN(\grant[41] ));
  NOR2_X1    g3000(.A1(new_n991_), .A2(new_n607_), .ZN(new_n3386_));
  OAI21_X1   g3001(.A1(new_n466_), .A2(new_n3386_), .B(new_n614_), .ZN(new_n3387_));
  AOI21_X1   g3002(.A1(new_n3387_), .A2(new_n462_), .B(new_n620_), .ZN(new_n3388_));
  OAI21_X1   g3003(.A1(new_n3388_), .A2(new_n625_), .B(new_n629_), .ZN(new_n3389_));
  AOI21_X1   g3004(.A1(new_n3389_), .A2(new_n457_), .B(new_n635_), .ZN(new_n3390_));
  OAI21_X1   g3005(.A1(new_n3390_), .A2(new_n452_), .B(new_n640_), .ZN(new_n3391_));
  AOI21_X1   g3006(.A1(new_n3391_), .A2(new_n646_), .B(new_n651_), .ZN(new_n3392_));
  OAI21_X1   g3007(.A1(new_n3392_), .A2(new_n448_), .B(new_n656_), .ZN(new_n3393_));
  AOI21_X1   g3008(.A1(new_n3393_), .A2(new_n444_), .B(new_n662_), .ZN(new_n3394_));
  OAI21_X1   g3009(.A1(new_n3394_), .A2(new_n667_), .B(new_n671_), .ZN(new_n3395_));
  AOI21_X1   g3010(.A1(new_n3395_), .A2(new_n439_), .B(new_n677_), .ZN(new_n3396_));
  OAI21_X1   g3011(.A1(new_n3396_), .A2(new_n434_), .B(new_n682_), .ZN(new_n3397_));
  AOI21_X1   g3012(.A1(new_n3397_), .A2(new_n688_), .B(new_n693_), .ZN(new_n3398_));
  OAI21_X1   g3013(.A1(new_n3398_), .A2(new_n430_), .B(new_n698_), .ZN(new_n3399_));
  AOI21_X1   g3014(.A1(new_n3399_), .A2(new_n426_), .B(new_n704_), .ZN(new_n3400_));
  OAI21_X1   g3015(.A1(new_n3400_), .A2(new_n709_), .B(new_n713_), .ZN(new_n3401_));
  AOI21_X1   g3016(.A1(new_n3401_), .A2(new_n421_), .B(new_n719_), .ZN(new_n3402_));
  OAI21_X1   g3017(.A1(new_n3402_), .A2(new_n416_), .B(new_n724_), .ZN(new_n3403_));
  AOI21_X1   g3018(.A1(new_n3403_), .A2(new_n730_), .B(new_n735_), .ZN(new_n3404_));
  OAI21_X1   g3019(.A1(new_n3404_), .A2(new_n412_), .B(new_n740_), .ZN(new_n3405_));
  AOI21_X1   g3020(.A1(new_n3405_), .A2(new_n408_), .B(new_n746_), .ZN(new_n3406_));
  OAI21_X1   g3021(.A1(new_n3406_), .A2(new_n751_), .B(new_n755_), .ZN(new_n3407_));
  AOI21_X1   g3022(.A1(new_n3407_), .A2(new_n403_), .B(new_n761_), .ZN(new_n3408_));
  OAI21_X1   g3023(.A1(new_n3408_), .A2(new_n398_), .B(new_n766_), .ZN(new_n3409_));
  AOI21_X1   g3024(.A1(new_n3409_), .A2(new_n772_), .B(new_n777_), .ZN(new_n3410_));
  OAI21_X1   g3025(.A1(new_n3410_), .A2(new_n394_), .B(new_n782_), .ZN(new_n3411_));
  AOI21_X1   g3026(.A1(new_n3411_), .A2(new_n390_), .B(new_n788_), .ZN(new_n3412_));
  OAI21_X1   g3027(.A1(new_n3412_), .A2(new_n793_), .B(new_n797_), .ZN(new_n3413_));
  AOI21_X1   g3028(.A1(new_n3413_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n3414_));
  OAI21_X1   g3029(.A1(new_n3414_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n3415_));
  AOI21_X1   g3030(.A1(new_n3415_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n3416_));
  OAI21_X1   g3031(.A1(new_n3416_), .A2(new_n912_), .B(new_n917_), .ZN(new_n3417_));
  AOI21_X1   g3032(.A1(new_n3417_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n3418_));
  OAI21_X1   g3033(.A1(new_n3418_), .A2(new_n893_), .B(new_n928_), .ZN(new_n3419_));
  AOI21_X1   g3034(.A1(new_n3419_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n3420_));
  OAI21_X1   g3035(.A1(new_n3420_), .A2(new_n889_), .B(new_n942_), .ZN(new_n3421_));
  AOI21_X1   g3036(.A1(new_n3421_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n3422_));
  OAI21_X1   g3037(.A1(new_n3422_), .A2(new_n952_), .B(new_n957_), .ZN(new_n3423_));
  AOI21_X1   g3038(.A1(new_n3423_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n3424_));
  OAI21_X1   g3039(.A1(new_n3424_), .A2(new_n879_), .B(new_n968_), .ZN(new_n3425_));
  AOI21_X1   g3040(.A1(new_n3425_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n3426_));
  OAI21_X1   g3041(.A1(new_n3426_), .A2(new_n875_), .B(new_n982_), .ZN(new_n3427_));
  OAI21_X1   g3042(.A1(new_n985_), .A2(\priority[42] ), .B(\req[42] ), .ZN(new_n3428_));
  AOI21_X1   g3043(.A1(new_n3427_), .A2(new_n1642_), .B(new_n3428_), .ZN(\grant[42] ));
  NOR2_X1    g3044(.A1(new_n1359_), .A2(new_n996_), .ZN(new_n3430_));
  OAI21_X1   g3045(.A1(new_n869_), .A2(new_n3430_), .B(new_n1003_), .ZN(new_n3431_));
  AOI21_X1   g3046(.A1(new_n3431_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n3432_));
  OAI21_X1   g3047(.A1(new_n3432_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n3433_));
  AOI21_X1   g3048(.A1(new_n3433_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n3434_));
  OAI21_X1   g3049(.A1(new_n3434_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n3435_));
  AOI21_X1   g3050(.A1(new_n3435_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n3436_));
  OAI21_X1   g3051(.A1(new_n3436_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n3437_));
  AOI21_X1   g3052(.A1(new_n3437_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n3438_));
  OAI21_X1   g3053(.A1(new_n3438_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n3439_));
  AOI21_X1   g3054(.A1(new_n3439_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n3440_));
  OAI21_X1   g3055(.A1(new_n3440_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n3441_));
  AOI21_X1   g3056(.A1(new_n3441_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n3442_));
  OAI21_X1   g3057(.A1(new_n3442_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n3443_));
  AOI21_X1   g3058(.A1(new_n3443_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n3444_));
  OAI21_X1   g3059(.A1(new_n3444_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n3445_));
  AOI21_X1   g3060(.A1(new_n3445_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n3446_));
  OAI21_X1   g3061(.A1(new_n3446_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n3447_));
  AOI21_X1   g3062(.A1(new_n3447_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n3448_));
  OAI21_X1   g3063(.A1(new_n3448_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n3449_));
  AOI21_X1   g3064(.A1(new_n3449_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n3450_));
  OAI21_X1   g3065(.A1(new_n3450_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n3451_));
  AOI21_X1   g3066(.A1(new_n3451_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n3452_));
  OAI21_X1   g3067(.A1(new_n3452_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n3453_));
  AOI21_X1   g3068(.A1(new_n3453_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n3454_));
  OAI21_X1   g3069(.A1(new_n3454_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n3455_));
  AOI21_X1   g3070(.A1(new_n3455_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n3456_));
  OAI21_X1   g3071(.A1(new_n3456_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n3457_));
  AOI21_X1   g3072(.A1(new_n3457_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n3458_));
  OAI21_X1   g3073(.A1(new_n3458_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n3459_));
  AOI21_X1   g3074(.A1(new_n3459_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n3460_));
  OAI21_X1   g3075(.A1(new_n3460_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n3461_));
  AOI21_X1   g3076(.A1(new_n3461_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n3462_));
  OAI21_X1   g3077(.A1(new_n3462_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n3463_));
  AOI21_X1   g3078(.A1(new_n3463_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n3464_));
  OAI21_X1   g3079(.A1(new_n3464_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n3465_));
  AOI21_X1   g3080(.A1(new_n3465_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n3466_));
  OAI21_X1   g3081(.A1(new_n3466_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n3467_));
  AOI21_X1   g3082(.A1(new_n3467_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n3468_));
  OAI21_X1   g3083(.A1(new_n3468_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n3469_));
  AOI21_X1   g3084(.A1(new_n3469_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n3470_));
  OAI21_X1   g3085(.A1(new_n3470_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n3471_));
  OAI21_X1   g3086(.A1(new_n601_), .A2(\priority[43] ), .B(\req[43] ), .ZN(new_n3472_));
  AOI21_X1   g3087(.A1(new_n3471_), .A2(new_n1730_), .B(new_n3472_), .ZN(\grant[43] ));
  NOR2_X1    g3088(.A1(new_n465_), .A2(new_n1363_), .ZN(new_n3474_));
  OAI21_X1   g3089(.A1(new_n1252_), .A2(new_n3474_), .B(new_n1369_), .ZN(new_n3475_));
  AOI21_X1   g3090(.A1(new_n3475_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n3476_));
  OAI21_X1   g3091(.A1(new_n3476_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n3477_));
  AOI21_X1   g3092(.A1(new_n3477_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n3478_));
  OAI21_X1   g3093(.A1(new_n3478_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n3479_));
  AOI21_X1   g3094(.A1(new_n3479_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n3480_));
  OAI21_X1   g3095(.A1(new_n3480_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n3481_));
  AOI21_X1   g3096(.A1(new_n3481_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n3482_));
  OAI21_X1   g3097(.A1(new_n3482_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n3483_));
  AOI21_X1   g3098(.A1(new_n3483_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n3484_));
  OAI21_X1   g3099(.A1(new_n3484_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n3485_));
  AOI21_X1   g3100(.A1(new_n3485_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n3486_));
  OAI21_X1   g3101(.A1(new_n3486_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n3487_));
  AOI21_X1   g3102(.A1(new_n3487_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n3488_));
  OAI21_X1   g3103(.A1(new_n3488_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n3489_));
  AOI21_X1   g3104(.A1(new_n3489_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n3490_));
  OAI21_X1   g3105(.A1(new_n3490_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n3491_));
  AOI21_X1   g3106(.A1(new_n3491_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n3492_));
  OAI21_X1   g3107(.A1(new_n3492_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n3493_));
  AOI21_X1   g3108(.A1(new_n3493_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n3494_));
  OAI21_X1   g3109(.A1(new_n3494_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n3495_));
  AOI21_X1   g3110(.A1(new_n3495_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n3496_));
  OAI21_X1   g3111(.A1(new_n3496_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n3497_));
  AOI21_X1   g3112(.A1(new_n3497_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n3498_));
  OAI21_X1   g3113(.A1(new_n3498_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n3499_));
  AOI21_X1   g3114(.A1(new_n3499_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n3500_));
  OAI21_X1   g3115(.A1(new_n3500_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n3501_));
  AOI21_X1   g3116(.A1(new_n3501_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n3502_));
  OAI21_X1   g3117(.A1(new_n3502_), .A2(new_n506_), .B(new_n514_), .ZN(new_n3503_));
  AOI21_X1   g3118(.A1(new_n3503_), .A2(new_n520_), .B(new_n525_), .ZN(new_n3504_));
  OAI21_X1   g3119(.A1(new_n3504_), .A2(new_n502_), .B(new_n530_), .ZN(new_n3505_));
  AOI21_X1   g3120(.A1(new_n3505_), .A2(new_n498_), .B(new_n536_), .ZN(new_n3506_));
  OAI21_X1   g3121(.A1(new_n3506_), .A2(new_n541_), .B(new_n545_), .ZN(new_n3507_));
  AOI21_X1   g3122(.A1(new_n3507_), .A2(new_n493_), .B(new_n551_), .ZN(new_n3508_));
  OAI21_X1   g3123(.A1(new_n3508_), .A2(new_n488_), .B(new_n556_), .ZN(new_n3509_));
  AOI21_X1   g3124(.A1(new_n3509_), .A2(new_n562_), .B(new_n567_), .ZN(new_n3510_));
  OAI21_X1   g3125(.A1(new_n3510_), .A2(new_n484_), .B(new_n572_), .ZN(new_n3511_));
  AOI21_X1   g3126(.A1(new_n3511_), .A2(new_n480_), .B(new_n578_), .ZN(new_n3512_));
  OAI21_X1   g3127(.A1(new_n3512_), .A2(new_n583_), .B(new_n587_), .ZN(new_n3513_));
  AOI21_X1   g3128(.A1(new_n3513_), .A2(new_n475_), .B(new_n593_), .ZN(new_n3514_));
  OAI21_X1   g3129(.A1(new_n3514_), .A2(new_n470_), .B(new_n598_), .ZN(new_n3515_));
  OAI21_X1   g3130(.A1(new_n605_), .A2(\priority[44] ), .B(\req[44] ), .ZN(new_n3516_));
  AOI21_X1   g3131(.A1(new_n3515_), .A2(new_n604_), .B(new_n3516_), .ZN(\grant[44] ));
  NOR2_X1    g3132(.A1(new_n868_), .A2(new_n613_), .ZN(new_n3518_));
  OAI21_X1   g3133(.A1(new_n461_), .A2(new_n3518_), .B(new_n619_), .ZN(new_n3519_));
  AOI21_X1   g3134(.A1(new_n3519_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n3520_));
  OAI21_X1   g3135(.A1(new_n3520_), .A2(new_n456_), .B(new_n634_), .ZN(new_n3521_));
  AOI21_X1   g3136(.A1(new_n3521_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n3522_));
  OAI21_X1   g3137(.A1(new_n3522_), .A2(new_n645_), .B(new_n650_), .ZN(new_n3523_));
  AOI21_X1   g3138(.A1(new_n3523_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n3524_));
  OAI21_X1   g3139(.A1(new_n3524_), .A2(new_n443_), .B(new_n661_), .ZN(new_n3525_));
  AOI21_X1   g3140(.A1(new_n3525_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n3526_));
  OAI21_X1   g3141(.A1(new_n3526_), .A2(new_n438_), .B(new_n676_), .ZN(new_n3527_));
  AOI21_X1   g3142(.A1(new_n3527_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n3528_));
  OAI21_X1   g3143(.A1(new_n3528_), .A2(new_n687_), .B(new_n692_), .ZN(new_n3529_));
  AOI21_X1   g3144(.A1(new_n3529_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n3530_));
  OAI21_X1   g3145(.A1(new_n3530_), .A2(new_n425_), .B(new_n703_), .ZN(new_n3531_));
  AOI21_X1   g3146(.A1(new_n3531_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n3532_));
  OAI21_X1   g3147(.A1(new_n3532_), .A2(new_n420_), .B(new_n718_), .ZN(new_n3533_));
  AOI21_X1   g3148(.A1(new_n3533_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n3534_));
  OAI21_X1   g3149(.A1(new_n3534_), .A2(new_n729_), .B(new_n734_), .ZN(new_n3535_));
  AOI21_X1   g3150(.A1(new_n3535_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n3536_));
  OAI21_X1   g3151(.A1(new_n3536_), .A2(new_n407_), .B(new_n745_), .ZN(new_n3537_));
  AOI21_X1   g3152(.A1(new_n3537_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n3538_));
  OAI21_X1   g3153(.A1(new_n3538_), .A2(new_n402_), .B(new_n760_), .ZN(new_n3539_));
  AOI21_X1   g3154(.A1(new_n3539_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n3540_));
  OAI21_X1   g3155(.A1(new_n3540_), .A2(new_n771_), .B(new_n776_), .ZN(new_n3541_));
  AOI21_X1   g3156(.A1(new_n3541_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n3542_));
  OAI21_X1   g3157(.A1(new_n3542_), .A2(new_n389_), .B(new_n787_), .ZN(new_n3543_));
  AOI21_X1   g3158(.A1(new_n3543_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n3544_));
  OAI21_X1   g3159(.A1(new_n3544_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n3545_));
  AOI21_X1   g3160(.A1(new_n3545_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n3546_));
  OAI21_X1   g3161(.A1(new_n3546_), .A2(new_n900_), .B(new_n908_), .ZN(new_n3547_));
  AOI21_X1   g3162(.A1(new_n3547_), .A2(new_n913_), .B(new_n918_), .ZN(new_n3548_));
  OAI21_X1   g3163(.A1(new_n3548_), .A2(new_n897_), .B(new_n923_), .ZN(new_n3549_));
  AOI21_X1   g3164(.A1(new_n3549_), .A2(new_n894_), .B(new_n929_), .ZN(new_n3550_));
  OAI21_X1   g3165(.A1(new_n3550_), .A2(new_n933_), .B(new_n937_), .ZN(new_n3551_));
  AOI21_X1   g3166(.A1(new_n3551_), .A2(new_n890_), .B(new_n943_), .ZN(new_n3552_));
  OAI21_X1   g3167(.A1(new_n3552_), .A2(new_n886_), .B(new_n948_), .ZN(new_n3553_));
  AOI21_X1   g3168(.A1(new_n3553_), .A2(new_n953_), .B(new_n958_), .ZN(new_n3554_));
  OAI21_X1   g3169(.A1(new_n3554_), .A2(new_n883_), .B(new_n963_), .ZN(new_n3555_));
  AOI21_X1   g3170(.A1(new_n3555_), .A2(new_n880_), .B(new_n969_), .ZN(new_n3556_));
  OAI21_X1   g3171(.A1(new_n3556_), .A2(new_n973_), .B(new_n977_), .ZN(new_n3557_));
  AOI21_X1   g3172(.A1(new_n3557_), .A2(new_n876_), .B(new_n983_), .ZN(new_n3558_));
  OAI21_X1   g3173(.A1(new_n3558_), .A2(new_n872_), .B(new_n988_), .ZN(new_n3559_));
  OAI21_X1   g3174(.A1(new_n994_), .A2(\priority[45] ), .B(\req[45] ), .ZN(new_n3560_));
  AOI21_X1   g3175(.A1(new_n3559_), .A2(new_n993_), .B(new_n3560_), .ZN(\grant[45] ));
  NOR2_X1    g3176(.A1(new_n1251_), .A2(new_n1002_), .ZN(new_n3562_));
  OAI21_X1   g3177(.A1(new_n865_), .A2(new_n3562_), .B(new_n1008_), .ZN(new_n3563_));
  AOI21_X1   g3178(.A1(new_n3563_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n3564_));
  OAI21_X1   g3179(.A1(new_n3564_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n3565_));
  AOI21_X1   g3180(.A1(new_n3565_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n3566_));
  OAI21_X1   g3181(.A1(new_n3566_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n3567_));
  AOI21_X1   g3182(.A1(new_n3567_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n3568_));
  OAI21_X1   g3183(.A1(new_n3568_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n3569_));
  AOI21_X1   g3184(.A1(new_n3569_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n3570_));
  OAI21_X1   g3185(.A1(new_n3570_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n3571_));
  AOI21_X1   g3186(.A1(new_n3571_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n3572_));
  OAI21_X1   g3187(.A1(new_n3572_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n3573_));
  AOI21_X1   g3188(.A1(new_n3573_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n3574_));
  OAI21_X1   g3189(.A1(new_n3574_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n3575_));
  AOI21_X1   g3190(.A1(new_n3575_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n3576_));
  OAI21_X1   g3191(.A1(new_n3576_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n3577_));
  AOI21_X1   g3192(.A1(new_n3577_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n3578_));
  OAI21_X1   g3193(.A1(new_n3578_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n3579_));
  AOI21_X1   g3194(.A1(new_n3579_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n3580_));
  OAI21_X1   g3195(.A1(new_n3580_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n3581_));
  AOI21_X1   g3196(.A1(new_n3581_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n3582_));
  OAI21_X1   g3197(.A1(new_n3582_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n3583_));
  AOI21_X1   g3198(.A1(new_n3583_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n3584_));
  OAI21_X1   g3199(.A1(new_n3584_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n3585_));
  AOI21_X1   g3200(.A1(new_n3585_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n3586_));
  OAI21_X1   g3201(.A1(new_n3586_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n3587_));
  AOI21_X1   g3202(.A1(new_n3587_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n3588_));
  OAI21_X1   g3203(.A1(new_n3588_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n3589_));
  AOI21_X1   g3204(.A1(new_n3589_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n3590_));
  OAI21_X1   g3205(.A1(new_n3590_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n3591_));
  AOI21_X1   g3206(.A1(new_n3591_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n3592_));
  OAI21_X1   g3207(.A1(new_n3592_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n3593_));
  AOI21_X1   g3208(.A1(new_n3593_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n3594_));
  OAI21_X1   g3209(.A1(new_n3594_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n3595_));
  AOI21_X1   g3210(.A1(new_n3595_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n3596_));
  OAI21_X1   g3211(.A1(new_n3596_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n3597_));
  AOI21_X1   g3212(.A1(new_n3597_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n3598_));
  OAI21_X1   g3213(.A1(new_n3598_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n3599_));
  AOI21_X1   g3214(.A1(new_n3599_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n3600_));
  OAI21_X1   g3215(.A1(new_n3600_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n3601_));
  AOI21_X1   g3216(.A1(new_n3601_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n3602_));
  OAI21_X1   g3217(.A1(new_n3602_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n3603_));
  OAI21_X1   g3218(.A1(new_n464_), .A2(\priority[46] ), .B(\req[46] ), .ZN(new_n3604_));
  AOI21_X1   g3219(.A1(new_n3603_), .A2(new_n1361_), .B(new_n3604_), .ZN(\grant[46] ));
  NOR2_X1    g3220(.A1(new_n460_), .A2(new_n1368_), .ZN(new_n3606_));
  OAI21_X1   g3221(.A1(new_n1248_), .A2(new_n3606_), .B(new_n1373_), .ZN(new_n3607_));
  AOI21_X1   g3222(.A1(new_n3607_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n3608_));
  OAI21_X1   g3223(.A1(new_n3608_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n3609_));
  AOI21_X1   g3224(.A1(new_n3609_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n3610_));
  OAI21_X1   g3225(.A1(new_n3610_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n3611_));
  AOI21_X1   g3226(.A1(new_n3611_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n3612_));
  OAI21_X1   g3227(.A1(new_n3612_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n3613_));
  AOI21_X1   g3228(.A1(new_n3613_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n3614_));
  OAI21_X1   g3229(.A1(new_n3614_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n3615_));
  AOI21_X1   g3230(.A1(new_n3615_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n3616_));
  OAI21_X1   g3231(.A1(new_n3616_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n3617_));
  AOI21_X1   g3232(.A1(new_n3617_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n3618_));
  OAI21_X1   g3233(.A1(new_n3618_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n3619_));
  AOI21_X1   g3234(.A1(new_n3619_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n3620_));
  OAI21_X1   g3235(.A1(new_n3620_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n3621_));
  AOI21_X1   g3236(.A1(new_n3621_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n3622_));
  OAI21_X1   g3237(.A1(new_n3622_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n3623_));
  AOI21_X1   g3238(.A1(new_n3623_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n3624_));
  OAI21_X1   g3239(.A1(new_n3624_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n3625_));
  AOI21_X1   g3240(.A1(new_n3625_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n3626_));
  OAI21_X1   g3241(.A1(new_n3626_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n3627_));
  AOI21_X1   g3242(.A1(new_n3627_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n3628_));
  OAI21_X1   g3243(.A1(new_n3628_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n3629_));
  AOI21_X1   g3244(.A1(new_n3629_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n3630_));
  OAI21_X1   g3245(.A1(new_n3630_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n3631_));
  AOI21_X1   g3246(.A1(new_n3631_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n3632_));
  OAI21_X1   g3247(.A1(new_n3632_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n3633_));
  AOI21_X1   g3248(.A1(new_n3633_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n3634_));
  OAI21_X1   g3249(.A1(new_n3634_), .A2(new_n519_), .B(new_n524_), .ZN(new_n3635_));
  AOI21_X1   g3250(.A1(new_n3635_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n3636_));
  OAI21_X1   g3251(.A1(new_n3636_), .A2(new_n497_), .B(new_n535_), .ZN(new_n3637_));
  AOI21_X1   g3252(.A1(new_n3637_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n3638_));
  OAI21_X1   g3253(.A1(new_n3638_), .A2(new_n492_), .B(new_n550_), .ZN(new_n3639_));
  AOI21_X1   g3254(.A1(new_n3639_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n3640_));
  OAI21_X1   g3255(.A1(new_n3640_), .A2(new_n561_), .B(new_n566_), .ZN(new_n3641_));
  AOI21_X1   g3256(.A1(new_n3641_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n3642_));
  OAI21_X1   g3257(.A1(new_n3642_), .A2(new_n479_), .B(new_n577_), .ZN(new_n3643_));
  AOI21_X1   g3258(.A1(new_n3643_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n3644_));
  OAI21_X1   g3259(.A1(new_n3644_), .A2(new_n474_), .B(new_n592_), .ZN(new_n3645_));
  AOI21_X1   g3260(.A1(new_n3645_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n3646_));
  OAI21_X1   g3261(.A1(new_n3646_), .A2(new_n603_), .B(new_n608_), .ZN(new_n3647_));
  OAI21_X1   g3262(.A1(new_n611_), .A2(\priority[47] ), .B(\req[47] ), .ZN(new_n3648_));
  AOI21_X1   g3263(.A1(new_n3647_), .A2(new_n1550_), .B(new_n3648_), .ZN(\grant[47] ));
  NOR2_X1    g3264(.A1(new_n864_), .A2(new_n618_), .ZN(new_n3650_));
  OAI21_X1   g3265(.A1(new_n625_), .A2(new_n3650_), .B(new_n629_), .ZN(new_n3651_));
  AOI21_X1   g3266(.A1(new_n3651_), .A2(new_n457_), .B(new_n635_), .ZN(new_n3652_));
  OAI21_X1   g3267(.A1(new_n3652_), .A2(new_n452_), .B(new_n640_), .ZN(new_n3653_));
  AOI21_X1   g3268(.A1(new_n3653_), .A2(new_n646_), .B(new_n651_), .ZN(new_n3654_));
  OAI21_X1   g3269(.A1(new_n3654_), .A2(new_n448_), .B(new_n656_), .ZN(new_n3655_));
  AOI21_X1   g3270(.A1(new_n3655_), .A2(new_n444_), .B(new_n662_), .ZN(new_n3656_));
  OAI21_X1   g3271(.A1(new_n3656_), .A2(new_n667_), .B(new_n671_), .ZN(new_n3657_));
  AOI21_X1   g3272(.A1(new_n3657_), .A2(new_n439_), .B(new_n677_), .ZN(new_n3658_));
  OAI21_X1   g3273(.A1(new_n3658_), .A2(new_n434_), .B(new_n682_), .ZN(new_n3659_));
  AOI21_X1   g3274(.A1(new_n3659_), .A2(new_n688_), .B(new_n693_), .ZN(new_n3660_));
  OAI21_X1   g3275(.A1(new_n3660_), .A2(new_n430_), .B(new_n698_), .ZN(new_n3661_));
  AOI21_X1   g3276(.A1(new_n3661_), .A2(new_n426_), .B(new_n704_), .ZN(new_n3662_));
  OAI21_X1   g3277(.A1(new_n3662_), .A2(new_n709_), .B(new_n713_), .ZN(new_n3663_));
  AOI21_X1   g3278(.A1(new_n3663_), .A2(new_n421_), .B(new_n719_), .ZN(new_n3664_));
  OAI21_X1   g3279(.A1(new_n3664_), .A2(new_n416_), .B(new_n724_), .ZN(new_n3665_));
  AOI21_X1   g3280(.A1(new_n3665_), .A2(new_n730_), .B(new_n735_), .ZN(new_n3666_));
  OAI21_X1   g3281(.A1(new_n3666_), .A2(new_n412_), .B(new_n740_), .ZN(new_n3667_));
  AOI21_X1   g3282(.A1(new_n3667_), .A2(new_n408_), .B(new_n746_), .ZN(new_n3668_));
  OAI21_X1   g3283(.A1(new_n3668_), .A2(new_n751_), .B(new_n755_), .ZN(new_n3669_));
  AOI21_X1   g3284(.A1(new_n3669_), .A2(new_n403_), .B(new_n761_), .ZN(new_n3670_));
  OAI21_X1   g3285(.A1(new_n3670_), .A2(new_n398_), .B(new_n766_), .ZN(new_n3671_));
  AOI21_X1   g3286(.A1(new_n3671_), .A2(new_n772_), .B(new_n777_), .ZN(new_n3672_));
  OAI21_X1   g3287(.A1(new_n3672_), .A2(new_n394_), .B(new_n782_), .ZN(new_n3673_));
  AOI21_X1   g3288(.A1(new_n3673_), .A2(new_n390_), .B(new_n788_), .ZN(new_n3674_));
  OAI21_X1   g3289(.A1(new_n3674_), .A2(new_n793_), .B(new_n797_), .ZN(new_n3675_));
  AOI21_X1   g3290(.A1(new_n3675_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n3676_));
  OAI21_X1   g3291(.A1(new_n3676_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n3677_));
  AOI21_X1   g3292(.A1(new_n3677_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n3678_));
  OAI21_X1   g3293(.A1(new_n3678_), .A2(new_n912_), .B(new_n917_), .ZN(new_n3679_));
  AOI21_X1   g3294(.A1(new_n3679_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n3680_));
  OAI21_X1   g3295(.A1(new_n3680_), .A2(new_n893_), .B(new_n928_), .ZN(new_n3681_));
  AOI21_X1   g3296(.A1(new_n3681_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n3682_));
  OAI21_X1   g3297(.A1(new_n3682_), .A2(new_n889_), .B(new_n942_), .ZN(new_n3683_));
  AOI21_X1   g3298(.A1(new_n3683_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n3684_));
  OAI21_X1   g3299(.A1(new_n3684_), .A2(new_n952_), .B(new_n957_), .ZN(new_n3685_));
  AOI21_X1   g3300(.A1(new_n3685_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n3686_));
  OAI21_X1   g3301(.A1(new_n3686_), .A2(new_n879_), .B(new_n968_), .ZN(new_n3687_));
  AOI21_X1   g3302(.A1(new_n3687_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n3688_));
  OAI21_X1   g3303(.A1(new_n3688_), .A2(new_n875_), .B(new_n982_), .ZN(new_n3689_));
  AOI21_X1   g3304(.A1(new_n3689_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n3690_));
  OAI21_X1   g3305(.A1(new_n3690_), .A2(new_n992_), .B(new_n997_), .ZN(new_n3691_));
  OAI21_X1   g3306(.A1(new_n1000_), .A2(\priority[48] ), .B(\req[48] ), .ZN(new_n3692_));
  AOI21_X1   g3307(.A1(new_n3691_), .A2(new_n1640_), .B(new_n3692_), .ZN(\grant[48] ));
  NOR2_X1    g3308(.A1(new_n1247_), .A2(new_n1007_), .ZN(new_n3694_));
  OAI21_X1   g3309(.A1(new_n1013_), .A2(new_n3694_), .B(new_n1017_), .ZN(new_n3695_));
  AOI21_X1   g3310(.A1(new_n3695_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n3696_));
  OAI21_X1   g3311(.A1(new_n3696_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n3697_));
  AOI21_X1   g3312(.A1(new_n3697_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n3698_));
  OAI21_X1   g3313(.A1(new_n3698_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n3699_));
  AOI21_X1   g3314(.A1(new_n3699_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n3700_));
  OAI21_X1   g3315(.A1(new_n3700_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n3701_));
  AOI21_X1   g3316(.A1(new_n3701_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n3702_));
  OAI21_X1   g3317(.A1(new_n3702_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n3703_));
  AOI21_X1   g3318(.A1(new_n3703_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n3704_));
  OAI21_X1   g3319(.A1(new_n3704_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n3705_));
  AOI21_X1   g3320(.A1(new_n3705_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n3706_));
  OAI21_X1   g3321(.A1(new_n3706_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n3707_));
  AOI21_X1   g3322(.A1(new_n3707_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n3708_));
  OAI21_X1   g3323(.A1(new_n3708_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n3709_));
  AOI21_X1   g3324(.A1(new_n3709_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n3710_));
  OAI21_X1   g3325(.A1(new_n3710_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n3711_));
  AOI21_X1   g3326(.A1(new_n3711_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n3712_));
  OAI21_X1   g3327(.A1(new_n3712_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n3713_));
  AOI21_X1   g3328(.A1(new_n3713_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n3714_));
  OAI21_X1   g3329(.A1(new_n3714_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n3715_));
  AOI21_X1   g3330(.A1(new_n3715_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n3716_));
  OAI21_X1   g3331(.A1(new_n3716_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n3717_));
  AOI21_X1   g3332(.A1(new_n3717_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n3718_));
  OAI21_X1   g3333(.A1(new_n3718_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n3719_));
  AOI21_X1   g3334(.A1(new_n3719_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n3720_));
  OAI21_X1   g3335(.A1(new_n3720_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n3721_));
  AOI21_X1   g3336(.A1(new_n3721_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n3722_));
  OAI21_X1   g3337(.A1(new_n3722_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n3723_));
  AOI21_X1   g3338(.A1(new_n3723_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n3724_));
  OAI21_X1   g3339(.A1(new_n3724_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n3725_));
  AOI21_X1   g3340(.A1(new_n3725_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n3726_));
  OAI21_X1   g3341(.A1(new_n3726_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n3727_));
  AOI21_X1   g3342(.A1(new_n3727_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n3728_));
  OAI21_X1   g3343(.A1(new_n3728_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n3729_));
  AOI21_X1   g3344(.A1(new_n3729_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n3730_));
  OAI21_X1   g3345(.A1(new_n3730_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n3731_));
  AOI21_X1   g3346(.A1(new_n3731_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n3732_));
  OAI21_X1   g3347(.A1(new_n3732_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n3733_));
  AOI21_X1   g3348(.A1(new_n3733_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n3734_));
  OAI21_X1   g3349(.A1(new_n3734_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n3735_));
  OAI21_X1   g3350(.A1(new_n459_), .A2(\priority[49] ), .B(\req[49] ), .ZN(new_n3736_));
  AOI21_X1   g3351(.A1(new_n3735_), .A2(new_n1728_), .B(new_n3736_), .ZN(\grant[49] ));
  NOR2_X1    g3352(.A1(new_n624_), .A2(new_n1372_), .ZN(new_n3738_));
  OAI21_X1   g3353(.A1(new_n1378_), .A2(new_n3738_), .B(new_n1381_), .ZN(new_n3739_));
  AOI21_X1   g3354(.A1(new_n3739_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n3740_));
  OAI21_X1   g3355(.A1(new_n3740_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n3741_));
  AOI21_X1   g3356(.A1(new_n3741_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n3742_));
  OAI21_X1   g3357(.A1(new_n3742_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n3743_));
  AOI21_X1   g3358(.A1(new_n3743_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n3744_));
  OAI21_X1   g3359(.A1(new_n3744_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n3745_));
  AOI21_X1   g3360(.A1(new_n3745_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n3746_));
  OAI21_X1   g3361(.A1(new_n3746_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n3747_));
  AOI21_X1   g3362(.A1(new_n3747_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n3748_));
  OAI21_X1   g3363(.A1(new_n3748_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n3749_));
  AOI21_X1   g3364(.A1(new_n3749_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n3750_));
  OAI21_X1   g3365(.A1(new_n3750_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n3751_));
  AOI21_X1   g3366(.A1(new_n3751_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n3752_));
  OAI21_X1   g3367(.A1(new_n3752_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n3753_));
  AOI21_X1   g3368(.A1(new_n3753_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n3754_));
  OAI21_X1   g3369(.A1(new_n3754_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n3755_));
  AOI21_X1   g3370(.A1(new_n3755_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n3756_));
  OAI21_X1   g3371(.A1(new_n3756_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n3757_));
  AOI21_X1   g3372(.A1(new_n3757_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n3758_));
  OAI21_X1   g3373(.A1(new_n3758_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n3759_));
  AOI21_X1   g3374(.A1(new_n3759_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n3760_));
  OAI21_X1   g3375(.A1(new_n3760_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n3761_));
  AOI21_X1   g3376(.A1(new_n3761_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n3762_));
  OAI21_X1   g3377(.A1(new_n3762_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n3763_));
  AOI21_X1   g3378(.A1(new_n3763_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n3764_));
  OAI21_X1   g3379(.A1(new_n3764_), .A2(new_n506_), .B(new_n514_), .ZN(new_n3765_));
  AOI21_X1   g3380(.A1(new_n3765_), .A2(new_n520_), .B(new_n525_), .ZN(new_n3766_));
  OAI21_X1   g3381(.A1(new_n3766_), .A2(new_n502_), .B(new_n530_), .ZN(new_n3767_));
  AOI21_X1   g3382(.A1(new_n3767_), .A2(new_n498_), .B(new_n536_), .ZN(new_n3768_));
  OAI21_X1   g3383(.A1(new_n3768_), .A2(new_n541_), .B(new_n545_), .ZN(new_n3769_));
  AOI21_X1   g3384(.A1(new_n3769_), .A2(new_n493_), .B(new_n551_), .ZN(new_n3770_));
  OAI21_X1   g3385(.A1(new_n3770_), .A2(new_n488_), .B(new_n556_), .ZN(new_n3771_));
  AOI21_X1   g3386(.A1(new_n3771_), .A2(new_n562_), .B(new_n567_), .ZN(new_n3772_));
  OAI21_X1   g3387(.A1(new_n3772_), .A2(new_n484_), .B(new_n572_), .ZN(new_n3773_));
  AOI21_X1   g3388(.A1(new_n3773_), .A2(new_n480_), .B(new_n578_), .ZN(new_n3774_));
  OAI21_X1   g3389(.A1(new_n3774_), .A2(new_n583_), .B(new_n587_), .ZN(new_n3775_));
  AOI21_X1   g3390(.A1(new_n3775_), .A2(new_n475_), .B(new_n593_), .ZN(new_n3776_));
  OAI21_X1   g3391(.A1(new_n3776_), .A2(new_n470_), .B(new_n598_), .ZN(new_n3777_));
  AOI21_X1   g3392(.A1(new_n3777_), .A2(new_n604_), .B(new_n609_), .ZN(new_n3778_));
  OAI21_X1   g3393(.A1(new_n3778_), .A2(new_n466_), .B(new_n614_), .ZN(new_n3779_));
  OAI21_X1   g3394(.A1(new_n616_), .A2(\priority[50] ), .B(\req[50] ), .ZN(new_n3780_));
  AOI21_X1   g3395(.A1(new_n3779_), .A2(new_n462_), .B(new_n3780_), .ZN(\grant[50] ));
  NOR2_X1    g3396(.A1(new_n1012_), .A2(new_n628_), .ZN(new_n3782_));
  OAI21_X1   g3397(.A1(new_n456_), .A2(new_n3782_), .B(new_n634_), .ZN(new_n3783_));
  AOI21_X1   g3398(.A1(new_n3783_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n3784_));
  OAI21_X1   g3399(.A1(new_n3784_), .A2(new_n645_), .B(new_n650_), .ZN(new_n3785_));
  AOI21_X1   g3400(.A1(new_n3785_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n3786_));
  OAI21_X1   g3401(.A1(new_n3786_), .A2(new_n443_), .B(new_n661_), .ZN(new_n3787_));
  AOI21_X1   g3402(.A1(new_n3787_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n3788_));
  OAI21_X1   g3403(.A1(new_n3788_), .A2(new_n438_), .B(new_n676_), .ZN(new_n3789_));
  AOI21_X1   g3404(.A1(new_n3789_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n3790_));
  OAI21_X1   g3405(.A1(new_n3790_), .A2(new_n687_), .B(new_n692_), .ZN(new_n3791_));
  AOI21_X1   g3406(.A1(new_n3791_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n3792_));
  OAI21_X1   g3407(.A1(new_n3792_), .A2(new_n425_), .B(new_n703_), .ZN(new_n3793_));
  AOI21_X1   g3408(.A1(new_n3793_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n3794_));
  OAI21_X1   g3409(.A1(new_n3794_), .A2(new_n420_), .B(new_n718_), .ZN(new_n3795_));
  AOI21_X1   g3410(.A1(new_n3795_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n3796_));
  OAI21_X1   g3411(.A1(new_n3796_), .A2(new_n729_), .B(new_n734_), .ZN(new_n3797_));
  AOI21_X1   g3412(.A1(new_n3797_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n3798_));
  OAI21_X1   g3413(.A1(new_n3798_), .A2(new_n407_), .B(new_n745_), .ZN(new_n3799_));
  AOI21_X1   g3414(.A1(new_n3799_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n3800_));
  OAI21_X1   g3415(.A1(new_n3800_), .A2(new_n402_), .B(new_n760_), .ZN(new_n3801_));
  AOI21_X1   g3416(.A1(new_n3801_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n3802_));
  OAI21_X1   g3417(.A1(new_n3802_), .A2(new_n771_), .B(new_n776_), .ZN(new_n3803_));
  AOI21_X1   g3418(.A1(new_n3803_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n3804_));
  OAI21_X1   g3419(.A1(new_n3804_), .A2(new_n389_), .B(new_n787_), .ZN(new_n3805_));
  AOI21_X1   g3420(.A1(new_n3805_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n3806_));
  OAI21_X1   g3421(.A1(new_n3806_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n3807_));
  AOI21_X1   g3422(.A1(new_n3807_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n3808_));
  OAI21_X1   g3423(.A1(new_n3808_), .A2(new_n900_), .B(new_n908_), .ZN(new_n3809_));
  AOI21_X1   g3424(.A1(new_n3809_), .A2(new_n913_), .B(new_n918_), .ZN(new_n3810_));
  OAI21_X1   g3425(.A1(new_n3810_), .A2(new_n897_), .B(new_n923_), .ZN(new_n3811_));
  AOI21_X1   g3426(.A1(new_n3811_), .A2(new_n894_), .B(new_n929_), .ZN(new_n3812_));
  OAI21_X1   g3427(.A1(new_n3812_), .A2(new_n933_), .B(new_n937_), .ZN(new_n3813_));
  AOI21_X1   g3428(.A1(new_n3813_), .A2(new_n890_), .B(new_n943_), .ZN(new_n3814_));
  OAI21_X1   g3429(.A1(new_n3814_), .A2(new_n886_), .B(new_n948_), .ZN(new_n3815_));
  AOI21_X1   g3430(.A1(new_n3815_), .A2(new_n953_), .B(new_n958_), .ZN(new_n3816_));
  OAI21_X1   g3431(.A1(new_n3816_), .A2(new_n883_), .B(new_n963_), .ZN(new_n3817_));
  AOI21_X1   g3432(.A1(new_n3817_), .A2(new_n880_), .B(new_n969_), .ZN(new_n3818_));
  OAI21_X1   g3433(.A1(new_n3818_), .A2(new_n973_), .B(new_n977_), .ZN(new_n3819_));
  AOI21_X1   g3434(.A1(new_n3819_), .A2(new_n876_), .B(new_n983_), .ZN(new_n3820_));
  OAI21_X1   g3435(.A1(new_n3820_), .A2(new_n872_), .B(new_n988_), .ZN(new_n3821_));
  AOI21_X1   g3436(.A1(new_n3821_), .A2(new_n993_), .B(new_n998_), .ZN(new_n3822_));
  OAI21_X1   g3437(.A1(new_n3822_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n3823_));
  OAI21_X1   g3438(.A1(new_n1005_), .A2(\priority[51] ), .B(\req[51] ), .ZN(new_n3824_));
  AOI21_X1   g3439(.A1(new_n3823_), .A2(new_n866_), .B(new_n3824_), .ZN(\grant[51] ));
  NOR2_X1    g3440(.A1(new_n1377_), .A2(new_n1016_), .ZN(new_n3826_));
  OAI21_X1   g3441(.A1(new_n861_), .A2(new_n3826_), .B(new_n1022_), .ZN(new_n3827_));
  AOI21_X1   g3442(.A1(new_n3827_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n3828_));
  OAI21_X1   g3443(.A1(new_n3828_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n3829_));
  AOI21_X1   g3444(.A1(new_n3829_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n3830_));
  OAI21_X1   g3445(.A1(new_n3830_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n3831_));
  AOI21_X1   g3446(.A1(new_n3831_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n3832_));
  OAI21_X1   g3447(.A1(new_n3832_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n3833_));
  AOI21_X1   g3448(.A1(new_n3833_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n3834_));
  OAI21_X1   g3449(.A1(new_n3834_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n3835_));
  AOI21_X1   g3450(.A1(new_n3835_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n3836_));
  OAI21_X1   g3451(.A1(new_n3836_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n3837_));
  AOI21_X1   g3452(.A1(new_n3837_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n3838_));
  OAI21_X1   g3453(.A1(new_n3838_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n3839_));
  AOI21_X1   g3454(.A1(new_n3839_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n3840_));
  OAI21_X1   g3455(.A1(new_n3840_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n3841_));
  AOI21_X1   g3456(.A1(new_n3841_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n3842_));
  OAI21_X1   g3457(.A1(new_n3842_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n3843_));
  AOI21_X1   g3458(.A1(new_n3843_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n3844_));
  OAI21_X1   g3459(.A1(new_n3844_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n3845_));
  AOI21_X1   g3460(.A1(new_n3845_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n3846_));
  OAI21_X1   g3461(.A1(new_n3846_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n3847_));
  AOI21_X1   g3462(.A1(new_n3847_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n3848_));
  OAI21_X1   g3463(.A1(new_n3848_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n3849_));
  AOI21_X1   g3464(.A1(new_n3849_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n3850_));
  OAI21_X1   g3465(.A1(new_n3850_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n3851_));
  AOI21_X1   g3466(.A1(new_n3851_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n3852_));
  OAI21_X1   g3467(.A1(new_n3852_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n3853_));
  AOI21_X1   g3468(.A1(new_n3853_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n3854_));
  OAI21_X1   g3469(.A1(new_n3854_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n3855_));
  AOI21_X1   g3470(.A1(new_n3855_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n3856_));
  OAI21_X1   g3471(.A1(new_n3856_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n3857_));
  AOI21_X1   g3472(.A1(new_n3857_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n3858_));
  OAI21_X1   g3473(.A1(new_n3858_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n3859_));
  AOI21_X1   g3474(.A1(new_n3859_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n3860_));
  OAI21_X1   g3475(.A1(new_n3860_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n3861_));
  AOI21_X1   g3476(.A1(new_n3861_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n3862_));
  OAI21_X1   g3477(.A1(new_n3862_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n3863_));
  AOI21_X1   g3478(.A1(new_n3863_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n3864_));
  OAI21_X1   g3479(.A1(new_n3864_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n3865_));
  AOI21_X1   g3480(.A1(new_n3865_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n3866_));
  OAI21_X1   g3481(.A1(new_n3866_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n3867_));
  OAI21_X1   g3482(.A1(new_n623_), .A2(\priority[52] ), .B(\req[52] ), .ZN(new_n3868_));
  AOI21_X1   g3483(.A1(new_n3867_), .A2(new_n1249_), .B(new_n3868_), .ZN(\grant[52] ));
  NOR2_X1    g3484(.A1(new_n455_), .A2(new_n1380_), .ZN(new_n3870_));
  OAI21_X1   g3485(.A1(new_n1244_), .A2(new_n3870_), .B(new_n1385_), .ZN(new_n3871_));
  AOI21_X1   g3486(.A1(new_n3871_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n3872_));
  OAI21_X1   g3487(.A1(new_n3872_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n3873_));
  AOI21_X1   g3488(.A1(new_n3873_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n3874_));
  OAI21_X1   g3489(.A1(new_n3874_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n3875_));
  AOI21_X1   g3490(.A1(new_n3875_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n3876_));
  OAI21_X1   g3491(.A1(new_n3876_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n3877_));
  AOI21_X1   g3492(.A1(new_n3877_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n3878_));
  OAI21_X1   g3493(.A1(new_n3878_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n3879_));
  AOI21_X1   g3494(.A1(new_n3879_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n3880_));
  OAI21_X1   g3495(.A1(new_n3880_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n3881_));
  AOI21_X1   g3496(.A1(new_n3881_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n3882_));
  OAI21_X1   g3497(.A1(new_n3882_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n3883_));
  AOI21_X1   g3498(.A1(new_n3883_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n3884_));
  OAI21_X1   g3499(.A1(new_n3884_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n3885_));
  AOI21_X1   g3500(.A1(new_n3885_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n3886_));
  OAI21_X1   g3501(.A1(new_n3886_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n3887_));
  AOI21_X1   g3502(.A1(new_n3887_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n3888_));
  OAI21_X1   g3503(.A1(new_n3888_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n3889_));
  AOI21_X1   g3504(.A1(new_n3889_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n3890_));
  OAI21_X1   g3505(.A1(new_n3890_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n3891_));
  AOI21_X1   g3506(.A1(new_n3891_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n3892_));
  OAI21_X1   g3507(.A1(new_n3892_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n3893_));
  AOI21_X1   g3508(.A1(new_n3893_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n3894_));
  OAI21_X1   g3509(.A1(new_n3894_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n3895_));
  AOI21_X1   g3510(.A1(new_n3895_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n3896_));
  OAI21_X1   g3511(.A1(new_n3896_), .A2(new_n519_), .B(new_n524_), .ZN(new_n3897_));
  AOI21_X1   g3512(.A1(new_n3897_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n3898_));
  OAI21_X1   g3513(.A1(new_n3898_), .A2(new_n497_), .B(new_n535_), .ZN(new_n3899_));
  AOI21_X1   g3514(.A1(new_n3899_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n3900_));
  OAI21_X1   g3515(.A1(new_n3900_), .A2(new_n492_), .B(new_n550_), .ZN(new_n3901_));
  AOI21_X1   g3516(.A1(new_n3901_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n3902_));
  OAI21_X1   g3517(.A1(new_n3902_), .A2(new_n561_), .B(new_n566_), .ZN(new_n3903_));
  AOI21_X1   g3518(.A1(new_n3903_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n3904_));
  OAI21_X1   g3519(.A1(new_n3904_), .A2(new_n479_), .B(new_n577_), .ZN(new_n3905_));
  AOI21_X1   g3520(.A1(new_n3905_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n3906_));
  OAI21_X1   g3521(.A1(new_n3906_), .A2(new_n474_), .B(new_n592_), .ZN(new_n3907_));
  AOI21_X1   g3522(.A1(new_n3907_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n3908_));
  OAI21_X1   g3523(.A1(new_n3908_), .A2(new_n603_), .B(new_n608_), .ZN(new_n3909_));
  AOI21_X1   g3524(.A1(new_n3909_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n3910_));
  OAI21_X1   g3525(.A1(new_n3910_), .A2(new_n461_), .B(new_n619_), .ZN(new_n3911_));
  OAI21_X1   g3526(.A1(new_n626_), .A2(\priority[53] ), .B(\req[53] ), .ZN(new_n3912_));
  AOI21_X1   g3527(.A1(new_n3911_), .A2(new_n1548_), .B(new_n3912_), .ZN(\grant[53] ));
  NOR2_X1    g3528(.A1(new_n860_), .A2(new_n633_), .ZN(new_n3914_));
  OAI21_X1   g3529(.A1(new_n452_), .A2(new_n3914_), .B(new_n640_), .ZN(new_n3915_));
  AOI21_X1   g3530(.A1(new_n3915_), .A2(new_n646_), .B(new_n651_), .ZN(new_n3916_));
  OAI21_X1   g3531(.A1(new_n3916_), .A2(new_n448_), .B(new_n656_), .ZN(new_n3917_));
  AOI21_X1   g3532(.A1(new_n3917_), .A2(new_n444_), .B(new_n662_), .ZN(new_n3918_));
  OAI21_X1   g3533(.A1(new_n3918_), .A2(new_n667_), .B(new_n671_), .ZN(new_n3919_));
  AOI21_X1   g3534(.A1(new_n3919_), .A2(new_n439_), .B(new_n677_), .ZN(new_n3920_));
  OAI21_X1   g3535(.A1(new_n3920_), .A2(new_n434_), .B(new_n682_), .ZN(new_n3921_));
  AOI21_X1   g3536(.A1(new_n3921_), .A2(new_n688_), .B(new_n693_), .ZN(new_n3922_));
  OAI21_X1   g3537(.A1(new_n3922_), .A2(new_n430_), .B(new_n698_), .ZN(new_n3923_));
  AOI21_X1   g3538(.A1(new_n3923_), .A2(new_n426_), .B(new_n704_), .ZN(new_n3924_));
  OAI21_X1   g3539(.A1(new_n3924_), .A2(new_n709_), .B(new_n713_), .ZN(new_n3925_));
  AOI21_X1   g3540(.A1(new_n3925_), .A2(new_n421_), .B(new_n719_), .ZN(new_n3926_));
  OAI21_X1   g3541(.A1(new_n3926_), .A2(new_n416_), .B(new_n724_), .ZN(new_n3927_));
  AOI21_X1   g3542(.A1(new_n3927_), .A2(new_n730_), .B(new_n735_), .ZN(new_n3928_));
  OAI21_X1   g3543(.A1(new_n3928_), .A2(new_n412_), .B(new_n740_), .ZN(new_n3929_));
  AOI21_X1   g3544(.A1(new_n3929_), .A2(new_n408_), .B(new_n746_), .ZN(new_n3930_));
  OAI21_X1   g3545(.A1(new_n3930_), .A2(new_n751_), .B(new_n755_), .ZN(new_n3931_));
  AOI21_X1   g3546(.A1(new_n3931_), .A2(new_n403_), .B(new_n761_), .ZN(new_n3932_));
  OAI21_X1   g3547(.A1(new_n3932_), .A2(new_n398_), .B(new_n766_), .ZN(new_n3933_));
  AOI21_X1   g3548(.A1(new_n3933_), .A2(new_n772_), .B(new_n777_), .ZN(new_n3934_));
  OAI21_X1   g3549(.A1(new_n3934_), .A2(new_n394_), .B(new_n782_), .ZN(new_n3935_));
  AOI21_X1   g3550(.A1(new_n3935_), .A2(new_n390_), .B(new_n788_), .ZN(new_n3936_));
  OAI21_X1   g3551(.A1(new_n3936_), .A2(new_n793_), .B(new_n797_), .ZN(new_n3937_));
  AOI21_X1   g3552(.A1(new_n3937_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n3938_));
  OAI21_X1   g3553(.A1(new_n3938_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n3939_));
  AOI21_X1   g3554(.A1(new_n3939_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n3940_));
  OAI21_X1   g3555(.A1(new_n3940_), .A2(new_n912_), .B(new_n917_), .ZN(new_n3941_));
  AOI21_X1   g3556(.A1(new_n3941_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n3942_));
  OAI21_X1   g3557(.A1(new_n3942_), .A2(new_n893_), .B(new_n928_), .ZN(new_n3943_));
  AOI21_X1   g3558(.A1(new_n3943_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n3944_));
  OAI21_X1   g3559(.A1(new_n3944_), .A2(new_n889_), .B(new_n942_), .ZN(new_n3945_));
  AOI21_X1   g3560(.A1(new_n3945_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n3946_));
  OAI21_X1   g3561(.A1(new_n3946_), .A2(new_n952_), .B(new_n957_), .ZN(new_n3947_));
  AOI21_X1   g3562(.A1(new_n3947_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n3948_));
  OAI21_X1   g3563(.A1(new_n3948_), .A2(new_n879_), .B(new_n968_), .ZN(new_n3949_));
  AOI21_X1   g3564(.A1(new_n3949_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n3950_));
  OAI21_X1   g3565(.A1(new_n3950_), .A2(new_n875_), .B(new_n982_), .ZN(new_n3951_));
  AOI21_X1   g3566(.A1(new_n3951_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n3952_));
  OAI21_X1   g3567(.A1(new_n3952_), .A2(new_n992_), .B(new_n997_), .ZN(new_n3953_));
  AOI21_X1   g3568(.A1(new_n3953_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n3954_));
  OAI21_X1   g3569(.A1(new_n3954_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n3955_));
  OAI21_X1   g3570(.A1(new_n1014_), .A2(\priority[54] ), .B(\req[54] ), .ZN(new_n3956_));
  AOI21_X1   g3571(.A1(new_n3955_), .A2(new_n1638_), .B(new_n3956_), .ZN(\grant[54] ));
  NOR2_X1    g3572(.A1(new_n1243_), .A2(new_n1021_), .ZN(new_n3958_));
  OAI21_X1   g3573(.A1(new_n858_), .A2(new_n3958_), .B(new_n1028_), .ZN(new_n3959_));
  AOI21_X1   g3574(.A1(new_n3959_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n3960_));
  OAI21_X1   g3575(.A1(new_n3960_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n3961_));
  AOI21_X1   g3576(.A1(new_n3961_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n3962_));
  OAI21_X1   g3577(.A1(new_n3962_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n3963_));
  AOI21_X1   g3578(.A1(new_n3963_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n3964_));
  OAI21_X1   g3579(.A1(new_n3964_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n3965_));
  AOI21_X1   g3580(.A1(new_n3965_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n3966_));
  OAI21_X1   g3581(.A1(new_n3966_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n3967_));
  AOI21_X1   g3582(.A1(new_n3967_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n3968_));
  OAI21_X1   g3583(.A1(new_n3968_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n3969_));
  AOI21_X1   g3584(.A1(new_n3969_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n3970_));
  OAI21_X1   g3585(.A1(new_n3970_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n3971_));
  AOI21_X1   g3586(.A1(new_n3971_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n3972_));
  OAI21_X1   g3587(.A1(new_n3972_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n3973_));
  AOI21_X1   g3588(.A1(new_n3973_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n3974_));
  OAI21_X1   g3589(.A1(new_n3974_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n3975_));
  AOI21_X1   g3590(.A1(new_n3975_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n3976_));
  OAI21_X1   g3591(.A1(new_n3976_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n3977_));
  AOI21_X1   g3592(.A1(new_n3977_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n3978_));
  OAI21_X1   g3593(.A1(new_n3978_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n3979_));
  AOI21_X1   g3594(.A1(new_n3979_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n3980_));
  OAI21_X1   g3595(.A1(new_n3980_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n3981_));
  AOI21_X1   g3596(.A1(new_n3981_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n3982_));
  OAI21_X1   g3597(.A1(new_n3982_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n3983_));
  AOI21_X1   g3598(.A1(new_n3983_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n3984_));
  OAI21_X1   g3599(.A1(new_n3984_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n3985_));
  AOI21_X1   g3600(.A1(new_n3985_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n3986_));
  OAI21_X1   g3601(.A1(new_n3986_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n3987_));
  AOI21_X1   g3602(.A1(new_n3987_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n3988_));
  OAI21_X1   g3603(.A1(new_n3988_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n3989_));
  AOI21_X1   g3604(.A1(new_n3989_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n3990_));
  OAI21_X1   g3605(.A1(new_n3990_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n3991_));
  AOI21_X1   g3606(.A1(new_n3991_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n3992_));
  OAI21_X1   g3607(.A1(new_n3992_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n3993_));
  AOI21_X1   g3608(.A1(new_n3993_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n3994_));
  OAI21_X1   g3609(.A1(new_n3994_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n3995_));
  AOI21_X1   g3610(.A1(new_n3995_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n3996_));
  OAI21_X1   g3611(.A1(new_n3996_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n3997_));
  AOI21_X1   g3612(.A1(new_n3997_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n3998_));
  OAI21_X1   g3613(.A1(new_n3998_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n3999_));
  OAI21_X1   g3614(.A1(new_n454_), .A2(\priority[55] ), .B(\req[55] ), .ZN(new_n4000_));
  AOI21_X1   g3615(.A1(new_n3999_), .A2(new_n1726_), .B(new_n4000_), .ZN(\grant[55] ));
  NOR2_X1    g3616(.A1(new_n451_), .A2(new_n1384_), .ZN(new_n4002_));
  OAI21_X1   g3617(.A1(new_n1241_), .A2(new_n4002_), .B(new_n1390_), .ZN(new_n4003_));
  AOI21_X1   g3618(.A1(new_n4003_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n4004_));
  OAI21_X1   g3619(.A1(new_n4004_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n4005_));
  AOI21_X1   g3620(.A1(new_n4005_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n4006_));
  OAI21_X1   g3621(.A1(new_n4006_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n4007_));
  AOI21_X1   g3622(.A1(new_n4007_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n4008_));
  OAI21_X1   g3623(.A1(new_n4008_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n4009_));
  AOI21_X1   g3624(.A1(new_n4009_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n4010_));
  OAI21_X1   g3625(.A1(new_n4010_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n4011_));
  AOI21_X1   g3626(.A1(new_n4011_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n4012_));
  OAI21_X1   g3627(.A1(new_n4012_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n4013_));
  AOI21_X1   g3628(.A1(new_n4013_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n4014_));
  OAI21_X1   g3629(.A1(new_n4014_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n4015_));
  AOI21_X1   g3630(.A1(new_n4015_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n4016_));
  OAI21_X1   g3631(.A1(new_n4016_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n4017_));
  AOI21_X1   g3632(.A1(new_n4017_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n4018_));
  OAI21_X1   g3633(.A1(new_n4018_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n4019_));
  AOI21_X1   g3634(.A1(new_n4019_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n4020_));
  OAI21_X1   g3635(.A1(new_n4020_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n4021_));
  AOI21_X1   g3636(.A1(new_n4021_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n4022_));
  OAI21_X1   g3637(.A1(new_n4022_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n4023_));
  AOI21_X1   g3638(.A1(new_n4023_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n4024_));
  OAI21_X1   g3639(.A1(new_n4024_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n4025_));
  AOI21_X1   g3640(.A1(new_n4025_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n4026_));
  OAI21_X1   g3641(.A1(new_n4026_), .A2(new_n506_), .B(new_n514_), .ZN(new_n4027_));
  AOI21_X1   g3642(.A1(new_n4027_), .A2(new_n520_), .B(new_n525_), .ZN(new_n4028_));
  OAI21_X1   g3643(.A1(new_n4028_), .A2(new_n502_), .B(new_n530_), .ZN(new_n4029_));
  AOI21_X1   g3644(.A1(new_n4029_), .A2(new_n498_), .B(new_n536_), .ZN(new_n4030_));
  OAI21_X1   g3645(.A1(new_n4030_), .A2(new_n541_), .B(new_n545_), .ZN(new_n4031_));
  AOI21_X1   g3646(.A1(new_n4031_), .A2(new_n493_), .B(new_n551_), .ZN(new_n4032_));
  OAI21_X1   g3647(.A1(new_n4032_), .A2(new_n488_), .B(new_n556_), .ZN(new_n4033_));
  AOI21_X1   g3648(.A1(new_n4033_), .A2(new_n562_), .B(new_n567_), .ZN(new_n4034_));
  OAI21_X1   g3649(.A1(new_n4034_), .A2(new_n484_), .B(new_n572_), .ZN(new_n4035_));
  AOI21_X1   g3650(.A1(new_n4035_), .A2(new_n480_), .B(new_n578_), .ZN(new_n4036_));
  OAI21_X1   g3651(.A1(new_n4036_), .A2(new_n583_), .B(new_n587_), .ZN(new_n4037_));
  AOI21_X1   g3652(.A1(new_n4037_), .A2(new_n475_), .B(new_n593_), .ZN(new_n4038_));
  OAI21_X1   g3653(.A1(new_n4038_), .A2(new_n470_), .B(new_n598_), .ZN(new_n4039_));
  AOI21_X1   g3654(.A1(new_n4039_), .A2(new_n604_), .B(new_n609_), .ZN(new_n4040_));
  OAI21_X1   g3655(.A1(new_n4040_), .A2(new_n466_), .B(new_n614_), .ZN(new_n4041_));
  AOI21_X1   g3656(.A1(new_n4041_), .A2(new_n462_), .B(new_n620_), .ZN(new_n4042_));
  OAI21_X1   g3657(.A1(new_n4042_), .A2(new_n625_), .B(new_n629_), .ZN(new_n4043_));
  OAI21_X1   g3658(.A1(new_n631_), .A2(\priority[56] ), .B(\req[56] ), .ZN(new_n4044_));
  AOI21_X1   g3659(.A1(new_n4043_), .A2(new_n457_), .B(new_n4044_), .ZN(\grant[56] ));
  NOR2_X1    g3660(.A1(new_n857_), .A2(new_n639_), .ZN(new_n4046_));
  OAI21_X1   g3661(.A1(new_n645_), .A2(new_n4046_), .B(new_n650_), .ZN(new_n4047_));
  AOI21_X1   g3662(.A1(new_n4047_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n4048_));
  OAI21_X1   g3663(.A1(new_n4048_), .A2(new_n443_), .B(new_n661_), .ZN(new_n4049_));
  AOI21_X1   g3664(.A1(new_n4049_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n4050_));
  OAI21_X1   g3665(.A1(new_n4050_), .A2(new_n438_), .B(new_n676_), .ZN(new_n4051_));
  AOI21_X1   g3666(.A1(new_n4051_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n4052_));
  OAI21_X1   g3667(.A1(new_n4052_), .A2(new_n687_), .B(new_n692_), .ZN(new_n4053_));
  AOI21_X1   g3668(.A1(new_n4053_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n4054_));
  OAI21_X1   g3669(.A1(new_n4054_), .A2(new_n425_), .B(new_n703_), .ZN(new_n4055_));
  AOI21_X1   g3670(.A1(new_n4055_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n4056_));
  OAI21_X1   g3671(.A1(new_n4056_), .A2(new_n420_), .B(new_n718_), .ZN(new_n4057_));
  AOI21_X1   g3672(.A1(new_n4057_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n4058_));
  OAI21_X1   g3673(.A1(new_n4058_), .A2(new_n729_), .B(new_n734_), .ZN(new_n4059_));
  AOI21_X1   g3674(.A1(new_n4059_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n4060_));
  OAI21_X1   g3675(.A1(new_n4060_), .A2(new_n407_), .B(new_n745_), .ZN(new_n4061_));
  AOI21_X1   g3676(.A1(new_n4061_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n4062_));
  OAI21_X1   g3677(.A1(new_n4062_), .A2(new_n402_), .B(new_n760_), .ZN(new_n4063_));
  AOI21_X1   g3678(.A1(new_n4063_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n4064_));
  OAI21_X1   g3679(.A1(new_n4064_), .A2(new_n771_), .B(new_n776_), .ZN(new_n4065_));
  AOI21_X1   g3680(.A1(new_n4065_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n4066_));
  OAI21_X1   g3681(.A1(new_n4066_), .A2(new_n389_), .B(new_n787_), .ZN(new_n4067_));
  AOI21_X1   g3682(.A1(new_n4067_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n4068_));
  OAI21_X1   g3683(.A1(new_n4068_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n4069_));
  AOI21_X1   g3684(.A1(new_n4069_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n4070_));
  OAI21_X1   g3685(.A1(new_n4070_), .A2(new_n900_), .B(new_n908_), .ZN(new_n4071_));
  AOI21_X1   g3686(.A1(new_n4071_), .A2(new_n913_), .B(new_n918_), .ZN(new_n4072_));
  OAI21_X1   g3687(.A1(new_n4072_), .A2(new_n897_), .B(new_n923_), .ZN(new_n4073_));
  AOI21_X1   g3688(.A1(new_n4073_), .A2(new_n894_), .B(new_n929_), .ZN(new_n4074_));
  OAI21_X1   g3689(.A1(new_n4074_), .A2(new_n933_), .B(new_n937_), .ZN(new_n4075_));
  AOI21_X1   g3690(.A1(new_n4075_), .A2(new_n890_), .B(new_n943_), .ZN(new_n4076_));
  OAI21_X1   g3691(.A1(new_n4076_), .A2(new_n886_), .B(new_n948_), .ZN(new_n4077_));
  AOI21_X1   g3692(.A1(new_n4077_), .A2(new_n953_), .B(new_n958_), .ZN(new_n4078_));
  OAI21_X1   g3693(.A1(new_n4078_), .A2(new_n883_), .B(new_n963_), .ZN(new_n4079_));
  AOI21_X1   g3694(.A1(new_n4079_), .A2(new_n880_), .B(new_n969_), .ZN(new_n4080_));
  OAI21_X1   g3695(.A1(new_n4080_), .A2(new_n973_), .B(new_n977_), .ZN(new_n4081_));
  AOI21_X1   g3696(.A1(new_n4081_), .A2(new_n876_), .B(new_n983_), .ZN(new_n4082_));
  OAI21_X1   g3697(.A1(new_n4082_), .A2(new_n872_), .B(new_n988_), .ZN(new_n4083_));
  AOI21_X1   g3698(.A1(new_n4083_), .A2(new_n993_), .B(new_n998_), .ZN(new_n4084_));
  OAI21_X1   g3699(.A1(new_n4084_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n4085_));
  AOI21_X1   g3700(.A1(new_n4085_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n4086_));
  OAI21_X1   g3701(.A1(new_n4086_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n4087_));
  OAI21_X1   g3702(.A1(new_n1019_), .A2(\priority[57] ), .B(\req[57] ), .ZN(new_n4088_));
  AOI21_X1   g3703(.A1(new_n4087_), .A2(new_n862_), .B(new_n4088_), .ZN(\grant[57] ));
  NOR2_X1    g3704(.A1(new_n1240_), .A2(new_n1027_), .ZN(new_n4090_));
  OAI21_X1   g3705(.A1(new_n1032_), .A2(new_n4090_), .B(new_n1037_), .ZN(new_n4091_));
  AOI21_X1   g3706(.A1(new_n4091_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n4092_));
  OAI21_X1   g3707(.A1(new_n4092_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n4093_));
  AOI21_X1   g3708(.A1(new_n4093_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n4094_));
  OAI21_X1   g3709(.A1(new_n4094_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n4095_));
  AOI21_X1   g3710(.A1(new_n4095_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n4096_));
  OAI21_X1   g3711(.A1(new_n4096_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n4097_));
  AOI21_X1   g3712(.A1(new_n4097_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n4098_));
  OAI21_X1   g3713(.A1(new_n4098_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n4099_));
  AOI21_X1   g3714(.A1(new_n4099_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n4100_));
  OAI21_X1   g3715(.A1(new_n4100_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n4101_));
  AOI21_X1   g3716(.A1(new_n4101_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n4102_));
  OAI21_X1   g3717(.A1(new_n4102_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n4103_));
  AOI21_X1   g3718(.A1(new_n4103_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n4104_));
  OAI21_X1   g3719(.A1(new_n4104_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n4105_));
  AOI21_X1   g3720(.A1(new_n4105_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n4106_));
  OAI21_X1   g3721(.A1(new_n4106_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n4107_));
  AOI21_X1   g3722(.A1(new_n4107_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n4108_));
  OAI21_X1   g3723(.A1(new_n4108_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n4109_));
  AOI21_X1   g3724(.A1(new_n4109_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n4110_));
  OAI21_X1   g3725(.A1(new_n4110_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n4111_));
  AOI21_X1   g3726(.A1(new_n4111_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n4112_));
  OAI21_X1   g3727(.A1(new_n4112_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n4113_));
  AOI21_X1   g3728(.A1(new_n4113_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n4114_));
  OAI21_X1   g3729(.A1(new_n4114_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n4115_));
  AOI21_X1   g3730(.A1(new_n4115_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n4116_));
  OAI21_X1   g3731(.A1(new_n4116_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n4117_));
  AOI21_X1   g3732(.A1(new_n4117_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n4118_));
  OAI21_X1   g3733(.A1(new_n4118_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n4119_));
  AOI21_X1   g3734(.A1(new_n4119_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n4120_));
  OAI21_X1   g3735(.A1(new_n4120_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n4121_));
  AOI21_X1   g3736(.A1(new_n4121_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n4122_));
  OAI21_X1   g3737(.A1(new_n4122_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n4123_));
  AOI21_X1   g3738(.A1(new_n4123_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n4124_));
  OAI21_X1   g3739(.A1(new_n4124_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n4125_));
  AOI21_X1   g3740(.A1(new_n4125_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n4126_));
  OAI21_X1   g3741(.A1(new_n4126_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n4127_));
  AOI21_X1   g3742(.A1(new_n4127_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n4128_));
  OAI21_X1   g3743(.A1(new_n4128_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n4129_));
  AOI21_X1   g3744(.A1(new_n4129_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n4130_));
  OAI21_X1   g3745(.A1(new_n4130_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n4131_));
  OAI21_X1   g3746(.A1(new_n450_), .A2(\priority[58] ), .B(\req[58] ), .ZN(new_n4132_));
  AOI21_X1   g3747(.A1(new_n4131_), .A2(new_n1245_), .B(new_n4132_), .ZN(\grant[58] ));
  NOR2_X1    g3748(.A1(new_n644_), .A2(new_n1389_), .ZN(new_n4134_));
  OAI21_X1   g3749(.A1(new_n1394_), .A2(new_n4134_), .B(new_n1398_), .ZN(new_n4135_));
  AOI21_X1   g3750(.A1(new_n4135_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n4136_));
  OAI21_X1   g3751(.A1(new_n4136_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n4137_));
  AOI21_X1   g3752(.A1(new_n4137_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n4138_));
  OAI21_X1   g3753(.A1(new_n4138_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n4139_));
  AOI21_X1   g3754(.A1(new_n4139_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n4140_));
  OAI21_X1   g3755(.A1(new_n4140_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n4141_));
  AOI21_X1   g3756(.A1(new_n4141_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n4142_));
  OAI21_X1   g3757(.A1(new_n4142_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n4143_));
  AOI21_X1   g3758(.A1(new_n4143_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n4144_));
  OAI21_X1   g3759(.A1(new_n4144_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n4145_));
  AOI21_X1   g3760(.A1(new_n4145_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n4146_));
  OAI21_X1   g3761(.A1(new_n4146_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n4147_));
  AOI21_X1   g3762(.A1(new_n4147_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n4148_));
  OAI21_X1   g3763(.A1(new_n4148_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n4149_));
  AOI21_X1   g3764(.A1(new_n4149_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n4150_));
  OAI21_X1   g3765(.A1(new_n4150_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n4151_));
  AOI21_X1   g3766(.A1(new_n4151_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n4152_));
  OAI21_X1   g3767(.A1(new_n4152_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n4153_));
  AOI21_X1   g3768(.A1(new_n4153_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n4154_));
  OAI21_X1   g3769(.A1(new_n4154_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n4155_));
  AOI21_X1   g3770(.A1(new_n4155_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n4156_));
  OAI21_X1   g3771(.A1(new_n4156_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n4157_));
  AOI21_X1   g3772(.A1(new_n4157_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n4158_));
  OAI21_X1   g3773(.A1(new_n4158_), .A2(new_n519_), .B(new_n524_), .ZN(new_n4159_));
  AOI21_X1   g3774(.A1(new_n4159_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n4160_));
  OAI21_X1   g3775(.A1(new_n4160_), .A2(new_n497_), .B(new_n535_), .ZN(new_n4161_));
  AOI21_X1   g3776(.A1(new_n4161_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n4162_));
  OAI21_X1   g3777(.A1(new_n4162_), .A2(new_n492_), .B(new_n550_), .ZN(new_n4163_));
  AOI21_X1   g3778(.A1(new_n4163_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n4164_));
  OAI21_X1   g3779(.A1(new_n4164_), .A2(new_n561_), .B(new_n566_), .ZN(new_n4165_));
  AOI21_X1   g3780(.A1(new_n4165_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n4166_));
  OAI21_X1   g3781(.A1(new_n4166_), .A2(new_n479_), .B(new_n577_), .ZN(new_n4167_));
  AOI21_X1   g3782(.A1(new_n4167_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n4168_));
  OAI21_X1   g3783(.A1(new_n4168_), .A2(new_n474_), .B(new_n592_), .ZN(new_n4169_));
  AOI21_X1   g3784(.A1(new_n4169_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n4170_));
  OAI21_X1   g3785(.A1(new_n4170_), .A2(new_n603_), .B(new_n608_), .ZN(new_n4171_));
  AOI21_X1   g3786(.A1(new_n4171_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n4172_));
  OAI21_X1   g3787(.A1(new_n4172_), .A2(new_n461_), .B(new_n619_), .ZN(new_n4173_));
  AOI21_X1   g3788(.A1(new_n4173_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n4174_));
  OAI21_X1   g3789(.A1(new_n4174_), .A2(new_n456_), .B(new_n634_), .ZN(new_n4175_));
  OAI21_X1   g3790(.A1(new_n637_), .A2(\priority[59] ), .B(\req[59] ), .ZN(new_n4176_));
  AOI21_X1   g3791(.A1(new_n4175_), .A2(new_n1546_), .B(new_n4176_), .ZN(\grant[59] ));
  NOR2_X1    g3792(.A1(new_n1031_), .A2(new_n649_), .ZN(new_n4178_));
  OAI21_X1   g3793(.A1(new_n448_), .A2(new_n4178_), .B(new_n656_), .ZN(new_n4179_));
  AOI21_X1   g3794(.A1(new_n4179_), .A2(new_n444_), .B(new_n662_), .ZN(new_n4180_));
  OAI21_X1   g3795(.A1(new_n4180_), .A2(new_n667_), .B(new_n671_), .ZN(new_n4181_));
  AOI21_X1   g3796(.A1(new_n4181_), .A2(new_n439_), .B(new_n677_), .ZN(new_n4182_));
  OAI21_X1   g3797(.A1(new_n4182_), .A2(new_n434_), .B(new_n682_), .ZN(new_n4183_));
  AOI21_X1   g3798(.A1(new_n4183_), .A2(new_n688_), .B(new_n693_), .ZN(new_n4184_));
  OAI21_X1   g3799(.A1(new_n4184_), .A2(new_n430_), .B(new_n698_), .ZN(new_n4185_));
  AOI21_X1   g3800(.A1(new_n4185_), .A2(new_n426_), .B(new_n704_), .ZN(new_n4186_));
  OAI21_X1   g3801(.A1(new_n4186_), .A2(new_n709_), .B(new_n713_), .ZN(new_n4187_));
  AOI21_X1   g3802(.A1(new_n4187_), .A2(new_n421_), .B(new_n719_), .ZN(new_n4188_));
  OAI21_X1   g3803(.A1(new_n4188_), .A2(new_n416_), .B(new_n724_), .ZN(new_n4189_));
  AOI21_X1   g3804(.A1(new_n4189_), .A2(new_n730_), .B(new_n735_), .ZN(new_n4190_));
  OAI21_X1   g3805(.A1(new_n4190_), .A2(new_n412_), .B(new_n740_), .ZN(new_n4191_));
  AOI21_X1   g3806(.A1(new_n4191_), .A2(new_n408_), .B(new_n746_), .ZN(new_n4192_));
  OAI21_X1   g3807(.A1(new_n4192_), .A2(new_n751_), .B(new_n755_), .ZN(new_n4193_));
  AOI21_X1   g3808(.A1(new_n4193_), .A2(new_n403_), .B(new_n761_), .ZN(new_n4194_));
  OAI21_X1   g3809(.A1(new_n4194_), .A2(new_n398_), .B(new_n766_), .ZN(new_n4195_));
  AOI21_X1   g3810(.A1(new_n4195_), .A2(new_n772_), .B(new_n777_), .ZN(new_n4196_));
  OAI21_X1   g3811(.A1(new_n4196_), .A2(new_n394_), .B(new_n782_), .ZN(new_n4197_));
  AOI21_X1   g3812(.A1(new_n4197_), .A2(new_n390_), .B(new_n788_), .ZN(new_n4198_));
  OAI21_X1   g3813(.A1(new_n4198_), .A2(new_n793_), .B(new_n797_), .ZN(new_n4199_));
  AOI21_X1   g3814(.A1(new_n4199_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n4200_));
  OAI21_X1   g3815(.A1(new_n4200_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n4201_));
  AOI21_X1   g3816(.A1(new_n4201_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n4202_));
  OAI21_X1   g3817(.A1(new_n4202_), .A2(new_n912_), .B(new_n917_), .ZN(new_n4203_));
  AOI21_X1   g3818(.A1(new_n4203_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n4204_));
  OAI21_X1   g3819(.A1(new_n4204_), .A2(new_n893_), .B(new_n928_), .ZN(new_n4205_));
  AOI21_X1   g3820(.A1(new_n4205_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n4206_));
  OAI21_X1   g3821(.A1(new_n4206_), .A2(new_n889_), .B(new_n942_), .ZN(new_n4207_));
  AOI21_X1   g3822(.A1(new_n4207_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n4208_));
  OAI21_X1   g3823(.A1(new_n4208_), .A2(new_n952_), .B(new_n957_), .ZN(new_n4209_));
  AOI21_X1   g3824(.A1(new_n4209_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n4210_));
  OAI21_X1   g3825(.A1(new_n4210_), .A2(new_n879_), .B(new_n968_), .ZN(new_n4211_));
  AOI21_X1   g3826(.A1(new_n4211_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n4212_));
  OAI21_X1   g3827(.A1(new_n4212_), .A2(new_n875_), .B(new_n982_), .ZN(new_n4213_));
  AOI21_X1   g3828(.A1(new_n4213_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n4214_));
  OAI21_X1   g3829(.A1(new_n4214_), .A2(new_n992_), .B(new_n997_), .ZN(new_n4215_));
  AOI21_X1   g3830(.A1(new_n4215_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n4216_));
  OAI21_X1   g3831(.A1(new_n4216_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n4217_));
  AOI21_X1   g3832(.A1(new_n4217_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n4218_));
  OAI21_X1   g3833(.A1(new_n4218_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n4219_));
  OAI21_X1   g3834(.A1(new_n1025_), .A2(\priority[60] ), .B(\req[60] ), .ZN(new_n4220_));
  AOI21_X1   g3835(.A1(new_n4219_), .A2(new_n1636_), .B(new_n4220_), .ZN(\grant[60] ));
  NOR2_X1    g3836(.A1(new_n1393_), .A2(new_n1036_), .ZN(new_n4222_));
  OAI21_X1   g3837(.A1(new_n855_), .A2(new_n4222_), .B(new_n1043_), .ZN(new_n4223_));
  AOI21_X1   g3838(.A1(new_n4223_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n4224_));
  OAI21_X1   g3839(.A1(new_n4224_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n4225_));
  AOI21_X1   g3840(.A1(new_n4225_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n4226_));
  OAI21_X1   g3841(.A1(new_n4226_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n4227_));
  AOI21_X1   g3842(.A1(new_n4227_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n4228_));
  OAI21_X1   g3843(.A1(new_n4228_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n4229_));
  AOI21_X1   g3844(.A1(new_n4229_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n4230_));
  OAI21_X1   g3845(.A1(new_n4230_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n4231_));
  AOI21_X1   g3846(.A1(new_n4231_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n4232_));
  OAI21_X1   g3847(.A1(new_n4232_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n4233_));
  AOI21_X1   g3848(.A1(new_n4233_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n4234_));
  OAI21_X1   g3849(.A1(new_n4234_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n4235_));
  AOI21_X1   g3850(.A1(new_n4235_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n4236_));
  OAI21_X1   g3851(.A1(new_n4236_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n4237_));
  AOI21_X1   g3852(.A1(new_n4237_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n4238_));
  OAI21_X1   g3853(.A1(new_n4238_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n4239_));
  AOI21_X1   g3854(.A1(new_n4239_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n4240_));
  OAI21_X1   g3855(.A1(new_n4240_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n4241_));
  AOI21_X1   g3856(.A1(new_n4241_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n4242_));
  OAI21_X1   g3857(.A1(new_n4242_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n4243_));
  AOI21_X1   g3858(.A1(new_n4243_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n4244_));
  OAI21_X1   g3859(.A1(new_n4244_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n4245_));
  AOI21_X1   g3860(.A1(new_n4245_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n4246_));
  OAI21_X1   g3861(.A1(new_n4246_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n4247_));
  AOI21_X1   g3862(.A1(new_n4247_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n4248_));
  OAI21_X1   g3863(.A1(new_n4248_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n4249_));
  AOI21_X1   g3864(.A1(new_n4249_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n4250_));
  OAI21_X1   g3865(.A1(new_n4250_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n4251_));
  AOI21_X1   g3866(.A1(new_n4251_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n4252_));
  OAI21_X1   g3867(.A1(new_n4252_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n4253_));
  AOI21_X1   g3868(.A1(new_n4253_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n4254_));
  OAI21_X1   g3869(.A1(new_n4254_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n4255_));
  AOI21_X1   g3870(.A1(new_n4255_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n4256_));
  OAI21_X1   g3871(.A1(new_n4256_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n4257_));
  AOI21_X1   g3872(.A1(new_n4257_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n4258_));
  OAI21_X1   g3873(.A1(new_n4258_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n4259_));
  AOI21_X1   g3874(.A1(new_n4259_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n4260_));
  OAI21_X1   g3875(.A1(new_n4260_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n4261_));
  AOI21_X1   g3876(.A1(new_n4261_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n4262_));
  OAI21_X1   g3877(.A1(new_n4262_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n4263_));
  OAI21_X1   g3878(.A1(new_n643_), .A2(\priority[61] ), .B(\req[61] ), .ZN(new_n4264_));
  AOI21_X1   g3879(.A1(new_n4263_), .A2(new_n1724_), .B(new_n4264_), .ZN(\grant[61] ));
  NOR2_X1    g3880(.A1(new_n447_), .A2(new_n1397_), .ZN(new_n4266_));
  OAI21_X1   g3881(.A1(new_n1238_), .A2(new_n4266_), .B(new_n1403_), .ZN(new_n4267_));
  AOI21_X1   g3882(.A1(new_n4267_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n4268_));
  OAI21_X1   g3883(.A1(new_n4268_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n4269_));
  AOI21_X1   g3884(.A1(new_n4269_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n4270_));
  OAI21_X1   g3885(.A1(new_n4270_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n4271_));
  AOI21_X1   g3886(.A1(new_n4271_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n4272_));
  OAI21_X1   g3887(.A1(new_n4272_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n4273_));
  AOI21_X1   g3888(.A1(new_n4273_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n4274_));
  OAI21_X1   g3889(.A1(new_n4274_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n4275_));
  AOI21_X1   g3890(.A1(new_n4275_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n4276_));
  OAI21_X1   g3891(.A1(new_n4276_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n4277_));
  AOI21_X1   g3892(.A1(new_n4277_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n4278_));
  OAI21_X1   g3893(.A1(new_n4278_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n4279_));
  AOI21_X1   g3894(.A1(new_n4279_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n4280_));
  OAI21_X1   g3895(.A1(new_n4280_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n4281_));
  AOI21_X1   g3896(.A1(new_n4281_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n4282_));
  OAI21_X1   g3897(.A1(new_n4282_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n4283_));
  AOI21_X1   g3898(.A1(new_n4283_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n4284_));
  OAI21_X1   g3899(.A1(new_n4284_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n4285_));
  AOI21_X1   g3900(.A1(new_n4285_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n4286_));
  OAI21_X1   g3901(.A1(new_n4286_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n4287_));
  AOI21_X1   g3902(.A1(new_n4287_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n4288_));
  OAI21_X1   g3903(.A1(new_n4288_), .A2(new_n506_), .B(new_n514_), .ZN(new_n4289_));
  AOI21_X1   g3904(.A1(new_n4289_), .A2(new_n520_), .B(new_n525_), .ZN(new_n4290_));
  OAI21_X1   g3905(.A1(new_n4290_), .A2(new_n502_), .B(new_n530_), .ZN(new_n4291_));
  AOI21_X1   g3906(.A1(new_n4291_), .A2(new_n498_), .B(new_n536_), .ZN(new_n4292_));
  OAI21_X1   g3907(.A1(new_n4292_), .A2(new_n541_), .B(new_n545_), .ZN(new_n4293_));
  AOI21_X1   g3908(.A1(new_n4293_), .A2(new_n493_), .B(new_n551_), .ZN(new_n4294_));
  OAI21_X1   g3909(.A1(new_n4294_), .A2(new_n488_), .B(new_n556_), .ZN(new_n4295_));
  AOI21_X1   g3910(.A1(new_n4295_), .A2(new_n562_), .B(new_n567_), .ZN(new_n4296_));
  OAI21_X1   g3911(.A1(new_n4296_), .A2(new_n484_), .B(new_n572_), .ZN(new_n4297_));
  AOI21_X1   g3912(.A1(new_n4297_), .A2(new_n480_), .B(new_n578_), .ZN(new_n4298_));
  OAI21_X1   g3913(.A1(new_n4298_), .A2(new_n583_), .B(new_n587_), .ZN(new_n4299_));
  AOI21_X1   g3914(.A1(new_n4299_), .A2(new_n475_), .B(new_n593_), .ZN(new_n4300_));
  OAI21_X1   g3915(.A1(new_n4300_), .A2(new_n470_), .B(new_n598_), .ZN(new_n4301_));
  AOI21_X1   g3916(.A1(new_n4301_), .A2(new_n604_), .B(new_n609_), .ZN(new_n4302_));
  OAI21_X1   g3917(.A1(new_n4302_), .A2(new_n466_), .B(new_n614_), .ZN(new_n4303_));
  AOI21_X1   g3918(.A1(new_n4303_), .A2(new_n462_), .B(new_n620_), .ZN(new_n4304_));
  OAI21_X1   g3919(.A1(new_n4304_), .A2(new_n625_), .B(new_n629_), .ZN(new_n4305_));
  AOI21_X1   g3920(.A1(new_n4305_), .A2(new_n457_), .B(new_n635_), .ZN(new_n4306_));
  OAI21_X1   g3921(.A1(new_n4306_), .A2(new_n452_), .B(new_n640_), .ZN(new_n4307_));
  OAI21_X1   g3922(.A1(new_n647_), .A2(\priority[62] ), .B(\req[62] ), .ZN(new_n4308_));
  AOI21_X1   g3923(.A1(new_n4307_), .A2(new_n646_), .B(new_n4308_), .ZN(\grant[62] ));
  NOR2_X1    g3924(.A1(new_n854_), .A2(new_n655_), .ZN(new_n4310_));
  OAI21_X1   g3925(.A1(new_n443_), .A2(new_n4310_), .B(new_n661_), .ZN(new_n4311_));
  AOI21_X1   g3926(.A1(new_n4311_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n4312_));
  OAI21_X1   g3927(.A1(new_n4312_), .A2(new_n438_), .B(new_n676_), .ZN(new_n4313_));
  AOI21_X1   g3928(.A1(new_n4313_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n4314_));
  OAI21_X1   g3929(.A1(new_n4314_), .A2(new_n687_), .B(new_n692_), .ZN(new_n4315_));
  AOI21_X1   g3930(.A1(new_n4315_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n4316_));
  OAI21_X1   g3931(.A1(new_n4316_), .A2(new_n425_), .B(new_n703_), .ZN(new_n4317_));
  AOI21_X1   g3932(.A1(new_n4317_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n4318_));
  OAI21_X1   g3933(.A1(new_n4318_), .A2(new_n420_), .B(new_n718_), .ZN(new_n4319_));
  AOI21_X1   g3934(.A1(new_n4319_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n4320_));
  OAI21_X1   g3935(.A1(new_n4320_), .A2(new_n729_), .B(new_n734_), .ZN(new_n4321_));
  AOI21_X1   g3936(.A1(new_n4321_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n4322_));
  OAI21_X1   g3937(.A1(new_n4322_), .A2(new_n407_), .B(new_n745_), .ZN(new_n4323_));
  AOI21_X1   g3938(.A1(new_n4323_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n4324_));
  OAI21_X1   g3939(.A1(new_n4324_), .A2(new_n402_), .B(new_n760_), .ZN(new_n4325_));
  AOI21_X1   g3940(.A1(new_n4325_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n4326_));
  OAI21_X1   g3941(.A1(new_n4326_), .A2(new_n771_), .B(new_n776_), .ZN(new_n4327_));
  AOI21_X1   g3942(.A1(new_n4327_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n4328_));
  OAI21_X1   g3943(.A1(new_n4328_), .A2(new_n389_), .B(new_n787_), .ZN(new_n4329_));
  AOI21_X1   g3944(.A1(new_n4329_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n4330_));
  OAI21_X1   g3945(.A1(new_n4330_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n4331_));
  AOI21_X1   g3946(.A1(new_n4331_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n4332_));
  OAI21_X1   g3947(.A1(new_n4332_), .A2(new_n900_), .B(new_n908_), .ZN(new_n4333_));
  AOI21_X1   g3948(.A1(new_n4333_), .A2(new_n913_), .B(new_n918_), .ZN(new_n4334_));
  OAI21_X1   g3949(.A1(new_n4334_), .A2(new_n897_), .B(new_n923_), .ZN(new_n4335_));
  AOI21_X1   g3950(.A1(new_n4335_), .A2(new_n894_), .B(new_n929_), .ZN(new_n4336_));
  OAI21_X1   g3951(.A1(new_n4336_), .A2(new_n933_), .B(new_n937_), .ZN(new_n4337_));
  AOI21_X1   g3952(.A1(new_n4337_), .A2(new_n890_), .B(new_n943_), .ZN(new_n4338_));
  OAI21_X1   g3953(.A1(new_n4338_), .A2(new_n886_), .B(new_n948_), .ZN(new_n4339_));
  AOI21_X1   g3954(.A1(new_n4339_), .A2(new_n953_), .B(new_n958_), .ZN(new_n4340_));
  OAI21_X1   g3955(.A1(new_n4340_), .A2(new_n883_), .B(new_n963_), .ZN(new_n4341_));
  AOI21_X1   g3956(.A1(new_n4341_), .A2(new_n880_), .B(new_n969_), .ZN(new_n4342_));
  OAI21_X1   g3957(.A1(new_n4342_), .A2(new_n973_), .B(new_n977_), .ZN(new_n4343_));
  AOI21_X1   g3958(.A1(new_n4343_), .A2(new_n876_), .B(new_n983_), .ZN(new_n4344_));
  OAI21_X1   g3959(.A1(new_n4344_), .A2(new_n872_), .B(new_n988_), .ZN(new_n4345_));
  AOI21_X1   g3960(.A1(new_n4345_), .A2(new_n993_), .B(new_n998_), .ZN(new_n4346_));
  OAI21_X1   g3961(.A1(new_n4346_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n4347_));
  AOI21_X1   g3962(.A1(new_n4347_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n4348_));
  OAI21_X1   g3963(.A1(new_n4348_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n4349_));
  AOI21_X1   g3964(.A1(new_n4349_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n4350_));
  OAI21_X1   g3965(.A1(new_n4350_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n4351_));
  OAI21_X1   g3966(.A1(new_n1034_), .A2(\priority[63] ), .B(\req[63] ), .ZN(new_n4352_));
  AOI21_X1   g3967(.A1(new_n4351_), .A2(new_n1033_), .B(new_n4352_), .ZN(\grant[63] ));
  NOR2_X1    g3968(.A1(new_n1237_), .A2(new_n1042_), .ZN(new_n4354_));
  OAI21_X1   g3969(.A1(new_n851_), .A2(new_n4354_), .B(new_n1048_), .ZN(new_n4355_));
  AOI21_X1   g3970(.A1(new_n4355_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n4356_));
  OAI21_X1   g3971(.A1(new_n4356_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n4357_));
  AOI21_X1   g3972(.A1(new_n4357_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n4358_));
  OAI21_X1   g3973(.A1(new_n4358_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n4359_));
  AOI21_X1   g3974(.A1(new_n4359_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n4360_));
  OAI21_X1   g3975(.A1(new_n4360_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n4361_));
  AOI21_X1   g3976(.A1(new_n4361_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n4362_));
  OAI21_X1   g3977(.A1(new_n4362_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n4363_));
  AOI21_X1   g3978(.A1(new_n4363_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n4364_));
  OAI21_X1   g3979(.A1(new_n4364_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n4365_));
  AOI21_X1   g3980(.A1(new_n4365_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n4366_));
  OAI21_X1   g3981(.A1(new_n4366_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n4367_));
  AOI21_X1   g3982(.A1(new_n4367_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n4368_));
  OAI21_X1   g3983(.A1(new_n4368_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n4369_));
  AOI21_X1   g3984(.A1(new_n4369_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n4370_));
  OAI21_X1   g3985(.A1(new_n4370_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n4371_));
  AOI21_X1   g3986(.A1(new_n4371_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n4372_));
  OAI21_X1   g3987(.A1(new_n4372_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n4373_));
  AOI21_X1   g3988(.A1(new_n4373_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n4374_));
  OAI21_X1   g3989(.A1(new_n4374_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n4375_));
  AOI21_X1   g3990(.A1(new_n4375_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n4376_));
  OAI21_X1   g3991(.A1(new_n4376_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n4377_));
  AOI21_X1   g3992(.A1(new_n4377_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n4378_));
  OAI21_X1   g3993(.A1(new_n4378_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n4379_));
  AOI21_X1   g3994(.A1(new_n4379_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n4380_));
  OAI21_X1   g3995(.A1(new_n4380_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n4381_));
  AOI21_X1   g3996(.A1(new_n4381_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n4382_));
  OAI21_X1   g3997(.A1(new_n4382_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n4383_));
  AOI21_X1   g3998(.A1(new_n4383_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n4384_));
  OAI21_X1   g3999(.A1(new_n4384_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n4385_));
  AOI21_X1   g4000(.A1(new_n4385_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n4386_));
  OAI21_X1   g4001(.A1(new_n4386_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n4387_));
  AOI21_X1   g4002(.A1(new_n4387_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n4388_));
  OAI21_X1   g4003(.A1(new_n4388_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n4389_));
  AOI21_X1   g4004(.A1(new_n4389_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n4390_));
  OAI21_X1   g4005(.A1(new_n4390_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n4391_));
  AOI21_X1   g4006(.A1(new_n4391_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n4392_));
  OAI21_X1   g4007(.A1(new_n4392_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n4393_));
  AOI21_X1   g4008(.A1(new_n4393_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n4394_));
  OAI21_X1   g4009(.A1(new_n4394_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n4395_));
  OAI21_X1   g4010(.A1(new_n446_), .A2(\priority[64] ), .B(\req[64] ), .ZN(new_n4396_));
  AOI21_X1   g4011(.A1(new_n4395_), .A2(new_n1395_), .B(new_n4396_), .ZN(\grant[64] ));
  NOR2_X1    g4012(.A1(new_n442_), .A2(new_n1402_), .ZN(new_n4398_));
  OAI21_X1   g4013(.A1(new_n1234_), .A2(new_n4398_), .B(new_n1407_), .ZN(new_n4399_));
  AOI21_X1   g4014(.A1(new_n4399_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n4400_));
  OAI21_X1   g4015(.A1(new_n4400_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n4401_));
  AOI21_X1   g4016(.A1(new_n4401_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n4402_));
  OAI21_X1   g4017(.A1(new_n4402_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n4403_));
  AOI21_X1   g4018(.A1(new_n4403_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n4404_));
  OAI21_X1   g4019(.A1(new_n4404_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n4405_));
  AOI21_X1   g4020(.A1(new_n4405_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n4406_));
  OAI21_X1   g4021(.A1(new_n4406_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n4407_));
  AOI21_X1   g4022(.A1(new_n4407_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n4408_));
  OAI21_X1   g4023(.A1(new_n4408_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n4409_));
  AOI21_X1   g4024(.A1(new_n4409_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n4410_));
  OAI21_X1   g4025(.A1(new_n4410_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n4411_));
  AOI21_X1   g4026(.A1(new_n4411_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n4412_));
  OAI21_X1   g4027(.A1(new_n4412_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n4413_));
  AOI21_X1   g4028(.A1(new_n4413_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n4414_));
  OAI21_X1   g4029(.A1(new_n4414_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n4415_));
  AOI21_X1   g4030(.A1(new_n4415_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n4416_));
  OAI21_X1   g4031(.A1(new_n4416_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n4417_));
  AOI21_X1   g4032(.A1(new_n4417_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n4418_));
  OAI21_X1   g4033(.A1(new_n4418_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n4419_));
  AOI21_X1   g4034(.A1(new_n4419_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n4420_));
  OAI21_X1   g4035(.A1(new_n4420_), .A2(new_n519_), .B(new_n524_), .ZN(new_n4421_));
  AOI21_X1   g4036(.A1(new_n4421_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n4422_));
  OAI21_X1   g4037(.A1(new_n4422_), .A2(new_n497_), .B(new_n535_), .ZN(new_n4423_));
  AOI21_X1   g4038(.A1(new_n4423_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n4424_));
  OAI21_X1   g4039(.A1(new_n4424_), .A2(new_n492_), .B(new_n550_), .ZN(new_n4425_));
  AOI21_X1   g4040(.A1(new_n4425_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n4426_));
  OAI21_X1   g4041(.A1(new_n4426_), .A2(new_n561_), .B(new_n566_), .ZN(new_n4427_));
  AOI21_X1   g4042(.A1(new_n4427_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n4428_));
  OAI21_X1   g4043(.A1(new_n4428_), .A2(new_n479_), .B(new_n577_), .ZN(new_n4429_));
  AOI21_X1   g4044(.A1(new_n4429_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n4430_));
  OAI21_X1   g4045(.A1(new_n4430_), .A2(new_n474_), .B(new_n592_), .ZN(new_n4431_));
  AOI21_X1   g4046(.A1(new_n4431_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n4432_));
  OAI21_X1   g4047(.A1(new_n4432_), .A2(new_n603_), .B(new_n608_), .ZN(new_n4433_));
  AOI21_X1   g4048(.A1(new_n4433_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n4434_));
  OAI21_X1   g4049(.A1(new_n4434_), .A2(new_n461_), .B(new_n619_), .ZN(new_n4435_));
  AOI21_X1   g4050(.A1(new_n4435_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n4436_));
  OAI21_X1   g4051(.A1(new_n4436_), .A2(new_n456_), .B(new_n634_), .ZN(new_n4437_));
  AOI21_X1   g4052(.A1(new_n4437_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n4438_));
  OAI21_X1   g4053(.A1(new_n4438_), .A2(new_n645_), .B(new_n650_), .ZN(new_n4439_));
  OAI21_X1   g4054(.A1(new_n653_), .A2(\priority[65] ), .B(\req[65] ), .ZN(new_n4440_));
  AOI21_X1   g4055(.A1(new_n4439_), .A2(new_n1544_), .B(new_n4440_), .ZN(\grant[65] ));
  NOR2_X1    g4056(.A1(new_n850_), .A2(new_n660_), .ZN(new_n4442_));
  OAI21_X1   g4057(.A1(new_n667_), .A2(new_n4442_), .B(new_n671_), .ZN(new_n4443_));
  AOI21_X1   g4058(.A1(new_n4443_), .A2(new_n439_), .B(new_n677_), .ZN(new_n4444_));
  OAI21_X1   g4059(.A1(new_n4444_), .A2(new_n434_), .B(new_n682_), .ZN(new_n4445_));
  AOI21_X1   g4060(.A1(new_n4445_), .A2(new_n688_), .B(new_n693_), .ZN(new_n4446_));
  OAI21_X1   g4061(.A1(new_n4446_), .A2(new_n430_), .B(new_n698_), .ZN(new_n4447_));
  AOI21_X1   g4062(.A1(new_n4447_), .A2(new_n426_), .B(new_n704_), .ZN(new_n4448_));
  OAI21_X1   g4063(.A1(new_n4448_), .A2(new_n709_), .B(new_n713_), .ZN(new_n4449_));
  AOI21_X1   g4064(.A1(new_n4449_), .A2(new_n421_), .B(new_n719_), .ZN(new_n4450_));
  OAI21_X1   g4065(.A1(new_n4450_), .A2(new_n416_), .B(new_n724_), .ZN(new_n4451_));
  AOI21_X1   g4066(.A1(new_n4451_), .A2(new_n730_), .B(new_n735_), .ZN(new_n4452_));
  OAI21_X1   g4067(.A1(new_n4452_), .A2(new_n412_), .B(new_n740_), .ZN(new_n4453_));
  AOI21_X1   g4068(.A1(new_n4453_), .A2(new_n408_), .B(new_n746_), .ZN(new_n4454_));
  OAI21_X1   g4069(.A1(new_n4454_), .A2(new_n751_), .B(new_n755_), .ZN(new_n4455_));
  AOI21_X1   g4070(.A1(new_n4455_), .A2(new_n403_), .B(new_n761_), .ZN(new_n4456_));
  OAI21_X1   g4071(.A1(new_n4456_), .A2(new_n398_), .B(new_n766_), .ZN(new_n4457_));
  AOI21_X1   g4072(.A1(new_n4457_), .A2(new_n772_), .B(new_n777_), .ZN(new_n4458_));
  OAI21_X1   g4073(.A1(new_n4458_), .A2(new_n394_), .B(new_n782_), .ZN(new_n4459_));
  AOI21_X1   g4074(.A1(new_n4459_), .A2(new_n390_), .B(new_n788_), .ZN(new_n4460_));
  OAI21_X1   g4075(.A1(new_n4460_), .A2(new_n793_), .B(new_n797_), .ZN(new_n4461_));
  AOI21_X1   g4076(.A1(new_n4461_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n4462_));
  OAI21_X1   g4077(.A1(new_n4462_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n4463_));
  AOI21_X1   g4078(.A1(new_n4463_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n4464_));
  OAI21_X1   g4079(.A1(new_n4464_), .A2(new_n912_), .B(new_n917_), .ZN(new_n4465_));
  AOI21_X1   g4080(.A1(new_n4465_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n4466_));
  OAI21_X1   g4081(.A1(new_n4466_), .A2(new_n893_), .B(new_n928_), .ZN(new_n4467_));
  AOI21_X1   g4082(.A1(new_n4467_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n4468_));
  OAI21_X1   g4083(.A1(new_n4468_), .A2(new_n889_), .B(new_n942_), .ZN(new_n4469_));
  AOI21_X1   g4084(.A1(new_n4469_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n4470_));
  OAI21_X1   g4085(.A1(new_n4470_), .A2(new_n952_), .B(new_n957_), .ZN(new_n4471_));
  AOI21_X1   g4086(.A1(new_n4471_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n4472_));
  OAI21_X1   g4087(.A1(new_n4472_), .A2(new_n879_), .B(new_n968_), .ZN(new_n4473_));
  AOI21_X1   g4088(.A1(new_n4473_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n4474_));
  OAI21_X1   g4089(.A1(new_n4474_), .A2(new_n875_), .B(new_n982_), .ZN(new_n4475_));
  AOI21_X1   g4090(.A1(new_n4475_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n4476_));
  OAI21_X1   g4091(.A1(new_n4476_), .A2(new_n992_), .B(new_n997_), .ZN(new_n4477_));
  AOI21_X1   g4092(.A1(new_n4477_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n4478_));
  OAI21_X1   g4093(.A1(new_n4478_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n4479_));
  AOI21_X1   g4094(.A1(new_n4479_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n4480_));
  OAI21_X1   g4095(.A1(new_n4480_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n4481_));
  AOI21_X1   g4096(.A1(new_n4481_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n4482_));
  OAI21_X1   g4097(.A1(new_n4482_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n4483_));
  OAI21_X1   g4098(.A1(new_n1040_), .A2(\priority[66] ), .B(\req[66] ), .ZN(new_n4484_));
  AOI21_X1   g4099(.A1(new_n4483_), .A2(new_n1634_), .B(new_n4484_), .ZN(\grant[66] ));
  NOR2_X1    g4100(.A1(new_n1233_), .A2(new_n1047_), .ZN(new_n4486_));
  OAI21_X1   g4101(.A1(new_n1053_), .A2(new_n4486_), .B(new_n1057_), .ZN(new_n4487_));
  AOI21_X1   g4102(.A1(new_n4487_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n4488_));
  OAI21_X1   g4103(.A1(new_n4488_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n4489_));
  AOI21_X1   g4104(.A1(new_n4489_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n4490_));
  OAI21_X1   g4105(.A1(new_n4490_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n4491_));
  AOI21_X1   g4106(.A1(new_n4491_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n4492_));
  OAI21_X1   g4107(.A1(new_n4492_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n4493_));
  AOI21_X1   g4108(.A1(new_n4493_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n4494_));
  OAI21_X1   g4109(.A1(new_n4494_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n4495_));
  AOI21_X1   g4110(.A1(new_n4495_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n4496_));
  OAI21_X1   g4111(.A1(new_n4496_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n4497_));
  AOI21_X1   g4112(.A1(new_n4497_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n4498_));
  OAI21_X1   g4113(.A1(new_n4498_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n4499_));
  AOI21_X1   g4114(.A1(new_n4499_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n4500_));
  OAI21_X1   g4115(.A1(new_n4500_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n4501_));
  AOI21_X1   g4116(.A1(new_n4501_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n4502_));
  OAI21_X1   g4117(.A1(new_n4502_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n4503_));
  AOI21_X1   g4118(.A1(new_n4503_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n4504_));
  OAI21_X1   g4119(.A1(new_n4504_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n4505_));
  AOI21_X1   g4120(.A1(new_n4505_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n4506_));
  OAI21_X1   g4121(.A1(new_n4506_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n4507_));
  AOI21_X1   g4122(.A1(new_n4507_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n4508_));
  OAI21_X1   g4123(.A1(new_n4508_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n4509_));
  AOI21_X1   g4124(.A1(new_n4509_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n4510_));
  OAI21_X1   g4125(.A1(new_n4510_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n4511_));
  AOI21_X1   g4126(.A1(new_n4511_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n4512_));
  OAI21_X1   g4127(.A1(new_n4512_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n4513_));
  AOI21_X1   g4128(.A1(new_n4513_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n4514_));
  OAI21_X1   g4129(.A1(new_n4514_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n4515_));
  AOI21_X1   g4130(.A1(new_n4515_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n4516_));
  OAI21_X1   g4131(.A1(new_n4516_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n4517_));
  AOI21_X1   g4132(.A1(new_n4517_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n4518_));
  OAI21_X1   g4133(.A1(new_n4518_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n4519_));
  AOI21_X1   g4134(.A1(new_n4519_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n4520_));
  OAI21_X1   g4135(.A1(new_n4520_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n4521_));
  AOI21_X1   g4136(.A1(new_n4521_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n4522_));
  OAI21_X1   g4137(.A1(new_n4522_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n4523_));
  AOI21_X1   g4138(.A1(new_n4523_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n4524_));
  OAI21_X1   g4139(.A1(new_n4524_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n4525_));
  AOI21_X1   g4140(.A1(new_n4525_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n4526_));
  OAI21_X1   g4141(.A1(new_n4526_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n4527_));
  OAI21_X1   g4142(.A1(new_n441_), .A2(\priority[67] ), .B(\req[67] ), .ZN(new_n4528_));
  AOI21_X1   g4143(.A1(new_n4527_), .A2(new_n1722_), .B(new_n4528_), .ZN(\grant[67] ));
  NOR2_X1    g4144(.A1(new_n666_), .A2(new_n1406_), .ZN(new_n4530_));
  OAI21_X1   g4145(.A1(new_n1412_), .A2(new_n4530_), .B(new_n1415_), .ZN(new_n4531_));
  AOI21_X1   g4146(.A1(new_n4531_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n4532_));
  OAI21_X1   g4147(.A1(new_n4532_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n4533_));
  AOI21_X1   g4148(.A1(new_n4533_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n4534_));
  OAI21_X1   g4149(.A1(new_n4534_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n4535_));
  AOI21_X1   g4150(.A1(new_n4535_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n4536_));
  OAI21_X1   g4151(.A1(new_n4536_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n4537_));
  AOI21_X1   g4152(.A1(new_n4537_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n4538_));
  OAI21_X1   g4153(.A1(new_n4538_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n4539_));
  AOI21_X1   g4154(.A1(new_n4539_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n4540_));
  OAI21_X1   g4155(.A1(new_n4540_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n4541_));
  AOI21_X1   g4156(.A1(new_n4541_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n4542_));
  OAI21_X1   g4157(.A1(new_n4542_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n4543_));
  AOI21_X1   g4158(.A1(new_n4543_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n4544_));
  OAI21_X1   g4159(.A1(new_n4544_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n4545_));
  AOI21_X1   g4160(.A1(new_n4545_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n4546_));
  OAI21_X1   g4161(.A1(new_n4546_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n4547_));
  AOI21_X1   g4162(.A1(new_n4547_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n4548_));
  OAI21_X1   g4163(.A1(new_n4548_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n4549_));
  AOI21_X1   g4164(.A1(new_n4549_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n4550_));
  OAI21_X1   g4165(.A1(new_n4550_), .A2(new_n506_), .B(new_n514_), .ZN(new_n4551_));
  AOI21_X1   g4166(.A1(new_n4551_), .A2(new_n520_), .B(new_n525_), .ZN(new_n4552_));
  OAI21_X1   g4167(.A1(new_n4552_), .A2(new_n502_), .B(new_n530_), .ZN(new_n4553_));
  AOI21_X1   g4168(.A1(new_n4553_), .A2(new_n498_), .B(new_n536_), .ZN(new_n4554_));
  OAI21_X1   g4169(.A1(new_n4554_), .A2(new_n541_), .B(new_n545_), .ZN(new_n4555_));
  AOI21_X1   g4170(.A1(new_n4555_), .A2(new_n493_), .B(new_n551_), .ZN(new_n4556_));
  OAI21_X1   g4171(.A1(new_n4556_), .A2(new_n488_), .B(new_n556_), .ZN(new_n4557_));
  AOI21_X1   g4172(.A1(new_n4557_), .A2(new_n562_), .B(new_n567_), .ZN(new_n4558_));
  OAI21_X1   g4173(.A1(new_n4558_), .A2(new_n484_), .B(new_n572_), .ZN(new_n4559_));
  AOI21_X1   g4174(.A1(new_n4559_), .A2(new_n480_), .B(new_n578_), .ZN(new_n4560_));
  OAI21_X1   g4175(.A1(new_n4560_), .A2(new_n583_), .B(new_n587_), .ZN(new_n4561_));
  AOI21_X1   g4176(.A1(new_n4561_), .A2(new_n475_), .B(new_n593_), .ZN(new_n4562_));
  OAI21_X1   g4177(.A1(new_n4562_), .A2(new_n470_), .B(new_n598_), .ZN(new_n4563_));
  AOI21_X1   g4178(.A1(new_n4563_), .A2(new_n604_), .B(new_n609_), .ZN(new_n4564_));
  OAI21_X1   g4179(.A1(new_n4564_), .A2(new_n466_), .B(new_n614_), .ZN(new_n4565_));
  AOI21_X1   g4180(.A1(new_n4565_), .A2(new_n462_), .B(new_n620_), .ZN(new_n4566_));
  OAI21_X1   g4181(.A1(new_n4566_), .A2(new_n625_), .B(new_n629_), .ZN(new_n4567_));
  AOI21_X1   g4182(.A1(new_n4567_), .A2(new_n457_), .B(new_n635_), .ZN(new_n4568_));
  OAI21_X1   g4183(.A1(new_n4568_), .A2(new_n452_), .B(new_n640_), .ZN(new_n4569_));
  AOI21_X1   g4184(.A1(new_n4569_), .A2(new_n646_), .B(new_n651_), .ZN(new_n4570_));
  OAI21_X1   g4185(.A1(new_n4570_), .A2(new_n448_), .B(new_n656_), .ZN(new_n4571_));
  OAI21_X1   g4186(.A1(new_n658_), .A2(\priority[68] ), .B(\req[68] ), .ZN(new_n4572_));
  AOI21_X1   g4187(.A1(new_n4571_), .A2(new_n444_), .B(new_n4572_), .ZN(\grant[68] ));
  NOR2_X1    g4188(.A1(new_n1052_), .A2(new_n670_), .ZN(new_n4574_));
  OAI21_X1   g4189(.A1(new_n438_), .A2(new_n4574_), .B(new_n676_), .ZN(new_n4575_));
  AOI21_X1   g4190(.A1(new_n4575_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n4576_));
  OAI21_X1   g4191(.A1(new_n4576_), .A2(new_n687_), .B(new_n692_), .ZN(new_n4577_));
  AOI21_X1   g4192(.A1(new_n4577_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n4578_));
  OAI21_X1   g4193(.A1(new_n4578_), .A2(new_n425_), .B(new_n703_), .ZN(new_n4579_));
  AOI21_X1   g4194(.A1(new_n4579_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n4580_));
  OAI21_X1   g4195(.A1(new_n4580_), .A2(new_n420_), .B(new_n718_), .ZN(new_n4581_));
  AOI21_X1   g4196(.A1(new_n4581_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n4582_));
  OAI21_X1   g4197(.A1(new_n4582_), .A2(new_n729_), .B(new_n734_), .ZN(new_n4583_));
  AOI21_X1   g4198(.A1(new_n4583_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n4584_));
  OAI21_X1   g4199(.A1(new_n4584_), .A2(new_n407_), .B(new_n745_), .ZN(new_n4585_));
  AOI21_X1   g4200(.A1(new_n4585_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n4586_));
  OAI21_X1   g4201(.A1(new_n4586_), .A2(new_n402_), .B(new_n760_), .ZN(new_n4587_));
  AOI21_X1   g4202(.A1(new_n4587_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n4588_));
  OAI21_X1   g4203(.A1(new_n4588_), .A2(new_n771_), .B(new_n776_), .ZN(new_n4589_));
  AOI21_X1   g4204(.A1(new_n4589_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n4590_));
  OAI21_X1   g4205(.A1(new_n4590_), .A2(new_n389_), .B(new_n787_), .ZN(new_n4591_));
  AOI21_X1   g4206(.A1(new_n4591_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n4592_));
  OAI21_X1   g4207(.A1(new_n4592_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n4593_));
  AOI21_X1   g4208(.A1(new_n4593_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n4594_));
  OAI21_X1   g4209(.A1(new_n4594_), .A2(new_n900_), .B(new_n908_), .ZN(new_n4595_));
  AOI21_X1   g4210(.A1(new_n4595_), .A2(new_n913_), .B(new_n918_), .ZN(new_n4596_));
  OAI21_X1   g4211(.A1(new_n4596_), .A2(new_n897_), .B(new_n923_), .ZN(new_n4597_));
  AOI21_X1   g4212(.A1(new_n4597_), .A2(new_n894_), .B(new_n929_), .ZN(new_n4598_));
  OAI21_X1   g4213(.A1(new_n4598_), .A2(new_n933_), .B(new_n937_), .ZN(new_n4599_));
  AOI21_X1   g4214(.A1(new_n4599_), .A2(new_n890_), .B(new_n943_), .ZN(new_n4600_));
  OAI21_X1   g4215(.A1(new_n4600_), .A2(new_n886_), .B(new_n948_), .ZN(new_n4601_));
  AOI21_X1   g4216(.A1(new_n4601_), .A2(new_n953_), .B(new_n958_), .ZN(new_n4602_));
  OAI21_X1   g4217(.A1(new_n4602_), .A2(new_n883_), .B(new_n963_), .ZN(new_n4603_));
  AOI21_X1   g4218(.A1(new_n4603_), .A2(new_n880_), .B(new_n969_), .ZN(new_n4604_));
  OAI21_X1   g4219(.A1(new_n4604_), .A2(new_n973_), .B(new_n977_), .ZN(new_n4605_));
  AOI21_X1   g4220(.A1(new_n4605_), .A2(new_n876_), .B(new_n983_), .ZN(new_n4606_));
  OAI21_X1   g4221(.A1(new_n4606_), .A2(new_n872_), .B(new_n988_), .ZN(new_n4607_));
  AOI21_X1   g4222(.A1(new_n4607_), .A2(new_n993_), .B(new_n998_), .ZN(new_n4608_));
  OAI21_X1   g4223(.A1(new_n4608_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n4609_));
  AOI21_X1   g4224(.A1(new_n4609_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n4610_));
  OAI21_X1   g4225(.A1(new_n4610_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n4611_));
  AOI21_X1   g4226(.A1(new_n4611_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n4612_));
  OAI21_X1   g4227(.A1(new_n4612_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n4613_));
  AOI21_X1   g4228(.A1(new_n4613_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n4614_));
  OAI21_X1   g4229(.A1(new_n4614_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n4615_));
  OAI21_X1   g4230(.A1(new_n1045_), .A2(\priority[69] ), .B(\req[69] ), .ZN(new_n4616_));
  AOI21_X1   g4231(.A1(new_n4615_), .A2(new_n852_), .B(new_n4616_), .ZN(\grant[69] ));
  NOR2_X1    g4232(.A1(new_n1411_), .A2(new_n1056_), .ZN(new_n4618_));
  OAI21_X1   g4233(.A1(new_n847_), .A2(new_n4618_), .B(new_n1062_), .ZN(new_n4619_));
  AOI21_X1   g4234(.A1(new_n4619_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n4620_));
  OAI21_X1   g4235(.A1(new_n4620_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n4621_));
  AOI21_X1   g4236(.A1(new_n4621_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n4622_));
  OAI21_X1   g4237(.A1(new_n4622_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n4623_));
  AOI21_X1   g4238(.A1(new_n4623_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n4624_));
  OAI21_X1   g4239(.A1(new_n4624_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n4625_));
  AOI21_X1   g4240(.A1(new_n4625_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n4626_));
  OAI21_X1   g4241(.A1(new_n4626_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n4627_));
  AOI21_X1   g4242(.A1(new_n4627_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n4628_));
  OAI21_X1   g4243(.A1(new_n4628_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n4629_));
  AOI21_X1   g4244(.A1(new_n4629_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n4630_));
  OAI21_X1   g4245(.A1(new_n4630_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n4631_));
  AOI21_X1   g4246(.A1(new_n4631_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n4632_));
  OAI21_X1   g4247(.A1(new_n4632_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n4633_));
  AOI21_X1   g4248(.A1(new_n4633_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n4634_));
  OAI21_X1   g4249(.A1(new_n4634_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n4635_));
  AOI21_X1   g4250(.A1(new_n4635_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n4636_));
  OAI21_X1   g4251(.A1(new_n4636_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n4637_));
  AOI21_X1   g4252(.A1(new_n4637_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n4638_));
  OAI21_X1   g4253(.A1(new_n4638_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n4639_));
  AOI21_X1   g4254(.A1(new_n4639_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n4640_));
  OAI21_X1   g4255(.A1(new_n4640_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n4641_));
  AOI21_X1   g4256(.A1(new_n4641_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n4642_));
  OAI21_X1   g4257(.A1(new_n4642_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n4643_));
  AOI21_X1   g4258(.A1(new_n4643_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n4644_));
  OAI21_X1   g4259(.A1(new_n4644_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n4645_));
  AOI21_X1   g4260(.A1(new_n4645_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n4646_));
  OAI21_X1   g4261(.A1(new_n4646_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n4647_));
  AOI21_X1   g4262(.A1(new_n4647_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n4648_));
  OAI21_X1   g4263(.A1(new_n4648_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n4649_));
  AOI21_X1   g4264(.A1(new_n4649_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n4650_));
  OAI21_X1   g4265(.A1(new_n4650_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n4651_));
  AOI21_X1   g4266(.A1(new_n4651_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n4652_));
  OAI21_X1   g4267(.A1(new_n4652_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n4653_));
  AOI21_X1   g4268(.A1(new_n4653_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n4654_));
  OAI21_X1   g4269(.A1(new_n4654_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n4655_));
  AOI21_X1   g4270(.A1(new_n4655_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n4656_));
  OAI21_X1   g4271(.A1(new_n4656_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n4657_));
  AOI21_X1   g4272(.A1(new_n4657_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n4658_));
  OAI21_X1   g4273(.A1(new_n4658_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n4659_));
  OAI21_X1   g4274(.A1(new_n665_), .A2(\priority[70] ), .B(\req[70] ), .ZN(new_n4660_));
  AOI21_X1   g4275(.A1(new_n4659_), .A2(new_n1235_), .B(new_n4660_), .ZN(\grant[70] ));
  NOR2_X1    g4276(.A1(new_n437_), .A2(new_n1414_), .ZN(new_n4662_));
  OAI21_X1   g4277(.A1(new_n1230_), .A2(new_n4662_), .B(new_n1419_), .ZN(new_n4663_));
  AOI21_X1   g4278(.A1(new_n4663_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n4664_));
  OAI21_X1   g4279(.A1(new_n4664_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n4665_));
  AOI21_X1   g4280(.A1(new_n4665_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n4666_));
  OAI21_X1   g4281(.A1(new_n4666_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n4667_));
  AOI21_X1   g4282(.A1(new_n4667_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n4668_));
  OAI21_X1   g4283(.A1(new_n4668_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n4669_));
  AOI21_X1   g4284(.A1(new_n4669_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n4670_));
  OAI21_X1   g4285(.A1(new_n4670_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n4671_));
  AOI21_X1   g4286(.A1(new_n4671_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n4672_));
  OAI21_X1   g4287(.A1(new_n4672_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n4673_));
  AOI21_X1   g4288(.A1(new_n4673_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n4674_));
  OAI21_X1   g4289(.A1(new_n4674_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n4675_));
  AOI21_X1   g4290(.A1(new_n4675_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n4676_));
  OAI21_X1   g4291(.A1(new_n4676_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n4677_));
  AOI21_X1   g4292(.A1(new_n4677_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n4678_));
  OAI21_X1   g4293(.A1(new_n4678_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n4679_));
  AOI21_X1   g4294(.A1(new_n4679_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n4680_));
  OAI21_X1   g4295(.A1(new_n4680_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n4681_));
  AOI21_X1   g4296(.A1(new_n4681_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n4682_));
  OAI21_X1   g4297(.A1(new_n4682_), .A2(new_n519_), .B(new_n524_), .ZN(new_n4683_));
  AOI21_X1   g4298(.A1(new_n4683_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n4684_));
  OAI21_X1   g4299(.A1(new_n4684_), .A2(new_n497_), .B(new_n535_), .ZN(new_n4685_));
  AOI21_X1   g4300(.A1(new_n4685_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n4686_));
  OAI21_X1   g4301(.A1(new_n4686_), .A2(new_n492_), .B(new_n550_), .ZN(new_n4687_));
  AOI21_X1   g4302(.A1(new_n4687_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n4688_));
  OAI21_X1   g4303(.A1(new_n4688_), .A2(new_n561_), .B(new_n566_), .ZN(new_n4689_));
  AOI21_X1   g4304(.A1(new_n4689_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n4690_));
  OAI21_X1   g4305(.A1(new_n4690_), .A2(new_n479_), .B(new_n577_), .ZN(new_n4691_));
  AOI21_X1   g4306(.A1(new_n4691_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n4692_));
  OAI21_X1   g4307(.A1(new_n4692_), .A2(new_n474_), .B(new_n592_), .ZN(new_n4693_));
  AOI21_X1   g4308(.A1(new_n4693_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n4694_));
  OAI21_X1   g4309(.A1(new_n4694_), .A2(new_n603_), .B(new_n608_), .ZN(new_n4695_));
  AOI21_X1   g4310(.A1(new_n4695_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n4696_));
  OAI21_X1   g4311(.A1(new_n4696_), .A2(new_n461_), .B(new_n619_), .ZN(new_n4697_));
  AOI21_X1   g4312(.A1(new_n4697_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n4698_));
  OAI21_X1   g4313(.A1(new_n4698_), .A2(new_n456_), .B(new_n634_), .ZN(new_n4699_));
  AOI21_X1   g4314(.A1(new_n4699_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n4700_));
  OAI21_X1   g4315(.A1(new_n4700_), .A2(new_n645_), .B(new_n650_), .ZN(new_n4701_));
  AOI21_X1   g4316(.A1(new_n4701_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n4702_));
  OAI21_X1   g4317(.A1(new_n4702_), .A2(new_n443_), .B(new_n661_), .ZN(new_n4703_));
  OAI21_X1   g4318(.A1(new_n668_), .A2(\priority[71] ), .B(\req[71] ), .ZN(new_n4704_));
  AOI21_X1   g4319(.A1(new_n4703_), .A2(new_n1542_), .B(new_n4704_), .ZN(\grant[71] ));
  NOR2_X1    g4320(.A1(new_n846_), .A2(new_n675_), .ZN(new_n4706_));
  OAI21_X1   g4321(.A1(new_n434_), .A2(new_n4706_), .B(new_n682_), .ZN(new_n4707_));
  AOI21_X1   g4322(.A1(new_n4707_), .A2(new_n688_), .B(new_n693_), .ZN(new_n4708_));
  OAI21_X1   g4323(.A1(new_n4708_), .A2(new_n430_), .B(new_n698_), .ZN(new_n4709_));
  AOI21_X1   g4324(.A1(new_n4709_), .A2(new_n426_), .B(new_n704_), .ZN(new_n4710_));
  OAI21_X1   g4325(.A1(new_n4710_), .A2(new_n709_), .B(new_n713_), .ZN(new_n4711_));
  AOI21_X1   g4326(.A1(new_n4711_), .A2(new_n421_), .B(new_n719_), .ZN(new_n4712_));
  OAI21_X1   g4327(.A1(new_n4712_), .A2(new_n416_), .B(new_n724_), .ZN(new_n4713_));
  AOI21_X1   g4328(.A1(new_n4713_), .A2(new_n730_), .B(new_n735_), .ZN(new_n4714_));
  OAI21_X1   g4329(.A1(new_n4714_), .A2(new_n412_), .B(new_n740_), .ZN(new_n4715_));
  AOI21_X1   g4330(.A1(new_n4715_), .A2(new_n408_), .B(new_n746_), .ZN(new_n4716_));
  OAI21_X1   g4331(.A1(new_n4716_), .A2(new_n751_), .B(new_n755_), .ZN(new_n4717_));
  AOI21_X1   g4332(.A1(new_n4717_), .A2(new_n403_), .B(new_n761_), .ZN(new_n4718_));
  OAI21_X1   g4333(.A1(new_n4718_), .A2(new_n398_), .B(new_n766_), .ZN(new_n4719_));
  AOI21_X1   g4334(.A1(new_n4719_), .A2(new_n772_), .B(new_n777_), .ZN(new_n4720_));
  OAI21_X1   g4335(.A1(new_n4720_), .A2(new_n394_), .B(new_n782_), .ZN(new_n4721_));
  AOI21_X1   g4336(.A1(new_n4721_), .A2(new_n390_), .B(new_n788_), .ZN(new_n4722_));
  OAI21_X1   g4337(.A1(new_n4722_), .A2(new_n793_), .B(new_n797_), .ZN(new_n4723_));
  AOI21_X1   g4338(.A1(new_n4723_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n4724_));
  OAI21_X1   g4339(.A1(new_n4724_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n4725_));
  AOI21_X1   g4340(.A1(new_n4725_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n4726_));
  OAI21_X1   g4341(.A1(new_n4726_), .A2(new_n912_), .B(new_n917_), .ZN(new_n4727_));
  AOI21_X1   g4342(.A1(new_n4727_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n4728_));
  OAI21_X1   g4343(.A1(new_n4728_), .A2(new_n893_), .B(new_n928_), .ZN(new_n4729_));
  AOI21_X1   g4344(.A1(new_n4729_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n4730_));
  OAI21_X1   g4345(.A1(new_n4730_), .A2(new_n889_), .B(new_n942_), .ZN(new_n4731_));
  AOI21_X1   g4346(.A1(new_n4731_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n4732_));
  OAI21_X1   g4347(.A1(new_n4732_), .A2(new_n952_), .B(new_n957_), .ZN(new_n4733_));
  AOI21_X1   g4348(.A1(new_n4733_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n4734_));
  OAI21_X1   g4349(.A1(new_n4734_), .A2(new_n879_), .B(new_n968_), .ZN(new_n4735_));
  AOI21_X1   g4350(.A1(new_n4735_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n4736_));
  OAI21_X1   g4351(.A1(new_n4736_), .A2(new_n875_), .B(new_n982_), .ZN(new_n4737_));
  AOI21_X1   g4352(.A1(new_n4737_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n4738_));
  OAI21_X1   g4353(.A1(new_n4738_), .A2(new_n992_), .B(new_n997_), .ZN(new_n4739_));
  AOI21_X1   g4354(.A1(new_n4739_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n4740_));
  OAI21_X1   g4355(.A1(new_n4740_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n4741_));
  AOI21_X1   g4356(.A1(new_n4741_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n4742_));
  OAI21_X1   g4357(.A1(new_n4742_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n4743_));
  AOI21_X1   g4358(.A1(new_n4743_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n4744_));
  OAI21_X1   g4359(.A1(new_n4744_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n4745_));
  AOI21_X1   g4360(.A1(new_n4745_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n4746_));
  OAI21_X1   g4361(.A1(new_n4746_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n4747_));
  OAI21_X1   g4362(.A1(new_n1054_), .A2(\priority[72] ), .B(\req[72] ), .ZN(new_n4748_));
  AOI21_X1   g4363(.A1(new_n4747_), .A2(new_n1632_), .B(new_n4748_), .ZN(\grant[72] ));
  NOR2_X1    g4364(.A1(new_n1229_), .A2(new_n1061_), .ZN(new_n4750_));
  OAI21_X1   g4365(.A1(new_n844_), .A2(new_n4750_), .B(new_n1068_), .ZN(new_n4751_));
  AOI21_X1   g4366(.A1(new_n4751_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n4752_));
  OAI21_X1   g4367(.A1(new_n4752_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n4753_));
  AOI21_X1   g4368(.A1(new_n4753_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n4754_));
  OAI21_X1   g4369(.A1(new_n4754_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n4755_));
  AOI21_X1   g4370(.A1(new_n4755_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n4756_));
  OAI21_X1   g4371(.A1(new_n4756_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n4757_));
  AOI21_X1   g4372(.A1(new_n4757_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n4758_));
  OAI21_X1   g4373(.A1(new_n4758_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n4759_));
  AOI21_X1   g4374(.A1(new_n4759_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n4760_));
  OAI21_X1   g4375(.A1(new_n4760_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n4761_));
  AOI21_X1   g4376(.A1(new_n4761_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n4762_));
  OAI21_X1   g4377(.A1(new_n4762_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n4763_));
  AOI21_X1   g4378(.A1(new_n4763_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n4764_));
  OAI21_X1   g4379(.A1(new_n4764_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n4765_));
  AOI21_X1   g4380(.A1(new_n4765_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n4766_));
  OAI21_X1   g4381(.A1(new_n4766_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n4767_));
  AOI21_X1   g4382(.A1(new_n4767_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n4768_));
  OAI21_X1   g4383(.A1(new_n4768_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n4769_));
  AOI21_X1   g4384(.A1(new_n4769_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n4770_));
  OAI21_X1   g4385(.A1(new_n4770_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n4771_));
  AOI21_X1   g4386(.A1(new_n4771_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n4772_));
  OAI21_X1   g4387(.A1(new_n4772_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n4773_));
  AOI21_X1   g4388(.A1(new_n4773_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n4774_));
  OAI21_X1   g4389(.A1(new_n4774_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n4775_));
  AOI21_X1   g4390(.A1(new_n4775_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n4776_));
  OAI21_X1   g4391(.A1(new_n4776_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n4777_));
  AOI21_X1   g4392(.A1(new_n4777_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n4778_));
  OAI21_X1   g4393(.A1(new_n4778_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n4779_));
  AOI21_X1   g4394(.A1(new_n4779_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n4780_));
  OAI21_X1   g4395(.A1(new_n4780_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n4781_));
  AOI21_X1   g4396(.A1(new_n4781_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n4782_));
  OAI21_X1   g4397(.A1(new_n4782_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n4783_));
  AOI21_X1   g4398(.A1(new_n4783_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n4784_));
  OAI21_X1   g4399(.A1(new_n4784_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n4785_));
  AOI21_X1   g4400(.A1(new_n4785_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n4786_));
  OAI21_X1   g4401(.A1(new_n4786_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n4787_));
  AOI21_X1   g4402(.A1(new_n4787_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n4788_));
  OAI21_X1   g4403(.A1(new_n4788_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n4789_));
  AOI21_X1   g4404(.A1(new_n4789_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n4790_));
  OAI21_X1   g4405(.A1(new_n4790_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n4791_));
  OAI21_X1   g4406(.A1(new_n436_), .A2(\priority[73] ), .B(\req[73] ), .ZN(new_n4792_));
  AOI21_X1   g4407(.A1(new_n4791_), .A2(new_n1720_), .B(new_n4792_), .ZN(\grant[73] ));
  NOR2_X1    g4408(.A1(new_n433_), .A2(new_n1418_), .ZN(new_n4794_));
  OAI21_X1   g4409(.A1(new_n1227_), .A2(new_n4794_), .B(new_n1424_), .ZN(new_n4795_));
  AOI21_X1   g4410(.A1(new_n4795_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n4796_));
  OAI21_X1   g4411(.A1(new_n4796_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n4797_));
  AOI21_X1   g4412(.A1(new_n4797_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n4798_));
  OAI21_X1   g4413(.A1(new_n4798_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n4799_));
  AOI21_X1   g4414(.A1(new_n4799_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n4800_));
  OAI21_X1   g4415(.A1(new_n4800_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n4801_));
  AOI21_X1   g4416(.A1(new_n4801_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n4802_));
  OAI21_X1   g4417(.A1(new_n4802_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n4803_));
  AOI21_X1   g4418(.A1(new_n4803_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n4804_));
  OAI21_X1   g4419(.A1(new_n4804_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n4805_));
  AOI21_X1   g4420(.A1(new_n4805_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n4806_));
  OAI21_X1   g4421(.A1(new_n4806_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n4807_));
  AOI21_X1   g4422(.A1(new_n4807_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n4808_));
  OAI21_X1   g4423(.A1(new_n4808_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n4809_));
  AOI21_X1   g4424(.A1(new_n4809_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n4810_));
  OAI21_X1   g4425(.A1(new_n4810_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n4811_));
  AOI21_X1   g4426(.A1(new_n4811_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n4812_));
  OAI21_X1   g4427(.A1(new_n4812_), .A2(new_n506_), .B(new_n514_), .ZN(new_n4813_));
  AOI21_X1   g4428(.A1(new_n4813_), .A2(new_n520_), .B(new_n525_), .ZN(new_n4814_));
  OAI21_X1   g4429(.A1(new_n4814_), .A2(new_n502_), .B(new_n530_), .ZN(new_n4815_));
  AOI21_X1   g4430(.A1(new_n4815_), .A2(new_n498_), .B(new_n536_), .ZN(new_n4816_));
  OAI21_X1   g4431(.A1(new_n4816_), .A2(new_n541_), .B(new_n545_), .ZN(new_n4817_));
  AOI21_X1   g4432(.A1(new_n4817_), .A2(new_n493_), .B(new_n551_), .ZN(new_n4818_));
  OAI21_X1   g4433(.A1(new_n4818_), .A2(new_n488_), .B(new_n556_), .ZN(new_n4819_));
  AOI21_X1   g4434(.A1(new_n4819_), .A2(new_n562_), .B(new_n567_), .ZN(new_n4820_));
  OAI21_X1   g4435(.A1(new_n4820_), .A2(new_n484_), .B(new_n572_), .ZN(new_n4821_));
  AOI21_X1   g4436(.A1(new_n4821_), .A2(new_n480_), .B(new_n578_), .ZN(new_n4822_));
  OAI21_X1   g4437(.A1(new_n4822_), .A2(new_n583_), .B(new_n587_), .ZN(new_n4823_));
  AOI21_X1   g4438(.A1(new_n4823_), .A2(new_n475_), .B(new_n593_), .ZN(new_n4824_));
  OAI21_X1   g4439(.A1(new_n4824_), .A2(new_n470_), .B(new_n598_), .ZN(new_n4825_));
  AOI21_X1   g4440(.A1(new_n4825_), .A2(new_n604_), .B(new_n609_), .ZN(new_n4826_));
  OAI21_X1   g4441(.A1(new_n4826_), .A2(new_n466_), .B(new_n614_), .ZN(new_n4827_));
  AOI21_X1   g4442(.A1(new_n4827_), .A2(new_n462_), .B(new_n620_), .ZN(new_n4828_));
  OAI21_X1   g4443(.A1(new_n4828_), .A2(new_n625_), .B(new_n629_), .ZN(new_n4829_));
  AOI21_X1   g4444(.A1(new_n4829_), .A2(new_n457_), .B(new_n635_), .ZN(new_n4830_));
  OAI21_X1   g4445(.A1(new_n4830_), .A2(new_n452_), .B(new_n640_), .ZN(new_n4831_));
  AOI21_X1   g4446(.A1(new_n4831_), .A2(new_n646_), .B(new_n651_), .ZN(new_n4832_));
  OAI21_X1   g4447(.A1(new_n4832_), .A2(new_n448_), .B(new_n656_), .ZN(new_n4833_));
  AOI21_X1   g4448(.A1(new_n4833_), .A2(new_n444_), .B(new_n662_), .ZN(new_n4834_));
  OAI21_X1   g4449(.A1(new_n4834_), .A2(new_n667_), .B(new_n671_), .ZN(new_n4835_));
  OAI21_X1   g4450(.A1(new_n673_), .A2(\priority[74] ), .B(\req[74] ), .ZN(new_n4836_));
  AOI21_X1   g4451(.A1(new_n4835_), .A2(new_n439_), .B(new_n4836_), .ZN(\grant[74] ));
  NOR2_X1    g4452(.A1(new_n843_), .A2(new_n681_), .ZN(new_n4838_));
  OAI21_X1   g4453(.A1(new_n687_), .A2(new_n4838_), .B(new_n692_), .ZN(new_n4839_));
  AOI21_X1   g4454(.A1(new_n4839_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n4840_));
  OAI21_X1   g4455(.A1(new_n4840_), .A2(new_n425_), .B(new_n703_), .ZN(new_n4841_));
  AOI21_X1   g4456(.A1(new_n4841_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n4842_));
  OAI21_X1   g4457(.A1(new_n4842_), .A2(new_n420_), .B(new_n718_), .ZN(new_n4843_));
  AOI21_X1   g4458(.A1(new_n4843_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n4844_));
  OAI21_X1   g4459(.A1(new_n4844_), .A2(new_n729_), .B(new_n734_), .ZN(new_n4845_));
  AOI21_X1   g4460(.A1(new_n4845_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n4846_));
  OAI21_X1   g4461(.A1(new_n4846_), .A2(new_n407_), .B(new_n745_), .ZN(new_n4847_));
  AOI21_X1   g4462(.A1(new_n4847_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n4848_));
  OAI21_X1   g4463(.A1(new_n4848_), .A2(new_n402_), .B(new_n760_), .ZN(new_n4849_));
  AOI21_X1   g4464(.A1(new_n4849_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n4850_));
  OAI21_X1   g4465(.A1(new_n4850_), .A2(new_n771_), .B(new_n776_), .ZN(new_n4851_));
  AOI21_X1   g4466(.A1(new_n4851_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n4852_));
  OAI21_X1   g4467(.A1(new_n4852_), .A2(new_n389_), .B(new_n787_), .ZN(new_n4853_));
  AOI21_X1   g4468(.A1(new_n4853_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n4854_));
  OAI21_X1   g4469(.A1(new_n4854_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n4855_));
  AOI21_X1   g4470(.A1(new_n4855_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n4856_));
  OAI21_X1   g4471(.A1(new_n4856_), .A2(new_n900_), .B(new_n908_), .ZN(new_n4857_));
  AOI21_X1   g4472(.A1(new_n4857_), .A2(new_n913_), .B(new_n918_), .ZN(new_n4858_));
  OAI21_X1   g4473(.A1(new_n4858_), .A2(new_n897_), .B(new_n923_), .ZN(new_n4859_));
  AOI21_X1   g4474(.A1(new_n4859_), .A2(new_n894_), .B(new_n929_), .ZN(new_n4860_));
  OAI21_X1   g4475(.A1(new_n4860_), .A2(new_n933_), .B(new_n937_), .ZN(new_n4861_));
  AOI21_X1   g4476(.A1(new_n4861_), .A2(new_n890_), .B(new_n943_), .ZN(new_n4862_));
  OAI21_X1   g4477(.A1(new_n4862_), .A2(new_n886_), .B(new_n948_), .ZN(new_n4863_));
  AOI21_X1   g4478(.A1(new_n4863_), .A2(new_n953_), .B(new_n958_), .ZN(new_n4864_));
  OAI21_X1   g4479(.A1(new_n4864_), .A2(new_n883_), .B(new_n963_), .ZN(new_n4865_));
  AOI21_X1   g4480(.A1(new_n4865_), .A2(new_n880_), .B(new_n969_), .ZN(new_n4866_));
  OAI21_X1   g4481(.A1(new_n4866_), .A2(new_n973_), .B(new_n977_), .ZN(new_n4867_));
  AOI21_X1   g4482(.A1(new_n4867_), .A2(new_n876_), .B(new_n983_), .ZN(new_n4868_));
  OAI21_X1   g4483(.A1(new_n4868_), .A2(new_n872_), .B(new_n988_), .ZN(new_n4869_));
  AOI21_X1   g4484(.A1(new_n4869_), .A2(new_n993_), .B(new_n998_), .ZN(new_n4870_));
  OAI21_X1   g4485(.A1(new_n4870_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n4871_));
  AOI21_X1   g4486(.A1(new_n4871_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n4872_));
  OAI21_X1   g4487(.A1(new_n4872_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n4873_));
  AOI21_X1   g4488(.A1(new_n4873_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n4874_));
  OAI21_X1   g4489(.A1(new_n4874_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n4875_));
  AOI21_X1   g4490(.A1(new_n4875_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n4876_));
  OAI21_X1   g4491(.A1(new_n4876_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n4877_));
  AOI21_X1   g4492(.A1(new_n4877_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n4878_));
  OAI21_X1   g4493(.A1(new_n4878_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n4879_));
  OAI21_X1   g4494(.A1(new_n1059_), .A2(\priority[75] ), .B(\req[75] ), .ZN(new_n4880_));
  AOI21_X1   g4495(.A1(new_n4879_), .A2(new_n848_), .B(new_n4880_), .ZN(\grant[75] ));
  NOR2_X1    g4496(.A1(new_n1226_), .A2(new_n1067_), .ZN(new_n4882_));
  OAI21_X1   g4497(.A1(new_n1072_), .A2(new_n4882_), .B(new_n1077_), .ZN(new_n4883_));
  AOI21_X1   g4498(.A1(new_n4883_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n4884_));
  OAI21_X1   g4499(.A1(new_n4884_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n4885_));
  AOI21_X1   g4500(.A1(new_n4885_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n4886_));
  OAI21_X1   g4501(.A1(new_n4886_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n4887_));
  AOI21_X1   g4502(.A1(new_n4887_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n4888_));
  OAI21_X1   g4503(.A1(new_n4888_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n4889_));
  AOI21_X1   g4504(.A1(new_n4889_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n4890_));
  OAI21_X1   g4505(.A1(new_n4890_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n4891_));
  AOI21_X1   g4506(.A1(new_n4891_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n4892_));
  OAI21_X1   g4507(.A1(new_n4892_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n4893_));
  AOI21_X1   g4508(.A1(new_n4893_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n4894_));
  OAI21_X1   g4509(.A1(new_n4894_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n4895_));
  AOI21_X1   g4510(.A1(new_n4895_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n4896_));
  OAI21_X1   g4511(.A1(new_n4896_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n4897_));
  AOI21_X1   g4512(.A1(new_n4897_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n4898_));
  OAI21_X1   g4513(.A1(new_n4898_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n4899_));
  AOI21_X1   g4514(.A1(new_n4899_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n4900_));
  OAI21_X1   g4515(.A1(new_n4900_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n4901_));
  AOI21_X1   g4516(.A1(new_n4901_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n4902_));
  OAI21_X1   g4517(.A1(new_n4902_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n4903_));
  AOI21_X1   g4518(.A1(new_n4903_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n4904_));
  OAI21_X1   g4519(.A1(new_n4904_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n4905_));
  AOI21_X1   g4520(.A1(new_n4905_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n4906_));
  OAI21_X1   g4521(.A1(new_n4906_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n4907_));
  AOI21_X1   g4522(.A1(new_n4907_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n4908_));
  OAI21_X1   g4523(.A1(new_n4908_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n4909_));
  AOI21_X1   g4524(.A1(new_n4909_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n4910_));
  OAI21_X1   g4525(.A1(new_n4910_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n4911_));
  AOI21_X1   g4526(.A1(new_n4911_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n4912_));
  OAI21_X1   g4527(.A1(new_n4912_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n4913_));
  AOI21_X1   g4528(.A1(new_n4913_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n4914_));
  OAI21_X1   g4529(.A1(new_n4914_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n4915_));
  AOI21_X1   g4530(.A1(new_n4915_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n4916_));
  OAI21_X1   g4531(.A1(new_n4916_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n4917_));
  AOI21_X1   g4532(.A1(new_n4917_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n4918_));
  OAI21_X1   g4533(.A1(new_n4918_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n4919_));
  AOI21_X1   g4534(.A1(new_n4919_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n4920_));
  OAI21_X1   g4535(.A1(new_n4920_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n4921_));
  AOI21_X1   g4536(.A1(new_n4921_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n4922_));
  OAI21_X1   g4537(.A1(new_n4922_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n4923_));
  OAI21_X1   g4538(.A1(new_n432_), .A2(\priority[76] ), .B(\req[76] ), .ZN(new_n4924_));
  AOI21_X1   g4539(.A1(new_n4923_), .A2(new_n1231_), .B(new_n4924_), .ZN(\grant[76] ));
  NOR2_X1    g4540(.A1(new_n686_), .A2(new_n1423_), .ZN(new_n4926_));
  OAI21_X1   g4541(.A1(new_n1428_), .A2(new_n4926_), .B(new_n1432_), .ZN(new_n4927_));
  AOI21_X1   g4542(.A1(new_n4927_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n4928_));
  OAI21_X1   g4543(.A1(new_n4928_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n4929_));
  AOI21_X1   g4544(.A1(new_n4929_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n4930_));
  OAI21_X1   g4545(.A1(new_n4930_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n4931_));
  AOI21_X1   g4546(.A1(new_n4931_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n4932_));
  OAI21_X1   g4547(.A1(new_n4932_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n4933_));
  AOI21_X1   g4548(.A1(new_n4933_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n4934_));
  OAI21_X1   g4549(.A1(new_n4934_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n4935_));
  AOI21_X1   g4550(.A1(new_n4935_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n4936_));
  OAI21_X1   g4551(.A1(new_n4936_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n4937_));
  AOI21_X1   g4552(.A1(new_n4937_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n4938_));
  OAI21_X1   g4553(.A1(new_n4938_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n4939_));
  AOI21_X1   g4554(.A1(new_n4939_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n4940_));
  OAI21_X1   g4555(.A1(new_n4940_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n4941_));
  AOI21_X1   g4556(.A1(new_n4941_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n4942_));
  OAI21_X1   g4557(.A1(new_n4942_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n4943_));
  AOI21_X1   g4558(.A1(new_n4943_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n4944_));
  OAI21_X1   g4559(.A1(new_n4944_), .A2(new_n519_), .B(new_n524_), .ZN(new_n4945_));
  AOI21_X1   g4560(.A1(new_n4945_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n4946_));
  OAI21_X1   g4561(.A1(new_n4946_), .A2(new_n497_), .B(new_n535_), .ZN(new_n4947_));
  AOI21_X1   g4562(.A1(new_n4947_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n4948_));
  OAI21_X1   g4563(.A1(new_n4948_), .A2(new_n492_), .B(new_n550_), .ZN(new_n4949_));
  AOI21_X1   g4564(.A1(new_n4949_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n4950_));
  OAI21_X1   g4565(.A1(new_n4950_), .A2(new_n561_), .B(new_n566_), .ZN(new_n4951_));
  AOI21_X1   g4566(.A1(new_n4951_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n4952_));
  OAI21_X1   g4567(.A1(new_n4952_), .A2(new_n479_), .B(new_n577_), .ZN(new_n4953_));
  AOI21_X1   g4568(.A1(new_n4953_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n4954_));
  OAI21_X1   g4569(.A1(new_n4954_), .A2(new_n474_), .B(new_n592_), .ZN(new_n4955_));
  AOI21_X1   g4570(.A1(new_n4955_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n4956_));
  OAI21_X1   g4571(.A1(new_n4956_), .A2(new_n603_), .B(new_n608_), .ZN(new_n4957_));
  AOI21_X1   g4572(.A1(new_n4957_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n4958_));
  OAI21_X1   g4573(.A1(new_n4958_), .A2(new_n461_), .B(new_n619_), .ZN(new_n4959_));
  AOI21_X1   g4574(.A1(new_n4959_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n4960_));
  OAI21_X1   g4575(.A1(new_n4960_), .A2(new_n456_), .B(new_n634_), .ZN(new_n4961_));
  AOI21_X1   g4576(.A1(new_n4961_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n4962_));
  OAI21_X1   g4577(.A1(new_n4962_), .A2(new_n645_), .B(new_n650_), .ZN(new_n4963_));
  AOI21_X1   g4578(.A1(new_n4963_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n4964_));
  OAI21_X1   g4579(.A1(new_n4964_), .A2(new_n443_), .B(new_n661_), .ZN(new_n4965_));
  AOI21_X1   g4580(.A1(new_n4965_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n4966_));
  OAI21_X1   g4581(.A1(new_n4966_), .A2(new_n438_), .B(new_n676_), .ZN(new_n4967_));
  OAI21_X1   g4582(.A1(new_n679_), .A2(\priority[77] ), .B(\req[77] ), .ZN(new_n4968_));
  AOI21_X1   g4583(.A1(new_n4967_), .A2(new_n1540_), .B(new_n4968_), .ZN(\grant[77] ));
  NOR2_X1    g4584(.A1(new_n1071_), .A2(new_n691_), .ZN(new_n4970_));
  OAI21_X1   g4585(.A1(new_n430_), .A2(new_n4970_), .B(new_n698_), .ZN(new_n4971_));
  AOI21_X1   g4586(.A1(new_n4971_), .A2(new_n426_), .B(new_n704_), .ZN(new_n4972_));
  OAI21_X1   g4587(.A1(new_n4972_), .A2(new_n709_), .B(new_n713_), .ZN(new_n4973_));
  AOI21_X1   g4588(.A1(new_n4973_), .A2(new_n421_), .B(new_n719_), .ZN(new_n4974_));
  OAI21_X1   g4589(.A1(new_n4974_), .A2(new_n416_), .B(new_n724_), .ZN(new_n4975_));
  AOI21_X1   g4590(.A1(new_n4975_), .A2(new_n730_), .B(new_n735_), .ZN(new_n4976_));
  OAI21_X1   g4591(.A1(new_n4976_), .A2(new_n412_), .B(new_n740_), .ZN(new_n4977_));
  AOI21_X1   g4592(.A1(new_n4977_), .A2(new_n408_), .B(new_n746_), .ZN(new_n4978_));
  OAI21_X1   g4593(.A1(new_n4978_), .A2(new_n751_), .B(new_n755_), .ZN(new_n4979_));
  AOI21_X1   g4594(.A1(new_n4979_), .A2(new_n403_), .B(new_n761_), .ZN(new_n4980_));
  OAI21_X1   g4595(.A1(new_n4980_), .A2(new_n398_), .B(new_n766_), .ZN(new_n4981_));
  AOI21_X1   g4596(.A1(new_n4981_), .A2(new_n772_), .B(new_n777_), .ZN(new_n4982_));
  OAI21_X1   g4597(.A1(new_n4982_), .A2(new_n394_), .B(new_n782_), .ZN(new_n4983_));
  AOI21_X1   g4598(.A1(new_n4983_), .A2(new_n390_), .B(new_n788_), .ZN(new_n4984_));
  OAI21_X1   g4599(.A1(new_n4984_), .A2(new_n793_), .B(new_n797_), .ZN(new_n4985_));
  AOI21_X1   g4600(.A1(new_n4985_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n4986_));
  OAI21_X1   g4601(.A1(new_n4986_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n4987_));
  AOI21_X1   g4602(.A1(new_n4987_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n4988_));
  OAI21_X1   g4603(.A1(new_n4988_), .A2(new_n912_), .B(new_n917_), .ZN(new_n4989_));
  AOI21_X1   g4604(.A1(new_n4989_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n4990_));
  OAI21_X1   g4605(.A1(new_n4990_), .A2(new_n893_), .B(new_n928_), .ZN(new_n4991_));
  AOI21_X1   g4606(.A1(new_n4991_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n4992_));
  OAI21_X1   g4607(.A1(new_n4992_), .A2(new_n889_), .B(new_n942_), .ZN(new_n4993_));
  AOI21_X1   g4608(.A1(new_n4993_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n4994_));
  OAI21_X1   g4609(.A1(new_n4994_), .A2(new_n952_), .B(new_n957_), .ZN(new_n4995_));
  AOI21_X1   g4610(.A1(new_n4995_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n4996_));
  OAI21_X1   g4611(.A1(new_n4996_), .A2(new_n879_), .B(new_n968_), .ZN(new_n4997_));
  AOI21_X1   g4612(.A1(new_n4997_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n4998_));
  OAI21_X1   g4613(.A1(new_n4998_), .A2(new_n875_), .B(new_n982_), .ZN(new_n4999_));
  AOI21_X1   g4614(.A1(new_n4999_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n5000_));
  OAI21_X1   g4615(.A1(new_n5000_), .A2(new_n992_), .B(new_n997_), .ZN(new_n5001_));
  AOI21_X1   g4616(.A1(new_n5001_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n5002_));
  OAI21_X1   g4617(.A1(new_n5002_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n5003_));
  AOI21_X1   g4618(.A1(new_n5003_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n5004_));
  OAI21_X1   g4619(.A1(new_n5004_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n5005_));
  AOI21_X1   g4620(.A1(new_n5005_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n5006_));
  OAI21_X1   g4621(.A1(new_n5006_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n5007_));
  AOI21_X1   g4622(.A1(new_n5007_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n5008_));
  OAI21_X1   g4623(.A1(new_n5008_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n5009_));
  AOI21_X1   g4624(.A1(new_n5009_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n5010_));
  OAI21_X1   g4625(.A1(new_n5010_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n5011_));
  OAI21_X1   g4626(.A1(new_n1065_), .A2(\priority[78] ), .B(\req[78] ), .ZN(new_n5012_));
  AOI21_X1   g4627(.A1(new_n5011_), .A2(new_n1630_), .B(new_n5012_), .ZN(\grant[78] ));
  NOR2_X1    g4628(.A1(new_n1427_), .A2(new_n1076_), .ZN(new_n5014_));
  OAI21_X1   g4629(.A1(new_n841_), .A2(new_n5014_), .B(new_n1083_), .ZN(new_n5015_));
  AOI21_X1   g4630(.A1(new_n5015_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n5016_));
  OAI21_X1   g4631(.A1(new_n5016_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n5017_));
  AOI21_X1   g4632(.A1(new_n5017_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n5018_));
  OAI21_X1   g4633(.A1(new_n5018_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n5019_));
  AOI21_X1   g4634(.A1(new_n5019_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n5020_));
  OAI21_X1   g4635(.A1(new_n5020_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n5021_));
  AOI21_X1   g4636(.A1(new_n5021_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n5022_));
  OAI21_X1   g4637(.A1(new_n5022_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n5023_));
  AOI21_X1   g4638(.A1(new_n5023_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n5024_));
  OAI21_X1   g4639(.A1(new_n5024_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n5025_));
  AOI21_X1   g4640(.A1(new_n5025_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n5026_));
  OAI21_X1   g4641(.A1(new_n5026_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n5027_));
  AOI21_X1   g4642(.A1(new_n5027_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n5028_));
  OAI21_X1   g4643(.A1(new_n5028_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n5029_));
  AOI21_X1   g4644(.A1(new_n5029_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n5030_));
  OAI21_X1   g4645(.A1(new_n5030_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n5031_));
  AOI21_X1   g4646(.A1(new_n5031_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n5032_));
  OAI21_X1   g4647(.A1(new_n5032_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n5033_));
  AOI21_X1   g4648(.A1(new_n5033_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n5034_));
  OAI21_X1   g4649(.A1(new_n5034_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n5035_));
  AOI21_X1   g4650(.A1(new_n5035_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n5036_));
  OAI21_X1   g4651(.A1(new_n5036_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n5037_));
  AOI21_X1   g4652(.A1(new_n5037_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n5038_));
  OAI21_X1   g4653(.A1(new_n5038_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n5039_));
  AOI21_X1   g4654(.A1(new_n5039_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n5040_));
  OAI21_X1   g4655(.A1(new_n5040_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n5041_));
  AOI21_X1   g4656(.A1(new_n5041_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n5042_));
  OAI21_X1   g4657(.A1(new_n5042_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n5043_));
  AOI21_X1   g4658(.A1(new_n5043_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n5044_));
  OAI21_X1   g4659(.A1(new_n5044_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n5045_));
  AOI21_X1   g4660(.A1(new_n5045_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n5046_));
  OAI21_X1   g4661(.A1(new_n5046_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n5047_));
  AOI21_X1   g4662(.A1(new_n5047_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n5048_));
  OAI21_X1   g4663(.A1(new_n5048_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n5049_));
  AOI21_X1   g4664(.A1(new_n5049_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n5050_));
  OAI21_X1   g4665(.A1(new_n5050_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n5051_));
  AOI21_X1   g4666(.A1(new_n5051_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n5052_));
  OAI21_X1   g4667(.A1(new_n5052_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n5053_));
  AOI21_X1   g4668(.A1(new_n5053_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n5054_));
  OAI21_X1   g4669(.A1(new_n5054_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n5055_));
  OAI21_X1   g4670(.A1(new_n685_), .A2(\priority[79] ), .B(\req[79] ), .ZN(new_n5056_));
  AOI21_X1   g4671(.A1(new_n5055_), .A2(new_n1718_), .B(new_n5056_), .ZN(\grant[79] ));
  NOR2_X1    g4672(.A1(new_n429_), .A2(new_n1431_), .ZN(new_n5058_));
  OAI21_X1   g4673(.A1(new_n1224_), .A2(new_n5058_), .B(new_n1437_), .ZN(new_n5059_));
  AOI21_X1   g4674(.A1(new_n5059_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n5060_));
  OAI21_X1   g4675(.A1(new_n5060_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n5061_));
  AOI21_X1   g4676(.A1(new_n5061_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n5062_));
  OAI21_X1   g4677(.A1(new_n5062_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n5063_));
  AOI21_X1   g4678(.A1(new_n5063_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n5064_));
  OAI21_X1   g4679(.A1(new_n5064_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n5065_));
  AOI21_X1   g4680(.A1(new_n5065_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n5066_));
  OAI21_X1   g4681(.A1(new_n5066_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n5067_));
  AOI21_X1   g4682(.A1(new_n5067_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n5068_));
  OAI21_X1   g4683(.A1(new_n5068_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n5069_));
  AOI21_X1   g4684(.A1(new_n5069_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n5070_));
  OAI21_X1   g4685(.A1(new_n5070_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n5071_));
  AOI21_X1   g4686(.A1(new_n5071_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n5072_));
  OAI21_X1   g4687(.A1(new_n5072_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n5073_));
  AOI21_X1   g4688(.A1(new_n5073_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n5074_));
  OAI21_X1   g4689(.A1(new_n5074_), .A2(new_n506_), .B(new_n514_), .ZN(new_n5075_));
  AOI21_X1   g4690(.A1(new_n5075_), .A2(new_n520_), .B(new_n525_), .ZN(new_n5076_));
  OAI21_X1   g4691(.A1(new_n5076_), .A2(new_n502_), .B(new_n530_), .ZN(new_n5077_));
  AOI21_X1   g4692(.A1(new_n5077_), .A2(new_n498_), .B(new_n536_), .ZN(new_n5078_));
  OAI21_X1   g4693(.A1(new_n5078_), .A2(new_n541_), .B(new_n545_), .ZN(new_n5079_));
  AOI21_X1   g4694(.A1(new_n5079_), .A2(new_n493_), .B(new_n551_), .ZN(new_n5080_));
  OAI21_X1   g4695(.A1(new_n5080_), .A2(new_n488_), .B(new_n556_), .ZN(new_n5081_));
  AOI21_X1   g4696(.A1(new_n5081_), .A2(new_n562_), .B(new_n567_), .ZN(new_n5082_));
  OAI21_X1   g4697(.A1(new_n5082_), .A2(new_n484_), .B(new_n572_), .ZN(new_n5083_));
  AOI21_X1   g4698(.A1(new_n5083_), .A2(new_n480_), .B(new_n578_), .ZN(new_n5084_));
  OAI21_X1   g4699(.A1(new_n5084_), .A2(new_n583_), .B(new_n587_), .ZN(new_n5085_));
  AOI21_X1   g4700(.A1(new_n5085_), .A2(new_n475_), .B(new_n593_), .ZN(new_n5086_));
  OAI21_X1   g4701(.A1(new_n5086_), .A2(new_n470_), .B(new_n598_), .ZN(new_n5087_));
  AOI21_X1   g4702(.A1(new_n5087_), .A2(new_n604_), .B(new_n609_), .ZN(new_n5088_));
  OAI21_X1   g4703(.A1(new_n5088_), .A2(new_n466_), .B(new_n614_), .ZN(new_n5089_));
  AOI21_X1   g4704(.A1(new_n5089_), .A2(new_n462_), .B(new_n620_), .ZN(new_n5090_));
  OAI21_X1   g4705(.A1(new_n5090_), .A2(new_n625_), .B(new_n629_), .ZN(new_n5091_));
  AOI21_X1   g4706(.A1(new_n5091_), .A2(new_n457_), .B(new_n635_), .ZN(new_n5092_));
  OAI21_X1   g4707(.A1(new_n5092_), .A2(new_n452_), .B(new_n640_), .ZN(new_n5093_));
  AOI21_X1   g4708(.A1(new_n5093_), .A2(new_n646_), .B(new_n651_), .ZN(new_n5094_));
  OAI21_X1   g4709(.A1(new_n5094_), .A2(new_n448_), .B(new_n656_), .ZN(new_n5095_));
  AOI21_X1   g4710(.A1(new_n5095_), .A2(new_n444_), .B(new_n662_), .ZN(new_n5096_));
  OAI21_X1   g4711(.A1(new_n5096_), .A2(new_n667_), .B(new_n671_), .ZN(new_n5097_));
  AOI21_X1   g4712(.A1(new_n5097_), .A2(new_n439_), .B(new_n677_), .ZN(new_n5098_));
  OAI21_X1   g4713(.A1(new_n5098_), .A2(new_n434_), .B(new_n682_), .ZN(new_n5099_));
  OAI21_X1   g4714(.A1(new_n689_), .A2(\priority[80] ), .B(\req[80] ), .ZN(new_n5100_));
  AOI21_X1   g4715(.A1(new_n5099_), .A2(new_n688_), .B(new_n5100_), .ZN(\grant[80] ));
  NOR2_X1    g4716(.A1(new_n840_), .A2(new_n697_), .ZN(new_n5102_));
  OAI21_X1   g4717(.A1(new_n425_), .A2(new_n5102_), .B(new_n703_), .ZN(new_n5103_));
  AOI21_X1   g4718(.A1(new_n5103_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n5104_));
  OAI21_X1   g4719(.A1(new_n5104_), .A2(new_n420_), .B(new_n718_), .ZN(new_n5105_));
  AOI21_X1   g4720(.A1(new_n5105_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n5106_));
  OAI21_X1   g4721(.A1(new_n5106_), .A2(new_n729_), .B(new_n734_), .ZN(new_n5107_));
  AOI21_X1   g4722(.A1(new_n5107_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n5108_));
  OAI21_X1   g4723(.A1(new_n5108_), .A2(new_n407_), .B(new_n745_), .ZN(new_n5109_));
  AOI21_X1   g4724(.A1(new_n5109_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n5110_));
  OAI21_X1   g4725(.A1(new_n5110_), .A2(new_n402_), .B(new_n760_), .ZN(new_n5111_));
  AOI21_X1   g4726(.A1(new_n5111_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n5112_));
  OAI21_X1   g4727(.A1(new_n5112_), .A2(new_n771_), .B(new_n776_), .ZN(new_n5113_));
  AOI21_X1   g4728(.A1(new_n5113_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n5114_));
  OAI21_X1   g4729(.A1(new_n5114_), .A2(new_n389_), .B(new_n787_), .ZN(new_n5115_));
  AOI21_X1   g4730(.A1(new_n5115_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n5116_));
  OAI21_X1   g4731(.A1(new_n5116_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n5117_));
  AOI21_X1   g4732(.A1(new_n5117_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n5118_));
  OAI21_X1   g4733(.A1(new_n5118_), .A2(new_n900_), .B(new_n908_), .ZN(new_n5119_));
  AOI21_X1   g4734(.A1(new_n5119_), .A2(new_n913_), .B(new_n918_), .ZN(new_n5120_));
  OAI21_X1   g4735(.A1(new_n5120_), .A2(new_n897_), .B(new_n923_), .ZN(new_n5121_));
  AOI21_X1   g4736(.A1(new_n5121_), .A2(new_n894_), .B(new_n929_), .ZN(new_n5122_));
  OAI21_X1   g4737(.A1(new_n5122_), .A2(new_n933_), .B(new_n937_), .ZN(new_n5123_));
  AOI21_X1   g4738(.A1(new_n5123_), .A2(new_n890_), .B(new_n943_), .ZN(new_n5124_));
  OAI21_X1   g4739(.A1(new_n5124_), .A2(new_n886_), .B(new_n948_), .ZN(new_n5125_));
  AOI21_X1   g4740(.A1(new_n5125_), .A2(new_n953_), .B(new_n958_), .ZN(new_n5126_));
  OAI21_X1   g4741(.A1(new_n5126_), .A2(new_n883_), .B(new_n963_), .ZN(new_n5127_));
  AOI21_X1   g4742(.A1(new_n5127_), .A2(new_n880_), .B(new_n969_), .ZN(new_n5128_));
  OAI21_X1   g4743(.A1(new_n5128_), .A2(new_n973_), .B(new_n977_), .ZN(new_n5129_));
  AOI21_X1   g4744(.A1(new_n5129_), .A2(new_n876_), .B(new_n983_), .ZN(new_n5130_));
  OAI21_X1   g4745(.A1(new_n5130_), .A2(new_n872_), .B(new_n988_), .ZN(new_n5131_));
  AOI21_X1   g4746(.A1(new_n5131_), .A2(new_n993_), .B(new_n998_), .ZN(new_n5132_));
  OAI21_X1   g4747(.A1(new_n5132_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n5133_));
  AOI21_X1   g4748(.A1(new_n5133_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n5134_));
  OAI21_X1   g4749(.A1(new_n5134_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n5135_));
  AOI21_X1   g4750(.A1(new_n5135_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n5136_));
  OAI21_X1   g4751(.A1(new_n5136_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n5137_));
  AOI21_X1   g4752(.A1(new_n5137_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n5138_));
  OAI21_X1   g4753(.A1(new_n5138_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n5139_));
  AOI21_X1   g4754(.A1(new_n5139_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n5140_));
  OAI21_X1   g4755(.A1(new_n5140_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n5141_));
  AOI21_X1   g4756(.A1(new_n5141_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n5142_));
  OAI21_X1   g4757(.A1(new_n5142_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n5143_));
  OAI21_X1   g4758(.A1(new_n1074_), .A2(\priority[81] ), .B(\req[81] ), .ZN(new_n5144_));
  AOI21_X1   g4759(.A1(new_n5143_), .A2(new_n1073_), .B(new_n5144_), .ZN(\grant[81] ));
  NOR2_X1    g4760(.A1(new_n1223_), .A2(new_n1082_), .ZN(new_n5146_));
  OAI21_X1   g4761(.A1(new_n837_), .A2(new_n5146_), .B(new_n1088_), .ZN(new_n5147_));
  AOI21_X1   g4762(.A1(new_n5147_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n5148_));
  OAI21_X1   g4763(.A1(new_n5148_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n5149_));
  AOI21_X1   g4764(.A1(new_n5149_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n5150_));
  OAI21_X1   g4765(.A1(new_n5150_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n5151_));
  AOI21_X1   g4766(.A1(new_n5151_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n5152_));
  OAI21_X1   g4767(.A1(new_n5152_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n5153_));
  AOI21_X1   g4768(.A1(new_n5153_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n5154_));
  OAI21_X1   g4769(.A1(new_n5154_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n5155_));
  AOI21_X1   g4770(.A1(new_n5155_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n5156_));
  OAI21_X1   g4771(.A1(new_n5156_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n5157_));
  AOI21_X1   g4772(.A1(new_n5157_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n5158_));
  OAI21_X1   g4773(.A1(new_n5158_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n5159_));
  AOI21_X1   g4774(.A1(new_n5159_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n5160_));
  OAI21_X1   g4775(.A1(new_n5160_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n5161_));
  AOI21_X1   g4776(.A1(new_n5161_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n5162_));
  OAI21_X1   g4777(.A1(new_n5162_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n5163_));
  AOI21_X1   g4778(.A1(new_n5163_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n5164_));
  OAI21_X1   g4779(.A1(new_n5164_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n5165_));
  AOI21_X1   g4780(.A1(new_n5165_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n5166_));
  OAI21_X1   g4781(.A1(new_n5166_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n5167_));
  AOI21_X1   g4782(.A1(new_n5167_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n5168_));
  OAI21_X1   g4783(.A1(new_n5168_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n5169_));
  AOI21_X1   g4784(.A1(new_n5169_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n5170_));
  OAI21_X1   g4785(.A1(new_n5170_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n5171_));
  AOI21_X1   g4786(.A1(new_n5171_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n5172_));
  OAI21_X1   g4787(.A1(new_n5172_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n5173_));
  AOI21_X1   g4788(.A1(new_n5173_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n5174_));
  OAI21_X1   g4789(.A1(new_n5174_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n5175_));
  AOI21_X1   g4790(.A1(new_n5175_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n5176_));
  OAI21_X1   g4791(.A1(new_n5176_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n5177_));
  AOI21_X1   g4792(.A1(new_n5177_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n5178_));
  OAI21_X1   g4793(.A1(new_n5178_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n5179_));
  AOI21_X1   g4794(.A1(new_n5179_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n5180_));
  OAI21_X1   g4795(.A1(new_n5180_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n5181_));
  AOI21_X1   g4796(.A1(new_n5181_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n5182_));
  OAI21_X1   g4797(.A1(new_n5182_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n5183_));
  AOI21_X1   g4798(.A1(new_n5183_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n5184_));
  OAI21_X1   g4799(.A1(new_n5184_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n5185_));
  AOI21_X1   g4800(.A1(new_n5185_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n5186_));
  OAI21_X1   g4801(.A1(new_n5186_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n5187_));
  OAI21_X1   g4802(.A1(new_n428_), .A2(\priority[82] ), .B(\req[82] ), .ZN(new_n5188_));
  AOI21_X1   g4803(.A1(new_n5187_), .A2(new_n1429_), .B(new_n5188_), .ZN(\grant[82] ));
  NOR2_X1    g4804(.A1(new_n424_), .A2(new_n1436_), .ZN(new_n5190_));
  OAI21_X1   g4805(.A1(new_n1220_), .A2(new_n5190_), .B(new_n1441_), .ZN(new_n5191_));
  AOI21_X1   g4806(.A1(new_n5191_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n5192_));
  OAI21_X1   g4807(.A1(new_n5192_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n5193_));
  AOI21_X1   g4808(.A1(new_n5193_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n5194_));
  OAI21_X1   g4809(.A1(new_n5194_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n5195_));
  AOI21_X1   g4810(.A1(new_n5195_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n5196_));
  OAI21_X1   g4811(.A1(new_n5196_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n5197_));
  AOI21_X1   g4812(.A1(new_n5197_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n5198_));
  OAI21_X1   g4813(.A1(new_n5198_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n5199_));
  AOI21_X1   g4814(.A1(new_n5199_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n5200_));
  OAI21_X1   g4815(.A1(new_n5200_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n5201_));
  AOI21_X1   g4816(.A1(new_n5201_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n5202_));
  OAI21_X1   g4817(.A1(new_n5202_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n5203_));
  AOI21_X1   g4818(.A1(new_n5203_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n5204_));
  OAI21_X1   g4819(.A1(new_n5204_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n5205_));
  AOI21_X1   g4820(.A1(new_n5205_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n5206_));
  OAI21_X1   g4821(.A1(new_n5206_), .A2(new_n519_), .B(new_n524_), .ZN(new_n5207_));
  AOI21_X1   g4822(.A1(new_n5207_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n5208_));
  OAI21_X1   g4823(.A1(new_n5208_), .A2(new_n497_), .B(new_n535_), .ZN(new_n5209_));
  AOI21_X1   g4824(.A1(new_n5209_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n5210_));
  OAI21_X1   g4825(.A1(new_n5210_), .A2(new_n492_), .B(new_n550_), .ZN(new_n5211_));
  AOI21_X1   g4826(.A1(new_n5211_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n5212_));
  OAI21_X1   g4827(.A1(new_n5212_), .A2(new_n561_), .B(new_n566_), .ZN(new_n5213_));
  AOI21_X1   g4828(.A1(new_n5213_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n5214_));
  OAI21_X1   g4829(.A1(new_n5214_), .A2(new_n479_), .B(new_n577_), .ZN(new_n5215_));
  AOI21_X1   g4830(.A1(new_n5215_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n5216_));
  OAI21_X1   g4831(.A1(new_n5216_), .A2(new_n474_), .B(new_n592_), .ZN(new_n5217_));
  AOI21_X1   g4832(.A1(new_n5217_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n5218_));
  OAI21_X1   g4833(.A1(new_n5218_), .A2(new_n603_), .B(new_n608_), .ZN(new_n5219_));
  AOI21_X1   g4834(.A1(new_n5219_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n5220_));
  OAI21_X1   g4835(.A1(new_n5220_), .A2(new_n461_), .B(new_n619_), .ZN(new_n5221_));
  AOI21_X1   g4836(.A1(new_n5221_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n5222_));
  OAI21_X1   g4837(.A1(new_n5222_), .A2(new_n456_), .B(new_n634_), .ZN(new_n5223_));
  AOI21_X1   g4838(.A1(new_n5223_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n5224_));
  OAI21_X1   g4839(.A1(new_n5224_), .A2(new_n645_), .B(new_n650_), .ZN(new_n5225_));
  AOI21_X1   g4840(.A1(new_n5225_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n5226_));
  OAI21_X1   g4841(.A1(new_n5226_), .A2(new_n443_), .B(new_n661_), .ZN(new_n5227_));
  AOI21_X1   g4842(.A1(new_n5227_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n5228_));
  OAI21_X1   g4843(.A1(new_n5228_), .A2(new_n438_), .B(new_n676_), .ZN(new_n5229_));
  AOI21_X1   g4844(.A1(new_n5229_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n5230_));
  OAI21_X1   g4845(.A1(new_n5230_), .A2(new_n687_), .B(new_n692_), .ZN(new_n5231_));
  OAI21_X1   g4846(.A1(new_n695_), .A2(\priority[83] ), .B(\req[83] ), .ZN(new_n5232_));
  AOI21_X1   g4847(.A1(new_n5231_), .A2(new_n1538_), .B(new_n5232_), .ZN(\grant[83] ));
  NOR2_X1    g4848(.A1(new_n836_), .A2(new_n702_), .ZN(new_n5234_));
  OAI21_X1   g4849(.A1(new_n709_), .A2(new_n5234_), .B(new_n713_), .ZN(new_n5235_));
  AOI21_X1   g4850(.A1(new_n5235_), .A2(new_n421_), .B(new_n719_), .ZN(new_n5236_));
  OAI21_X1   g4851(.A1(new_n5236_), .A2(new_n416_), .B(new_n724_), .ZN(new_n5237_));
  AOI21_X1   g4852(.A1(new_n5237_), .A2(new_n730_), .B(new_n735_), .ZN(new_n5238_));
  OAI21_X1   g4853(.A1(new_n5238_), .A2(new_n412_), .B(new_n740_), .ZN(new_n5239_));
  AOI21_X1   g4854(.A1(new_n5239_), .A2(new_n408_), .B(new_n746_), .ZN(new_n5240_));
  OAI21_X1   g4855(.A1(new_n5240_), .A2(new_n751_), .B(new_n755_), .ZN(new_n5241_));
  AOI21_X1   g4856(.A1(new_n5241_), .A2(new_n403_), .B(new_n761_), .ZN(new_n5242_));
  OAI21_X1   g4857(.A1(new_n5242_), .A2(new_n398_), .B(new_n766_), .ZN(new_n5243_));
  AOI21_X1   g4858(.A1(new_n5243_), .A2(new_n772_), .B(new_n777_), .ZN(new_n5244_));
  OAI21_X1   g4859(.A1(new_n5244_), .A2(new_n394_), .B(new_n782_), .ZN(new_n5245_));
  AOI21_X1   g4860(.A1(new_n5245_), .A2(new_n390_), .B(new_n788_), .ZN(new_n5246_));
  OAI21_X1   g4861(.A1(new_n5246_), .A2(new_n793_), .B(new_n797_), .ZN(new_n5247_));
  AOI21_X1   g4862(.A1(new_n5247_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n5248_));
  OAI21_X1   g4863(.A1(new_n5248_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n5249_));
  AOI21_X1   g4864(.A1(new_n5249_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n5250_));
  OAI21_X1   g4865(.A1(new_n5250_), .A2(new_n912_), .B(new_n917_), .ZN(new_n5251_));
  AOI21_X1   g4866(.A1(new_n5251_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n5252_));
  OAI21_X1   g4867(.A1(new_n5252_), .A2(new_n893_), .B(new_n928_), .ZN(new_n5253_));
  AOI21_X1   g4868(.A1(new_n5253_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n5254_));
  OAI21_X1   g4869(.A1(new_n5254_), .A2(new_n889_), .B(new_n942_), .ZN(new_n5255_));
  AOI21_X1   g4870(.A1(new_n5255_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n5256_));
  OAI21_X1   g4871(.A1(new_n5256_), .A2(new_n952_), .B(new_n957_), .ZN(new_n5257_));
  AOI21_X1   g4872(.A1(new_n5257_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n5258_));
  OAI21_X1   g4873(.A1(new_n5258_), .A2(new_n879_), .B(new_n968_), .ZN(new_n5259_));
  AOI21_X1   g4874(.A1(new_n5259_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n5260_));
  OAI21_X1   g4875(.A1(new_n5260_), .A2(new_n875_), .B(new_n982_), .ZN(new_n5261_));
  AOI21_X1   g4876(.A1(new_n5261_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n5262_));
  OAI21_X1   g4877(.A1(new_n5262_), .A2(new_n992_), .B(new_n997_), .ZN(new_n5263_));
  AOI21_X1   g4878(.A1(new_n5263_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n5264_));
  OAI21_X1   g4879(.A1(new_n5264_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n5265_));
  AOI21_X1   g4880(.A1(new_n5265_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n5266_));
  OAI21_X1   g4881(.A1(new_n5266_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n5267_));
  AOI21_X1   g4882(.A1(new_n5267_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n5268_));
  OAI21_X1   g4883(.A1(new_n5268_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n5269_));
  AOI21_X1   g4884(.A1(new_n5269_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n5270_));
  OAI21_X1   g4885(.A1(new_n5270_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n5271_));
  AOI21_X1   g4886(.A1(new_n5271_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n5272_));
  OAI21_X1   g4887(.A1(new_n5272_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n5273_));
  AOI21_X1   g4888(.A1(new_n5273_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n5274_));
  OAI21_X1   g4889(.A1(new_n5274_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n5275_));
  OAI21_X1   g4890(.A1(new_n1080_), .A2(\priority[84] ), .B(\req[84] ), .ZN(new_n5276_));
  AOI21_X1   g4891(.A1(new_n5275_), .A2(new_n1628_), .B(new_n5276_), .ZN(\grant[84] ));
  NOR2_X1    g4892(.A1(new_n1219_), .A2(new_n1087_), .ZN(new_n5278_));
  OAI21_X1   g4893(.A1(new_n1093_), .A2(new_n5278_), .B(new_n1097_), .ZN(new_n5279_));
  AOI21_X1   g4894(.A1(new_n5279_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n5280_));
  OAI21_X1   g4895(.A1(new_n5280_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n5281_));
  AOI21_X1   g4896(.A1(new_n5281_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n5282_));
  OAI21_X1   g4897(.A1(new_n5282_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n5283_));
  AOI21_X1   g4898(.A1(new_n5283_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n5284_));
  OAI21_X1   g4899(.A1(new_n5284_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n5285_));
  AOI21_X1   g4900(.A1(new_n5285_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n5286_));
  OAI21_X1   g4901(.A1(new_n5286_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n5287_));
  AOI21_X1   g4902(.A1(new_n5287_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n5288_));
  OAI21_X1   g4903(.A1(new_n5288_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n5289_));
  AOI21_X1   g4904(.A1(new_n5289_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n5290_));
  OAI21_X1   g4905(.A1(new_n5290_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n5291_));
  AOI21_X1   g4906(.A1(new_n5291_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n5292_));
  OAI21_X1   g4907(.A1(new_n5292_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n5293_));
  AOI21_X1   g4908(.A1(new_n5293_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n5294_));
  OAI21_X1   g4909(.A1(new_n5294_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n5295_));
  AOI21_X1   g4910(.A1(new_n5295_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n5296_));
  OAI21_X1   g4911(.A1(new_n5296_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n5297_));
  AOI21_X1   g4912(.A1(new_n5297_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n5298_));
  OAI21_X1   g4913(.A1(new_n5298_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n5299_));
  AOI21_X1   g4914(.A1(new_n5299_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n5300_));
  OAI21_X1   g4915(.A1(new_n5300_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n5301_));
  AOI21_X1   g4916(.A1(new_n5301_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n5302_));
  OAI21_X1   g4917(.A1(new_n5302_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n5303_));
  AOI21_X1   g4918(.A1(new_n5303_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n5304_));
  OAI21_X1   g4919(.A1(new_n5304_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n5305_));
  AOI21_X1   g4920(.A1(new_n5305_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n5306_));
  OAI21_X1   g4921(.A1(new_n5306_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n5307_));
  AOI21_X1   g4922(.A1(new_n5307_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n5308_));
  OAI21_X1   g4923(.A1(new_n5308_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n5309_));
  AOI21_X1   g4924(.A1(new_n5309_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n5310_));
  OAI21_X1   g4925(.A1(new_n5310_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n5311_));
  AOI21_X1   g4926(.A1(new_n5311_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n5312_));
  OAI21_X1   g4927(.A1(new_n5312_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n5313_));
  AOI21_X1   g4928(.A1(new_n5313_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n5314_));
  OAI21_X1   g4929(.A1(new_n5314_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n5315_));
  AOI21_X1   g4930(.A1(new_n5315_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n5316_));
  OAI21_X1   g4931(.A1(new_n5316_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n5317_));
  AOI21_X1   g4932(.A1(new_n5317_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n5318_));
  OAI21_X1   g4933(.A1(new_n5318_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n5319_));
  OAI21_X1   g4934(.A1(new_n423_), .A2(\priority[85] ), .B(\req[85] ), .ZN(new_n5320_));
  AOI21_X1   g4935(.A1(new_n5319_), .A2(new_n1716_), .B(new_n5320_), .ZN(\grant[85] ));
  NOR2_X1    g4936(.A1(new_n708_), .A2(new_n1440_), .ZN(new_n5322_));
  OAI21_X1   g4937(.A1(new_n1446_), .A2(new_n5322_), .B(new_n1449_), .ZN(new_n5323_));
  AOI21_X1   g4938(.A1(new_n5323_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n5324_));
  OAI21_X1   g4939(.A1(new_n5324_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n5325_));
  AOI21_X1   g4940(.A1(new_n5325_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n5326_));
  OAI21_X1   g4941(.A1(new_n5326_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n5327_));
  AOI21_X1   g4942(.A1(new_n5327_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n5328_));
  OAI21_X1   g4943(.A1(new_n5328_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n5329_));
  AOI21_X1   g4944(.A1(new_n5329_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n5330_));
  OAI21_X1   g4945(.A1(new_n5330_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n5331_));
  AOI21_X1   g4946(.A1(new_n5331_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n5332_));
  OAI21_X1   g4947(.A1(new_n5332_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n5333_));
  AOI21_X1   g4948(.A1(new_n5333_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n5334_));
  OAI21_X1   g4949(.A1(new_n5334_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n5335_));
  AOI21_X1   g4950(.A1(new_n5335_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n5336_));
  OAI21_X1   g4951(.A1(new_n5336_), .A2(new_n506_), .B(new_n514_), .ZN(new_n5337_));
  AOI21_X1   g4952(.A1(new_n5337_), .A2(new_n520_), .B(new_n525_), .ZN(new_n5338_));
  OAI21_X1   g4953(.A1(new_n5338_), .A2(new_n502_), .B(new_n530_), .ZN(new_n5339_));
  AOI21_X1   g4954(.A1(new_n5339_), .A2(new_n498_), .B(new_n536_), .ZN(new_n5340_));
  OAI21_X1   g4955(.A1(new_n5340_), .A2(new_n541_), .B(new_n545_), .ZN(new_n5341_));
  AOI21_X1   g4956(.A1(new_n5341_), .A2(new_n493_), .B(new_n551_), .ZN(new_n5342_));
  OAI21_X1   g4957(.A1(new_n5342_), .A2(new_n488_), .B(new_n556_), .ZN(new_n5343_));
  AOI21_X1   g4958(.A1(new_n5343_), .A2(new_n562_), .B(new_n567_), .ZN(new_n5344_));
  OAI21_X1   g4959(.A1(new_n5344_), .A2(new_n484_), .B(new_n572_), .ZN(new_n5345_));
  AOI21_X1   g4960(.A1(new_n5345_), .A2(new_n480_), .B(new_n578_), .ZN(new_n5346_));
  OAI21_X1   g4961(.A1(new_n5346_), .A2(new_n583_), .B(new_n587_), .ZN(new_n5347_));
  AOI21_X1   g4962(.A1(new_n5347_), .A2(new_n475_), .B(new_n593_), .ZN(new_n5348_));
  OAI21_X1   g4963(.A1(new_n5348_), .A2(new_n470_), .B(new_n598_), .ZN(new_n5349_));
  AOI21_X1   g4964(.A1(new_n5349_), .A2(new_n604_), .B(new_n609_), .ZN(new_n5350_));
  OAI21_X1   g4965(.A1(new_n5350_), .A2(new_n466_), .B(new_n614_), .ZN(new_n5351_));
  AOI21_X1   g4966(.A1(new_n5351_), .A2(new_n462_), .B(new_n620_), .ZN(new_n5352_));
  OAI21_X1   g4967(.A1(new_n5352_), .A2(new_n625_), .B(new_n629_), .ZN(new_n5353_));
  AOI21_X1   g4968(.A1(new_n5353_), .A2(new_n457_), .B(new_n635_), .ZN(new_n5354_));
  OAI21_X1   g4969(.A1(new_n5354_), .A2(new_n452_), .B(new_n640_), .ZN(new_n5355_));
  AOI21_X1   g4970(.A1(new_n5355_), .A2(new_n646_), .B(new_n651_), .ZN(new_n5356_));
  OAI21_X1   g4971(.A1(new_n5356_), .A2(new_n448_), .B(new_n656_), .ZN(new_n5357_));
  AOI21_X1   g4972(.A1(new_n5357_), .A2(new_n444_), .B(new_n662_), .ZN(new_n5358_));
  OAI21_X1   g4973(.A1(new_n5358_), .A2(new_n667_), .B(new_n671_), .ZN(new_n5359_));
  AOI21_X1   g4974(.A1(new_n5359_), .A2(new_n439_), .B(new_n677_), .ZN(new_n5360_));
  OAI21_X1   g4975(.A1(new_n5360_), .A2(new_n434_), .B(new_n682_), .ZN(new_n5361_));
  AOI21_X1   g4976(.A1(new_n5361_), .A2(new_n688_), .B(new_n693_), .ZN(new_n5362_));
  OAI21_X1   g4977(.A1(new_n5362_), .A2(new_n430_), .B(new_n698_), .ZN(new_n5363_));
  OAI21_X1   g4978(.A1(new_n700_), .A2(\priority[86] ), .B(\req[86] ), .ZN(new_n5364_));
  AOI21_X1   g4979(.A1(new_n5363_), .A2(new_n426_), .B(new_n5364_), .ZN(\grant[86] ));
  NOR2_X1    g4980(.A1(new_n1092_), .A2(new_n712_), .ZN(new_n5366_));
  OAI21_X1   g4981(.A1(new_n420_), .A2(new_n5366_), .B(new_n718_), .ZN(new_n5367_));
  AOI21_X1   g4982(.A1(new_n5367_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n5368_));
  OAI21_X1   g4983(.A1(new_n5368_), .A2(new_n729_), .B(new_n734_), .ZN(new_n5369_));
  AOI21_X1   g4984(.A1(new_n5369_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n5370_));
  OAI21_X1   g4985(.A1(new_n5370_), .A2(new_n407_), .B(new_n745_), .ZN(new_n5371_));
  AOI21_X1   g4986(.A1(new_n5371_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n5372_));
  OAI21_X1   g4987(.A1(new_n5372_), .A2(new_n402_), .B(new_n760_), .ZN(new_n5373_));
  AOI21_X1   g4988(.A1(new_n5373_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n5374_));
  OAI21_X1   g4989(.A1(new_n5374_), .A2(new_n771_), .B(new_n776_), .ZN(new_n5375_));
  AOI21_X1   g4990(.A1(new_n5375_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n5376_));
  OAI21_X1   g4991(.A1(new_n5376_), .A2(new_n389_), .B(new_n787_), .ZN(new_n5377_));
  AOI21_X1   g4992(.A1(new_n5377_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n5378_));
  OAI21_X1   g4993(.A1(new_n5378_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n5379_));
  AOI21_X1   g4994(.A1(new_n5379_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n5380_));
  OAI21_X1   g4995(.A1(new_n5380_), .A2(new_n900_), .B(new_n908_), .ZN(new_n5381_));
  AOI21_X1   g4996(.A1(new_n5381_), .A2(new_n913_), .B(new_n918_), .ZN(new_n5382_));
  OAI21_X1   g4997(.A1(new_n5382_), .A2(new_n897_), .B(new_n923_), .ZN(new_n5383_));
  AOI21_X1   g4998(.A1(new_n5383_), .A2(new_n894_), .B(new_n929_), .ZN(new_n5384_));
  OAI21_X1   g4999(.A1(new_n5384_), .A2(new_n933_), .B(new_n937_), .ZN(new_n5385_));
  AOI21_X1   g5000(.A1(new_n5385_), .A2(new_n890_), .B(new_n943_), .ZN(new_n5386_));
  OAI21_X1   g5001(.A1(new_n5386_), .A2(new_n886_), .B(new_n948_), .ZN(new_n5387_));
  AOI21_X1   g5002(.A1(new_n5387_), .A2(new_n953_), .B(new_n958_), .ZN(new_n5388_));
  OAI21_X1   g5003(.A1(new_n5388_), .A2(new_n883_), .B(new_n963_), .ZN(new_n5389_));
  AOI21_X1   g5004(.A1(new_n5389_), .A2(new_n880_), .B(new_n969_), .ZN(new_n5390_));
  OAI21_X1   g5005(.A1(new_n5390_), .A2(new_n973_), .B(new_n977_), .ZN(new_n5391_));
  AOI21_X1   g5006(.A1(new_n5391_), .A2(new_n876_), .B(new_n983_), .ZN(new_n5392_));
  OAI21_X1   g5007(.A1(new_n5392_), .A2(new_n872_), .B(new_n988_), .ZN(new_n5393_));
  AOI21_X1   g5008(.A1(new_n5393_), .A2(new_n993_), .B(new_n998_), .ZN(new_n5394_));
  OAI21_X1   g5009(.A1(new_n5394_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n5395_));
  AOI21_X1   g5010(.A1(new_n5395_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n5396_));
  OAI21_X1   g5011(.A1(new_n5396_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n5397_));
  AOI21_X1   g5012(.A1(new_n5397_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n5398_));
  OAI21_X1   g5013(.A1(new_n5398_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n5399_));
  AOI21_X1   g5014(.A1(new_n5399_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n5400_));
  OAI21_X1   g5015(.A1(new_n5400_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n5401_));
  AOI21_X1   g5016(.A1(new_n5401_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n5402_));
  OAI21_X1   g5017(.A1(new_n5402_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n5403_));
  AOI21_X1   g5018(.A1(new_n5403_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n5404_));
  OAI21_X1   g5019(.A1(new_n5404_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n5405_));
  AOI21_X1   g5020(.A1(new_n5405_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n5406_));
  OAI21_X1   g5021(.A1(new_n5406_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n5407_));
  OAI21_X1   g5022(.A1(new_n1085_), .A2(\priority[87] ), .B(\req[87] ), .ZN(new_n5408_));
  AOI21_X1   g5023(.A1(new_n5407_), .A2(new_n838_), .B(new_n5408_), .ZN(\grant[87] ));
  NOR2_X1    g5024(.A1(new_n1445_), .A2(new_n1096_), .ZN(new_n5410_));
  OAI21_X1   g5025(.A1(new_n833_), .A2(new_n5410_), .B(new_n1102_), .ZN(new_n5411_));
  AOI21_X1   g5026(.A1(new_n5411_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n5412_));
  OAI21_X1   g5027(.A1(new_n5412_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n5413_));
  AOI21_X1   g5028(.A1(new_n5413_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n5414_));
  OAI21_X1   g5029(.A1(new_n5414_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n5415_));
  AOI21_X1   g5030(.A1(new_n5415_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n5416_));
  OAI21_X1   g5031(.A1(new_n5416_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n5417_));
  AOI21_X1   g5032(.A1(new_n5417_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n5418_));
  OAI21_X1   g5033(.A1(new_n5418_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n5419_));
  AOI21_X1   g5034(.A1(new_n5419_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n5420_));
  OAI21_X1   g5035(.A1(new_n5420_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n5421_));
  AOI21_X1   g5036(.A1(new_n5421_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n5422_));
  OAI21_X1   g5037(.A1(new_n5422_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n5423_));
  AOI21_X1   g5038(.A1(new_n5423_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n5424_));
  OAI21_X1   g5039(.A1(new_n5424_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n5425_));
  AOI21_X1   g5040(.A1(new_n5425_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n5426_));
  OAI21_X1   g5041(.A1(new_n5426_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n5427_));
  AOI21_X1   g5042(.A1(new_n5427_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n5428_));
  OAI21_X1   g5043(.A1(new_n5428_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n5429_));
  AOI21_X1   g5044(.A1(new_n5429_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n5430_));
  OAI21_X1   g5045(.A1(new_n5430_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n5431_));
  AOI21_X1   g5046(.A1(new_n5431_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n5432_));
  OAI21_X1   g5047(.A1(new_n5432_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n5433_));
  AOI21_X1   g5048(.A1(new_n5433_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n5434_));
  OAI21_X1   g5049(.A1(new_n5434_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n5435_));
  AOI21_X1   g5050(.A1(new_n5435_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n5436_));
  OAI21_X1   g5051(.A1(new_n5436_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n5437_));
  AOI21_X1   g5052(.A1(new_n5437_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n5438_));
  OAI21_X1   g5053(.A1(new_n5438_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n5439_));
  AOI21_X1   g5054(.A1(new_n5439_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n5440_));
  OAI21_X1   g5055(.A1(new_n5440_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n5441_));
  AOI21_X1   g5056(.A1(new_n5441_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n5442_));
  OAI21_X1   g5057(.A1(new_n5442_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n5443_));
  AOI21_X1   g5058(.A1(new_n5443_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n5444_));
  OAI21_X1   g5059(.A1(new_n5444_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n5445_));
  AOI21_X1   g5060(.A1(new_n5445_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n5446_));
  OAI21_X1   g5061(.A1(new_n5446_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n5447_));
  AOI21_X1   g5062(.A1(new_n5447_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n5448_));
  OAI21_X1   g5063(.A1(new_n5448_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n5449_));
  AOI21_X1   g5064(.A1(new_n5449_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n5450_));
  OAI21_X1   g5065(.A1(new_n5450_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n5451_));
  OAI21_X1   g5066(.A1(new_n707_), .A2(\priority[88] ), .B(\req[88] ), .ZN(new_n5452_));
  AOI21_X1   g5067(.A1(new_n5451_), .A2(new_n1221_), .B(new_n5452_), .ZN(\grant[88] ));
  NOR2_X1    g5068(.A1(new_n419_), .A2(new_n1448_), .ZN(new_n5454_));
  OAI21_X1   g5069(.A1(new_n1216_), .A2(new_n5454_), .B(new_n1453_), .ZN(new_n5455_));
  AOI21_X1   g5070(.A1(new_n5455_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n5456_));
  OAI21_X1   g5071(.A1(new_n5456_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n5457_));
  AOI21_X1   g5072(.A1(new_n5457_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n5458_));
  OAI21_X1   g5073(.A1(new_n5458_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n5459_));
  AOI21_X1   g5074(.A1(new_n5459_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n5460_));
  OAI21_X1   g5075(.A1(new_n5460_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n5461_));
  AOI21_X1   g5076(.A1(new_n5461_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n5462_));
  OAI21_X1   g5077(.A1(new_n5462_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n5463_));
  AOI21_X1   g5078(.A1(new_n5463_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n5464_));
  OAI21_X1   g5079(.A1(new_n5464_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n5465_));
  AOI21_X1   g5080(.A1(new_n5465_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n5466_));
  OAI21_X1   g5081(.A1(new_n5466_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n5467_));
  AOI21_X1   g5082(.A1(new_n5467_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n5468_));
  OAI21_X1   g5083(.A1(new_n5468_), .A2(new_n519_), .B(new_n524_), .ZN(new_n5469_));
  AOI21_X1   g5084(.A1(new_n5469_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n5470_));
  OAI21_X1   g5085(.A1(new_n5470_), .A2(new_n497_), .B(new_n535_), .ZN(new_n5471_));
  AOI21_X1   g5086(.A1(new_n5471_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n5472_));
  OAI21_X1   g5087(.A1(new_n5472_), .A2(new_n492_), .B(new_n550_), .ZN(new_n5473_));
  AOI21_X1   g5088(.A1(new_n5473_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n5474_));
  OAI21_X1   g5089(.A1(new_n5474_), .A2(new_n561_), .B(new_n566_), .ZN(new_n5475_));
  AOI21_X1   g5090(.A1(new_n5475_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n5476_));
  OAI21_X1   g5091(.A1(new_n5476_), .A2(new_n479_), .B(new_n577_), .ZN(new_n5477_));
  AOI21_X1   g5092(.A1(new_n5477_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n5478_));
  OAI21_X1   g5093(.A1(new_n5478_), .A2(new_n474_), .B(new_n592_), .ZN(new_n5479_));
  AOI21_X1   g5094(.A1(new_n5479_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n5480_));
  OAI21_X1   g5095(.A1(new_n5480_), .A2(new_n603_), .B(new_n608_), .ZN(new_n5481_));
  AOI21_X1   g5096(.A1(new_n5481_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n5482_));
  OAI21_X1   g5097(.A1(new_n5482_), .A2(new_n461_), .B(new_n619_), .ZN(new_n5483_));
  AOI21_X1   g5098(.A1(new_n5483_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n5484_));
  OAI21_X1   g5099(.A1(new_n5484_), .A2(new_n456_), .B(new_n634_), .ZN(new_n5485_));
  AOI21_X1   g5100(.A1(new_n5485_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n5486_));
  OAI21_X1   g5101(.A1(new_n5486_), .A2(new_n645_), .B(new_n650_), .ZN(new_n5487_));
  AOI21_X1   g5102(.A1(new_n5487_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n5488_));
  OAI21_X1   g5103(.A1(new_n5488_), .A2(new_n443_), .B(new_n661_), .ZN(new_n5489_));
  AOI21_X1   g5104(.A1(new_n5489_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n5490_));
  OAI21_X1   g5105(.A1(new_n5490_), .A2(new_n438_), .B(new_n676_), .ZN(new_n5491_));
  AOI21_X1   g5106(.A1(new_n5491_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n5492_));
  OAI21_X1   g5107(.A1(new_n5492_), .A2(new_n687_), .B(new_n692_), .ZN(new_n5493_));
  AOI21_X1   g5108(.A1(new_n5493_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n5494_));
  OAI21_X1   g5109(.A1(new_n5494_), .A2(new_n425_), .B(new_n703_), .ZN(new_n5495_));
  OAI21_X1   g5110(.A1(new_n710_), .A2(\priority[89] ), .B(\req[89] ), .ZN(new_n5496_));
  AOI21_X1   g5111(.A1(new_n5495_), .A2(new_n1536_), .B(new_n5496_), .ZN(\grant[89] ));
  NOR2_X1    g5112(.A1(new_n832_), .A2(new_n717_), .ZN(new_n5498_));
  OAI21_X1   g5113(.A1(new_n416_), .A2(new_n5498_), .B(new_n724_), .ZN(new_n5499_));
  AOI21_X1   g5114(.A1(new_n5499_), .A2(new_n730_), .B(new_n735_), .ZN(new_n5500_));
  OAI21_X1   g5115(.A1(new_n5500_), .A2(new_n412_), .B(new_n740_), .ZN(new_n5501_));
  AOI21_X1   g5116(.A1(new_n5501_), .A2(new_n408_), .B(new_n746_), .ZN(new_n5502_));
  OAI21_X1   g5117(.A1(new_n5502_), .A2(new_n751_), .B(new_n755_), .ZN(new_n5503_));
  AOI21_X1   g5118(.A1(new_n5503_), .A2(new_n403_), .B(new_n761_), .ZN(new_n5504_));
  OAI21_X1   g5119(.A1(new_n5504_), .A2(new_n398_), .B(new_n766_), .ZN(new_n5505_));
  AOI21_X1   g5120(.A1(new_n5505_), .A2(new_n772_), .B(new_n777_), .ZN(new_n5506_));
  OAI21_X1   g5121(.A1(new_n5506_), .A2(new_n394_), .B(new_n782_), .ZN(new_n5507_));
  AOI21_X1   g5122(.A1(new_n5507_), .A2(new_n390_), .B(new_n788_), .ZN(new_n5508_));
  OAI21_X1   g5123(.A1(new_n5508_), .A2(new_n793_), .B(new_n797_), .ZN(new_n5509_));
  AOI21_X1   g5124(.A1(new_n5509_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n5510_));
  OAI21_X1   g5125(.A1(new_n5510_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n5511_));
  AOI21_X1   g5126(.A1(new_n5511_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n5512_));
  OAI21_X1   g5127(.A1(new_n5512_), .A2(new_n912_), .B(new_n917_), .ZN(new_n5513_));
  AOI21_X1   g5128(.A1(new_n5513_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n5514_));
  OAI21_X1   g5129(.A1(new_n5514_), .A2(new_n893_), .B(new_n928_), .ZN(new_n5515_));
  AOI21_X1   g5130(.A1(new_n5515_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n5516_));
  OAI21_X1   g5131(.A1(new_n5516_), .A2(new_n889_), .B(new_n942_), .ZN(new_n5517_));
  AOI21_X1   g5132(.A1(new_n5517_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n5518_));
  OAI21_X1   g5133(.A1(new_n5518_), .A2(new_n952_), .B(new_n957_), .ZN(new_n5519_));
  AOI21_X1   g5134(.A1(new_n5519_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n5520_));
  OAI21_X1   g5135(.A1(new_n5520_), .A2(new_n879_), .B(new_n968_), .ZN(new_n5521_));
  AOI21_X1   g5136(.A1(new_n5521_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n5522_));
  OAI21_X1   g5137(.A1(new_n5522_), .A2(new_n875_), .B(new_n982_), .ZN(new_n5523_));
  AOI21_X1   g5138(.A1(new_n5523_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n5524_));
  OAI21_X1   g5139(.A1(new_n5524_), .A2(new_n992_), .B(new_n997_), .ZN(new_n5525_));
  AOI21_X1   g5140(.A1(new_n5525_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n5526_));
  OAI21_X1   g5141(.A1(new_n5526_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n5527_));
  AOI21_X1   g5142(.A1(new_n5527_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n5528_));
  OAI21_X1   g5143(.A1(new_n5528_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n5529_));
  AOI21_X1   g5144(.A1(new_n5529_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n5530_));
  OAI21_X1   g5145(.A1(new_n5530_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n5531_));
  AOI21_X1   g5146(.A1(new_n5531_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n5532_));
  OAI21_X1   g5147(.A1(new_n5532_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n5533_));
  AOI21_X1   g5148(.A1(new_n5533_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n5534_));
  OAI21_X1   g5149(.A1(new_n5534_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n5535_));
  AOI21_X1   g5150(.A1(new_n5535_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n5536_));
  OAI21_X1   g5151(.A1(new_n5536_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n5537_));
  AOI21_X1   g5152(.A1(new_n5537_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n5538_));
  OAI21_X1   g5153(.A1(new_n5538_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n5539_));
  OAI21_X1   g5154(.A1(new_n1094_), .A2(\priority[90] ), .B(\req[90] ), .ZN(new_n5540_));
  AOI21_X1   g5155(.A1(new_n5539_), .A2(new_n1626_), .B(new_n5540_), .ZN(\grant[90] ));
  NOR2_X1    g5156(.A1(new_n1215_), .A2(new_n1101_), .ZN(new_n5542_));
  OAI21_X1   g5157(.A1(new_n830_), .A2(new_n5542_), .B(new_n1108_), .ZN(new_n5543_));
  AOI21_X1   g5158(.A1(new_n5543_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n5544_));
  OAI21_X1   g5159(.A1(new_n5544_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n5545_));
  AOI21_X1   g5160(.A1(new_n5545_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n5546_));
  OAI21_X1   g5161(.A1(new_n5546_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n5547_));
  AOI21_X1   g5162(.A1(new_n5547_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n5548_));
  OAI21_X1   g5163(.A1(new_n5548_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n5549_));
  AOI21_X1   g5164(.A1(new_n5549_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n5550_));
  OAI21_X1   g5165(.A1(new_n5550_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n5551_));
  AOI21_X1   g5166(.A1(new_n5551_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n5552_));
  OAI21_X1   g5167(.A1(new_n5552_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n5553_));
  AOI21_X1   g5168(.A1(new_n5553_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n5554_));
  OAI21_X1   g5169(.A1(new_n5554_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n5555_));
  AOI21_X1   g5170(.A1(new_n5555_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n5556_));
  OAI21_X1   g5171(.A1(new_n5556_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n5557_));
  AOI21_X1   g5172(.A1(new_n5557_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n5558_));
  OAI21_X1   g5173(.A1(new_n5558_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n5559_));
  AOI21_X1   g5174(.A1(new_n5559_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n5560_));
  OAI21_X1   g5175(.A1(new_n5560_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n5561_));
  AOI21_X1   g5176(.A1(new_n5561_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n5562_));
  OAI21_X1   g5177(.A1(new_n5562_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n5563_));
  AOI21_X1   g5178(.A1(new_n5563_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n5564_));
  OAI21_X1   g5179(.A1(new_n5564_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n5565_));
  AOI21_X1   g5180(.A1(new_n5565_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n5566_));
  OAI21_X1   g5181(.A1(new_n5566_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n5567_));
  AOI21_X1   g5182(.A1(new_n5567_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n5568_));
  OAI21_X1   g5183(.A1(new_n5568_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n5569_));
  AOI21_X1   g5184(.A1(new_n5569_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n5570_));
  OAI21_X1   g5185(.A1(new_n5570_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n5571_));
  AOI21_X1   g5186(.A1(new_n5571_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n5572_));
  OAI21_X1   g5187(.A1(new_n5572_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n5573_));
  AOI21_X1   g5188(.A1(new_n5573_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n5574_));
  OAI21_X1   g5189(.A1(new_n5574_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n5575_));
  AOI21_X1   g5190(.A1(new_n5575_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n5576_));
  OAI21_X1   g5191(.A1(new_n5576_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n5577_));
  AOI21_X1   g5192(.A1(new_n5577_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n5578_));
  OAI21_X1   g5193(.A1(new_n5578_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n5579_));
  AOI21_X1   g5194(.A1(new_n5579_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n5580_));
  OAI21_X1   g5195(.A1(new_n5580_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n5581_));
  AOI21_X1   g5196(.A1(new_n5581_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n5582_));
  OAI21_X1   g5197(.A1(new_n5582_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n5583_));
  OAI21_X1   g5198(.A1(new_n418_), .A2(\priority[91] ), .B(\req[91] ), .ZN(new_n5584_));
  AOI21_X1   g5199(.A1(new_n5583_), .A2(new_n1714_), .B(new_n5584_), .ZN(\grant[91] ));
  NOR2_X1    g5200(.A1(new_n415_), .A2(new_n1452_), .ZN(new_n5586_));
  OAI21_X1   g5201(.A1(new_n1213_), .A2(new_n5586_), .B(new_n1458_), .ZN(new_n5587_));
  AOI21_X1   g5202(.A1(new_n5587_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n5588_));
  OAI21_X1   g5203(.A1(new_n5588_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n5589_));
  AOI21_X1   g5204(.A1(new_n5589_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n5590_));
  OAI21_X1   g5205(.A1(new_n5590_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n5591_));
  AOI21_X1   g5206(.A1(new_n5591_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n5592_));
  OAI21_X1   g5207(.A1(new_n5592_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n5593_));
  AOI21_X1   g5208(.A1(new_n5593_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n5594_));
  OAI21_X1   g5209(.A1(new_n5594_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n5595_));
  AOI21_X1   g5210(.A1(new_n5595_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n5596_));
  OAI21_X1   g5211(.A1(new_n5596_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n5597_));
  AOI21_X1   g5212(.A1(new_n5597_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n5598_));
  OAI21_X1   g5213(.A1(new_n5598_), .A2(new_n506_), .B(new_n514_), .ZN(new_n5599_));
  AOI21_X1   g5214(.A1(new_n5599_), .A2(new_n520_), .B(new_n525_), .ZN(new_n5600_));
  OAI21_X1   g5215(.A1(new_n5600_), .A2(new_n502_), .B(new_n530_), .ZN(new_n5601_));
  AOI21_X1   g5216(.A1(new_n5601_), .A2(new_n498_), .B(new_n536_), .ZN(new_n5602_));
  OAI21_X1   g5217(.A1(new_n5602_), .A2(new_n541_), .B(new_n545_), .ZN(new_n5603_));
  AOI21_X1   g5218(.A1(new_n5603_), .A2(new_n493_), .B(new_n551_), .ZN(new_n5604_));
  OAI21_X1   g5219(.A1(new_n5604_), .A2(new_n488_), .B(new_n556_), .ZN(new_n5605_));
  AOI21_X1   g5220(.A1(new_n5605_), .A2(new_n562_), .B(new_n567_), .ZN(new_n5606_));
  OAI21_X1   g5221(.A1(new_n5606_), .A2(new_n484_), .B(new_n572_), .ZN(new_n5607_));
  AOI21_X1   g5222(.A1(new_n5607_), .A2(new_n480_), .B(new_n578_), .ZN(new_n5608_));
  OAI21_X1   g5223(.A1(new_n5608_), .A2(new_n583_), .B(new_n587_), .ZN(new_n5609_));
  AOI21_X1   g5224(.A1(new_n5609_), .A2(new_n475_), .B(new_n593_), .ZN(new_n5610_));
  OAI21_X1   g5225(.A1(new_n5610_), .A2(new_n470_), .B(new_n598_), .ZN(new_n5611_));
  AOI21_X1   g5226(.A1(new_n5611_), .A2(new_n604_), .B(new_n609_), .ZN(new_n5612_));
  OAI21_X1   g5227(.A1(new_n5612_), .A2(new_n466_), .B(new_n614_), .ZN(new_n5613_));
  AOI21_X1   g5228(.A1(new_n5613_), .A2(new_n462_), .B(new_n620_), .ZN(new_n5614_));
  OAI21_X1   g5229(.A1(new_n5614_), .A2(new_n625_), .B(new_n629_), .ZN(new_n5615_));
  AOI21_X1   g5230(.A1(new_n5615_), .A2(new_n457_), .B(new_n635_), .ZN(new_n5616_));
  OAI21_X1   g5231(.A1(new_n5616_), .A2(new_n452_), .B(new_n640_), .ZN(new_n5617_));
  AOI21_X1   g5232(.A1(new_n5617_), .A2(new_n646_), .B(new_n651_), .ZN(new_n5618_));
  OAI21_X1   g5233(.A1(new_n5618_), .A2(new_n448_), .B(new_n656_), .ZN(new_n5619_));
  AOI21_X1   g5234(.A1(new_n5619_), .A2(new_n444_), .B(new_n662_), .ZN(new_n5620_));
  OAI21_X1   g5235(.A1(new_n5620_), .A2(new_n667_), .B(new_n671_), .ZN(new_n5621_));
  AOI21_X1   g5236(.A1(new_n5621_), .A2(new_n439_), .B(new_n677_), .ZN(new_n5622_));
  OAI21_X1   g5237(.A1(new_n5622_), .A2(new_n434_), .B(new_n682_), .ZN(new_n5623_));
  AOI21_X1   g5238(.A1(new_n5623_), .A2(new_n688_), .B(new_n693_), .ZN(new_n5624_));
  OAI21_X1   g5239(.A1(new_n5624_), .A2(new_n430_), .B(new_n698_), .ZN(new_n5625_));
  AOI21_X1   g5240(.A1(new_n5625_), .A2(new_n426_), .B(new_n704_), .ZN(new_n5626_));
  OAI21_X1   g5241(.A1(new_n5626_), .A2(new_n709_), .B(new_n713_), .ZN(new_n5627_));
  OAI21_X1   g5242(.A1(new_n715_), .A2(\priority[92] ), .B(\req[92] ), .ZN(new_n5628_));
  AOI21_X1   g5243(.A1(new_n5627_), .A2(new_n421_), .B(new_n5628_), .ZN(\grant[92] ));
  NOR2_X1    g5244(.A1(new_n829_), .A2(new_n723_), .ZN(new_n5630_));
  OAI21_X1   g5245(.A1(new_n729_), .A2(new_n5630_), .B(new_n734_), .ZN(new_n5631_));
  AOI21_X1   g5246(.A1(new_n5631_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n5632_));
  OAI21_X1   g5247(.A1(new_n5632_), .A2(new_n407_), .B(new_n745_), .ZN(new_n5633_));
  AOI21_X1   g5248(.A1(new_n5633_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n5634_));
  OAI21_X1   g5249(.A1(new_n5634_), .A2(new_n402_), .B(new_n760_), .ZN(new_n5635_));
  AOI21_X1   g5250(.A1(new_n5635_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n5636_));
  OAI21_X1   g5251(.A1(new_n5636_), .A2(new_n771_), .B(new_n776_), .ZN(new_n5637_));
  AOI21_X1   g5252(.A1(new_n5637_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n5638_));
  OAI21_X1   g5253(.A1(new_n5638_), .A2(new_n389_), .B(new_n787_), .ZN(new_n5639_));
  AOI21_X1   g5254(.A1(new_n5639_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n5640_));
  OAI21_X1   g5255(.A1(new_n5640_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n5641_));
  AOI21_X1   g5256(.A1(new_n5641_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n5642_));
  OAI21_X1   g5257(.A1(new_n5642_), .A2(new_n900_), .B(new_n908_), .ZN(new_n5643_));
  AOI21_X1   g5258(.A1(new_n5643_), .A2(new_n913_), .B(new_n918_), .ZN(new_n5644_));
  OAI21_X1   g5259(.A1(new_n5644_), .A2(new_n897_), .B(new_n923_), .ZN(new_n5645_));
  AOI21_X1   g5260(.A1(new_n5645_), .A2(new_n894_), .B(new_n929_), .ZN(new_n5646_));
  OAI21_X1   g5261(.A1(new_n5646_), .A2(new_n933_), .B(new_n937_), .ZN(new_n5647_));
  AOI21_X1   g5262(.A1(new_n5647_), .A2(new_n890_), .B(new_n943_), .ZN(new_n5648_));
  OAI21_X1   g5263(.A1(new_n5648_), .A2(new_n886_), .B(new_n948_), .ZN(new_n5649_));
  AOI21_X1   g5264(.A1(new_n5649_), .A2(new_n953_), .B(new_n958_), .ZN(new_n5650_));
  OAI21_X1   g5265(.A1(new_n5650_), .A2(new_n883_), .B(new_n963_), .ZN(new_n5651_));
  AOI21_X1   g5266(.A1(new_n5651_), .A2(new_n880_), .B(new_n969_), .ZN(new_n5652_));
  OAI21_X1   g5267(.A1(new_n5652_), .A2(new_n973_), .B(new_n977_), .ZN(new_n5653_));
  AOI21_X1   g5268(.A1(new_n5653_), .A2(new_n876_), .B(new_n983_), .ZN(new_n5654_));
  OAI21_X1   g5269(.A1(new_n5654_), .A2(new_n872_), .B(new_n988_), .ZN(new_n5655_));
  AOI21_X1   g5270(.A1(new_n5655_), .A2(new_n993_), .B(new_n998_), .ZN(new_n5656_));
  OAI21_X1   g5271(.A1(new_n5656_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n5657_));
  AOI21_X1   g5272(.A1(new_n5657_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n5658_));
  OAI21_X1   g5273(.A1(new_n5658_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n5659_));
  AOI21_X1   g5274(.A1(new_n5659_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n5660_));
  OAI21_X1   g5275(.A1(new_n5660_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n5661_));
  AOI21_X1   g5276(.A1(new_n5661_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n5662_));
  OAI21_X1   g5277(.A1(new_n5662_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n5663_));
  AOI21_X1   g5278(.A1(new_n5663_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n5664_));
  OAI21_X1   g5279(.A1(new_n5664_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n5665_));
  AOI21_X1   g5280(.A1(new_n5665_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n5666_));
  OAI21_X1   g5281(.A1(new_n5666_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n5667_));
  AOI21_X1   g5282(.A1(new_n5667_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n5668_));
  OAI21_X1   g5283(.A1(new_n5668_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n5669_));
  AOI21_X1   g5284(.A1(new_n5669_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n5670_));
  OAI21_X1   g5285(.A1(new_n5670_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n5671_));
  OAI21_X1   g5286(.A1(new_n1099_), .A2(\priority[93] ), .B(\req[93] ), .ZN(new_n5672_));
  AOI21_X1   g5287(.A1(new_n5671_), .A2(new_n834_), .B(new_n5672_), .ZN(\grant[93] ));
  NOR2_X1    g5288(.A1(new_n1212_), .A2(new_n1107_), .ZN(new_n5674_));
  OAI21_X1   g5289(.A1(new_n1112_), .A2(new_n5674_), .B(new_n1117_), .ZN(new_n5675_));
  AOI21_X1   g5290(.A1(new_n5675_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n5676_));
  OAI21_X1   g5291(.A1(new_n5676_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n5677_));
  AOI21_X1   g5292(.A1(new_n5677_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n5678_));
  OAI21_X1   g5293(.A1(new_n5678_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n5679_));
  AOI21_X1   g5294(.A1(new_n5679_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n5680_));
  OAI21_X1   g5295(.A1(new_n5680_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n5681_));
  AOI21_X1   g5296(.A1(new_n5681_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n5682_));
  OAI21_X1   g5297(.A1(new_n5682_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n5683_));
  AOI21_X1   g5298(.A1(new_n5683_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n5684_));
  OAI21_X1   g5299(.A1(new_n5684_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n5685_));
  AOI21_X1   g5300(.A1(new_n5685_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n5686_));
  OAI21_X1   g5301(.A1(new_n5686_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n5687_));
  AOI21_X1   g5302(.A1(new_n5687_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n5688_));
  OAI21_X1   g5303(.A1(new_n5688_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n5689_));
  AOI21_X1   g5304(.A1(new_n5689_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n5690_));
  OAI21_X1   g5305(.A1(new_n5690_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n5691_));
  AOI21_X1   g5306(.A1(new_n5691_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n5692_));
  OAI21_X1   g5307(.A1(new_n5692_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n5693_));
  AOI21_X1   g5308(.A1(new_n5693_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n5694_));
  OAI21_X1   g5309(.A1(new_n5694_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n5695_));
  AOI21_X1   g5310(.A1(new_n5695_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n5696_));
  OAI21_X1   g5311(.A1(new_n5696_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n5697_));
  AOI21_X1   g5312(.A1(new_n5697_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n5698_));
  OAI21_X1   g5313(.A1(new_n5698_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n5699_));
  AOI21_X1   g5314(.A1(new_n5699_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n5700_));
  OAI21_X1   g5315(.A1(new_n5700_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n5701_));
  AOI21_X1   g5316(.A1(new_n5701_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n5702_));
  OAI21_X1   g5317(.A1(new_n5702_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n5703_));
  AOI21_X1   g5318(.A1(new_n5703_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n5704_));
  OAI21_X1   g5319(.A1(new_n5704_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n5705_));
  AOI21_X1   g5320(.A1(new_n5705_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n5706_));
  OAI21_X1   g5321(.A1(new_n5706_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n5707_));
  AOI21_X1   g5322(.A1(new_n5707_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n5708_));
  OAI21_X1   g5323(.A1(new_n5708_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n5709_));
  AOI21_X1   g5324(.A1(new_n5709_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n5710_));
  OAI21_X1   g5325(.A1(new_n5710_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n5711_));
  AOI21_X1   g5326(.A1(new_n5711_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n5712_));
  OAI21_X1   g5327(.A1(new_n5712_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n5713_));
  AOI21_X1   g5328(.A1(new_n5713_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n5714_));
  OAI21_X1   g5329(.A1(new_n5714_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n5715_));
  OAI21_X1   g5330(.A1(new_n414_), .A2(\priority[94] ), .B(\req[94] ), .ZN(new_n5716_));
  AOI21_X1   g5331(.A1(new_n5715_), .A2(new_n1217_), .B(new_n5716_), .ZN(\grant[94] ));
  NOR2_X1    g5332(.A1(new_n728_), .A2(new_n1457_), .ZN(new_n5718_));
  OAI21_X1   g5333(.A1(new_n1462_), .A2(new_n5718_), .B(new_n1466_), .ZN(new_n5719_));
  AOI21_X1   g5334(.A1(new_n5719_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n5720_));
  OAI21_X1   g5335(.A1(new_n5720_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n5721_));
  AOI21_X1   g5336(.A1(new_n5721_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n5722_));
  OAI21_X1   g5337(.A1(new_n5722_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n5723_));
  AOI21_X1   g5338(.A1(new_n5723_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n5724_));
  OAI21_X1   g5339(.A1(new_n5724_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n5725_));
  AOI21_X1   g5340(.A1(new_n5725_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n5726_));
  OAI21_X1   g5341(.A1(new_n5726_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n5727_));
  AOI21_X1   g5342(.A1(new_n5727_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n5728_));
  OAI21_X1   g5343(.A1(new_n5728_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n5729_));
  AOI21_X1   g5344(.A1(new_n5729_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n5730_));
  OAI21_X1   g5345(.A1(new_n5730_), .A2(new_n519_), .B(new_n524_), .ZN(new_n5731_));
  AOI21_X1   g5346(.A1(new_n5731_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n5732_));
  OAI21_X1   g5347(.A1(new_n5732_), .A2(new_n497_), .B(new_n535_), .ZN(new_n5733_));
  AOI21_X1   g5348(.A1(new_n5733_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n5734_));
  OAI21_X1   g5349(.A1(new_n5734_), .A2(new_n492_), .B(new_n550_), .ZN(new_n5735_));
  AOI21_X1   g5350(.A1(new_n5735_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n5736_));
  OAI21_X1   g5351(.A1(new_n5736_), .A2(new_n561_), .B(new_n566_), .ZN(new_n5737_));
  AOI21_X1   g5352(.A1(new_n5737_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n5738_));
  OAI21_X1   g5353(.A1(new_n5738_), .A2(new_n479_), .B(new_n577_), .ZN(new_n5739_));
  AOI21_X1   g5354(.A1(new_n5739_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n5740_));
  OAI21_X1   g5355(.A1(new_n5740_), .A2(new_n474_), .B(new_n592_), .ZN(new_n5741_));
  AOI21_X1   g5356(.A1(new_n5741_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n5742_));
  OAI21_X1   g5357(.A1(new_n5742_), .A2(new_n603_), .B(new_n608_), .ZN(new_n5743_));
  AOI21_X1   g5358(.A1(new_n5743_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n5744_));
  OAI21_X1   g5359(.A1(new_n5744_), .A2(new_n461_), .B(new_n619_), .ZN(new_n5745_));
  AOI21_X1   g5360(.A1(new_n5745_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n5746_));
  OAI21_X1   g5361(.A1(new_n5746_), .A2(new_n456_), .B(new_n634_), .ZN(new_n5747_));
  AOI21_X1   g5362(.A1(new_n5747_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n5748_));
  OAI21_X1   g5363(.A1(new_n5748_), .A2(new_n645_), .B(new_n650_), .ZN(new_n5749_));
  AOI21_X1   g5364(.A1(new_n5749_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n5750_));
  OAI21_X1   g5365(.A1(new_n5750_), .A2(new_n443_), .B(new_n661_), .ZN(new_n5751_));
  AOI21_X1   g5366(.A1(new_n5751_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n5752_));
  OAI21_X1   g5367(.A1(new_n5752_), .A2(new_n438_), .B(new_n676_), .ZN(new_n5753_));
  AOI21_X1   g5368(.A1(new_n5753_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n5754_));
  OAI21_X1   g5369(.A1(new_n5754_), .A2(new_n687_), .B(new_n692_), .ZN(new_n5755_));
  AOI21_X1   g5370(.A1(new_n5755_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n5756_));
  OAI21_X1   g5371(.A1(new_n5756_), .A2(new_n425_), .B(new_n703_), .ZN(new_n5757_));
  AOI21_X1   g5372(.A1(new_n5757_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n5758_));
  OAI21_X1   g5373(.A1(new_n5758_), .A2(new_n420_), .B(new_n718_), .ZN(new_n5759_));
  OAI21_X1   g5374(.A1(new_n721_), .A2(\priority[95] ), .B(\req[95] ), .ZN(new_n5760_));
  AOI21_X1   g5375(.A1(new_n5759_), .A2(new_n1534_), .B(new_n5760_), .ZN(\grant[95] ));
  NOR2_X1    g5376(.A1(new_n1111_), .A2(new_n733_), .ZN(new_n5762_));
  OAI21_X1   g5377(.A1(new_n412_), .A2(new_n5762_), .B(new_n740_), .ZN(new_n5763_));
  AOI21_X1   g5378(.A1(new_n5763_), .A2(new_n408_), .B(new_n746_), .ZN(new_n5764_));
  OAI21_X1   g5379(.A1(new_n5764_), .A2(new_n751_), .B(new_n755_), .ZN(new_n5765_));
  AOI21_X1   g5380(.A1(new_n5765_), .A2(new_n403_), .B(new_n761_), .ZN(new_n5766_));
  OAI21_X1   g5381(.A1(new_n5766_), .A2(new_n398_), .B(new_n766_), .ZN(new_n5767_));
  AOI21_X1   g5382(.A1(new_n5767_), .A2(new_n772_), .B(new_n777_), .ZN(new_n5768_));
  OAI21_X1   g5383(.A1(new_n5768_), .A2(new_n394_), .B(new_n782_), .ZN(new_n5769_));
  AOI21_X1   g5384(.A1(new_n5769_), .A2(new_n390_), .B(new_n788_), .ZN(new_n5770_));
  OAI21_X1   g5385(.A1(new_n5770_), .A2(new_n793_), .B(new_n797_), .ZN(new_n5771_));
  AOI21_X1   g5386(.A1(new_n5771_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n5772_));
  OAI21_X1   g5387(.A1(new_n5772_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n5773_));
  AOI21_X1   g5388(.A1(new_n5773_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n5774_));
  OAI21_X1   g5389(.A1(new_n5774_), .A2(new_n912_), .B(new_n917_), .ZN(new_n5775_));
  AOI21_X1   g5390(.A1(new_n5775_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n5776_));
  OAI21_X1   g5391(.A1(new_n5776_), .A2(new_n893_), .B(new_n928_), .ZN(new_n5777_));
  AOI21_X1   g5392(.A1(new_n5777_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n5778_));
  OAI21_X1   g5393(.A1(new_n5778_), .A2(new_n889_), .B(new_n942_), .ZN(new_n5779_));
  AOI21_X1   g5394(.A1(new_n5779_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n5780_));
  OAI21_X1   g5395(.A1(new_n5780_), .A2(new_n952_), .B(new_n957_), .ZN(new_n5781_));
  AOI21_X1   g5396(.A1(new_n5781_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n5782_));
  OAI21_X1   g5397(.A1(new_n5782_), .A2(new_n879_), .B(new_n968_), .ZN(new_n5783_));
  AOI21_X1   g5398(.A1(new_n5783_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n5784_));
  OAI21_X1   g5399(.A1(new_n5784_), .A2(new_n875_), .B(new_n982_), .ZN(new_n5785_));
  AOI21_X1   g5400(.A1(new_n5785_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n5786_));
  OAI21_X1   g5401(.A1(new_n5786_), .A2(new_n992_), .B(new_n997_), .ZN(new_n5787_));
  AOI21_X1   g5402(.A1(new_n5787_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n5788_));
  OAI21_X1   g5403(.A1(new_n5788_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n5789_));
  AOI21_X1   g5404(.A1(new_n5789_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n5790_));
  OAI21_X1   g5405(.A1(new_n5790_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n5791_));
  AOI21_X1   g5406(.A1(new_n5791_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n5792_));
  OAI21_X1   g5407(.A1(new_n5792_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n5793_));
  AOI21_X1   g5408(.A1(new_n5793_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n5794_));
  OAI21_X1   g5409(.A1(new_n5794_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n5795_));
  AOI21_X1   g5410(.A1(new_n5795_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n5796_));
  OAI21_X1   g5411(.A1(new_n5796_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n5797_));
  AOI21_X1   g5412(.A1(new_n5797_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n5798_));
  OAI21_X1   g5413(.A1(new_n5798_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n5799_));
  AOI21_X1   g5414(.A1(new_n5799_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n5800_));
  OAI21_X1   g5415(.A1(new_n5800_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n5801_));
  AOI21_X1   g5416(.A1(new_n5801_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n5802_));
  OAI21_X1   g5417(.A1(new_n5802_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n5803_));
  OAI21_X1   g5418(.A1(new_n1105_), .A2(\priority[96] ), .B(\req[96] ), .ZN(new_n5804_));
  AOI21_X1   g5419(.A1(new_n5803_), .A2(new_n1624_), .B(new_n5804_), .ZN(\grant[96] ));
  NOR2_X1    g5420(.A1(new_n1461_), .A2(new_n1116_), .ZN(new_n5806_));
  OAI21_X1   g5421(.A1(new_n827_), .A2(new_n5806_), .B(new_n1123_), .ZN(new_n5807_));
  AOI21_X1   g5422(.A1(new_n5807_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n5808_));
  OAI21_X1   g5423(.A1(new_n5808_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n5809_));
  AOI21_X1   g5424(.A1(new_n5809_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n5810_));
  OAI21_X1   g5425(.A1(new_n5810_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n5811_));
  AOI21_X1   g5426(.A1(new_n5811_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n5812_));
  OAI21_X1   g5427(.A1(new_n5812_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n5813_));
  AOI21_X1   g5428(.A1(new_n5813_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n5814_));
  OAI21_X1   g5429(.A1(new_n5814_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n5815_));
  AOI21_X1   g5430(.A1(new_n5815_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n5816_));
  OAI21_X1   g5431(.A1(new_n5816_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n5817_));
  AOI21_X1   g5432(.A1(new_n5817_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n5818_));
  OAI21_X1   g5433(.A1(new_n5818_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n5819_));
  AOI21_X1   g5434(.A1(new_n5819_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n5820_));
  OAI21_X1   g5435(.A1(new_n5820_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n5821_));
  AOI21_X1   g5436(.A1(new_n5821_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n5822_));
  OAI21_X1   g5437(.A1(new_n5822_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n5823_));
  AOI21_X1   g5438(.A1(new_n5823_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n5824_));
  OAI21_X1   g5439(.A1(new_n5824_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n5825_));
  AOI21_X1   g5440(.A1(new_n5825_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n5826_));
  OAI21_X1   g5441(.A1(new_n5826_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n5827_));
  AOI21_X1   g5442(.A1(new_n5827_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n5828_));
  OAI21_X1   g5443(.A1(new_n5828_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n5829_));
  AOI21_X1   g5444(.A1(new_n5829_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n5830_));
  OAI21_X1   g5445(.A1(new_n5830_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n5831_));
  AOI21_X1   g5446(.A1(new_n5831_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n5832_));
  OAI21_X1   g5447(.A1(new_n5832_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n5833_));
  AOI21_X1   g5448(.A1(new_n5833_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n5834_));
  OAI21_X1   g5449(.A1(new_n5834_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n5835_));
  AOI21_X1   g5450(.A1(new_n5835_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n5836_));
  OAI21_X1   g5451(.A1(new_n5836_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n5837_));
  AOI21_X1   g5452(.A1(new_n5837_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n5838_));
  OAI21_X1   g5453(.A1(new_n5838_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n5839_));
  AOI21_X1   g5454(.A1(new_n5839_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n5840_));
  OAI21_X1   g5455(.A1(new_n5840_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n5841_));
  AOI21_X1   g5456(.A1(new_n5841_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n5842_));
  OAI21_X1   g5457(.A1(new_n5842_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n5843_));
  AOI21_X1   g5458(.A1(new_n5843_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n5844_));
  OAI21_X1   g5459(.A1(new_n5844_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n5845_));
  AOI21_X1   g5460(.A1(new_n5845_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n5846_));
  OAI21_X1   g5461(.A1(new_n5846_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n5847_));
  OAI21_X1   g5462(.A1(new_n727_), .A2(\priority[97] ), .B(\req[97] ), .ZN(new_n5848_));
  AOI21_X1   g5463(.A1(new_n5847_), .A2(new_n1712_), .B(new_n5848_), .ZN(\grant[97] ));
  NOR2_X1    g5464(.A1(new_n411_), .A2(new_n1465_), .ZN(new_n5850_));
  OAI21_X1   g5465(.A1(new_n1210_), .A2(new_n5850_), .B(new_n1471_), .ZN(new_n5851_));
  AOI21_X1   g5466(.A1(new_n5851_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n5852_));
  OAI21_X1   g5467(.A1(new_n5852_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n5853_));
  AOI21_X1   g5468(.A1(new_n5853_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n5854_));
  OAI21_X1   g5469(.A1(new_n5854_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n5855_));
  AOI21_X1   g5470(.A1(new_n5855_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n5856_));
  OAI21_X1   g5471(.A1(new_n5856_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n5857_));
  AOI21_X1   g5472(.A1(new_n5857_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n5858_));
  OAI21_X1   g5473(.A1(new_n5858_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n5859_));
  AOI21_X1   g5474(.A1(new_n5859_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n5860_));
  OAI21_X1   g5475(.A1(new_n5860_), .A2(new_n506_), .B(new_n514_), .ZN(new_n5861_));
  AOI21_X1   g5476(.A1(new_n5861_), .A2(new_n520_), .B(new_n525_), .ZN(new_n5862_));
  OAI21_X1   g5477(.A1(new_n5862_), .A2(new_n502_), .B(new_n530_), .ZN(new_n5863_));
  AOI21_X1   g5478(.A1(new_n5863_), .A2(new_n498_), .B(new_n536_), .ZN(new_n5864_));
  OAI21_X1   g5479(.A1(new_n5864_), .A2(new_n541_), .B(new_n545_), .ZN(new_n5865_));
  AOI21_X1   g5480(.A1(new_n5865_), .A2(new_n493_), .B(new_n551_), .ZN(new_n5866_));
  OAI21_X1   g5481(.A1(new_n5866_), .A2(new_n488_), .B(new_n556_), .ZN(new_n5867_));
  AOI21_X1   g5482(.A1(new_n5867_), .A2(new_n562_), .B(new_n567_), .ZN(new_n5868_));
  OAI21_X1   g5483(.A1(new_n5868_), .A2(new_n484_), .B(new_n572_), .ZN(new_n5869_));
  AOI21_X1   g5484(.A1(new_n5869_), .A2(new_n480_), .B(new_n578_), .ZN(new_n5870_));
  OAI21_X1   g5485(.A1(new_n5870_), .A2(new_n583_), .B(new_n587_), .ZN(new_n5871_));
  AOI21_X1   g5486(.A1(new_n5871_), .A2(new_n475_), .B(new_n593_), .ZN(new_n5872_));
  OAI21_X1   g5487(.A1(new_n5872_), .A2(new_n470_), .B(new_n598_), .ZN(new_n5873_));
  AOI21_X1   g5488(.A1(new_n5873_), .A2(new_n604_), .B(new_n609_), .ZN(new_n5874_));
  OAI21_X1   g5489(.A1(new_n5874_), .A2(new_n466_), .B(new_n614_), .ZN(new_n5875_));
  AOI21_X1   g5490(.A1(new_n5875_), .A2(new_n462_), .B(new_n620_), .ZN(new_n5876_));
  OAI21_X1   g5491(.A1(new_n5876_), .A2(new_n625_), .B(new_n629_), .ZN(new_n5877_));
  AOI21_X1   g5492(.A1(new_n5877_), .A2(new_n457_), .B(new_n635_), .ZN(new_n5878_));
  OAI21_X1   g5493(.A1(new_n5878_), .A2(new_n452_), .B(new_n640_), .ZN(new_n5879_));
  AOI21_X1   g5494(.A1(new_n5879_), .A2(new_n646_), .B(new_n651_), .ZN(new_n5880_));
  OAI21_X1   g5495(.A1(new_n5880_), .A2(new_n448_), .B(new_n656_), .ZN(new_n5881_));
  AOI21_X1   g5496(.A1(new_n5881_), .A2(new_n444_), .B(new_n662_), .ZN(new_n5882_));
  OAI21_X1   g5497(.A1(new_n5882_), .A2(new_n667_), .B(new_n671_), .ZN(new_n5883_));
  AOI21_X1   g5498(.A1(new_n5883_), .A2(new_n439_), .B(new_n677_), .ZN(new_n5884_));
  OAI21_X1   g5499(.A1(new_n5884_), .A2(new_n434_), .B(new_n682_), .ZN(new_n5885_));
  AOI21_X1   g5500(.A1(new_n5885_), .A2(new_n688_), .B(new_n693_), .ZN(new_n5886_));
  OAI21_X1   g5501(.A1(new_n5886_), .A2(new_n430_), .B(new_n698_), .ZN(new_n5887_));
  AOI21_X1   g5502(.A1(new_n5887_), .A2(new_n426_), .B(new_n704_), .ZN(new_n5888_));
  OAI21_X1   g5503(.A1(new_n5888_), .A2(new_n709_), .B(new_n713_), .ZN(new_n5889_));
  AOI21_X1   g5504(.A1(new_n5889_), .A2(new_n421_), .B(new_n719_), .ZN(new_n5890_));
  OAI21_X1   g5505(.A1(new_n5890_), .A2(new_n416_), .B(new_n724_), .ZN(new_n5891_));
  OAI21_X1   g5506(.A1(new_n731_), .A2(\priority[98] ), .B(\req[98] ), .ZN(new_n5892_));
  AOI21_X1   g5507(.A1(new_n5891_), .A2(new_n730_), .B(new_n5892_), .ZN(\grant[98] ));
  NOR2_X1    g5508(.A1(new_n826_), .A2(new_n739_), .ZN(new_n5894_));
  OAI21_X1   g5509(.A1(new_n407_), .A2(new_n5894_), .B(new_n745_), .ZN(new_n5895_));
  AOI21_X1   g5510(.A1(new_n5895_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n5896_));
  OAI21_X1   g5511(.A1(new_n5896_), .A2(new_n402_), .B(new_n760_), .ZN(new_n5897_));
  AOI21_X1   g5512(.A1(new_n5897_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n5898_));
  OAI21_X1   g5513(.A1(new_n5898_), .A2(new_n771_), .B(new_n776_), .ZN(new_n5899_));
  AOI21_X1   g5514(.A1(new_n5899_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n5900_));
  OAI21_X1   g5515(.A1(new_n5900_), .A2(new_n389_), .B(new_n787_), .ZN(new_n5901_));
  AOI21_X1   g5516(.A1(new_n5901_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n5902_));
  OAI21_X1   g5517(.A1(new_n5902_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n5903_));
  AOI21_X1   g5518(.A1(new_n5903_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n5904_));
  OAI21_X1   g5519(.A1(new_n5904_), .A2(new_n900_), .B(new_n908_), .ZN(new_n5905_));
  AOI21_X1   g5520(.A1(new_n5905_), .A2(new_n913_), .B(new_n918_), .ZN(new_n5906_));
  OAI21_X1   g5521(.A1(new_n5906_), .A2(new_n897_), .B(new_n923_), .ZN(new_n5907_));
  AOI21_X1   g5522(.A1(new_n5907_), .A2(new_n894_), .B(new_n929_), .ZN(new_n5908_));
  OAI21_X1   g5523(.A1(new_n5908_), .A2(new_n933_), .B(new_n937_), .ZN(new_n5909_));
  AOI21_X1   g5524(.A1(new_n5909_), .A2(new_n890_), .B(new_n943_), .ZN(new_n5910_));
  OAI21_X1   g5525(.A1(new_n5910_), .A2(new_n886_), .B(new_n948_), .ZN(new_n5911_));
  AOI21_X1   g5526(.A1(new_n5911_), .A2(new_n953_), .B(new_n958_), .ZN(new_n5912_));
  OAI21_X1   g5527(.A1(new_n5912_), .A2(new_n883_), .B(new_n963_), .ZN(new_n5913_));
  AOI21_X1   g5528(.A1(new_n5913_), .A2(new_n880_), .B(new_n969_), .ZN(new_n5914_));
  OAI21_X1   g5529(.A1(new_n5914_), .A2(new_n973_), .B(new_n977_), .ZN(new_n5915_));
  AOI21_X1   g5530(.A1(new_n5915_), .A2(new_n876_), .B(new_n983_), .ZN(new_n5916_));
  OAI21_X1   g5531(.A1(new_n5916_), .A2(new_n872_), .B(new_n988_), .ZN(new_n5917_));
  AOI21_X1   g5532(.A1(new_n5917_), .A2(new_n993_), .B(new_n998_), .ZN(new_n5918_));
  OAI21_X1   g5533(.A1(new_n5918_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n5919_));
  AOI21_X1   g5534(.A1(new_n5919_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n5920_));
  OAI21_X1   g5535(.A1(new_n5920_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n5921_));
  AOI21_X1   g5536(.A1(new_n5921_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n5922_));
  OAI21_X1   g5537(.A1(new_n5922_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n5923_));
  AOI21_X1   g5538(.A1(new_n5923_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n5924_));
  OAI21_X1   g5539(.A1(new_n5924_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n5925_));
  AOI21_X1   g5540(.A1(new_n5925_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n5926_));
  OAI21_X1   g5541(.A1(new_n5926_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n5927_));
  AOI21_X1   g5542(.A1(new_n5927_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n5928_));
  OAI21_X1   g5543(.A1(new_n5928_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n5929_));
  AOI21_X1   g5544(.A1(new_n5929_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n5930_));
  OAI21_X1   g5545(.A1(new_n5930_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n5931_));
  AOI21_X1   g5546(.A1(new_n5931_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n5932_));
  OAI21_X1   g5547(.A1(new_n5932_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n5933_));
  AOI21_X1   g5548(.A1(new_n5933_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n5934_));
  OAI21_X1   g5549(.A1(new_n5934_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n5935_));
  OAI21_X1   g5550(.A1(new_n1114_), .A2(\priority[99] ), .B(\req[99] ), .ZN(new_n5936_));
  AOI21_X1   g5551(.A1(new_n5935_), .A2(new_n1113_), .B(new_n5936_), .ZN(\grant[99] ));
  NOR2_X1    g5552(.A1(new_n1209_), .A2(new_n1122_), .ZN(new_n5938_));
  OAI21_X1   g5553(.A1(new_n823_), .A2(new_n5938_), .B(new_n1128_), .ZN(new_n5939_));
  AOI21_X1   g5554(.A1(new_n5939_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n5940_));
  OAI21_X1   g5555(.A1(new_n5940_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n5941_));
  AOI21_X1   g5556(.A1(new_n5941_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n5942_));
  OAI21_X1   g5557(.A1(new_n5942_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n5943_));
  AOI21_X1   g5558(.A1(new_n5943_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n5944_));
  OAI21_X1   g5559(.A1(new_n5944_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n5945_));
  AOI21_X1   g5560(.A1(new_n5945_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n5946_));
  OAI21_X1   g5561(.A1(new_n5946_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n5947_));
  AOI21_X1   g5562(.A1(new_n5947_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n5948_));
  OAI21_X1   g5563(.A1(new_n5948_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n5949_));
  AOI21_X1   g5564(.A1(new_n5949_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n5950_));
  OAI21_X1   g5565(.A1(new_n5950_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n5951_));
  AOI21_X1   g5566(.A1(new_n5951_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n5952_));
  OAI21_X1   g5567(.A1(new_n5952_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n5953_));
  AOI21_X1   g5568(.A1(new_n5953_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n5954_));
  OAI21_X1   g5569(.A1(new_n5954_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n5955_));
  AOI21_X1   g5570(.A1(new_n5955_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n5956_));
  OAI21_X1   g5571(.A1(new_n5956_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n5957_));
  AOI21_X1   g5572(.A1(new_n5957_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n5958_));
  OAI21_X1   g5573(.A1(new_n5958_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n5959_));
  AOI21_X1   g5574(.A1(new_n5959_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n5960_));
  OAI21_X1   g5575(.A1(new_n5960_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n5961_));
  AOI21_X1   g5576(.A1(new_n5961_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n5962_));
  OAI21_X1   g5577(.A1(new_n5962_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n5963_));
  AOI21_X1   g5578(.A1(new_n5963_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n5964_));
  OAI21_X1   g5579(.A1(new_n5964_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n5965_));
  AOI21_X1   g5580(.A1(new_n5965_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n5966_));
  OAI21_X1   g5581(.A1(new_n5966_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n5967_));
  AOI21_X1   g5582(.A1(new_n5967_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n5968_));
  OAI21_X1   g5583(.A1(new_n5968_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n5969_));
  AOI21_X1   g5584(.A1(new_n5969_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n5970_));
  OAI21_X1   g5585(.A1(new_n5970_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n5971_));
  AOI21_X1   g5586(.A1(new_n5971_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n5972_));
  OAI21_X1   g5587(.A1(new_n5972_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n5973_));
  AOI21_X1   g5588(.A1(new_n5973_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n5974_));
  OAI21_X1   g5589(.A1(new_n5974_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n5975_));
  AOI21_X1   g5590(.A1(new_n5975_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n5976_));
  OAI21_X1   g5591(.A1(new_n5976_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n5977_));
  AOI21_X1   g5592(.A1(new_n5977_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n5978_));
  OAI21_X1   g5593(.A1(new_n5978_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n5979_));
  OAI21_X1   g5594(.A1(new_n410_), .A2(\priority[100] ), .B(\req[100] ), .ZN(new_n5980_));
  AOI21_X1   g5595(.A1(new_n5979_), .A2(new_n1463_), .B(new_n5980_), .ZN(\grant[100] ));
  NOR2_X1    g5596(.A1(new_n406_), .A2(new_n1470_), .ZN(new_n5982_));
  OAI21_X1   g5597(.A1(new_n1206_), .A2(new_n5982_), .B(new_n1475_), .ZN(new_n5983_));
  AOI21_X1   g5598(.A1(new_n5983_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n5984_));
  OAI21_X1   g5599(.A1(new_n5984_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n5985_));
  AOI21_X1   g5600(.A1(new_n5985_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n5986_));
  OAI21_X1   g5601(.A1(new_n5986_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n5987_));
  AOI21_X1   g5602(.A1(new_n5987_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n5988_));
  OAI21_X1   g5603(.A1(new_n5988_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n5989_));
  AOI21_X1   g5604(.A1(new_n5989_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n5990_));
  OAI21_X1   g5605(.A1(new_n5990_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n5991_));
  AOI21_X1   g5606(.A1(new_n5991_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n5992_));
  OAI21_X1   g5607(.A1(new_n5992_), .A2(new_n519_), .B(new_n524_), .ZN(new_n5993_));
  AOI21_X1   g5608(.A1(new_n5993_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n5994_));
  OAI21_X1   g5609(.A1(new_n5994_), .A2(new_n497_), .B(new_n535_), .ZN(new_n5995_));
  AOI21_X1   g5610(.A1(new_n5995_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n5996_));
  OAI21_X1   g5611(.A1(new_n5996_), .A2(new_n492_), .B(new_n550_), .ZN(new_n5997_));
  AOI21_X1   g5612(.A1(new_n5997_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n5998_));
  OAI21_X1   g5613(.A1(new_n5998_), .A2(new_n561_), .B(new_n566_), .ZN(new_n5999_));
  AOI21_X1   g5614(.A1(new_n5999_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n6000_));
  OAI21_X1   g5615(.A1(new_n6000_), .A2(new_n479_), .B(new_n577_), .ZN(new_n6001_));
  AOI21_X1   g5616(.A1(new_n6001_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n6002_));
  OAI21_X1   g5617(.A1(new_n6002_), .A2(new_n474_), .B(new_n592_), .ZN(new_n6003_));
  AOI21_X1   g5618(.A1(new_n6003_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n6004_));
  OAI21_X1   g5619(.A1(new_n6004_), .A2(new_n603_), .B(new_n608_), .ZN(new_n6005_));
  AOI21_X1   g5620(.A1(new_n6005_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n6006_));
  OAI21_X1   g5621(.A1(new_n6006_), .A2(new_n461_), .B(new_n619_), .ZN(new_n6007_));
  AOI21_X1   g5622(.A1(new_n6007_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n6008_));
  OAI21_X1   g5623(.A1(new_n6008_), .A2(new_n456_), .B(new_n634_), .ZN(new_n6009_));
  AOI21_X1   g5624(.A1(new_n6009_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n6010_));
  OAI21_X1   g5625(.A1(new_n6010_), .A2(new_n645_), .B(new_n650_), .ZN(new_n6011_));
  AOI21_X1   g5626(.A1(new_n6011_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n6012_));
  OAI21_X1   g5627(.A1(new_n6012_), .A2(new_n443_), .B(new_n661_), .ZN(new_n6013_));
  AOI21_X1   g5628(.A1(new_n6013_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n6014_));
  OAI21_X1   g5629(.A1(new_n6014_), .A2(new_n438_), .B(new_n676_), .ZN(new_n6015_));
  AOI21_X1   g5630(.A1(new_n6015_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n6016_));
  OAI21_X1   g5631(.A1(new_n6016_), .A2(new_n687_), .B(new_n692_), .ZN(new_n6017_));
  AOI21_X1   g5632(.A1(new_n6017_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n6018_));
  OAI21_X1   g5633(.A1(new_n6018_), .A2(new_n425_), .B(new_n703_), .ZN(new_n6019_));
  AOI21_X1   g5634(.A1(new_n6019_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n6020_));
  OAI21_X1   g5635(.A1(new_n6020_), .A2(new_n420_), .B(new_n718_), .ZN(new_n6021_));
  AOI21_X1   g5636(.A1(new_n6021_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n6022_));
  OAI21_X1   g5637(.A1(new_n6022_), .A2(new_n729_), .B(new_n734_), .ZN(new_n6023_));
  OAI21_X1   g5638(.A1(new_n737_), .A2(\priority[101] ), .B(\req[101] ), .ZN(new_n6024_));
  AOI21_X1   g5639(.A1(new_n6023_), .A2(new_n1532_), .B(new_n6024_), .ZN(\grant[101] ));
  NOR2_X1    g5640(.A1(new_n822_), .A2(new_n744_), .ZN(new_n6026_));
  OAI21_X1   g5641(.A1(new_n751_), .A2(new_n6026_), .B(new_n755_), .ZN(new_n6027_));
  AOI21_X1   g5642(.A1(new_n6027_), .A2(new_n403_), .B(new_n761_), .ZN(new_n6028_));
  OAI21_X1   g5643(.A1(new_n6028_), .A2(new_n398_), .B(new_n766_), .ZN(new_n6029_));
  AOI21_X1   g5644(.A1(new_n6029_), .A2(new_n772_), .B(new_n777_), .ZN(new_n6030_));
  OAI21_X1   g5645(.A1(new_n6030_), .A2(new_n394_), .B(new_n782_), .ZN(new_n6031_));
  AOI21_X1   g5646(.A1(new_n6031_), .A2(new_n390_), .B(new_n788_), .ZN(new_n6032_));
  OAI21_X1   g5647(.A1(new_n6032_), .A2(new_n793_), .B(new_n797_), .ZN(new_n6033_));
  AOI21_X1   g5648(.A1(new_n6033_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n6034_));
  OAI21_X1   g5649(.A1(new_n6034_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n6035_));
  AOI21_X1   g5650(.A1(new_n6035_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n6036_));
  OAI21_X1   g5651(.A1(new_n6036_), .A2(new_n912_), .B(new_n917_), .ZN(new_n6037_));
  AOI21_X1   g5652(.A1(new_n6037_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n6038_));
  OAI21_X1   g5653(.A1(new_n6038_), .A2(new_n893_), .B(new_n928_), .ZN(new_n6039_));
  AOI21_X1   g5654(.A1(new_n6039_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n6040_));
  OAI21_X1   g5655(.A1(new_n6040_), .A2(new_n889_), .B(new_n942_), .ZN(new_n6041_));
  AOI21_X1   g5656(.A1(new_n6041_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n6042_));
  OAI21_X1   g5657(.A1(new_n6042_), .A2(new_n952_), .B(new_n957_), .ZN(new_n6043_));
  AOI21_X1   g5658(.A1(new_n6043_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n6044_));
  OAI21_X1   g5659(.A1(new_n6044_), .A2(new_n879_), .B(new_n968_), .ZN(new_n6045_));
  AOI21_X1   g5660(.A1(new_n6045_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n6046_));
  OAI21_X1   g5661(.A1(new_n6046_), .A2(new_n875_), .B(new_n982_), .ZN(new_n6047_));
  AOI21_X1   g5662(.A1(new_n6047_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n6048_));
  OAI21_X1   g5663(.A1(new_n6048_), .A2(new_n992_), .B(new_n997_), .ZN(new_n6049_));
  AOI21_X1   g5664(.A1(new_n6049_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n6050_));
  OAI21_X1   g5665(.A1(new_n6050_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n6051_));
  AOI21_X1   g5666(.A1(new_n6051_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n6052_));
  OAI21_X1   g5667(.A1(new_n6052_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n6053_));
  AOI21_X1   g5668(.A1(new_n6053_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n6054_));
  OAI21_X1   g5669(.A1(new_n6054_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n6055_));
  AOI21_X1   g5670(.A1(new_n6055_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n6056_));
  OAI21_X1   g5671(.A1(new_n6056_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n6057_));
  AOI21_X1   g5672(.A1(new_n6057_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n6058_));
  OAI21_X1   g5673(.A1(new_n6058_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n6059_));
  AOI21_X1   g5674(.A1(new_n6059_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n6060_));
  OAI21_X1   g5675(.A1(new_n6060_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n6061_));
  AOI21_X1   g5676(.A1(new_n6061_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n6062_));
  OAI21_X1   g5677(.A1(new_n6062_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n6063_));
  AOI21_X1   g5678(.A1(new_n6063_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n6064_));
  OAI21_X1   g5679(.A1(new_n6064_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n6065_));
  AOI21_X1   g5680(.A1(new_n6065_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n6066_));
  OAI21_X1   g5681(.A1(new_n6066_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n6067_));
  OAI21_X1   g5682(.A1(new_n1120_), .A2(\priority[102] ), .B(\req[102] ), .ZN(new_n6068_));
  AOI21_X1   g5683(.A1(new_n6067_), .A2(new_n1622_), .B(new_n6068_), .ZN(\grant[102] ));
  NOR2_X1    g5684(.A1(new_n1205_), .A2(new_n1127_), .ZN(new_n6070_));
  OAI21_X1   g5685(.A1(new_n1133_), .A2(new_n6070_), .B(new_n1137_), .ZN(new_n6071_));
  AOI21_X1   g5686(.A1(new_n6071_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n6072_));
  OAI21_X1   g5687(.A1(new_n6072_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n6073_));
  AOI21_X1   g5688(.A1(new_n6073_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n6074_));
  OAI21_X1   g5689(.A1(new_n6074_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n6075_));
  AOI21_X1   g5690(.A1(new_n6075_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n6076_));
  OAI21_X1   g5691(.A1(new_n6076_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n6077_));
  AOI21_X1   g5692(.A1(new_n6077_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n6078_));
  OAI21_X1   g5693(.A1(new_n6078_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n6079_));
  AOI21_X1   g5694(.A1(new_n6079_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n6080_));
  OAI21_X1   g5695(.A1(new_n6080_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n6081_));
  AOI21_X1   g5696(.A1(new_n6081_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n6082_));
  OAI21_X1   g5697(.A1(new_n6082_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n6083_));
  AOI21_X1   g5698(.A1(new_n6083_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n6084_));
  OAI21_X1   g5699(.A1(new_n6084_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n6085_));
  AOI21_X1   g5700(.A1(new_n6085_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n6086_));
  OAI21_X1   g5701(.A1(new_n6086_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n6087_));
  AOI21_X1   g5702(.A1(new_n6087_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n6088_));
  OAI21_X1   g5703(.A1(new_n6088_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n6089_));
  AOI21_X1   g5704(.A1(new_n6089_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n6090_));
  OAI21_X1   g5705(.A1(new_n6090_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n6091_));
  AOI21_X1   g5706(.A1(new_n6091_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n6092_));
  OAI21_X1   g5707(.A1(new_n6092_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n6093_));
  AOI21_X1   g5708(.A1(new_n6093_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n6094_));
  OAI21_X1   g5709(.A1(new_n6094_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n6095_));
  AOI21_X1   g5710(.A1(new_n6095_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n6096_));
  OAI21_X1   g5711(.A1(new_n6096_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n6097_));
  AOI21_X1   g5712(.A1(new_n6097_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n6098_));
  OAI21_X1   g5713(.A1(new_n6098_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n6099_));
  AOI21_X1   g5714(.A1(new_n6099_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n6100_));
  OAI21_X1   g5715(.A1(new_n6100_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n6101_));
  AOI21_X1   g5716(.A1(new_n6101_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n6102_));
  OAI21_X1   g5717(.A1(new_n6102_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n6103_));
  AOI21_X1   g5718(.A1(new_n6103_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n6104_));
  OAI21_X1   g5719(.A1(new_n6104_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n6105_));
  AOI21_X1   g5720(.A1(new_n6105_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n6106_));
  OAI21_X1   g5721(.A1(new_n6106_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n6107_));
  AOI21_X1   g5722(.A1(new_n6107_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n6108_));
  OAI21_X1   g5723(.A1(new_n6108_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n6109_));
  AOI21_X1   g5724(.A1(new_n6109_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n6110_));
  OAI21_X1   g5725(.A1(new_n6110_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n6111_));
  OAI21_X1   g5726(.A1(new_n405_), .A2(\priority[103] ), .B(\req[103] ), .ZN(new_n6112_));
  AOI21_X1   g5727(.A1(new_n6111_), .A2(new_n1710_), .B(new_n6112_), .ZN(\grant[103] ));
  NOR2_X1    g5728(.A1(new_n750_), .A2(new_n1474_), .ZN(new_n6114_));
  OAI21_X1   g5729(.A1(new_n1480_), .A2(new_n6114_), .B(new_n1483_), .ZN(new_n6115_));
  AOI21_X1   g5730(.A1(new_n6115_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n6116_));
  OAI21_X1   g5731(.A1(new_n6116_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n6117_));
  AOI21_X1   g5732(.A1(new_n6117_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n6118_));
  OAI21_X1   g5733(.A1(new_n6118_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n6119_));
  AOI21_X1   g5734(.A1(new_n6119_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n6120_));
  OAI21_X1   g5735(.A1(new_n6120_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n6121_));
  AOI21_X1   g5736(.A1(new_n6121_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n6122_));
  OAI21_X1   g5737(.A1(new_n6122_), .A2(new_n506_), .B(new_n514_), .ZN(new_n6123_));
  AOI21_X1   g5738(.A1(new_n6123_), .A2(new_n520_), .B(new_n525_), .ZN(new_n6124_));
  OAI21_X1   g5739(.A1(new_n6124_), .A2(new_n502_), .B(new_n530_), .ZN(new_n6125_));
  AOI21_X1   g5740(.A1(new_n6125_), .A2(new_n498_), .B(new_n536_), .ZN(new_n6126_));
  OAI21_X1   g5741(.A1(new_n6126_), .A2(new_n541_), .B(new_n545_), .ZN(new_n6127_));
  AOI21_X1   g5742(.A1(new_n6127_), .A2(new_n493_), .B(new_n551_), .ZN(new_n6128_));
  OAI21_X1   g5743(.A1(new_n6128_), .A2(new_n488_), .B(new_n556_), .ZN(new_n6129_));
  AOI21_X1   g5744(.A1(new_n6129_), .A2(new_n562_), .B(new_n567_), .ZN(new_n6130_));
  OAI21_X1   g5745(.A1(new_n6130_), .A2(new_n484_), .B(new_n572_), .ZN(new_n6131_));
  AOI21_X1   g5746(.A1(new_n6131_), .A2(new_n480_), .B(new_n578_), .ZN(new_n6132_));
  OAI21_X1   g5747(.A1(new_n6132_), .A2(new_n583_), .B(new_n587_), .ZN(new_n6133_));
  AOI21_X1   g5748(.A1(new_n6133_), .A2(new_n475_), .B(new_n593_), .ZN(new_n6134_));
  OAI21_X1   g5749(.A1(new_n6134_), .A2(new_n470_), .B(new_n598_), .ZN(new_n6135_));
  AOI21_X1   g5750(.A1(new_n6135_), .A2(new_n604_), .B(new_n609_), .ZN(new_n6136_));
  OAI21_X1   g5751(.A1(new_n6136_), .A2(new_n466_), .B(new_n614_), .ZN(new_n6137_));
  AOI21_X1   g5752(.A1(new_n6137_), .A2(new_n462_), .B(new_n620_), .ZN(new_n6138_));
  OAI21_X1   g5753(.A1(new_n6138_), .A2(new_n625_), .B(new_n629_), .ZN(new_n6139_));
  AOI21_X1   g5754(.A1(new_n6139_), .A2(new_n457_), .B(new_n635_), .ZN(new_n6140_));
  OAI21_X1   g5755(.A1(new_n6140_), .A2(new_n452_), .B(new_n640_), .ZN(new_n6141_));
  AOI21_X1   g5756(.A1(new_n6141_), .A2(new_n646_), .B(new_n651_), .ZN(new_n6142_));
  OAI21_X1   g5757(.A1(new_n6142_), .A2(new_n448_), .B(new_n656_), .ZN(new_n6143_));
  AOI21_X1   g5758(.A1(new_n6143_), .A2(new_n444_), .B(new_n662_), .ZN(new_n6144_));
  OAI21_X1   g5759(.A1(new_n6144_), .A2(new_n667_), .B(new_n671_), .ZN(new_n6145_));
  AOI21_X1   g5760(.A1(new_n6145_), .A2(new_n439_), .B(new_n677_), .ZN(new_n6146_));
  OAI21_X1   g5761(.A1(new_n6146_), .A2(new_n434_), .B(new_n682_), .ZN(new_n6147_));
  AOI21_X1   g5762(.A1(new_n6147_), .A2(new_n688_), .B(new_n693_), .ZN(new_n6148_));
  OAI21_X1   g5763(.A1(new_n6148_), .A2(new_n430_), .B(new_n698_), .ZN(new_n6149_));
  AOI21_X1   g5764(.A1(new_n6149_), .A2(new_n426_), .B(new_n704_), .ZN(new_n6150_));
  OAI21_X1   g5765(.A1(new_n6150_), .A2(new_n709_), .B(new_n713_), .ZN(new_n6151_));
  AOI21_X1   g5766(.A1(new_n6151_), .A2(new_n421_), .B(new_n719_), .ZN(new_n6152_));
  OAI21_X1   g5767(.A1(new_n6152_), .A2(new_n416_), .B(new_n724_), .ZN(new_n6153_));
  AOI21_X1   g5768(.A1(new_n6153_), .A2(new_n730_), .B(new_n735_), .ZN(new_n6154_));
  OAI21_X1   g5769(.A1(new_n6154_), .A2(new_n412_), .B(new_n740_), .ZN(new_n6155_));
  OAI21_X1   g5770(.A1(new_n742_), .A2(\priority[104] ), .B(\req[104] ), .ZN(new_n6156_));
  AOI21_X1   g5771(.A1(new_n6155_), .A2(new_n408_), .B(new_n6156_), .ZN(\grant[104] ));
  NOR2_X1    g5772(.A1(new_n1132_), .A2(new_n754_), .ZN(new_n6158_));
  OAI21_X1   g5773(.A1(new_n402_), .A2(new_n6158_), .B(new_n760_), .ZN(new_n6159_));
  AOI21_X1   g5774(.A1(new_n6159_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n6160_));
  OAI21_X1   g5775(.A1(new_n6160_), .A2(new_n771_), .B(new_n776_), .ZN(new_n6161_));
  AOI21_X1   g5776(.A1(new_n6161_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n6162_));
  OAI21_X1   g5777(.A1(new_n6162_), .A2(new_n389_), .B(new_n787_), .ZN(new_n6163_));
  AOI21_X1   g5778(.A1(new_n6163_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n6164_));
  OAI21_X1   g5779(.A1(new_n6164_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n6165_));
  AOI21_X1   g5780(.A1(new_n6165_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n6166_));
  OAI21_X1   g5781(.A1(new_n6166_), .A2(new_n900_), .B(new_n908_), .ZN(new_n6167_));
  AOI21_X1   g5782(.A1(new_n6167_), .A2(new_n913_), .B(new_n918_), .ZN(new_n6168_));
  OAI21_X1   g5783(.A1(new_n6168_), .A2(new_n897_), .B(new_n923_), .ZN(new_n6169_));
  AOI21_X1   g5784(.A1(new_n6169_), .A2(new_n894_), .B(new_n929_), .ZN(new_n6170_));
  OAI21_X1   g5785(.A1(new_n6170_), .A2(new_n933_), .B(new_n937_), .ZN(new_n6171_));
  AOI21_X1   g5786(.A1(new_n6171_), .A2(new_n890_), .B(new_n943_), .ZN(new_n6172_));
  OAI21_X1   g5787(.A1(new_n6172_), .A2(new_n886_), .B(new_n948_), .ZN(new_n6173_));
  AOI21_X1   g5788(.A1(new_n6173_), .A2(new_n953_), .B(new_n958_), .ZN(new_n6174_));
  OAI21_X1   g5789(.A1(new_n6174_), .A2(new_n883_), .B(new_n963_), .ZN(new_n6175_));
  AOI21_X1   g5790(.A1(new_n6175_), .A2(new_n880_), .B(new_n969_), .ZN(new_n6176_));
  OAI21_X1   g5791(.A1(new_n6176_), .A2(new_n973_), .B(new_n977_), .ZN(new_n6177_));
  AOI21_X1   g5792(.A1(new_n6177_), .A2(new_n876_), .B(new_n983_), .ZN(new_n6178_));
  OAI21_X1   g5793(.A1(new_n6178_), .A2(new_n872_), .B(new_n988_), .ZN(new_n6179_));
  AOI21_X1   g5794(.A1(new_n6179_), .A2(new_n993_), .B(new_n998_), .ZN(new_n6180_));
  OAI21_X1   g5795(.A1(new_n6180_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n6181_));
  AOI21_X1   g5796(.A1(new_n6181_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n6182_));
  OAI21_X1   g5797(.A1(new_n6182_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n6183_));
  AOI21_X1   g5798(.A1(new_n6183_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n6184_));
  OAI21_X1   g5799(.A1(new_n6184_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n6185_));
  AOI21_X1   g5800(.A1(new_n6185_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n6186_));
  OAI21_X1   g5801(.A1(new_n6186_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n6187_));
  AOI21_X1   g5802(.A1(new_n6187_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n6188_));
  OAI21_X1   g5803(.A1(new_n6188_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n6189_));
  AOI21_X1   g5804(.A1(new_n6189_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n6190_));
  OAI21_X1   g5805(.A1(new_n6190_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n6191_));
  AOI21_X1   g5806(.A1(new_n6191_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n6192_));
  OAI21_X1   g5807(.A1(new_n6192_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n6193_));
  AOI21_X1   g5808(.A1(new_n6193_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n6194_));
  OAI21_X1   g5809(.A1(new_n6194_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n6195_));
  AOI21_X1   g5810(.A1(new_n6195_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n6196_));
  OAI21_X1   g5811(.A1(new_n6196_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n6197_));
  AOI21_X1   g5812(.A1(new_n6197_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n6198_));
  OAI21_X1   g5813(.A1(new_n6198_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n6199_));
  OAI21_X1   g5814(.A1(new_n1125_), .A2(\priority[105] ), .B(\req[105] ), .ZN(new_n6200_));
  AOI21_X1   g5815(.A1(new_n6199_), .A2(new_n824_), .B(new_n6200_), .ZN(\grant[105] ));
  NOR2_X1    g5816(.A1(new_n1479_), .A2(new_n1136_), .ZN(new_n6202_));
  OAI21_X1   g5817(.A1(new_n819_), .A2(new_n6202_), .B(new_n1142_), .ZN(new_n6203_));
  AOI21_X1   g5818(.A1(new_n6203_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n6204_));
  OAI21_X1   g5819(.A1(new_n6204_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n6205_));
  AOI21_X1   g5820(.A1(new_n6205_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n6206_));
  OAI21_X1   g5821(.A1(new_n6206_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n6207_));
  AOI21_X1   g5822(.A1(new_n6207_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n6208_));
  OAI21_X1   g5823(.A1(new_n6208_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n6209_));
  AOI21_X1   g5824(.A1(new_n6209_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n6210_));
  OAI21_X1   g5825(.A1(new_n6210_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n6211_));
  AOI21_X1   g5826(.A1(new_n6211_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n6212_));
  OAI21_X1   g5827(.A1(new_n6212_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n6213_));
  AOI21_X1   g5828(.A1(new_n6213_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n6214_));
  OAI21_X1   g5829(.A1(new_n6214_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n6215_));
  AOI21_X1   g5830(.A1(new_n6215_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n6216_));
  OAI21_X1   g5831(.A1(new_n6216_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n6217_));
  AOI21_X1   g5832(.A1(new_n6217_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n6218_));
  OAI21_X1   g5833(.A1(new_n6218_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n6219_));
  AOI21_X1   g5834(.A1(new_n6219_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n6220_));
  OAI21_X1   g5835(.A1(new_n6220_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n6221_));
  AOI21_X1   g5836(.A1(new_n6221_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n6222_));
  OAI21_X1   g5837(.A1(new_n6222_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n6223_));
  AOI21_X1   g5838(.A1(new_n6223_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n6224_));
  OAI21_X1   g5839(.A1(new_n6224_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n6225_));
  AOI21_X1   g5840(.A1(new_n6225_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n6226_));
  OAI21_X1   g5841(.A1(new_n6226_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n6227_));
  AOI21_X1   g5842(.A1(new_n6227_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n6228_));
  OAI21_X1   g5843(.A1(new_n6228_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n6229_));
  AOI21_X1   g5844(.A1(new_n6229_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n6230_));
  OAI21_X1   g5845(.A1(new_n6230_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n6231_));
  AOI21_X1   g5846(.A1(new_n6231_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n6232_));
  OAI21_X1   g5847(.A1(new_n6232_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n6233_));
  AOI21_X1   g5848(.A1(new_n6233_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n6234_));
  OAI21_X1   g5849(.A1(new_n6234_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n6235_));
  AOI21_X1   g5850(.A1(new_n6235_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n6236_));
  OAI21_X1   g5851(.A1(new_n6236_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n6237_));
  AOI21_X1   g5852(.A1(new_n6237_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n6238_));
  OAI21_X1   g5853(.A1(new_n6238_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n6239_));
  AOI21_X1   g5854(.A1(new_n6239_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n6240_));
  OAI21_X1   g5855(.A1(new_n6240_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n6241_));
  AOI21_X1   g5856(.A1(new_n6241_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n6242_));
  OAI21_X1   g5857(.A1(new_n6242_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n6243_));
  OAI21_X1   g5858(.A1(new_n749_), .A2(\priority[106] ), .B(\req[106] ), .ZN(new_n6244_));
  AOI21_X1   g5859(.A1(new_n6243_), .A2(new_n1207_), .B(new_n6244_), .ZN(\grant[106] ));
  NOR2_X1    g5860(.A1(new_n401_), .A2(new_n1482_), .ZN(new_n6246_));
  OAI21_X1   g5861(.A1(new_n1202_), .A2(new_n6246_), .B(new_n1487_), .ZN(new_n6247_));
  AOI21_X1   g5862(.A1(new_n6247_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n6248_));
  OAI21_X1   g5863(.A1(new_n6248_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n6249_));
  AOI21_X1   g5864(.A1(new_n6249_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n6250_));
  OAI21_X1   g5865(.A1(new_n6250_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n6251_));
  AOI21_X1   g5866(.A1(new_n6251_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n6252_));
  OAI21_X1   g5867(.A1(new_n6252_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n6253_));
  AOI21_X1   g5868(.A1(new_n6253_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n6254_));
  OAI21_X1   g5869(.A1(new_n6254_), .A2(new_n519_), .B(new_n524_), .ZN(new_n6255_));
  AOI21_X1   g5870(.A1(new_n6255_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n6256_));
  OAI21_X1   g5871(.A1(new_n6256_), .A2(new_n497_), .B(new_n535_), .ZN(new_n6257_));
  AOI21_X1   g5872(.A1(new_n6257_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n6258_));
  OAI21_X1   g5873(.A1(new_n6258_), .A2(new_n492_), .B(new_n550_), .ZN(new_n6259_));
  AOI21_X1   g5874(.A1(new_n6259_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n6260_));
  OAI21_X1   g5875(.A1(new_n6260_), .A2(new_n561_), .B(new_n566_), .ZN(new_n6261_));
  AOI21_X1   g5876(.A1(new_n6261_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n6262_));
  OAI21_X1   g5877(.A1(new_n6262_), .A2(new_n479_), .B(new_n577_), .ZN(new_n6263_));
  AOI21_X1   g5878(.A1(new_n6263_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n6264_));
  OAI21_X1   g5879(.A1(new_n6264_), .A2(new_n474_), .B(new_n592_), .ZN(new_n6265_));
  AOI21_X1   g5880(.A1(new_n6265_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n6266_));
  OAI21_X1   g5881(.A1(new_n6266_), .A2(new_n603_), .B(new_n608_), .ZN(new_n6267_));
  AOI21_X1   g5882(.A1(new_n6267_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n6268_));
  OAI21_X1   g5883(.A1(new_n6268_), .A2(new_n461_), .B(new_n619_), .ZN(new_n6269_));
  AOI21_X1   g5884(.A1(new_n6269_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n6270_));
  OAI21_X1   g5885(.A1(new_n6270_), .A2(new_n456_), .B(new_n634_), .ZN(new_n6271_));
  AOI21_X1   g5886(.A1(new_n6271_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n6272_));
  OAI21_X1   g5887(.A1(new_n6272_), .A2(new_n645_), .B(new_n650_), .ZN(new_n6273_));
  AOI21_X1   g5888(.A1(new_n6273_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n6274_));
  OAI21_X1   g5889(.A1(new_n6274_), .A2(new_n443_), .B(new_n661_), .ZN(new_n6275_));
  AOI21_X1   g5890(.A1(new_n6275_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n6276_));
  OAI21_X1   g5891(.A1(new_n6276_), .A2(new_n438_), .B(new_n676_), .ZN(new_n6277_));
  AOI21_X1   g5892(.A1(new_n6277_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n6278_));
  OAI21_X1   g5893(.A1(new_n6278_), .A2(new_n687_), .B(new_n692_), .ZN(new_n6279_));
  AOI21_X1   g5894(.A1(new_n6279_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n6280_));
  OAI21_X1   g5895(.A1(new_n6280_), .A2(new_n425_), .B(new_n703_), .ZN(new_n6281_));
  AOI21_X1   g5896(.A1(new_n6281_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n6282_));
  OAI21_X1   g5897(.A1(new_n6282_), .A2(new_n420_), .B(new_n718_), .ZN(new_n6283_));
  AOI21_X1   g5898(.A1(new_n6283_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n6284_));
  OAI21_X1   g5899(.A1(new_n6284_), .A2(new_n729_), .B(new_n734_), .ZN(new_n6285_));
  AOI21_X1   g5900(.A1(new_n6285_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n6286_));
  OAI21_X1   g5901(.A1(new_n6286_), .A2(new_n407_), .B(new_n745_), .ZN(new_n6287_));
  OAI21_X1   g5902(.A1(new_n752_), .A2(\priority[107] ), .B(\req[107] ), .ZN(new_n6288_));
  AOI21_X1   g5903(.A1(new_n6287_), .A2(new_n1530_), .B(new_n6288_), .ZN(\grant[107] ));
  NOR2_X1    g5904(.A1(new_n818_), .A2(new_n759_), .ZN(new_n6290_));
  OAI21_X1   g5905(.A1(new_n398_), .A2(new_n6290_), .B(new_n766_), .ZN(new_n6291_));
  AOI21_X1   g5906(.A1(new_n6291_), .A2(new_n772_), .B(new_n777_), .ZN(new_n6292_));
  OAI21_X1   g5907(.A1(new_n6292_), .A2(new_n394_), .B(new_n782_), .ZN(new_n6293_));
  AOI21_X1   g5908(.A1(new_n6293_), .A2(new_n390_), .B(new_n788_), .ZN(new_n6294_));
  OAI21_X1   g5909(.A1(new_n6294_), .A2(new_n793_), .B(new_n797_), .ZN(new_n6295_));
  AOI21_X1   g5910(.A1(new_n6295_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n6296_));
  OAI21_X1   g5911(.A1(new_n6296_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n6297_));
  AOI21_X1   g5912(.A1(new_n6297_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n6298_));
  OAI21_X1   g5913(.A1(new_n6298_), .A2(new_n912_), .B(new_n917_), .ZN(new_n6299_));
  AOI21_X1   g5914(.A1(new_n6299_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n6300_));
  OAI21_X1   g5915(.A1(new_n6300_), .A2(new_n893_), .B(new_n928_), .ZN(new_n6301_));
  AOI21_X1   g5916(.A1(new_n6301_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n6302_));
  OAI21_X1   g5917(.A1(new_n6302_), .A2(new_n889_), .B(new_n942_), .ZN(new_n6303_));
  AOI21_X1   g5918(.A1(new_n6303_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n6304_));
  OAI21_X1   g5919(.A1(new_n6304_), .A2(new_n952_), .B(new_n957_), .ZN(new_n6305_));
  AOI21_X1   g5920(.A1(new_n6305_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n6306_));
  OAI21_X1   g5921(.A1(new_n6306_), .A2(new_n879_), .B(new_n968_), .ZN(new_n6307_));
  AOI21_X1   g5922(.A1(new_n6307_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n6308_));
  OAI21_X1   g5923(.A1(new_n6308_), .A2(new_n875_), .B(new_n982_), .ZN(new_n6309_));
  AOI21_X1   g5924(.A1(new_n6309_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n6310_));
  OAI21_X1   g5925(.A1(new_n6310_), .A2(new_n992_), .B(new_n997_), .ZN(new_n6311_));
  AOI21_X1   g5926(.A1(new_n6311_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n6312_));
  OAI21_X1   g5927(.A1(new_n6312_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n6313_));
  AOI21_X1   g5928(.A1(new_n6313_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n6314_));
  OAI21_X1   g5929(.A1(new_n6314_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n6315_));
  AOI21_X1   g5930(.A1(new_n6315_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n6316_));
  OAI21_X1   g5931(.A1(new_n6316_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n6317_));
  AOI21_X1   g5932(.A1(new_n6317_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n6318_));
  OAI21_X1   g5933(.A1(new_n6318_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n6319_));
  AOI21_X1   g5934(.A1(new_n6319_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n6320_));
  OAI21_X1   g5935(.A1(new_n6320_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n6321_));
  AOI21_X1   g5936(.A1(new_n6321_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n6322_));
  OAI21_X1   g5937(.A1(new_n6322_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n6323_));
  AOI21_X1   g5938(.A1(new_n6323_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n6324_));
  OAI21_X1   g5939(.A1(new_n6324_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n6325_));
  AOI21_X1   g5940(.A1(new_n6325_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n6326_));
  OAI21_X1   g5941(.A1(new_n6326_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n6327_));
  AOI21_X1   g5942(.A1(new_n6327_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n6328_));
  OAI21_X1   g5943(.A1(new_n6328_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n6329_));
  AOI21_X1   g5944(.A1(new_n6329_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n6330_));
  OAI21_X1   g5945(.A1(new_n6330_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n6331_));
  OAI21_X1   g5946(.A1(new_n1134_), .A2(\priority[108] ), .B(\req[108] ), .ZN(new_n6332_));
  AOI21_X1   g5947(.A1(new_n6331_), .A2(new_n1620_), .B(new_n6332_), .ZN(\grant[108] ));
  NOR2_X1    g5948(.A1(new_n1201_), .A2(new_n1141_), .ZN(new_n6334_));
  OAI21_X1   g5949(.A1(new_n816_), .A2(new_n6334_), .B(new_n1148_), .ZN(new_n6335_));
  AOI21_X1   g5950(.A1(new_n6335_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n6336_));
  OAI21_X1   g5951(.A1(new_n6336_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n6337_));
  AOI21_X1   g5952(.A1(new_n6337_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n6338_));
  OAI21_X1   g5953(.A1(new_n6338_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n6339_));
  AOI21_X1   g5954(.A1(new_n6339_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n6340_));
  OAI21_X1   g5955(.A1(new_n6340_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n6341_));
  AOI21_X1   g5956(.A1(new_n6341_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n6342_));
  OAI21_X1   g5957(.A1(new_n6342_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n6343_));
  AOI21_X1   g5958(.A1(new_n6343_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n6344_));
  OAI21_X1   g5959(.A1(new_n6344_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n6345_));
  AOI21_X1   g5960(.A1(new_n6345_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n6346_));
  OAI21_X1   g5961(.A1(new_n6346_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n6347_));
  AOI21_X1   g5962(.A1(new_n6347_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n6348_));
  OAI21_X1   g5963(.A1(new_n6348_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n6349_));
  AOI21_X1   g5964(.A1(new_n6349_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n6350_));
  OAI21_X1   g5965(.A1(new_n6350_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n6351_));
  AOI21_X1   g5966(.A1(new_n6351_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n6352_));
  OAI21_X1   g5967(.A1(new_n6352_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n6353_));
  AOI21_X1   g5968(.A1(new_n6353_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n6354_));
  OAI21_X1   g5969(.A1(new_n6354_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n6355_));
  AOI21_X1   g5970(.A1(new_n6355_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n6356_));
  OAI21_X1   g5971(.A1(new_n6356_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n6357_));
  AOI21_X1   g5972(.A1(new_n6357_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n6358_));
  OAI21_X1   g5973(.A1(new_n6358_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n6359_));
  AOI21_X1   g5974(.A1(new_n6359_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n6360_));
  OAI21_X1   g5975(.A1(new_n6360_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n6361_));
  AOI21_X1   g5976(.A1(new_n6361_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n6362_));
  OAI21_X1   g5977(.A1(new_n6362_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n6363_));
  AOI21_X1   g5978(.A1(new_n6363_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n6364_));
  OAI21_X1   g5979(.A1(new_n6364_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n6365_));
  AOI21_X1   g5980(.A1(new_n6365_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n6366_));
  OAI21_X1   g5981(.A1(new_n6366_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n6367_));
  AOI21_X1   g5982(.A1(new_n6367_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n6368_));
  OAI21_X1   g5983(.A1(new_n6368_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n6369_));
  AOI21_X1   g5984(.A1(new_n6369_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n6370_));
  OAI21_X1   g5985(.A1(new_n6370_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n6371_));
  AOI21_X1   g5986(.A1(new_n6371_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n6372_));
  OAI21_X1   g5987(.A1(new_n6372_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n6373_));
  AOI21_X1   g5988(.A1(new_n6373_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n6374_));
  OAI21_X1   g5989(.A1(new_n6374_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n6375_));
  OAI21_X1   g5990(.A1(new_n400_), .A2(\priority[109] ), .B(\req[109] ), .ZN(new_n6376_));
  AOI21_X1   g5991(.A1(new_n6375_), .A2(new_n1708_), .B(new_n6376_), .ZN(\grant[109] ));
  NOR2_X1    g5992(.A1(new_n397_), .A2(new_n1486_), .ZN(new_n6378_));
  OAI21_X1   g5993(.A1(new_n1199_), .A2(new_n6378_), .B(new_n1492_), .ZN(new_n6379_));
  AOI21_X1   g5994(.A1(new_n6379_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n6380_));
  OAI21_X1   g5995(.A1(new_n6380_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n6381_));
  AOI21_X1   g5996(.A1(new_n6381_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n6382_));
  OAI21_X1   g5997(.A1(new_n6382_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n6383_));
  AOI21_X1   g5998(.A1(new_n6383_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n6384_));
  OAI21_X1   g5999(.A1(new_n6384_), .A2(new_n506_), .B(new_n514_), .ZN(new_n6385_));
  AOI21_X1   g6000(.A1(new_n6385_), .A2(new_n520_), .B(new_n525_), .ZN(new_n6386_));
  OAI21_X1   g6001(.A1(new_n6386_), .A2(new_n502_), .B(new_n530_), .ZN(new_n6387_));
  AOI21_X1   g6002(.A1(new_n6387_), .A2(new_n498_), .B(new_n536_), .ZN(new_n6388_));
  OAI21_X1   g6003(.A1(new_n6388_), .A2(new_n541_), .B(new_n545_), .ZN(new_n6389_));
  AOI21_X1   g6004(.A1(new_n6389_), .A2(new_n493_), .B(new_n551_), .ZN(new_n6390_));
  OAI21_X1   g6005(.A1(new_n6390_), .A2(new_n488_), .B(new_n556_), .ZN(new_n6391_));
  AOI21_X1   g6006(.A1(new_n6391_), .A2(new_n562_), .B(new_n567_), .ZN(new_n6392_));
  OAI21_X1   g6007(.A1(new_n6392_), .A2(new_n484_), .B(new_n572_), .ZN(new_n6393_));
  AOI21_X1   g6008(.A1(new_n6393_), .A2(new_n480_), .B(new_n578_), .ZN(new_n6394_));
  OAI21_X1   g6009(.A1(new_n6394_), .A2(new_n583_), .B(new_n587_), .ZN(new_n6395_));
  AOI21_X1   g6010(.A1(new_n6395_), .A2(new_n475_), .B(new_n593_), .ZN(new_n6396_));
  OAI21_X1   g6011(.A1(new_n6396_), .A2(new_n470_), .B(new_n598_), .ZN(new_n6397_));
  AOI21_X1   g6012(.A1(new_n6397_), .A2(new_n604_), .B(new_n609_), .ZN(new_n6398_));
  OAI21_X1   g6013(.A1(new_n6398_), .A2(new_n466_), .B(new_n614_), .ZN(new_n6399_));
  AOI21_X1   g6014(.A1(new_n6399_), .A2(new_n462_), .B(new_n620_), .ZN(new_n6400_));
  OAI21_X1   g6015(.A1(new_n6400_), .A2(new_n625_), .B(new_n629_), .ZN(new_n6401_));
  AOI21_X1   g6016(.A1(new_n6401_), .A2(new_n457_), .B(new_n635_), .ZN(new_n6402_));
  OAI21_X1   g6017(.A1(new_n6402_), .A2(new_n452_), .B(new_n640_), .ZN(new_n6403_));
  AOI21_X1   g6018(.A1(new_n6403_), .A2(new_n646_), .B(new_n651_), .ZN(new_n6404_));
  OAI21_X1   g6019(.A1(new_n6404_), .A2(new_n448_), .B(new_n656_), .ZN(new_n6405_));
  AOI21_X1   g6020(.A1(new_n6405_), .A2(new_n444_), .B(new_n662_), .ZN(new_n6406_));
  OAI21_X1   g6021(.A1(new_n6406_), .A2(new_n667_), .B(new_n671_), .ZN(new_n6407_));
  AOI21_X1   g6022(.A1(new_n6407_), .A2(new_n439_), .B(new_n677_), .ZN(new_n6408_));
  OAI21_X1   g6023(.A1(new_n6408_), .A2(new_n434_), .B(new_n682_), .ZN(new_n6409_));
  AOI21_X1   g6024(.A1(new_n6409_), .A2(new_n688_), .B(new_n693_), .ZN(new_n6410_));
  OAI21_X1   g6025(.A1(new_n6410_), .A2(new_n430_), .B(new_n698_), .ZN(new_n6411_));
  AOI21_X1   g6026(.A1(new_n6411_), .A2(new_n426_), .B(new_n704_), .ZN(new_n6412_));
  OAI21_X1   g6027(.A1(new_n6412_), .A2(new_n709_), .B(new_n713_), .ZN(new_n6413_));
  AOI21_X1   g6028(.A1(new_n6413_), .A2(new_n421_), .B(new_n719_), .ZN(new_n6414_));
  OAI21_X1   g6029(.A1(new_n6414_), .A2(new_n416_), .B(new_n724_), .ZN(new_n6415_));
  AOI21_X1   g6030(.A1(new_n6415_), .A2(new_n730_), .B(new_n735_), .ZN(new_n6416_));
  OAI21_X1   g6031(.A1(new_n6416_), .A2(new_n412_), .B(new_n740_), .ZN(new_n6417_));
  AOI21_X1   g6032(.A1(new_n6417_), .A2(new_n408_), .B(new_n746_), .ZN(new_n6418_));
  OAI21_X1   g6033(.A1(new_n6418_), .A2(new_n751_), .B(new_n755_), .ZN(new_n6419_));
  OAI21_X1   g6034(.A1(new_n757_), .A2(\priority[110] ), .B(\req[110] ), .ZN(new_n6420_));
  AOI21_X1   g6035(.A1(new_n6419_), .A2(new_n403_), .B(new_n6420_), .ZN(\grant[110] ));
  NOR2_X1    g6036(.A1(new_n815_), .A2(new_n765_), .ZN(new_n6422_));
  OAI21_X1   g6037(.A1(new_n771_), .A2(new_n6422_), .B(new_n776_), .ZN(new_n6423_));
  AOI21_X1   g6038(.A1(new_n6423_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n6424_));
  OAI21_X1   g6039(.A1(new_n6424_), .A2(new_n389_), .B(new_n787_), .ZN(new_n6425_));
  AOI21_X1   g6040(.A1(new_n6425_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n6426_));
  OAI21_X1   g6041(.A1(new_n6426_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n6427_));
  AOI21_X1   g6042(.A1(new_n6427_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n6428_));
  OAI21_X1   g6043(.A1(new_n6428_), .A2(new_n900_), .B(new_n908_), .ZN(new_n6429_));
  AOI21_X1   g6044(.A1(new_n6429_), .A2(new_n913_), .B(new_n918_), .ZN(new_n6430_));
  OAI21_X1   g6045(.A1(new_n6430_), .A2(new_n897_), .B(new_n923_), .ZN(new_n6431_));
  AOI21_X1   g6046(.A1(new_n6431_), .A2(new_n894_), .B(new_n929_), .ZN(new_n6432_));
  OAI21_X1   g6047(.A1(new_n6432_), .A2(new_n933_), .B(new_n937_), .ZN(new_n6433_));
  AOI21_X1   g6048(.A1(new_n6433_), .A2(new_n890_), .B(new_n943_), .ZN(new_n6434_));
  OAI21_X1   g6049(.A1(new_n6434_), .A2(new_n886_), .B(new_n948_), .ZN(new_n6435_));
  AOI21_X1   g6050(.A1(new_n6435_), .A2(new_n953_), .B(new_n958_), .ZN(new_n6436_));
  OAI21_X1   g6051(.A1(new_n6436_), .A2(new_n883_), .B(new_n963_), .ZN(new_n6437_));
  AOI21_X1   g6052(.A1(new_n6437_), .A2(new_n880_), .B(new_n969_), .ZN(new_n6438_));
  OAI21_X1   g6053(.A1(new_n6438_), .A2(new_n973_), .B(new_n977_), .ZN(new_n6439_));
  AOI21_X1   g6054(.A1(new_n6439_), .A2(new_n876_), .B(new_n983_), .ZN(new_n6440_));
  OAI21_X1   g6055(.A1(new_n6440_), .A2(new_n872_), .B(new_n988_), .ZN(new_n6441_));
  AOI21_X1   g6056(.A1(new_n6441_), .A2(new_n993_), .B(new_n998_), .ZN(new_n6442_));
  OAI21_X1   g6057(.A1(new_n6442_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n6443_));
  AOI21_X1   g6058(.A1(new_n6443_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n6444_));
  OAI21_X1   g6059(.A1(new_n6444_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n6445_));
  AOI21_X1   g6060(.A1(new_n6445_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n6446_));
  OAI21_X1   g6061(.A1(new_n6446_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n6447_));
  AOI21_X1   g6062(.A1(new_n6447_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n6448_));
  OAI21_X1   g6063(.A1(new_n6448_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n6449_));
  AOI21_X1   g6064(.A1(new_n6449_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n6450_));
  OAI21_X1   g6065(.A1(new_n6450_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n6451_));
  AOI21_X1   g6066(.A1(new_n6451_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n6452_));
  OAI21_X1   g6067(.A1(new_n6452_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n6453_));
  AOI21_X1   g6068(.A1(new_n6453_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n6454_));
  OAI21_X1   g6069(.A1(new_n6454_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n6455_));
  AOI21_X1   g6070(.A1(new_n6455_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n6456_));
  OAI21_X1   g6071(.A1(new_n6456_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n6457_));
  AOI21_X1   g6072(.A1(new_n6457_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n6458_));
  OAI21_X1   g6073(.A1(new_n6458_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n6459_));
  AOI21_X1   g6074(.A1(new_n6459_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n6460_));
  OAI21_X1   g6075(.A1(new_n6460_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n6461_));
  AOI21_X1   g6076(.A1(new_n6461_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n6462_));
  OAI21_X1   g6077(.A1(new_n6462_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n6463_));
  OAI21_X1   g6078(.A1(new_n1139_), .A2(\priority[111] ), .B(\req[111] ), .ZN(new_n6464_));
  AOI21_X1   g6079(.A1(new_n6463_), .A2(new_n820_), .B(new_n6464_), .ZN(\grant[111] ));
  NOR2_X1    g6080(.A1(new_n1198_), .A2(new_n1147_), .ZN(new_n6466_));
  OAI21_X1   g6081(.A1(new_n1152_), .A2(new_n6466_), .B(new_n1157_), .ZN(new_n6467_));
  AOI21_X1   g6082(.A1(new_n6467_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n6468_));
  OAI21_X1   g6083(.A1(new_n6468_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n6469_));
  AOI21_X1   g6084(.A1(new_n6469_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n6470_));
  OAI21_X1   g6085(.A1(new_n6470_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n6471_));
  AOI21_X1   g6086(.A1(new_n6471_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n6472_));
  OAI21_X1   g6087(.A1(new_n6472_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n6473_));
  AOI21_X1   g6088(.A1(new_n6473_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n6474_));
  OAI21_X1   g6089(.A1(new_n6474_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n6475_));
  AOI21_X1   g6090(.A1(new_n6475_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n6476_));
  OAI21_X1   g6091(.A1(new_n6476_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n6477_));
  AOI21_X1   g6092(.A1(new_n6477_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n6478_));
  OAI21_X1   g6093(.A1(new_n6478_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n6479_));
  AOI21_X1   g6094(.A1(new_n6479_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n6480_));
  OAI21_X1   g6095(.A1(new_n6480_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n6481_));
  AOI21_X1   g6096(.A1(new_n6481_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n6482_));
  OAI21_X1   g6097(.A1(new_n6482_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n6483_));
  AOI21_X1   g6098(.A1(new_n6483_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n6484_));
  OAI21_X1   g6099(.A1(new_n6484_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n6485_));
  AOI21_X1   g6100(.A1(new_n6485_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n6486_));
  OAI21_X1   g6101(.A1(new_n6486_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n6487_));
  AOI21_X1   g6102(.A1(new_n6487_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n6488_));
  OAI21_X1   g6103(.A1(new_n6488_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n6489_));
  AOI21_X1   g6104(.A1(new_n6489_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n6490_));
  OAI21_X1   g6105(.A1(new_n6490_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n6491_));
  AOI21_X1   g6106(.A1(new_n6491_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n6492_));
  OAI21_X1   g6107(.A1(new_n6492_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n6493_));
  AOI21_X1   g6108(.A1(new_n6493_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n6494_));
  OAI21_X1   g6109(.A1(new_n6494_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n6495_));
  AOI21_X1   g6110(.A1(new_n6495_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n6496_));
  OAI21_X1   g6111(.A1(new_n6496_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n6497_));
  AOI21_X1   g6112(.A1(new_n6497_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n6498_));
  OAI21_X1   g6113(.A1(new_n6498_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n6499_));
  AOI21_X1   g6114(.A1(new_n6499_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n6500_));
  OAI21_X1   g6115(.A1(new_n6500_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n6501_));
  AOI21_X1   g6116(.A1(new_n6501_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n6502_));
  OAI21_X1   g6117(.A1(new_n6502_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n6503_));
  AOI21_X1   g6118(.A1(new_n6503_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n6504_));
  OAI21_X1   g6119(.A1(new_n6504_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n6505_));
  AOI21_X1   g6120(.A1(new_n6505_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n6506_));
  OAI21_X1   g6121(.A1(new_n6506_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n6507_));
  OAI21_X1   g6122(.A1(new_n396_), .A2(\priority[112] ), .B(\req[112] ), .ZN(new_n6508_));
  AOI21_X1   g6123(.A1(new_n6507_), .A2(new_n1203_), .B(new_n6508_), .ZN(\grant[112] ));
  NOR2_X1    g6124(.A1(new_n770_), .A2(new_n1491_), .ZN(new_n6510_));
  OAI21_X1   g6125(.A1(new_n1496_), .A2(new_n6510_), .B(new_n1500_), .ZN(new_n6511_));
  AOI21_X1   g6126(.A1(new_n6511_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n6512_));
  OAI21_X1   g6127(.A1(new_n6512_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n6513_));
  AOI21_X1   g6128(.A1(new_n6513_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n6514_));
  OAI21_X1   g6129(.A1(new_n6514_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n6515_));
  AOI21_X1   g6130(.A1(new_n6515_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n6516_));
  OAI21_X1   g6131(.A1(new_n6516_), .A2(new_n519_), .B(new_n524_), .ZN(new_n6517_));
  AOI21_X1   g6132(.A1(new_n6517_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n6518_));
  OAI21_X1   g6133(.A1(new_n6518_), .A2(new_n497_), .B(new_n535_), .ZN(new_n6519_));
  AOI21_X1   g6134(.A1(new_n6519_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n6520_));
  OAI21_X1   g6135(.A1(new_n6520_), .A2(new_n492_), .B(new_n550_), .ZN(new_n6521_));
  AOI21_X1   g6136(.A1(new_n6521_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n6522_));
  OAI21_X1   g6137(.A1(new_n6522_), .A2(new_n561_), .B(new_n566_), .ZN(new_n6523_));
  AOI21_X1   g6138(.A1(new_n6523_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n6524_));
  OAI21_X1   g6139(.A1(new_n6524_), .A2(new_n479_), .B(new_n577_), .ZN(new_n6525_));
  AOI21_X1   g6140(.A1(new_n6525_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n6526_));
  OAI21_X1   g6141(.A1(new_n6526_), .A2(new_n474_), .B(new_n592_), .ZN(new_n6527_));
  AOI21_X1   g6142(.A1(new_n6527_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n6528_));
  OAI21_X1   g6143(.A1(new_n6528_), .A2(new_n603_), .B(new_n608_), .ZN(new_n6529_));
  AOI21_X1   g6144(.A1(new_n6529_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n6530_));
  OAI21_X1   g6145(.A1(new_n6530_), .A2(new_n461_), .B(new_n619_), .ZN(new_n6531_));
  AOI21_X1   g6146(.A1(new_n6531_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n6532_));
  OAI21_X1   g6147(.A1(new_n6532_), .A2(new_n456_), .B(new_n634_), .ZN(new_n6533_));
  AOI21_X1   g6148(.A1(new_n6533_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n6534_));
  OAI21_X1   g6149(.A1(new_n6534_), .A2(new_n645_), .B(new_n650_), .ZN(new_n6535_));
  AOI21_X1   g6150(.A1(new_n6535_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n6536_));
  OAI21_X1   g6151(.A1(new_n6536_), .A2(new_n443_), .B(new_n661_), .ZN(new_n6537_));
  AOI21_X1   g6152(.A1(new_n6537_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n6538_));
  OAI21_X1   g6153(.A1(new_n6538_), .A2(new_n438_), .B(new_n676_), .ZN(new_n6539_));
  AOI21_X1   g6154(.A1(new_n6539_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n6540_));
  OAI21_X1   g6155(.A1(new_n6540_), .A2(new_n687_), .B(new_n692_), .ZN(new_n6541_));
  AOI21_X1   g6156(.A1(new_n6541_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n6542_));
  OAI21_X1   g6157(.A1(new_n6542_), .A2(new_n425_), .B(new_n703_), .ZN(new_n6543_));
  AOI21_X1   g6158(.A1(new_n6543_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n6544_));
  OAI21_X1   g6159(.A1(new_n6544_), .A2(new_n420_), .B(new_n718_), .ZN(new_n6545_));
  AOI21_X1   g6160(.A1(new_n6545_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n6546_));
  OAI21_X1   g6161(.A1(new_n6546_), .A2(new_n729_), .B(new_n734_), .ZN(new_n6547_));
  AOI21_X1   g6162(.A1(new_n6547_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n6548_));
  OAI21_X1   g6163(.A1(new_n6548_), .A2(new_n407_), .B(new_n745_), .ZN(new_n6549_));
  AOI21_X1   g6164(.A1(new_n6549_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n6550_));
  OAI21_X1   g6165(.A1(new_n6550_), .A2(new_n402_), .B(new_n760_), .ZN(new_n6551_));
  OAI21_X1   g6166(.A1(new_n763_), .A2(\priority[113] ), .B(\req[113] ), .ZN(new_n6552_));
  AOI21_X1   g6167(.A1(new_n6551_), .A2(new_n1528_), .B(new_n6552_), .ZN(\grant[113] ));
  NOR2_X1    g6168(.A1(new_n1151_), .A2(new_n775_), .ZN(new_n6554_));
  OAI21_X1   g6169(.A1(new_n394_), .A2(new_n6554_), .B(new_n782_), .ZN(new_n6555_));
  AOI21_X1   g6170(.A1(new_n6555_), .A2(new_n390_), .B(new_n788_), .ZN(new_n6556_));
  OAI21_X1   g6171(.A1(new_n6556_), .A2(new_n793_), .B(new_n797_), .ZN(new_n6557_));
  AOI21_X1   g6172(.A1(new_n6557_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n6558_));
  OAI21_X1   g6173(.A1(new_n6558_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n6559_));
  AOI21_X1   g6174(.A1(new_n6559_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n6560_));
  OAI21_X1   g6175(.A1(new_n6560_), .A2(new_n912_), .B(new_n917_), .ZN(new_n6561_));
  AOI21_X1   g6176(.A1(new_n6561_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n6562_));
  OAI21_X1   g6177(.A1(new_n6562_), .A2(new_n893_), .B(new_n928_), .ZN(new_n6563_));
  AOI21_X1   g6178(.A1(new_n6563_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n6564_));
  OAI21_X1   g6179(.A1(new_n6564_), .A2(new_n889_), .B(new_n942_), .ZN(new_n6565_));
  AOI21_X1   g6180(.A1(new_n6565_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n6566_));
  OAI21_X1   g6181(.A1(new_n6566_), .A2(new_n952_), .B(new_n957_), .ZN(new_n6567_));
  AOI21_X1   g6182(.A1(new_n6567_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n6568_));
  OAI21_X1   g6183(.A1(new_n6568_), .A2(new_n879_), .B(new_n968_), .ZN(new_n6569_));
  AOI21_X1   g6184(.A1(new_n6569_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n6570_));
  OAI21_X1   g6185(.A1(new_n6570_), .A2(new_n875_), .B(new_n982_), .ZN(new_n6571_));
  AOI21_X1   g6186(.A1(new_n6571_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n6572_));
  OAI21_X1   g6187(.A1(new_n6572_), .A2(new_n992_), .B(new_n997_), .ZN(new_n6573_));
  AOI21_X1   g6188(.A1(new_n6573_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n6574_));
  OAI21_X1   g6189(.A1(new_n6574_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n6575_));
  AOI21_X1   g6190(.A1(new_n6575_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n6576_));
  OAI21_X1   g6191(.A1(new_n6576_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n6577_));
  AOI21_X1   g6192(.A1(new_n6577_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n6578_));
  OAI21_X1   g6193(.A1(new_n6578_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n6579_));
  AOI21_X1   g6194(.A1(new_n6579_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n6580_));
  OAI21_X1   g6195(.A1(new_n6580_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n6581_));
  AOI21_X1   g6196(.A1(new_n6581_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n6582_));
  OAI21_X1   g6197(.A1(new_n6582_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n6583_));
  AOI21_X1   g6198(.A1(new_n6583_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n6584_));
  OAI21_X1   g6199(.A1(new_n6584_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n6585_));
  AOI21_X1   g6200(.A1(new_n6585_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n6586_));
  OAI21_X1   g6201(.A1(new_n6586_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n6587_));
  AOI21_X1   g6202(.A1(new_n6587_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n6588_));
  OAI21_X1   g6203(.A1(new_n6588_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n6589_));
  AOI21_X1   g6204(.A1(new_n6589_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n6590_));
  OAI21_X1   g6205(.A1(new_n6590_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n6591_));
  AOI21_X1   g6206(.A1(new_n6591_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n6592_));
  OAI21_X1   g6207(.A1(new_n6592_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n6593_));
  AOI21_X1   g6208(.A1(new_n6593_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n6594_));
  OAI21_X1   g6209(.A1(new_n6594_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n6595_));
  OAI21_X1   g6210(.A1(new_n1145_), .A2(\priority[114] ), .B(\req[114] ), .ZN(new_n6596_));
  AOI21_X1   g6211(.A1(new_n6595_), .A2(new_n1618_), .B(new_n6596_), .ZN(\grant[114] ));
  NOR2_X1    g6212(.A1(new_n1495_), .A2(new_n1156_), .ZN(new_n6598_));
  OAI21_X1   g6213(.A1(new_n813_), .A2(new_n6598_), .B(new_n1163_), .ZN(new_n6599_));
  AOI21_X1   g6214(.A1(new_n6599_), .A2(new_n810_), .B(new_n1169_), .ZN(new_n6600_));
  OAI21_X1   g6215(.A1(new_n6600_), .A2(new_n1173_), .B(new_n1177_), .ZN(new_n6601_));
  AOI21_X1   g6216(.A1(new_n6601_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n6602_));
  OAI21_X1   g6217(.A1(new_n6602_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n6603_));
  AOI21_X1   g6218(.A1(new_n6603_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n6604_));
  OAI21_X1   g6219(.A1(new_n6604_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n6605_));
  AOI21_X1   g6220(.A1(new_n6605_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n6606_));
  OAI21_X1   g6221(.A1(new_n6606_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n6607_));
  AOI21_X1   g6222(.A1(new_n6607_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n6608_));
  OAI21_X1   g6223(.A1(new_n6608_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n6609_));
  AOI21_X1   g6224(.A1(new_n6609_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n6610_));
  OAI21_X1   g6225(.A1(new_n6610_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n6611_));
  AOI21_X1   g6226(.A1(new_n6611_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n6612_));
  OAI21_X1   g6227(.A1(new_n6612_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n6613_));
  AOI21_X1   g6228(.A1(new_n6613_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n6614_));
  OAI21_X1   g6229(.A1(new_n6614_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n6615_));
  AOI21_X1   g6230(.A1(new_n6615_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n6616_));
  OAI21_X1   g6231(.A1(new_n6616_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n6617_));
  AOI21_X1   g6232(.A1(new_n6617_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n6618_));
  OAI21_X1   g6233(.A1(new_n6618_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n6619_));
  AOI21_X1   g6234(.A1(new_n6619_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n6620_));
  OAI21_X1   g6235(.A1(new_n6620_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n6621_));
  AOI21_X1   g6236(.A1(new_n6621_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n6622_));
  OAI21_X1   g6237(.A1(new_n6622_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n6623_));
  AOI21_X1   g6238(.A1(new_n6623_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n6624_));
  OAI21_X1   g6239(.A1(new_n6624_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n6625_));
  AOI21_X1   g6240(.A1(new_n6625_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n6626_));
  OAI21_X1   g6241(.A1(new_n6626_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n6627_));
  AOI21_X1   g6242(.A1(new_n6627_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n6628_));
  OAI21_X1   g6243(.A1(new_n6628_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n6629_));
  AOI21_X1   g6244(.A1(new_n6629_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n6630_));
  OAI21_X1   g6245(.A1(new_n6630_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n6631_));
  AOI21_X1   g6246(.A1(new_n6631_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n6632_));
  OAI21_X1   g6247(.A1(new_n6632_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n6633_));
  AOI21_X1   g6248(.A1(new_n6633_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n6634_));
  OAI21_X1   g6249(.A1(new_n6634_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n6635_));
  AOI21_X1   g6250(.A1(new_n6635_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n6636_));
  OAI21_X1   g6251(.A1(new_n6636_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n6637_));
  AOI21_X1   g6252(.A1(new_n6637_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n6638_));
  OAI21_X1   g6253(.A1(new_n6638_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n6639_));
  OAI21_X1   g6254(.A1(new_n769_), .A2(\priority[115] ), .B(\req[115] ), .ZN(new_n6640_));
  AOI21_X1   g6255(.A1(new_n6639_), .A2(new_n1706_), .B(new_n6640_), .ZN(\grant[115] ));
  NOR2_X1    g6256(.A1(new_n393_), .A2(new_n1499_), .ZN(new_n6642_));
  OAI21_X1   g6257(.A1(new_n1196_), .A2(new_n6642_), .B(new_n1505_), .ZN(new_n6643_));
  AOI21_X1   g6258(.A1(new_n6643_), .A2(new_n1193_), .B(new_n1510_), .ZN(new_n6644_));
  OAI21_X1   g6259(.A1(new_n6644_), .A2(new_n1514_), .B(new_n1517_), .ZN(new_n6645_));
  AOI21_X1   g6260(.A1(new_n6645_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n6646_));
  OAI21_X1   g6261(.A1(new_n6646_), .A2(new_n506_), .B(new_n514_), .ZN(new_n6647_));
  AOI21_X1   g6262(.A1(new_n6647_), .A2(new_n520_), .B(new_n525_), .ZN(new_n6648_));
  OAI21_X1   g6263(.A1(new_n6648_), .A2(new_n502_), .B(new_n530_), .ZN(new_n6649_));
  AOI21_X1   g6264(.A1(new_n6649_), .A2(new_n498_), .B(new_n536_), .ZN(new_n6650_));
  OAI21_X1   g6265(.A1(new_n6650_), .A2(new_n541_), .B(new_n545_), .ZN(new_n6651_));
  AOI21_X1   g6266(.A1(new_n6651_), .A2(new_n493_), .B(new_n551_), .ZN(new_n6652_));
  OAI21_X1   g6267(.A1(new_n6652_), .A2(new_n488_), .B(new_n556_), .ZN(new_n6653_));
  AOI21_X1   g6268(.A1(new_n6653_), .A2(new_n562_), .B(new_n567_), .ZN(new_n6654_));
  OAI21_X1   g6269(.A1(new_n6654_), .A2(new_n484_), .B(new_n572_), .ZN(new_n6655_));
  AOI21_X1   g6270(.A1(new_n6655_), .A2(new_n480_), .B(new_n578_), .ZN(new_n6656_));
  OAI21_X1   g6271(.A1(new_n6656_), .A2(new_n583_), .B(new_n587_), .ZN(new_n6657_));
  AOI21_X1   g6272(.A1(new_n6657_), .A2(new_n475_), .B(new_n593_), .ZN(new_n6658_));
  OAI21_X1   g6273(.A1(new_n6658_), .A2(new_n470_), .B(new_n598_), .ZN(new_n6659_));
  AOI21_X1   g6274(.A1(new_n6659_), .A2(new_n604_), .B(new_n609_), .ZN(new_n6660_));
  OAI21_X1   g6275(.A1(new_n6660_), .A2(new_n466_), .B(new_n614_), .ZN(new_n6661_));
  AOI21_X1   g6276(.A1(new_n6661_), .A2(new_n462_), .B(new_n620_), .ZN(new_n6662_));
  OAI21_X1   g6277(.A1(new_n6662_), .A2(new_n625_), .B(new_n629_), .ZN(new_n6663_));
  AOI21_X1   g6278(.A1(new_n6663_), .A2(new_n457_), .B(new_n635_), .ZN(new_n6664_));
  OAI21_X1   g6279(.A1(new_n6664_), .A2(new_n452_), .B(new_n640_), .ZN(new_n6665_));
  AOI21_X1   g6280(.A1(new_n6665_), .A2(new_n646_), .B(new_n651_), .ZN(new_n6666_));
  OAI21_X1   g6281(.A1(new_n6666_), .A2(new_n448_), .B(new_n656_), .ZN(new_n6667_));
  AOI21_X1   g6282(.A1(new_n6667_), .A2(new_n444_), .B(new_n662_), .ZN(new_n6668_));
  OAI21_X1   g6283(.A1(new_n6668_), .A2(new_n667_), .B(new_n671_), .ZN(new_n6669_));
  AOI21_X1   g6284(.A1(new_n6669_), .A2(new_n439_), .B(new_n677_), .ZN(new_n6670_));
  OAI21_X1   g6285(.A1(new_n6670_), .A2(new_n434_), .B(new_n682_), .ZN(new_n6671_));
  AOI21_X1   g6286(.A1(new_n6671_), .A2(new_n688_), .B(new_n693_), .ZN(new_n6672_));
  OAI21_X1   g6287(.A1(new_n6672_), .A2(new_n430_), .B(new_n698_), .ZN(new_n6673_));
  AOI21_X1   g6288(.A1(new_n6673_), .A2(new_n426_), .B(new_n704_), .ZN(new_n6674_));
  OAI21_X1   g6289(.A1(new_n6674_), .A2(new_n709_), .B(new_n713_), .ZN(new_n6675_));
  AOI21_X1   g6290(.A1(new_n6675_), .A2(new_n421_), .B(new_n719_), .ZN(new_n6676_));
  OAI21_X1   g6291(.A1(new_n6676_), .A2(new_n416_), .B(new_n724_), .ZN(new_n6677_));
  AOI21_X1   g6292(.A1(new_n6677_), .A2(new_n730_), .B(new_n735_), .ZN(new_n6678_));
  OAI21_X1   g6293(.A1(new_n6678_), .A2(new_n412_), .B(new_n740_), .ZN(new_n6679_));
  AOI21_X1   g6294(.A1(new_n6679_), .A2(new_n408_), .B(new_n746_), .ZN(new_n6680_));
  OAI21_X1   g6295(.A1(new_n6680_), .A2(new_n751_), .B(new_n755_), .ZN(new_n6681_));
  AOI21_X1   g6296(.A1(new_n6681_), .A2(new_n403_), .B(new_n761_), .ZN(new_n6682_));
  OAI21_X1   g6297(.A1(new_n6682_), .A2(new_n398_), .B(new_n766_), .ZN(new_n6683_));
  OAI21_X1   g6298(.A1(new_n773_), .A2(\priority[116] ), .B(\req[116] ), .ZN(new_n6684_));
  AOI21_X1   g6299(.A1(new_n6683_), .A2(new_n772_), .B(new_n6684_), .ZN(\grant[116] ));
  NOR2_X1    g6300(.A1(new_n812_), .A2(new_n781_), .ZN(new_n6686_));
  OAI21_X1   g6301(.A1(new_n389_), .A2(new_n6686_), .B(new_n787_), .ZN(new_n6687_));
  AOI21_X1   g6302(.A1(new_n6687_), .A2(new_n1524_), .B(new_n1525_), .ZN(new_n6688_));
  OAI21_X1   g6303(.A1(new_n6688_), .A2(new_n802_), .B(new_n1607_), .ZN(new_n6689_));
  AOI21_X1   g6304(.A1(new_n6689_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n6690_));
  OAI21_X1   g6305(.A1(new_n6690_), .A2(new_n900_), .B(new_n908_), .ZN(new_n6691_));
  AOI21_X1   g6306(.A1(new_n6691_), .A2(new_n913_), .B(new_n918_), .ZN(new_n6692_));
  OAI21_X1   g6307(.A1(new_n6692_), .A2(new_n897_), .B(new_n923_), .ZN(new_n6693_));
  AOI21_X1   g6308(.A1(new_n6693_), .A2(new_n894_), .B(new_n929_), .ZN(new_n6694_));
  OAI21_X1   g6309(.A1(new_n6694_), .A2(new_n933_), .B(new_n937_), .ZN(new_n6695_));
  AOI21_X1   g6310(.A1(new_n6695_), .A2(new_n890_), .B(new_n943_), .ZN(new_n6696_));
  OAI21_X1   g6311(.A1(new_n6696_), .A2(new_n886_), .B(new_n948_), .ZN(new_n6697_));
  AOI21_X1   g6312(.A1(new_n6697_), .A2(new_n953_), .B(new_n958_), .ZN(new_n6698_));
  OAI21_X1   g6313(.A1(new_n6698_), .A2(new_n883_), .B(new_n963_), .ZN(new_n6699_));
  AOI21_X1   g6314(.A1(new_n6699_), .A2(new_n880_), .B(new_n969_), .ZN(new_n6700_));
  OAI21_X1   g6315(.A1(new_n6700_), .A2(new_n973_), .B(new_n977_), .ZN(new_n6701_));
  AOI21_X1   g6316(.A1(new_n6701_), .A2(new_n876_), .B(new_n983_), .ZN(new_n6702_));
  OAI21_X1   g6317(.A1(new_n6702_), .A2(new_n872_), .B(new_n988_), .ZN(new_n6703_));
  AOI21_X1   g6318(.A1(new_n6703_), .A2(new_n993_), .B(new_n998_), .ZN(new_n6704_));
  OAI21_X1   g6319(.A1(new_n6704_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n6705_));
  AOI21_X1   g6320(.A1(new_n6705_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n6706_));
  OAI21_X1   g6321(.A1(new_n6706_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n6707_));
  AOI21_X1   g6322(.A1(new_n6707_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n6708_));
  OAI21_X1   g6323(.A1(new_n6708_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n6709_));
  AOI21_X1   g6324(.A1(new_n6709_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n6710_));
  OAI21_X1   g6325(.A1(new_n6710_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n6711_));
  AOI21_X1   g6326(.A1(new_n6711_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n6712_));
  OAI21_X1   g6327(.A1(new_n6712_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n6713_));
  AOI21_X1   g6328(.A1(new_n6713_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n6714_));
  OAI21_X1   g6329(.A1(new_n6714_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n6715_));
  AOI21_X1   g6330(.A1(new_n6715_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n6716_));
  OAI21_X1   g6331(.A1(new_n6716_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n6717_));
  AOI21_X1   g6332(.A1(new_n6717_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n6718_));
  OAI21_X1   g6333(.A1(new_n6718_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n6719_));
  AOI21_X1   g6334(.A1(new_n6719_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n6720_));
  OAI21_X1   g6335(.A1(new_n6720_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n6721_));
  AOI21_X1   g6336(.A1(new_n6721_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n6722_));
  OAI21_X1   g6337(.A1(new_n6722_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n6723_));
  AOI21_X1   g6338(.A1(new_n6723_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n6724_));
  OAI21_X1   g6339(.A1(new_n6724_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n6725_));
  AOI21_X1   g6340(.A1(new_n6725_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n6726_));
  OAI21_X1   g6341(.A1(new_n6726_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n6727_));
  OAI21_X1   g6342(.A1(new_n1154_), .A2(\priority[117] ), .B(\req[117] ), .ZN(new_n6728_));
  AOI21_X1   g6343(.A1(new_n6727_), .A2(new_n1153_), .B(new_n6728_), .ZN(\grant[117] ));
  NOR2_X1    g6344(.A1(new_n1195_), .A2(new_n1162_), .ZN(new_n6730_));
  OAI21_X1   g6345(.A1(new_n809_), .A2(new_n6730_), .B(new_n1168_), .ZN(new_n6731_));
  AOI21_X1   g6346(.A1(new_n6731_), .A2(new_n1614_), .B(new_n1615_), .ZN(new_n6732_));
  OAI21_X1   g6347(.A1(new_n6732_), .A2(new_n1181_), .B(new_n1697_), .ZN(new_n6733_));
  AOI21_X1   g6348(.A1(new_n6733_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n6734_));
  OAI21_X1   g6349(.A1(new_n6734_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n6735_));
  AOI21_X1   g6350(.A1(new_n6735_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n6736_));
  OAI21_X1   g6351(.A1(new_n6736_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n6737_));
  AOI21_X1   g6352(.A1(new_n6737_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n6738_));
  OAI21_X1   g6353(.A1(new_n6738_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n6739_));
  AOI21_X1   g6354(.A1(new_n6739_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n6740_));
  OAI21_X1   g6355(.A1(new_n6740_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n6741_));
  AOI21_X1   g6356(.A1(new_n6741_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n6742_));
  OAI21_X1   g6357(.A1(new_n6742_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n6743_));
  AOI21_X1   g6358(.A1(new_n6743_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n6744_));
  OAI21_X1   g6359(.A1(new_n6744_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n6745_));
  AOI21_X1   g6360(.A1(new_n6745_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n6746_));
  OAI21_X1   g6361(.A1(new_n6746_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n6747_));
  AOI21_X1   g6362(.A1(new_n6747_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n6748_));
  OAI21_X1   g6363(.A1(new_n6748_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n6749_));
  AOI21_X1   g6364(.A1(new_n6749_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n6750_));
  OAI21_X1   g6365(.A1(new_n6750_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n6751_));
  AOI21_X1   g6366(.A1(new_n6751_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n6752_));
  OAI21_X1   g6367(.A1(new_n6752_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n6753_));
  AOI21_X1   g6368(.A1(new_n6753_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n6754_));
  OAI21_X1   g6369(.A1(new_n6754_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n6755_));
  AOI21_X1   g6370(.A1(new_n6755_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n6756_));
  OAI21_X1   g6371(.A1(new_n6756_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n6757_));
  AOI21_X1   g6372(.A1(new_n6757_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n6758_));
  OAI21_X1   g6373(.A1(new_n6758_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n6759_));
  AOI21_X1   g6374(.A1(new_n6759_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n6760_));
  OAI21_X1   g6375(.A1(new_n6760_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n6761_));
  AOI21_X1   g6376(.A1(new_n6761_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n6762_));
  OAI21_X1   g6377(.A1(new_n6762_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n6763_));
  AOI21_X1   g6378(.A1(new_n6763_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n6764_));
  OAI21_X1   g6379(.A1(new_n6764_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n6765_));
  AOI21_X1   g6380(.A1(new_n6765_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n6766_));
  OAI21_X1   g6381(.A1(new_n6766_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n6767_));
  AOI21_X1   g6382(.A1(new_n6767_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n6768_));
  OAI21_X1   g6383(.A1(new_n6768_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n6769_));
  AOI21_X1   g6384(.A1(new_n6769_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n6770_));
  OAI21_X1   g6385(.A1(new_n6770_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n6771_));
  OAI21_X1   g6386(.A1(new_n392_), .A2(\priority[118] ), .B(\req[118] ), .ZN(new_n6772_));
  AOI21_X1   g6387(.A1(new_n6771_), .A2(new_n1497_), .B(new_n6772_), .ZN(\grant[118] ));
  NOR2_X1    g6388(.A1(new_n388_), .A2(new_n1504_), .ZN(new_n6774_));
  OAI21_X1   g6389(.A1(new_n1192_), .A2(new_n6774_), .B(new_n1509_), .ZN(new_n6775_));
  AOI21_X1   g6390(.A1(new_n6775_), .A2(new_n1702_), .B(new_n1703_), .ZN(new_n6776_));
  OAI21_X1   g6391(.A1(new_n6776_), .A2(new_n1188_), .B(new_n1784_), .ZN(new_n6777_));
  AOI21_X1   g6392(.A1(new_n6777_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n6778_));
  OAI21_X1   g6393(.A1(new_n6778_), .A2(new_n519_), .B(new_n524_), .ZN(new_n6779_));
  AOI21_X1   g6394(.A1(new_n6779_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n6780_));
  OAI21_X1   g6395(.A1(new_n6780_), .A2(new_n497_), .B(new_n535_), .ZN(new_n6781_));
  AOI21_X1   g6396(.A1(new_n6781_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n6782_));
  OAI21_X1   g6397(.A1(new_n6782_), .A2(new_n492_), .B(new_n550_), .ZN(new_n6783_));
  AOI21_X1   g6398(.A1(new_n6783_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n6784_));
  OAI21_X1   g6399(.A1(new_n6784_), .A2(new_n561_), .B(new_n566_), .ZN(new_n6785_));
  AOI21_X1   g6400(.A1(new_n6785_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n6786_));
  OAI21_X1   g6401(.A1(new_n6786_), .A2(new_n479_), .B(new_n577_), .ZN(new_n6787_));
  AOI21_X1   g6402(.A1(new_n6787_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n6788_));
  OAI21_X1   g6403(.A1(new_n6788_), .A2(new_n474_), .B(new_n592_), .ZN(new_n6789_));
  AOI21_X1   g6404(.A1(new_n6789_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n6790_));
  OAI21_X1   g6405(.A1(new_n6790_), .A2(new_n603_), .B(new_n608_), .ZN(new_n6791_));
  AOI21_X1   g6406(.A1(new_n6791_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n6792_));
  OAI21_X1   g6407(.A1(new_n6792_), .A2(new_n461_), .B(new_n619_), .ZN(new_n6793_));
  AOI21_X1   g6408(.A1(new_n6793_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n6794_));
  OAI21_X1   g6409(.A1(new_n6794_), .A2(new_n456_), .B(new_n634_), .ZN(new_n6795_));
  AOI21_X1   g6410(.A1(new_n6795_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n6796_));
  OAI21_X1   g6411(.A1(new_n6796_), .A2(new_n645_), .B(new_n650_), .ZN(new_n6797_));
  AOI21_X1   g6412(.A1(new_n6797_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n6798_));
  OAI21_X1   g6413(.A1(new_n6798_), .A2(new_n443_), .B(new_n661_), .ZN(new_n6799_));
  AOI21_X1   g6414(.A1(new_n6799_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n6800_));
  OAI21_X1   g6415(.A1(new_n6800_), .A2(new_n438_), .B(new_n676_), .ZN(new_n6801_));
  AOI21_X1   g6416(.A1(new_n6801_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n6802_));
  OAI21_X1   g6417(.A1(new_n6802_), .A2(new_n687_), .B(new_n692_), .ZN(new_n6803_));
  AOI21_X1   g6418(.A1(new_n6803_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n6804_));
  OAI21_X1   g6419(.A1(new_n6804_), .A2(new_n425_), .B(new_n703_), .ZN(new_n6805_));
  AOI21_X1   g6420(.A1(new_n6805_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n6806_));
  OAI21_X1   g6421(.A1(new_n6806_), .A2(new_n420_), .B(new_n718_), .ZN(new_n6807_));
  AOI21_X1   g6422(.A1(new_n6807_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n6808_));
  OAI21_X1   g6423(.A1(new_n6808_), .A2(new_n729_), .B(new_n734_), .ZN(new_n6809_));
  AOI21_X1   g6424(.A1(new_n6809_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n6810_));
  OAI21_X1   g6425(.A1(new_n6810_), .A2(new_n407_), .B(new_n745_), .ZN(new_n6811_));
  AOI21_X1   g6426(.A1(new_n6811_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n6812_));
  OAI21_X1   g6427(.A1(new_n6812_), .A2(new_n402_), .B(new_n760_), .ZN(new_n6813_));
  AOI21_X1   g6428(.A1(new_n6813_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n6814_));
  OAI21_X1   g6429(.A1(new_n6814_), .A2(new_n771_), .B(new_n776_), .ZN(new_n6815_));
  OAI21_X1   g6430(.A1(new_n779_), .A2(\priority[119] ), .B(\req[119] ), .ZN(new_n6816_));
  AOI21_X1   g6431(.A1(new_n6815_), .A2(new_n1526_), .B(new_n6816_), .ZN(\grant[119] ));
  NOR2_X1    g6432(.A1(new_n808_), .A2(new_n786_), .ZN(new_n6818_));
  OAI21_X1   g6433(.A1(new_n793_), .A2(new_n6818_), .B(new_n797_), .ZN(new_n6819_));
  AOI21_X1   g6434(.A1(new_n6819_), .A2(new_n803_), .B(new_n1789_), .ZN(new_n6820_));
  OAI21_X1   g6435(.A1(new_n6820_), .A2(new_n1522_), .B(new_n1832_), .ZN(new_n6821_));
  AOI21_X1   g6436(.A1(new_n6821_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n6822_));
  OAI21_X1   g6437(.A1(new_n6822_), .A2(new_n912_), .B(new_n917_), .ZN(new_n6823_));
  AOI21_X1   g6438(.A1(new_n6823_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n6824_));
  OAI21_X1   g6439(.A1(new_n6824_), .A2(new_n893_), .B(new_n928_), .ZN(new_n6825_));
  AOI21_X1   g6440(.A1(new_n6825_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n6826_));
  OAI21_X1   g6441(.A1(new_n6826_), .A2(new_n889_), .B(new_n942_), .ZN(new_n6827_));
  AOI21_X1   g6442(.A1(new_n6827_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n6828_));
  OAI21_X1   g6443(.A1(new_n6828_), .A2(new_n952_), .B(new_n957_), .ZN(new_n6829_));
  AOI21_X1   g6444(.A1(new_n6829_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n6830_));
  OAI21_X1   g6445(.A1(new_n6830_), .A2(new_n879_), .B(new_n968_), .ZN(new_n6831_));
  AOI21_X1   g6446(.A1(new_n6831_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n6832_));
  OAI21_X1   g6447(.A1(new_n6832_), .A2(new_n875_), .B(new_n982_), .ZN(new_n6833_));
  AOI21_X1   g6448(.A1(new_n6833_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n6834_));
  OAI21_X1   g6449(.A1(new_n6834_), .A2(new_n992_), .B(new_n997_), .ZN(new_n6835_));
  AOI21_X1   g6450(.A1(new_n6835_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n6836_));
  OAI21_X1   g6451(.A1(new_n6836_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n6837_));
  AOI21_X1   g6452(.A1(new_n6837_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n6838_));
  OAI21_X1   g6453(.A1(new_n6838_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n6839_));
  AOI21_X1   g6454(.A1(new_n6839_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n6840_));
  OAI21_X1   g6455(.A1(new_n6840_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n6841_));
  AOI21_X1   g6456(.A1(new_n6841_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n6842_));
  OAI21_X1   g6457(.A1(new_n6842_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n6843_));
  AOI21_X1   g6458(.A1(new_n6843_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n6844_));
  OAI21_X1   g6459(.A1(new_n6844_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n6845_));
  AOI21_X1   g6460(.A1(new_n6845_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n6846_));
  OAI21_X1   g6461(.A1(new_n6846_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n6847_));
  AOI21_X1   g6462(.A1(new_n6847_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n6848_));
  OAI21_X1   g6463(.A1(new_n6848_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n6849_));
  AOI21_X1   g6464(.A1(new_n6849_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n6850_));
  OAI21_X1   g6465(.A1(new_n6850_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n6851_));
  AOI21_X1   g6466(.A1(new_n6851_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n6852_));
  OAI21_X1   g6467(.A1(new_n6852_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n6853_));
  AOI21_X1   g6468(.A1(new_n6853_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n6854_));
  OAI21_X1   g6469(.A1(new_n6854_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n6855_));
  AOI21_X1   g6470(.A1(new_n6855_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n6856_));
  OAI21_X1   g6471(.A1(new_n6856_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n6857_));
  AOI21_X1   g6472(.A1(new_n6857_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n6858_));
  OAI21_X1   g6473(.A1(new_n6858_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n6859_));
  OAI21_X1   g6474(.A1(new_n1160_), .A2(\priority[120] ), .B(\req[120] ), .ZN(new_n6860_));
  AOI21_X1   g6475(.A1(new_n6859_), .A2(new_n1616_), .B(new_n6860_), .ZN(\grant[120] ));
  NOR2_X1    g6476(.A1(new_n1191_), .A2(new_n1167_), .ZN(new_n6862_));
  OAI21_X1   g6477(.A1(new_n1173_), .A2(new_n6862_), .B(new_n1177_), .ZN(new_n6863_));
  AOI21_X1   g6478(.A1(new_n6863_), .A2(new_n1182_), .B(new_n1837_), .ZN(new_n6864_));
  OAI21_X1   g6479(.A1(new_n6864_), .A2(new_n1612_), .B(new_n1880_), .ZN(new_n6865_));
  AOI21_X1   g6480(.A1(new_n6865_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n6866_));
  OAI21_X1   g6481(.A1(new_n6866_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n6867_));
  AOI21_X1   g6482(.A1(new_n6867_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n6868_));
  OAI21_X1   g6483(.A1(new_n6868_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n6869_));
  AOI21_X1   g6484(.A1(new_n6869_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n6870_));
  OAI21_X1   g6485(.A1(new_n6870_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n6871_));
  AOI21_X1   g6486(.A1(new_n6871_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n6872_));
  OAI21_X1   g6487(.A1(new_n6872_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n6873_));
  AOI21_X1   g6488(.A1(new_n6873_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n6874_));
  OAI21_X1   g6489(.A1(new_n6874_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n6875_));
  AOI21_X1   g6490(.A1(new_n6875_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n6876_));
  OAI21_X1   g6491(.A1(new_n6876_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n6877_));
  AOI21_X1   g6492(.A1(new_n6877_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n6878_));
  OAI21_X1   g6493(.A1(new_n6878_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n6879_));
  AOI21_X1   g6494(.A1(new_n6879_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n6880_));
  OAI21_X1   g6495(.A1(new_n6880_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n6881_));
  AOI21_X1   g6496(.A1(new_n6881_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n6882_));
  OAI21_X1   g6497(.A1(new_n6882_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n6883_));
  AOI21_X1   g6498(.A1(new_n6883_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n6884_));
  OAI21_X1   g6499(.A1(new_n6884_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n6885_));
  AOI21_X1   g6500(.A1(new_n6885_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n6886_));
  OAI21_X1   g6501(.A1(new_n6886_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n6887_));
  AOI21_X1   g6502(.A1(new_n6887_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n6888_));
  OAI21_X1   g6503(.A1(new_n6888_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n6889_));
  AOI21_X1   g6504(.A1(new_n6889_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n6890_));
  OAI21_X1   g6505(.A1(new_n6890_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n6891_));
  AOI21_X1   g6506(.A1(new_n6891_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n6892_));
  OAI21_X1   g6507(.A1(new_n6892_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n6893_));
  AOI21_X1   g6508(.A1(new_n6893_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n6894_));
  OAI21_X1   g6509(.A1(new_n6894_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n6895_));
  AOI21_X1   g6510(.A1(new_n6895_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n6896_));
  OAI21_X1   g6511(.A1(new_n6896_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n6897_));
  AOI21_X1   g6512(.A1(new_n6897_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n6898_));
  OAI21_X1   g6513(.A1(new_n6898_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n6899_));
  AOI21_X1   g6514(.A1(new_n6899_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n6900_));
  OAI21_X1   g6515(.A1(new_n6900_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n6901_));
  AOI21_X1   g6516(.A1(new_n6901_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n6902_));
  OAI21_X1   g6517(.A1(new_n6902_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n6903_));
  OAI21_X1   g6518(.A1(new_n387_), .A2(\priority[121] ), .B(\req[121] ), .ZN(new_n6904_));
  AOI21_X1   g6519(.A1(new_n6903_), .A2(new_n1704_), .B(new_n6904_), .ZN(\grant[121] ));
  NOR2_X1    g6520(.A1(new_n792_), .A2(new_n1508_), .ZN(new_n6906_));
  OAI21_X1   g6521(.A1(new_n1514_), .A2(new_n6906_), .B(new_n1517_), .ZN(new_n6907_));
  AOI21_X1   g6522(.A1(new_n6907_), .A2(new_n1189_), .B(new_n1884_), .ZN(new_n6908_));
  OAI21_X1   g6523(.A1(new_n6908_), .A2(new_n506_), .B(new_n514_), .ZN(new_n6909_));
  AOI21_X1   g6524(.A1(new_n6909_), .A2(new_n520_), .B(new_n525_), .ZN(new_n6910_));
  OAI21_X1   g6525(.A1(new_n6910_), .A2(new_n502_), .B(new_n530_), .ZN(new_n6911_));
  AOI21_X1   g6526(.A1(new_n6911_), .A2(new_n498_), .B(new_n536_), .ZN(new_n6912_));
  OAI21_X1   g6527(.A1(new_n6912_), .A2(new_n541_), .B(new_n545_), .ZN(new_n6913_));
  AOI21_X1   g6528(.A1(new_n6913_), .A2(new_n493_), .B(new_n551_), .ZN(new_n6914_));
  OAI21_X1   g6529(.A1(new_n6914_), .A2(new_n488_), .B(new_n556_), .ZN(new_n6915_));
  AOI21_X1   g6530(.A1(new_n6915_), .A2(new_n562_), .B(new_n567_), .ZN(new_n6916_));
  OAI21_X1   g6531(.A1(new_n6916_), .A2(new_n484_), .B(new_n572_), .ZN(new_n6917_));
  AOI21_X1   g6532(.A1(new_n6917_), .A2(new_n480_), .B(new_n578_), .ZN(new_n6918_));
  OAI21_X1   g6533(.A1(new_n6918_), .A2(new_n583_), .B(new_n587_), .ZN(new_n6919_));
  AOI21_X1   g6534(.A1(new_n6919_), .A2(new_n475_), .B(new_n593_), .ZN(new_n6920_));
  OAI21_X1   g6535(.A1(new_n6920_), .A2(new_n470_), .B(new_n598_), .ZN(new_n6921_));
  AOI21_X1   g6536(.A1(new_n6921_), .A2(new_n604_), .B(new_n609_), .ZN(new_n6922_));
  OAI21_X1   g6537(.A1(new_n6922_), .A2(new_n466_), .B(new_n614_), .ZN(new_n6923_));
  AOI21_X1   g6538(.A1(new_n6923_), .A2(new_n462_), .B(new_n620_), .ZN(new_n6924_));
  OAI21_X1   g6539(.A1(new_n6924_), .A2(new_n625_), .B(new_n629_), .ZN(new_n6925_));
  AOI21_X1   g6540(.A1(new_n6925_), .A2(new_n457_), .B(new_n635_), .ZN(new_n6926_));
  OAI21_X1   g6541(.A1(new_n6926_), .A2(new_n452_), .B(new_n640_), .ZN(new_n6927_));
  AOI21_X1   g6542(.A1(new_n6927_), .A2(new_n646_), .B(new_n651_), .ZN(new_n6928_));
  OAI21_X1   g6543(.A1(new_n6928_), .A2(new_n448_), .B(new_n656_), .ZN(new_n6929_));
  AOI21_X1   g6544(.A1(new_n6929_), .A2(new_n444_), .B(new_n662_), .ZN(new_n6930_));
  OAI21_X1   g6545(.A1(new_n6930_), .A2(new_n667_), .B(new_n671_), .ZN(new_n6931_));
  AOI21_X1   g6546(.A1(new_n6931_), .A2(new_n439_), .B(new_n677_), .ZN(new_n6932_));
  OAI21_X1   g6547(.A1(new_n6932_), .A2(new_n434_), .B(new_n682_), .ZN(new_n6933_));
  AOI21_X1   g6548(.A1(new_n6933_), .A2(new_n688_), .B(new_n693_), .ZN(new_n6934_));
  OAI21_X1   g6549(.A1(new_n6934_), .A2(new_n430_), .B(new_n698_), .ZN(new_n6935_));
  AOI21_X1   g6550(.A1(new_n6935_), .A2(new_n426_), .B(new_n704_), .ZN(new_n6936_));
  OAI21_X1   g6551(.A1(new_n6936_), .A2(new_n709_), .B(new_n713_), .ZN(new_n6937_));
  AOI21_X1   g6552(.A1(new_n6937_), .A2(new_n421_), .B(new_n719_), .ZN(new_n6938_));
  OAI21_X1   g6553(.A1(new_n6938_), .A2(new_n416_), .B(new_n724_), .ZN(new_n6939_));
  AOI21_X1   g6554(.A1(new_n6939_), .A2(new_n730_), .B(new_n735_), .ZN(new_n6940_));
  OAI21_X1   g6555(.A1(new_n6940_), .A2(new_n412_), .B(new_n740_), .ZN(new_n6941_));
  AOI21_X1   g6556(.A1(new_n6941_), .A2(new_n408_), .B(new_n746_), .ZN(new_n6942_));
  OAI21_X1   g6557(.A1(new_n6942_), .A2(new_n751_), .B(new_n755_), .ZN(new_n6943_));
  AOI21_X1   g6558(.A1(new_n6943_), .A2(new_n403_), .B(new_n761_), .ZN(new_n6944_));
  OAI21_X1   g6559(.A1(new_n6944_), .A2(new_n398_), .B(new_n766_), .ZN(new_n6945_));
  AOI21_X1   g6560(.A1(new_n6945_), .A2(new_n772_), .B(new_n777_), .ZN(new_n6946_));
  OAI21_X1   g6561(.A1(new_n6946_), .A2(new_n394_), .B(new_n782_), .ZN(new_n6947_));
  OAI21_X1   g6562(.A1(new_n784_), .A2(\priority[122] ), .B(\req[122] ), .ZN(new_n6948_));
  AOI21_X1   g6563(.A1(new_n6947_), .A2(new_n390_), .B(new_n6948_), .ZN(\grant[122] ));
  NOR2_X1    g6564(.A1(new_n1172_), .A2(new_n796_), .ZN(new_n6950_));
  OAI21_X1   g6565(.A1(new_n802_), .A2(new_n6950_), .B(new_n1607_), .ZN(new_n6951_));
  AOI21_X1   g6566(.A1(new_n6951_), .A2(new_n1523_), .B(new_n1929_), .ZN(new_n6952_));
  OAI21_X1   g6567(.A1(new_n6952_), .A2(new_n900_), .B(new_n908_), .ZN(new_n6953_));
  AOI21_X1   g6568(.A1(new_n6953_), .A2(new_n913_), .B(new_n918_), .ZN(new_n6954_));
  OAI21_X1   g6569(.A1(new_n6954_), .A2(new_n897_), .B(new_n923_), .ZN(new_n6955_));
  AOI21_X1   g6570(.A1(new_n6955_), .A2(new_n894_), .B(new_n929_), .ZN(new_n6956_));
  OAI21_X1   g6571(.A1(new_n6956_), .A2(new_n933_), .B(new_n937_), .ZN(new_n6957_));
  AOI21_X1   g6572(.A1(new_n6957_), .A2(new_n890_), .B(new_n943_), .ZN(new_n6958_));
  OAI21_X1   g6573(.A1(new_n6958_), .A2(new_n886_), .B(new_n948_), .ZN(new_n6959_));
  AOI21_X1   g6574(.A1(new_n6959_), .A2(new_n953_), .B(new_n958_), .ZN(new_n6960_));
  OAI21_X1   g6575(.A1(new_n6960_), .A2(new_n883_), .B(new_n963_), .ZN(new_n6961_));
  AOI21_X1   g6576(.A1(new_n6961_), .A2(new_n880_), .B(new_n969_), .ZN(new_n6962_));
  OAI21_X1   g6577(.A1(new_n6962_), .A2(new_n973_), .B(new_n977_), .ZN(new_n6963_));
  AOI21_X1   g6578(.A1(new_n6963_), .A2(new_n876_), .B(new_n983_), .ZN(new_n6964_));
  OAI21_X1   g6579(.A1(new_n6964_), .A2(new_n872_), .B(new_n988_), .ZN(new_n6965_));
  AOI21_X1   g6580(.A1(new_n6965_), .A2(new_n993_), .B(new_n998_), .ZN(new_n6966_));
  OAI21_X1   g6581(.A1(new_n6966_), .A2(new_n869_), .B(new_n1003_), .ZN(new_n6967_));
  AOI21_X1   g6582(.A1(new_n6967_), .A2(new_n866_), .B(new_n1009_), .ZN(new_n6968_));
  OAI21_X1   g6583(.A1(new_n6968_), .A2(new_n1013_), .B(new_n1017_), .ZN(new_n6969_));
  AOI21_X1   g6584(.A1(new_n6969_), .A2(new_n862_), .B(new_n1023_), .ZN(new_n6970_));
  OAI21_X1   g6585(.A1(new_n6970_), .A2(new_n858_), .B(new_n1028_), .ZN(new_n6971_));
  AOI21_X1   g6586(.A1(new_n6971_), .A2(new_n1033_), .B(new_n1038_), .ZN(new_n6972_));
  OAI21_X1   g6587(.A1(new_n6972_), .A2(new_n855_), .B(new_n1043_), .ZN(new_n6973_));
  AOI21_X1   g6588(.A1(new_n6973_), .A2(new_n852_), .B(new_n1049_), .ZN(new_n6974_));
  OAI21_X1   g6589(.A1(new_n6974_), .A2(new_n1053_), .B(new_n1057_), .ZN(new_n6975_));
  AOI21_X1   g6590(.A1(new_n6975_), .A2(new_n848_), .B(new_n1063_), .ZN(new_n6976_));
  OAI21_X1   g6591(.A1(new_n6976_), .A2(new_n844_), .B(new_n1068_), .ZN(new_n6977_));
  AOI21_X1   g6592(.A1(new_n6977_), .A2(new_n1073_), .B(new_n1078_), .ZN(new_n6978_));
  OAI21_X1   g6593(.A1(new_n6978_), .A2(new_n841_), .B(new_n1083_), .ZN(new_n6979_));
  AOI21_X1   g6594(.A1(new_n6979_), .A2(new_n838_), .B(new_n1089_), .ZN(new_n6980_));
  OAI21_X1   g6595(.A1(new_n6980_), .A2(new_n1093_), .B(new_n1097_), .ZN(new_n6981_));
  AOI21_X1   g6596(.A1(new_n6981_), .A2(new_n834_), .B(new_n1103_), .ZN(new_n6982_));
  OAI21_X1   g6597(.A1(new_n6982_), .A2(new_n830_), .B(new_n1108_), .ZN(new_n6983_));
  AOI21_X1   g6598(.A1(new_n6983_), .A2(new_n1113_), .B(new_n1118_), .ZN(new_n6984_));
  OAI21_X1   g6599(.A1(new_n6984_), .A2(new_n827_), .B(new_n1123_), .ZN(new_n6985_));
  AOI21_X1   g6600(.A1(new_n6985_), .A2(new_n824_), .B(new_n1129_), .ZN(new_n6986_));
  OAI21_X1   g6601(.A1(new_n6986_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n6987_));
  AOI21_X1   g6602(.A1(new_n6987_), .A2(new_n820_), .B(new_n1143_), .ZN(new_n6988_));
  OAI21_X1   g6603(.A1(new_n6988_), .A2(new_n816_), .B(new_n1148_), .ZN(new_n6989_));
  AOI21_X1   g6604(.A1(new_n6989_), .A2(new_n1153_), .B(new_n1158_), .ZN(new_n6990_));
  OAI21_X1   g6605(.A1(new_n6990_), .A2(new_n813_), .B(new_n1163_), .ZN(new_n6991_));
  OAI21_X1   g6606(.A1(new_n1165_), .A2(\priority[123] ), .B(\req[123] ), .ZN(new_n6992_));
  AOI21_X1   g6607(.A1(new_n6991_), .A2(new_n810_), .B(new_n6992_), .ZN(\grant[123] ));
  NOR2_X1    g6608(.A1(new_n1513_), .A2(new_n1176_), .ZN(new_n6994_));
  OAI21_X1   g6609(.A1(new_n1181_), .A2(new_n6994_), .B(new_n1697_), .ZN(new_n6995_));
  AOI21_X1   g6610(.A1(new_n6995_), .A2(new_n1613_), .B(new_n1974_), .ZN(new_n6996_));
  OAI21_X1   g6611(.A1(new_n6996_), .A2(new_n1283_), .B(new_n1288_), .ZN(new_n6997_));
  AOI21_X1   g6612(.A1(new_n6997_), .A2(new_n1293_), .B(new_n1297_), .ZN(new_n6998_));
  OAI21_X1   g6613(.A1(new_n6998_), .A2(new_n1280_), .B(new_n1301_), .ZN(new_n6999_));
  AOI21_X1   g6614(.A1(new_n6999_), .A2(new_n1277_), .B(new_n1306_), .ZN(new_n7000_));
  OAI21_X1   g6615(.A1(new_n7000_), .A2(new_n1310_), .B(new_n1313_), .ZN(new_n7001_));
  AOI21_X1   g6616(.A1(new_n7001_), .A2(new_n1273_), .B(new_n1318_), .ZN(new_n7002_));
  OAI21_X1   g6617(.A1(new_n7002_), .A2(new_n1269_), .B(new_n1322_), .ZN(new_n7003_));
  AOI21_X1   g6618(.A1(new_n7003_), .A2(new_n1327_), .B(new_n1331_), .ZN(new_n7004_));
  OAI21_X1   g6619(.A1(new_n7004_), .A2(new_n1266_), .B(new_n1335_), .ZN(new_n7005_));
  AOI21_X1   g6620(.A1(new_n7005_), .A2(new_n1263_), .B(new_n1340_), .ZN(new_n7006_));
  OAI21_X1   g6621(.A1(new_n7006_), .A2(new_n1344_), .B(new_n1347_), .ZN(new_n7007_));
  AOI21_X1   g6622(.A1(new_n7007_), .A2(new_n1259_), .B(new_n1352_), .ZN(new_n7008_));
  OAI21_X1   g6623(.A1(new_n7008_), .A2(new_n1255_), .B(new_n1356_), .ZN(new_n7009_));
  AOI21_X1   g6624(.A1(new_n7009_), .A2(new_n1361_), .B(new_n1365_), .ZN(new_n7010_));
  OAI21_X1   g6625(.A1(new_n7010_), .A2(new_n1252_), .B(new_n1369_), .ZN(new_n7011_));
  AOI21_X1   g6626(.A1(new_n7011_), .A2(new_n1249_), .B(new_n1374_), .ZN(new_n7012_));
  OAI21_X1   g6627(.A1(new_n7012_), .A2(new_n1378_), .B(new_n1381_), .ZN(new_n7013_));
  AOI21_X1   g6628(.A1(new_n7013_), .A2(new_n1245_), .B(new_n1386_), .ZN(new_n7014_));
  OAI21_X1   g6629(.A1(new_n7014_), .A2(new_n1241_), .B(new_n1390_), .ZN(new_n7015_));
  AOI21_X1   g6630(.A1(new_n7015_), .A2(new_n1395_), .B(new_n1399_), .ZN(new_n7016_));
  OAI21_X1   g6631(.A1(new_n7016_), .A2(new_n1238_), .B(new_n1403_), .ZN(new_n7017_));
  AOI21_X1   g6632(.A1(new_n7017_), .A2(new_n1235_), .B(new_n1408_), .ZN(new_n7018_));
  OAI21_X1   g6633(.A1(new_n7018_), .A2(new_n1412_), .B(new_n1415_), .ZN(new_n7019_));
  AOI21_X1   g6634(.A1(new_n7019_), .A2(new_n1231_), .B(new_n1420_), .ZN(new_n7020_));
  OAI21_X1   g6635(.A1(new_n7020_), .A2(new_n1227_), .B(new_n1424_), .ZN(new_n7021_));
  AOI21_X1   g6636(.A1(new_n7021_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n7022_));
  OAI21_X1   g6637(.A1(new_n7022_), .A2(new_n1224_), .B(new_n1437_), .ZN(new_n7023_));
  AOI21_X1   g6638(.A1(new_n7023_), .A2(new_n1221_), .B(new_n1442_), .ZN(new_n7024_));
  OAI21_X1   g6639(.A1(new_n7024_), .A2(new_n1446_), .B(new_n1449_), .ZN(new_n7025_));
  AOI21_X1   g6640(.A1(new_n7025_), .A2(new_n1217_), .B(new_n1454_), .ZN(new_n7026_));
  OAI21_X1   g6641(.A1(new_n7026_), .A2(new_n1213_), .B(new_n1458_), .ZN(new_n7027_));
  AOI21_X1   g6642(.A1(new_n7027_), .A2(new_n1463_), .B(new_n1467_), .ZN(new_n7028_));
  OAI21_X1   g6643(.A1(new_n7028_), .A2(new_n1210_), .B(new_n1471_), .ZN(new_n7029_));
  AOI21_X1   g6644(.A1(new_n7029_), .A2(new_n1207_), .B(new_n1476_), .ZN(new_n7030_));
  OAI21_X1   g6645(.A1(new_n7030_), .A2(new_n1480_), .B(new_n1483_), .ZN(new_n7031_));
  AOI21_X1   g6646(.A1(new_n7031_), .A2(new_n1203_), .B(new_n1488_), .ZN(new_n7032_));
  OAI21_X1   g6647(.A1(new_n7032_), .A2(new_n1199_), .B(new_n1492_), .ZN(new_n7033_));
  AOI21_X1   g6648(.A1(new_n7033_), .A2(new_n1497_), .B(new_n1501_), .ZN(new_n7034_));
  OAI21_X1   g6649(.A1(new_n7034_), .A2(new_n1196_), .B(new_n1505_), .ZN(new_n7035_));
  OAI21_X1   g6650(.A1(new_n791_), .A2(\priority[124] ), .B(\req[124] ), .ZN(new_n7036_));
  AOI21_X1   g6651(.A1(new_n7035_), .A2(new_n1193_), .B(new_n7036_), .ZN(\grant[124] ));
  NOR2_X1    g6652(.A1(new_n801_), .A2(new_n1516_), .ZN(new_n7038_));
  OAI21_X1   g6653(.A1(new_n1188_), .A2(new_n7038_), .B(new_n1784_), .ZN(new_n7039_));
  AOI21_X1   g6654(.A1(new_n7039_), .A2(new_n1701_), .B(new_n2019_), .ZN(new_n7040_));
  OAI21_X1   g6655(.A1(new_n7040_), .A2(new_n519_), .B(new_n524_), .ZN(new_n7041_));
  AOI21_X1   g6656(.A1(new_n7041_), .A2(new_n1562_), .B(new_n1563_), .ZN(new_n7042_));
  OAI21_X1   g6657(.A1(new_n7042_), .A2(new_n497_), .B(new_n535_), .ZN(new_n7043_));
  AOI21_X1   g6658(.A1(new_n7043_), .A2(new_n1560_), .B(new_n1561_), .ZN(new_n7044_));
  OAI21_X1   g6659(.A1(new_n7044_), .A2(new_n492_), .B(new_n550_), .ZN(new_n7045_));
  AOI21_X1   g6660(.A1(new_n7045_), .A2(new_n1558_), .B(new_n1559_), .ZN(new_n7046_));
  OAI21_X1   g6661(.A1(new_n7046_), .A2(new_n561_), .B(new_n566_), .ZN(new_n7047_));
  AOI21_X1   g6662(.A1(new_n7047_), .A2(new_n1556_), .B(new_n1557_), .ZN(new_n7048_));
  OAI21_X1   g6663(.A1(new_n7048_), .A2(new_n479_), .B(new_n577_), .ZN(new_n7049_));
  AOI21_X1   g6664(.A1(new_n7049_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n7050_));
  OAI21_X1   g6665(.A1(new_n7050_), .A2(new_n474_), .B(new_n592_), .ZN(new_n7051_));
  AOI21_X1   g6666(.A1(new_n7051_), .A2(new_n1552_), .B(new_n1553_), .ZN(new_n7052_));
  OAI21_X1   g6667(.A1(new_n7052_), .A2(new_n603_), .B(new_n608_), .ZN(new_n7053_));
  AOI21_X1   g6668(.A1(new_n7053_), .A2(new_n1550_), .B(new_n1551_), .ZN(new_n7054_));
  OAI21_X1   g6669(.A1(new_n7054_), .A2(new_n461_), .B(new_n619_), .ZN(new_n7055_));
  AOI21_X1   g6670(.A1(new_n7055_), .A2(new_n1548_), .B(new_n1549_), .ZN(new_n7056_));
  OAI21_X1   g6671(.A1(new_n7056_), .A2(new_n456_), .B(new_n634_), .ZN(new_n7057_));
  AOI21_X1   g6672(.A1(new_n7057_), .A2(new_n1546_), .B(new_n1547_), .ZN(new_n7058_));
  OAI21_X1   g6673(.A1(new_n7058_), .A2(new_n645_), .B(new_n650_), .ZN(new_n7059_));
  AOI21_X1   g6674(.A1(new_n7059_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n7060_));
  OAI21_X1   g6675(.A1(new_n7060_), .A2(new_n443_), .B(new_n661_), .ZN(new_n7061_));
  AOI21_X1   g6676(.A1(new_n7061_), .A2(new_n1542_), .B(new_n1543_), .ZN(new_n7062_));
  OAI21_X1   g6677(.A1(new_n7062_), .A2(new_n438_), .B(new_n676_), .ZN(new_n7063_));
  AOI21_X1   g6678(.A1(new_n7063_), .A2(new_n1540_), .B(new_n1541_), .ZN(new_n7064_));
  OAI21_X1   g6679(.A1(new_n7064_), .A2(new_n687_), .B(new_n692_), .ZN(new_n7065_));
  AOI21_X1   g6680(.A1(new_n7065_), .A2(new_n1538_), .B(new_n1539_), .ZN(new_n7066_));
  OAI21_X1   g6681(.A1(new_n7066_), .A2(new_n425_), .B(new_n703_), .ZN(new_n7067_));
  AOI21_X1   g6682(.A1(new_n7067_), .A2(new_n1536_), .B(new_n1537_), .ZN(new_n7068_));
  OAI21_X1   g6683(.A1(new_n7068_), .A2(new_n420_), .B(new_n718_), .ZN(new_n7069_));
  AOI21_X1   g6684(.A1(new_n7069_), .A2(new_n1534_), .B(new_n1535_), .ZN(new_n7070_));
  OAI21_X1   g6685(.A1(new_n7070_), .A2(new_n729_), .B(new_n734_), .ZN(new_n7071_));
  AOI21_X1   g6686(.A1(new_n7071_), .A2(new_n1532_), .B(new_n1533_), .ZN(new_n7072_));
  OAI21_X1   g6687(.A1(new_n7072_), .A2(new_n407_), .B(new_n745_), .ZN(new_n7073_));
  AOI21_X1   g6688(.A1(new_n7073_), .A2(new_n1530_), .B(new_n1531_), .ZN(new_n7074_));
  OAI21_X1   g6689(.A1(new_n7074_), .A2(new_n402_), .B(new_n760_), .ZN(new_n7075_));
  AOI21_X1   g6690(.A1(new_n7075_), .A2(new_n1528_), .B(new_n1529_), .ZN(new_n7076_));
  OAI21_X1   g6691(.A1(new_n7076_), .A2(new_n771_), .B(new_n776_), .ZN(new_n7077_));
  AOI21_X1   g6692(.A1(new_n7077_), .A2(new_n1526_), .B(new_n1527_), .ZN(new_n7078_));
  OAI21_X1   g6693(.A1(new_n7078_), .A2(new_n389_), .B(new_n787_), .ZN(new_n7079_));
  OAI21_X1   g6694(.A1(new_n794_), .A2(\priority[125] ), .B(\req[125] ), .ZN(new_n7080_));
  AOI21_X1   g6695(.A1(new_n7079_), .A2(new_n1524_), .B(new_n7080_), .ZN(\grant[125] ));
  NOR2_X1    g6696(.A1(new_n1180_), .A2(new_n1606_), .ZN(new_n7082_));
  OAI21_X1   g6697(.A1(new_n1522_), .A2(new_n7082_), .B(new_n1832_), .ZN(new_n7083_));
  AOI21_X1   g6698(.A1(new_n7083_), .A2(new_n1788_), .B(new_n2064_), .ZN(new_n7084_));
  OAI21_X1   g6699(.A1(new_n7084_), .A2(new_n912_), .B(new_n917_), .ZN(new_n7085_));
  AOI21_X1   g6700(.A1(new_n7085_), .A2(new_n1652_), .B(new_n1653_), .ZN(new_n7086_));
  OAI21_X1   g6701(.A1(new_n7086_), .A2(new_n893_), .B(new_n928_), .ZN(new_n7087_));
  AOI21_X1   g6702(.A1(new_n7087_), .A2(new_n1650_), .B(new_n1651_), .ZN(new_n7088_));
  OAI21_X1   g6703(.A1(new_n7088_), .A2(new_n889_), .B(new_n942_), .ZN(new_n7089_));
  AOI21_X1   g6704(.A1(new_n7089_), .A2(new_n1648_), .B(new_n1649_), .ZN(new_n7090_));
  OAI21_X1   g6705(.A1(new_n7090_), .A2(new_n952_), .B(new_n957_), .ZN(new_n7091_));
  AOI21_X1   g6706(.A1(new_n7091_), .A2(new_n1646_), .B(new_n1647_), .ZN(new_n7092_));
  OAI21_X1   g6707(.A1(new_n7092_), .A2(new_n879_), .B(new_n968_), .ZN(new_n7093_));
  AOI21_X1   g6708(.A1(new_n7093_), .A2(new_n1644_), .B(new_n1645_), .ZN(new_n7094_));
  OAI21_X1   g6709(.A1(new_n7094_), .A2(new_n875_), .B(new_n982_), .ZN(new_n7095_));
  AOI21_X1   g6710(.A1(new_n7095_), .A2(new_n1642_), .B(new_n1643_), .ZN(new_n7096_));
  OAI21_X1   g6711(.A1(new_n7096_), .A2(new_n992_), .B(new_n997_), .ZN(new_n7097_));
  AOI21_X1   g6712(.A1(new_n7097_), .A2(new_n1640_), .B(new_n1641_), .ZN(new_n7098_));
  OAI21_X1   g6713(.A1(new_n7098_), .A2(new_n865_), .B(new_n1008_), .ZN(new_n7099_));
  AOI21_X1   g6714(.A1(new_n7099_), .A2(new_n1638_), .B(new_n1639_), .ZN(new_n7100_));
  OAI21_X1   g6715(.A1(new_n7100_), .A2(new_n861_), .B(new_n1022_), .ZN(new_n7101_));
  AOI21_X1   g6716(.A1(new_n7101_), .A2(new_n1636_), .B(new_n1637_), .ZN(new_n7102_));
  OAI21_X1   g6717(.A1(new_n7102_), .A2(new_n1032_), .B(new_n1037_), .ZN(new_n7103_));
  AOI21_X1   g6718(.A1(new_n7103_), .A2(new_n1634_), .B(new_n1635_), .ZN(new_n7104_));
  OAI21_X1   g6719(.A1(new_n7104_), .A2(new_n851_), .B(new_n1048_), .ZN(new_n7105_));
  AOI21_X1   g6720(.A1(new_n7105_), .A2(new_n1632_), .B(new_n1633_), .ZN(new_n7106_));
  OAI21_X1   g6721(.A1(new_n7106_), .A2(new_n847_), .B(new_n1062_), .ZN(new_n7107_));
  AOI21_X1   g6722(.A1(new_n7107_), .A2(new_n1630_), .B(new_n1631_), .ZN(new_n7108_));
  OAI21_X1   g6723(.A1(new_n7108_), .A2(new_n1072_), .B(new_n1077_), .ZN(new_n7109_));
  AOI21_X1   g6724(.A1(new_n7109_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n7110_));
  OAI21_X1   g6725(.A1(new_n7110_), .A2(new_n837_), .B(new_n1088_), .ZN(new_n7111_));
  AOI21_X1   g6726(.A1(new_n7111_), .A2(new_n1626_), .B(new_n1627_), .ZN(new_n7112_));
  OAI21_X1   g6727(.A1(new_n7112_), .A2(new_n833_), .B(new_n1102_), .ZN(new_n7113_));
  AOI21_X1   g6728(.A1(new_n7113_), .A2(new_n1624_), .B(new_n1625_), .ZN(new_n7114_));
  OAI21_X1   g6729(.A1(new_n7114_), .A2(new_n1112_), .B(new_n1117_), .ZN(new_n7115_));
  AOI21_X1   g6730(.A1(new_n7115_), .A2(new_n1622_), .B(new_n1623_), .ZN(new_n7116_));
  OAI21_X1   g6731(.A1(new_n7116_), .A2(new_n823_), .B(new_n1128_), .ZN(new_n7117_));
  AOI21_X1   g6732(.A1(new_n7117_), .A2(new_n1620_), .B(new_n1621_), .ZN(new_n7118_));
  OAI21_X1   g6733(.A1(new_n7118_), .A2(new_n819_), .B(new_n1142_), .ZN(new_n7119_));
  AOI21_X1   g6734(.A1(new_n7119_), .A2(new_n1618_), .B(new_n1619_), .ZN(new_n7120_));
  OAI21_X1   g6735(.A1(new_n7120_), .A2(new_n1152_), .B(new_n1157_), .ZN(new_n7121_));
  AOI21_X1   g6736(.A1(new_n7121_), .A2(new_n1616_), .B(new_n1617_), .ZN(new_n7122_));
  OAI21_X1   g6737(.A1(new_n7122_), .A2(new_n809_), .B(new_n1168_), .ZN(new_n7123_));
  OAI21_X1   g6738(.A1(new_n1174_), .A2(\priority[126] ), .B(\req[126] ), .ZN(new_n7124_));
  AOI21_X1   g6739(.A1(new_n7123_), .A2(new_n1614_), .B(new_n7124_), .ZN(\grant[126] ));
  NOR2_X1    g6740(.A1(new_n1187_), .A2(new_n1696_), .ZN(new_n7126_));
  OAI21_X1   g6741(.A1(new_n1612_), .A2(new_n7126_), .B(new_n1880_), .ZN(new_n7127_));
  AOI21_X1   g6742(.A1(new_n7127_), .A2(new_n1836_), .B(new_n2109_), .ZN(new_n7128_));
  OAI21_X1   g6743(.A1(new_n7128_), .A2(new_n1292_), .B(new_n1296_), .ZN(new_n7129_));
  AOI21_X1   g6744(.A1(new_n7129_), .A2(new_n1740_), .B(new_n1741_), .ZN(new_n7130_));
  OAI21_X1   g6745(.A1(new_n7130_), .A2(new_n1276_), .B(new_n1305_), .ZN(new_n7131_));
  AOI21_X1   g6746(.A1(new_n7131_), .A2(new_n1738_), .B(new_n1739_), .ZN(new_n7132_));
  OAI21_X1   g6747(.A1(new_n7132_), .A2(new_n1272_), .B(new_n1317_), .ZN(new_n7133_));
  AOI21_X1   g6748(.A1(new_n7133_), .A2(new_n1736_), .B(new_n1737_), .ZN(new_n7134_));
  OAI21_X1   g6749(.A1(new_n7134_), .A2(new_n1326_), .B(new_n1330_), .ZN(new_n7135_));
  AOI21_X1   g6750(.A1(new_n7135_), .A2(new_n1734_), .B(new_n1735_), .ZN(new_n7136_));
  OAI21_X1   g6751(.A1(new_n7136_), .A2(new_n1262_), .B(new_n1339_), .ZN(new_n7137_));
  AOI21_X1   g6752(.A1(new_n7137_), .A2(new_n1732_), .B(new_n1733_), .ZN(new_n7138_));
  OAI21_X1   g6753(.A1(new_n7138_), .A2(new_n1258_), .B(new_n1351_), .ZN(new_n7139_));
  AOI21_X1   g6754(.A1(new_n7139_), .A2(new_n1730_), .B(new_n1731_), .ZN(new_n7140_));
  OAI21_X1   g6755(.A1(new_n7140_), .A2(new_n1360_), .B(new_n1364_), .ZN(new_n7141_));
  AOI21_X1   g6756(.A1(new_n7141_), .A2(new_n1728_), .B(new_n1729_), .ZN(new_n7142_));
  OAI21_X1   g6757(.A1(new_n7142_), .A2(new_n1248_), .B(new_n1373_), .ZN(new_n7143_));
  AOI21_X1   g6758(.A1(new_n7143_), .A2(new_n1726_), .B(new_n1727_), .ZN(new_n7144_));
  OAI21_X1   g6759(.A1(new_n7144_), .A2(new_n1244_), .B(new_n1385_), .ZN(new_n7145_));
  AOI21_X1   g6760(.A1(new_n7145_), .A2(new_n1724_), .B(new_n1725_), .ZN(new_n7146_));
  OAI21_X1   g6761(.A1(new_n7146_), .A2(new_n1394_), .B(new_n1398_), .ZN(new_n7147_));
  AOI21_X1   g6762(.A1(new_n7147_), .A2(new_n1722_), .B(new_n1723_), .ZN(new_n7148_));
  OAI21_X1   g6763(.A1(new_n7148_), .A2(new_n1234_), .B(new_n1407_), .ZN(new_n7149_));
  AOI21_X1   g6764(.A1(new_n7149_), .A2(new_n1720_), .B(new_n1721_), .ZN(new_n7150_));
  OAI21_X1   g6765(.A1(new_n7150_), .A2(new_n1230_), .B(new_n1419_), .ZN(new_n7151_));
  AOI21_X1   g6766(.A1(new_n7151_), .A2(new_n1718_), .B(new_n1719_), .ZN(new_n7152_));
  OAI21_X1   g6767(.A1(new_n7152_), .A2(new_n1428_), .B(new_n1432_), .ZN(new_n7153_));
  AOI21_X1   g6768(.A1(new_n7153_), .A2(new_n1716_), .B(new_n1717_), .ZN(new_n7154_));
  OAI21_X1   g6769(.A1(new_n7154_), .A2(new_n1220_), .B(new_n1441_), .ZN(new_n7155_));
  AOI21_X1   g6770(.A1(new_n7155_), .A2(new_n1714_), .B(new_n1715_), .ZN(new_n7156_));
  OAI21_X1   g6771(.A1(new_n7156_), .A2(new_n1216_), .B(new_n1453_), .ZN(new_n7157_));
  AOI21_X1   g6772(.A1(new_n7157_), .A2(new_n1712_), .B(new_n1713_), .ZN(new_n7158_));
  OAI21_X1   g6773(.A1(new_n7158_), .A2(new_n1462_), .B(new_n1466_), .ZN(new_n7159_));
  AOI21_X1   g6774(.A1(new_n7159_), .A2(new_n1710_), .B(new_n1711_), .ZN(new_n7160_));
  OAI21_X1   g6775(.A1(new_n7160_), .A2(new_n1206_), .B(new_n1475_), .ZN(new_n7161_));
  AOI21_X1   g6776(.A1(new_n7161_), .A2(new_n1708_), .B(new_n1709_), .ZN(new_n7162_));
  OAI21_X1   g6777(.A1(new_n7162_), .A2(new_n1202_), .B(new_n1487_), .ZN(new_n7163_));
  AOI21_X1   g6778(.A1(new_n7163_), .A2(new_n1706_), .B(new_n1707_), .ZN(new_n7164_));
  OAI21_X1   g6779(.A1(new_n7164_), .A2(new_n1496_), .B(new_n1500_), .ZN(new_n7165_));
  AOI21_X1   g6780(.A1(new_n7165_), .A2(new_n1704_), .B(new_n1705_), .ZN(new_n7166_));
  OAI21_X1   g6781(.A1(new_n7166_), .A2(new_n1192_), .B(new_n1509_), .ZN(new_n7167_));
  OAI21_X1   g6782(.A1(new_n800_), .A2(\priority[127] ), .B(\req[127] ), .ZN(new_n7168_));
  AOI21_X1   g6783(.A1(new_n7167_), .A2(new_n1702_), .B(new_n7168_), .ZN(\grant[127] ));
  NOR4_X1    g6784(.A1(new_n1162_), .A2(new_n1176_), .A3(new_n1284_), .A4(new_n1295_), .ZN(new_n7170_));
  NOR4_X1    g6785(.A1(new_n1304_), .A2(new_n1316_), .A3(new_n1329_), .A4(new_n1338_), .ZN(new_n7171_));
  NOR4_X1    g6786(.A1(new_n1107_), .A2(new_n1122_), .A3(new_n1136_), .A4(new_n1147_), .ZN(new_n7172_));
  NOR4_X1    g6787(.A1(new_n1056_), .A2(new_n1067_), .A3(new_n1082_), .A4(new_n1096_), .ZN(new_n7173_));
  AND4_X2    g6788(.A1(new_n7170_), .A2(new_n7171_), .A3(new_n7172_), .A4(new_n7173_), .Z(new_n7174_));
  NOR4_X1    g6789(.A1(new_n1440_), .A2(new_n1452_), .A3(new_n1465_), .A4(new_n1474_), .ZN(new_n7175_));
  NOR4_X1    g6790(.A1(new_n1486_), .A2(new_n1499_), .A3(new_n1508_), .A4(new_n1606_), .ZN(new_n7176_));
  NOR4_X1    g6791(.A1(new_n1397_), .A2(new_n1406_), .A3(new_n1418_), .A4(new_n1431_), .ZN(new_n7177_));
  NOR4_X1    g6792(.A1(new_n1350_), .A2(new_n1363_), .A3(new_n1372_), .A4(new_n1384_), .ZN(new_n7178_));
  AND4_X2    g6793(.A1(new_n7175_), .A2(new_n7176_), .A3(new_n7177_), .A4(new_n7178_), .Z(new_n7179_));
  NOR4_X1    g6794(.A1(new_n947_), .A2(new_n962_), .A3(new_n976_), .A4(new_n987_), .ZN(new_n7180_));
  NOR4_X1    g6795(.A1(new_n1002_), .A2(new_n1016_), .A3(new_n1027_), .A4(new_n1042_), .ZN(new_n7181_));
  NOR4_X1    g6796(.A1(new_n786_), .A2(new_n907_), .A3(new_n922_), .A4(new_n936_), .ZN(new_n7182_));
  NOR4_X1    g6797(.A1(new_n733_), .A2(new_n744_), .A3(new_n759_), .A4(new_n775_), .ZN(new_n7183_));
  AND4_X2    g6798(.A1(new_n7180_), .A2(new_n7181_), .A3(new_n7182_), .A4(new_n7183_), .Z(new_n7184_));
  NOR4_X1    g6799(.A1(new_n618_), .A2(new_n633_), .A3(new_n649_), .A4(new_n660_), .ZN(new_n7185_));
  NOR4_X1    g6800(.A1(new_n675_), .A2(new_n691_), .A3(new_n702_), .A4(new_n717_), .ZN(new_n7186_));
  NOR4_X1    g6801(.A1(new_n565_), .A2(new_n576_), .A3(new_n591_), .A4(new_n607_), .ZN(new_n7187_));
  NOR4_X1    g6802(.A1(new_n509_), .A2(new_n523_), .A3(new_n534_), .A4(new_n549_), .ZN(new_n7188_));
  AND4_X2    g6803(.A1(new_n7185_), .A2(new_n7186_), .A3(new_n7187_), .A4(new_n7188_), .Z(new_n7189_));
  NAND4_X1   g6804(.A1(new_n7174_), .A2(new_n7179_), .A3(new_n7184_), .A4(new_n7189_), .ZN(anyGrant));
endmodule


