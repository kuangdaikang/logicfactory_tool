// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:58 2022

module ex4  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43,
    v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57,
    v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71,
    v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85,
    v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99,
    v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111,
    v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123,
    v124, v125, v126, v127,
    \v128.0 , \v128.1 , \v128.2 , \v128.3 , \v128.4 , \v128.5 , \v128.6 ,
    \v128.7 , \v128.8 , \v128.9 , \v128.10 , \v128.11 , \v128.12 ,
    \v128.13 , \v128.14 , \v128.15 , \v128.16 , \v128.17 , \v128.18 ,
    \v128.19 , \v128.20 , \v128.21 , \v128.22 , \v128.23 , \v128.24 ,
    \v128.25 , \v128.26 , \v128.27   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42,
    v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56,
    v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70,
    v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84,
    v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98,
    v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110,
    v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122,
    v123, v124, v125, v126, v127;
  output \v128.0 , \v128.1 , \v128.2 , \v128.3 , \v128.4 , \v128.5 , \v128.6 ,
    \v128.7 , \v128.8 , \v128.9 , \v128.10 , \v128.11 , \v128.12 ,
    \v128.13 , \v128.14 , \v128.15 , \v128.16 , \v128.17 , \v128.18 ,
    \v128.19 , \v128.20 , \v128.21 , \v128.22 , \v128.23 , \v128.24 ,
    \v128.25 , \v128.26 , \v128.27 ;
  wire new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_;
  assign new_n158_ = ~v32 & ~v72;
  assign new_n159_ = ~v8 & ~v48;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~v80 & new_n160_;
  assign new_n162_ = ~v0 & new_n161_;
  assign new_n163_ = ~v48 & ~v72;
  assign new_n164_ = ~v8 & ~v32;
  assign new_n165_ = ~new_n163_ & ~new_n164_;
  assign new_n166_ = ~v64 & new_n165_;
  assign new_n167_ = ~v16 & new_n166_;
  assign new_n168_ = ~v32 & ~v48;
  assign new_n169_ = ~v8 & ~v72;
  assign new_n170_ = ~new_n168_ & ~new_n169_;
  assign new_n171_ = ~new_n167_ & new_n170_;
  assign new_n172_ = ~new_n162_ & new_n171_;
  assign \v128.0  = v40 & ~new_n172_;
  assign new_n174_ = ~v33 & ~v73;
  assign new_n175_ = ~v9 & ~v49;
  assign new_n176_ = ~new_n174_ & ~new_n175_;
  assign new_n177_ = ~v81 & new_n176_;
  assign new_n178_ = ~v1 & new_n177_;
  assign new_n179_ = ~v49 & ~v73;
  assign new_n180_ = ~v9 & ~v33;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign new_n182_ = ~v65 & new_n181_;
  assign new_n183_ = ~v17 & new_n182_;
  assign new_n184_ = ~v33 & ~v49;
  assign new_n185_ = ~v9 & ~v73;
  assign new_n186_ = ~new_n184_ & ~new_n185_;
  assign new_n187_ = ~new_n183_ & new_n186_;
  assign new_n188_ = ~new_n178_ & new_n187_;
  assign \v128.1  = v41 & ~new_n188_;
  assign new_n190_ = ~v34 & ~v74;
  assign new_n191_ = ~v10 & ~v50;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = ~v82 & new_n192_;
  assign new_n194_ = ~v2 & new_n193_;
  assign new_n195_ = ~v50 & ~v74;
  assign new_n196_ = ~v10 & ~v34;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = ~v66 & new_n197_;
  assign new_n199_ = ~v18 & new_n198_;
  assign new_n200_ = ~v34 & ~v50;
  assign new_n201_ = ~v10 & ~v74;
  assign new_n202_ = ~new_n200_ & ~new_n201_;
  assign new_n203_ = ~new_n199_ & new_n202_;
  assign new_n204_ = ~new_n194_ & new_n203_;
  assign \v128.2  = v42 & ~new_n204_;
  assign new_n206_ = ~v35 & ~v75;
  assign new_n207_ = ~v11 & ~v51;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = ~v83 & new_n208_;
  assign new_n210_ = ~v3 & new_n209_;
  assign new_n211_ = ~v51 & ~v75;
  assign new_n212_ = ~v11 & ~v35;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~v67 & new_n213_;
  assign new_n215_ = ~v19 & new_n214_;
  assign new_n216_ = ~v35 & ~v51;
  assign new_n217_ = ~v11 & ~v75;
  assign new_n218_ = ~new_n216_ & ~new_n217_;
  assign new_n219_ = ~new_n215_ & new_n218_;
  assign new_n220_ = ~new_n210_ & new_n219_;
  assign \v128.3  = v43 & ~new_n220_;
  assign new_n222_ = ~v36 & ~v76;
  assign new_n223_ = ~v12 & ~v52;
  assign new_n224_ = ~new_n222_ & ~new_n223_;
  assign new_n225_ = ~v84 & new_n224_;
  assign new_n226_ = ~v4 & new_n225_;
  assign new_n227_ = ~v52 & ~v76;
  assign new_n228_ = ~v12 & ~v36;
  assign new_n229_ = ~new_n227_ & ~new_n228_;
  assign new_n230_ = ~v68 & new_n229_;
  assign new_n231_ = ~v20 & new_n230_;
  assign new_n232_ = ~v36 & ~v52;
  assign new_n233_ = ~v12 & ~v76;
  assign new_n234_ = ~new_n232_ & ~new_n233_;
  assign new_n235_ = ~new_n231_ & new_n234_;
  assign new_n236_ = ~new_n226_ & new_n235_;
  assign \v128.4  = v44 & ~new_n236_;
  assign new_n238_ = v109 & v117;
  assign new_n239_ = ~v37 & ~v69;
  assign new_n240_ = ~v13 & ~v21;
  assign new_n241_ = ~v61 & ~v93;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = ~new_n239_ & ~new_n242_;
  assign new_n244_ = ~v5 & new_n243_;
  assign new_n245_ = ~new_n240_ & ~new_n241_;
  assign new_n246_ = ~v29 & new_n245_;
  assign new_n247_ = v13 & v21;
  assign new_n248_ = ~new_n246_ & new_n247_;
  assign new_n249_ = ~new_n244_ & new_n248_;
  assign new_n250_ = ~new_n238_ & ~new_n249_;
  assign new_n251_ = v101 & v125;
  assign new_n252_ = ~v5 & ~new_n239_;
  assign new_n253_ = ~v29 & ~new_n240_;
  assign new_n254_ = ~new_n252_ & ~new_n253_;
  assign new_n255_ = ~new_n251_ & ~new_n254_;
  assign new_n256_ = v37 & v69;
  assign new_n257_ = v5 & new_n256_;
  assign new_n258_ = ~new_n240_ & ~new_n257_;
  assign new_n259_ = ~v29 & new_n258_;
  assign new_n260_ = ~new_n255_ & ~new_n259_;
  assign new_n261_ = ~new_n241_ & ~new_n260_;
  assign new_n262_ = v61 & v93;
  assign new_n263_ = ~v109 & ~v117;
  assign new_n264_ = new_n239_ & new_n263_;
  assign new_n265_ = ~new_n240_ & ~new_n264_;
  assign new_n266_ = ~v5 & new_n265_;
  assign new_n267_ = new_n256_ & ~new_n266_;
  assign new_n268_ = ~new_n262_ & ~new_n267_;
  assign new_n269_ = v29 & new_n251_;
  assign new_n270_ = ~new_n240_ & ~new_n269_;
  assign new_n271_ = ~new_n239_ & new_n270_;
  assign new_n272_ = v29 & v125;
  assign new_n273_ = ~new_n240_ & ~new_n272_;
  assign new_n274_ = ~new_n263_ & new_n273_;
  assign new_n275_ = ~new_n271_ & ~new_n274_;
  assign new_n276_ = ~v5 & ~new_n275_;
  assign new_n277_ = ~new_n268_ & ~new_n276_;
  assign new_n278_ = ~new_n261_ & new_n277_;
  assign new_n279_ = ~new_n250_ & new_n278_;
  assign new_n280_ = v85 & ~new_n279_;
  assign new_n281_ = ~v5 & ~v85;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = v77 & ~new_n282_;
  assign new_n284_ = ~v13 & ~v37;
  assign new_n285_ = ~v69 & ~new_n284_;
  assign new_n286_ = ~v21 & new_n285_;
  assign new_n287_ = v37 & ~v85;
  assign new_n288_ = ~v5 & new_n287_;
  assign new_n289_ = ~new_n286_ & ~new_n288_;
  assign new_n290_ = ~new_n283_ & new_n289_;
  assign new_n291_ = v53 & ~new_n290_;
  assign new_n292_ = ~v37 & ~v77;
  assign new_n293_ = ~v85 & ~new_n292_;
  assign new_n294_ = ~v5 & new_n293_;
  assign new_n295_ = ~v69 & v77;
  assign new_n296_ = ~v21 & new_n295_;
  assign new_n297_ = ~new_n294_ & ~new_n296_;
  assign new_n298_ = v13 & ~new_n297_;
  assign new_n299_ = ~v37 & ~v53;
  assign new_n300_ = ~v21 & v37;
  assign new_n301_ = new_n295_ & new_n300_;
  assign new_n302_ = ~v13 & ~v77;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = ~new_n299_ & new_n303_;
  assign new_n305_ = ~new_n298_ & new_n304_;
  assign new_n306_ = ~new_n291_ & new_n305_;
  assign \v128.5  = v45 & ~new_n306_;
  assign new_n308_ = v110 & v118;
  assign new_n309_ = ~v38 & ~v70;
  assign new_n310_ = ~v14 & ~v22;
  assign new_n311_ = ~v62 & ~v94;
  assign new_n312_ = new_n310_ & new_n311_;
  assign new_n313_ = ~new_n309_ & ~new_n312_;
  assign new_n314_ = ~v6 & new_n313_;
  assign new_n315_ = ~new_n310_ & ~new_n311_;
  assign new_n316_ = ~v30 & new_n315_;
  assign new_n317_ = v14 & v22;
  assign new_n318_ = ~new_n316_ & new_n317_;
  assign new_n319_ = ~new_n314_ & new_n318_;
  assign new_n320_ = ~new_n308_ & ~new_n319_;
  assign new_n321_ = v102 & v126;
  assign new_n322_ = ~v6 & ~new_n309_;
  assign new_n323_ = ~v30 & ~new_n310_;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign new_n325_ = ~new_n321_ & ~new_n324_;
  assign new_n326_ = v38 & v70;
  assign new_n327_ = v6 & new_n326_;
  assign new_n328_ = ~new_n310_ & ~new_n327_;
  assign new_n329_ = ~v30 & new_n328_;
  assign new_n330_ = ~new_n325_ & ~new_n329_;
  assign new_n331_ = ~new_n311_ & ~new_n330_;
  assign new_n332_ = v62 & v94;
  assign new_n333_ = ~v110 & ~v118;
  assign new_n334_ = new_n309_ & new_n333_;
  assign new_n335_ = ~new_n310_ & ~new_n334_;
  assign new_n336_ = ~v6 & new_n335_;
  assign new_n337_ = new_n326_ & ~new_n336_;
  assign new_n338_ = ~new_n332_ & ~new_n337_;
  assign new_n339_ = v30 & new_n321_;
  assign new_n340_ = ~new_n310_ & ~new_n339_;
  assign new_n341_ = ~new_n309_ & new_n340_;
  assign new_n342_ = v30 & v126;
  assign new_n343_ = ~new_n310_ & ~new_n342_;
  assign new_n344_ = ~new_n333_ & new_n343_;
  assign new_n345_ = ~new_n341_ & ~new_n344_;
  assign new_n346_ = ~v6 & ~new_n345_;
  assign new_n347_ = ~new_n338_ & ~new_n346_;
  assign new_n348_ = ~new_n331_ & new_n347_;
  assign new_n349_ = ~new_n320_ & new_n348_;
  assign new_n350_ = v86 & ~new_n349_;
  assign new_n351_ = ~v6 & ~v86;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = v78 & ~new_n352_;
  assign new_n354_ = ~v14 & ~v38;
  assign new_n355_ = ~v70 & ~new_n354_;
  assign new_n356_ = ~v22 & new_n355_;
  assign new_n357_ = v38 & ~v86;
  assign new_n358_ = ~v6 & new_n357_;
  assign new_n359_ = ~new_n356_ & ~new_n358_;
  assign new_n360_ = ~new_n353_ & new_n359_;
  assign new_n361_ = v54 & ~new_n360_;
  assign new_n362_ = ~v38 & ~v78;
  assign new_n363_ = ~v86 & ~new_n362_;
  assign new_n364_ = ~v6 & new_n363_;
  assign new_n365_ = ~v70 & v78;
  assign new_n366_ = ~v22 & new_n365_;
  assign new_n367_ = ~new_n364_ & ~new_n366_;
  assign new_n368_ = v14 & ~new_n367_;
  assign new_n369_ = ~v38 & ~v54;
  assign new_n370_ = ~v22 & v38;
  assign new_n371_ = new_n365_ & new_n370_;
  assign new_n372_ = ~v14 & ~v78;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = ~new_n369_ & new_n373_;
  assign new_n375_ = ~new_n368_ & new_n374_;
  assign new_n376_ = ~new_n361_ & new_n375_;
  assign \v128.6  = v46 & ~new_n376_;
  assign new_n378_ = ~v104 & ~v112;
  assign new_n379_ = v32 & v64;
  assign new_n380_ = v8 & v16;
  assign new_n381_ = v56 & v88;
  assign new_n382_ = new_n380_ & new_n381_;
  assign new_n383_ = ~new_n379_ & ~new_n382_;
  assign new_n384_ = v0 & new_n383_;
  assign new_n385_ = ~v8 & ~v16;
  assign new_n386_ = ~new_n380_ & ~new_n381_;
  assign new_n387_ = v24 & new_n386_;
  assign new_n388_ = new_n385_ & ~new_n387_;
  assign new_n389_ = ~new_n384_ & new_n388_;
  assign new_n390_ = ~new_n378_ & ~new_n389_;
  assign new_n391_ = ~v0 & ~v32;
  assign new_n392_ = ~v96 & ~v120;
  assign new_n393_ = ~v64 & new_n392_;
  assign new_n394_ = new_n391_ & new_n393_;
  assign new_n395_ = ~new_n380_ & ~new_n394_;
  assign new_n396_ = v24 & new_n395_;
  assign new_n397_ = ~new_n379_ & ~new_n392_;
  assign new_n398_ = v0 & new_n397_;
  assign new_n399_ = ~new_n396_ & ~new_n398_;
  assign new_n400_ = ~new_n381_ & ~new_n399_;
  assign new_n401_ = ~v56 & ~v88;
  assign new_n402_ = ~v32 & ~v64;
  assign new_n403_ = v104 & v112;
  assign new_n404_ = new_n379_ & new_n403_;
  assign new_n405_ = ~new_n380_ & ~new_n404_;
  assign new_n406_ = v0 & new_n405_;
  assign new_n407_ = new_n402_ & ~new_n406_;
  assign new_n408_ = ~new_n401_ & ~new_n407_;
  assign new_n409_ = ~v24 & new_n392_;
  assign new_n410_ = ~new_n380_ & ~new_n409_;
  assign new_n411_ = ~new_n379_ & new_n410_;
  assign new_n412_ = ~v24 & ~v120;
  assign new_n413_ = ~new_n380_ & ~new_n412_;
  assign new_n414_ = ~new_n403_ & new_n413_;
  assign new_n415_ = ~new_n411_ & ~new_n414_;
  assign new_n416_ = v0 & ~new_n415_;
  assign new_n417_ = ~new_n408_ & ~new_n416_;
  assign new_n418_ = ~new_n400_ & new_n417_;
  assign new_n419_ = ~new_n390_ & new_n418_;
  assign new_n420_ = ~v80 & ~new_n419_;
  assign new_n421_ = v0 & v80;
  assign new_n422_ = ~new_n420_ & ~new_n421_;
  assign new_n423_ = ~v72 & ~new_n422_;
  assign new_n424_ = v8 & v32;
  assign new_n425_ = v64 & ~new_n424_;
  assign new_n426_ = v16 & new_n425_;
  assign new_n427_ = ~v32 & v80;
  assign new_n428_ = v0 & new_n427_;
  assign new_n429_ = ~new_n426_ & ~new_n428_;
  assign new_n430_ = ~new_n423_ & new_n429_;
  assign new_n431_ = ~v48 & ~new_n430_;
  assign new_n432_ = v32 & v72;
  assign new_n433_ = v80 & ~new_n432_;
  assign new_n434_ = v0 & new_n433_;
  assign new_n435_ = v64 & ~v72;
  assign new_n436_ = v16 & new_n435_;
  assign new_n437_ = ~new_n434_ & ~new_n436_;
  assign new_n438_ = ~v8 & ~new_n437_;
  assign new_n439_ = v32 & v48;
  assign new_n440_ = v16 & ~v32;
  assign new_n441_ = new_n435_ & new_n440_;
  assign new_n442_ = v8 & v72;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign new_n444_ = ~new_n439_ & new_n443_;
  assign new_n445_ = ~new_n438_ & new_n444_;
  assign new_n446_ = ~new_n431_ & new_n445_;
  assign \v128.8  = ~v40 & ~new_n446_;
  assign new_n448_ = v33 & v73;
  assign new_n449_ = v9 & v49;
  assign new_n450_ = ~new_n448_ & ~new_n449_;
  assign new_n451_ = v81 & new_n450_;
  assign new_n452_ = v1 & new_n451_;
  assign new_n453_ = v49 & v73;
  assign new_n454_ = v9 & v33;
  assign new_n455_ = ~new_n453_ & ~new_n454_;
  assign new_n456_ = v65 & new_n455_;
  assign new_n457_ = v17 & new_n456_;
  assign new_n458_ = v33 & v49;
  assign new_n459_ = v9 & v73;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~new_n457_ & new_n460_;
  assign new_n462_ = ~new_n452_ & new_n461_;
  assign \v128.9  = ~v41 & ~new_n462_;
  assign new_n464_ = v34 & v74;
  assign new_n465_ = v10 & v50;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign new_n467_ = v82 & new_n466_;
  assign new_n468_ = v2 & new_n467_;
  assign new_n469_ = v50 & v74;
  assign new_n470_ = v10 & v34;
  assign new_n471_ = ~new_n469_ & ~new_n470_;
  assign new_n472_ = v66 & new_n471_;
  assign new_n473_ = v18 & new_n472_;
  assign new_n474_ = v34 & v50;
  assign new_n475_ = v10 & v74;
  assign new_n476_ = ~new_n474_ & ~new_n475_;
  assign new_n477_ = ~new_n473_ & new_n476_;
  assign new_n478_ = ~new_n468_ & new_n477_;
  assign \v128.10  = ~v42 & ~new_n478_;
  assign new_n480_ = v35 & v75;
  assign new_n481_ = v11 & v51;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = v83 & new_n482_;
  assign new_n484_ = v3 & new_n483_;
  assign new_n485_ = v51 & v75;
  assign new_n486_ = v11 & v35;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = v67 & new_n487_;
  assign new_n489_ = v19 & new_n488_;
  assign new_n490_ = v35 & v51;
  assign new_n491_ = v11 & v75;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = ~new_n489_ & new_n492_;
  assign new_n494_ = ~new_n484_ & new_n493_;
  assign \v128.11  = ~v43 & ~new_n494_;
  assign new_n496_ = v36 & v76;
  assign new_n497_ = v12 & v52;
  assign new_n498_ = ~new_n496_ & ~new_n497_;
  assign new_n499_ = v84 & new_n498_;
  assign new_n500_ = v4 & new_n499_;
  assign new_n501_ = v52 & v76;
  assign new_n502_ = v12 & v36;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign new_n504_ = v68 & new_n503_;
  assign new_n505_ = v20 & new_n504_;
  assign new_n506_ = v36 & v52;
  assign new_n507_ = v12 & v76;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = ~new_n505_ & new_n508_;
  assign new_n510_ = ~new_n500_ & new_n509_;
  assign \v128.12  = ~v44 & ~new_n510_;
  assign new_n512_ = new_n247_ & new_n262_;
  assign new_n513_ = ~new_n256_ & ~new_n512_;
  assign new_n514_ = v5 & new_n513_;
  assign new_n515_ = ~new_n247_ & ~new_n262_;
  assign new_n516_ = v29 & new_n515_;
  assign new_n517_ = new_n240_ & ~new_n516_;
  assign new_n518_ = ~new_n514_ & new_n517_;
  assign new_n519_ = ~new_n263_ & ~new_n518_;
  assign new_n520_ = ~v5 & ~v37;
  assign new_n521_ = ~v101 & ~v125;
  assign new_n522_ = ~v69 & new_n521_;
  assign new_n523_ = new_n520_ & new_n522_;
  assign new_n524_ = ~new_n247_ & ~new_n523_;
  assign new_n525_ = v29 & new_n524_;
  assign new_n526_ = ~new_n256_ & ~new_n521_;
  assign new_n527_ = v5 & new_n526_;
  assign new_n528_ = ~new_n525_ & ~new_n527_;
  assign new_n529_ = ~new_n262_ & ~new_n528_;
  assign new_n530_ = new_n238_ & new_n256_;
  assign new_n531_ = ~new_n247_ & ~new_n530_;
  assign new_n532_ = v5 & new_n531_;
  assign new_n533_ = new_n239_ & ~new_n532_;
  assign new_n534_ = ~new_n241_ & ~new_n533_;
  assign new_n535_ = ~v29 & new_n521_;
  assign new_n536_ = ~new_n247_ & ~new_n535_;
  assign new_n537_ = ~new_n256_ & new_n536_;
  assign new_n538_ = ~v29 & ~v125;
  assign new_n539_ = ~new_n247_ & ~new_n538_;
  assign new_n540_ = ~new_n238_ & new_n539_;
  assign new_n541_ = ~new_n537_ & ~new_n540_;
  assign new_n542_ = v5 & ~new_n541_;
  assign new_n543_ = ~new_n534_ & ~new_n542_;
  assign new_n544_ = ~new_n529_ & new_n543_;
  assign new_n545_ = ~new_n519_ & new_n544_;
  assign new_n546_ = ~v85 & ~new_n545_;
  assign new_n547_ = v5 & v85;
  assign new_n548_ = ~new_n546_ & ~new_n547_;
  assign new_n549_ = ~v77 & ~new_n548_;
  assign new_n550_ = v13 & v37;
  assign new_n551_ = v69 & ~new_n550_;
  assign new_n552_ = v21 & new_n551_;
  assign new_n553_ = ~v37 & v85;
  assign new_n554_ = v5 & new_n553_;
  assign new_n555_ = ~new_n552_ & ~new_n554_;
  assign new_n556_ = ~new_n549_ & new_n555_;
  assign new_n557_ = ~v53 & ~new_n556_;
  assign new_n558_ = v37 & v77;
  assign new_n559_ = v85 & ~new_n558_;
  assign new_n560_ = v5 & new_n559_;
  assign new_n561_ = v69 & ~v77;
  assign new_n562_ = v21 & new_n561_;
  assign new_n563_ = ~new_n560_ & ~new_n562_;
  assign new_n564_ = ~v13 & ~new_n563_;
  assign new_n565_ = v37 & v53;
  assign new_n566_ = v21 & ~v37;
  assign new_n567_ = new_n561_ & new_n566_;
  assign new_n568_ = v13 & v77;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = ~new_n565_ & new_n569_;
  assign new_n571_ = ~new_n564_ & new_n570_;
  assign new_n572_ = ~new_n557_ & new_n571_;
  assign \v128.13  = ~v45 & ~new_n572_;
  assign new_n574_ = new_n317_ & new_n332_;
  assign new_n575_ = ~new_n326_ & ~new_n574_;
  assign new_n576_ = v6 & new_n575_;
  assign new_n577_ = ~new_n317_ & ~new_n332_;
  assign new_n578_ = v30 & new_n577_;
  assign new_n579_ = new_n310_ & ~new_n578_;
  assign new_n580_ = ~new_n576_ & new_n579_;
  assign new_n581_ = ~new_n333_ & ~new_n580_;
  assign new_n582_ = ~v6 & ~v38;
  assign new_n583_ = ~v102 & ~v126;
  assign new_n584_ = ~v70 & new_n583_;
  assign new_n585_ = new_n582_ & new_n584_;
  assign new_n586_ = ~new_n317_ & ~new_n585_;
  assign new_n587_ = v30 & new_n586_;
  assign new_n588_ = ~new_n326_ & ~new_n583_;
  assign new_n589_ = v6 & new_n588_;
  assign new_n590_ = ~new_n587_ & ~new_n589_;
  assign new_n591_ = ~new_n332_ & ~new_n590_;
  assign new_n592_ = new_n308_ & new_n326_;
  assign new_n593_ = ~new_n317_ & ~new_n592_;
  assign new_n594_ = v6 & new_n593_;
  assign new_n595_ = new_n309_ & ~new_n594_;
  assign new_n596_ = ~new_n311_ & ~new_n595_;
  assign new_n597_ = ~v30 & new_n583_;
  assign new_n598_ = ~new_n317_ & ~new_n597_;
  assign new_n599_ = ~new_n326_ & new_n598_;
  assign new_n600_ = ~v30 & ~v126;
  assign new_n601_ = ~new_n317_ & ~new_n600_;
  assign new_n602_ = ~new_n308_ & new_n601_;
  assign new_n603_ = ~new_n599_ & ~new_n602_;
  assign new_n604_ = v6 & ~new_n603_;
  assign new_n605_ = ~new_n596_ & ~new_n604_;
  assign new_n606_ = ~new_n591_ & new_n605_;
  assign new_n607_ = ~new_n581_ & new_n606_;
  assign new_n608_ = ~v86 & ~new_n607_;
  assign new_n609_ = v6 & v86;
  assign new_n610_ = ~new_n608_ & ~new_n609_;
  assign new_n611_ = ~v78 & ~new_n610_;
  assign new_n612_ = v14 & v38;
  assign new_n613_ = v70 & ~new_n612_;
  assign new_n614_ = v22 & new_n613_;
  assign new_n615_ = ~v38 & v86;
  assign new_n616_ = v6 & new_n615_;
  assign new_n617_ = ~new_n614_ & ~new_n616_;
  assign new_n618_ = ~new_n611_ & new_n617_;
  assign new_n619_ = ~v54 & ~new_n618_;
  assign new_n620_ = v38 & v78;
  assign new_n621_ = v86 & ~new_n620_;
  assign new_n622_ = v6 & new_n621_;
  assign new_n623_ = v70 & ~v78;
  assign new_n624_ = v22 & new_n623_;
  assign new_n625_ = ~new_n622_ & ~new_n624_;
  assign new_n626_ = ~v14 & ~new_n625_;
  assign new_n627_ = v38 & v54;
  assign new_n628_ = v22 & ~v38;
  assign new_n629_ = new_n623_ & new_n628_;
  assign new_n630_ = v14 & v78;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = ~new_n627_ & new_n631_;
  assign new_n633_ = ~new_n626_ & new_n632_;
  assign new_n634_ = ~new_n619_ & new_n633_;
  assign \v128.14  = ~v46 & ~new_n634_;
  assign \v128.7  = 1'b0;
  assign \v128.15  = 1'b0;
  assign \v128.16  = 1'b0;
  assign \v128.17  = 1'b0;
  assign \v128.18  = 1'b0;
  assign \v128.19  = 1'b0;
  assign \v128.20  = 1'b0;
  assign \v128.21  = 1'b0;
  assign \v128.22  = 1'b0;
  assign \v128.23  = 1'b0;
  assign \v128.24  = 1'b0;
  assign \v128.25  = 1'b0;
  assign \v128.26  = 1'b0;
  assign \v128.27  = 1'b0;
endmodule


