// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:35 2022

module b4  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32,
    \v33.0 , \v33.1 , \v33.2 , \v33.3 , \v33.4 , \v33.5 , \v33.6 , \v33.7 ,
    \v33.8 , \v33.9 , \v33.10 , \v33.11 , \v33.12 , \v33.13 , \v33.14 ,
    \v33.15 , \v33.16 , \v33.17 , \v33.18 , \v33.19 , \v33.20 , \v33.21 ,
    \v33.22   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32;
  output \v33.0 , \v33.1 , \v33.2 , \v33.3 , \v33.4 , \v33.5 , \v33.6 ,
    \v33.7 , \v33.8 , \v33.9 , \v33.10 , \v33.11 , \v33.12 , \v33.13 ,
    \v33.14 , \v33.15 , \v33.16 , \v33.17 , \v33.18 , \v33.19 , \v33.20 ,
    \v33.21 , \v33.22 ;
  wire new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n73_,
    new_n74_, new_n76_, new_n77_, new_n78_, new_n79_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n112_, new_n113_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n339_, new_n340_, new_n342_,
    new_n343_, new_n344_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_;
  assign new_n58_ = ~v16 & v31;
  assign new_n59_ = ~v15 & new_n58_;
  assign new_n60_ = v1 & v22;
  assign new_n61_ = v30 & ~v31;
  assign new_n62_ = v28 & new_n61_;
  assign new_n63_ = new_n60_ & new_n62_;
  assign new_n64_ = ~new_n59_ & ~new_n63_;
  assign \v33.1  = ~v0 & ~new_n64_;
  assign new_n66_ = ~v4 & v32;
  assign new_n67_ = v1 & v24;
  assign new_n68_ = v29 & ~v32;
  assign new_n69_ = v28 & new_n68_;
  assign new_n70_ = new_n67_ & new_n69_;
  assign new_n71_ = ~new_n66_ & ~new_n70_;
  assign \v33.2  = ~v0 & ~new_n71_;
  assign new_n73_ = ~v28 & ~v30;
  assign new_n74_ = v3 & new_n73_;
  assign \v33.3  = ~v0 & new_n74_;
  assign new_n76_ = ~v0 & v3;
  assign new_n77_ = v29 & ~v30;
  assign new_n78_ = ~v28 & new_n77_;
  assign new_n79_ = new_n76_ & new_n78_;
  assign \v33.4  = v0 | new_n79_;
  assign new_n81_ = ~v11 & ~v12;
  assign new_n82_ = v11 & v12;
  assign new_n83_ = v21 & v29;
  assign new_n84_ = new_n82_ & new_n83_;
  assign new_n85_ = ~new_n81_ & ~new_n84_;
  assign new_n86_ = ~v9 & ~new_n85_;
  assign new_n87_ = v12 & v20;
  assign new_n88_ = ~v12 & v21;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = v29 & ~new_n89_;
  assign new_n91_ = v19 & new_n90_;
  assign new_n92_ = v11 & new_n91_;
  assign new_n93_ = ~v11 & v12;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = v9 & ~new_n94_;
  assign new_n96_ = ~new_n86_ & ~new_n95_;
  assign new_n97_ = v10 & ~new_n96_;
  assign new_n98_ = v10 & ~new_n81_;
  assign new_n99_ = v29 & ~new_n98_;
  assign new_n100_ = v21 & new_n99_;
  assign new_n101_ = v20 & new_n100_;
  assign new_n102_ = v19 & new_n101_;
  assign new_n103_ = v9 & new_n102_;
  assign new_n104_ = ~v9 & ~v10;
  assign new_n105_ = v11 & ~v12;
  assign new_n106_ = new_n104_ & new_n105_;
  assign new_n107_ = ~new_n103_ & ~new_n106_;
  assign new_n108_ = ~new_n97_ & new_n107_;
  assign new_n109_ = v30 & ~new_n108_;
  assign new_n110_ = ~v28 & new_n109_;
  assign \v33.5  = ~v0 & new_n110_;
  assign new_n112_ = ~v15 & v17;
  assign new_n113_ = v15 & ~v17;
  assign new_n114_ = v7 & new_n113_;
  assign new_n115_ = ~new_n112_ & ~new_n114_;
  assign new_n116_ = ~v6 & ~new_n115_;
  assign new_n117_ = v15 & v17;
  assign new_n118_ = ~v14 & new_n117_;
  assign new_n119_ = ~new_n116_ & ~new_n118_;
  assign new_n120_ = v28 & ~new_n119_;
  assign new_n121_ = v23 & new_n120_;
  assign new_n122_ = v1 & new_n121_;
  assign new_n123_ = ~v9 & v10;
  assign new_n124_ = new_n81_ & new_n123_;
  assign new_n125_ = ~v14 & v15;
  assign new_n126_ = v17 & ~v28;
  assign new_n127_ = new_n125_ & new_n126_;
  assign new_n128_ = new_n124_ & new_n127_;
  assign new_n129_ = ~new_n122_ & ~new_n128_;
  assign new_n130_ = v30 & ~new_n129_;
  assign new_n131_ = ~v18 & new_n130_;
  assign new_n132_ = ~v16 & new_n131_;
  assign \v33.6  = ~v0 & new_n132_;
  assign new_n134_ = ~v17 & v18;
  assign new_n135_ = v16 & new_n134_;
  assign new_n136_ = ~v6 & ~v16;
  assign new_n137_ = v17 & ~v18;
  assign new_n138_ = new_n136_ & new_n137_;
  assign new_n139_ = ~new_n135_ & ~new_n138_;
  assign new_n140_ = v23 & v28;
  assign new_n141_ = v1 & new_n140_;
  assign new_n142_ = ~v12 & ~v28;
  assign new_n143_ = ~v11 & new_n142_;
  assign new_n144_ = new_n123_ & new_n143_;
  assign new_n145_ = ~new_n141_ & ~new_n144_;
  assign new_n146_ = ~new_n139_ & ~new_n145_;
  assign new_n147_ = ~v8 & v18;
  assign new_n148_ = ~v6 & new_n147_;
  assign new_n149_ = ~v6 & ~new_n148_;
  assign new_n150_ = v17 & ~new_n149_;
  assign new_n151_ = ~v17 & ~v18;
  assign new_n152_ = ~new_n150_ & ~new_n151_;
  assign new_n153_ = ~v28 & ~new_n152_;
  assign new_n154_ = v23 & new_n153_;
  assign new_n155_ = ~v16 & new_n154_;
  assign new_n156_ = v12 & new_n155_;
  assign new_n157_ = v11 & new_n156_;
  assign new_n158_ = ~v10 & new_n157_;
  assign new_n159_ = ~v9 & new_n158_;
  assign new_n160_ = v1 & new_n159_;
  assign new_n161_ = ~new_n146_ & ~new_n160_;
  assign new_n162_ = v30 & ~new_n161_;
  assign new_n163_ = ~v15 & new_n162_;
  assign \v33.7  = ~v0 & new_n163_;
  assign new_n165_ = v22 & v28;
  assign new_n166_ = v1 & new_n165_;
  assign new_n167_ = ~new_n144_ & ~new_n166_;
  assign new_n168_ = v18 & ~new_n167_;
  assign new_n169_ = ~v15 & new_n168_;
  assign new_n170_ = ~v0 & new_n169_;
  assign new_n171_ = new_n82_ & new_n104_;
  assign new_n172_ = ~v28 & ~new_n171_;
  assign new_n173_ = v22 & ~new_n172_;
  assign new_n174_ = ~v18 & new_n173_;
  assign new_n175_ = v15 & new_n174_;
  assign new_n176_ = v1 & new_n175_;
  assign new_n177_ = ~new_n170_ & ~new_n176_;
  assign new_n178_ = v30 & ~new_n177_;
  assign new_n179_ = ~v17 & new_n178_;
  assign new_n180_ = v16 & new_n179_;
  assign \v33.8  = v0 | new_n180_;
  assign new_n182_ = v10 & new_n81_;
  assign new_n183_ = ~v16 & v17;
  assign new_n184_ = ~v14 & new_n183_;
  assign new_n185_ = new_n182_ & new_n184_;
  assign new_n186_ = v1 & ~v6;
  assign new_n187_ = v8 & ~v10;
  assign new_n188_ = new_n186_ & new_n187_;
  assign new_n189_ = ~v17 & v22;
  assign new_n190_ = v16 & new_n189_;
  assign new_n191_ = new_n82_ & new_n190_;
  assign new_n192_ = new_n188_ & new_n191_;
  assign new_n193_ = ~new_n185_ & ~new_n192_;
  assign new_n194_ = ~v0 & ~new_n193_;
  assign new_n195_ = v7 & v10;
  assign new_n196_ = ~v6 & new_n195_;
  assign new_n197_ = ~v16 & ~v17;
  assign new_n198_ = new_n81_ & new_n197_;
  assign new_n199_ = new_n196_ & new_n198_;
  assign new_n200_ = ~new_n194_ & ~new_n199_;
  assign new_n201_ = ~v28 & ~new_n200_;
  assign new_n202_ = ~v9 & new_n201_;
  assign new_n203_ = v16 & ~v17;
  assign new_n204_ = v16 & ~new_n203_;
  assign new_n205_ = v28 & ~new_n204_;
  assign new_n206_ = v22 & new_n205_;
  assign new_n207_ = v1 & new_n206_;
  assign new_n208_ = ~new_n202_ & ~new_n207_;
  assign new_n209_ = v30 & ~new_n208_;
  assign new_n210_ = ~v18 & new_n209_;
  assign new_n211_ = v15 & new_n210_;
  assign \v33.9  = v0 | new_n211_;
  assign new_n213_ = ~v6 & ~v15;
  assign new_n214_ = ~new_n125_ & ~new_n213_;
  assign new_n215_ = v17 & ~new_n214_;
  assign new_n216_ = ~v0 & new_n215_;
  assign new_n217_ = ~v6 & v7;
  assign new_n218_ = new_n113_ & new_n217_;
  assign new_n219_ = ~new_n216_ & ~new_n218_;
  assign new_n220_ = v28 & ~new_n219_;
  assign new_n221_ = v22 & new_n220_;
  assign new_n222_ = v1 & new_n221_;
  assign new_n223_ = v10 & ~v11;
  assign new_n224_ = ~v0 & ~v9;
  assign new_n225_ = new_n223_ & new_n224_;
  assign new_n226_ = ~v12 & ~v14;
  assign new_n227_ = v15 & new_n126_;
  assign new_n228_ = new_n226_ & new_n227_;
  assign new_n229_ = new_n225_ & new_n228_;
  assign new_n230_ = ~new_n222_ & ~new_n229_;
  assign new_n231_ = v30 & ~new_n230_;
  assign new_n232_ = ~v18 & new_n231_;
  assign new_n233_ = ~v16 & new_n232_;
  assign new_n234_ = v0 & v7;
  assign \v33.10  = new_n233_ | new_n234_;
  assign new_n236_ = ~v15 & v16;
  assign new_n237_ = v6 & ~new_n236_;
  assign new_n238_ = ~v6 & v8;
  assign new_n239_ = v15 & v16;
  assign new_n240_ = new_n238_ & new_n239_;
  assign new_n241_ = ~new_n237_ & ~new_n240_;
  assign new_n242_ = ~v0 & ~new_n241_;
  assign new_n243_ = ~v15 & ~v16;
  assign new_n244_ = v7 & new_n243_;
  assign new_n245_ = ~new_n242_ & ~new_n244_;
  assign new_n246_ = ~v28 & ~new_n245_;
  assign new_n247_ = v12 & new_n246_;
  assign new_n248_ = v11 & new_n247_;
  assign new_n249_ = ~v10 & new_n248_;
  assign new_n250_ = ~v9 & new_n249_;
  assign new_n251_ = ~v16 & v28;
  assign new_n252_ = v15 & new_n251_;
  assign new_n253_ = new_n217_ & new_n252_;
  assign new_n254_ = ~new_n250_ & ~new_n253_;
  assign new_n255_ = ~v18 & ~new_n254_;
  assign new_n256_ = ~v0 & ~v15;
  assign new_n257_ = v18 & v28;
  assign new_n258_ = v16 & new_n257_;
  assign new_n259_ = new_n256_ & new_n258_;
  assign new_n260_ = ~new_n255_ & ~new_n259_;
  assign new_n261_ = v22 & ~new_n260_;
  assign new_n262_ = v1 & new_n261_;
  assign new_n263_ = v16 & v18;
  assign new_n264_ = new_n256_ & new_n263_;
  assign new_n265_ = ~v16 & ~v18;
  assign new_n266_ = v15 & new_n265_;
  assign new_n267_ = new_n217_ & new_n266_;
  assign new_n268_ = ~new_n264_ & ~new_n267_;
  assign new_n269_ = ~v28 & ~new_n268_;
  assign new_n270_ = ~v12 & new_n269_;
  assign new_n271_ = ~v11 & new_n270_;
  assign new_n272_ = v10 & new_n271_;
  assign new_n273_ = ~v9 & new_n272_;
  assign new_n274_ = ~new_n262_ & ~new_n273_;
  assign new_n275_ = v30 & ~new_n274_;
  assign new_n276_ = ~v17 & new_n275_;
  assign \v33.11  = new_n234_ | new_n276_;
  assign new_n278_ = ~v10 & v11;
  assign new_n279_ = v1 & new_n278_;
  assign new_n280_ = v17 & v23;
  assign new_n281_ = v12 & ~v16;
  assign new_n282_ = new_n280_ & new_n281_;
  assign new_n283_ = new_n279_ & new_n282_;
  assign new_n284_ = ~v17 & ~v28;
  assign new_n285_ = v16 & new_n284_;
  assign new_n286_ = new_n182_ & new_n285_;
  assign new_n287_ = ~new_n283_ & ~new_n286_;
  assign new_n288_ = ~v9 & ~new_n287_;
  assign new_n289_ = ~new_n183_ & ~new_n203_;
  assign new_n290_ = v28 & ~new_n289_;
  assign new_n291_ = v23 & new_n290_;
  assign new_n292_ = v1 & new_n291_;
  assign new_n293_ = ~new_n288_ & ~new_n292_;
  assign new_n294_ = v30 & ~new_n293_;
  assign new_n295_ = v18 & new_n294_;
  assign new_n296_ = ~v15 & new_n295_;
  assign new_n297_ = ~v0 & new_n296_;
  assign new_n298_ = v0 & ~v7;
  assign \v33.12  = new_n297_ | new_n298_;
  assign new_n300_ = ~v12 & ~v18;
  assign new_n301_ = new_n223_ & new_n300_;
  assign new_n302_ = ~v8 & ~v10;
  assign new_n303_ = v1 & new_n302_;
  assign new_n304_ = v18 & v23;
  assign new_n305_ = new_n82_ & new_n304_;
  assign new_n306_ = new_n303_ & new_n305_;
  assign new_n307_ = ~new_n301_ & ~new_n306_;
  assign new_n308_ = ~v15 & ~new_n307_;
  assign new_n309_ = ~v6 & new_n308_;
  assign new_n310_ = v15 & ~v18;
  assign new_n311_ = ~v14 & new_n310_;
  assign new_n312_ = new_n182_ & new_n311_;
  assign new_n313_ = ~new_n309_ & ~new_n312_;
  assign new_n314_ = ~v28 & ~new_n313_;
  assign new_n315_ = ~v9 & new_n314_;
  assign new_n316_ = ~v15 & v18;
  assign new_n317_ = v18 & ~new_n316_;
  assign new_n318_ = v28 & ~new_n317_;
  assign new_n319_ = v23 & new_n318_;
  assign new_n320_ = v1 & new_n319_;
  assign new_n321_ = ~new_n315_ & ~new_n320_;
  assign new_n322_ = v30 & ~new_n321_;
  assign new_n323_ = v17 & new_n322_;
  assign new_n324_ = ~v16 & new_n323_;
  assign new_n325_ = ~v0 & new_n324_;
  assign \v33.13  = new_n298_ | new_n325_;
  assign new_n327_ = ~v0 & v24;
  assign new_n328_ = ~v25 & ~new_n327_;
  assign new_n329_ = v29 & ~new_n328_;
  assign new_n330_ = v28 & new_n329_;
  assign new_n331_ = v1 & new_n330_;
  assign \v33.14  = v0 | new_n331_;
  assign new_n333_ = ~v0 & v1;
  assign new_n334_ = v13 & new_n333_;
  assign new_n335_ = ~v22 & new_n334_;
  assign new_n336_ = v24 & new_n335_;
  assign new_n337_ = v28 & new_n336_;
  assign \v33.15  = v29 & new_n337_;
  assign new_n339_ = v24 & new_n333_;
  assign new_n340_ = v28 & new_n339_;
  assign \v33.16  = v29 & new_n340_;
  assign new_n342_ = v28 & v30;
  assign new_n343_ = v22 & new_n342_;
  assign new_n344_ = ~v5 & ~new_n343_;
  assign \v33.17  = ~v0 & ~new_n344_;
  assign new_n346_ = v3 & ~v27;
  assign new_n347_ = v26 & ~new_n346_;
  assign new_n348_ = ~v0 & new_n123_;
  assign new_n349_ = ~v28 & v30;
  assign new_n350_ = new_n81_ & new_n349_;
  assign new_n351_ = new_n348_ & new_n350_;
  assign new_n352_ = ~new_n347_ & ~new_n351_;
  assign \v33.18  = v0 | ~new_n352_;
  assign new_n354_ = ~v3 & v27;
  assign new_n355_ = v26 & ~v27;
  assign new_n356_ = v3 & new_n355_;
  assign new_n357_ = ~new_n351_ & ~new_n356_;
  assign new_n358_ = ~new_n354_ & new_n357_;
  assign \v33.19  = v0 | ~new_n358_;
  assign new_n360_ = v19 & ~new_n89_;
  assign new_n361_ = v9 & new_n360_;
  assign new_n362_ = v12 & v21;
  assign new_n363_ = ~v9 & new_n362_;
  assign new_n364_ = ~new_n361_ & ~new_n363_;
  assign new_n365_ = v29 & ~new_n364_;
  assign new_n366_ = v10 & new_n365_;
  assign new_n367_ = ~v10 & ~v12;
  assign new_n368_ = ~v9 & new_n367_;
  assign new_n369_ = ~new_n366_ & ~new_n368_;
  assign new_n370_ = v11 & ~new_n369_;
  assign new_n371_ = v10 & new_n93_;
  assign new_n372_ = ~new_n102_ & ~new_n371_;
  assign new_n373_ = v9 & ~new_n372_;
  assign new_n374_ = ~new_n370_ & ~new_n373_;
  assign new_n375_ = v30 & ~new_n374_;
  assign new_n376_ = ~v28 & new_n375_;
  assign \v33.20  = ~v0 & new_n376_;
  assign new_n378_ = v19 & new_n83_;
  assign new_n379_ = new_n105_ & new_n378_;
  assign new_n380_ = ~new_n93_ & ~new_n379_;
  assign new_n381_ = v10 & ~new_n380_;
  assign new_n382_ = v12 & ~new_n82_;
  assign new_n383_ = v29 & ~new_n382_;
  assign new_n384_ = v21 & new_n383_;
  assign new_n385_ = v20 & new_n384_;
  assign new_n386_ = v19 & new_n385_;
  assign new_n387_ = ~v10 & new_n386_;
  assign new_n388_ = ~new_n381_ & ~new_n387_;
  assign new_n389_ = v9 & ~new_n388_;
  assign new_n390_ = v10 & v11;
  assign new_n391_ = ~v9 & new_n390_;
  assign new_n392_ = v12 & new_n83_;
  assign new_n393_ = new_n391_ & new_n392_;
  assign new_n394_ = ~new_n389_ & ~new_n393_;
  assign new_n395_ = v30 & ~new_n394_;
  assign new_n396_ = ~v29 & ~v30;
  assign new_n397_ = v3 & new_n396_;
  assign new_n398_ = ~new_n395_ & ~new_n397_;
  assign new_n399_ = ~v0 & ~new_n398_;
  assign new_n400_ = ~v3 & v29;
  assign new_n401_ = v2 & ~v29;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign new_n403_ = ~v30 & ~new_n402_;
  assign new_n404_ = ~new_n399_ & ~new_n403_;
  assign new_n405_ = ~v28 & ~new_n404_;
  assign \v33.21  = v0 | new_n405_;
  assign new_n407_ = v3 & ~v30;
  assign new_n408_ = ~v9 & new_n105_;
  assign new_n409_ = v12 & v19;
  assign new_n410_ = v9 & new_n409_;
  assign new_n411_ = v20 & new_n83_;
  assign new_n412_ = new_n410_ & new_n411_;
  assign new_n413_ = ~new_n408_ & ~new_n412_;
  assign new_n414_ = ~v10 & ~new_n413_;
  assign new_n415_ = v10 & new_n82_;
  assign new_n416_ = ~v11 & new_n88_;
  assign new_n417_ = ~new_n415_ & ~new_n416_;
  assign new_n418_ = v29 & ~new_n417_;
  assign new_n419_ = v20 & new_n418_;
  assign new_n420_ = v19 & new_n419_;
  assign new_n421_ = v9 & new_n420_;
  assign new_n422_ = ~new_n414_ & ~new_n421_;
  assign new_n423_ = v30 & ~new_n422_;
  assign new_n424_ = ~new_n407_ & ~new_n423_;
  assign new_n425_ = ~v28 & ~new_n424_;
  assign \v33.22  = ~v0 & new_n425_;
  assign \v33.0  = 1'b0;
endmodule


