// Benchmark "voter" written by ABC on Mon Sep 11 23:43:35 2023

module voter ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_,
    new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_,
    new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_,
    new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_,
    new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_,
    new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_,
    new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_,
    new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_,
    new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_,
    new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_,
    new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4537_, new_n4538_, new_n4539_, new_n4540_,
    new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_,
    new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_,
    new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_,
    new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_,
    new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_,
    new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_,
    new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_,
    new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_,
    new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_,
    new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_,
    new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_,
    new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_,
    new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_,
    new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_,
    new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_,
    new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_,
    new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_,
    new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_,
    new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_,
    new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_,
    new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_,
    new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_,
    new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_,
    new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_,
    new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_,
    new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_,
    new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_,
    new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_,
    new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_,
    new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_,
    new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_,
    new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_,
    new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_,
    new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_,
    new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_,
    new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_,
    new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_,
    new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_,
    new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_,
    new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_,
    new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_,
    new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_,
    new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_,
    new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_,
    new_n6091_, new_n6092_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6106_, new_n6107_, new_n6108_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_,
    new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_,
    new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_,
    new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_,
    new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_,
    new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_,
    new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_,
    new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_,
    new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_,
    new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_,
    new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_,
    new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_,
    new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_,
    new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_,
    new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_,
    new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_,
    new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_,
    new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_,
    new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_,
    new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_,
    new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_,
    new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_,
    new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_,
    new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_,
    new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_,
    new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_,
    new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_,
    new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_,
    new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_,
    new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_,
    new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_,
    new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_,
    new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_,
    new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_,
    new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_,
    new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_,
    new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_,
    new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_,
    new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6867_, new_n6868_,
    new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_,
    new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_,
    new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_,
    new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_,
    new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_,
    new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_,
    new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_,
    new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_,
    new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_,
    new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_,
    new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_,
    new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_,
    new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_,
    new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_,
    new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_,
    new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_,
    new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_,
    new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_,
    new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_,
    new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_,
    new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_,
    new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_,
    new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_,
    new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_,
    new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_,
    new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_,
    new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_,
    new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_,
    new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_,
    new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_,
    new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_,
    new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_,
    new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_,
    new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_,
    new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_,
    new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_,
    new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_,
    new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_,
    new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_,
    new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_,
    new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_,
    new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_,
    new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_,
    new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_,
    new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_,
    new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_,
    new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_,
    new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_,
    new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_,
    new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_,
    new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_,
    new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_,
    new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_,
    new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_,
    new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_,
    new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_,
    new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_,
    new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_,
    new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_,
    new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_,
    new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_,
    new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_,
    new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_,
    new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_,
    new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_,
    new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_,
    new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_,
    new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_,
    new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_,
    new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_,
    new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_,
    new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_,
    new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_,
    new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_,
    new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_,
    new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_,
    new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_,
    new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_,
    new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_,
    new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_,
    new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_,
    new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_,
    new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_,
    new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_,
    new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_,
    new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_,
    new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_,
    new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_,
    new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_,
    new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_,
    new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_,
    new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_,
    new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_,
    new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_,
    new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_,
    new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_,
    new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_,
    new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_,
    new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_,
    new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_,
    new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_,
    new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_,
    new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_,
    new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_,
    new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_,
    new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_,
    new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_,
    new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_,
    new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_,
    new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_,
    new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_,
    new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9018_, new_n9019_, new_n9020_,
    new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_,
    new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_,
    new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_,
    new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_,
    new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_,
    new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_,
    new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_,
    new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_,
    new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_,
    new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_,
    new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_,
    new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_,
    new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_,
    new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_,
    new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_,
    new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_,
    new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_,
    new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_,
    new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_,
    new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_,
    new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_,
    new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_,
    new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_,
    new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_,
    new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_,
    new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_,
    new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_,
    new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_,
    new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_,
    new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_,
    new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_,
    new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_,
    new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_,
    new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_,
    new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_,
    new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_,
    new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_,
    new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_,
    new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_,
    new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_,
    new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_,
    new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_,
    new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_,
    new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_,
    new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_,
    new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_,
    new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_,
    new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_,
    new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_,
    new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_,
    new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_,
    new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_,
    new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_,
    new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_,
    new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_,
    new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_,
    new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_,
    new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_,
    new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_,
    new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_,
    new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_,
    new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_,
    new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_,
    new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_,
    new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_,
    new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_,
    new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_,
    new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_,
    new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_,
    new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_,
    new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_,
    new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_,
    new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_,
    new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_,
    new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_,
    new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_,
    new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_,
    new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_,
    new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_,
    new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_,
    new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_,
    new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_,
    new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_,
    new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_,
    new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_,
    new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_,
    new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_,
    new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_,
    new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_,
    new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_,
    new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_,
    new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_,
    new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_,
    new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_,
    new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_,
    new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_,
    new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_,
    new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_,
    new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_,
    new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_,
    new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_,
    new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10892_, new_n10893_, new_n10894_, new_n10895_, new_n10896_,
    new_n10897_, new_n10898_, new_n10899_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11221_,
    new_n11222_, new_n11223_, new_n11224_, new_n11225_, new_n11226_,
    new_n11227_, new_n11228_, new_n11229_, new_n11230_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11371_,
    new_n11372_, new_n11373_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11392_, new_n11393_, new_n11394_, new_n11395_, new_n11396_,
    new_n11397_, new_n11398_, new_n11399_, new_n11400_, new_n11401_,
    new_n11402_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11415_, new_n11416_,
    new_n11417_, new_n11418_, new_n11419_, new_n11420_, new_n11421_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11440_, new_n11441_,
    new_n11442_, new_n11443_, new_n11444_, new_n11445_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11460_, new_n11461_,
    new_n11462_, new_n11463_, new_n11464_, new_n11465_, new_n11466_,
    new_n11467_, new_n11468_, new_n11469_, new_n11470_, new_n11471_,
    new_n11472_, new_n11473_, new_n11474_, new_n11475_, new_n11476_,
    new_n11477_, new_n11478_, new_n11479_, new_n11480_, new_n11481_,
    new_n11482_, new_n11483_, new_n11484_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11499_, new_n11500_, new_n11501_,
    new_n11502_, new_n11503_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11510_, new_n11511_,
    new_n11512_, new_n11513_, new_n11514_, new_n11515_, new_n11516_,
    new_n11517_, new_n11518_, new_n11519_, new_n11520_, new_n11521_,
    new_n11522_, new_n11523_, new_n11524_, new_n11525_, new_n11526_,
    new_n11527_, new_n11528_, new_n11529_, new_n11530_, new_n11531_,
    new_n11532_, new_n11533_, new_n11534_, new_n11535_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11543_, new_n11544_, new_n11545_, new_n11546_,
    new_n11547_, new_n11548_, new_n11549_, new_n11550_, new_n11551_,
    new_n11552_, new_n11553_, new_n11554_, new_n11555_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11566_,
    new_n11567_, new_n11568_, new_n11569_, new_n11570_, new_n11571_,
    new_n11572_, new_n11573_, new_n11574_, new_n11575_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12100_, new_n12101_,
    new_n12102_, new_n12103_, new_n12104_, new_n12105_, new_n12106_,
    new_n12107_, new_n12108_, new_n12109_, new_n12110_, new_n12111_,
    new_n12112_, new_n12113_, new_n12114_, new_n12115_, new_n12116_,
    new_n12117_, new_n12118_, new_n12119_, new_n12120_, new_n12121_,
    new_n12122_, new_n12123_, new_n12124_, new_n12125_, new_n12126_,
    new_n12127_, new_n12128_, new_n12129_, new_n12130_, new_n12131_,
    new_n12132_, new_n12133_, new_n12134_, new_n12135_, new_n12136_,
    new_n12137_, new_n12138_, new_n12139_, new_n12140_, new_n12141_,
    new_n12142_, new_n12143_, new_n12144_, new_n12145_, new_n12146_,
    new_n12147_, new_n12148_, new_n12149_, new_n12150_, new_n12151_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12158_, new_n12159_, new_n12160_, new_n12161_,
    new_n12162_, new_n12163_, new_n12164_, new_n12165_, new_n12166_,
    new_n12167_, new_n12168_, new_n12169_, new_n12170_, new_n12171_,
    new_n12172_, new_n12173_, new_n12174_, new_n12175_, new_n12176_,
    new_n12177_, new_n12178_, new_n12179_, new_n12180_, new_n12181_,
    new_n12182_, new_n12183_, new_n12184_, new_n12185_, new_n12186_,
    new_n12187_, new_n12188_, new_n12189_, new_n12190_, new_n12191_,
    new_n12192_, new_n12193_, new_n12194_, new_n12195_, new_n12196_,
    new_n12197_, new_n12198_, new_n12199_, new_n12200_, new_n12201_,
    new_n12202_, new_n12203_, new_n12204_, new_n12205_, new_n12206_,
    new_n12207_, new_n12208_, new_n12209_, new_n12210_, new_n12211_,
    new_n12212_, new_n12213_, new_n12214_, new_n12215_, new_n12216_,
    new_n12217_, new_n12218_, new_n12219_, new_n12220_, new_n12221_,
    new_n12222_, new_n12223_, new_n12224_, new_n12225_, new_n12226_,
    new_n12227_, new_n12228_, new_n12229_, new_n12230_, new_n12231_,
    new_n12232_, new_n12233_, new_n12234_, new_n12235_, new_n12236_,
    new_n12237_, new_n12238_, new_n12239_, new_n12240_, new_n12241_,
    new_n12242_, new_n12243_, new_n12244_, new_n12245_, new_n12246_,
    new_n12247_, new_n12248_, new_n12249_, new_n12250_, new_n12251_,
    new_n12252_, new_n12253_, new_n12254_, new_n12255_, new_n12256_,
    new_n12257_, new_n12258_, new_n12259_, new_n12260_, new_n12261_,
    new_n12262_, new_n12263_, new_n12264_, new_n12265_, new_n12266_,
    new_n12267_, new_n12268_, new_n12269_, new_n12270_, new_n12271_,
    new_n12272_, new_n12273_, new_n12274_, new_n12275_, new_n12276_,
    new_n12277_, new_n12278_, new_n12279_, new_n12280_, new_n12281_,
    new_n12282_, new_n12283_, new_n12284_, new_n12285_, new_n12286_,
    new_n12287_, new_n12288_, new_n12289_, new_n12290_, new_n12291_,
    new_n12292_, new_n12293_, new_n12294_, new_n12295_, new_n12296_,
    new_n12297_, new_n12298_, new_n12299_, new_n12300_, new_n12301_,
    new_n12302_, new_n12303_, new_n12304_, new_n12305_, new_n12306_,
    new_n12307_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12327_, new_n12328_, new_n12329_, new_n12330_, new_n12331_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12353_, new_n12354_, new_n12355_, new_n12356_,
    new_n12357_, new_n12358_, new_n12359_, new_n12360_, new_n12361_,
    new_n12362_, new_n12363_, new_n12364_, new_n12365_, new_n12366_,
    new_n12367_, new_n12368_, new_n12369_, new_n12370_, new_n12371_,
    new_n12372_, new_n12373_, new_n12374_, new_n12375_, new_n12376_,
    new_n12377_, new_n12378_, new_n12379_, new_n12380_, new_n12381_,
    new_n12382_, new_n12383_, new_n12384_, new_n12385_, new_n12386_,
    new_n12387_, new_n12388_, new_n12389_, new_n12390_, new_n12391_,
    new_n12392_, new_n12393_, new_n12394_, new_n12395_, new_n12396_,
    new_n12397_, new_n12398_, new_n12399_, new_n12400_, new_n12401_,
    new_n12402_, new_n12403_, new_n12404_, new_n12405_, new_n12406_,
    new_n12407_, new_n12408_, new_n12409_, new_n12410_, new_n12411_,
    new_n12412_, new_n12413_, new_n12414_, new_n12415_, new_n12416_,
    new_n12417_, new_n12418_, new_n12419_, new_n12420_, new_n12421_,
    new_n12422_, new_n12423_, new_n12424_, new_n12425_, new_n12426_,
    new_n12427_, new_n12428_, new_n12429_, new_n12430_, new_n12431_,
    new_n12432_, new_n12433_, new_n12434_, new_n12435_, new_n12436_,
    new_n12437_, new_n12438_, new_n12439_, new_n12440_, new_n12441_,
    new_n12442_, new_n12443_, new_n12444_, new_n12445_, new_n12446_,
    new_n12447_, new_n12448_, new_n12449_, new_n12450_, new_n12451_,
    new_n12452_, new_n12453_, new_n12454_, new_n12455_, new_n12456_,
    new_n12457_, new_n12458_, new_n12459_, new_n12460_, new_n12461_,
    new_n12462_, new_n12463_, new_n12464_, new_n12465_, new_n12466_,
    new_n12467_, new_n12468_, new_n12469_, new_n12470_, new_n12471_,
    new_n12472_, new_n12473_, new_n12474_, new_n12475_, new_n12476_,
    new_n12477_, new_n12478_, new_n12479_, new_n12480_, new_n12481_,
    new_n12482_, new_n12483_, new_n12484_, new_n12485_, new_n12486_,
    new_n12487_, new_n12488_, new_n12489_, new_n12490_, new_n12491_,
    new_n12492_, new_n12493_, new_n12494_, new_n12495_, new_n12496_,
    new_n12497_, new_n12498_, new_n12499_, new_n12500_, new_n12501_,
    new_n12502_, new_n12503_, new_n12504_, new_n12505_, new_n12506_,
    new_n12507_, new_n12508_, new_n12509_, new_n12510_, new_n12511_,
    new_n12512_, new_n12513_, new_n12514_, new_n12515_, new_n12516_,
    new_n12517_, new_n12518_, new_n12519_, new_n12520_, new_n12521_,
    new_n12522_, new_n12523_, new_n12524_, new_n12525_, new_n12526_,
    new_n12527_, new_n12528_, new_n12529_, new_n12530_, new_n12531_,
    new_n12532_, new_n12533_, new_n12534_, new_n12535_, new_n12536_,
    new_n12537_, new_n12538_, new_n12539_, new_n12540_, new_n12541_,
    new_n12542_, new_n12543_, new_n12544_, new_n12545_, new_n12546_,
    new_n12547_, new_n12548_, new_n12549_, new_n12550_, new_n12551_,
    new_n12552_, new_n12553_, new_n12554_, new_n12555_, new_n12556_,
    new_n12557_, new_n12558_, new_n12559_, new_n12560_, new_n12561_,
    new_n12562_, new_n12563_, new_n12564_, new_n12565_, new_n12566_,
    new_n12567_, new_n12568_, new_n12569_, new_n12570_, new_n12571_,
    new_n12572_, new_n12573_, new_n12574_, new_n12575_, new_n12576_,
    new_n12577_, new_n12578_, new_n12579_, new_n12580_, new_n12581_,
    new_n12582_, new_n12583_, new_n12584_, new_n12585_, new_n12586_,
    new_n12587_, new_n12588_, new_n12589_, new_n12590_, new_n12591_,
    new_n12592_, new_n12593_, new_n12594_, new_n12595_, new_n12596_,
    new_n12597_, new_n12598_, new_n12599_, new_n12600_, new_n12601_,
    new_n12602_, new_n12603_, new_n12604_, new_n12605_, new_n12606_,
    new_n12607_, new_n12608_, new_n12609_, new_n12610_, new_n12611_,
    new_n12612_, new_n12613_, new_n12614_, new_n12615_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12629_, new_n12630_, new_n12631_,
    new_n12632_, new_n12633_, new_n12634_, new_n12635_, new_n12636_,
    new_n12637_, new_n12638_, new_n12639_, new_n12640_, new_n12641_,
    new_n12642_, new_n12643_, new_n12644_, new_n12645_, new_n12646_,
    new_n12647_, new_n12648_, new_n12649_, new_n12650_, new_n12651_,
    new_n12652_, new_n12653_, new_n12654_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12664_, new_n12665_, new_n12666_,
    new_n12667_, new_n12668_, new_n12669_, new_n12670_, new_n12671_,
    new_n12672_, new_n12673_, new_n12674_, new_n12675_, new_n12676_,
    new_n12677_, new_n12678_, new_n12679_, new_n12680_, new_n12681_,
    new_n12682_, new_n12683_, new_n12684_, new_n12685_, new_n12686_,
    new_n12687_, new_n12688_, new_n12689_, new_n12690_, new_n12691_,
    new_n12692_, new_n12693_, new_n12694_, new_n12695_, new_n12696_,
    new_n12697_, new_n12698_, new_n12699_, new_n12700_, new_n12701_,
    new_n12702_, new_n12703_, new_n12704_, new_n12705_, new_n12706_,
    new_n12707_, new_n12708_, new_n12709_, new_n12710_, new_n12711_,
    new_n12712_, new_n12713_, new_n12714_, new_n12715_, new_n12716_,
    new_n12717_, new_n12718_, new_n12719_, new_n12720_, new_n12721_,
    new_n12722_, new_n12723_, new_n12724_, new_n12725_, new_n12726_,
    new_n12727_, new_n12728_, new_n12729_, new_n12730_, new_n12731_,
    new_n12732_, new_n12733_, new_n12734_, new_n12735_, new_n12736_,
    new_n12737_, new_n12738_, new_n12739_, new_n12740_, new_n12741_,
    new_n12742_, new_n12743_, new_n12744_, new_n12745_, new_n12746_,
    new_n12747_, new_n12748_, new_n12749_, new_n12750_, new_n12751_,
    new_n12752_, new_n12753_, new_n12754_, new_n12755_, new_n12756_,
    new_n12757_, new_n12758_, new_n12759_, new_n12760_, new_n12761_,
    new_n12762_, new_n12763_, new_n12764_, new_n12765_, new_n12766_,
    new_n12767_, new_n12768_, new_n12769_, new_n12770_, new_n12771_,
    new_n12772_, new_n12773_, new_n12774_, new_n12775_, new_n12776_,
    new_n12777_, new_n12778_, new_n12779_, new_n12780_, new_n12781_,
    new_n12782_, new_n12783_, new_n12784_, new_n12785_, new_n12786_,
    new_n12787_, new_n12788_, new_n12789_, new_n12790_, new_n12791_,
    new_n12792_, new_n12793_, new_n12794_, new_n12795_, new_n12796_,
    new_n12797_, new_n12798_, new_n12799_, new_n12800_, new_n12801_,
    new_n12802_, new_n12803_, new_n12804_, new_n12805_, new_n12806_,
    new_n12807_, new_n12808_, new_n12809_, new_n12810_, new_n12811_,
    new_n12812_, new_n12813_, new_n12814_, new_n12815_, new_n12816_,
    new_n12817_, new_n12818_, new_n12819_, new_n12820_, new_n12821_,
    new_n12822_, new_n12823_, new_n12824_, new_n12825_, new_n12826_,
    new_n12827_, new_n12828_, new_n12829_, new_n12830_, new_n12831_,
    new_n12832_, new_n12833_, new_n12834_, new_n12835_, new_n12836_,
    new_n12837_, new_n12838_, new_n12839_, new_n12840_, new_n12841_,
    new_n12842_, new_n12843_, new_n12844_, new_n12845_, new_n12846_,
    new_n12847_, new_n12848_, new_n12849_, new_n12850_, new_n12851_,
    new_n12852_, new_n12853_, new_n12854_, new_n12855_, new_n12856_,
    new_n12857_, new_n12858_, new_n12859_, new_n12860_, new_n12861_,
    new_n12862_, new_n12863_, new_n12864_, new_n12865_, new_n12866_,
    new_n12867_, new_n12868_, new_n12869_, new_n12870_, new_n12871_,
    new_n12872_, new_n12873_, new_n12874_, new_n12875_, new_n12876_,
    new_n12877_, new_n12878_, new_n12879_, new_n12880_, new_n12881_,
    new_n12882_, new_n12883_, new_n12884_, new_n12885_, new_n12886_,
    new_n12887_, new_n12888_, new_n12889_, new_n12890_, new_n12891_,
    new_n12892_, new_n12893_, new_n12894_, new_n12895_, new_n12896_,
    new_n12897_, new_n12898_, new_n12899_, new_n12900_, new_n12901_,
    new_n12902_, new_n12903_, new_n12904_, new_n12905_, new_n12906_,
    new_n12907_, new_n12908_, new_n12909_, new_n12910_, new_n12911_,
    new_n12912_, new_n12913_, new_n12914_, new_n12915_, new_n12916_,
    new_n12917_, new_n12918_, new_n12919_, new_n12920_, new_n12921_,
    new_n12922_, new_n12923_, new_n12924_, new_n12925_, new_n12926_,
    new_n12927_, new_n12928_, new_n12929_, new_n12930_, new_n12931_,
    new_n12932_, new_n12933_, new_n12934_, new_n12935_, new_n12936_,
    new_n12937_, new_n12938_, new_n12939_, new_n12940_, new_n12941_,
    new_n12942_, new_n12943_, new_n12944_, new_n12945_, new_n12946_,
    new_n12947_, new_n12948_, new_n12949_, new_n12950_, new_n12951_,
    new_n12952_, new_n12953_, new_n12954_, new_n12955_, new_n12956_,
    new_n12957_, new_n12958_, new_n12959_, new_n12960_, new_n12961_,
    new_n12962_, new_n12963_, new_n12964_, new_n12965_, new_n12966_,
    new_n12967_, new_n12968_, new_n12969_, new_n12970_, new_n12971_,
    new_n12972_, new_n12973_, new_n12974_, new_n12975_, new_n12976_,
    new_n12977_, new_n12978_, new_n12979_, new_n12980_, new_n12981_,
    new_n12982_, new_n12983_, new_n12984_, new_n12985_, new_n12986_,
    new_n12987_, new_n12988_, new_n12989_, new_n12990_, new_n12991_,
    new_n12992_, new_n12993_, new_n12994_, new_n12995_, new_n12996_,
    new_n12997_, new_n12998_, new_n12999_, new_n13000_, new_n13001_,
    new_n13002_, new_n13003_, new_n13004_, new_n13005_, new_n13006_,
    new_n13007_, new_n13008_, new_n13009_, new_n13010_, new_n13011_,
    new_n13012_, new_n13013_, new_n13014_, new_n13015_, new_n13016_,
    new_n13017_, new_n13018_, new_n13019_, new_n13020_, new_n13021_,
    new_n13022_, new_n13023_, new_n13024_, new_n13025_, new_n13026_,
    new_n13027_, new_n13028_, new_n13029_, new_n13030_, new_n13031_,
    new_n13032_, new_n13033_, new_n13034_, new_n13035_, new_n13036_,
    new_n13037_, new_n13038_, new_n13039_, new_n13040_, new_n13041_,
    new_n13042_, new_n13043_, new_n13044_, new_n13045_, new_n13046_,
    new_n13047_, new_n13048_, new_n13049_, new_n13050_, new_n13051_,
    new_n13052_, new_n13053_, new_n13054_, new_n13055_, new_n13056_,
    new_n13057_, new_n13058_, new_n13059_, new_n13060_, new_n13061_,
    new_n13062_, new_n13063_, new_n13064_, new_n13065_, new_n13066_,
    new_n13067_, new_n13068_, new_n13069_, new_n13070_, new_n13071_,
    new_n13072_, new_n13073_, new_n13074_, new_n13075_, new_n13076_,
    new_n13077_, new_n13078_, new_n13079_, new_n13080_, new_n13081_,
    new_n13082_, new_n13083_, new_n13084_, new_n13085_, new_n13086_,
    new_n13087_, new_n13088_, new_n13089_, new_n13090_, new_n13091_,
    new_n13092_, new_n13093_, new_n13094_, new_n13095_, new_n13096_,
    new_n13097_, new_n13098_, new_n13099_, new_n13100_, new_n13101_,
    new_n13102_, new_n13103_, new_n13104_, new_n13105_, new_n13106_,
    new_n13107_, new_n13108_, new_n13109_, new_n13110_, new_n13111_,
    new_n13112_, new_n13113_, new_n13114_, new_n13115_, new_n13116_,
    new_n13117_, new_n13118_, new_n13119_, new_n13120_, new_n13121_,
    new_n13122_, new_n13123_, new_n13124_, new_n13125_, new_n13126_,
    new_n13127_, new_n13128_, new_n13129_, new_n13130_, new_n13131_,
    new_n13132_, new_n13133_, new_n13134_, new_n13135_, new_n13136_,
    new_n13137_, new_n13138_, new_n13139_, new_n13140_, new_n13141_,
    new_n13142_, new_n13143_, new_n13144_, new_n13145_, new_n13146_,
    new_n13147_, new_n13148_, new_n13149_, new_n13150_, new_n13151_,
    new_n13152_, new_n13153_, new_n13154_, new_n13155_, new_n13156_,
    new_n13157_, new_n13158_, new_n13159_, new_n13160_, new_n13161_,
    new_n13162_, new_n13163_, new_n13164_, new_n13165_, new_n13166_,
    new_n13167_, new_n13168_, new_n13169_, new_n13170_, new_n13171_,
    new_n13172_, new_n13173_, new_n13174_, new_n13175_, new_n13176_,
    new_n13177_, new_n13178_, new_n13179_, new_n13180_, new_n13181_,
    new_n13182_, new_n13183_, new_n13184_, new_n13185_, new_n13186_,
    new_n13187_, new_n13188_, new_n13189_, new_n13190_, new_n13191_,
    new_n13192_, new_n13193_, new_n13194_, new_n13195_, new_n13196_,
    new_n13197_, new_n13198_, new_n13199_, new_n13200_, new_n13201_,
    new_n13202_, new_n13203_, new_n13204_, new_n13205_, new_n13206_,
    new_n13207_, new_n13208_, new_n13209_, new_n13210_, new_n13211_,
    new_n13212_, new_n13213_, new_n13214_, new_n13215_, new_n13216_,
    new_n13217_, new_n13218_, new_n13219_, new_n13220_, new_n13221_,
    new_n13222_, new_n13223_, new_n13224_, new_n13225_, new_n13226_,
    new_n13227_, new_n13228_, new_n13229_, new_n13230_, new_n13231_,
    new_n13232_, new_n13233_, new_n13234_, new_n13235_, new_n13236_,
    new_n13237_, new_n13238_, new_n13239_, new_n13240_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13245_, new_n13246_,
    new_n13247_, new_n13248_, new_n13249_, new_n13250_, new_n13251_,
    new_n13252_, new_n13253_, new_n13254_, new_n13255_, new_n13256_,
    new_n13257_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13262_, new_n13263_, new_n13264_, new_n13265_, new_n13266_,
    new_n13267_, new_n13268_, new_n13269_, new_n13270_, new_n13271_,
    new_n13272_, new_n13273_, new_n13274_, new_n13275_, new_n13276_,
    new_n13277_, new_n13278_, new_n13279_, new_n13280_, new_n13281_,
    new_n13282_, new_n13283_, new_n13284_, new_n13285_, new_n13286_,
    new_n13287_, new_n13288_, new_n13289_, new_n13290_, new_n13291_,
    new_n13292_, new_n13293_, new_n13294_, new_n13295_, new_n13296_,
    new_n13297_, new_n13298_, new_n13299_, new_n13300_, new_n13301_,
    new_n13302_, new_n13303_, new_n13304_, new_n13305_, new_n13306_,
    new_n13307_, new_n13308_, new_n13309_, new_n13310_, new_n13311_,
    new_n13312_, new_n13313_, new_n13314_, new_n13315_, new_n13316_,
    new_n13317_, new_n13318_, new_n13319_, new_n13320_, new_n13321_,
    new_n13322_, new_n13323_, new_n13324_, new_n13325_, new_n13326_,
    new_n13327_, new_n13328_, new_n13329_, new_n13330_, new_n13331_,
    new_n13332_, new_n13333_, new_n13334_, new_n13335_, new_n13336_,
    new_n13337_, new_n13338_, new_n13339_, new_n13340_, new_n13341_,
    new_n13342_, new_n13343_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13354_, new_n13355_, new_n13356_,
    new_n13357_, new_n13358_, new_n13359_, new_n13360_, new_n13361_,
    new_n13362_, new_n13363_, new_n13364_, new_n13365_, new_n13366_,
    new_n13367_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13373_, new_n13374_, new_n13375_, new_n13376_,
    new_n13377_, new_n13378_, new_n13379_, new_n13380_, new_n13381_,
    new_n13382_, new_n13383_, new_n13384_, new_n13385_, new_n13386_,
    new_n13387_, new_n13388_, new_n13389_, new_n13390_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13395_, new_n13396_,
    new_n13397_, new_n13398_, new_n13399_, new_n13400_, new_n13401_,
    new_n13402_, new_n13403_, new_n13404_, new_n13405_, new_n13406_,
    new_n13407_, new_n13408_, new_n13409_, new_n13410_, new_n13411_,
    new_n13412_, new_n13413_, new_n13414_, new_n13415_, new_n13416_,
    new_n13417_, new_n13418_, new_n13419_, new_n13420_, new_n13421_,
    new_n13422_, new_n13423_, new_n13424_, new_n13425_, new_n13426_,
    new_n13427_, new_n13428_, new_n13429_, new_n13430_, new_n13431_,
    new_n13432_, new_n13433_, new_n13434_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13473_, new_n13474_, new_n13475_, new_n13476_,
    new_n13477_, new_n13478_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14445_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14456_,
    new_n14457_, new_n14458_, new_n14459_, new_n14460_, new_n14461_,
    new_n14462_, new_n14463_, new_n14464_, new_n14465_, new_n14466_,
    new_n14467_, new_n14468_, new_n14469_, new_n14470_, new_n14471_,
    new_n14472_, new_n14473_, new_n14474_, new_n14475_, new_n14476_,
    new_n14477_, new_n14478_, new_n14479_, new_n14480_, new_n14481_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14487_, new_n14488_, new_n14489_, new_n14490_, new_n14491_,
    new_n14492_, new_n14493_, new_n14494_, new_n14495_, new_n14496_,
    new_n14497_, new_n14498_, new_n14499_, new_n14500_, new_n14501_,
    new_n14502_, new_n14503_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14522_, new_n14523_, new_n14524_, new_n14525_, new_n14526_,
    new_n14527_, new_n14528_, new_n14529_, new_n14530_, new_n14531_,
    new_n14532_, new_n14533_, new_n14534_, new_n14535_, new_n14536_,
    new_n14537_, new_n14538_, new_n14539_, new_n14540_, new_n14541_,
    new_n14542_, new_n14543_, new_n14544_, new_n14545_, new_n14546_,
    new_n14547_, new_n14548_, new_n14549_, new_n14550_, new_n14551_,
    new_n14552_, new_n14553_, new_n14554_, new_n14555_, new_n14556_,
    new_n14557_, new_n14558_, new_n14559_, new_n14560_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14575_, new_n14576_,
    new_n14577_, new_n14578_, new_n14579_, new_n14580_, new_n14581_,
    new_n14582_, new_n14583_, new_n14584_, new_n14585_, new_n14586_,
    new_n14587_, new_n14588_, new_n14589_, new_n14590_, new_n14591_,
    new_n14592_, new_n14593_, new_n14594_, new_n14595_, new_n14596_,
    new_n14597_, new_n14598_, new_n14599_, new_n14600_, new_n14601_,
    new_n14602_, new_n14603_, new_n14604_, new_n14605_, new_n14606_,
    new_n14607_, new_n14608_, new_n14609_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14620_, new_n14621_,
    new_n14622_, new_n14623_, new_n14624_, new_n14625_, new_n14626_,
    new_n14627_, new_n14628_, new_n14629_, new_n14630_, new_n14631_,
    new_n14632_, new_n14633_, new_n14634_, new_n14635_, new_n14636_,
    new_n14637_, new_n14638_, new_n14639_, new_n14640_, new_n14641_,
    new_n14642_, new_n14643_, new_n14644_, new_n14645_, new_n14646_,
    new_n14647_, new_n14648_, new_n14649_, new_n14650_, new_n14651_,
    new_n14652_, new_n14653_, new_n14654_, new_n14655_, new_n14656_,
    new_n14657_, new_n14658_, new_n14659_, new_n14660_, new_n14661_,
    new_n14662_, new_n14663_, new_n14664_, new_n14665_, new_n14666_,
    new_n14667_, new_n14668_, new_n14669_, new_n14670_, new_n14671_,
    new_n14672_, new_n14673_, new_n14674_, new_n14675_, new_n14676_,
    new_n14677_, new_n14678_, new_n14679_, new_n14680_, new_n14681_,
    new_n14682_, new_n14683_, new_n14684_, new_n14685_, new_n14686_,
    new_n14687_, new_n14688_, new_n14689_, new_n14690_, new_n14691_,
    new_n14692_, new_n14693_, new_n14694_, new_n14695_, new_n14696_,
    new_n14697_, new_n14698_, new_n14699_, new_n14700_, new_n14701_,
    new_n14702_, new_n14703_, new_n14704_, new_n14705_, new_n14706_,
    new_n14707_, new_n14708_, new_n14709_, new_n14710_, new_n14711_,
    new_n14712_, new_n14713_, new_n14714_, new_n14715_, new_n14716_,
    new_n14717_, new_n14718_, new_n14719_, new_n14720_, new_n14721_,
    new_n14722_, new_n14723_, new_n14724_, new_n14725_, new_n14726_,
    new_n14727_, new_n14728_, new_n14729_, new_n14730_, new_n14731_,
    new_n14732_, new_n14733_, new_n14734_, new_n14735_, new_n14736_,
    new_n14737_, new_n14738_, new_n14739_, new_n14740_, new_n14741_,
    new_n14742_, new_n14743_, new_n14744_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14781_,
    new_n14782_, new_n14783_, new_n14784_, new_n14785_, new_n14786_,
    new_n14787_, new_n14788_, new_n14789_, new_n14790_, new_n14791_,
    new_n14792_, new_n14793_, new_n14794_, new_n14795_, new_n14796_,
    new_n14797_, new_n14798_, new_n14799_, new_n14800_, new_n14801_,
    new_n14802_, new_n14803_, new_n14804_, new_n14805_, new_n14806_,
    new_n14807_, new_n14808_, new_n14809_, new_n14810_, new_n14811_,
    new_n14812_, new_n14813_, new_n14814_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14958_, new_n14959_, new_n14960_, new_n14961_,
    new_n14962_, new_n14963_, new_n14964_, new_n14965_, new_n14966_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14976_,
    new_n14977_, new_n14978_, new_n14979_, new_n14980_, new_n14981_,
    new_n14982_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15113_, new_n15114_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15127_, new_n15128_, new_n15129_, new_n15130_, new_n15131_,
    new_n15132_, new_n15133_, new_n15134_, new_n15135_, new_n15136_,
    new_n15137_, new_n15138_, new_n15139_, new_n15140_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15179_, new_n15180_, new_n15181_,
    new_n15182_, new_n15183_, new_n15184_, new_n15185_, new_n15186_,
    new_n15187_, new_n15188_, new_n15189_, new_n15190_, new_n15191_,
    new_n15192_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15206_,
    new_n15207_, new_n15208_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15213_, new_n15214_, new_n15215_, new_n15216_,
    new_n15217_, new_n15218_, new_n15219_, new_n15220_, new_n15221_,
    new_n15222_, new_n15223_, new_n15224_, new_n15225_, new_n15226_,
    new_n15227_, new_n15228_, new_n15229_, new_n15230_, new_n15231_,
    new_n15232_, new_n15233_, new_n15234_, new_n15235_, new_n15236_,
    new_n15237_, new_n15238_, new_n15239_, new_n15240_, new_n15241_,
    new_n15242_, new_n15243_, new_n15244_, new_n15245_, new_n15246_,
    new_n15247_, new_n15248_, new_n15249_, new_n15250_, new_n15251_,
    new_n15252_, new_n15253_, new_n15254_, new_n15255_, new_n15256_,
    new_n15257_, new_n15258_, new_n15259_, new_n15260_, new_n15261_,
    new_n15262_, new_n15263_, new_n15264_, new_n15265_, new_n15266_,
    new_n15267_, new_n15268_, new_n15269_, new_n15270_, new_n15271_,
    new_n15272_, new_n15273_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15280_, new_n15281_,
    new_n15282_, new_n15283_, new_n15284_, new_n15285_, new_n15286_,
    new_n15287_, new_n15288_, new_n15289_, new_n15290_, new_n15291_,
    new_n15292_, new_n15293_, new_n15294_, new_n15295_, new_n15296_,
    new_n15297_, new_n15298_, new_n15299_, new_n15300_, new_n15301_,
    new_n15302_, new_n15303_, new_n15304_, new_n15305_, new_n15306_,
    new_n15307_, new_n15308_, new_n15309_, new_n15310_, new_n15311_,
    new_n15312_, new_n15313_, new_n15314_, new_n15315_, new_n15316_,
    new_n15317_, new_n15318_, new_n15319_, new_n15320_, new_n15321_,
    new_n15322_, new_n15323_, new_n15324_, new_n15325_, new_n15326_,
    new_n15327_, new_n15328_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15434_, new_n15435_, new_n15436_,
    new_n15437_, new_n15438_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15470_, new_n15471_,
    new_n15472_, new_n15473_, new_n15474_, new_n15475_, new_n15476_,
    new_n15477_, new_n15478_, new_n15479_, new_n15480_, new_n15481_,
    new_n15482_, new_n15483_, new_n15484_, new_n15485_, new_n15486_,
    new_n15487_, new_n15488_, new_n15489_, new_n15490_, new_n15491_,
    new_n15492_, new_n15493_, new_n15494_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15544_, new_n15545_, new_n15546_,
    new_n15547_, new_n15548_, new_n15549_, new_n15550_, new_n15551_,
    new_n15552_, new_n15553_, new_n15554_, new_n15555_, new_n15556_,
    new_n15557_, new_n15558_, new_n15559_, new_n15560_, new_n15561_,
    new_n15562_, new_n15563_, new_n15564_, new_n15565_, new_n15566_,
    new_n15567_, new_n15568_, new_n15569_, new_n15570_, new_n15571_,
    new_n15572_, new_n15573_, new_n15574_, new_n15575_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15580_, new_n15581_,
    new_n15582_, new_n15583_, new_n15584_, new_n15585_, new_n15586_,
    new_n15587_, new_n15588_, new_n15589_, new_n15590_, new_n15591_,
    new_n15592_, new_n15593_, new_n15594_, new_n15595_, new_n15596_,
    new_n15597_, new_n15598_, new_n15599_, new_n15600_, new_n15601_,
    new_n15602_, new_n15603_, new_n15604_, new_n15605_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15611_,
    new_n15612_, new_n15613_, new_n15614_, new_n15615_, new_n15616_,
    new_n15617_, new_n15618_, new_n15619_, new_n15620_, new_n15621_,
    new_n15622_, new_n15623_, new_n15624_, new_n15625_, new_n15626_,
    new_n15627_, new_n15628_, new_n15629_, new_n15630_, new_n15631_,
    new_n15632_, new_n15633_, new_n15634_, new_n15635_, new_n15636_,
    new_n15637_, new_n15638_, new_n15639_, new_n15640_, new_n15641_,
    new_n15642_, new_n15643_, new_n15644_, new_n15645_, new_n15646_,
    new_n15647_, new_n15648_, new_n15649_, new_n15650_, new_n15651_,
    new_n15652_, new_n15653_, new_n15654_, new_n15655_, new_n15656_,
    new_n15657_, new_n15658_, new_n15659_, new_n15660_, new_n15661_,
    new_n15662_, new_n15663_, new_n15664_, new_n15665_, new_n15666_,
    new_n15667_, new_n15668_, new_n15669_, new_n15670_, new_n15671_,
    new_n15672_, new_n15673_, new_n15674_, new_n15675_, new_n15676_,
    new_n15677_, new_n15678_, new_n15679_, new_n15680_, new_n15681_,
    new_n15682_, new_n15683_, new_n15684_, new_n15685_, new_n15686_,
    new_n15687_, new_n15688_, new_n15689_, new_n15690_, new_n15691_,
    new_n15692_, new_n15693_, new_n15694_, new_n15695_, new_n15696_,
    new_n15697_, new_n15698_, new_n15699_, new_n15700_, new_n15701_,
    new_n15702_, new_n15703_, new_n15704_, new_n15705_, new_n15706_,
    new_n15707_, new_n15708_, new_n15709_, new_n15710_, new_n15711_,
    new_n15712_, new_n15713_, new_n15714_, new_n15715_, new_n15716_,
    new_n15717_, new_n15718_, new_n15719_, new_n15720_, new_n15721_,
    new_n15722_, new_n15723_, new_n15724_, new_n15725_, new_n15726_,
    new_n15727_, new_n15728_, new_n15729_, new_n15730_, new_n15731_,
    new_n15732_, new_n15733_, new_n15734_, new_n15735_, new_n15736_,
    new_n15737_, new_n15738_, new_n15739_, new_n15740_, new_n15741_,
    new_n15742_, new_n15743_, new_n15744_, new_n15745_, new_n15746_,
    new_n15747_, new_n15748_, new_n15749_, new_n15750_, new_n15751_,
    new_n15752_, new_n15753_, new_n15754_, new_n15755_, new_n15756_,
    new_n15757_, new_n15758_, new_n15759_, new_n15760_, new_n15761_,
    new_n15762_, new_n15763_, new_n15764_, new_n15765_, new_n15766_,
    new_n15767_, new_n15768_, new_n15769_, new_n15770_, new_n15771_,
    new_n15772_, new_n15773_, new_n15774_, new_n15775_, new_n15776_,
    new_n15777_, new_n15778_, new_n15779_, new_n15780_, new_n15781_,
    new_n15782_, new_n15783_, new_n15784_, new_n15785_, new_n15786_,
    new_n15787_, new_n15788_, new_n15789_, new_n15790_, new_n15791_,
    new_n15792_, new_n15793_, new_n15794_, new_n15795_, new_n15796_,
    new_n15797_, new_n15798_, new_n15799_, new_n15800_, new_n15801_,
    new_n15802_, new_n15803_, new_n15804_, new_n15805_, new_n15806_,
    new_n15807_, new_n15808_, new_n15809_, new_n15810_, new_n15811_,
    new_n15812_, new_n15813_, new_n15814_, new_n15815_, new_n15816_,
    new_n15817_, new_n15818_, new_n15819_, new_n15820_, new_n15821_,
    new_n15822_, new_n15823_, new_n15824_, new_n15825_, new_n15826_,
    new_n15827_, new_n15828_, new_n15829_, new_n15830_, new_n15831_,
    new_n15832_, new_n15833_, new_n15834_, new_n15835_, new_n15836_,
    new_n15837_, new_n15838_, new_n15839_, new_n15840_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15850_, new_n15851_,
    new_n15852_, new_n15853_, new_n15854_, new_n15855_, new_n15856_,
    new_n15857_, new_n15858_, new_n15859_, new_n15860_, new_n15861_,
    new_n15862_, new_n15863_, new_n15864_, new_n15865_, new_n15866_,
    new_n15867_, new_n15868_, new_n15869_, new_n15870_, new_n15871_,
    new_n15872_, new_n15873_, new_n15874_, new_n15875_, new_n15876_,
    new_n15877_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15889_, new_n15890_, new_n15891_,
    new_n15892_, new_n15893_, new_n15894_, new_n15895_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15925_, new_n15926_,
    new_n15927_, new_n15928_, new_n15929_, new_n15930_, new_n15931_,
    new_n15932_, new_n15933_, new_n15934_, new_n15935_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16011_,
    new_n16012_, new_n16013_, new_n16014_, new_n16015_, new_n16016_,
    new_n16017_, new_n16018_, new_n16019_, new_n16020_, new_n16021_,
    new_n16022_, new_n16023_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16040_, new_n16041_,
    new_n16042_, new_n16043_, new_n16044_, new_n16045_, new_n16046_,
    new_n16047_, new_n16048_, new_n16049_, new_n16050_, new_n16051_,
    new_n16052_, new_n16053_, new_n16054_, new_n16055_, new_n16056_,
    new_n16057_, new_n16058_, new_n16059_, new_n16060_, new_n16061_,
    new_n16062_, new_n16063_, new_n16064_, new_n16065_, new_n16066_,
    new_n16067_, new_n16068_, new_n16069_, new_n16070_, new_n16071_,
    new_n16072_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16082_, new_n16083_, new_n16084_, new_n16085_, new_n16086_,
    new_n16087_, new_n16088_, new_n16089_, new_n16090_, new_n16091_,
    new_n16092_, new_n16093_, new_n16094_, new_n16095_, new_n16096_,
    new_n16097_, new_n16098_, new_n16099_, new_n16100_, new_n16101_,
    new_n16102_, new_n16103_, new_n16104_, new_n16105_, new_n16106_,
    new_n16107_, new_n16108_, new_n16109_, new_n16110_, new_n16111_,
    new_n16112_, new_n16113_, new_n16114_, new_n16115_, new_n16116_,
    new_n16117_, new_n16118_, new_n16119_, new_n16120_, new_n16121_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16164_, new_n16165_, new_n16166_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16295_, new_n16296_,
    new_n16297_, new_n16298_, new_n16299_, new_n16300_, new_n16301_,
    new_n16302_, new_n16303_, new_n16304_, new_n16305_, new_n16306_,
    new_n16307_, new_n16308_, new_n16309_, new_n16310_, new_n16311_,
    new_n16312_, new_n16313_, new_n16314_, new_n16315_, new_n16316_,
    new_n16317_, new_n16318_, new_n16319_, new_n16320_, new_n16321_,
    new_n16322_, new_n16323_, new_n16324_, new_n16325_, new_n16326_,
    new_n16327_, new_n16328_, new_n16329_, new_n16330_, new_n16331_,
    new_n16332_, new_n16333_, new_n16334_, new_n16335_, new_n16336_,
    new_n16337_, new_n16338_, new_n16339_, new_n16340_, new_n16341_,
    new_n16342_, new_n16343_, new_n16344_, new_n16345_, new_n16346_,
    new_n16347_, new_n16348_, new_n16349_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17283_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17328_, new_n17329_, new_n17330_, new_n17331_,
    new_n17332_, new_n17333_, new_n17334_, new_n17335_, new_n17336_,
    new_n17337_, new_n17338_, new_n17339_, new_n17340_, new_n17341_,
    new_n17342_, new_n17343_, new_n17344_, new_n17345_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17361_,
    new_n17362_, new_n17363_, new_n17364_, new_n17365_, new_n17366_,
    new_n17367_, new_n17368_, new_n17369_, new_n17370_, new_n17371_,
    new_n17372_, new_n17373_, new_n17374_, new_n17375_, new_n17376_,
    new_n17377_, new_n17378_, new_n17379_, new_n17380_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17398_, new_n17399_, new_n17400_, new_n17401_,
    new_n17402_, new_n17403_, new_n17404_, new_n17405_, new_n17406_,
    new_n17407_, new_n17408_, new_n17409_, new_n17410_, new_n17411_,
    new_n17412_, new_n17413_, new_n17414_, new_n17415_, new_n17416_,
    new_n17417_, new_n17418_, new_n17419_, new_n17420_, new_n17421_,
    new_n17422_, new_n17423_, new_n17424_, new_n17425_, new_n17426_,
    new_n17427_, new_n17428_, new_n17429_, new_n17430_, new_n17431_,
    new_n17432_, new_n17433_, new_n17434_, new_n17435_, new_n17436_,
    new_n17437_, new_n17438_, new_n17439_, new_n17440_, new_n17441_,
    new_n17442_, new_n17443_, new_n17444_, new_n17445_, new_n17446_,
    new_n17447_, new_n17448_, new_n17449_, new_n17450_, new_n17451_,
    new_n17452_, new_n17453_, new_n17454_, new_n17455_, new_n17456_,
    new_n17457_, new_n17458_, new_n17459_, new_n17460_, new_n17461_,
    new_n17462_, new_n17463_, new_n17464_, new_n17465_, new_n17466_,
    new_n17467_, new_n17468_, new_n17469_, new_n17470_, new_n17471_,
    new_n17472_, new_n17473_, new_n17474_, new_n17475_, new_n17476_,
    new_n17477_, new_n17478_, new_n17479_, new_n17480_, new_n17481_,
    new_n17482_, new_n17483_, new_n17484_, new_n17485_, new_n17486_,
    new_n17487_, new_n17488_, new_n17489_, new_n17490_, new_n17491_,
    new_n17492_, new_n17493_, new_n17494_, new_n17495_, new_n17496_,
    new_n17497_, new_n17498_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17504_, new_n17505_, new_n17506_,
    new_n17507_, new_n17508_, new_n17509_, new_n17510_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17516_,
    new_n17517_, new_n17518_, new_n17519_, new_n17520_, new_n17521_,
    new_n17522_, new_n17523_, new_n17524_, new_n17525_, new_n17526_,
    new_n17527_, new_n17528_, new_n17529_, new_n17530_, new_n17531_,
    new_n17532_, new_n17533_, new_n17534_, new_n17535_, new_n17536_,
    new_n17537_, new_n17538_, new_n17539_, new_n17540_, new_n17541_,
    new_n17542_, new_n17543_, new_n17544_, new_n17545_, new_n17546_,
    new_n17547_, new_n17548_, new_n17549_, new_n17550_, new_n17551_,
    new_n17552_, new_n17553_, new_n17554_, new_n17555_, new_n17556_,
    new_n17557_, new_n17558_, new_n17559_, new_n17560_, new_n17561_,
    new_n17562_, new_n17563_, new_n17564_, new_n17565_, new_n17566_,
    new_n17567_, new_n17568_, new_n17569_, new_n17570_, new_n17571_,
    new_n17572_, new_n17573_, new_n17574_, new_n17575_, new_n17576_,
    new_n17577_, new_n17578_, new_n17579_, new_n17580_, new_n17581_,
    new_n17582_, new_n17583_, new_n17584_, new_n17585_, new_n17586_,
    new_n17587_, new_n17588_, new_n17589_, new_n17590_, new_n17591_,
    new_n17592_, new_n17593_, new_n17594_, new_n17595_, new_n17596_,
    new_n17597_, new_n17598_, new_n17599_, new_n17600_, new_n17601_,
    new_n17602_, new_n17603_, new_n17604_, new_n17605_, new_n17606_,
    new_n17607_, new_n17608_, new_n17609_, new_n17610_, new_n17611_,
    new_n17612_, new_n17613_, new_n17614_, new_n17615_, new_n17616_,
    new_n17617_, new_n17618_, new_n17619_, new_n17620_, new_n17621_,
    new_n17622_, new_n17623_, new_n17624_, new_n17625_, new_n17626_,
    new_n17627_, new_n17628_, new_n17629_, new_n17630_, new_n17631_,
    new_n17632_, new_n17633_, new_n17634_, new_n17635_, new_n17636_,
    new_n17637_, new_n17638_, new_n17639_, new_n17640_, new_n17641_,
    new_n17642_, new_n17643_, new_n17644_, new_n17645_, new_n17648_,
    new_n17649_, new_n17650_, new_n17651_, new_n17652_, new_n17653_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17663_,
    new_n17664_, new_n17665_, new_n17666_, new_n17667_, new_n17668_,
    new_n17669_, new_n17670_, new_n17671_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17691_, new_n17692_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17700_, new_n17701_, new_n17702_, new_n17703_,
    new_n17704_, new_n17705_, new_n17706_, new_n17707_, new_n17708_,
    new_n17709_, new_n17710_, new_n17711_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17729_, new_n17730_, new_n17731_, new_n17732_, new_n17733_,
    new_n17734_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17741_, new_n17742_, new_n17743_,
    new_n17744_, new_n17745_, new_n17746_, new_n17747_, new_n17748_,
    new_n17749_, new_n17750_, new_n17751_, new_n17752_, new_n17753_,
    new_n17754_, new_n17755_, new_n17756_, new_n17757_, new_n17758_,
    new_n17759_, new_n17760_, new_n17761_, new_n17762_, new_n17763_,
    new_n17764_, new_n17765_, new_n17766_, new_n17767_, new_n17768_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17802_, new_n17803_,
    new_n17804_, new_n17805_, new_n17806_, new_n17807_, new_n17808_,
    new_n17809_, new_n17810_, new_n17811_, new_n17812_, new_n17813_,
    new_n17814_, new_n17815_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17834_, new_n17835_, new_n17836_, new_n17837_, new_n17838_,
    new_n17839_, new_n17840_, new_n17841_, new_n17842_, new_n17843_,
    new_n17844_, new_n17845_, new_n17846_, new_n17847_, new_n17848_,
    new_n17849_, new_n17850_, new_n17851_, new_n17852_, new_n17853_,
    new_n17854_, new_n17855_, new_n17856_, new_n17857_, new_n17858_,
    new_n17859_, new_n17860_, new_n17861_, new_n17862_, new_n17863_,
    new_n17864_, new_n17865_, new_n17866_, new_n17867_, new_n17868_,
    new_n17869_, new_n17870_, new_n17871_, new_n17872_, new_n17873_,
    new_n17874_, new_n17875_, new_n17876_, new_n17877_, new_n17878_,
    new_n17879_, new_n17880_, new_n17881_, new_n17882_, new_n17883_,
    new_n17884_, new_n17885_, new_n17886_, new_n17887_, new_n17888_,
    new_n17889_, new_n17890_, new_n17891_, new_n17892_, new_n17893_,
    new_n17894_, new_n17895_, new_n17896_, new_n17897_, new_n17898_,
    new_n17899_, new_n17900_, new_n17901_, new_n17902_, new_n17903_,
    new_n17904_, new_n17905_, new_n17906_, new_n17907_, new_n17908_,
    new_n17909_, new_n17910_, new_n17911_, new_n17912_, new_n17913_,
    new_n17914_, new_n17915_, new_n17916_, new_n17917_, new_n17918_,
    new_n17919_, new_n17920_, new_n17921_, new_n17922_, new_n17923_,
    new_n17924_, new_n17925_, new_n17926_, new_n17927_, new_n17928_,
    new_n17929_, new_n17930_, new_n17931_, new_n17932_, new_n17933_,
    new_n17934_, new_n17935_, new_n17936_, new_n17937_, new_n17938_,
    new_n17939_, new_n17940_, new_n17941_, new_n17942_, new_n17943_,
    new_n17944_, new_n17945_, new_n17946_, new_n17947_, new_n17948_,
    new_n17949_, new_n17950_, new_n17951_, new_n17952_, new_n17953_,
    new_n17954_, new_n17955_, new_n17956_, new_n17957_, new_n17958_,
    new_n17959_, new_n17960_, new_n17961_, new_n17962_, new_n17963_,
    new_n17964_, new_n17965_, new_n17966_, new_n17967_, new_n17968_,
    new_n17969_, new_n17970_, new_n17971_, new_n17972_, new_n17973_,
    new_n17974_, new_n17975_, new_n17976_, new_n17977_, new_n17978_,
    new_n17979_, new_n17980_, new_n17981_, new_n17982_, new_n17983_,
    new_n17984_, new_n17985_, new_n17986_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17993_,
    new_n17994_, new_n17995_, new_n17996_, new_n17997_, new_n17998_,
    new_n17999_, new_n18000_, new_n18001_, new_n18002_, new_n18003_,
    new_n18004_, new_n18005_, new_n18006_, new_n18007_, new_n18008_,
    new_n18009_, new_n18010_, new_n18011_, new_n18012_, new_n18013_,
    new_n18014_, new_n18015_, new_n18016_, new_n18017_, new_n18018_,
    new_n18019_, new_n18020_, new_n18021_, new_n18022_, new_n18023_,
    new_n18024_, new_n18025_, new_n18026_, new_n18027_, new_n18028_,
    new_n18029_, new_n18030_, new_n18031_, new_n18032_, new_n18033_,
    new_n18034_, new_n18035_, new_n18036_, new_n18037_, new_n18038_,
    new_n18039_, new_n18040_, new_n18041_, new_n18042_, new_n18043_,
    new_n18044_, new_n18045_, new_n18046_, new_n18047_, new_n18048_,
    new_n18049_, new_n18050_, new_n18051_;
  INV_X1     g00000(.I(\A[334] ), .ZN(new_n1003_));
  NOR2_X1    g00001(.A1(\A[335] ), .A2(\A[336] ), .ZN(new_n1004_));
  NAND2_X1   g00002(.A1(\A[335] ), .A2(\A[336] ), .ZN(new_n1005_));
  AOI21_X1   g00003(.A1(new_n1003_), .A2(new_n1005_), .B(new_n1004_), .ZN(new_n1006_));
  INV_X1     g00004(.I(new_n1006_), .ZN(new_n1007_));
  INV_X1     g00005(.I(\A[331] ), .ZN(new_n1008_));
  NOR2_X1    g00006(.A1(\A[332] ), .A2(\A[333] ), .ZN(new_n1009_));
  NAND2_X1   g00007(.A1(\A[332] ), .A2(\A[333] ), .ZN(new_n1010_));
  AOI21_X1   g00008(.A1(new_n1008_), .A2(new_n1010_), .B(new_n1009_), .ZN(new_n1011_));
  INV_X1     g00009(.I(\A[333] ), .ZN(new_n1012_));
  NOR2_X1    g00010(.A1(new_n1012_), .A2(\A[332] ), .ZN(new_n1013_));
  INV_X1     g00011(.I(\A[332] ), .ZN(new_n1014_));
  NOR2_X1    g00012(.A1(new_n1014_), .A2(\A[333] ), .ZN(new_n1015_));
  OAI21_X1   g00013(.A1(new_n1013_), .A2(new_n1015_), .B(\A[331] ), .ZN(new_n1016_));
  INV_X1     g00014(.I(new_n1010_), .ZN(new_n1017_));
  OAI21_X1   g00015(.A1(new_n1017_), .A2(new_n1009_), .B(new_n1008_), .ZN(new_n1018_));
  NAND2_X1   g00016(.A1(new_n1016_), .A2(new_n1018_), .ZN(new_n1019_));
  INV_X1     g00017(.I(\A[336] ), .ZN(new_n1020_));
  NOR2_X1    g00018(.A1(new_n1020_), .A2(\A[335] ), .ZN(new_n1021_));
  INV_X1     g00019(.I(\A[335] ), .ZN(new_n1022_));
  NOR2_X1    g00020(.A1(new_n1022_), .A2(\A[336] ), .ZN(new_n1023_));
  OAI21_X1   g00021(.A1(new_n1021_), .A2(new_n1023_), .B(\A[334] ), .ZN(new_n1024_));
  AND2_X2    g00022(.A1(\A[335] ), .A2(\A[336] ), .Z(new_n1025_));
  OAI21_X1   g00023(.A1(new_n1025_), .A2(new_n1004_), .B(new_n1003_), .ZN(new_n1026_));
  NAND2_X1   g00024(.A1(new_n1024_), .A2(new_n1026_), .ZN(new_n1027_));
  OAI21_X1   g00025(.A1(new_n1019_), .A2(new_n1027_), .B(new_n1011_), .ZN(new_n1028_));
  INV_X1     g00026(.I(new_n1011_), .ZN(new_n1029_));
  NAND2_X1   g00027(.A1(new_n1014_), .A2(\A[333] ), .ZN(new_n1030_));
  NAND2_X1   g00028(.A1(new_n1012_), .A2(\A[332] ), .ZN(new_n1031_));
  AOI21_X1   g00029(.A1(new_n1030_), .A2(new_n1031_), .B(new_n1008_), .ZN(new_n1032_));
  INV_X1     g00030(.I(new_n1009_), .ZN(new_n1033_));
  AOI21_X1   g00031(.A1(new_n1033_), .A2(new_n1010_), .B(\A[331] ), .ZN(new_n1034_));
  NOR2_X1    g00032(.A1(new_n1034_), .A2(new_n1032_), .ZN(new_n1035_));
  NAND2_X1   g00033(.A1(new_n1022_), .A2(\A[336] ), .ZN(new_n1036_));
  NAND2_X1   g00034(.A1(new_n1020_), .A2(\A[335] ), .ZN(new_n1037_));
  AOI21_X1   g00035(.A1(new_n1036_), .A2(new_n1037_), .B(new_n1003_), .ZN(new_n1038_));
  OR2_X2     g00036(.A1(\A[335] ), .A2(\A[336] ), .Z(new_n1039_));
  AOI21_X1   g00037(.A1(new_n1039_), .A2(new_n1005_), .B(\A[334] ), .ZN(new_n1040_));
  NOR2_X1    g00038(.A1(new_n1038_), .A2(new_n1040_), .ZN(new_n1041_));
  NAND3_X1   g00039(.A1(new_n1035_), .A2(new_n1041_), .A3(new_n1029_), .ZN(new_n1042_));
  AOI21_X1   g00040(.A1(new_n1028_), .A2(new_n1042_), .B(new_n1007_), .ZN(new_n1043_));
  AOI21_X1   g00041(.A1(new_n1035_), .A2(new_n1041_), .B(new_n1029_), .ZN(new_n1044_));
  NOR3_X1    g00042(.A1(new_n1019_), .A2(new_n1027_), .A3(new_n1011_), .ZN(new_n1045_));
  NOR3_X1    g00043(.A1(new_n1044_), .A2(new_n1045_), .A3(new_n1006_), .ZN(new_n1046_));
  NOR2_X1    g00044(.A1(new_n1043_), .A2(new_n1046_), .ZN(new_n1047_));
  INV_X1     g00045(.I(\A[340] ), .ZN(new_n1048_));
  NOR2_X1    g00046(.A1(\A[341] ), .A2(\A[342] ), .ZN(new_n1049_));
  NAND2_X1   g00047(.A1(\A[341] ), .A2(\A[342] ), .ZN(new_n1050_));
  AOI21_X1   g00048(.A1(new_n1048_), .A2(new_n1050_), .B(new_n1049_), .ZN(new_n1051_));
  INV_X1     g00049(.I(\A[337] ), .ZN(new_n1052_));
  NOR2_X1    g00050(.A1(\A[338] ), .A2(\A[339] ), .ZN(new_n1053_));
  NAND2_X1   g00051(.A1(\A[338] ), .A2(\A[339] ), .ZN(new_n1054_));
  AOI21_X1   g00052(.A1(new_n1052_), .A2(new_n1054_), .B(new_n1053_), .ZN(new_n1055_));
  INV_X1     g00053(.I(new_n1055_), .ZN(new_n1056_));
  INV_X1     g00054(.I(\A[341] ), .ZN(new_n1057_));
  NAND2_X1   g00055(.A1(new_n1057_), .A2(\A[342] ), .ZN(new_n1058_));
  INV_X1     g00056(.I(\A[342] ), .ZN(new_n1059_));
  NAND2_X1   g00057(.A1(new_n1059_), .A2(\A[341] ), .ZN(new_n1060_));
  AOI21_X1   g00058(.A1(new_n1058_), .A2(new_n1060_), .B(new_n1048_), .ZN(new_n1061_));
  INV_X1     g00059(.I(new_n1049_), .ZN(new_n1062_));
  AOI21_X1   g00060(.A1(new_n1062_), .A2(new_n1050_), .B(\A[340] ), .ZN(new_n1063_));
  NOR2_X1    g00061(.A1(new_n1063_), .A2(new_n1061_), .ZN(new_n1064_));
  INV_X1     g00062(.I(\A[338] ), .ZN(new_n1065_));
  NAND2_X1   g00063(.A1(new_n1065_), .A2(\A[339] ), .ZN(new_n1066_));
  INV_X1     g00064(.I(\A[339] ), .ZN(new_n1067_));
  NAND2_X1   g00065(.A1(new_n1067_), .A2(\A[338] ), .ZN(new_n1068_));
  AOI21_X1   g00066(.A1(new_n1066_), .A2(new_n1068_), .B(new_n1052_), .ZN(new_n1069_));
  INV_X1     g00067(.I(new_n1053_), .ZN(new_n1070_));
  AOI21_X1   g00068(.A1(new_n1070_), .A2(new_n1054_), .B(\A[337] ), .ZN(new_n1071_));
  NOR2_X1    g00069(.A1(new_n1071_), .A2(new_n1069_), .ZN(new_n1072_));
  AOI21_X1   g00070(.A1(new_n1064_), .A2(new_n1072_), .B(new_n1056_), .ZN(new_n1073_));
  NOR2_X1    g00071(.A1(new_n1059_), .A2(\A[341] ), .ZN(new_n1074_));
  NOR2_X1    g00072(.A1(new_n1057_), .A2(\A[342] ), .ZN(new_n1075_));
  OAI21_X1   g00073(.A1(new_n1074_), .A2(new_n1075_), .B(\A[340] ), .ZN(new_n1076_));
  INV_X1     g00074(.I(new_n1050_), .ZN(new_n1077_));
  OAI21_X1   g00075(.A1(new_n1077_), .A2(new_n1049_), .B(new_n1048_), .ZN(new_n1078_));
  NOR2_X1    g00076(.A1(new_n1067_), .A2(\A[338] ), .ZN(new_n1079_));
  NOR2_X1    g00077(.A1(new_n1065_), .A2(\A[339] ), .ZN(new_n1080_));
  OAI21_X1   g00078(.A1(new_n1079_), .A2(new_n1080_), .B(\A[337] ), .ZN(new_n1081_));
  AND2_X2    g00079(.A1(\A[338] ), .A2(\A[339] ), .Z(new_n1082_));
  OAI21_X1   g00080(.A1(new_n1082_), .A2(new_n1053_), .B(new_n1052_), .ZN(new_n1083_));
  NAND4_X1   g00081(.A1(new_n1076_), .A2(new_n1081_), .A3(new_n1078_), .A4(new_n1083_), .ZN(new_n1084_));
  NOR2_X1    g00082(.A1(new_n1084_), .A2(new_n1055_), .ZN(new_n1085_));
  OAI21_X1   g00083(.A1(new_n1085_), .A2(new_n1073_), .B(new_n1051_), .ZN(new_n1086_));
  INV_X1     g00084(.I(new_n1051_), .ZN(new_n1087_));
  NAND2_X1   g00085(.A1(new_n1084_), .A2(new_n1055_), .ZN(new_n1088_));
  NAND3_X1   g00086(.A1(new_n1064_), .A2(new_n1072_), .A3(new_n1056_), .ZN(new_n1089_));
  NAND3_X1   g00087(.A1(new_n1088_), .A2(new_n1089_), .A3(new_n1087_), .ZN(new_n1090_));
  NAND2_X1   g00088(.A1(new_n1086_), .A2(new_n1090_), .ZN(new_n1091_));
  NAND2_X1   g00089(.A1(new_n1035_), .A2(new_n1041_), .ZN(new_n1092_));
  NAND4_X1   g00090(.A1(new_n1035_), .A2(new_n1041_), .A3(new_n1006_), .A4(new_n1011_), .ZN(new_n1093_));
  OAI22_X1   g00091(.A1(new_n1061_), .A2(new_n1063_), .B1(new_n1071_), .B2(new_n1069_), .ZN(new_n1094_));
  NAND2_X1   g00092(.A1(new_n1094_), .A2(new_n1084_), .ZN(new_n1095_));
  NOR2_X1    g00093(.A1(new_n1095_), .A2(new_n1093_), .ZN(new_n1096_));
  NAND2_X1   g00094(.A1(new_n1019_), .A2(new_n1027_), .ZN(new_n1097_));
  NAND2_X1   g00095(.A1(new_n1076_), .A2(new_n1078_), .ZN(new_n1098_));
  NAND2_X1   g00096(.A1(new_n1081_), .A2(new_n1083_), .ZN(new_n1099_));
  NAND2_X1   g00097(.A1(new_n1051_), .A2(new_n1055_), .ZN(new_n1100_));
  NOR3_X1    g00098(.A1(new_n1098_), .A2(new_n1099_), .A3(new_n1100_), .ZN(new_n1101_));
  NAND4_X1   g00099(.A1(new_n1096_), .A2(new_n1092_), .A3(new_n1097_), .A4(new_n1101_), .ZN(new_n1102_));
  NAND2_X1   g00100(.A1(new_n1006_), .A2(new_n1011_), .ZN(new_n1103_));
  NOR3_X1    g00101(.A1(new_n1019_), .A2(new_n1027_), .A3(new_n1103_), .ZN(new_n1104_));
  NAND3_X1   g00102(.A1(new_n1104_), .A2(new_n1084_), .A3(new_n1094_), .ZN(new_n1105_));
  NAND2_X1   g00103(.A1(new_n1092_), .A2(new_n1097_), .ZN(new_n1106_));
  AOI21_X1   g00104(.A1(new_n1098_), .A2(new_n1099_), .B(new_n1100_), .ZN(new_n1107_));
  NOR3_X1    g00105(.A1(new_n1105_), .A2(new_n1106_), .A3(new_n1107_), .ZN(new_n1108_));
  OAI21_X1   g00106(.A1(new_n1102_), .A2(new_n1091_), .B(new_n1047_), .ZN(new_n1109_));
  NAND3_X1   g00107(.A1(new_n1101_), .A2(new_n1084_), .A3(new_n1094_), .ZN(new_n1110_));
  NOR2_X1    g00108(.A1(new_n1019_), .A2(new_n1027_), .ZN(new_n1111_));
  NOR2_X1    g00109(.A1(new_n1035_), .A2(new_n1041_), .ZN(new_n1112_));
  NOR3_X1    g00110(.A1(new_n1093_), .A2(new_n1111_), .A3(new_n1112_), .ZN(new_n1113_));
  NAND2_X1   g00111(.A1(new_n1113_), .A2(new_n1110_), .ZN(new_n1114_));
  NAND4_X1   g00112(.A1(new_n1064_), .A2(new_n1072_), .A3(new_n1051_), .A4(new_n1055_), .ZN(new_n1115_));
  NOR2_X1    g00113(.A1(new_n1095_), .A2(new_n1115_), .ZN(new_n1116_));
  NAND3_X1   g00114(.A1(new_n1104_), .A2(new_n1092_), .A3(new_n1097_), .ZN(new_n1117_));
  NAND2_X1   g00115(.A1(new_n1116_), .A2(new_n1117_), .ZN(new_n1118_));
  INV_X1     g00116(.I(\A[325] ), .ZN(new_n1119_));
  INV_X1     g00117(.I(\A[326] ), .ZN(new_n1120_));
  NAND2_X1   g00118(.A1(new_n1120_), .A2(\A[327] ), .ZN(new_n1121_));
  INV_X1     g00119(.I(\A[327] ), .ZN(new_n1122_));
  NAND2_X1   g00120(.A1(new_n1122_), .A2(\A[326] ), .ZN(new_n1123_));
  AOI21_X1   g00121(.A1(new_n1121_), .A2(new_n1123_), .B(new_n1119_), .ZN(new_n1124_));
  NAND2_X1   g00122(.A1(\A[326] ), .A2(\A[327] ), .ZN(new_n1125_));
  NOR2_X1    g00123(.A1(\A[326] ), .A2(\A[327] ), .ZN(new_n1126_));
  INV_X1     g00124(.I(new_n1126_), .ZN(new_n1127_));
  AOI21_X1   g00125(.A1(new_n1127_), .A2(new_n1125_), .B(\A[325] ), .ZN(new_n1128_));
  NOR2_X1    g00126(.A1(new_n1128_), .A2(new_n1124_), .ZN(new_n1129_));
  INV_X1     g00127(.I(\A[328] ), .ZN(new_n1130_));
  INV_X1     g00128(.I(\A[329] ), .ZN(new_n1131_));
  NAND2_X1   g00129(.A1(new_n1131_), .A2(\A[330] ), .ZN(new_n1132_));
  INV_X1     g00130(.I(\A[330] ), .ZN(new_n1133_));
  NAND2_X1   g00131(.A1(new_n1133_), .A2(\A[329] ), .ZN(new_n1134_));
  AOI21_X1   g00132(.A1(new_n1132_), .A2(new_n1134_), .B(new_n1130_), .ZN(new_n1135_));
  NAND2_X1   g00133(.A1(\A[329] ), .A2(\A[330] ), .ZN(new_n1136_));
  NOR2_X1    g00134(.A1(\A[329] ), .A2(\A[330] ), .ZN(new_n1137_));
  INV_X1     g00135(.I(new_n1137_), .ZN(new_n1138_));
  AOI21_X1   g00136(.A1(new_n1138_), .A2(new_n1136_), .B(\A[328] ), .ZN(new_n1139_));
  NOR2_X1    g00137(.A1(new_n1139_), .A2(new_n1135_), .ZN(new_n1140_));
  NOR2_X1    g00138(.A1(new_n1129_), .A2(new_n1140_), .ZN(new_n1141_));
  NOR4_X1    g00139(.A1(new_n1124_), .A2(new_n1128_), .A3(new_n1139_), .A4(new_n1135_), .ZN(new_n1142_));
  NOR2_X1    g00140(.A1(new_n1141_), .A2(new_n1142_), .ZN(new_n1143_));
  NOR2_X1    g00141(.A1(new_n1122_), .A2(\A[326] ), .ZN(new_n1144_));
  NOR2_X1    g00142(.A1(new_n1120_), .A2(\A[327] ), .ZN(new_n1145_));
  OAI21_X1   g00143(.A1(new_n1144_), .A2(new_n1145_), .B(\A[325] ), .ZN(new_n1146_));
  INV_X1     g00144(.I(new_n1125_), .ZN(new_n1147_));
  OAI21_X1   g00145(.A1(new_n1147_), .A2(new_n1126_), .B(new_n1119_), .ZN(new_n1148_));
  NAND2_X1   g00146(.A1(new_n1146_), .A2(new_n1148_), .ZN(new_n1149_));
  NOR2_X1    g00147(.A1(new_n1133_), .A2(\A[329] ), .ZN(new_n1150_));
  NOR2_X1    g00148(.A1(new_n1131_), .A2(\A[330] ), .ZN(new_n1151_));
  OAI21_X1   g00149(.A1(new_n1150_), .A2(new_n1151_), .B(\A[328] ), .ZN(new_n1152_));
  INV_X1     g00150(.I(new_n1136_), .ZN(new_n1153_));
  OAI21_X1   g00151(.A1(new_n1153_), .A2(new_n1137_), .B(new_n1130_), .ZN(new_n1154_));
  NAND2_X1   g00152(.A1(new_n1152_), .A2(new_n1154_), .ZN(new_n1155_));
  AOI21_X1   g00153(.A1(new_n1130_), .A2(new_n1136_), .B(new_n1137_), .ZN(new_n1156_));
  AOI21_X1   g00154(.A1(new_n1119_), .A2(new_n1125_), .B(new_n1126_), .ZN(new_n1157_));
  NAND2_X1   g00155(.A1(new_n1156_), .A2(new_n1157_), .ZN(new_n1158_));
  NOR3_X1    g00156(.A1(new_n1149_), .A2(new_n1155_), .A3(new_n1158_), .ZN(new_n1159_));
  INV_X1     g00157(.I(\A[319] ), .ZN(new_n1160_));
  INV_X1     g00158(.I(\A[320] ), .ZN(new_n1161_));
  NAND2_X1   g00159(.A1(new_n1161_), .A2(\A[321] ), .ZN(new_n1162_));
  INV_X1     g00160(.I(\A[321] ), .ZN(new_n1163_));
  NAND2_X1   g00161(.A1(new_n1163_), .A2(\A[320] ), .ZN(new_n1164_));
  AOI21_X1   g00162(.A1(new_n1162_), .A2(new_n1164_), .B(new_n1160_), .ZN(new_n1165_));
  NOR2_X1    g00163(.A1(\A[320] ), .A2(\A[321] ), .ZN(new_n1166_));
  INV_X1     g00164(.I(new_n1166_), .ZN(new_n1167_));
  NAND2_X1   g00165(.A1(\A[320] ), .A2(\A[321] ), .ZN(new_n1168_));
  AOI21_X1   g00166(.A1(new_n1167_), .A2(new_n1168_), .B(\A[319] ), .ZN(new_n1169_));
  NOR2_X1    g00167(.A1(new_n1169_), .A2(new_n1165_), .ZN(new_n1170_));
  INV_X1     g00168(.I(\A[322] ), .ZN(new_n1171_));
  INV_X1     g00169(.I(\A[323] ), .ZN(new_n1172_));
  NAND2_X1   g00170(.A1(new_n1172_), .A2(\A[324] ), .ZN(new_n1173_));
  INV_X1     g00171(.I(\A[324] ), .ZN(new_n1174_));
  NAND2_X1   g00172(.A1(new_n1174_), .A2(\A[323] ), .ZN(new_n1175_));
  AOI21_X1   g00173(.A1(new_n1173_), .A2(new_n1175_), .B(new_n1171_), .ZN(new_n1176_));
  NOR2_X1    g00174(.A1(\A[323] ), .A2(\A[324] ), .ZN(new_n1177_));
  INV_X1     g00175(.I(new_n1177_), .ZN(new_n1178_));
  NAND2_X1   g00176(.A1(\A[323] ), .A2(\A[324] ), .ZN(new_n1179_));
  AOI21_X1   g00177(.A1(new_n1178_), .A2(new_n1179_), .B(\A[322] ), .ZN(new_n1180_));
  NOR2_X1    g00178(.A1(new_n1180_), .A2(new_n1176_), .ZN(new_n1181_));
  AOI21_X1   g00179(.A1(new_n1171_), .A2(new_n1179_), .B(new_n1177_), .ZN(new_n1182_));
  AOI21_X1   g00180(.A1(new_n1160_), .A2(new_n1168_), .B(new_n1166_), .ZN(new_n1183_));
  NAND2_X1   g00181(.A1(new_n1182_), .A2(new_n1183_), .ZN(new_n1184_));
  NAND2_X1   g00182(.A1(new_n1143_), .A2(new_n1159_), .ZN(new_n1186_));
  AOI21_X1   g00183(.A1(new_n1118_), .A2(new_n1114_), .B(new_n1186_), .ZN(new_n1187_));
  NOR2_X1    g00184(.A1(new_n1109_), .A2(new_n1187_), .ZN(new_n1188_));
  OAI21_X1   g00185(.A1(new_n1044_), .A2(new_n1045_), .B(new_n1006_), .ZN(new_n1189_));
  NAND3_X1   g00186(.A1(new_n1028_), .A2(new_n1042_), .A3(new_n1007_), .ZN(new_n1190_));
  NAND2_X1   g00187(.A1(new_n1189_), .A2(new_n1190_), .ZN(new_n1191_));
  AOI21_X1   g00188(.A1(new_n1088_), .A2(new_n1089_), .B(new_n1087_), .ZN(new_n1192_));
  NOR3_X1    g00189(.A1(new_n1085_), .A2(new_n1073_), .A3(new_n1051_), .ZN(new_n1193_));
  NOR2_X1    g00190(.A1(new_n1193_), .A2(new_n1192_), .ZN(new_n1194_));
  NOR3_X1    g00191(.A1(new_n1105_), .A2(new_n1106_), .A3(new_n1115_), .ZN(new_n1195_));
  AOI21_X1   g00192(.A1(new_n1194_), .A2(new_n1195_), .B(new_n1191_), .ZN(new_n1196_));
  NOR2_X1    g00193(.A1(new_n1116_), .A2(new_n1117_), .ZN(new_n1197_));
  NOR2_X1    g00194(.A1(new_n1113_), .A2(new_n1110_), .ZN(new_n1198_));
  NAND2_X1   g00195(.A1(new_n1149_), .A2(new_n1155_), .ZN(new_n1199_));
  INV_X1     g00196(.I(new_n1142_), .ZN(new_n1200_));
  NAND2_X1   g00197(.A1(new_n1200_), .A2(new_n1199_), .ZN(new_n1201_));
  INV_X1     g00198(.I(new_n1159_), .ZN(new_n1202_));
  NOR2_X1    g00199(.A1(new_n1201_), .A2(new_n1202_), .ZN(new_n1203_));
  OAI21_X1   g00200(.A1(new_n1197_), .A2(new_n1198_), .B(new_n1203_), .ZN(new_n1204_));
  NOR2_X1    g00201(.A1(new_n1196_), .A2(new_n1204_), .ZN(new_n1205_));
  NOR2_X1    g00202(.A1(new_n1188_), .A2(new_n1205_), .ZN(new_n1206_));
  NAND2_X1   g00203(.A1(new_n1109_), .A2(new_n1187_), .ZN(new_n1207_));
  INV_X1     g00204(.I(new_n1156_), .ZN(new_n1208_));
  OAI21_X1   g00205(.A1(new_n1149_), .A2(new_n1155_), .B(new_n1157_), .ZN(new_n1209_));
  INV_X1     g00206(.I(new_n1157_), .ZN(new_n1210_));
  NAND3_X1   g00207(.A1(new_n1129_), .A2(new_n1140_), .A3(new_n1210_), .ZN(new_n1211_));
  AOI21_X1   g00208(.A1(new_n1209_), .A2(new_n1211_), .B(new_n1208_), .ZN(new_n1212_));
  NOR2_X1    g00209(.A1(new_n1142_), .A2(new_n1210_), .ZN(new_n1213_));
  NOR3_X1    g00210(.A1(new_n1149_), .A2(new_n1155_), .A3(new_n1157_), .ZN(new_n1214_));
  NOR3_X1    g00211(.A1(new_n1213_), .A2(new_n1214_), .A3(new_n1156_), .ZN(new_n1215_));
  NOR2_X1    g00212(.A1(new_n1163_), .A2(\A[320] ), .ZN(new_n1216_));
  NOR2_X1    g00213(.A1(new_n1161_), .A2(\A[321] ), .ZN(new_n1217_));
  OAI21_X1   g00214(.A1(new_n1216_), .A2(new_n1217_), .B(\A[319] ), .ZN(new_n1218_));
  INV_X1     g00215(.I(new_n1168_), .ZN(new_n1219_));
  OAI21_X1   g00216(.A1(new_n1219_), .A2(new_n1166_), .B(new_n1160_), .ZN(new_n1220_));
  NAND2_X1   g00217(.A1(new_n1218_), .A2(new_n1220_), .ZN(new_n1221_));
  NOR2_X1    g00218(.A1(new_n1174_), .A2(\A[323] ), .ZN(new_n1222_));
  NOR2_X1    g00219(.A1(new_n1172_), .A2(\A[324] ), .ZN(new_n1223_));
  OAI21_X1   g00220(.A1(new_n1222_), .A2(new_n1223_), .B(\A[322] ), .ZN(new_n1224_));
  INV_X1     g00221(.I(new_n1179_), .ZN(new_n1225_));
  OAI21_X1   g00222(.A1(new_n1225_), .A2(new_n1177_), .B(new_n1171_), .ZN(new_n1226_));
  NAND2_X1   g00223(.A1(new_n1224_), .A2(new_n1226_), .ZN(new_n1227_));
  NOR3_X1    g00224(.A1(new_n1221_), .A2(new_n1227_), .A3(new_n1184_), .ZN(new_n1228_));
  NOR4_X1    g00225(.A1(new_n1165_), .A2(new_n1169_), .A3(new_n1180_), .A4(new_n1176_), .ZN(new_n1229_));
  NOR2_X1    g00226(.A1(new_n1170_), .A2(new_n1181_), .ZN(new_n1230_));
  NOR2_X1    g00227(.A1(new_n1230_), .A2(new_n1229_), .ZN(new_n1231_));
  INV_X1     g00228(.I(new_n1158_), .ZN(new_n1232_));
  NAND2_X1   g00229(.A1(new_n1208_), .A2(new_n1210_), .ZN(new_n1233_));
  AOI21_X1   g00230(.A1(new_n1142_), .A2(new_n1233_), .B(new_n1232_), .ZN(new_n1234_));
  NAND4_X1   g00231(.A1(new_n1143_), .A2(new_n1231_), .A3(new_n1234_), .A4(new_n1228_), .ZN(new_n1235_));
  NOR3_X1    g00232(.A1(new_n1235_), .A2(new_n1212_), .A3(new_n1215_), .ZN(new_n1236_));
  INV_X1     g00233(.I(new_n1183_), .ZN(new_n1237_));
  NOR2_X1    g00234(.A1(new_n1229_), .A2(new_n1237_), .ZN(new_n1238_));
  NOR3_X1    g00235(.A1(new_n1221_), .A2(new_n1227_), .A3(new_n1183_), .ZN(new_n1239_));
  OAI21_X1   g00236(.A1(new_n1238_), .A2(new_n1239_), .B(new_n1182_), .ZN(new_n1240_));
  INV_X1     g00237(.I(new_n1182_), .ZN(new_n1241_));
  OAI21_X1   g00238(.A1(new_n1221_), .A2(new_n1227_), .B(new_n1183_), .ZN(new_n1242_));
  NAND3_X1   g00239(.A1(new_n1170_), .A2(new_n1181_), .A3(new_n1237_), .ZN(new_n1243_));
  NAND3_X1   g00240(.A1(new_n1242_), .A2(new_n1243_), .A3(new_n1241_), .ZN(new_n1244_));
  NAND2_X1   g00241(.A1(new_n1240_), .A2(new_n1244_), .ZN(new_n1245_));
  NAND2_X1   g00242(.A1(new_n1236_), .A2(new_n1245_), .ZN(new_n1246_));
  NAND4_X1   g00243(.A1(new_n1143_), .A2(new_n1231_), .A3(new_n1159_), .A4(new_n1228_), .ZN(new_n1247_));
  NAND2_X1   g00244(.A1(new_n1245_), .A2(new_n1247_), .ZN(new_n1248_));
  NOR2_X1    g00245(.A1(new_n1215_), .A2(new_n1212_), .ZN(new_n1249_));
  NAND4_X1   g00246(.A1(new_n1200_), .A2(new_n1199_), .A3(new_n1156_), .A4(new_n1157_), .ZN(new_n1250_));
  AOI21_X1   g00247(.A1(new_n1242_), .A2(new_n1243_), .B(new_n1241_), .ZN(new_n1251_));
  NOR3_X1    g00248(.A1(new_n1238_), .A2(new_n1239_), .A3(new_n1182_), .ZN(new_n1252_));
  NOR2_X1    g00249(.A1(new_n1252_), .A2(new_n1251_), .ZN(new_n1253_));
  NAND3_X1   g00250(.A1(new_n1200_), .A2(new_n1159_), .A3(new_n1199_), .ZN(new_n1254_));
  INV_X1     g00251(.I(new_n1228_), .ZN(new_n1255_));
  INV_X1     g00252(.I(new_n1229_), .ZN(new_n1256_));
  NAND2_X1   g00253(.A1(new_n1221_), .A2(new_n1227_), .ZN(new_n1257_));
  NAND2_X1   g00254(.A1(new_n1256_), .A2(new_n1257_), .ZN(new_n1258_));
  NOR3_X1    g00255(.A1(new_n1254_), .A2(new_n1255_), .A3(new_n1258_), .ZN(new_n1259_));
  AOI22_X1   g00256(.A1(new_n1253_), .A2(new_n1259_), .B1(new_n1249_), .B2(new_n1250_), .ZN(new_n1260_));
  OAI21_X1   g00257(.A1(new_n1213_), .A2(new_n1214_), .B(new_n1156_), .ZN(new_n1261_));
  NAND3_X1   g00258(.A1(new_n1209_), .A2(new_n1211_), .A3(new_n1208_), .ZN(new_n1262_));
  NAND3_X1   g00259(.A1(new_n1261_), .A2(new_n1250_), .A3(new_n1262_), .ZN(new_n1263_));
  NOR3_X1    g00260(.A1(new_n1263_), .A2(new_n1245_), .A3(new_n1247_), .ZN(new_n1264_));
  OAI21_X1   g00261(.A1(new_n1260_), .A2(new_n1264_), .B(new_n1248_), .ZN(new_n1265_));
  NAND2_X1   g00262(.A1(new_n1265_), .A2(new_n1246_), .ZN(new_n1266_));
  OAI21_X1   g00263(.A1(new_n1266_), .A2(new_n1206_), .B(new_n1207_), .ZN(new_n1267_));
  NOR4_X1    g00264(.A1(new_n1091_), .A2(new_n1105_), .A3(new_n1106_), .A4(new_n1107_), .ZN(new_n1268_));
  AOI21_X1   g00265(.A1(new_n1194_), .A2(new_n1195_), .B(new_n1047_), .ZN(new_n1269_));
  NOR2_X1    g00266(.A1(new_n1051_), .A2(new_n1055_), .ZN(new_n1270_));
  OAI21_X1   g00267(.A1(new_n1084_), .A2(new_n1270_), .B(new_n1100_), .ZN(new_n1271_));
  NOR2_X1    g00268(.A1(new_n1006_), .A2(new_n1011_), .ZN(new_n1272_));
  OAI21_X1   g00269(.A1(new_n1092_), .A2(new_n1272_), .B(new_n1103_), .ZN(new_n1273_));
  XOR2_X1    g00270(.A1(new_n1273_), .A2(new_n1271_), .Z(new_n1274_));
  NOR3_X1    g00271(.A1(new_n1269_), .A2(new_n1268_), .A3(new_n1274_), .ZN(new_n1275_));
  INV_X1     g00272(.I(new_n1234_), .ZN(new_n1276_));
  NOR4_X1    g00273(.A1(new_n1276_), .A2(new_n1201_), .A3(new_n1258_), .A4(new_n1255_), .ZN(new_n1277_));
  NAND2_X1   g00274(.A1(new_n1277_), .A2(new_n1249_), .ZN(new_n1278_));
  NOR4_X1    g00275(.A1(new_n1141_), .A2(new_n1142_), .A3(new_n1208_), .A4(new_n1210_), .ZN(new_n1279_));
  NOR3_X1    g00276(.A1(new_n1215_), .A2(new_n1212_), .A3(new_n1279_), .ZN(new_n1280_));
  OAI21_X1   g00277(.A1(new_n1280_), .A2(new_n1247_), .B(new_n1245_), .ZN(new_n1281_));
  NOR3_X1    g00278(.A1(new_n1215_), .A2(new_n1212_), .A3(new_n1201_), .ZN(new_n1282_));
  NOR2_X1    g00279(.A1(new_n1182_), .A2(new_n1183_), .ZN(new_n1283_));
  OAI21_X1   g00280(.A1(new_n1256_), .A2(new_n1283_), .B(new_n1184_), .ZN(new_n1284_));
  INV_X1     g00281(.I(new_n1284_), .ZN(new_n1285_));
  OAI21_X1   g00282(.A1(new_n1282_), .A2(new_n1234_), .B(new_n1285_), .ZN(new_n1286_));
  NAND3_X1   g00283(.A1(new_n1261_), .A2(new_n1262_), .A3(new_n1143_), .ZN(new_n1287_));
  NAND3_X1   g00284(.A1(new_n1287_), .A2(new_n1276_), .A3(new_n1284_), .ZN(new_n1288_));
  NAND4_X1   g00285(.A1(new_n1281_), .A2(new_n1286_), .A3(new_n1288_), .A4(new_n1278_), .ZN(new_n1289_));
  NAND2_X1   g00286(.A1(new_n1289_), .A2(new_n1275_), .ZN(new_n1290_));
  NAND2_X1   g00287(.A1(new_n1194_), .A2(new_n1108_), .ZN(new_n1291_));
  OAI21_X1   g00288(.A1(new_n1102_), .A2(new_n1091_), .B(new_n1191_), .ZN(new_n1292_));
  XNOR2_X1   g00289(.A1(new_n1273_), .A2(new_n1271_), .ZN(new_n1293_));
  NAND3_X1   g00290(.A1(new_n1292_), .A2(new_n1293_), .A3(new_n1291_), .ZN(new_n1294_));
  NAND2_X1   g00291(.A1(new_n1263_), .A2(new_n1259_), .ZN(new_n1295_));
  AOI21_X1   g00292(.A1(new_n1295_), .A2(new_n1245_), .B(new_n1236_), .ZN(new_n1296_));
  AOI21_X1   g00293(.A1(new_n1287_), .A2(new_n1276_), .B(new_n1284_), .ZN(new_n1297_));
  NOR3_X1    g00294(.A1(new_n1282_), .A2(new_n1234_), .A3(new_n1285_), .ZN(new_n1298_));
  NOR2_X1    g00295(.A1(new_n1298_), .A2(new_n1297_), .ZN(new_n1299_));
  NAND3_X1   g00296(.A1(new_n1296_), .A2(new_n1299_), .A3(new_n1294_), .ZN(new_n1300_));
  NAND2_X1   g00297(.A1(new_n1290_), .A2(new_n1300_), .ZN(new_n1301_));
  NAND2_X1   g00298(.A1(new_n1301_), .A2(new_n1267_), .ZN(new_n1302_));
  NAND2_X1   g00299(.A1(new_n1196_), .A2(new_n1204_), .ZN(new_n1303_));
  NAND2_X1   g00300(.A1(new_n1109_), .A2(new_n1187_), .ZN(new_n1304_));
  NAND2_X1   g00301(.A1(new_n1304_), .A2(new_n1303_), .ZN(new_n1305_));
  NOR2_X1    g00302(.A1(new_n1278_), .A2(new_n1253_), .ZN(new_n1306_));
  OAI21_X1   g00303(.A1(new_n1245_), .A2(new_n1247_), .B(new_n1263_), .ZN(new_n1307_));
  NAND3_X1   g00304(.A1(new_n1280_), .A2(new_n1253_), .A3(new_n1259_), .ZN(new_n1308_));
  NAND2_X1   g00305(.A1(new_n1307_), .A2(new_n1308_), .ZN(new_n1309_));
  AOI21_X1   g00306(.A1(new_n1309_), .A2(new_n1248_), .B(new_n1306_), .ZN(new_n1310_));
  OAI21_X1   g00307(.A1(new_n1310_), .A2(new_n1109_), .B(new_n1305_), .ZN(new_n1311_));
  NAND2_X1   g00308(.A1(new_n1289_), .A2(new_n1294_), .ZN(new_n1312_));
  NAND3_X1   g00309(.A1(new_n1275_), .A2(new_n1299_), .A3(new_n1296_), .ZN(new_n1313_));
  NAND2_X1   g00310(.A1(new_n1313_), .A2(new_n1312_), .ZN(new_n1314_));
  NAND2_X1   g00311(.A1(new_n1314_), .A2(new_n1311_), .ZN(new_n1315_));
  NAND2_X1   g00312(.A1(new_n1302_), .A2(new_n1315_), .ZN(new_n1316_));
  INV_X1     g00313(.I(\A[364] ), .ZN(new_n1317_));
  NOR2_X1    g00314(.A1(\A[365] ), .A2(\A[366] ), .ZN(new_n1318_));
  NAND2_X1   g00315(.A1(\A[365] ), .A2(\A[366] ), .ZN(new_n1319_));
  AOI21_X1   g00316(.A1(new_n1317_), .A2(new_n1319_), .B(new_n1318_), .ZN(new_n1320_));
  INV_X1     g00317(.I(new_n1320_), .ZN(new_n1321_));
  INV_X1     g00318(.I(\A[361] ), .ZN(new_n1322_));
  NOR2_X1    g00319(.A1(\A[362] ), .A2(\A[363] ), .ZN(new_n1323_));
  NAND2_X1   g00320(.A1(\A[362] ), .A2(\A[363] ), .ZN(new_n1324_));
  AOI21_X1   g00321(.A1(new_n1322_), .A2(new_n1324_), .B(new_n1323_), .ZN(new_n1325_));
  INV_X1     g00322(.I(\A[363] ), .ZN(new_n1326_));
  NOR2_X1    g00323(.A1(new_n1326_), .A2(\A[362] ), .ZN(new_n1327_));
  INV_X1     g00324(.I(\A[362] ), .ZN(new_n1328_));
  NOR2_X1    g00325(.A1(new_n1328_), .A2(\A[363] ), .ZN(new_n1329_));
  OAI21_X1   g00326(.A1(new_n1327_), .A2(new_n1329_), .B(\A[361] ), .ZN(new_n1330_));
  INV_X1     g00327(.I(new_n1324_), .ZN(new_n1331_));
  OAI21_X1   g00328(.A1(new_n1331_), .A2(new_n1323_), .B(new_n1322_), .ZN(new_n1332_));
  NAND2_X1   g00329(.A1(new_n1330_), .A2(new_n1332_), .ZN(new_n1333_));
  INV_X1     g00330(.I(\A[366] ), .ZN(new_n1334_));
  NOR2_X1    g00331(.A1(new_n1334_), .A2(\A[365] ), .ZN(new_n1335_));
  INV_X1     g00332(.I(\A[365] ), .ZN(new_n1336_));
  NOR2_X1    g00333(.A1(new_n1336_), .A2(\A[366] ), .ZN(new_n1337_));
  OAI21_X1   g00334(.A1(new_n1335_), .A2(new_n1337_), .B(\A[364] ), .ZN(new_n1338_));
  AND2_X2    g00335(.A1(\A[365] ), .A2(\A[366] ), .Z(new_n1339_));
  OAI21_X1   g00336(.A1(new_n1339_), .A2(new_n1318_), .B(new_n1317_), .ZN(new_n1340_));
  NAND2_X1   g00337(.A1(new_n1338_), .A2(new_n1340_), .ZN(new_n1341_));
  OAI21_X1   g00338(.A1(new_n1333_), .A2(new_n1341_), .B(new_n1325_), .ZN(new_n1342_));
  INV_X1     g00339(.I(new_n1325_), .ZN(new_n1343_));
  NAND2_X1   g00340(.A1(new_n1328_), .A2(\A[363] ), .ZN(new_n1344_));
  NAND2_X1   g00341(.A1(new_n1326_), .A2(\A[362] ), .ZN(new_n1345_));
  AOI21_X1   g00342(.A1(new_n1344_), .A2(new_n1345_), .B(new_n1322_), .ZN(new_n1346_));
  INV_X1     g00343(.I(new_n1323_), .ZN(new_n1347_));
  AOI21_X1   g00344(.A1(new_n1347_), .A2(new_n1324_), .B(\A[361] ), .ZN(new_n1348_));
  NOR2_X1    g00345(.A1(new_n1348_), .A2(new_n1346_), .ZN(new_n1349_));
  NAND2_X1   g00346(.A1(new_n1336_), .A2(\A[366] ), .ZN(new_n1350_));
  NAND2_X1   g00347(.A1(new_n1334_), .A2(\A[365] ), .ZN(new_n1351_));
  AOI21_X1   g00348(.A1(new_n1350_), .A2(new_n1351_), .B(new_n1317_), .ZN(new_n1352_));
  INV_X1     g00349(.I(new_n1318_), .ZN(new_n1353_));
  AOI21_X1   g00350(.A1(new_n1353_), .A2(new_n1319_), .B(\A[364] ), .ZN(new_n1354_));
  NOR2_X1    g00351(.A1(new_n1354_), .A2(new_n1352_), .ZN(new_n1355_));
  NAND3_X1   g00352(.A1(new_n1349_), .A2(new_n1355_), .A3(new_n1343_), .ZN(new_n1356_));
  AOI21_X1   g00353(.A1(new_n1356_), .A2(new_n1342_), .B(new_n1321_), .ZN(new_n1357_));
  AOI21_X1   g00354(.A1(new_n1349_), .A2(new_n1355_), .B(new_n1343_), .ZN(new_n1358_));
  NOR3_X1    g00355(.A1(new_n1333_), .A2(new_n1341_), .A3(new_n1325_), .ZN(new_n1359_));
  NOR3_X1    g00356(.A1(new_n1358_), .A2(new_n1359_), .A3(new_n1320_), .ZN(new_n1360_));
  INV_X1     g00357(.I(\A[357] ), .ZN(new_n1361_));
  NOR2_X1    g00358(.A1(new_n1361_), .A2(\A[356] ), .ZN(new_n1362_));
  INV_X1     g00359(.I(\A[356] ), .ZN(new_n1363_));
  NOR2_X1    g00360(.A1(new_n1363_), .A2(\A[357] ), .ZN(new_n1364_));
  OAI21_X1   g00361(.A1(new_n1362_), .A2(new_n1364_), .B(\A[355] ), .ZN(new_n1365_));
  INV_X1     g00362(.I(\A[355] ), .ZN(new_n1366_));
  NOR2_X1    g00363(.A1(\A[356] ), .A2(\A[357] ), .ZN(new_n1367_));
  NAND2_X1   g00364(.A1(\A[356] ), .A2(\A[357] ), .ZN(new_n1368_));
  INV_X1     g00365(.I(new_n1368_), .ZN(new_n1369_));
  OAI21_X1   g00366(.A1(new_n1369_), .A2(new_n1367_), .B(new_n1366_), .ZN(new_n1370_));
  NAND2_X1   g00367(.A1(new_n1365_), .A2(new_n1370_), .ZN(new_n1371_));
  INV_X1     g00368(.I(\A[358] ), .ZN(new_n1372_));
  INV_X1     g00369(.I(\A[359] ), .ZN(new_n1373_));
  NAND2_X1   g00370(.A1(new_n1373_), .A2(\A[360] ), .ZN(new_n1374_));
  INV_X1     g00371(.I(\A[360] ), .ZN(new_n1375_));
  NAND2_X1   g00372(.A1(new_n1375_), .A2(\A[359] ), .ZN(new_n1376_));
  AOI21_X1   g00373(.A1(new_n1374_), .A2(new_n1376_), .B(new_n1372_), .ZN(new_n1377_));
  NOR2_X1    g00374(.A1(\A[359] ), .A2(\A[360] ), .ZN(new_n1378_));
  INV_X1     g00375(.I(new_n1378_), .ZN(new_n1379_));
  NAND2_X1   g00376(.A1(\A[359] ), .A2(\A[360] ), .ZN(new_n1380_));
  AOI21_X1   g00377(.A1(new_n1379_), .A2(new_n1380_), .B(\A[358] ), .ZN(new_n1381_));
  NOR2_X1    g00378(.A1(new_n1381_), .A2(new_n1377_), .ZN(new_n1382_));
  NOR2_X1    g00379(.A1(new_n1382_), .A2(new_n1371_), .ZN(new_n1383_));
  NAND2_X1   g00380(.A1(new_n1363_), .A2(\A[357] ), .ZN(new_n1384_));
  NAND2_X1   g00381(.A1(new_n1361_), .A2(\A[356] ), .ZN(new_n1385_));
  AOI21_X1   g00382(.A1(new_n1384_), .A2(new_n1385_), .B(new_n1366_), .ZN(new_n1386_));
  INV_X1     g00383(.I(new_n1367_), .ZN(new_n1387_));
  AOI21_X1   g00384(.A1(new_n1387_), .A2(new_n1368_), .B(\A[355] ), .ZN(new_n1388_));
  NOR2_X1    g00385(.A1(new_n1388_), .A2(new_n1386_), .ZN(new_n1389_));
  NOR2_X1    g00386(.A1(new_n1375_), .A2(\A[359] ), .ZN(new_n1390_));
  NOR2_X1    g00387(.A1(new_n1373_), .A2(\A[360] ), .ZN(new_n1391_));
  OAI21_X1   g00388(.A1(new_n1390_), .A2(new_n1391_), .B(\A[358] ), .ZN(new_n1392_));
  INV_X1     g00389(.I(new_n1380_), .ZN(new_n1393_));
  OAI21_X1   g00390(.A1(new_n1393_), .A2(new_n1378_), .B(new_n1372_), .ZN(new_n1394_));
  NAND2_X1   g00391(.A1(new_n1392_), .A2(new_n1394_), .ZN(new_n1395_));
  NOR2_X1    g00392(.A1(new_n1389_), .A2(new_n1395_), .ZN(new_n1396_));
  NOR2_X1    g00393(.A1(new_n1355_), .A2(new_n1333_), .ZN(new_n1397_));
  NOR2_X1    g00394(.A1(new_n1349_), .A2(new_n1341_), .ZN(new_n1398_));
  OAI22_X1   g00395(.A1(new_n1383_), .A2(new_n1396_), .B1(new_n1397_), .B2(new_n1398_), .ZN(new_n1399_));
  NAND4_X1   g00396(.A1(new_n1365_), .A2(new_n1370_), .A3(new_n1392_), .A4(new_n1394_), .ZN(new_n1400_));
  AOI21_X1   g00397(.A1(new_n1372_), .A2(new_n1380_), .B(new_n1378_), .ZN(new_n1401_));
  AOI21_X1   g00398(.A1(new_n1366_), .A2(new_n1368_), .B(new_n1367_), .ZN(new_n1402_));
  NAND2_X1   g00399(.A1(new_n1401_), .A2(new_n1402_), .ZN(new_n1403_));
  NAND2_X1   g00400(.A1(new_n1320_), .A2(new_n1325_), .ZN(new_n1404_));
  AOI21_X1   g00401(.A1(new_n1333_), .A2(new_n1341_), .B(new_n1404_), .ZN(new_n1405_));
  OR3_X2     g00402(.A1(new_n1405_), .A2(new_n1400_), .A3(new_n1403_), .Z(new_n1406_));
  NOR4_X1    g00403(.A1(new_n1406_), .A2(new_n1399_), .A3(new_n1357_), .A4(new_n1360_), .ZN(new_n1407_));
  NOR4_X1    g00404(.A1(new_n1386_), .A2(new_n1388_), .A3(new_n1381_), .A4(new_n1377_), .ZN(new_n1408_));
  INV_X1     g00405(.I(new_n1402_), .ZN(new_n1409_));
  NOR2_X1    g00406(.A1(new_n1408_), .A2(new_n1409_), .ZN(new_n1410_));
  NOR2_X1    g00407(.A1(new_n1400_), .A2(new_n1402_), .ZN(new_n1411_));
  OAI21_X1   g00408(.A1(new_n1410_), .A2(new_n1411_), .B(new_n1401_), .ZN(new_n1412_));
  INV_X1     g00409(.I(new_n1401_), .ZN(new_n1413_));
  NAND2_X1   g00410(.A1(new_n1400_), .A2(new_n1402_), .ZN(new_n1414_));
  NAND3_X1   g00411(.A1(new_n1389_), .A2(new_n1382_), .A3(new_n1409_), .ZN(new_n1415_));
  NAND3_X1   g00412(.A1(new_n1414_), .A2(new_n1415_), .A3(new_n1413_), .ZN(new_n1416_));
  NAND2_X1   g00413(.A1(new_n1412_), .A2(new_n1416_), .ZN(new_n1417_));
  OAI21_X1   g00414(.A1(new_n1358_), .A2(new_n1359_), .B(new_n1320_), .ZN(new_n1418_));
  NAND3_X1   g00415(.A1(new_n1356_), .A2(new_n1342_), .A3(new_n1321_), .ZN(new_n1419_));
  NAND2_X1   g00416(.A1(new_n1418_), .A2(new_n1419_), .ZN(new_n1420_));
  NOR2_X1    g00417(.A1(new_n1383_), .A2(new_n1396_), .ZN(new_n1421_));
  NOR2_X1    g00418(.A1(new_n1397_), .A2(new_n1398_), .ZN(new_n1422_));
  NOR4_X1    g00419(.A1(new_n1346_), .A2(new_n1348_), .A3(new_n1354_), .A4(new_n1352_), .ZN(new_n1423_));
  INV_X1     g00420(.I(new_n1403_), .ZN(new_n1424_));
  INV_X1     g00421(.I(new_n1404_), .ZN(new_n1425_));
  NAND4_X1   g00422(.A1(new_n1423_), .A2(new_n1408_), .A3(new_n1424_), .A4(new_n1425_), .ZN(new_n1426_));
  NOR3_X1    g00423(.A1(new_n1421_), .A2(new_n1422_), .A3(new_n1426_), .ZN(new_n1427_));
  NOR2_X1    g00424(.A1(new_n1420_), .A2(new_n1427_), .ZN(new_n1428_));
  NOR3_X1    g00425(.A1(new_n1428_), .A2(new_n1407_), .A3(new_n1417_), .ZN(new_n1429_));
  OAI22_X1   g00426(.A1(new_n1399_), .A2(new_n1426_), .B1(new_n1360_), .B2(new_n1357_), .ZN(new_n1430_));
  NAND2_X1   g00427(.A1(new_n1389_), .A2(new_n1395_), .ZN(new_n1431_));
  NAND2_X1   g00428(.A1(new_n1382_), .A2(new_n1371_), .ZN(new_n1432_));
  NAND2_X1   g00429(.A1(new_n1349_), .A2(new_n1341_), .ZN(new_n1433_));
  NAND2_X1   g00430(.A1(new_n1355_), .A2(new_n1333_), .ZN(new_n1434_));
  AOI22_X1   g00431(.A1(new_n1431_), .A2(new_n1432_), .B1(new_n1434_), .B2(new_n1433_), .ZN(new_n1435_));
  INV_X1     g00432(.I(new_n1426_), .ZN(new_n1436_));
  NAND4_X1   g00433(.A1(new_n1436_), .A2(new_n1435_), .A3(new_n1418_), .A4(new_n1419_), .ZN(new_n1437_));
  AOI21_X1   g00434(.A1(new_n1430_), .A2(new_n1437_), .B(new_n1417_), .ZN(new_n1438_));
  NOR2_X1    g00435(.A1(new_n1429_), .A2(new_n1438_), .ZN(new_n1439_));
  NAND2_X1   g00436(.A1(new_n1408_), .A2(new_n1424_), .ZN(new_n1440_));
  NOR2_X1    g00437(.A1(new_n1440_), .A2(new_n1405_), .ZN(new_n1441_));
  NAND4_X1   g00438(.A1(new_n1435_), .A2(new_n1418_), .A3(new_n1441_), .A4(new_n1419_), .ZN(new_n1442_));
  AOI21_X1   g00439(.A1(new_n1414_), .A2(new_n1415_), .B(new_n1413_), .ZN(new_n1443_));
  NOR3_X1    g00440(.A1(new_n1410_), .A2(new_n1411_), .A3(new_n1401_), .ZN(new_n1444_));
  NOR2_X1    g00441(.A1(new_n1444_), .A2(new_n1443_), .ZN(new_n1445_));
  NOR2_X1    g00442(.A1(new_n1360_), .A2(new_n1357_), .ZN(new_n1446_));
  NAND2_X1   g00443(.A1(new_n1431_), .A2(new_n1432_), .ZN(new_n1447_));
  NAND2_X1   g00444(.A1(new_n1434_), .A2(new_n1433_), .ZN(new_n1448_));
  NOR2_X1    g00445(.A1(new_n1400_), .A2(new_n1403_), .ZN(new_n1449_));
  NOR3_X1    g00446(.A1(new_n1333_), .A2(new_n1341_), .A3(new_n1404_), .ZN(new_n1450_));
  NAND4_X1   g00447(.A1(new_n1447_), .A2(new_n1448_), .A3(new_n1449_), .A4(new_n1450_), .ZN(new_n1451_));
  NAND2_X1   g00448(.A1(new_n1446_), .A2(new_n1451_), .ZN(new_n1452_));
  NAND3_X1   g00449(.A1(new_n1452_), .A2(new_n1442_), .A3(new_n1445_), .ZN(new_n1453_));
  AOI22_X1   g00450(.A1(new_n1436_), .A2(new_n1435_), .B1(new_n1418_), .B2(new_n1419_), .ZN(new_n1454_));
  NOR4_X1    g00451(.A1(new_n1399_), .A2(new_n1357_), .A3(new_n1360_), .A4(new_n1426_), .ZN(new_n1455_));
  OAI21_X1   g00452(.A1(new_n1454_), .A2(new_n1455_), .B(new_n1445_), .ZN(new_n1456_));
  NAND2_X1   g00453(.A1(new_n1448_), .A2(new_n1450_), .ZN(new_n1457_));
  NOR2_X1    g00454(.A1(new_n1421_), .A2(new_n1440_), .ZN(new_n1458_));
  NAND2_X1   g00455(.A1(new_n1458_), .A2(new_n1457_), .ZN(new_n1459_));
  INV_X1     g00456(.I(new_n1450_), .ZN(new_n1460_));
  NOR2_X1    g00457(.A1(new_n1422_), .A2(new_n1460_), .ZN(new_n1461_));
  OAI21_X1   g00458(.A1(new_n1383_), .A2(new_n1396_), .B(new_n1449_), .ZN(new_n1462_));
  NAND2_X1   g00459(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1463_));
  INV_X1     g00460(.I(\A[354] ), .ZN(new_n1464_));
  NOR2_X1    g00461(.A1(new_n1464_), .A2(\A[353] ), .ZN(new_n1465_));
  INV_X1     g00462(.I(\A[353] ), .ZN(new_n1466_));
  NOR2_X1    g00463(.A1(new_n1466_), .A2(\A[354] ), .ZN(new_n1467_));
  OAI21_X1   g00464(.A1(new_n1465_), .A2(new_n1467_), .B(\A[352] ), .ZN(new_n1468_));
  INV_X1     g00465(.I(\A[352] ), .ZN(new_n1469_));
  NOR2_X1    g00466(.A1(\A[353] ), .A2(\A[354] ), .ZN(new_n1470_));
  NAND2_X1   g00467(.A1(\A[353] ), .A2(\A[354] ), .ZN(new_n1471_));
  INV_X1     g00468(.I(new_n1471_), .ZN(new_n1472_));
  OAI21_X1   g00469(.A1(new_n1472_), .A2(new_n1470_), .B(new_n1469_), .ZN(new_n1473_));
  NAND2_X1   g00470(.A1(new_n1468_), .A2(new_n1473_), .ZN(new_n1474_));
  AOI21_X1   g00471(.A1(new_n1469_), .A2(new_n1471_), .B(new_n1470_), .ZN(new_n1475_));
  NAND4_X1   g00472(.A1(new_n1475_), .A2(\A[349] ), .A3(\A[350] ), .A4(\A[351] ), .ZN(new_n1476_));
  NOR2_X1    g00473(.A1(new_n1474_), .A2(new_n1476_), .ZN(new_n1477_));
  INV_X1     g00474(.I(\A[351] ), .ZN(new_n1478_));
  NOR2_X1    g00475(.A1(new_n1478_), .A2(\A[350] ), .ZN(new_n1479_));
  INV_X1     g00476(.I(\A[350] ), .ZN(new_n1480_));
  NOR2_X1    g00477(.A1(new_n1480_), .A2(\A[351] ), .ZN(new_n1481_));
  OAI21_X1   g00478(.A1(new_n1479_), .A2(new_n1481_), .B(\A[349] ), .ZN(new_n1482_));
  INV_X1     g00479(.I(\A[349] ), .ZN(new_n1483_));
  NOR2_X1    g00480(.A1(\A[350] ), .A2(\A[351] ), .ZN(new_n1484_));
  AND2_X2    g00481(.A1(\A[350] ), .A2(\A[351] ), .Z(new_n1485_));
  OAI21_X1   g00482(.A1(new_n1485_), .A2(new_n1484_), .B(new_n1483_), .ZN(new_n1486_));
  NAND2_X1   g00483(.A1(new_n1482_), .A2(new_n1486_), .ZN(new_n1487_));
  XOR2_X1    g00484(.A1(new_n1474_), .A2(new_n1487_), .Z(new_n1488_));
  INV_X1     g00485(.I(\A[343] ), .ZN(new_n1489_));
  INV_X1     g00486(.I(\A[344] ), .ZN(new_n1490_));
  NAND2_X1   g00487(.A1(new_n1490_), .A2(\A[345] ), .ZN(new_n1491_));
  INV_X1     g00488(.I(\A[345] ), .ZN(new_n1492_));
  NAND2_X1   g00489(.A1(new_n1492_), .A2(\A[344] ), .ZN(new_n1493_));
  AOI21_X1   g00490(.A1(new_n1491_), .A2(new_n1493_), .B(new_n1489_), .ZN(new_n1494_));
  NOR2_X1    g00491(.A1(\A[344] ), .A2(\A[345] ), .ZN(new_n1495_));
  INV_X1     g00492(.I(new_n1495_), .ZN(new_n1496_));
  NAND2_X1   g00493(.A1(\A[344] ), .A2(\A[345] ), .ZN(new_n1497_));
  AOI21_X1   g00494(.A1(new_n1496_), .A2(new_n1497_), .B(\A[343] ), .ZN(new_n1498_));
  NOR2_X1    g00495(.A1(new_n1498_), .A2(new_n1494_), .ZN(new_n1499_));
  INV_X1     g00496(.I(\A[346] ), .ZN(new_n1500_));
  INV_X1     g00497(.I(\A[347] ), .ZN(new_n1501_));
  NAND2_X1   g00498(.A1(new_n1501_), .A2(\A[348] ), .ZN(new_n1502_));
  INV_X1     g00499(.I(\A[348] ), .ZN(new_n1503_));
  NAND2_X1   g00500(.A1(new_n1503_), .A2(\A[347] ), .ZN(new_n1504_));
  AOI21_X1   g00501(.A1(new_n1502_), .A2(new_n1504_), .B(new_n1500_), .ZN(new_n1505_));
  OR2_X2     g00502(.A1(\A[347] ), .A2(\A[348] ), .Z(new_n1506_));
  NAND2_X1   g00503(.A1(\A[347] ), .A2(\A[348] ), .ZN(new_n1507_));
  AOI21_X1   g00504(.A1(new_n1506_), .A2(new_n1507_), .B(\A[346] ), .ZN(new_n1508_));
  NOR2_X1    g00505(.A1(new_n1505_), .A2(new_n1508_), .ZN(new_n1509_));
  NOR2_X1    g00506(.A1(\A[347] ), .A2(\A[348] ), .ZN(new_n1510_));
  AOI21_X1   g00507(.A1(new_n1500_), .A2(new_n1507_), .B(new_n1510_), .ZN(new_n1511_));
  AOI21_X1   g00508(.A1(new_n1489_), .A2(new_n1497_), .B(new_n1495_), .ZN(new_n1512_));
  NAND2_X1   g00509(.A1(new_n1511_), .A2(new_n1512_), .ZN(new_n1513_));
  INV_X1     g00510(.I(new_n1513_), .ZN(new_n1514_));
  NAND2_X1   g00511(.A1(new_n1488_), .A2(new_n1477_), .ZN(new_n1515_));
  AOI21_X1   g00512(.A1(new_n1459_), .A2(new_n1463_), .B(new_n1515_), .ZN(new_n1516_));
  AOI21_X1   g00513(.A1(new_n1453_), .A2(new_n1456_), .B(new_n1516_), .ZN(new_n1517_));
  NOR2_X1    g00514(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1518_));
  NOR2_X1    g00515(.A1(new_n1458_), .A2(new_n1457_), .ZN(new_n1519_));
  INV_X1     g00516(.I(new_n1515_), .ZN(new_n1520_));
  OAI21_X1   g00517(.A1(new_n1519_), .A2(new_n1518_), .B(new_n1520_), .ZN(new_n1521_));
  NOR3_X1    g00518(.A1(new_n1429_), .A2(new_n1521_), .A3(new_n1438_), .ZN(new_n1522_));
  NOR4_X1    g00519(.A1(new_n1494_), .A2(new_n1498_), .A3(new_n1505_), .A4(new_n1508_), .ZN(new_n1523_));
  INV_X1     g00520(.I(new_n1512_), .ZN(new_n1524_));
  NOR2_X1    g00521(.A1(new_n1523_), .A2(new_n1524_), .ZN(new_n1525_));
  NOR2_X1    g00522(.A1(new_n1492_), .A2(\A[344] ), .ZN(new_n1526_));
  NOR2_X1    g00523(.A1(new_n1490_), .A2(\A[345] ), .ZN(new_n1527_));
  OAI21_X1   g00524(.A1(new_n1526_), .A2(new_n1527_), .B(\A[343] ), .ZN(new_n1528_));
  INV_X1     g00525(.I(new_n1497_), .ZN(new_n1529_));
  OAI21_X1   g00526(.A1(new_n1529_), .A2(new_n1495_), .B(new_n1489_), .ZN(new_n1530_));
  NAND2_X1   g00527(.A1(new_n1528_), .A2(new_n1530_), .ZN(new_n1531_));
  NOR2_X1    g00528(.A1(new_n1503_), .A2(\A[347] ), .ZN(new_n1532_));
  NOR2_X1    g00529(.A1(new_n1501_), .A2(\A[348] ), .ZN(new_n1533_));
  OAI21_X1   g00530(.A1(new_n1532_), .A2(new_n1533_), .B(\A[346] ), .ZN(new_n1534_));
  AND2_X2    g00531(.A1(\A[347] ), .A2(\A[348] ), .Z(new_n1535_));
  OAI21_X1   g00532(.A1(new_n1535_), .A2(new_n1510_), .B(new_n1500_), .ZN(new_n1536_));
  NAND2_X1   g00533(.A1(new_n1534_), .A2(new_n1536_), .ZN(new_n1537_));
  NOR3_X1    g00534(.A1(new_n1531_), .A2(new_n1537_), .A3(new_n1512_), .ZN(new_n1538_));
  OAI21_X1   g00535(.A1(new_n1525_), .A2(new_n1538_), .B(new_n1511_), .ZN(new_n1539_));
  INV_X1     g00536(.I(new_n1511_), .ZN(new_n1540_));
  OAI21_X1   g00537(.A1(new_n1531_), .A2(new_n1537_), .B(new_n1512_), .ZN(new_n1541_));
  NAND3_X1   g00538(.A1(new_n1499_), .A2(new_n1509_), .A3(new_n1524_), .ZN(new_n1542_));
  NAND3_X1   g00539(.A1(new_n1541_), .A2(new_n1542_), .A3(new_n1540_), .ZN(new_n1543_));
  NAND2_X1   g00540(.A1(new_n1539_), .A2(new_n1543_), .ZN(new_n1544_));
  NAND2_X1   g00541(.A1(new_n1466_), .A2(\A[354] ), .ZN(new_n1545_));
  NAND2_X1   g00542(.A1(new_n1464_), .A2(\A[353] ), .ZN(new_n1546_));
  AOI21_X1   g00543(.A1(new_n1545_), .A2(new_n1546_), .B(new_n1469_), .ZN(new_n1547_));
  INV_X1     g00544(.I(new_n1470_), .ZN(new_n1548_));
  AOI21_X1   g00545(.A1(new_n1548_), .A2(new_n1471_), .B(\A[352] ), .ZN(new_n1549_));
  NOR2_X1    g00546(.A1(new_n1549_), .A2(new_n1547_), .ZN(new_n1550_));
  XOR2_X1    g00547(.A1(new_n1550_), .A2(new_n1487_), .Z(new_n1551_));
  NOR2_X1    g00548(.A1(new_n1531_), .A2(new_n1509_), .ZN(new_n1552_));
  NOR2_X1    g00549(.A1(new_n1499_), .A2(new_n1537_), .ZN(new_n1553_));
  NOR2_X1    g00550(.A1(new_n1552_), .A2(new_n1553_), .ZN(new_n1554_));
  NAND2_X1   g00551(.A1(new_n1480_), .A2(\A[351] ), .ZN(new_n1555_));
  NAND2_X1   g00552(.A1(new_n1478_), .A2(\A[350] ), .ZN(new_n1556_));
  AOI21_X1   g00553(.A1(new_n1555_), .A2(new_n1556_), .B(new_n1483_), .ZN(new_n1557_));
  INV_X1     g00554(.I(new_n1484_), .ZN(new_n1558_));
  NAND2_X1   g00555(.A1(\A[350] ), .A2(\A[351] ), .ZN(new_n1559_));
  AOI21_X1   g00556(.A1(new_n1558_), .A2(new_n1559_), .B(\A[349] ), .ZN(new_n1560_));
  NOR2_X1    g00557(.A1(new_n1560_), .A2(new_n1557_), .ZN(new_n1561_));
  AOI21_X1   g00558(.A1(new_n1483_), .A2(new_n1559_), .B(new_n1484_), .ZN(new_n1562_));
  INV_X1     g00559(.I(new_n1562_), .ZN(new_n1563_));
  AOI21_X1   g00560(.A1(new_n1550_), .A2(new_n1561_), .B(new_n1563_), .ZN(new_n1564_));
  NOR3_X1    g00561(.A1(new_n1474_), .A2(new_n1487_), .A3(new_n1562_), .ZN(new_n1565_));
  OAI21_X1   g00562(.A1(new_n1564_), .A2(new_n1565_), .B(new_n1475_), .ZN(new_n1566_));
  INV_X1     g00563(.I(new_n1475_), .ZN(new_n1567_));
  OAI21_X1   g00564(.A1(new_n1474_), .A2(new_n1487_), .B(new_n1562_), .ZN(new_n1568_));
  NAND3_X1   g00565(.A1(new_n1550_), .A2(new_n1561_), .A3(new_n1563_), .ZN(new_n1569_));
  NAND3_X1   g00566(.A1(new_n1569_), .A2(new_n1568_), .A3(new_n1567_), .ZN(new_n1570_));
  NAND2_X1   g00567(.A1(new_n1566_), .A2(new_n1570_), .ZN(new_n1571_));
  NAND2_X1   g00568(.A1(new_n1523_), .A2(new_n1514_), .ZN(new_n1572_));
  NAND2_X1   g00569(.A1(new_n1475_), .A2(new_n1562_), .ZN(new_n1573_));
  AOI21_X1   g00570(.A1(new_n1474_), .A2(new_n1487_), .B(new_n1573_), .ZN(new_n1574_));
  NOR2_X1    g00571(.A1(new_n1572_), .A2(new_n1574_), .ZN(new_n1575_));
  INV_X1     g00572(.I(new_n1575_), .ZN(new_n1576_));
  NOR4_X1    g00573(.A1(new_n1571_), .A2(new_n1551_), .A3(new_n1554_), .A4(new_n1576_), .ZN(new_n1577_));
  NOR3_X1    g00574(.A1(new_n1531_), .A2(new_n1537_), .A3(new_n1513_), .ZN(new_n1578_));
  NAND2_X1   g00575(.A1(new_n1578_), .A2(new_n1477_), .ZN(new_n1579_));
  NOR3_X1    g00576(.A1(new_n1551_), .A2(new_n1554_), .A3(new_n1579_), .ZN(new_n1580_));
  NAND2_X1   g00577(.A1(new_n1580_), .A2(new_n1544_), .ZN(new_n1581_));
  AOI21_X1   g00578(.A1(new_n1569_), .A2(new_n1568_), .B(new_n1567_), .ZN(new_n1582_));
  NOR3_X1    g00579(.A1(new_n1564_), .A2(new_n1565_), .A3(new_n1475_), .ZN(new_n1583_));
  NOR2_X1    g00580(.A1(new_n1583_), .A2(new_n1582_), .ZN(new_n1584_));
  OAI21_X1   g00581(.A1(new_n1544_), .A2(new_n1580_), .B(new_n1584_), .ZN(new_n1585_));
  AOI21_X1   g00582(.A1(new_n1541_), .A2(new_n1542_), .B(new_n1540_), .ZN(new_n1586_));
  NOR3_X1    g00583(.A1(new_n1525_), .A2(new_n1538_), .A3(new_n1511_), .ZN(new_n1587_));
  NOR2_X1    g00584(.A1(new_n1587_), .A2(new_n1586_), .ZN(new_n1588_));
  XOR2_X1    g00585(.A1(new_n1531_), .A2(new_n1537_), .Z(new_n1589_));
  NAND4_X1   g00586(.A1(new_n1488_), .A2(new_n1589_), .A3(new_n1477_), .A4(new_n1578_), .ZN(new_n1590_));
  NAND3_X1   g00587(.A1(new_n1590_), .A2(new_n1588_), .A3(new_n1571_), .ZN(new_n1591_));
  NAND2_X1   g00588(.A1(new_n1585_), .A2(new_n1591_), .ZN(new_n1592_));
  AOI22_X1   g00589(.A1(new_n1592_), .A2(new_n1581_), .B1(new_n1544_), .B2(new_n1577_), .ZN(new_n1593_));
  OAI22_X1   g00590(.A1(new_n1593_), .A2(new_n1439_), .B1(new_n1522_), .B2(new_n1517_), .ZN(new_n1594_));
  OAI21_X1   g00591(.A1(new_n1320_), .A2(new_n1325_), .B(new_n1423_), .ZN(new_n1595_));
  NAND2_X1   g00592(.A1(new_n1595_), .A2(new_n1404_), .ZN(new_n1596_));
  OAI21_X1   g00593(.A1(new_n1401_), .A2(new_n1402_), .B(new_n1408_), .ZN(new_n1597_));
  NAND2_X1   g00594(.A1(new_n1597_), .A2(new_n1403_), .ZN(new_n1598_));
  INV_X1     g00595(.I(new_n1598_), .ZN(new_n1599_));
  OAI21_X1   g00596(.A1(new_n1420_), .A2(new_n1427_), .B(new_n1417_), .ZN(new_n1600_));
  AOI21_X1   g00597(.A1(new_n1600_), .A2(new_n1442_), .B(new_n1599_), .ZN(new_n1601_));
  AOI21_X1   g00598(.A1(new_n1446_), .A2(new_n1451_), .B(new_n1445_), .ZN(new_n1602_));
  NOR3_X1    g00599(.A1(new_n1602_), .A2(new_n1407_), .A3(new_n1598_), .ZN(new_n1603_));
  OAI21_X1   g00600(.A1(new_n1603_), .A2(new_n1601_), .B(new_n1596_), .ZN(new_n1604_));
  INV_X1     g00601(.I(new_n1596_), .ZN(new_n1605_));
  OAI21_X1   g00602(.A1(new_n1602_), .A2(new_n1407_), .B(new_n1598_), .ZN(new_n1606_));
  NAND3_X1   g00603(.A1(new_n1600_), .A2(new_n1442_), .A3(new_n1599_), .ZN(new_n1607_));
  NAND3_X1   g00604(.A1(new_n1606_), .A2(new_n1607_), .A3(new_n1605_), .ZN(new_n1608_));
  NAND2_X1   g00605(.A1(new_n1604_), .A2(new_n1608_), .ZN(new_n1609_));
  NAND2_X1   g00606(.A1(new_n1567_), .A2(new_n1563_), .ZN(new_n1610_));
  NAND3_X1   g00607(.A1(new_n1610_), .A2(new_n1550_), .A3(new_n1561_), .ZN(new_n1611_));
  NAND2_X1   g00608(.A1(new_n1611_), .A2(new_n1573_), .ZN(new_n1612_));
  INV_X1     g00609(.I(new_n1612_), .ZN(new_n1613_));
  OAI21_X1   g00610(.A1(new_n1511_), .A2(new_n1512_), .B(new_n1523_), .ZN(new_n1614_));
  NAND2_X1   g00611(.A1(new_n1614_), .A2(new_n1513_), .ZN(new_n1615_));
  AOI21_X1   g00612(.A1(new_n1590_), .A2(new_n1584_), .B(new_n1588_), .ZN(new_n1616_));
  OAI21_X1   g00613(.A1(new_n1616_), .A2(new_n1577_), .B(new_n1615_), .ZN(new_n1617_));
  NOR2_X1    g00614(.A1(new_n1551_), .A2(new_n1554_), .ZN(new_n1618_));
  NAND3_X1   g00615(.A1(new_n1584_), .A2(new_n1618_), .A3(new_n1575_), .ZN(new_n1619_));
  INV_X1     g00616(.I(new_n1615_), .ZN(new_n1620_));
  OAI21_X1   g00617(.A1(new_n1571_), .A2(new_n1580_), .B(new_n1544_), .ZN(new_n1621_));
  NAND3_X1   g00618(.A1(new_n1621_), .A2(new_n1619_), .A3(new_n1620_), .ZN(new_n1622_));
  AOI21_X1   g00619(.A1(new_n1617_), .A2(new_n1622_), .B(new_n1613_), .ZN(new_n1623_));
  AOI21_X1   g00620(.A1(new_n1621_), .A2(new_n1619_), .B(new_n1620_), .ZN(new_n1624_));
  NOR3_X1    g00621(.A1(new_n1616_), .A2(new_n1577_), .A3(new_n1615_), .ZN(new_n1625_));
  NOR3_X1    g00622(.A1(new_n1625_), .A2(new_n1624_), .A3(new_n1612_), .ZN(new_n1626_));
  NOR2_X1    g00623(.A1(new_n1626_), .A2(new_n1623_), .ZN(new_n1627_));
  NAND2_X1   g00624(.A1(new_n1609_), .A2(new_n1627_), .ZN(new_n1628_));
  OAI21_X1   g00625(.A1(new_n1625_), .A2(new_n1624_), .B(new_n1612_), .ZN(new_n1629_));
  NAND3_X1   g00626(.A1(new_n1617_), .A2(new_n1622_), .A3(new_n1613_), .ZN(new_n1630_));
  NAND2_X1   g00627(.A1(new_n1629_), .A2(new_n1630_), .ZN(new_n1631_));
  NAND3_X1   g00628(.A1(new_n1631_), .A2(new_n1604_), .A3(new_n1608_), .ZN(new_n1632_));
  AOI21_X1   g00629(.A1(new_n1628_), .A2(new_n1632_), .B(new_n1594_), .ZN(new_n1633_));
  NAND2_X1   g00630(.A1(new_n1453_), .A2(new_n1456_), .ZN(new_n1634_));
  OAI21_X1   g00631(.A1(new_n1429_), .A2(new_n1438_), .B(new_n1521_), .ZN(new_n1635_));
  NAND3_X1   g00632(.A1(new_n1453_), .A2(new_n1456_), .A3(new_n1516_), .ZN(new_n1636_));
  NAND2_X1   g00633(.A1(new_n1577_), .A2(new_n1544_), .ZN(new_n1637_));
  AOI21_X1   g00634(.A1(new_n1590_), .A2(new_n1588_), .B(new_n1571_), .ZN(new_n1638_));
  NOR3_X1    g00635(.A1(new_n1584_), .A2(new_n1580_), .A3(new_n1544_), .ZN(new_n1639_));
  OAI21_X1   g00636(.A1(new_n1638_), .A2(new_n1639_), .B(new_n1581_), .ZN(new_n1640_));
  NAND2_X1   g00637(.A1(new_n1640_), .A2(new_n1637_), .ZN(new_n1641_));
  AOI22_X1   g00638(.A1(new_n1641_), .A2(new_n1634_), .B1(new_n1635_), .B2(new_n1636_), .ZN(new_n1642_));
  NAND4_X1   g00639(.A1(new_n1604_), .A2(new_n1608_), .A3(new_n1629_), .A4(new_n1630_), .ZN(new_n1643_));
  AOI21_X1   g00640(.A1(new_n1606_), .A2(new_n1607_), .B(new_n1605_), .ZN(new_n1644_));
  NOR3_X1    g00641(.A1(new_n1603_), .A2(new_n1601_), .A3(new_n1596_), .ZN(new_n1645_));
  OAI22_X1   g00642(.A1(new_n1645_), .A2(new_n1644_), .B1(new_n1623_), .B2(new_n1626_), .ZN(new_n1646_));
  AOI21_X1   g00643(.A1(new_n1646_), .A2(new_n1643_), .B(new_n1642_), .ZN(new_n1647_));
  NOR3_X1    g00644(.A1(new_n1633_), .A2(new_n1316_), .A3(new_n1647_), .ZN(new_n1648_));
  NOR3_X1    g00645(.A1(new_n1641_), .A2(new_n1517_), .A3(new_n1522_), .ZN(new_n1649_));
  INV_X1     g00646(.I(new_n1649_), .ZN(new_n1650_));
  NOR2_X1    g00647(.A1(new_n1519_), .A2(new_n1518_), .ZN(new_n1651_));
  INV_X1     g00648(.I(new_n1477_), .ZN(new_n1652_));
  NOR2_X1    g00649(.A1(new_n1551_), .A2(new_n1652_), .ZN(new_n1653_));
  NOR2_X1    g00650(.A1(new_n1651_), .A2(new_n1653_), .ZN(new_n1654_));
  NAND2_X1   g00651(.A1(new_n1459_), .A2(new_n1463_), .ZN(new_n1655_));
  INV_X1     g00652(.I(new_n1653_), .ZN(new_n1656_));
  NOR2_X1    g00653(.A1(new_n1655_), .A2(new_n1656_), .ZN(new_n1657_));
  NOR2_X1    g00654(.A1(new_n1197_), .A2(new_n1198_), .ZN(new_n1658_));
  INV_X1     g00655(.I(new_n1254_), .ZN(new_n1659_));
  NOR2_X1    g00656(.A1(new_n1658_), .A2(new_n1659_), .ZN(new_n1660_));
  NAND2_X1   g00657(.A1(new_n1118_), .A2(new_n1114_), .ZN(new_n1661_));
  NOR2_X1    g00658(.A1(new_n1661_), .A2(new_n1254_), .ZN(new_n1662_));
  NOR4_X1    g00659(.A1(new_n1654_), .A2(new_n1657_), .A3(new_n1660_), .A4(new_n1662_), .ZN(new_n1663_));
  NOR2_X1    g00660(.A1(new_n1649_), .A2(new_n1663_), .ZN(new_n1664_));
  INV_X1     g00661(.I(new_n1664_), .ZN(new_n1665_));
  NAND2_X1   g00662(.A1(new_n1649_), .A2(new_n1663_), .ZN(new_n1666_));
  NAND3_X1   g00663(.A1(new_n1305_), .A2(new_n1246_), .A3(new_n1265_), .ZN(new_n1667_));
  NAND2_X1   g00664(.A1(new_n1266_), .A2(new_n1206_), .ZN(new_n1668_));
  NAND2_X1   g00665(.A1(new_n1668_), .A2(new_n1667_), .ZN(new_n1669_));
  AOI22_X1   g00666(.A1(new_n1665_), .A2(new_n1666_), .B1(new_n1650_), .B2(new_n1669_), .ZN(new_n1670_));
  OAI21_X1   g00667(.A1(new_n1633_), .A2(new_n1647_), .B(new_n1316_), .ZN(new_n1671_));
  AOI21_X1   g00668(.A1(new_n1671_), .A2(new_n1670_), .B(new_n1648_), .ZN(new_n1672_));
  NOR2_X1    g00669(.A1(new_n1605_), .A2(new_n1599_), .ZN(new_n1673_));
  NAND2_X1   g00670(.A1(new_n1600_), .A2(new_n1442_), .ZN(new_n1674_));
  AOI21_X1   g00671(.A1(new_n1605_), .A2(new_n1599_), .B(new_n1674_), .ZN(new_n1675_));
  NOR2_X1    g00672(.A1(new_n1675_), .A2(new_n1673_), .ZN(new_n1676_));
  NOR2_X1    g00673(.A1(new_n1645_), .A2(new_n1644_), .ZN(new_n1677_));
  AOI21_X1   g00674(.A1(new_n1677_), .A2(new_n1627_), .B(new_n1642_), .ZN(new_n1678_));
  NAND2_X1   g00675(.A1(new_n1621_), .A2(new_n1619_), .ZN(new_n1679_));
  XOR2_X1    g00676(.A1(new_n1598_), .A2(new_n1596_), .Z(new_n1680_));
  XOR2_X1    g00677(.A1(new_n1615_), .A2(new_n1612_), .Z(new_n1681_));
  NOR4_X1    g00678(.A1(new_n1674_), .A2(new_n1679_), .A3(new_n1680_), .A4(new_n1681_), .ZN(new_n1682_));
  INV_X1     g00679(.I(new_n1682_), .ZN(new_n1683_));
  NOR2_X1    g00680(.A1(new_n1620_), .A2(new_n1613_), .ZN(new_n1684_));
  AOI21_X1   g00681(.A1(new_n1613_), .A2(new_n1620_), .B(new_n1679_), .ZN(new_n1685_));
  NOR2_X1    g00682(.A1(new_n1685_), .A2(new_n1684_), .ZN(new_n1686_));
  INV_X1     g00683(.I(new_n1686_), .ZN(new_n1687_));
  OAI21_X1   g00684(.A1(new_n1678_), .A2(new_n1683_), .B(new_n1687_), .ZN(new_n1688_));
  NAND2_X1   g00685(.A1(new_n1643_), .A2(new_n1594_), .ZN(new_n1689_));
  NAND3_X1   g00686(.A1(new_n1689_), .A2(new_n1682_), .A3(new_n1686_), .ZN(new_n1690_));
  AOI21_X1   g00687(.A1(new_n1688_), .A2(new_n1690_), .B(new_n1676_), .ZN(new_n1691_));
  INV_X1     g00688(.I(new_n1676_), .ZN(new_n1692_));
  AOI21_X1   g00689(.A1(new_n1689_), .A2(new_n1682_), .B(new_n1686_), .ZN(new_n1693_));
  NOR3_X1    g00690(.A1(new_n1678_), .A2(new_n1683_), .A3(new_n1687_), .ZN(new_n1694_));
  NOR3_X1    g00691(.A1(new_n1694_), .A2(new_n1693_), .A3(new_n1692_), .ZN(new_n1695_));
  NAND2_X1   g00692(.A1(new_n1273_), .A2(new_n1271_), .ZN(new_n1696_));
  NOR2_X1    g00693(.A1(new_n1269_), .A2(new_n1268_), .ZN(new_n1697_));
  OAI21_X1   g00694(.A1(new_n1271_), .A2(new_n1273_), .B(new_n1697_), .ZN(new_n1698_));
  NAND2_X1   g00695(.A1(new_n1698_), .A2(new_n1696_), .ZN(new_n1699_));
  INV_X1     g00696(.I(new_n1699_), .ZN(new_n1700_));
  INV_X1     g00697(.I(new_n1289_), .ZN(new_n1701_));
  NAND3_X1   g00698(.A1(new_n1267_), .A2(new_n1275_), .A3(new_n1701_), .ZN(new_n1702_));
  OAI21_X1   g00699(.A1(new_n1282_), .A2(new_n1234_), .B(new_n1284_), .ZN(new_n1703_));
  NAND3_X1   g00700(.A1(new_n1287_), .A2(new_n1276_), .A3(new_n1285_), .ZN(new_n1704_));
  NAND2_X1   g00701(.A1(new_n1296_), .A2(new_n1704_), .ZN(new_n1705_));
  NAND2_X1   g00702(.A1(new_n1705_), .A2(new_n1703_), .ZN(new_n1706_));
  NAND2_X1   g00703(.A1(new_n1702_), .A2(new_n1706_), .ZN(new_n1707_));
  INV_X1     g00704(.I(new_n1313_), .ZN(new_n1708_));
  NAND3_X1   g00705(.A1(new_n1667_), .A2(new_n1207_), .A3(new_n1312_), .ZN(new_n1709_));
  INV_X1     g00706(.I(new_n1706_), .ZN(new_n1710_));
  NAND3_X1   g00707(.A1(new_n1709_), .A2(new_n1708_), .A3(new_n1710_), .ZN(new_n1711_));
  AOI21_X1   g00708(.A1(new_n1707_), .A2(new_n1711_), .B(new_n1700_), .ZN(new_n1712_));
  AOI21_X1   g00709(.A1(new_n1709_), .A2(new_n1708_), .B(new_n1710_), .ZN(new_n1713_));
  NOR4_X1    g00710(.A1(new_n1311_), .A2(new_n1294_), .A3(new_n1289_), .A4(new_n1706_), .ZN(new_n1714_));
  NOR3_X1    g00711(.A1(new_n1713_), .A2(new_n1699_), .A3(new_n1714_), .ZN(new_n1715_));
  NOR2_X1    g00712(.A1(new_n1712_), .A2(new_n1715_), .ZN(new_n1716_));
  OAI21_X1   g00713(.A1(new_n1691_), .A2(new_n1695_), .B(new_n1716_), .ZN(new_n1717_));
  OAI21_X1   g00714(.A1(new_n1694_), .A2(new_n1693_), .B(new_n1692_), .ZN(new_n1718_));
  NAND3_X1   g00715(.A1(new_n1688_), .A2(new_n1690_), .A3(new_n1676_), .ZN(new_n1719_));
  OAI21_X1   g00716(.A1(new_n1713_), .A2(new_n1714_), .B(new_n1699_), .ZN(new_n1720_));
  NAND3_X1   g00717(.A1(new_n1707_), .A2(new_n1700_), .A3(new_n1711_), .ZN(new_n1721_));
  NAND2_X1   g00718(.A1(new_n1721_), .A2(new_n1720_), .ZN(new_n1722_));
  NAND3_X1   g00719(.A1(new_n1722_), .A2(new_n1718_), .A3(new_n1719_), .ZN(new_n1723_));
  AOI21_X1   g00720(.A1(new_n1717_), .A2(new_n1723_), .B(new_n1672_), .ZN(new_n1724_));
  XOR2_X1    g00721(.A1(new_n1289_), .A2(new_n1275_), .Z(new_n1725_));
  NOR2_X1    g00722(.A1(new_n1725_), .A2(new_n1311_), .ZN(new_n1726_));
  XOR2_X1    g00723(.A1(new_n1289_), .A2(new_n1294_), .Z(new_n1727_));
  NOR2_X1    g00724(.A1(new_n1727_), .A2(new_n1267_), .ZN(new_n1728_));
  NOR2_X1    g00725(.A1(new_n1728_), .A2(new_n1726_), .ZN(new_n1729_));
  NOR2_X1    g00726(.A1(new_n1677_), .A2(new_n1631_), .ZN(new_n1730_));
  NOR2_X1    g00727(.A1(new_n1609_), .A2(new_n1627_), .ZN(new_n1731_));
  OAI21_X1   g00728(.A1(new_n1730_), .A2(new_n1731_), .B(new_n1642_), .ZN(new_n1732_));
  INV_X1     g00729(.I(new_n1643_), .ZN(new_n1733_));
  AOI22_X1   g00730(.A1(new_n1604_), .A2(new_n1608_), .B1(new_n1629_), .B2(new_n1630_), .ZN(new_n1734_));
  OAI21_X1   g00731(.A1(new_n1733_), .A2(new_n1734_), .B(new_n1594_), .ZN(new_n1735_));
  NAND3_X1   g00732(.A1(new_n1729_), .A2(new_n1732_), .A3(new_n1735_), .ZN(new_n1736_));
  INV_X1     g00733(.I(new_n1670_), .ZN(new_n1737_));
  AOI21_X1   g00734(.A1(new_n1732_), .A2(new_n1735_), .B(new_n1729_), .ZN(new_n1738_));
  OAI21_X1   g00735(.A1(new_n1738_), .A2(new_n1737_), .B(new_n1736_), .ZN(new_n1739_));
  NAND4_X1   g00736(.A1(new_n1718_), .A2(new_n1719_), .A3(new_n1720_), .A4(new_n1721_), .ZN(new_n1740_));
  OAI21_X1   g00737(.A1(new_n1691_), .A2(new_n1695_), .B(new_n1722_), .ZN(new_n1741_));
  AOI21_X1   g00738(.A1(new_n1741_), .A2(new_n1740_), .B(new_n1739_), .ZN(new_n1742_));
  INV_X1     g00739(.I(\A[286] ), .ZN(new_n1743_));
  NOR2_X1    g00740(.A1(\A[287] ), .A2(\A[288] ), .ZN(new_n1744_));
  NAND2_X1   g00741(.A1(\A[287] ), .A2(\A[288] ), .ZN(new_n1745_));
  AOI21_X1   g00742(.A1(new_n1743_), .A2(new_n1745_), .B(new_n1744_), .ZN(new_n1746_));
  INV_X1     g00743(.I(new_n1746_), .ZN(new_n1747_));
  INV_X1     g00744(.I(\A[283] ), .ZN(new_n1748_));
  NOR2_X1    g00745(.A1(\A[284] ), .A2(\A[285] ), .ZN(new_n1749_));
  NAND2_X1   g00746(.A1(\A[284] ), .A2(\A[285] ), .ZN(new_n1750_));
  AOI21_X1   g00747(.A1(new_n1748_), .A2(new_n1750_), .B(new_n1749_), .ZN(new_n1751_));
  INV_X1     g00748(.I(\A[284] ), .ZN(new_n1752_));
  NAND2_X1   g00749(.A1(new_n1752_), .A2(\A[285] ), .ZN(new_n1753_));
  INV_X1     g00750(.I(new_n1753_), .ZN(new_n1754_));
  NOR2_X1    g00751(.A1(new_n1752_), .A2(\A[285] ), .ZN(new_n1755_));
  OAI21_X1   g00752(.A1(new_n1754_), .A2(new_n1755_), .B(\A[283] ), .ZN(new_n1756_));
  INV_X1     g00753(.I(new_n1750_), .ZN(new_n1757_));
  OAI21_X1   g00754(.A1(new_n1757_), .A2(new_n1749_), .B(new_n1748_), .ZN(new_n1758_));
  INV_X1     g00755(.I(\A[288] ), .ZN(new_n1759_));
  NOR2_X1    g00756(.A1(new_n1759_), .A2(\A[287] ), .ZN(new_n1760_));
  INV_X1     g00757(.I(\A[287] ), .ZN(new_n1761_));
  NOR2_X1    g00758(.A1(new_n1761_), .A2(\A[288] ), .ZN(new_n1762_));
  OAI21_X1   g00759(.A1(new_n1760_), .A2(new_n1762_), .B(\A[286] ), .ZN(new_n1763_));
  INV_X1     g00760(.I(new_n1745_), .ZN(new_n1764_));
  OAI21_X1   g00761(.A1(new_n1764_), .A2(new_n1744_), .B(new_n1743_), .ZN(new_n1765_));
  NAND4_X1   g00762(.A1(new_n1756_), .A2(new_n1758_), .A3(new_n1765_), .A4(new_n1763_), .ZN(new_n1766_));
  NAND2_X1   g00763(.A1(new_n1766_), .A2(new_n1751_), .ZN(new_n1767_));
  INV_X1     g00764(.I(new_n1751_), .ZN(new_n1768_));
  INV_X1     g00765(.I(\A[285] ), .ZN(new_n1769_));
  NAND2_X1   g00766(.A1(new_n1769_), .A2(\A[284] ), .ZN(new_n1770_));
  AOI21_X1   g00767(.A1(new_n1753_), .A2(new_n1770_), .B(new_n1748_), .ZN(new_n1771_));
  INV_X1     g00768(.I(new_n1749_), .ZN(new_n1772_));
  AOI21_X1   g00769(.A1(new_n1772_), .A2(new_n1750_), .B(\A[283] ), .ZN(new_n1773_));
  NAND2_X1   g00770(.A1(new_n1761_), .A2(\A[288] ), .ZN(new_n1774_));
  NAND2_X1   g00771(.A1(new_n1759_), .A2(\A[287] ), .ZN(new_n1775_));
  AOI21_X1   g00772(.A1(new_n1774_), .A2(new_n1775_), .B(new_n1743_), .ZN(new_n1776_));
  INV_X1     g00773(.I(new_n1744_), .ZN(new_n1777_));
  AOI21_X1   g00774(.A1(new_n1777_), .A2(new_n1745_), .B(\A[286] ), .ZN(new_n1778_));
  NOR4_X1    g00775(.A1(new_n1771_), .A2(new_n1773_), .A3(new_n1778_), .A4(new_n1776_), .ZN(new_n1779_));
  NAND2_X1   g00776(.A1(new_n1779_), .A2(new_n1768_), .ZN(new_n1780_));
  AOI21_X1   g00777(.A1(new_n1767_), .A2(new_n1780_), .B(new_n1747_), .ZN(new_n1781_));
  NOR2_X1    g00778(.A1(new_n1779_), .A2(new_n1768_), .ZN(new_n1782_));
  NOR2_X1    g00779(.A1(new_n1766_), .A2(new_n1751_), .ZN(new_n1783_));
  NOR3_X1    g00780(.A1(new_n1783_), .A2(new_n1782_), .A3(new_n1746_), .ZN(new_n1784_));
  OR2_X2     g00781(.A1(new_n1781_), .A2(new_n1784_), .Z(new_n1785_));
  INV_X1     g00782(.I(\A[292] ), .ZN(new_n1786_));
  NOR2_X1    g00783(.A1(\A[293] ), .A2(\A[294] ), .ZN(new_n1787_));
  NAND2_X1   g00784(.A1(\A[293] ), .A2(\A[294] ), .ZN(new_n1788_));
  AOI21_X1   g00785(.A1(new_n1786_), .A2(new_n1788_), .B(new_n1787_), .ZN(new_n1789_));
  INV_X1     g00786(.I(\A[289] ), .ZN(new_n1790_));
  NOR2_X1    g00787(.A1(\A[290] ), .A2(\A[291] ), .ZN(new_n1791_));
  NAND2_X1   g00788(.A1(\A[290] ), .A2(\A[291] ), .ZN(new_n1792_));
  AOI21_X1   g00789(.A1(new_n1790_), .A2(new_n1792_), .B(new_n1791_), .ZN(new_n1793_));
  NAND2_X1   g00790(.A1(new_n1789_), .A2(new_n1793_), .ZN(new_n1794_));
  INV_X1     g00791(.I(\A[290] ), .ZN(new_n1795_));
  NAND2_X1   g00792(.A1(new_n1795_), .A2(\A[291] ), .ZN(new_n1796_));
  INV_X1     g00793(.I(\A[291] ), .ZN(new_n1797_));
  NAND2_X1   g00794(.A1(new_n1797_), .A2(\A[290] ), .ZN(new_n1798_));
  AOI21_X1   g00795(.A1(new_n1796_), .A2(new_n1798_), .B(new_n1790_), .ZN(new_n1799_));
  INV_X1     g00796(.I(new_n1791_), .ZN(new_n1800_));
  AOI21_X1   g00797(.A1(new_n1800_), .A2(new_n1792_), .B(\A[289] ), .ZN(new_n1801_));
  NOR2_X1    g00798(.A1(new_n1801_), .A2(new_n1799_), .ZN(new_n1802_));
  INV_X1     g00799(.I(\A[294] ), .ZN(new_n1803_));
  NOR2_X1    g00800(.A1(new_n1803_), .A2(\A[293] ), .ZN(new_n1804_));
  INV_X1     g00801(.I(\A[293] ), .ZN(new_n1805_));
  NOR2_X1    g00802(.A1(new_n1805_), .A2(\A[294] ), .ZN(new_n1806_));
  OAI21_X1   g00803(.A1(new_n1804_), .A2(new_n1806_), .B(\A[292] ), .ZN(new_n1807_));
  AND2_X2    g00804(.A1(\A[293] ), .A2(\A[294] ), .Z(new_n1808_));
  OAI21_X1   g00805(.A1(new_n1808_), .A2(new_n1787_), .B(new_n1786_), .ZN(new_n1809_));
  NAND2_X1   g00806(.A1(new_n1807_), .A2(new_n1809_), .ZN(new_n1810_));
  NAND2_X1   g00807(.A1(new_n1802_), .A2(new_n1810_), .ZN(new_n1811_));
  NOR2_X1    g00808(.A1(new_n1797_), .A2(\A[290] ), .ZN(new_n1812_));
  NOR2_X1    g00809(.A1(new_n1795_), .A2(\A[291] ), .ZN(new_n1813_));
  OAI21_X1   g00810(.A1(new_n1812_), .A2(new_n1813_), .B(\A[289] ), .ZN(new_n1814_));
  INV_X1     g00811(.I(new_n1792_), .ZN(new_n1815_));
  OAI21_X1   g00812(.A1(new_n1815_), .A2(new_n1791_), .B(new_n1790_), .ZN(new_n1816_));
  NAND2_X1   g00813(.A1(new_n1814_), .A2(new_n1816_), .ZN(new_n1817_));
  NAND2_X1   g00814(.A1(new_n1805_), .A2(\A[294] ), .ZN(new_n1818_));
  NAND2_X1   g00815(.A1(new_n1803_), .A2(\A[293] ), .ZN(new_n1819_));
  AOI21_X1   g00816(.A1(new_n1818_), .A2(new_n1819_), .B(new_n1786_), .ZN(new_n1820_));
  INV_X1     g00817(.I(new_n1787_), .ZN(new_n1821_));
  AOI21_X1   g00818(.A1(new_n1821_), .A2(new_n1788_), .B(\A[292] ), .ZN(new_n1822_));
  NOR2_X1    g00819(.A1(new_n1822_), .A2(new_n1820_), .ZN(new_n1823_));
  NAND2_X1   g00820(.A1(new_n1823_), .A2(new_n1817_), .ZN(new_n1824_));
  AOI21_X1   g00821(.A1(new_n1824_), .A2(new_n1811_), .B(new_n1794_), .ZN(new_n1825_));
  INV_X1     g00822(.I(new_n1789_), .ZN(new_n1826_));
  NAND4_X1   g00823(.A1(new_n1814_), .A2(new_n1807_), .A3(new_n1816_), .A4(new_n1809_), .ZN(new_n1827_));
  NAND2_X1   g00824(.A1(new_n1827_), .A2(new_n1793_), .ZN(new_n1828_));
  INV_X1     g00825(.I(new_n1793_), .ZN(new_n1829_));
  NAND3_X1   g00826(.A1(new_n1802_), .A2(new_n1823_), .A3(new_n1829_), .ZN(new_n1830_));
  AOI21_X1   g00827(.A1(new_n1828_), .A2(new_n1830_), .B(new_n1826_), .ZN(new_n1831_));
  AOI21_X1   g00828(.A1(new_n1802_), .A2(new_n1823_), .B(new_n1829_), .ZN(new_n1832_));
  NOR3_X1    g00829(.A1(new_n1817_), .A2(new_n1810_), .A3(new_n1793_), .ZN(new_n1833_));
  NOR3_X1    g00830(.A1(new_n1832_), .A2(new_n1833_), .A3(new_n1789_), .ZN(new_n1834_));
  NOR3_X1    g00831(.A1(new_n1831_), .A2(new_n1834_), .A3(new_n1825_), .ZN(new_n1835_));
  INV_X1     g00832(.I(new_n1794_), .ZN(new_n1836_));
  NOR4_X1    g00833(.A1(new_n1799_), .A2(new_n1801_), .A3(new_n1822_), .A4(new_n1820_), .ZN(new_n1837_));
  NAND2_X1   g00834(.A1(new_n1837_), .A2(new_n1836_), .ZN(new_n1838_));
  NAND2_X1   g00835(.A1(new_n1817_), .A2(new_n1810_), .ZN(new_n1839_));
  NAND2_X1   g00836(.A1(new_n1839_), .A2(new_n1827_), .ZN(new_n1840_));
  OAI22_X1   g00837(.A1(new_n1771_), .A2(new_n1773_), .B1(new_n1778_), .B2(new_n1776_), .ZN(new_n1841_));
  NAND2_X1   g00838(.A1(new_n1766_), .A2(new_n1841_), .ZN(new_n1842_));
  NAND2_X1   g00839(.A1(new_n1746_), .A2(new_n1751_), .ZN(new_n1843_));
  INV_X1     g00840(.I(new_n1843_), .ZN(new_n1844_));
  NAND2_X1   g00841(.A1(new_n1779_), .A2(new_n1844_), .ZN(new_n1845_));
  NOR4_X1    g00842(.A1(new_n1840_), .A2(new_n1842_), .A3(new_n1845_), .A4(new_n1838_), .ZN(new_n1846_));
  NAND2_X1   g00843(.A1(new_n1835_), .A2(new_n1846_), .ZN(new_n1847_));
  NOR2_X1    g00844(.A1(new_n1823_), .A2(new_n1817_), .ZN(new_n1848_));
  NOR2_X1    g00845(.A1(new_n1802_), .A2(new_n1810_), .ZN(new_n1849_));
  OAI21_X1   g00846(.A1(new_n1848_), .A2(new_n1849_), .B(new_n1836_), .ZN(new_n1850_));
  OAI21_X1   g00847(.A1(new_n1832_), .A2(new_n1833_), .B(new_n1789_), .ZN(new_n1851_));
  NAND3_X1   g00848(.A1(new_n1828_), .A2(new_n1830_), .A3(new_n1826_), .ZN(new_n1852_));
  NAND3_X1   g00849(.A1(new_n1852_), .A2(new_n1851_), .A3(new_n1850_), .ZN(new_n1853_));
  NOR2_X1    g00850(.A1(new_n1827_), .A2(new_n1794_), .ZN(new_n1854_));
  AOI22_X1   g00851(.A1(new_n1814_), .A2(new_n1816_), .B1(new_n1807_), .B2(new_n1809_), .ZN(new_n1855_));
  NOR2_X1    g00852(.A1(new_n1837_), .A2(new_n1855_), .ZN(new_n1856_));
  AOI22_X1   g00853(.A1(new_n1756_), .A2(new_n1758_), .B1(new_n1765_), .B2(new_n1763_), .ZN(new_n1857_));
  NOR2_X1    g00854(.A1(new_n1857_), .A2(new_n1779_), .ZN(new_n1858_));
  NOR2_X1    g00855(.A1(new_n1766_), .A2(new_n1843_), .ZN(new_n1859_));
  NAND4_X1   g00856(.A1(new_n1858_), .A2(new_n1859_), .A3(new_n1856_), .A4(new_n1854_), .ZN(new_n1860_));
  NAND2_X1   g00857(.A1(new_n1853_), .A2(new_n1860_), .ZN(new_n1861_));
  AOI21_X1   g00858(.A1(new_n1847_), .A2(new_n1861_), .B(new_n1785_), .ZN(new_n1862_));
  NOR2_X1    g00859(.A1(new_n1835_), .A2(new_n1860_), .ZN(new_n1863_));
  NOR2_X1    g00860(.A1(new_n1831_), .A2(new_n1834_), .ZN(new_n1864_));
  NAND3_X1   g00861(.A1(new_n1858_), .A2(new_n1856_), .A3(new_n1854_), .ZN(new_n1865_));
  INV_X1     g00862(.I(new_n1865_), .ZN(new_n1866_));
  NAND2_X1   g00863(.A1(new_n1850_), .A2(new_n1859_), .ZN(new_n1867_));
  AOI21_X1   g00864(.A1(new_n1866_), .A2(new_n1864_), .B(new_n1867_), .ZN(new_n1868_));
  NOR3_X1    g00865(.A1(new_n1868_), .A2(new_n1863_), .A3(new_n1785_), .ZN(new_n1869_));
  NOR2_X1    g00866(.A1(new_n1869_), .A2(new_n1862_), .ZN(new_n1870_));
  NOR2_X1    g00867(.A1(new_n1781_), .A2(new_n1784_), .ZN(new_n1871_));
  NOR4_X1    g00868(.A1(new_n1860_), .A2(new_n1825_), .A3(new_n1831_), .A4(new_n1834_), .ZN(new_n1872_));
  NOR2_X1    g00869(.A1(new_n1835_), .A2(new_n1846_), .ZN(new_n1873_));
  OAI21_X1   g00870(.A1(new_n1873_), .A2(new_n1872_), .B(new_n1871_), .ZN(new_n1874_));
  NAND2_X1   g00871(.A1(new_n1853_), .A2(new_n1846_), .ZN(new_n1875_));
  NAND2_X1   g00872(.A1(new_n1852_), .A2(new_n1851_), .ZN(new_n1876_));
  NOR2_X1    g00873(.A1(new_n1825_), .A2(new_n1845_), .ZN(new_n1877_));
  OAI21_X1   g00874(.A1(new_n1876_), .A2(new_n1865_), .B(new_n1877_), .ZN(new_n1878_));
  NAND3_X1   g00875(.A1(new_n1878_), .A2(new_n1875_), .A3(new_n1871_), .ZN(new_n1879_));
  NAND2_X1   g00876(.A1(new_n1856_), .A2(new_n1854_), .ZN(new_n1880_));
  NOR2_X1    g00877(.A1(new_n1842_), .A2(new_n1845_), .ZN(new_n1881_));
  NAND2_X1   g00878(.A1(new_n1881_), .A2(new_n1880_), .ZN(new_n1882_));
  NOR2_X1    g00879(.A1(new_n1840_), .A2(new_n1838_), .ZN(new_n1883_));
  NAND2_X1   g00880(.A1(new_n1858_), .A2(new_n1859_), .ZN(new_n1884_));
  NAND2_X1   g00881(.A1(new_n1883_), .A2(new_n1884_), .ZN(new_n1885_));
  NAND2_X1   g00882(.A1(new_n1885_), .A2(new_n1882_), .ZN(new_n1886_));
  INV_X1     g00883(.I(\A[279] ), .ZN(new_n1887_));
  NOR2_X1    g00884(.A1(new_n1887_), .A2(\A[278] ), .ZN(new_n1888_));
  INV_X1     g00885(.I(\A[278] ), .ZN(new_n1889_));
  NOR2_X1    g00886(.A1(new_n1889_), .A2(\A[279] ), .ZN(new_n1890_));
  OAI21_X1   g00887(.A1(new_n1888_), .A2(new_n1890_), .B(\A[277] ), .ZN(new_n1891_));
  INV_X1     g00888(.I(\A[277] ), .ZN(new_n1892_));
  NOR2_X1    g00889(.A1(\A[278] ), .A2(\A[279] ), .ZN(new_n1893_));
  NAND2_X1   g00890(.A1(\A[278] ), .A2(\A[279] ), .ZN(new_n1894_));
  INV_X1     g00891(.I(new_n1894_), .ZN(new_n1895_));
  OAI21_X1   g00892(.A1(new_n1895_), .A2(new_n1893_), .B(new_n1892_), .ZN(new_n1896_));
  NAND2_X1   g00893(.A1(new_n1891_), .A2(new_n1896_), .ZN(new_n1897_));
  INV_X1     g00894(.I(\A[282] ), .ZN(new_n1898_));
  NOR2_X1    g00895(.A1(new_n1898_), .A2(\A[281] ), .ZN(new_n1899_));
  INV_X1     g00896(.I(\A[281] ), .ZN(new_n1900_));
  NOR2_X1    g00897(.A1(new_n1900_), .A2(\A[282] ), .ZN(new_n1901_));
  OAI21_X1   g00898(.A1(new_n1899_), .A2(new_n1901_), .B(\A[280] ), .ZN(new_n1902_));
  INV_X1     g00899(.I(\A[280] ), .ZN(new_n1903_));
  NOR2_X1    g00900(.A1(\A[281] ), .A2(\A[282] ), .ZN(new_n1904_));
  AND2_X2    g00901(.A1(\A[281] ), .A2(\A[282] ), .Z(new_n1905_));
  OAI21_X1   g00902(.A1(new_n1905_), .A2(new_n1904_), .B(new_n1903_), .ZN(new_n1906_));
  NAND2_X1   g00903(.A1(new_n1902_), .A2(new_n1906_), .ZN(new_n1907_));
  NAND2_X1   g00904(.A1(\A[281] ), .A2(\A[282] ), .ZN(new_n1908_));
  AOI21_X1   g00905(.A1(new_n1903_), .A2(new_n1908_), .B(new_n1904_), .ZN(new_n1909_));
  AOI21_X1   g00906(.A1(new_n1892_), .A2(new_n1894_), .B(new_n1893_), .ZN(new_n1910_));
  NAND2_X1   g00907(.A1(new_n1909_), .A2(new_n1910_), .ZN(new_n1911_));
  NOR3_X1    g00908(.A1(new_n1897_), .A2(new_n1907_), .A3(new_n1911_), .ZN(new_n1912_));
  NOR2_X1    g00909(.A1(new_n1897_), .A2(new_n1907_), .ZN(new_n1913_));
  NAND2_X1   g00910(.A1(new_n1889_), .A2(\A[279] ), .ZN(new_n1914_));
  NAND2_X1   g00911(.A1(new_n1887_), .A2(\A[278] ), .ZN(new_n1915_));
  AOI21_X1   g00912(.A1(new_n1914_), .A2(new_n1915_), .B(new_n1892_), .ZN(new_n1916_));
  INV_X1     g00913(.I(new_n1893_), .ZN(new_n1917_));
  AOI21_X1   g00914(.A1(new_n1917_), .A2(new_n1894_), .B(\A[277] ), .ZN(new_n1918_));
  NOR2_X1    g00915(.A1(new_n1918_), .A2(new_n1916_), .ZN(new_n1919_));
  NAND2_X1   g00916(.A1(new_n1900_), .A2(\A[282] ), .ZN(new_n1920_));
  NAND2_X1   g00917(.A1(new_n1898_), .A2(\A[281] ), .ZN(new_n1921_));
  AOI21_X1   g00918(.A1(new_n1920_), .A2(new_n1921_), .B(new_n1903_), .ZN(new_n1922_));
  NAND2_X1   g00919(.A1(new_n1900_), .A2(new_n1898_), .ZN(new_n1923_));
  AOI21_X1   g00920(.A1(new_n1923_), .A2(new_n1908_), .B(\A[280] ), .ZN(new_n1924_));
  NOR2_X1    g00921(.A1(new_n1924_), .A2(new_n1922_), .ZN(new_n1925_));
  NOR2_X1    g00922(.A1(new_n1919_), .A2(new_n1925_), .ZN(new_n1926_));
  NOR2_X1    g00923(.A1(new_n1926_), .A2(new_n1913_), .ZN(new_n1927_));
  INV_X1     g00924(.I(\A[271] ), .ZN(new_n1928_));
  INV_X1     g00925(.I(\A[272] ), .ZN(new_n1929_));
  NAND2_X1   g00926(.A1(new_n1929_), .A2(\A[273] ), .ZN(new_n1930_));
  INV_X1     g00927(.I(\A[273] ), .ZN(new_n1931_));
  NAND2_X1   g00928(.A1(new_n1931_), .A2(\A[272] ), .ZN(new_n1932_));
  AOI21_X1   g00929(.A1(new_n1930_), .A2(new_n1932_), .B(new_n1928_), .ZN(new_n1933_));
  NOR2_X1    g00930(.A1(\A[272] ), .A2(\A[273] ), .ZN(new_n1934_));
  INV_X1     g00931(.I(new_n1934_), .ZN(new_n1935_));
  NAND2_X1   g00932(.A1(\A[272] ), .A2(\A[273] ), .ZN(new_n1936_));
  AOI21_X1   g00933(.A1(new_n1935_), .A2(new_n1936_), .B(\A[271] ), .ZN(new_n1937_));
  NOR2_X1    g00934(.A1(new_n1937_), .A2(new_n1933_), .ZN(new_n1938_));
  INV_X1     g00935(.I(\A[274] ), .ZN(new_n1939_));
  INV_X1     g00936(.I(\A[275] ), .ZN(new_n1940_));
  NAND2_X1   g00937(.A1(new_n1940_), .A2(\A[276] ), .ZN(new_n1941_));
  INV_X1     g00938(.I(\A[276] ), .ZN(new_n1942_));
  NAND2_X1   g00939(.A1(new_n1942_), .A2(\A[275] ), .ZN(new_n1943_));
  AOI21_X1   g00940(.A1(new_n1941_), .A2(new_n1943_), .B(new_n1939_), .ZN(new_n1944_));
  OR2_X2     g00941(.A1(\A[275] ), .A2(\A[276] ), .Z(new_n1945_));
  NAND2_X1   g00942(.A1(\A[275] ), .A2(\A[276] ), .ZN(new_n1946_));
  AOI21_X1   g00943(.A1(new_n1945_), .A2(new_n1946_), .B(\A[274] ), .ZN(new_n1947_));
  NOR2_X1    g00944(.A1(new_n1944_), .A2(new_n1947_), .ZN(new_n1948_));
  NOR2_X1    g00945(.A1(\A[275] ), .A2(\A[276] ), .ZN(new_n1949_));
  AOI21_X1   g00946(.A1(new_n1939_), .A2(new_n1946_), .B(new_n1949_), .ZN(new_n1950_));
  AOI21_X1   g00947(.A1(new_n1928_), .A2(new_n1936_), .B(new_n1934_), .ZN(new_n1951_));
  NAND2_X1   g00948(.A1(new_n1950_), .A2(new_n1951_), .ZN(new_n1952_));
  NAND2_X1   g00949(.A1(new_n1927_), .A2(new_n1912_), .ZN(new_n1954_));
  INV_X1     g00950(.I(new_n1954_), .ZN(new_n1955_));
  NOR2_X1    g00951(.A1(new_n1886_), .A2(new_n1955_), .ZN(new_n1956_));
  AOI21_X1   g00952(.A1(new_n1879_), .A2(new_n1874_), .B(new_n1956_), .ZN(new_n1957_));
  NOR2_X1    g00953(.A1(new_n1883_), .A2(new_n1884_), .ZN(new_n1958_));
  NOR2_X1    g00954(.A1(new_n1881_), .A2(new_n1880_), .ZN(new_n1959_));
  NOR2_X1    g00955(.A1(new_n1958_), .A2(new_n1959_), .ZN(new_n1960_));
  NAND2_X1   g00956(.A1(new_n1960_), .A2(new_n1954_), .ZN(new_n1961_));
  NOR3_X1    g00957(.A1(new_n1869_), .A2(new_n1862_), .A3(new_n1961_), .ZN(new_n1962_));
  INV_X1     g00958(.I(new_n1910_), .ZN(new_n1963_));
  AOI21_X1   g00959(.A1(new_n1919_), .A2(new_n1925_), .B(new_n1963_), .ZN(new_n1964_));
  NOR3_X1    g00960(.A1(new_n1897_), .A2(new_n1907_), .A3(new_n1910_), .ZN(new_n1965_));
  OAI21_X1   g00961(.A1(new_n1964_), .A2(new_n1965_), .B(new_n1909_), .ZN(new_n1966_));
  INV_X1     g00962(.I(new_n1909_), .ZN(new_n1967_));
  OAI21_X1   g00963(.A1(new_n1897_), .A2(new_n1907_), .B(new_n1910_), .ZN(new_n1968_));
  NAND3_X1   g00964(.A1(new_n1919_), .A2(new_n1925_), .A3(new_n1963_), .ZN(new_n1969_));
  NAND3_X1   g00965(.A1(new_n1969_), .A2(new_n1968_), .A3(new_n1967_), .ZN(new_n1970_));
  NAND2_X1   g00966(.A1(new_n1966_), .A2(new_n1970_), .ZN(new_n1971_));
  NOR4_X1    g00967(.A1(new_n1933_), .A2(new_n1937_), .A3(new_n1944_), .A4(new_n1947_), .ZN(new_n1972_));
  NOR2_X1    g00968(.A1(new_n1938_), .A2(new_n1948_), .ZN(new_n1973_));
  NOR2_X1    g00969(.A1(new_n1973_), .A2(new_n1972_), .ZN(new_n1974_));
  NAND3_X1   g00970(.A1(new_n1927_), .A2(new_n1974_), .A3(new_n1912_), .ZN(new_n1975_));
  NAND2_X1   g00971(.A1(new_n1938_), .A2(new_n1948_), .ZN(new_n1976_));
  NAND2_X1   g00972(.A1(new_n1919_), .A2(new_n1907_), .ZN(new_n1977_));
  NAND2_X1   g00973(.A1(new_n1925_), .A2(new_n1897_), .ZN(new_n1978_));
  AOI21_X1   g00974(.A1(new_n1978_), .A2(new_n1977_), .B(new_n1911_), .ZN(new_n1979_));
  NOR3_X1    g00975(.A1(new_n1979_), .A2(new_n1976_), .A3(new_n1952_), .ZN(new_n1980_));
  OAI21_X1   g00976(.A1(new_n1975_), .A2(new_n1971_), .B(new_n1980_), .ZN(new_n1981_));
  INV_X1     g00977(.I(new_n1950_), .ZN(new_n1982_));
  NOR2_X1    g00978(.A1(new_n1931_), .A2(\A[272] ), .ZN(new_n1983_));
  NOR2_X1    g00979(.A1(new_n1929_), .A2(\A[273] ), .ZN(new_n1984_));
  OAI21_X1   g00980(.A1(new_n1983_), .A2(new_n1984_), .B(\A[271] ), .ZN(new_n1985_));
  INV_X1     g00981(.I(new_n1936_), .ZN(new_n1986_));
  OAI21_X1   g00982(.A1(new_n1986_), .A2(new_n1934_), .B(new_n1928_), .ZN(new_n1987_));
  NAND2_X1   g00983(.A1(new_n1985_), .A2(new_n1987_), .ZN(new_n1988_));
  NOR2_X1    g00984(.A1(new_n1942_), .A2(\A[275] ), .ZN(new_n1989_));
  NOR2_X1    g00985(.A1(new_n1940_), .A2(\A[276] ), .ZN(new_n1990_));
  OAI21_X1   g00986(.A1(new_n1989_), .A2(new_n1990_), .B(\A[274] ), .ZN(new_n1991_));
  AND2_X2    g00987(.A1(\A[275] ), .A2(\A[276] ), .Z(new_n1992_));
  OAI21_X1   g00988(.A1(new_n1992_), .A2(new_n1949_), .B(new_n1939_), .ZN(new_n1993_));
  NAND2_X1   g00989(.A1(new_n1991_), .A2(new_n1993_), .ZN(new_n1994_));
  OAI21_X1   g00990(.A1(new_n1988_), .A2(new_n1994_), .B(new_n1951_), .ZN(new_n1995_));
  INV_X1     g00991(.I(new_n1951_), .ZN(new_n1996_));
  NAND3_X1   g00992(.A1(new_n1938_), .A2(new_n1948_), .A3(new_n1996_), .ZN(new_n1997_));
  AOI21_X1   g00993(.A1(new_n1995_), .A2(new_n1997_), .B(new_n1982_), .ZN(new_n1998_));
  NOR2_X1    g00994(.A1(new_n1972_), .A2(new_n1996_), .ZN(new_n1999_));
  NOR3_X1    g00995(.A1(new_n1988_), .A2(new_n1994_), .A3(new_n1951_), .ZN(new_n2000_));
  NOR3_X1    g00996(.A1(new_n1999_), .A2(new_n1950_), .A3(new_n2000_), .ZN(new_n2001_));
  NOR2_X1    g00997(.A1(new_n2001_), .A2(new_n1998_), .ZN(new_n2002_));
  NOR2_X1    g00998(.A1(new_n1981_), .A2(new_n2002_), .ZN(new_n2003_));
  OAI21_X1   g00999(.A1(new_n1999_), .A2(new_n2000_), .B(new_n1950_), .ZN(new_n2004_));
  NAND3_X1   g01000(.A1(new_n1995_), .A2(new_n1997_), .A3(new_n1982_), .ZN(new_n2005_));
  NAND2_X1   g01001(.A1(new_n2004_), .A2(new_n2005_), .ZN(new_n2006_));
  NOR3_X1    g01002(.A1(new_n1988_), .A2(new_n1994_), .A3(new_n1952_), .ZN(new_n2007_));
  NAND4_X1   g01003(.A1(new_n1927_), .A2(new_n1974_), .A3(new_n1912_), .A4(new_n2007_), .ZN(new_n2008_));
  NAND2_X1   g01004(.A1(new_n2006_), .A2(new_n2008_), .ZN(new_n2009_));
  INV_X1     g01005(.I(new_n1911_), .ZN(new_n2010_));
  NOR2_X1    g01006(.A1(new_n1925_), .A2(new_n1897_), .ZN(new_n2011_));
  NOR2_X1    g01007(.A1(new_n1919_), .A2(new_n1907_), .ZN(new_n2012_));
  OAI21_X1   g01008(.A1(new_n2011_), .A2(new_n2012_), .B(new_n2010_), .ZN(new_n2013_));
  NAND3_X1   g01009(.A1(new_n1966_), .A2(new_n1970_), .A3(new_n2013_), .ZN(new_n2014_));
  OAI21_X1   g01010(.A1(new_n2006_), .A2(new_n2008_), .B(new_n2014_), .ZN(new_n2015_));
  AOI21_X1   g01011(.A1(new_n1969_), .A2(new_n1968_), .B(new_n1967_), .ZN(new_n2016_));
  NOR3_X1    g01012(.A1(new_n1964_), .A2(new_n1965_), .A3(new_n1909_), .ZN(new_n2017_));
  NOR3_X1    g01013(.A1(new_n2017_), .A2(new_n2016_), .A3(new_n1979_), .ZN(new_n2018_));
  NAND2_X1   g01014(.A1(new_n1919_), .A2(new_n1925_), .ZN(new_n2019_));
  NAND2_X1   g01015(.A1(new_n1897_), .A2(new_n1907_), .ZN(new_n2020_));
  NAND3_X1   g01016(.A1(new_n1912_), .A2(new_n2019_), .A3(new_n2020_), .ZN(new_n2021_));
  NAND2_X1   g01017(.A1(new_n1988_), .A2(new_n1994_), .ZN(new_n2022_));
  NAND3_X1   g01018(.A1(new_n2007_), .A2(new_n1976_), .A3(new_n2022_), .ZN(new_n2023_));
  NOR4_X1    g01019(.A1(new_n2021_), .A2(new_n2001_), .A3(new_n1998_), .A4(new_n2023_), .ZN(new_n2024_));
  NAND2_X1   g01020(.A1(new_n2024_), .A2(new_n2018_), .ZN(new_n2025_));
  NAND2_X1   g01021(.A1(new_n2015_), .A2(new_n2025_), .ZN(new_n2026_));
  AOI21_X1   g01022(.A1(new_n2026_), .A2(new_n2009_), .B(new_n2003_), .ZN(new_n2027_));
  OAI22_X1   g01023(.A1(new_n1957_), .A2(new_n1962_), .B1(new_n2027_), .B2(new_n1870_), .ZN(new_n2028_));
  AOI21_X1   g01024(.A1(new_n1853_), .A2(new_n1846_), .B(new_n1871_), .ZN(new_n2029_));
  NOR2_X1    g01025(.A1(new_n1789_), .A2(new_n1793_), .ZN(new_n2030_));
  OAI21_X1   g01026(.A1(new_n1827_), .A2(new_n2030_), .B(new_n1794_), .ZN(new_n2031_));
  NAND2_X1   g01027(.A1(new_n1747_), .A2(new_n1768_), .ZN(new_n2032_));
  AOI21_X1   g01028(.A1(new_n1779_), .A2(new_n2032_), .B(new_n1844_), .ZN(new_n2033_));
  XOR2_X1    g01029(.A1(new_n2033_), .A2(new_n2031_), .Z(new_n2034_));
  INV_X1     g01030(.I(new_n2034_), .ZN(new_n2035_));
  NOR3_X1    g01031(.A1(new_n2029_), .A2(new_n1868_), .A3(new_n2035_), .ZN(new_n2036_));
  OAI21_X1   g01032(.A1(new_n2018_), .A2(new_n2008_), .B(new_n2006_), .ZN(new_n2037_));
  NOR2_X1    g01033(.A1(new_n1909_), .A2(new_n1910_), .ZN(new_n2038_));
  OAI21_X1   g01034(.A1(new_n2019_), .A2(new_n2038_), .B(new_n1911_), .ZN(new_n2039_));
  NOR2_X1    g01035(.A1(new_n1950_), .A2(new_n1951_), .ZN(new_n2040_));
  OAI21_X1   g01036(.A1(new_n1976_), .A2(new_n2040_), .B(new_n1952_), .ZN(new_n2041_));
  XNOR2_X1   g01037(.A1(new_n2039_), .A2(new_n2041_), .ZN(new_n2042_));
  NAND3_X1   g01038(.A1(new_n1981_), .A2(new_n2037_), .A3(new_n2042_), .ZN(new_n2043_));
  XOR2_X1    g01039(.A1(new_n2036_), .A2(new_n2043_), .Z(new_n2044_));
  NOR2_X1    g01040(.A1(new_n2044_), .A2(new_n2028_), .ZN(new_n2045_));
  NAND2_X1   g01041(.A1(new_n1879_), .A2(new_n1874_), .ZN(new_n2046_));
  OAI21_X1   g01042(.A1(new_n1869_), .A2(new_n1862_), .B(new_n1961_), .ZN(new_n2047_));
  NAND3_X1   g01043(.A1(new_n1879_), .A2(new_n1874_), .A3(new_n1956_), .ZN(new_n2048_));
  NOR2_X1    g01044(.A1(new_n2017_), .A2(new_n2016_), .ZN(new_n2049_));
  NOR3_X1    g01045(.A1(new_n2021_), .A2(new_n1972_), .A3(new_n1973_), .ZN(new_n2050_));
  NAND2_X1   g01046(.A1(new_n2013_), .A2(new_n2007_), .ZN(new_n2051_));
  AOI21_X1   g01047(.A1(new_n2049_), .A2(new_n2050_), .B(new_n2051_), .ZN(new_n2052_));
  NAND2_X1   g01048(.A1(new_n2052_), .A2(new_n2006_), .ZN(new_n2053_));
  NOR2_X1    g01049(.A1(new_n2024_), .A2(new_n2018_), .ZN(new_n2054_));
  NOR3_X1    g01050(.A1(new_n2014_), .A2(new_n2006_), .A3(new_n2008_), .ZN(new_n2055_));
  OAI21_X1   g01051(.A1(new_n2054_), .A2(new_n2055_), .B(new_n2009_), .ZN(new_n2056_));
  NAND2_X1   g01052(.A1(new_n2056_), .A2(new_n2053_), .ZN(new_n2057_));
  AOI22_X1   g01053(.A1(new_n2047_), .A2(new_n2048_), .B1(new_n2057_), .B2(new_n2046_), .ZN(new_n2058_));
  INV_X1     g01054(.I(new_n2043_), .ZN(new_n2059_));
  NOR2_X1    g01055(.A1(new_n2059_), .A2(new_n2036_), .ZN(new_n2060_));
  NAND2_X1   g01056(.A1(new_n1875_), .A2(new_n1785_), .ZN(new_n2061_));
  NAND3_X1   g01057(.A1(new_n2061_), .A2(new_n1878_), .A3(new_n2034_), .ZN(new_n2062_));
  NOR2_X1    g01058(.A1(new_n2062_), .A2(new_n2043_), .ZN(new_n2063_));
  NOR2_X1    g01059(.A1(new_n2060_), .A2(new_n2063_), .ZN(new_n2064_));
  NOR2_X1    g01060(.A1(new_n2064_), .A2(new_n2058_), .ZN(new_n2065_));
  INV_X1     g01061(.I(\A[310] ), .ZN(new_n2066_));
  NOR2_X1    g01062(.A1(\A[311] ), .A2(\A[312] ), .ZN(new_n2067_));
  NAND2_X1   g01063(.A1(\A[311] ), .A2(\A[312] ), .ZN(new_n2068_));
  AOI21_X1   g01064(.A1(new_n2066_), .A2(new_n2068_), .B(new_n2067_), .ZN(new_n2069_));
  INV_X1     g01065(.I(\A[307] ), .ZN(new_n2070_));
  NOR2_X1    g01066(.A1(\A[308] ), .A2(\A[309] ), .ZN(new_n2071_));
  NAND2_X1   g01067(.A1(\A[308] ), .A2(\A[309] ), .ZN(new_n2072_));
  AOI21_X1   g01068(.A1(new_n2070_), .A2(new_n2072_), .B(new_n2071_), .ZN(new_n2073_));
  INV_X1     g01069(.I(new_n2073_), .ZN(new_n2074_));
  INV_X1     g01070(.I(\A[308] ), .ZN(new_n2075_));
  NAND2_X1   g01071(.A1(new_n2075_), .A2(\A[309] ), .ZN(new_n2076_));
  INV_X1     g01072(.I(\A[309] ), .ZN(new_n2077_));
  NAND2_X1   g01073(.A1(new_n2077_), .A2(\A[308] ), .ZN(new_n2078_));
  AOI21_X1   g01074(.A1(new_n2076_), .A2(new_n2078_), .B(new_n2070_), .ZN(new_n2079_));
  INV_X1     g01075(.I(new_n2071_), .ZN(new_n2080_));
  AOI21_X1   g01076(.A1(new_n2080_), .A2(new_n2072_), .B(\A[307] ), .ZN(new_n2081_));
  INV_X1     g01077(.I(\A[311] ), .ZN(new_n2082_));
  NAND2_X1   g01078(.A1(new_n2082_), .A2(\A[312] ), .ZN(new_n2083_));
  INV_X1     g01079(.I(\A[312] ), .ZN(new_n2084_));
  NAND2_X1   g01080(.A1(new_n2084_), .A2(\A[311] ), .ZN(new_n2085_));
  AOI21_X1   g01081(.A1(new_n2083_), .A2(new_n2085_), .B(new_n2066_), .ZN(new_n2086_));
  INV_X1     g01082(.I(new_n2067_), .ZN(new_n2087_));
  AOI21_X1   g01083(.A1(new_n2087_), .A2(new_n2068_), .B(\A[310] ), .ZN(new_n2088_));
  NOR4_X1    g01084(.A1(new_n2079_), .A2(new_n2081_), .A3(new_n2088_), .A4(new_n2086_), .ZN(new_n2089_));
  NOR2_X1    g01085(.A1(new_n2089_), .A2(new_n2074_), .ZN(new_n2090_));
  NOR2_X1    g01086(.A1(new_n2077_), .A2(\A[308] ), .ZN(new_n2091_));
  NOR2_X1    g01087(.A1(new_n2075_), .A2(\A[309] ), .ZN(new_n2092_));
  OAI21_X1   g01088(.A1(new_n2091_), .A2(new_n2092_), .B(\A[307] ), .ZN(new_n2093_));
  INV_X1     g01089(.I(new_n2072_), .ZN(new_n2094_));
  OAI21_X1   g01090(.A1(new_n2094_), .A2(new_n2071_), .B(new_n2070_), .ZN(new_n2095_));
  NAND2_X1   g01091(.A1(new_n2093_), .A2(new_n2095_), .ZN(new_n2096_));
  NOR2_X1    g01092(.A1(new_n2084_), .A2(\A[311] ), .ZN(new_n2097_));
  NOR2_X1    g01093(.A1(new_n2082_), .A2(\A[312] ), .ZN(new_n2098_));
  OAI21_X1   g01094(.A1(new_n2097_), .A2(new_n2098_), .B(\A[310] ), .ZN(new_n2099_));
  INV_X1     g01095(.I(new_n2068_), .ZN(new_n2100_));
  OAI21_X1   g01096(.A1(new_n2100_), .A2(new_n2067_), .B(new_n2066_), .ZN(new_n2101_));
  NAND2_X1   g01097(.A1(new_n2099_), .A2(new_n2101_), .ZN(new_n2102_));
  NOR3_X1    g01098(.A1(new_n2096_), .A2(new_n2102_), .A3(new_n2073_), .ZN(new_n2103_));
  OAI21_X1   g01099(.A1(new_n2090_), .A2(new_n2103_), .B(new_n2069_), .ZN(new_n2104_));
  INV_X1     g01100(.I(new_n2069_), .ZN(new_n2105_));
  OAI21_X1   g01101(.A1(new_n2096_), .A2(new_n2102_), .B(new_n2073_), .ZN(new_n2106_));
  NOR2_X1    g01102(.A1(new_n2081_), .A2(new_n2079_), .ZN(new_n2107_));
  NOR2_X1    g01103(.A1(new_n2088_), .A2(new_n2086_), .ZN(new_n2108_));
  NAND3_X1   g01104(.A1(new_n2107_), .A2(new_n2108_), .A3(new_n2074_), .ZN(new_n2109_));
  NAND3_X1   g01105(.A1(new_n2106_), .A2(new_n2109_), .A3(new_n2105_), .ZN(new_n2110_));
  NAND2_X1   g01106(.A1(new_n2104_), .A2(new_n2110_), .ZN(new_n2111_));
  INV_X1     g01107(.I(\A[316] ), .ZN(new_n2112_));
  NOR2_X1    g01108(.A1(\A[317] ), .A2(\A[318] ), .ZN(new_n2113_));
  NAND2_X1   g01109(.A1(\A[317] ), .A2(\A[318] ), .ZN(new_n2114_));
  AOI21_X1   g01110(.A1(new_n2112_), .A2(new_n2114_), .B(new_n2113_), .ZN(new_n2115_));
  INV_X1     g01111(.I(\A[313] ), .ZN(new_n2116_));
  NOR2_X1    g01112(.A1(\A[314] ), .A2(\A[315] ), .ZN(new_n2117_));
  NAND2_X1   g01113(.A1(\A[314] ), .A2(\A[315] ), .ZN(new_n2118_));
  AOI21_X1   g01114(.A1(new_n2116_), .A2(new_n2118_), .B(new_n2117_), .ZN(new_n2119_));
  NAND2_X1   g01115(.A1(new_n2115_), .A2(new_n2119_), .ZN(new_n2120_));
  INV_X1     g01116(.I(\A[314] ), .ZN(new_n2121_));
  NAND2_X1   g01117(.A1(new_n2121_), .A2(\A[315] ), .ZN(new_n2122_));
  INV_X1     g01118(.I(\A[315] ), .ZN(new_n2123_));
  NAND2_X1   g01119(.A1(new_n2123_), .A2(\A[314] ), .ZN(new_n2124_));
  AOI21_X1   g01120(.A1(new_n2122_), .A2(new_n2124_), .B(new_n2116_), .ZN(new_n2125_));
  INV_X1     g01121(.I(new_n2117_), .ZN(new_n2126_));
  AOI21_X1   g01122(.A1(new_n2126_), .A2(new_n2118_), .B(\A[313] ), .ZN(new_n2127_));
  NOR2_X1    g01123(.A1(new_n2127_), .A2(new_n2125_), .ZN(new_n2128_));
  INV_X1     g01124(.I(\A[318] ), .ZN(new_n2129_));
  NOR2_X1    g01125(.A1(new_n2129_), .A2(\A[317] ), .ZN(new_n2130_));
  INV_X1     g01126(.I(\A[317] ), .ZN(new_n2131_));
  NOR2_X1    g01127(.A1(new_n2131_), .A2(\A[318] ), .ZN(new_n2132_));
  OAI21_X1   g01128(.A1(new_n2130_), .A2(new_n2132_), .B(\A[316] ), .ZN(new_n2133_));
  AND2_X2    g01129(.A1(\A[317] ), .A2(\A[318] ), .Z(new_n2134_));
  OAI21_X1   g01130(.A1(new_n2134_), .A2(new_n2113_), .B(new_n2112_), .ZN(new_n2135_));
  NAND2_X1   g01131(.A1(new_n2133_), .A2(new_n2135_), .ZN(new_n2136_));
  NAND2_X1   g01132(.A1(new_n2128_), .A2(new_n2136_), .ZN(new_n2137_));
  NOR2_X1    g01133(.A1(new_n2123_), .A2(\A[314] ), .ZN(new_n2138_));
  NOR2_X1    g01134(.A1(new_n2121_), .A2(\A[315] ), .ZN(new_n2139_));
  OAI21_X1   g01135(.A1(new_n2138_), .A2(new_n2139_), .B(\A[313] ), .ZN(new_n2140_));
  AND2_X2    g01136(.A1(\A[314] ), .A2(\A[315] ), .Z(new_n2141_));
  OAI21_X1   g01137(.A1(new_n2141_), .A2(new_n2117_), .B(new_n2116_), .ZN(new_n2142_));
  NAND2_X1   g01138(.A1(new_n2140_), .A2(new_n2142_), .ZN(new_n2143_));
  NAND2_X1   g01139(.A1(new_n2131_), .A2(\A[318] ), .ZN(new_n2144_));
  NAND2_X1   g01140(.A1(new_n2129_), .A2(\A[317] ), .ZN(new_n2145_));
  AOI21_X1   g01141(.A1(new_n2144_), .A2(new_n2145_), .B(new_n2112_), .ZN(new_n2146_));
  OR2_X2     g01142(.A1(\A[317] ), .A2(\A[318] ), .Z(new_n2147_));
  AOI21_X1   g01143(.A1(new_n2147_), .A2(new_n2114_), .B(\A[316] ), .ZN(new_n2148_));
  NOR2_X1    g01144(.A1(new_n2146_), .A2(new_n2148_), .ZN(new_n2149_));
  NAND2_X1   g01145(.A1(new_n2149_), .A2(new_n2143_), .ZN(new_n2150_));
  AOI21_X1   g01146(.A1(new_n2137_), .A2(new_n2150_), .B(new_n2120_), .ZN(new_n2151_));
  INV_X1     g01147(.I(new_n2115_), .ZN(new_n2152_));
  NAND4_X1   g01148(.A1(new_n2140_), .A2(new_n2133_), .A3(new_n2142_), .A4(new_n2135_), .ZN(new_n2153_));
  NAND2_X1   g01149(.A1(new_n2153_), .A2(new_n2119_), .ZN(new_n2154_));
  INV_X1     g01150(.I(new_n2119_), .ZN(new_n2155_));
  NAND3_X1   g01151(.A1(new_n2128_), .A2(new_n2149_), .A3(new_n2155_), .ZN(new_n2156_));
  AOI21_X1   g01152(.A1(new_n2154_), .A2(new_n2156_), .B(new_n2152_), .ZN(new_n2157_));
  AOI21_X1   g01153(.A1(new_n2128_), .A2(new_n2149_), .B(new_n2155_), .ZN(new_n2158_));
  NOR3_X1    g01154(.A1(new_n2143_), .A2(new_n2136_), .A3(new_n2119_), .ZN(new_n2159_));
  NOR3_X1    g01155(.A1(new_n2158_), .A2(new_n2159_), .A3(new_n2115_), .ZN(new_n2160_));
  NOR3_X1    g01156(.A1(new_n2157_), .A2(new_n2160_), .A3(new_n2151_), .ZN(new_n2161_));
  INV_X1     g01157(.I(new_n2120_), .ZN(new_n2162_));
  NOR4_X1    g01158(.A1(new_n2125_), .A2(new_n2127_), .A3(new_n2146_), .A4(new_n2148_), .ZN(new_n2163_));
  NAND2_X1   g01159(.A1(new_n2163_), .A2(new_n2162_), .ZN(new_n2164_));
  AOI22_X1   g01160(.A1(new_n2140_), .A2(new_n2142_), .B1(new_n2133_), .B2(new_n2135_), .ZN(new_n2165_));
  OR2_X2     g01161(.A1(new_n2165_), .A2(new_n2163_), .Z(new_n2166_));
  NAND4_X1   g01162(.A1(new_n2093_), .A2(new_n2095_), .A3(new_n2099_), .A4(new_n2101_), .ZN(new_n2167_));
  NAND2_X1   g01163(.A1(new_n2096_), .A2(new_n2102_), .ZN(new_n2168_));
  NAND2_X1   g01164(.A1(new_n2168_), .A2(new_n2167_), .ZN(new_n2169_));
  NAND2_X1   g01165(.A1(new_n2069_), .A2(new_n2073_), .ZN(new_n2170_));
  INV_X1     g01166(.I(new_n2170_), .ZN(new_n2171_));
  NAND2_X1   g01167(.A1(new_n2089_), .A2(new_n2171_), .ZN(new_n2172_));
  NOR4_X1    g01168(.A1(new_n2166_), .A2(new_n2169_), .A3(new_n2172_), .A4(new_n2164_), .ZN(new_n2173_));
  NAND2_X1   g01169(.A1(new_n2161_), .A2(new_n2173_), .ZN(new_n2174_));
  NOR2_X1    g01170(.A1(new_n2149_), .A2(new_n2143_), .ZN(new_n2175_));
  NOR2_X1    g01171(.A1(new_n2128_), .A2(new_n2136_), .ZN(new_n2176_));
  OAI21_X1   g01172(.A1(new_n2175_), .A2(new_n2176_), .B(new_n2162_), .ZN(new_n2177_));
  OAI21_X1   g01173(.A1(new_n2158_), .A2(new_n2159_), .B(new_n2115_), .ZN(new_n2178_));
  NAND3_X1   g01174(.A1(new_n2154_), .A2(new_n2156_), .A3(new_n2152_), .ZN(new_n2179_));
  NAND3_X1   g01175(.A1(new_n2178_), .A2(new_n2179_), .A3(new_n2177_), .ZN(new_n2180_));
  NOR2_X1    g01176(.A1(new_n2153_), .A2(new_n2120_), .ZN(new_n2181_));
  NOR2_X1    g01177(.A1(new_n2165_), .A2(new_n2163_), .ZN(new_n2182_));
  AOI22_X1   g01178(.A1(new_n2093_), .A2(new_n2095_), .B1(new_n2099_), .B2(new_n2101_), .ZN(new_n2183_));
  NOR2_X1    g01179(.A1(new_n2183_), .A2(new_n2089_), .ZN(new_n2184_));
  NOR2_X1    g01180(.A1(new_n2167_), .A2(new_n2170_), .ZN(new_n2185_));
  NAND4_X1   g01181(.A1(new_n2184_), .A2(new_n2182_), .A3(new_n2185_), .A4(new_n2181_), .ZN(new_n2186_));
  NAND2_X1   g01182(.A1(new_n2180_), .A2(new_n2186_), .ZN(new_n2187_));
  AOI21_X1   g01183(.A1(new_n2174_), .A2(new_n2187_), .B(new_n2111_), .ZN(new_n2188_));
  NOR2_X1    g01184(.A1(new_n2161_), .A2(new_n2186_), .ZN(new_n2189_));
  NOR2_X1    g01185(.A1(new_n2157_), .A2(new_n2160_), .ZN(new_n2190_));
  NAND3_X1   g01186(.A1(new_n2184_), .A2(new_n2182_), .A3(new_n2181_), .ZN(new_n2191_));
  INV_X1     g01187(.I(new_n2191_), .ZN(new_n2192_));
  NAND2_X1   g01188(.A1(new_n2177_), .A2(new_n2185_), .ZN(new_n2193_));
  AOI21_X1   g01189(.A1(new_n2192_), .A2(new_n2190_), .B(new_n2193_), .ZN(new_n2194_));
  NOR3_X1    g01190(.A1(new_n2194_), .A2(new_n2189_), .A3(new_n2111_), .ZN(new_n2195_));
  NOR2_X1    g01191(.A1(new_n2195_), .A2(new_n2188_), .ZN(new_n2196_));
  AOI21_X1   g01192(.A1(new_n2106_), .A2(new_n2109_), .B(new_n2105_), .ZN(new_n2197_));
  NOR3_X1    g01193(.A1(new_n2090_), .A2(new_n2103_), .A3(new_n2069_), .ZN(new_n2198_));
  NOR2_X1    g01194(.A1(new_n2198_), .A2(new_n2197_), .ZN(new_n2199_));
  NOR4_X1    g01195(.A1(new_n2186_), .A2(new_n2151_), .A3(new_n2157_), .A4(new_n2160_), .ZN(new_n2200_));
  NOR2_X1    g01196(.A1(new_n2161_), .A2(new_n2173_), .ZN(new_n2201_));
  OAI21_X1   g01197(.A1(new_n2201_), .A2(new_n2200_), .B(new_n2199_), .ZN(new_n2202_));
  NAND2_X1   g01198(.A1(new_n2180_), .A2(new_n2173_), .ZN(new_n2203_));
  NAND2_X1   g01199(.A1(new_n2178_), .A2(new_n2179_), .ZN(new_n2204_));
  NOR2_X1    g01200(.A1(new_n2151_), .A2(new_n2172_), .ZN(new_n2205_));
  OAI21_X1   g01201(.A1(new_n2204_), .A2(new_n2191_), .B(new_n2205_), .ZN(new_n2206_));
  NAND3_X1   g01202(.A1(new_n2206_), .A2(new_n2203_), .A3(new_n2199_), .ZN(new_n2207_));
  NAND2_X1   g01203(.A1(new_n2182_), .A2(new_n2181_), .ZN(new_n2208_));
  INV_X1     g01204(.I(new_n2208_), .ZN(new_n2209_));
  NAND2_X1   g01205(.A1(new_n2184_), .A2(new_n2185_), .ZN(new_n2210_));
  NOR2_X1    g01206(.A1(new_n2209_), .A2(new_n2210_), .ZN(new_n2211_));
  INV_X1     g01207(.I(new_n2210_), .ZN(new_n2212_));
  NOR2_X1    g01208(.A1(new_n2212_), .A2(new_n2208_), .ZN(new_n2213_));
  INV_X1     g01209(.I(\A[303] ), .ZN(new_n2214_));
  NOR2_X1    g01210(.A1(new_n2214_), .A2(\A[302] ), .ZN(new_n2215_));
  INV_X1     g01211(.I(\A[302] ), .ZN(new_n2216_));
  NOR2_X1    g01212(.A1(new_n2216_), .A2(\A[303] ), .ZN(new_n2217_));
  OAI21_X1   g01213(.A1(new_n2215_), .A2(new_n2217_), .B(\A[301] ), .ZN(new_n2218_));
  INV_X1     g01214(.I(\A[301] ), .ZN(new_n2219_));
  NOR2_X1    g01215(.A1(\A[302] ), .A2(\A[303] ), .ZN(new_n2220_));
  AND2_X2    g01216(.A1(\A[302] ), .A2(\A[303] ), .Z(new_n2221_));
  OAI21_X1   g01217(.A1(new_n2221_), .A2(new_n2220_), .B(new_n2219_), .ZN(new_n2222_));
  NAND2_X1   g01218(.A1(new_n2218_), .A2(new_n2222_), .ZN(new_n2223_));
  INV_X1     g01219(.I(\A[306] ), .ZN(new_n2224_));
  NOR2_X1    g01220(.A1(new_n2224_), .A2(\A[305] ), .ZN(new_n2225_));
  INV_X1     g01221(.I(\A[305] ), .ZN(new_n2226_));
  NOR2_X1    g01222(.A1(new_n2226_), .A2(\A[306] ), .ZN(new_n2227_));
  OAI21_X1   g01223(.A1(new_n2225_), .A2(new_n2227_), .B(\A[304] ), .ZN(new_n2228_));
  INV_X1     g01224(.I(\A[304] ), .ZN(new_n2229_));
  NOR2_X1    g01225(.A1(\A[305] ), .A2(\A[306] ), .ZN(new_n2230_));
  AND2_X2    g01226(.A1(\A[305] ), .A2(\A[306] ), .Z(new_n2231_));
  OAI21_X1   g01227(.A1(new_n2231_), .A2(new_n2230_), .B(new_n2229_), .ZN(new_n2232_));
  NAND2_X1   g01228(.A1(new_n2228_), .A2(new_n2232_), .ZN(new_n2233_));
  NAND2_X1   g01229(.A1(\A[305] ), .A2(\A[306] ), .ZN(new_n2234_));
  AOI21_X1   g01230(.A1(new_n2229_), .A2(new_n2234_), .B(new_n2230_), .ZN(new_n2235_));
  NAND2_X1   g01231(.A1(\A[302] ), .A2(\A[303] ), .ZN(new_n2236_));
  AOI21_X1   g01232(.A1(new_n2219_), .A2(new_n2236_), .B(new_n2220_), .ZN(new_n2237_));
  NAND2_X1   g01233(.A1(new_n2235_), .A2(new_n2237_), .ZN(new_n2238_));
  NOR3_X1    g01234(.A1(new_n2223_), .A2(new_n2233_), .A3(new_n2238_), .ZN(new_n2239_));
  NOR2_X1    g01235(.A1(new_n2223_), .A2(new_n2233_), .ZN(new_n2240_));
  NAND2_X1   g01236(.A1(new_n2216_), .A2(\A[303] ), .ZN(new_n2241_));
  NAND2_X1   g01237(.A1(new_n2214_), .A2(\A[302] ), .ZN(new_n2242_));
  AOI21_X1   g01238(.A1(new_n2241_), .A2(new_n2242_), .B(new_n2219_), .ZN(new_n2243_));
  INV_X1     g01239(.I(new_n2220_), .ZN(new_n2244_));
  AOI21_X1   g01240(.A1(new_n2244_), .A2(new_n2236_), .B(\A[301] ), .ZN(new_n2245_));
  NOR2_X1    g01241(.A1(new_n2245_), .A2(new_n2243_), .ZN(new_n2246_));
  NAND2_X1   g01242(.A1(new_n2226_), .A2(\A[306] ), .ZN(new_n2247_));
  NAND2_X1   g01243(.A1(new_n2224_), .A2(\A[305] ), .ZN(new_n2248_));
  AOI21_X1   g01244(.A1(new_n2247_), .A2(new_n2248_), .B(new_n2229_), .ZN(new_n2249_));
  OR2_X2     g01245(.A1(\A[305] ), .A2(\A[306] ), .Z(new_n2250_));
  AOI21_X1   g01246(.A1(new_n2250_), .A2(new_n2234_), .B(\A[304] ), .ZN(new_n2251_));
  NOR2_X1    g01247(.A1(new_n2249_), .A2(new_n2251_), .ZN(new_n2252_));
  NOR2_X1    g01248(.A1(new_n2246_), .A2(new_n2252_), .ZN(new_n2253_));
  NOR2_X1    g01249(.A1(new_n2253_), .A2(new_n2240_), .ZN(new_n2254_));
  INV_X1     g01250(.I(\A[295] ), .ZN(new_n2255_));
  INV_X1     g01251(.I(\A[296] ), .ZN(new_n2256_));
  NAND2_X1   g01252(.A1(new_n2256_), .A2(\A[297] ), .ZN(new_n2257_));
  INV_X1     g01253(.I(\A[297] ), .ZN(new_n2258_));
  NAND2_X1   g01254(.A1(new_n2258_), .A2(\A[296] ), .ZN(new_n2259_));
  AOI21_X1   g01255(.A1(new_n2257_), .A2(new_n2259_), .B(new_n2255_), .ZN(new_n2260_));
  NOR2_X1    g01256(.A1(\A[296] ), .A2(\A[297] ), .ZN(new_n2261_));
  INV_X1     g01257(.I(new_n2261_), .ZN(new_n2262_));
  NAND2_X1   g01258(.A1(\A[296] ), .A2(\A[297] ), .ZN(new_n2263_));
  AOI21_X1   g01259(.A1(new_n2262_), .A2(new_n2263_), .B(\A[295] ), .ZN(new_n2264_));
  NOR2_X1    g01260(.A1(new_n2264_), .A2(new_n2260_), .ZN(new_n2265_));
  INV_X1     g01261(.I(\A[298] ), .ZN(new_n2266_));
  INV_X1     g01262(.I(\A[299] ), .ZN(new_n2267_));
  NAND2_X1   g01263(.A1(new_n2267_), .A2(\A[300] ), .ZN(new_n2268_));
  INV_X1     g01264(.I(\A[300] ), .ZN(new_n2269_));
  NAND2_X1   g01265(.A1(new_n2269_), .A2(\A[299] ), .ZN(new_n2270_));
  AOI21_X1   g01266(.A1(new_n2268_), .A2(new_n2270_), .B(new_n2266_), .ZN(new_n2271_));
  OR2_X2     g01267(.A1(\A[299] ), .A2(\A[300] ), .Z(new_n2272_));
  NAND2_X1   g01268(.A1(\A[299] ), .A2(\A[300] ), .ZN(new_n2273_));
  AOI21_X1   g01269(.A1(new_n2272_), .A2(new_n2273_), .B(\A[298] ), .ZN(new_n2274_));
  NOR2_X1    g01270(.A1(new_n2271_), .A2(new_n2274_), .ZN(new_n2275_));
  NOR2_X1    g01271(.A1(\A[299] ), .A2(\A[300] ), .ZN(new_n2276_));
  AOI21_X1   g01272(.A1(new_n2266_), .A2(new_n2273_), .B(new_n2276_), .ZN(new_n2277_));
  AOI21_X1   g01273(.A1(new_n2255_), .A2(new_n2263_), .B(new_n2261_), .ZN(new_n2278_));
  NAND2_X1   g01274(.A1(new_n2277_), .A2(new_n2278_), .ZN(new_n2279_));
  INV_X1     g01275(.I(new_n2279_), .ZN(new_n2280_));
  NAND2_X1   g01276(.A1(new_n2254_), .A2(new_n2239_), .ZN(new_n2281_));
  INV_X1     g01277(.I(new_n2281_), .ZN(new_n2282_));
  NOR3_X1    g01278(.A1(new_n2213_), .A2(new_n2211_), .A3(new_n2282_), .ZN(new_n2283_));
  AOI21_X1   g01279(.A1(new_n2207_), .A2(new_n2202_), .B(new_n2283_), .ZN(new_n2284_));
  NAND2_X1   g01280(.A1(new_n2212_), .A2(new_n2208_), .ZN(new_n2285_));
  NAND2_X1   g01281(.A1(new_n2209_), .A2(new_n2210_), .ZN(new_n2286_));
  NAND3_X1   g01282(.A1(new_n2285_), .A2(new_n2286_), .A3(new_n2281_), .ZN(new_n2287_));
  NOR3_X1    g01283(.A1(new_n2195_), .A2(new_n2188_), .A3(new_n2287_), .ZN(new_n2288_));
  INV_X1     g01284(.I(new_n2237_), .ZN(new_n2289_));
  AOI21_X1   g01285(.A1(new_n2246_), .A2(new_n2252_), .B(new_n2289_), .ZN(new_n2290_));
  NOR3_X1    g01286(.A1(new_n2223_), .A2(new_n2233_), .A3(new_n2237_), .ZN(new_n2291_));
  OAI21_X1   g01287(.A1(new_n2290_), .A2(new_n2291_), .B(new_n2235_), .ZN(new_n2292_));
  INV_X1     g01288(.I(new_n2235_), .ZN(new_n2293_));
  OAI21_X1   g01289(.A1(new_n2223_), .A2(new_n2233_), .B(new_n2237_), .ZN(new_n2294_));
  NAND3_X1   g01290(.A1(new_n2246_), .A2(new_n2252_), .A3(new_n2289_), .ZN(new_n2295_));
  NAND3_X1   g01291(.A1(new_n2294_), .A2(new_n2295_), .A3(new_n2293_), .ZN(new_n2296_));
  NAND2_X1   g01292(.A1(new_n2292_), .A2(new_n2296_), .ZN(new_n2297_));
  NOR4_X1    g01293(.A1(new_n2260_), .A2(new_n2264_), .A3(new_n2271_), .A4(new_n2274_), .ZN(new_n2298_));
  NOR2_X1    g01294(.A1(new_n2265_), .A2(new_n2275_), .ZN(new_n2299_));
  NOR2_X1    g01295(.A1(new_n2299_), .A2(new_n2298_), .ZN(new_n2300_));
  NAND3_X1   g01296(.A1(new_n2254_), .A2(new_n2300_), .A3(new_n2239_), .ZN(new_n2301_));
  NAND2_X1   g01297(.A1(new_n2265_), .A2(new_n2275_), .ZN(new_n2302_));
  NAND2_X1   g01298(.A1(new_n2246_), .A2(new_n2233_), .ZN(new_n2303_));
  NAND2_X1   g01299(.A1(new_n2252_), .A2(new_n2223_), .ZN(new_n2304_));
  AOI21_X1   g01300(.A1(new_n2303_), .A2(new_n2304_), .B(new_n2238_), .ZN(new_n2305_));
  NOR3_X1    g01301(.A1(new_n2305_), .A2(new_n2302_), .A3(new_n2279_), .ZN(new_n2306_));
  OAI21_X1   g01302(.A1(new_n2301_), .A2(new_n2297_), .B(new_n2306_), .ZN(new_n2307_));
  INV_X1     g01303(.I(new_n2277_), .ZN(new_n2308_));
  NOR2_X1    g01304(.A1(new_n2258_), .A2(\A[296] ), .ZN(new_n2309_));
  NOR2_X1    g01305(.A1(new_n2256_), .A2(\A[297] ), .ZN(new_n2310_));
  OAI21_X1   g01306(.A1(new_n2309_), .A2(new_n2310_), .B(\A[295] ), .ZN(new_n2311_));
  INV_X1     g01307(.I(new_n2263_), .ZN(new_n2312_));
  OAI21_X1   g01308(.A1(new_n2312_), .A2(new_n2261_), .B(new_n2255_), .ZN(new_n2313_));
  NAND2_X1   g01309(.A1(new_n2311_), .A2(new_n2313_), .ZN(new_n2314_));
  NOR2_X1    g01310(.A1(new_n2269_), .A2(\A[299] ), .ZN(new_n2315_));
  NOR2_X1    g01311(.A1(new_n2267_), .A2(\A[300] ), .ZN(new_n2316_));
  OAI21_X1   g01312(.A1(new_n2315_), .A2(new_n2316_), .B(\A[298] ), .ZN(new_n2317_));
  AND2_X2    g01313(.A1(\A[299] ), .A2(\A[300] ), .Z(new_n2318_));
  OAI21_X1   g01314(.A1(new_n2318_), .A2(new_n2276_), .B(new_n2266_), .ZN(new_n2319_));
  NAND2_X1   g01315(.A1(new_n2317_), .A2(new_n2319_), .ZN(new_n2320_));
  OAI21_X1   g01316(.A1(new_n2314_), .A2(new_n2320_), .B(new_n2278_), .ZN(new_n2321_));
  INV_X1     g01317(.I(new_n2278_), .ZN(new_n2322_));
  NAND3_X1   g01318(.A1(new_n2265_), .A2(new_n2275_), .A3(new_n2322_), .ZN(new_n2323_));
  AOI21_X1   g01319(.A1(new_n2321_), .A2(new_n2323_), .B(new_n2308_), .ZN(new_n2324_));
  AOI21_X1   g01320(.A1(new_n2265_), .A2(new_n2275_), .B(new_n2322_), .ZN(new_n2325_));
  NOR3_X1    g01321(.A1(new_n2314_), .A2(new_n2320_), .A3(new_n2278_), .ZN(new_n2326_));
  NOR3_X1    g01322(.A1(new_n2325_), .A2(new_n2326_), .A3(new_n2277_), .ZN(new_n2327_));
  NOR2_X1    g01323(.A1(new_n2324_), .A2(new_n2327_), .ZN(new_n2328_));
  NOR2_X1    g01324(.A1(new_n2307_), .A2(new_n2328_), .ZN(new_n2329_));
  OAI21_X1   g01325(.A1(new_n2325_), .A2(new_n2326_), .B(new_n2277_), .ZN(new_n2330_));
  NAND3_X1   g01326(.A1(new_n2321_), .A2(new_n2323_), .A3(new_n2308_), .ZN(new_n2331_));
  NAND2_X1   g01327(.A1(new_n2330_), .A2(new_n2331_), .ZN(new_n2332_));
  NOR3_X1    g01328(.A1(new_n2314_), .A2(new_n2320_), .A3(new_n2279_), .ZN(new_n2333_));
  NAND4_X1   g01329(.A1(new_n2254_), .A2(new_n2300_), .A3(new_n2239_), .A4(new_n2333_), .ZN(new_n2334_));
  NAND2_X1   g01330(.A1(new_n2332_), .A2(new_n2334_), .ZN(new_n2335_));
  INV_X1     g01331(.I(new_n2238_), .ZN(new_n2336_));
  NOR2_X1    g01332(.A1(new_n2252_), .A2(new_n2223_), .ZN(new_n2337_));
  NOR2_X1    g01333(.A1(new_n2246_), .A2(new_n2233_), .ZN(new_n2338_));
  OAI21_X1   g01334(.A1(new_n2337_), .A2(new_n2338_), .B(new_n2336_), .ZN(new_n2339_));
  NAND3_X1   g01335(.A1(new_n2292_), .A2(new_n2296_), .A3(new_n2339_), .ZN(new_n2340_));
  OAI21_X1   g01336(.A1(new_n2332_), .A2(new_n2334_), .B(new_n2340_), .ZN(new_n2341_));
  AOI21_X1   g01337(.A1(new_n2294_), .A2(new_n2295_), .B(new_n2293_), .ZN(new_n2342_));
  NOR3_X1    g01338(.A1(new_n2290_), .A2(new_n2291_), .A3(new_n2235_), .ZN(new_n2343_));
  NOR3_X1    g01339(.A1(new_n2342_), .A2(new_n2343_), .A3(new_n2305_), .ZN(new_n2344_));
  NAND2_X1   g01340(.A1(new_n2246_), .A2(new_n2252_), .ZN(new_n2345_));
  NAND2_X1   g01341(.A1(new_n2223_), .A2(new_n2233_), .ZN(new_n2346_));
  NAND3_X1   g01342(.A1(new_n2239_), .A2(new_n2345_), .A3(new_n2346_), .ZN(new_n2347_));
  OAI22_X1   g01343(.A1(new_n2260_), .A2(new_n2264_), .B1(new_n2271_), .B2(new_n2274_), .ZN(new_n2348_));
  NAND3_X1   g01344(.A1(new_n2333_), .A2(new_n2302_), .A3(new_n2348_), .ZN(new_n2349_));
  NOR4_X1    g01345(.A1(new_n2324_), .A2(new_n2327_), .A3(new_n2347_), .A4(new_n2349_), .ZN(new_n2350_));
  NAND2_X1   g01346(.A1(new_n2350_), .A2(new_n2344_), .ZN(new_n2351_));
  NAND2_X1   g01347(.A1(new_n2341_), .A2(new_n2351_), .ZN(new_n2352_));
  AOI21_X1   g01348(.A1(new_n2352_), .A2(new_n2335_), .B(new_n2329_), .ZN(new_n2353_));
  OAI22_X1   g01349(.A1(new_n2284_), .A2(new_n2288_), .B1(new_n2353_), .B2(new_n2196_), .ZN(new_n2354_));
  AOI21_X1   g01350(.A1(new_n2180_), .A2(new_n2173_), .B(new_n2199_), .ZN(new_n2355_));
  NAND2_X1   g01351(.A1(new_n2155_), .A2(new_n2152_), .ZN(new_n2356_));
  AOI21_X1   g01352(.A1(new_n2163_), .A2(new_n2356_), .B(new_n2162_), .ZN(new_n2357_));
  NAND2_X1   g01353(.A1(new_n2105_), .A2(new_n2074_), .ZN(new_n2358_));
  AOI21_X1   g01354(.A1(new_n2089_), .A2(new_n2358_), .B(new_n2171_), .ZN(new_n2359_));
  XOR2_X1    g01355(.A1(new_n2359_), .A2(new_n2357_), .Z(new_n2360_));
  NOR3_X1    g01356(.A1(new_n2355_), .A2(new_n2194_), .A3(new_n2360_), .ZN(new_n2361_));
  OAI21_X1   g01357(.A1(new_n2344_), .A2(new_n2334_), .B(new_n2332_), .ZN(new_n2362_));
  NOR2_X1    g01358(.A1(new_n2235_), .A2(new_n2237_), .ZN(new_n2363_));
  OAI21_X1   g01359(.A1(new_n2345_), .A2(new_n2363_), .B(new_n2238_), .ZN(new_n2364_));
  NAND2_X1   g01360(.A1(new_n2322_), .A2(new_n2308_), .ZN(new_n2365_));
  AOI21_X1   g01361(.A1(new_n2298_), .A2(new_n2365_), .B(new_n2280_), .ZN(new_n2366_));
  XOR2_X1    g01362(.A1(new_n2364_), .A2(new_n2366_), .Z(new_n2367_));
  NAND3_X1   g01363(.A1(new_n2362_), .A2(new_n2307_), .A3(new_n2367_), .ZN(new_n2368_));
  XOR2_X1    g01364(.A1(new_n2361_), .A2(new_n2368_), .Z(new_n2369_));
  NOR2_X1    g01365(.A1(new_n2354_), .A2(new_n2369_), .ZN(new_n2370_));
  NAND2_X1   g01366(.A1(new_n2207_), .A2(new_n2202_), .ZN(new_n2371_));
  OAI21_X1   g01367(.A1(new_n2195_), .A2(new_n2188_), .B(new_n2287_), .ZN(new_n2372_));
  NAND3_X1   g01368(.A1(new_n2207_), .A2(new_n2202_), .A3(new_n2283_), .ZN(new_n2373_));
  NOR2_X1    g01369(.A1(new_n2342_), .A2(new_n2343_), .ZN(new_n2374_));
  NOR3_X1    g01370(.A1(new_n2347_), .A2(new_n2298_), .A3(new_n2299_), .ZN(new_n2375_));
  NAND2_X1   g01371(.A1(new_n2339_), .A2(new_n2333_), .ZN(new_n2376_));
  AOI21_X1   g01372(.A1(new_n2374_), .A2(new_n2375_), .B(new_n2376_), .ZN(new_n2377_));
  NAND2_X1   g01373(.A1(new_n2377_), .A2(new_n2332_), .ZN(new_n2378_));
  NOR2_X1    g01374(.A1(new_n2350_), .A2(new_n2344_), .ZN(new_n2379_));
  NOR3_X1    g01375(.A1(new_n2340_), .A2(new_n2332_), .A3(new_n2334_), .ZN(new_n2380_));
  OAI21_X1   g01376(.A1(new_n2379_), .A2(new_n2380_), .B(new_n2335_), .ZN(new_n2381_));
  NAND2_X1   g01377(.A1(new_n2381_), .A2(new_n2378_), .ZN(new_n2382_));
  AOI22_X1   g01378(.A1(new_n2372_), .A2(new_n2373_), .B1(new_n2382_), .B2(new_n2371_), .ZN(new_n2383_));
  NOR2_X1    g01379(.A1(new_n2347_), .A2(new_n2349_), .ZN(new_n2384_));
  AOI21_X1   g01380(.A1(new_n2340_), .A2(new_n2384_), .B(new_n2328_), .ZN(new_n2385_));
  XNOR2_X1   g01381(.A1(new_n2364_), .A2(new_n2366_), .ZN(new_n2386_));
  NOR3_X1    g01382(.A1(new_n2385_), .A2(new_n2377_), .A3(new_n2386_), .ZN(new_n2387_));
  NOR2_X1    g01383(.A1(new_n2361_), .A2(new_n2387_), .ZN(new_n2388_));
  OAI21_X1   g01384(.A1(new_n2161_), .A2(new_n2186_), .B(new_n2111_), .ZN(new_n2389_));
  XNOR2_X1   g01385(.A1(new_n2359_), .A2(new_n2357_), .ZN(new_n2390_));
  NAND3_X1   g01386(.A1(new_n2389_), .A2(new_n2206_), .A3(new_n2390_), .ZN(new_n2391_));
  NOR2_X1    g01387(.A1(new_n2391_), .A2(new_n2368_), .ZN(new_n2392_));
  NOR2_X1    g01388(.A1(new_n2388_), .A2(new_n2392_), .ZN(new_n2393_));
  NOR2_X1    g01389(.A1(new_n2383_), .A2(new_n2393_), .ZN(new_n2394_));
  NOR4_X1    g01390(.A1(new_n2045_), .A2(new_n2065_), .A3(new_n2370_), .A4(new_n2394_), .ZN(new_n2395_));
  NOR3_X1    g01391(.A1(new_n2288_), .A2(new_n2284_), .A3(new_n2382_), .ZN(new_n2396_));
  INV_X1     g01392(.I(new_n2396_), .ZN(new_n2397_));
  AOI21_X1   g01393(.A1(new_n2286_), .A2(new_n2285_), .B(new_n2281_), .ZN(new_n2398_));
  NOR2_X1    g01394(.A1(new_n2398_), .A2(new_n2283_), .ZN(new_n2399_));
  NAND2_X1   g01395(.A1(new_n1886_), .A2(new_n1955_), .ZN(new_n2400_));
  NAND3_X1   g01396(.A1(new_n2399_), .A2(new_n1961_), .A3(new_n2400_), .ZN(new_n2401_));
  NAND2_X1   g01397(.A1(new_n2397_), .A2(new_n2401_), .ZN(new_n2402_));
  INV_X1     g01398(.I(new_n2401_), .ZN(new_n2403_));
  NAND2_X1   g01399(.A1(new_n2403_), .A2(new_n2396_), .ZN(new_n2404_));
  OAI21_X1   g01400(.A1(new_n1957_), .A2(new_n1962_), .B(new_n2027_), .ZN(new_n2405_));
  NAND3_X1   g01401(.A1(new_n2047_), .A2(new_n2048_), .A3(new_n2057_), .ZN(new_n2406_));
  NAND2_X1   g01402(.A1(new_n2405_), .A2(new_n2406_), .ZN(new_n2407_));
  AOI22_X1   g01403(.A1(new_n2402_), .A2(new_n2404_), .B1(new_n2407_), .B2(new_n2397_), .ZN(new_n2408_));
  OAI22_X1   g01404(.A1(new_n2045_), .A2(new_n2065_), .B1(new_n2370_), .B2(new_n2394_), .ZN(new_n2409_));
  AOI21_X1   g01405(.A1(new_n2408_), .A2(new_n2409_), .B(new_n2395_), .ZN(new_n2410_));
  INV_X1     g01406(.I(new_n2033_), .ZN(new_n2411_));
  NAND2_X1   g01407(.A1(new_n2411_), .A2(new_n2031_), .ZN(new_n2412_));
  NOR2_X1    g01408(.A1(new_n2029_), .A2(new_n1868_), .ZN(new_n2413_));
  OAI21_X1   g01409(.A1(new_n2031_), .A2(new_n2411_), .B(new_n2413_), .ZN(new_n2414_));
  NAND2_X1   g01410(.A1(new_n2414_), .A2(new_n2412_), .ZN(new_n2415_));
  NAND2_X1   g01411(.A1(new_n2062_), .A2(new_n2043_), .ZN(new_n2416_));
  NAND2_X1   g01412(.A1(new_n2059_), .A2(new_n2036_), .ZN(new_n2417_));
  AOI21_X1   g01413(.A1(new_n2028_), .A2(new_n2416_), .B(new_n2417_), .ZN(new_n2418_));
  NAND2_X1   g01414(.A1(new_n2039_), .A2(new_n2041_), .ZN(new_n2419_));
  OR2_X2     g01415(.A1(new_n2039_), .A2(new_n2041_), .Z(new_n2420_));
  NAND3_X1   g01416(.A1(new_n2037_), .A2(new_n1981_), .A3(new_n2420_), .ZN(new_n2421_));
  NAND2_X1   g01417(.A1(new_n2421_), .A2(new_n2419_), .ZN(new_n2422_));
  INV_X1     g01418(.I(new_n2422_), .ZN(new_n2423_));
  NOR2_X1    g01419(.A1(new_n2418_), .A2(new_n2423_), .ZN(new_n2424_));
  NOR4_X1    g01420(.A1(new_n2028_), .A2(new_n2422_), .A3(new_n2062_), .A4(new_n2043_), .ZN(new_n2425_));
  OAI21_X1   g01421(.A1(new_n2424_), .A2(new_n2425_), .B(new_n2415_), .ZN(new_n2426_));
  INV_X1     g01422(.I(new_n2415_), .ZN(new_n2427_));
  NAND3_X1   g01423(.A1(new_n2058_), .A2(new_n2036_), .A3(new_n2059_), .ZN(new_n2428_));
  NAND2_X1   g01424(.A1(new_n2428_), .A2(new_n2422_), .ZN(new_n2429_));
  NAND4_X1   g01425(.A1(new_n2058_), .A2(new_n2423_), .A3(new_n2036_), .A4(new_n2059_), .ZN(new_n2430_));
  NAND3_X1   g01426(.A1(new_n2429_), .A2(new_n2427_), .A3(new_n2430_), .ZN(new_n2431_));
  NAND2_X1   g01427(.A1(new_n2426_), .A2(new_n2431_), .ZN(new_n2432_));
  OR2_X2     g01428(.A1(new_n2359_), .A2(new_n2357_), .Z(new_n2433_));
  NAND2_X1   g01429(.A1(new_n2359_), .A2(new_n2357_), .ZN(new_n2434_));
  NAND3_X1   g01430(.A1(new_n2389_), .A2(new_n2206_), .A3(new_n2434_), .ZN(new_n2435_));
  NAND2_X1   g01431(.A1(new_n2435_), .A2(new_n2433_), .ZN(new_n2436_));
  INV_X1     g01432(.I(new_n2436_), .ZN(new_n2437_));
  NAND3_X1   g01433(.A1(new_n2383_), .A2(new_n2361_), .A3(new_n2387_), .ZN(new_n2438_));
  INV_X1     g01434(.I(new_n2366_), .ZN(new_n2439_));
  NAND2_X1   g01435(.A1(new_n2439_), .A2(new_n2364_), .ZN(new_n2440_));
  NOR2_X1    g01436(.A1(new_n2385_), .A2(new_n2377_), .ZN(new_n2441_));
  OAI21_X1   g01437(.A1(new_n2364_), .A2(new_n2439_), .B(new_n2441_), .ZN(new_n2442_));
  NAND2_X1   g01438(.A1(new_n2442_), .A2(new_n2440_), .ZN(new_n2443_));
  NAND2_X1   g01439(.A1(new_n2438_), .A2(new_n2443_), .ZN(new_n2444_));
  AND2_X2    g01440(.A1(new_n2442_), .A2(new_n2440_), .Z(new_n2445_));
  NAND4_X1   g01441(.A1(new_n2445_), .A2(new_n2383_), .A3(new_n2361_), .A4(new_n2387_), .ZN(new_n2446_));
  AOI21_X1   g01442(.A1(new_n2444_), .A2(new_n2446_), .B(new_n2437_), .ZN(new_n2447_));
  NAND2_X1   g01443(.A1(new_n2196_), .A2(new_n2283_), .ZN(new_n2448_));
  OAI21_X1   g01444(.A1(new_n2284_), .A2(new_n2288_), .B(new_n2353_), .ZN(new_n2449_));
  NAND2_X1   g01445(.A1(new_n2391_), .A2(new_n2368_), .ZN(new_n2450_));
  NAND3_X1   g01446(.A1(new_n2449_), .A2(new_n2448_), .A3(new_n2450_), .ZN(new_n2451_));
  AOI21_X1   g01447(.A1(new_n2451_), .A2(new_n2392_), .B(new_n2445_), .ZN(new_n2452_));
  NOR4_X1    g01448(.A1(new_n2354_), .A2(new_n2391_), .A3(new_n2368_), .A4(new_n2443_), .ZN(new_n2453_));
  NOR3_X1    g01449(.A1(new_n2452_), .A2(new_n2436_), .A3(new_n2453_), .ZN(new_n2454_));
  NOR2_X1    g01450(.A1(new_n2454_), .A2(new_n2447_), .ZN(new_n2455_));
  NAND2_X1   g01451(.A1(new_n2432_), .A2(new_n2455_), .ZN(new_n2456_));
  AOI21_X1   g01452(.A1(new_n2429_), .A2(new_n2430_), .B(new_n2427_), .ZN(new_n2457_));
  NOR3_X1    g01453(.A1(new_n2424_), .A2(new_n2415_), .A3(new_n2425_), .ZN(new_n2458_));
  NOR2_X1    g01454(.A1(new_n2458_), .A2(new_n2457_), .ZN(new_n2459_));
  OAI21_X1   g01455(.A1(new_n2452_), .A2(new_n2453_), .B(new_n2436_), .ZN(new_n2460_));
  NAND3_X1   g01456(.A1(new_n2444_), .A2(new_n2437_), .A3(new_n2446_), .ZN(new_n2461_));
  NAND2_X1   g01457(.A1(new_n2460_), .A2(new_n2461_), .ZN(new_n2462_));
  NAND2_X1   g01458(.A1(new_n2459_), .A2(new_n2462_), .ZN(new_n2463_));
  AOI21_X1   g01459(.A1(new_n2456_), .A2(new_n2463_), .B(new_n2410_), .ZN(new_n2464_));
  XNOR2_X1   g01460(.A1(new_n2036_), .A2(new_n2043_), .ZN(new_n2465_));
  NAND2_X1   g01461(.A1(new_n2465_), .A2(new_n2058_), .ZN(new_n2466_));
  NAND2_X1   g01462(.A1(new_n2417_), .A2(new_n2416_), .ZN(new_n2467_));
  NAND2_X1   g01463(.A1(new_n2028_), .A2(new_n2467_), .ZN(new_n2468_));
  XOR2_X1    g01464(.A1(new_n2391_), .A2(new_n2368_), .Z(new_n2469_));
  NAND2_X1   g01465(.A1(new_n2383_), .A2(new_n2469_), .ZN(new_n2470_));
  INV_X1     g01466(.I(new_n2392_), .ZN(new_n2471_));
  NAND2_X1   g01467(.A1(new_n2471_), .A2(new_n2450_), .ZN(new_n2472_));
  NAND2_X1   g01468(.A1(new_n2472_), .A2(new_n2354_), .ZN(new_n2473_));
  NAND4_X1   g01469(.A1(new_n2466_), .A2(new_n2468_), .A3(new_n2473_), .A4(new_n2470_), .ZN(new_n2474_));
  NOR2_X1    g01470(.A1(new_n2403_), .A2(new_n2396_), .ZN(new_n2475_));
  INV_X1     g01471(.I(new_n2404_), .ZN(new_n2476_));
  AOI21_X1   g01472(.A1(new_n2047_), .A2(new_n2048_), .B(new_n2057_), .ZN(new_n2477_));
  NOR3_X1    g01473(.A1(new_n1962_), .A2(new_n2027_), .A3(new_n1957_), .ZN(new_n2478_));
  NOR2_X1    g01474(.A1(new_n2478_), .A2(new_n2477_), .ZN(new_n2479_));
  OAI22_X1   g01475(.A1(new_n2476_), .A2(new_n2475_), .B1(new_n2396_), .B2(new_n2479_), .ZN(new_n2480_));
  AOI22_X1   g01476(.A1(new_n2466_), .A2(new_n2468_), .B1(new_n2473_), .B2(new_n2470_), .ZN(new_n2481_));
  OAI21_X1   g01477(.A1(new_n2480_), .A2(new_n2481_), .B(new_n2474_), .ZN(new_n2482_));
  NAND4_X1   g01478(.A1(new_n2426_), .A2(new_n2460_), .A3(new_n2431_), .A4(new_n2461_), .ZN(new_n2483_));
  OAI22_X1   g01479(.A1(new_n2458_), .A2(new_n2457_), .B1(new_n2454_), .B2(new_n2447_), .ZN(new_n2484_));
  AOI21_X1   g01480(.A1(new_n2484_), .A2(new_n2483_), .B(new_n2482_), .ZN(new_n2485_));
  NOR4_X1    g01481(.A1(new_n2464_), .A2(new_n1724_), .A3(new_n1742_), .A4(new_n2485_), .ZN(new_n2486_));
  NOR2_X1    g01482(.A1(new_n2370_), .A2(new_n2394_), .ZN(new_n2487_));
  NOR3_X1    g01483(.A1(new_n2487_), .A2(new_n2045_), .A3(new_n2065_), .ZN(new_n2488_));
  NOR2_X1    g01484(.A1(new_n2045_), .A2(new_n2065_), .ZN(new_n2489_));
  NOR3_X1    g01485(.A1(new_n2489_), .A2(new_n2370_), .A3(new_n2394_), .ZN(new_n2490_));
  OAI21_X1   g01486(.A1(new_n2490_), .A2(new_n2488_), .B(new_n2408_), .ZN(new_n2491_));
  OAI21_X1   g01487(.A1(new_n2395_), .A2(new_n2481_), .B(new_n2480_), .ZN(new_n2492_));
  AOI21_X1   g01488(.A1(new_n1732_), .A2(new_n1735_), .B(new_n1316_), .ZN(new_n2493_));
  NOR3_X1    g01489(.A1(new_n1729_), .A2(new_n1633_), .A3(new_n1647_), .ZN(new_n2494_));
  OAI21_X1   g01490(.A1(new_n2493_), .A2(new_n2494_), .B(new_n1670_), .ZN(new_n2495_));
  OAI21_X1   g01491(.A1(new_n1738_), .A2(new_n1648_), .B(new_n1737_), .ZN(new_n2496_));
  NAND4_X1   g01492(.A1(new_n2496_), .A2(new_n2495_), .A3(new_n2491_), .A4(new_n2492_), .ZN(new_n2497_));
  NAND2_X1   g01493(.A1(new_n1665_), .A2(new_n1666_), .ZN(new_n2498_));
  NOR2_X1    g01494(.A1(new_n2498_), .A2(new_n1669_), .ZN(new_n2499_));
  NOR2_X1    g01495(.A1(new_n1654_), .A2(new_n1657_), .ZN(new_n2500_));
  NOR2_X1    g01496(.A1(new_n1660_), .A2(new_n1662_), .ZN(new_n2501_));
  NOR2_X1    g01497(.A1(new_n2500_), .A2(new_n2501_), .ZN(new_n2502_));
  NOR2_X1    g01498(.A1(new_n2502_), .A2(new_n1663_), .ZN(new_n2503_));
  INV_X1     g01499(.I(new_n2503_), .ZN(new_n2504_));
  NAND2_X1   g01500(.A1(new_n1961_), .A2(new_n2400_), .ZN(new_n2505_));
  OAI21_X1   g01501(.A1(new_n2283_), .A2(new_n2398_), .B(new_n2505_), .ZN(new_n2506_));
  NAND2_X1   g01502(.A1(new_n2506_), .A2(new_n2401_), .ZN(new_n2507_));
  OAI22_X1   g01503(.A1(new_n2498_), .A2(new_n1669_), .B1(new_n2504_), .B2(new_n2507_), .ZN(new_n2508_));
  INV_X1     g01504(.I(new_n1669_), .ZN(new_n2509_));
  NOR3_X1    g01505(.A1(new_n2507_), .A2(new_n1663_), .A3(new_n2502_), .ZN(new_n2510_));
  NAND4_X1   g01506(.A1(new_n2510_), .A2(new_n1665_), .A3(new_n1666_), .A4(new_n2509_), .ZN(new_n2511_));
  NAND2_X1   g01507(.A1(new_n2508_), .A2(new_n2511_), .ZN(new_n2512_));
  NOR2_X1    g01508(.A1(new_n2476_), .A2(new_n2475_), .ZN(new_n2513_));
  XOR2_X1    g01509(.A1(new_n2513_), .A2(new_n2407_), .Z(new_n2514_));
  OAI21_X1   g01510(.A1(new_n2514_), .A2(new_n2499_), .B(new_n2512_), .ZN(new_n2515_));
  AOI22_X1   g01511(.A1(new_n2496_), .A2(new_n2495_), .B1(new_n2491_), .B2(new_n2492_), .ZN(new_n2516_));
  OAI21_X1   g01512(.A1(new_n2516_), .A2(new_n2515_), .B(new_n2497_), .ZN(new_n2517_));
  OAI22_X1   g01513(.A1(new_n2464_), .A2(new_n2485_), .B1(new_n1724_), .B2(new_n1742_), .ZN(new_n2518_));
  AOI21_X1   g01514(.A1(new_n2518_), .A2(new_n2517_), .B(new_n2486_), .ZN(new_n2519_));
  NOR3_X1    g01515(.A1(new_n1722_), .A2(new_n1691_), .A3(new_n1695_), .ZN(new_n2520_));
  NAND2_X1   g01516(.A1(new_n1689_), .A2(new_n1682_), .ZN(new_n2521_));
  XOR2_X1    g01517(.A1(new_n1699_), .A2(new_n1706_), .Z(new_n2522_));
  XOR2_X1    g01518(.A1(new_n1676_), .A2(new_n1686_), .Z(new_n2523_));
  NOR4_X1    g01519(.A1(new_n2522_), .A2(new_n2523_), .A3(new_n2521_), .A4(new_n1702_), .ZN(new_n2524_));
  OAI21_X1   g01520(.A1(new_n2520_), .A2(new_n1739_), .B(new_n2524_), .ZN(new_n2525_));
  NOR2_X1    g01521(.A1(new_n1692_), .A2(new_n1687_), .ZN(new_n2526_));
  INV_X1     g01522(.I(new_n2526_), .ZN(new_n2527_));
  NOR2_X1    g01523(.A1(new_n1676_), .A2(new_n1686_), .ZN(new_n2528_));
  OR3_X2     g01524(.A1(new_n1678_), .A2(new_n1683_), .A3(new_n2528_), .Z(new_n2529_));
  NAND2_X1   g01525(.A1(new_n1699_), .A2(new_n1706_), .ZN(new_n2530_));
  NAND4_X1   g01526(.A1(new_n1698_), .A2(new_n1696_), .A3(new_n1703_), .A4(new_n1705_), .ZN(new_n2531_));
  NAND3_X1   g01527(.A1(new_n1709_), .A2(new_n1708_), .A3(new_n2531_), .ZN(new_n2532_));
  NAND2_X1   g01528(.A1(new_n2532_), .A2(new_n2530_), .ZN(new_n2533_));
  INV_X1     g01529(.I(new_n2533_), .ZN(new_n2534_));
  NAND3_X1   g01530(.A1(new_n2534_), .A2(new_n2529_), .A3(new_n2527_), .ZN(new_n2535_));
  NOR2_X1    g01531(.A1(new_n2521_), .A2(new_n2528_), .ZN(new_n2536_));
  OAI21_X1   g01532(.A1(new_n2536_), .A2(new_n2526_), .B(new_n2533_), .ZN(new_n2537_));
  NAND2_X1   g01533(.A1(new_n2535_), .A2(new_n2537_), .ZN(new_n2538_));
  INV_X1     g01534(.I(new_n2538_), .ZN(new_n2539_));
  NAND2_X1   g01535(.A1(new_n2525_), .A2(new_n2539_), .ZN(new_n2540_));
  NAND2_X1   g01536(.A1(new_n1740_), .A2(new_n1672_), .ZN(new_n2541_));
  NAND3_X1   g01537(.A1(new_n2541_), .A2(new_n2524_), .A3(new_n2538_), .ZN(new_n2542_));
  NAND2_X1   g01538(.A1(new_n2540_), .A2(new_n2542_), .ZN(new_n2543_));
  NAND2_X1   g01539(.A1(new_n2445_), .A2(new_n2437_), .ZN(new_n2544_));
  NAND2_X1   g01540(.A1(new_n2443_), .A2(new_n2436_), .ZN(new_n2545_));
  NAND3_X1   g01541(.A1(new_n2451_), .A2(new_n2392_), .A3(new_n2545_), .ZN(new_n2546_));
  NAND2_X1   g01542(.A1(new_n2546_), .A2(new_n2544_), .ZN(new_n2547_));
  INV_X1     g01543(.I(new_n2547_), .ZN(new_n2548_));
  NAND2_X1   g01544(.A1(new_n2427_), .A2(new_n2423_), .ZN(new_n2549_));
  NAND2_X1   g01545(.A1(new_n2415_), .A2(new_n2422_), .ZN(new_n2550_));
  NAND2_X1   g01546(.A1(new_n2418_), .A2(new_n2550_), .ZN(new_n2551_));
  AND2_X2    g01547(.A1(new_n2551_), .A2(new_n2549_), .Z(new_n2552_));
  INV_X1     g01548(.I(new_n2552_), .ZN(new_n2553_));
  OAI21_X1   g01549(.A1(new_n2432_), .A2(new_n2462_), .B(new_n2410_), .ZN(new_n2554_));
  XOR2_X1    g01550(.A1(new_n2415_), .A2(new_n2422_), .Z(new_n2555_));
  XOR2_X1    g01551(.A1(new_n2443_), .A2(new_n2436_), .Z(new_n2556_));
  NOR4_X1    g01552(.A1(new_n2555_), .A2(new_n2556_), .A3(new_n2428_), .A4(new_n2438_), .ZN(new_n2557_));
  AOI21_X1   g01553(.A1(new_n2554_), .A2(new_n2557_), .B(new_n2553_), .ZN(new_n2558_));
  AOI21_X1   g01554(.A1(new_n2459_), .A2(new_n2455_), .B(new_n2482_), .ZN(new_n2559_));
  INV_X1     g01555(.I(new_n2557_), .ZN(new_n2560_));
  NOR3_X1    g01556(.A1(new_n2559_), .A2(new_n2552_), .A3(new_n2560_), .ZN(new_n2561_));
  OAI21_X1   g01557(.A1(new_n2561_), .A2(new_n2558_), .B(new_n2548_), .ZN(new_n2562_));
  OAI21_X1   g01558(.A1(new_n2559_), .A2(new_n2560_), .B(new_n2552_), .ZN(new_n2563_));
  NAND3_X1   g01559(.A1(new_n2554_), .A2(new_n2553_), .A3(new_n2557_), .ZN(new_n2564_));
  NAND3_X1   g01560(.A1(new_n2563_), .A2(new_n2564_), .A3(new_n2547_), .ZN(new_n2565_));
  NAND3_X1   g01561(.A1(new_n2543_), .A2(new_n2562_), .A3(new_n2565_), .ZN(new_n2566_));
  AOI21_X1   g01562(.A1(new_n2541_), .A2(new_n2524_), .B(new_n2538_), .ZN(new_n2567_));
  NOR2_X1    g01563(.A1(new_n2525_), .A2(new_n2539_), .ZN(new_n2568_));
  NOR2_X1    g01564(.A1(new_n2568_), .A2(new_n2567_), .ZN(new_n2569_));
  AOI21_X1   g01565(.A1(new_n2563_), .A2(new_n2564_), .B(new_n2547_), .ZN(new_n2570_));
  NOR3_X1    g01566(.A1(new_n2561_), .A2(new_n2558_), .A3(new_n2548_), .ZN(new_n2571_));
  OAI21_X1   g01567(.A1(new_n2570_), .A2(new_n2571_), .B(new_n2569_), .ZN(new_n2572_));
  AOI21_X1   g01568(.A1(new_n2572_), .A2(new_n2566_), .B(new_n2519_), .ZN(new_n2573_));
  AOI21_X1   g01569(.A1(new_n1718_), .A2(new_n1719_), .B(new_n1722_), .ZN(new_n2574_));
  NOR3_X1    g01570(.A1(new_n1716_), .A2(new_n1691_), .A3(new_n1695_), .ZN(new_n2575_));
  OAI21_X1   g01571(.A1(new_n2574_), .A2(new_n2575_), .B(new_n1739_), .ZN(new_n2576_));
  AOI22_X1   g01572(.A1(new_n1718_), .A2(new_n1719_), .B1(new_n1720_), .B2(new_n1721_), .ZN(new_n2577_));
  OAI21_X1   g01573(.A1(new_n2520_), .A2(new_n2577_), .B(new_n1672_), .ZN(new_n2578_));
  NOR2_X1    g01574(.A1(new_n2459_), .A2(new_n2462_), .ZN(new_n2579_));
  NOR2_X1    g01575(.A1(new_n2432_), .A2(new_n2455_), .ZN(new_n2580_));
  OAI21_X1   g01576(.A1(new_n2580_), .A2(new_n2579_), .B(new_n2482_), .ZN(new_n2581_));
  NOR4_X1    g01577(.A1(new_n2458_), .A2(new_n2454_), .A3(new_n2457_), .A4(new_n2447_), .ZN(new_n2582_));
  AOI22_X1   g01578(.A1(new_n2426_), .A2(new_n2431_), .B1(new_n2460_), .B2(new_n2461_), .ZN(new_n2583_));
  OAI21_X1   g01579(.A1(new_n2583_), .A2(new_n2582_), .B(new_n2410_), .ZN(new_n2584_));
  NAND4_X1   g01580(.A1(new_n2581_), .A2(new_n2576_), .A3(new_n2578_), .A4(new_n2584_), .ZN(new_n2585_));
  NAND2_X1   g01581(.A1(new_n2491_), .A2(new_n2492_), .ZN(new_n2586_));
  NAND2_X1   g01582(.A1(new_n2496_), .A2(new_n2495_), .ZN(new_n2587_));
  NOR2_X1    g01583(.A1(new_n2587_), .A2(new_n2586_), .ZN(new_n2588_));
  INV_X1     g01584(.I(new_n2515_), .ZN(new_n2589_));
  NAND2_X1   g01585(.A1(new_n2587_), .A2(new_n2586_), .ZN(new_n2590_));
  AOI21_X1   g01586(.A1(new_n2589_), .A2(new_n2590_), .B(new_n2588_), .ZN(new_n2591_));
  AOI22_X1   g01587(.A1(new_n2581_), .A2(new_n2584_), .B1(new_n2576_), .B2(new_n2578_), .ZN(new_n2592_));
  OAI21_X1   g01588(.A1(new_n2591_), .A2(new_n2592_), .B(new_n2585_), .ZN(new_n2593_));
  NAND3_X1   g01589(.A1(new_n2569_), .A2(new_n2562_), .A3(new_n2565_), .ZN(new_n2594_));
  OAI21_X1   g01590(.A1(new_n2570_), .A2(new_n2571_), .B(new_n2543_), .ZN(new_n2595_));
  AOI21_X1   g01591(.A1(new_n2595_), .A2(new_n2594_), .B(new_n2593_), .ZN(new_n2596_));
  INV_X1     g01592(.I(\A[430] ), .ZN(new_n2597_));
  NOR2_X1    g01593(.A1(\A[431] ), .A2(\A[432] ), .ZN(new_n2598_));
  NAND2_X1   g01594(.A1(\A[431] ), .A2(\A[432] ), .ZN(new_n2599_));
  AOI21_X1   g01595(.A1(new_n2597_), .A2(new_n2599_), .B(new_n2598_), .ZN(new_n2600_));
  INV_X1     g01596(.I(new_n2600_), .ZN(new_n2601_));
  INV_X1     g01597(.I(\A[427] ), .ZN(new_n2602_));
  NOR2_X1    g01598(.A1(\A[428] ), .A2(\A[429] ), .ZN(new_n2603_));
  NAND2_X1   g01599(.A1(\A[428] ), .A2(\A[429] ), .ZN(new_n2604_));
  AOI21_X1   g01600(.A1(new_n2602_), .A2(new_n2604_), .B(new_n2603_), .ZN(new_n2605_));
  INV_X1     g01601(.I(\A[429] ), .ZN(new_n2606_));
  NOR2_X1    g01602(.A1(new_n2606_), .A2(\A[428] ), .ZN(new_n2607_));
  INV_X1     g01603(.I(\A[428] ), .ZN(new_n2608_));
  NOR2_X1    g01604(.A1(new_n2608_), .A2(\A[429] ), .ZN(new_n2609_));
  OAI21_X1   g01605(.A1(new_n2607_), .A2(new_n2609_), .B(\A[427] ), .ZN(new_n2610_));
  INV_X1     g01606(.I(new_n2604_), .ZN(new_n2611_));
  OAI21_X1   g01607(.A1(new_n2611_), .A2(new_n2603_), .B(new_n2602_), .ZN(new_n2612_));
  NAND2_X1   g01608(.A1(new_n2610_), .A2(new_n2612_), .ZN(new_n2613_));
  INV_X1     g01609(.I(\A[432] ), .ZN(new_n2614_));
  NOR2_X1    g01610(.A1(new_n2614_), .A2(\A[431] ), .ZN(new_n2615_));
  INV_X1     g01611(.I(\A[431] ), .ZN(new_n2616_));
  NOR2_X1    g01612(.A1(new_n2616_), .A2(\A[432] ), .ZN(new_n2617_));
  OAI21_X1   g01613(.A1(new_n2615_), .A2(new_n2617_), .B(\A[430] ), .ZN(new_n2618_));
  INV_X1     g01614(.I(new_n2599_), .ZN(new_n2619_));
  OAI21_X1   g01615(.A1(new_n2619_), .A2(new_n2598_), .B(new_n2597_), .ZN(new_n2620_));
  NAND2_X1   g01616(.A1(new_n2618_), .A2(new_n2620_), .ZN(new_n2621_));
  OAI21_X1   g01617(.A1(new_n2613_), .A2(new_n2621_), .B(new_n2605_), .ZN(new_n2622_));
  INV_X1     g01618(.I(new_n2605_), .ZN(new_n2623_));
  NAND2_X1   g01619(.A1(new_n2608_), .A2(\A[429] ), .ZN(new_n2624_));
  NAND2_X1   g01620(.A1(new_n2606_), .A2(\A[428] ), .ZN(new_n2625_));
  AOI21_X1   g01621(.A1(new_n2624_), .A2(new_n2625_), .B(new_n2602_), .ZN(new_n2626_));
  INV_X1     g01622(.I(new_n2603_), .ZN(new_n2627_));
  AOI21_X1   g01623(.A1(new_n2627_), .A2(new_n2604_), .B(\A[427] ), .ZN(new_n2628_));
  NOR2_X1    g01624(.A1(new_n2628_), .A2(new_n2626_), .ZN(new_n2629_));
  NAND2_X1   g01625(.A1(new_n2616_), .A2(\A[432] ), .ZN(new_n2630_));
  NAND2_X1   g01626(.A1(new_n2614_), .A2(\A[431] ), .ZN(new_n2631_));
  AOI21_X1   g01627(.A1(new_n2630_), .A2(new_n2631_), .B(new_n2597_), .ZN(new_n2632_));
  INV_X1     g01628(.I(new_n2598_), .ZN(new_n2633_));
  AOI21_X1   g01629(.A1(new_n2633_), .A2(new_n2599_), .B(\A[430] ), .ZN(new_n2634_));
  NOR2_X1    g01630(.A1(new_n2634_), .A2(new_n2632_), .ZN(new_n2635_));
  NAND3_X1   g01631(.A1(new_n2629_), .A2(new_n2635_), .A3(new_n2623_), .ZN(new_n2636_));
  AOI21_X1   g01632(.A1(new_n2622_), .A2(new_n2636_), .B(new_n2601_), .ZN(new_n2637_));
  AOI21_X1   g01633(.A1(new_n2629_), .A2(new_n2635_), .B(new_n2623_), .ZN(new_n2638_));
  NOR3_X1    g01634(.A1(new_n2613_), .A2(new_n2621_), .A3(new_n2605_), .ZN(new_n2639_));
  NOR3_X1    g01635(.A1(new_n2638_), .A2(new_n2639_), .A3(new_n2600_), .ZN(new_n2640_));
  NOR2_X1    g01636(.A1(new_n2640_), .A2(new_n2637_), .ZN(new_n2641_));
  INV_X1     g01637(.I(\A[436] ), .ZN(new_n2642_));
  NOR2_X1    g01638(.A1(\A[437] ), .A2(\A[438] ), .ZN(new_n2643_));
  NAND2_X1   g01639(.A1(\A[437] ), .A2(\A[438] ), .ZN(new_n2644_));
  AOI21_X1   g01640(.A1(new_n2642_), .A2(new_n2644_), .B(new_n2643_), .ZN(new_n2645_));
  INV_X1     g01641(.I(\A[433] ), .ZN(new_n2646_));
  NOR2_X1    g01642(.A1(\A[434] ), .A2(\A[435] ), .ZN(new_n2647_));
  NAND2_X1   g01643(.A1(\A[434] ), .A2(\A[435] ), .ZN(new_n2648_));
  AOI21_X1   g01644(.A1(new_n2646_), .A2(new_n2648_), .B(new_n2647_), .ZN(new_n2649_));
  INV_X1     g01645(.I(new_n2649_), .ZN(new_n2650_));
  INV_X1     g01646(.I(\A[437] ), .ZN(new_n2651_));
  NAND2_X1   g01647(.A1(new_n2651_), .A2(\A[438] ), .ZN(new_n2652_));
  INV_X1     g01648(.I(\A[438] ), .ZN(new_n2653_));
  NAND2_X1   g01649(.A1(new_n2653_), .A2(\A[437] ), .ZN(new_n2654_));
  AOI21_X1   g01650(.A1(new_n2652_), .A2(new_n2654_), .B(new_n2642_), .ZN(new_n2655_));
  INV_X1     g01651(.I(new_n2643_), .ZN(new_n2656_));
  AOI21_X1   g01652(.A1(new_n2656_), .A2(new_n2644_), .B(\A[436] ), .ZN(new_n2657_));
  NOR2_X1    g01653(.A1(new_n2657_), .A2(new_n2655_), .ZN(new_n2658_));
  INV_X1     g01654(.I(\A[434] ), .ZN(new_n2659_));
  NAND2_X1   g01655(.A1(new_n2659_), .A2(\A[435] ), .ZN(new_n2660_));
  INV_X1     g01656(.I(\A[435] ), .ZN(new_n2661_));
  NAND2_X1   g01657(.A1(new_n2661_), .A2(\A[434] ), .ZN(new_n2662_));
  AOI21_X1   g01658(.A1(new_n2660_), .A2(new_n2662_), .B(new_n2646_), .ZN(new_n2663_));
  INV_X1     g01659(.I(new_n2647_), .ZN(new_n2664_));
  AOI21_X1   g01660(.A1(new_n2664_), .A2(new_n2648_), .B(\A[433] ), .ZN(new_n2665_));
  NOR2_X1    g01661(.A1(new_n2665_), .A2(new_n2663_), .ZN(new_n2666_));
  AOI21_X1   g01662(.A1(new_n2658_), .A2(new_n2666_), .B(new_n2650_), .ZN(new_n2667_));
  NOR2_X1    g01663(.A1(new_n2653_), .A2(\A[437] ), .ZN(new_n2668_));
  NOR2_X1    g01664(.A1(new_n2651_), .A2(\A[438] ), .ZN(new_n2669_));
  OAI21_X1   g01665(.A1(new_n2668_), .A2(new_n2669_), .B(\A[436] ), .ZN(new_n2670_));
  INV_X1     g01666(.I(new_n2644_), .ZN(new_n2671_));
  OAI21_X1   g01667(.A1(new_n2671_), .A2(new_n2643_), .B(new_n2642_), .ZN(new_n2672_));
  NOR2_X1    g01668(.A1(new_n2661_), .A2(\A[434] ), .ZN(new_n2673_));
  NOR2_X1    g01669(.A1(new_n2659_), .A2(\A[435] ), .ZN(new_n2674_));
  OAI21_X1   g01670(.A1(new_n2673_), .A2(new_n2674_), .B(\A[433] ), .ZN(new_n2675_));
  INV_X1     g01671(.I(new_n2648_), .ZN(new_n2676_));
  OAI21_X1   g01672(.A1(new_n2676_), .A2(new_n2647_), .B(new_n2646_), .ZN(new_n2677_));
  NAND4_X1   g01673(.A1(new_n2670_), .A2(new_n2672_), .A3(new_n2675_), .A4(new_n2677_), .ZN(new_n2678_));
  NOR2_X1    g01674(.A1(new_n2678_), .A2(new_n2649_), .ZN(new_n2679_));
  OAI21_X1   g01675(.A1(new_n2679_), .A2(new_n2667_), .B(new_n2645_), .ZN(new_n2680_));
  INV_X1     g01676(.I(new_n2645_), .ZN(new_n2681_));
  NAND2_X1   g01677(.A1(new_n2678_), .A2(new_n2649_), .ZN(new_n2682_));
  NAND3_X1   g01678(.A1(new_n2658_), .A2(new_n2666_), .A3(new_n2650_), .ZN(new_n2683_));
  NAND3_X1   g01679(.A1(new_n2682_), .A2(new_n2683_), .A3(new_n2681_), .ZN(new_n2684_));
  NAND2_X1   g01680(.A1(new_n2680_), .A2(new_n2684_), .ZN(new_n2685_));
  NAND2_X1   g01681(.A1(new_n2629_), .A2(new_n2635_), .ZN(new_n2686_));
  INV_X1     g01682(.I(new_n2678_), .ZN(new_n2687_));
  NAND4_X1   g01683(.A1(new_n2629_), .A2(new_n2635_), .A3(new_n2600_), .A4(new_n2605_), .ZN(new_n2688_));
  NOR2_X1    g01684(.A1(new_n2658_), .A2(new_n2666_), .ZN(new_n2689_));
  NOR3_X1    g01685(.A1(new_n2688_), .A2(new_n2687_), .A3(new_n2689_), .ZN(new_n2690_));
  NAND2_X1   g01686(.A1(new_n2613_), .A2(new_n2621_), .ZN(new_n2691_));
  NAND2_X1   g01687(.A1(new_n2670_), .A2(new_n2672_), .ZN(new_n2692_));
  NAND2_X1   g01688(.A1(new_n2675_), .A2(new_n2677_), .ZN(new_n2693_));
  NAND2_X1   g01689(.A1(new_n2645_), .A2(new_n2649_), .ZN(new_n2694_));
  NOR3_X1    g01690(.A1(new_n2692_), .A2(new_n2693_), .A3(new_n2694_), .ZN(new_n2695_));
  NAND4_X1   g01691(.A1(new_n2690_), .A2(new_n2686_), .A3(new_n2691_), .A4(new_n2695_), .ZN(new_n2696_));
  NAND2_X1   g01692(.A1(new_n2600_), .A2(new_n2605_), .ZN(new_n2697_));
  NOR3_X1    g01693(.A1(new_n2613_), .A2(new_n2621_), .A3(new_n2697_), .ZN(new_n2698_));
  NAND2_X1   g01694(.A1(new_n2692_), .A2(new_n2693_), .ZN(new_n2699_));
  NAND3_X1   g01695(.A1(new_n2698_), .A2(new_n2699_), .A3(new_n2678_), .ZN(new_n2700_));
  NAND2_X1   g01696(.A1(new_n2686_), .A2(new_n2691_), .ZN(new_n2701_));
  NOR2_X1    g01697(.A1(new_n2689_), .A2(new_n2694_), .ZN(new_n2702_));
  NOR3_X1    g01698(.A1(new_n2700_), .A2(new_n2701_), .A3(new_n2702_), .ZN(new_n2703_));
  OAI21_X1   g01699(.A1(new_n2696_), .A2(new_n2685_), .B(new_n2641_), .ZN(new_n2704_));
  NAND3_X1   g01700(.A1(new_n2695_), .A2(new_n2699_), .A3(new_n2678_), .ZN(new_n2705_));
  NOR2_X1    g01701(.A1(new_n2613_), .A2(new_n2621_), .ZN(new_n2706_));
  NOR2_X1    g01702(.A1(new_n2629_), .A2(new_n2635_), .ZN(new_n2707_));
  NOR3_X1    g01703(.A1(new_n2688_), .A2(new_n2707_), .A3(new_n2706_), .ZN(new_n2708_));
  NAND2_X1   g01704(.A1(new_n2708_), .A2(new_n2705_), .ZN(new_n2709_));
  NAND4_X1   g01705(.A1(new_n2658_), .A2(new_n2666_), .A3(new_n2645_), .A4(new_n2649_), .ZN(new_n2710_));
  NOR3_X1    g01706(.A1(new_n2710_), .A2(new_n2687_), .A3(new_n2689_), .ZN(new_n2711_));
  NAND3_X1   g01707(.A1(new_n2698_), .A2(new_n2686_), .A3(new_n2691_), .ZN(new_n2712_));
  NAND2_X1   g01708(.A1(new_n2711_), .A2(new_n2712_), .ZN(new_n2713_));
  INV_X1     g01709(.I(\A[421] ), .ZN(new_n2714_));
  INV_X1     g01710(.I(\A[422] ), .ZN(new_n2715_));
  NAND2_X1   g01711(.A1(new_n2715_), .A2(\A[423] ), .ZN(new_n2716_));
  INV_X1     g01712(.I(\A[423] ), .ZN(new_n2717_));
  NAND2_X1   g01713(.A1(new_n2717_), .A2(\A[422] ), .ZN(new_n2718_));
  AOI21_X1   g01714(.A1(new_n2716_), .A2(new_n2718_), .B(new_n2714_), .ZN(new_n2719_));
  NAND2_X1   g01715(.A1(\A[422] ), .A2(\A[423] ), .ZN(new_n2720_));
  NOR2_X1    g01716(.A1(\A[422] ), .A2(\A[423] ), .ZN(new_n2721_));
  INV_X1     g01717(.I(new_n2721_), .ZN(new_n2722_));
  AOI21_X1   g01718(.A1(new_n2722_), .A2(new_n2720_), .B(\A[421] ), .ZN(new_n2723_));
  NOR2_X1    g01719(.A1(new_n2723_), .A2(new_n2719_), .ZN(new_n2724_));
  INV_X1     g01720(.I(\A[424] ), .ZN(new_n2725_));
  INV_X1     g01721(.I(\A[425] ), .ZN(new_n2726_));
  NAND2_X1   g01722(.A1(new_n2726_), .A2(\A[426] ), .ZN(new_n2727_));
  INV_X1     g01723(.I(\A[426] ), .ZN(new_n2728_));
  NAND2_X1   g01724(.A1(new_n2728_), .A2(\A[425] ), .ZN(new_n2729_));
  AOI21_X1   g01725(.A1(new_n2727_), .A2(new_n2729_), .B(new_n2725_), .ZN(new_n2730_));
  NAND2_X1   g01726(.A1(\A[425] ), .A2(\A[426] ), .ZN(new_n2731_));
  NOR2_X1    g01727(.A1(\A[425] ), .A2(\A[426] ), .ZN(new_n2732_));
  INV_X1     g01728(.I(new_n2732_), .ZN(new_n2733_));
  AOI21_X1   g01729(.A1(new_n2733_), .A2(new_n2731_), .B(\A[424] ), .ZN(new_n2734_));
  NOR2_X1    g01730(.A1(new_n2734_), .A2(new_n2730_), .ZN(new_n2735_));
  NOR2_X1    g01731(.A1(new_n2724_), .A2(new_n2735_), .ZN(new_n2736_));
  NOR4_X1    g01732(.A1(new_n2719_), .A2(new_n2723_), .A3(new_n2734_), .A4(new_n2730_), .ZN(new_n2737_));
  NOR2_X1    g01733(.A1(new_n2736_), .A2(new_n2737_), .ZN(new_n2738_));
  NOR2_X1    g01734(.A1(new_n2717_), .A2(\A[422] ), .ZN(new_n2739_));
  NOR2_X1    g01735(.A1(new_n2715_), .A2(\A[423] ), .ZN(new_n2740_));
  OAI21_X1   g01736(.A1(new_n2739_), .A2(new_n2740_), .B(\A[421] ), .ZN(new_n2741_));
  INV_X1     g01737(.I(new_n2720_), .ZN(new_n2742_));
  OAI21_X1   g01738(.A1(new_n2742_), .A2(new_n2721_), .B(new_n2714_), .ZN(new_n2743_));
  NAND2_X1   g01739(.A1(new_n2741_), .A2(new_n2743_), .ZN(new_n2744_));
  NOR2_X1    g01740(.A1(new_n2728_), .A2(\A[425] ), .ZN(new_n2745_));
  NOR2_X1    g01741(.A1(new_n2726_), .A2(\A[426] ), .ZN(new_n2746_));
  OAI21_X1   g01742(.A1(new_n2745_), .A2(new_n2746_), .B(\A[424] ), .ZN(new_n2747_));
  INV_X1     g01743(.I(new_n2731_), .ZN(new_n2748_));
  OAI21_X1   g01744(.A1(new_n2748_), .A2(new_n2732_), .B(new_n2725_), .ZN(new_n2749_));
  NAND2_X1   g01745(.A1(new_n2747_), .A2(new_n2749_), .ZN(new_n2750_));
  AOI21_X1   g01746(.A1(new_n2725_), .A2(new_n2731_), .B(new_n2732_), .ZN(new_n2751_));
  AOI21_X1   g01747(.A1(new_n2714_), .A2(new_n2720_), .B(new_n2721_), .ZN(new_n2752_));
  NAND2_X1   g01748(.A1(new_n2751_), .A2(new_n2752_), .ZN(new_n2753_));
  NOR3_X1    g01749(.A1(new_n2744_), .A2(new_n2750_), .A3(new_n2753_), .ZN(new_n2754_));
  INV_X1     g01750(.I(\A[415] ), .ZN(new_n2755_));
  INV_X1     g01751(.I(\A[416] ), .ZN(new_n2756_));
  NAND2_X1   g01752(.A1(new_n2756_), .A2(\A[417] ), .ZN(new_n2757_));
  INV_X1     g01753(.I(\A[417] ), .ZN(new_n2758_));
  NAND2_X1   g01754(.A1(new_n2758_), .A2(\A[416] ), .ZN(new_n2759_));
  AOI21_X1   g01755(.A1(new_n2757_), .A2(new_n2759_), .B(new_n2755_), .ZN(new_n2760_));
  NOR2_X1    g01756(.A1(\A[416] ), .A2(\A[417] ), .ZN(new_n2761_));
  INV_X1     g01757(.I(new_n2761_), .ZN(new_n2762_));
  NAND2_X1   g01758(.A1(\A[416] ), .A2(\A[417] ), .ZN(new_n2763_));
  AOI21_X1   g01759(.A1(new_n2762_), .A2(new_n2763_), .B(\A[415] ), .ZN(new_n2764_));
  NOR2_X1    g01760(.A1(new_n2764_), .A2(new_n2760_), .ZN(new_n2765_));
  INV_X1     g01761(.I(\A[418] ), .ZN(new_n2766_));
  INV_X1     g01762(.I(\A[419] ), .ZN(new_n2767_));
  NAND2_X1   g01763(.A1(new_n2767_), .A2(\A[420] ), .ZN(new_n2768_));
  INV_X1     g01764(.I(\A[420] ), .ZN(new_n2769_));
  NAND2_X1   g01765(.A1(new_n2769_), .A2(\A[419] ), .ZN(new_n2770_));
  AOI21_X1   g01766(.A1(new_n2768_), .A2(new_n2770_), .B(new_n2766_), .ZN(new_n2771_));
  NOR2_X1    g01767(.A1(\A[419] ), .A2(\A[420] ), .ZN(new_n2772_));
  INV_X1     g01768(.I(new_n2772_), .ZN(new_n2773_));
  NAND2_X1   g01769(.A1(\A[419] ), .A2(\A[420] ), .ZN(new_n2774_));
  AOI21_X1   g01770(.A1(new_n2773_), .A2(new_n2774_), .B(\A[418] ), .ZN(new_n2775_));
  NOR2_X1    g01771(.A1(new_n2775_), .A2(new_n2771_), .ZN(new_n2776_));
  AOI21_X1   g01772(.A1(new_n2766_), .A2(new_n2774_), .B(new_n2772_), .ZN(new_n2777_));
  AOI21_X1   g01773(.A1(new_n2755_), .A2(new_n2763_), .B(new_n2761_), .ZN(new_n2778_));
  NAND2_X1   g01774(.A1(new_n2777_), .A2(new_n2778_), .ZN(new_n2779_));
  INV_X1     g01775(.I(new_n2779_), .ZN(new_n2780_));
  NAND2_X1   g01776(.A1(new_n2738_), .A2(new_n2754_), .ZN(new_n2781_));
  AOI21_X1   g01777(.A1(new_n2713_), .A2(new_n2709_), .B(new_n2781_), .ZN(new_n2782_));
  NOR2_X1    g01778(.A1(new_n2704_), .A2(new_n2782_), .ZN(new_n2783_));
  OAI21_X1   g01779(.A1(new_n2638_), .A2(new_n2639_), .B(new_n2600_), .ZN(new_n2784_));
  NAND3_X1   g01780(.A1(new_n2622_), .A2(new_n2636_), .A3(new_n2601_), .ZN(new_n2785_));
  NAND2_X1   g01781(.A1(new_n2784_), .A2(new_n2785_), .ZN(new_n2786_));
  AOI21_X1   g01782(.A1(new_n2682_), .A2(new_n2683_), .B(new_n2681_), .ZN(new_n2787_));
  NOR3_X1    g01783(.A1(new_n2679_), .A2(new_n2667_), .A3(new_n2645_), .ZN(new_n2788_));
  NOR2_X1    g01784(.A1(new_n2788_), .A2(new_n2787_), .ZN(new_n2789_));
  NOR3_X1    g01785(.A1(new_n2700_), .A2(new_n2701_), .A3(new_n2710_), .ZN(new_n2790_));
  AOI21_X1   g01786(.A1(new_n2789_), .A2(new_n2790_), .B(new_n2786_), .ZN(new_n2791_));
  NOR2_X1    g01787(.A1(new_n2711_), .A2(new_n2712_), .ZN(new_n2792_));
  NOR2_X1    g01788(.A1(new_n2708_), .A2(new_n2705_), .ZN(new_n2793_));
  NAND2_X1   g01789(.A1(new_n2744_), .A2(new_n2750_), .ZN(new_n2794_));
  INV_X1     g01790(.I(new_n2737_), .ZN(new_n2795_));
  NAND2_X1   g01791(.A1(new_n2795_), .A2(new_n2794_), .ZN(new_n2796_));
  INV_X1     g01792(.I(new_n2754_), .ZN(new_n2797_));
  NOR2_X1    g01793(.A1(new_n2796_), .A2(new_n2797_), .ZN(new_n2798_));
  OAI21_X1   g01794(.A1(new_n2792_), .A2(new_n2793_), .B(new_n2798_), .ZN(new_n2799_));
  NOR2_X1    g01795(.A1(new_n2791_), .A2(new_n2799_), .ZN(new_n2800_));
  NOR2_X1    g01796(.A1(new_n2783_), .A2(new_n2800_), .ZN(new_n2801_));
  NAND2_X1   g01797(.A1(new_n2704_), .A2(new_n2782_), .ZN(new_n2802_));
  INV_X1     g01798(.I(new_n2752_), .ZN(new_n2803_));
  NOR2_X1    g01799(.A1(new_n2737_), .A2(new_n2803_), .ZN(new_n2804_));
  NOR3_X1    g01800(.A1(new_n2744_), .A2(new_n2750_), .A3(new_n2752_), .ZN(new_n2805_));
  OAI21_X1   g01801(.A1(new_n2804_), .A2(new_n2805_), .B(new_n2751_), .ZN(new_n2806_));
  INV_X1     g01802(.I(new_n2751_), .ZN(new_n2807_));
  OAI21_X1   g01803(.A1(new_n2744_), .A2(new_n2750_), .B(new_n2752_), .ZN(new_n2808_));
  NAND3_X1   g01804(.A1(new_n2724_), .A2(new_n2735_), .A3(new_n2803_), .ZN(new_n2809_));
  NAND3_X1   g01805(.A1(new_n2808_), .A2(new_n2809_), .A3(new_n2807_), .ZN(new_n2810_));
  NAND2_X1   g01806(.A1(new_n2806_), .A2(new_n2810_), .ZN(new_n2811_));
  NOR2_X1    g01807(.A1(new_n2758_), .A2(\A[416] ), .ZN(new_n2812_));
  NOR2_X1    g01808(.A1(new_n2756_), .A2(\A[417] ), .ZN(new_n2813_));
  OAI21_X1   g01809(.A1(new_n2812_), .A2(new_n2813_), .B(\A[415] ), .ZN(new_n2814_));
  INV_X1     g01810(.I(new_n2763_), .ZN(new_n2815_));
  OAI21_X1   g01811(.A1(new_n2815_), .A2(new_n2761_), .B(new_n2755_), .ZN(new_n2816_));
  NAND2_X1   g01812(.A1(new_n2814_), .A2(new_n2816_), .ZN(new_n2817_));
  NOR2_X1    g01813(.A1(new_n2769_), .A2(\A[419] ), .ZN(new_n2818_));
  NOR2_X1    g01814(.A1(new_n2767_), .A2(\A[420] ), .ZN(new_n2819_));
  OAI21_X1   g01815(.A1(new_n2818_), .A2(new_n2819_), .B(\A[418] ), .ZN(new_n2820_));
  INV_X1     g01816(.I(new_n2774_), .ZN(new_n2821_));
  OAI21_X1   g01817(.A1(new_n2821_), .A2(new_n2772_), .B(new_n2766_), .ZN(new_n2822_));
  NAND2_X1   g01818(.A1(new_n2820_), .A2(new_n2822_), .ZN(new_n2823_));
  NOR3_X1    g01819(.A1(new_n2817_), .A2(new_n2823_), .A3(new_n2779_), .ZN(new_n2824_));
  NOR4_X1    g01820(.A1(new_n2760_), .A2(new_n2764_), .A3(new_n2775_), .A4(new_n2771_), .ZN(new_n2825_));
  NOR2_X1    g01821(.A1(new_n2765_), .A2(new_n2776_), .ZN(new_n2826_));
  NOR2_X1    g01822(.A1(new_n2826_), .A2(new_n2825_), .ZN(new_n2827_));
  INV_X1     g01823(.I(new_n2753_), .ZN(new_n2828_));
  NAND2_X1   g01824(.A1(new_n2807_), .A2(new_n2803_), .ZN(new_n2829_));
  AOI21_X1   g01825(.A1(new_n2737_), .A2(new_n2829_), .B(new_n2828_), .ZN(new_n2830_));
  NAND4_X1   g01826(.A1(new_n2738_), .A2(new_n2827_), .A3(new_n2830_), .A4(new_n2824_), .ZN(new_n2831_));
  NOR2_X1    g01827(.A1(new_n2811_), .A2(new_n2831_), .ZN(new_n2832_));
  INV_X1     g01828(.I(new_n2778_), .ZN(new_n2833_));
  NOR2_X1    g01829(.A1(new_n2825_), .A2(new_n2833_), .ZN(new_n2834_));
  NOR3_X1    g01830(.A1(new_n2817_), .A2(new_n2823_), .A3(new_n2778_), .ZN(new_n2835_));
  OAI21_X1   g01831(.A1(new_n2834_), .A2(new_n2835_), .B(new_n2777_), .ZN(new_n2836_));
  INV_X1     g01832(.I(new_n2777_), .ZN(new_n2837_));
  OAI21_X1   g01833(.A1(new_n2817_), .A2(new_n2823_), .B(new_n2778_), .ZN(new_n2838_));
  NAND2_X1   g01834(.A1(new_n2825_), .A2(new_n2833_), .ZN(new_n2839_));
  NAND3_X1   g01835(.A1(new_n2839_), .A2(new_n2838_), .A3(new_n2837_), .ZN(new_n2840_));
  NAND2_X1   g01836(.A1(new_n2836_), .A2(new_n2840_), .ZN(new_n2841_));
  NAND2_X1   g01837(.A1(new_n2832_), .A2(new_n2841_), .ZN(new_n2842_));
  NAND4_X1   g01838(.A1(new_n2738_), .A2(new_n2827_), .A3(new_n2754_), .A4(new_n2824_), .ZN(new_n2843_));
  NAND2_X1   g01839(.A1(new_n2841_), .A2(new_n2843_), .ZN(new_n2844_));
  AOI21_X1   g01840(.A1(new_n2839_), .A2(new_n2838_), .B(new_n2837_), .ZN(new_n2845_));
  NOR3_X1    g01841(.A1(new_n2834_), .A2(new_n2835_), .A3(new_n2777_), .ZN(new_n2846_));
  NOR2_X1    g01842(.A1(new_n2846_), .A2(new_n2845_), .ZN(new_n2847_));
  NAND3_X1   g01843(.A1(new_n2795_), .A2(new_n2754_), .A3(new_n2794_), .ZN(new_n2848_));
  NAND2_X1   g01844(.A1(new_n2825_), .A2(new_n2780_), .ZN(new_n2849_));
  NOR4_X1    g01845(.A1(new_n2848_), .A2(new_n2825_), .A3(new_n2849_), .A4(new_n2826_), .ZN(new_n2850_));
  AOI21_X1   g01846(.A1(new_n2808_), .A2(new_n2809_), .B(new_n2807_), .ZN(new_n2851_));
  NOR3_X1    g01847(.A1(new_n2804_), .A2(new_n2805_), .A3(new_n2751_), .ZN(new_n2852_));
  NOR4_X1    g01848(.A1(new_n2736_), .A2(new_n2737_), .A3(new_n2807_), .A4(new_n2803_), .ZN(new_n2853_));
  NOR3_X1    g01849(.A1(new_n2852_), .A2(new_n2851_), .A3(new_n2853_), .ZN(new_n2854_));
  AOI21_X1   g01850(.A1(new_n2847_), .A2(new_n2850_), .B(new_n2854_), .ZN(new_n2855_));
  NAND4_X1   g01851(.A1(new_n2795_), .A2(new_n2794_), .A3(new_n2751_), .A4(new_n2752_), .ZN(new_n2856_));
  NAND3_X1   g01852(.A1(new_n2806_), .A2(new_n2856_), .A3(new_n2810_), .ZN(new_n2857_));
  NOR3_X1    g01853(.A1(new_n2857_), .A2(new_n2841_), .A3(new_n2843_), .ZN(new_n2858_));
  OAI21_X1   g01854(.A1(new_n2855_), .A2(new_n2858_), .B(new_n2844_), .ZN(new_n2859_));
  NAND2_X1   g01855(.A1(new_n2859_), .A2(new_n2842_), .ZN(new_n2860_));
  OAI21_X1   g01856(.A1(new_n2860_), .A2(new_n2801_), .B(new_n2802_), .ZN(new_n2861_));
  NOR4_X1    g01857(.A1(new_n2685_), .A2(new_n2700_), .A3(new_n2701_), .A4(new_n2702_), .ZN(new_n2862_));
  AOI21_X1   g01858(.A1(new_n2789_), .A2(new_n2790_), .B(new_n2641_), .ZN(new_n2863_));
  NOR2_X1    g01859(.A1(new_n2645_), .A2(new_n2649_), .ZN(new_n2864_));
  OAI21_X1   g01860(.A1(new_n2678_), .A2(new_n2864_), .B(new_n2694_), .ZN(new_n2865_));
  NOR2_X1    g01861(.A1(new_n2600_), .A2(new_n2605_), .ZN(new_n2866_));
  OAI21_X1   g01862(.A1(new_n2686_), .A2(new_n2866_), .B(new_n2697_), .ZN(new_n2867_));
  XOR2_X1    g01863(.A1(new_n2867_), .A2(new_n2865_), .Z(new_n2868_));
  NOR3_X1    g01864(.A1(new_n2863_), .A2(new_n2862_), .A3(new_n2868_), .ZN(new_n2869_));
  OR2_X2     g01865(.A1(new_n2811_), .A2(new_n2831_), .Z(new_n2870_));
  OAI21_X1   g01866(.A1(new_n2854_), .A2(new_n2843_), .B(new_n2841_), .ZN(new_n2871_));
  NOR3_X1    g01867(.A1(new_n2852_), .A2(new_n2851_), .A3(new_n2796_), .ZN(new_n2872_));
  INV_X1     g01868(.I(new_n2825_), .ZN(new_n2873_));
  NOR2_X1    g01869(.A1(new_n2777_), .A2(new_n2778_), .ZN(new_n2874_));
  OAI21_X1   g01870(.A1(new_n2873_), .A2(new_n2874_), .B(new_n2779_), .ZN(new_n2875_));
  INV_X1     g01871(.I(new_n2875_), .ZN(new_n2876_));
  OAI21_X1   g01872(.A1(new_n2872_), .A2(new_n2830_), .B(new_n2876_), .ZN(new_n2877_));
  INV_X1     g01873(.I(new_n2830_), .ZN(new_n2878_));
  NAND3_X1   g01874(.A1(new_n2806_), .A2(new_n2810_), .A3(new_n2738_), .ZN(new_n2879_));
  NAND3_X1   g01875(.A1(new_n2879_), .A2(new_n2878_), .A3(new_n2875_), .ZN(new_n2880_));
  NAND4_X1   g01876(.A1(new_n2870_), .A2(new_n2871_), .A3(new_n2877_), .A4(new_n2880_), .ZN(new_n2881_));
  NAND2_X1   g01877(.A1(new_n2881_), .A2(new_n2869_), .ZN(new_n2882_));
  NAND2_X1   g01878(.A1(new_n2789_), .A2(new_n2703_), .ZN(new_n2883_));
  OAI21_X1   g01879(.A1(new_n2696_), .A2(new_n2685_), .B(new_n2786_), .ZN(new_n2884_));
  XNOR2_X1   g01880(.A1(new_n2867_), .A2(new_n2865_), .ZN(new_n2885_));
  NAND3_X1   g01881(.A1(new_n2884_), .A2(new_n2885_), .A3(new_n2883_), .ZN(new_n2886_));
  NAND2_X1   g01882(.A1(new_n2857_), .A2(new_n2850_), .ZN(new_n2887_));
  AOI21_X1   g01883(.A1(new_n2887_), .A2(new_n2841_), .B(new_n2832_), .ZN(new_n2888_));
  AOI21_X1   g01884(.A1(new_n2879_), .A2(new_n2878_), .B(new_n2875_), .ZN(new_n2889_));
  NOR3_X1    g01885(.A1(new_n2872_), .A2(new_n2830_), .A3(new_n2876_), .ZN(new_n2890_));
  NOR2_X1    g01886(.A1(new_n2890_), .A2(new_n2889_), .ZN(new_n2891_));
  NAND3_X1   g01887(.A1(new_n2886_), .A2(new_n2888_), .A3(new_n2891_), .ZN(new_n2892_));
  NAND2_X1   g01888(.A1(new_n2882_), .A2(new_n2892_), .ZN(new_n2893_));
  NAND2_X1   g01889(.A1(new_n2893_), .A2(new_n2861_), .ZN(new_n2894_));
  NAND2_X1   g01890(.A1(new_n2791_), .A2(new_n2799_), .ZN(new_n2895_));
  NAND2_X1   g01891(.A1(new_n2704_), .A2(new_n2782_), .ZN(new_n2896_));
  NAND2_X1   g01892(.A1(new_n2896_), .A2(new_n2895_), .ZN(new_n2897_));
  OAI21_X1   g01893(.A1(new_n2841_), .A2(new_n2843_), .B(new_n2857_), .ZN(new_n2898_));
  NAND3_X1   g01894(.A1(new_n2850_), .A2(new_n2854_), .A3(new_n2847_), .ZN(new_n2899_));
  NAND2_X1   g01895(.A1(new_n2898_), .A2(new_n2899_), .ZN(new_n2900_));
  AOI22_X1   g01896(.A1(new_n2900_), .A2(new_n2844_), .B1(new_n2832_), .B2(new_n2841_), .ZN(new_n2901_));
  OAI21_X1   g01897(.A1(new_n2901_), .A2(new_n2704_), .B(new_n2897_), .ZN(new_n2902_));
  NAND2_X1   g01898(.A1(new_n2881_), .A2(new_n2886_), .ZN(new_n2903_));
  NAND3_X1   g01899(.A1(new_n2869_), .A2(new_n2888_), .A3(new_n2891_), .ZN(new_n2904_));
  NAND2_X1   g01900(.A1(new_n2903_), .A2(new_n2904_), .ZN(new_n2905_));
  NAND2_X1   g01901(.A1(new_n2902_), .A2(new_n2905_), .ZN(new_n2906_));
  NAND2_X1   g01902(.A1(new_n2906_), .A2(new_n2894_), .ZN(new_n2907_));
  INV_X1     g01903(.I(\A[460] ), .ZN(new_n2908_));
  NOR2_X1    g01904(.A1(\A[461] ), .A2(\A[462] ), .ZN(new_n2909_));
  NAND2_X1   g01905(.A1(\A[461] ), .A2(\A[462] ), .ZN(new_n2910_));
  AOI21_X1   g01906(.A1(new_n2908_), .A2(new_n2910_), .B(new_n2909_), .ZN(new_n2911_));
  INV_X1     g01907(.I(new_n2911_), .ZN(new_n2912_));
  INV_X1     g01908(.I(\A[457] ), .ZN(new_n2913_));
  NOR2_X1    g01909(.A1(\A[458] ), .A2(\A[459] ), .ZN(new_n2914_));
  NAND2_X1   g01910(.A1(\A[458] ), .A2(\A[459] ), .ZN(new_n2915_));
  AOI21_X1   g01911(.A1(new_n2913_), .A2(new_n2915_), .B(new_n2914_), .ZN(new_n2916_));
  INV_X1     g01912(.I(\A[459] ), .ZN(new_n2917_));
  NOR2_X1    g01913(.A1(new_n2917_), .A2(\A[458] ), .ZN(new_n2918_));
  INV_X1     g01914(.I(\A[458] ), .ZN(new_n2919_));
  NOR2_X1    g01915(.A1(new_n2919_), .A2(\A[459] ), .ZN(new_n2920_));
  OAI21_X1   g01916(.A1(new_n2918_), .A2(new_n2920_), .B(\A[457] ), .ZN(new_n2921_));
  INV_X1     g01917(.I(new_n2915_), .ZN(new_n2922_));
  OAI21_X1   g01918(.A1(new_n2922_), .A2(new_n2914_), .B(new_n2913_), .ZN(new_n2923_));
  INV_X1     g01919(.I(\A[462] ), .ZN(new_n2924_));
  NOR2_X1    g01920(.A1(new_n2924_), .A2(\A[461] ), .ZN(new_n2925_));
  INV_X1     g01921(.I(\A[461] ), .ZN(new_n2926_));
  NOR2_X1    g01922(.A1(new_n2926_), .A2(\A[462] ), .ZN(new_n2927_));
  OAI21_X1   g01923(.A1(new_n2925_), .A2(new_n2927_), .B(\A[460] ), .ZN(new_n2928_));
  INV_X1     g01924(.I(new_n2910_), .ZN(new_n2929_));
  OAI21_X1   g01925(.A1(new_n2929_), .A2(new_n2909_), .B(new_n2908_), .ZN(new_n2930_));
  NAND4_X1   g01926(.A1(new_n2921_), .A2(new_n2923_), .A3(new_n2928_), .A4(new_n2930_), .ZN(new_n2931_));
  NAND2_X1   g01927(.A1(new_n2931_), .A2(new_n2916_), .ZN(new_n2932_));
  INV_X1     g01928(.I(new_n2916_), .ZN(new_n2933_));
  NAND2_X1   g01929(.A1(new_n2919_), .A2(\A[459] ), .ZN(new_n2934_));
  NAND2_X1   g01930(.A1(new_n2917_), .A2(\A[458] ), .ZN(new_n2935_));
  AOI21_X1   g01931(.A1(new_n2934_), .A2(new_n2935_), .B(new_n2913_), .ZN(new_n2936_));
  INV_X1     g01932(.I(new_n2914_), .ZN(new_n2937_));
  AOI21_X1   g01933(.A1(new_n2937_), .A2(new_n2915_), .B(\A[457] ), .ZN(new_n2938_));
  NOR2_X1    g01934(.A1(new_n2938_), .A2(new_n2936_), .ZN(new_n2939_));
  NAND2_X1   g01935(.A1(new_n2926_), .A2(\A[462] ), .ZN(new_n2940_));
  NAND2_X1   g01936(.A1(new_n2924_), .A2(\A[461] ), .ZN(new_n2941_));
  AOI21_X1   g01937(.A1(new_n2940_), .A2(new_n2941_), .B(new_n2908_), .ZN(new_n2942_));
  INV_X1     g01938(.I(new_n2909_), .ZN(new_n2943_));
  AOI21_X1   g01939(.A1(new_n2943_), .A2(new_n2910_), .B(\A[460] ), .ZN(new_n2944_));
  NOR2_X1    g01940(.A1(new_n2944_), .A2(new_n2942_), .ZN(new_n2945_));
  NAND3_X1   g01941(.A1(new_n2939_), .A2(new_n2945_), .A3(new_n2933_), .ZN(new_n2946_));
  AOI21_X1   g01942(.A1(new_n2932_), .A2(new_n2946_), .B(new_n2912_), .ZN(new_n2947_));
  NOR4_X1    g01943(.A1(new_n2936_), .A2(new_n2938_), .A3(new_n2944_), .A4(new_n2942_), .ZN(new_n2948_));
  NOR2_X1    g01944(.A1(new_n2948_), .A2(new_n2933_), .ZN(new_n2949_));
  NAND2_X1   g01945(.A1(new_n2921_), .A2(new_n2923_), .ZN(new_n2950_));
  NAND2_X1   g01946(.A1(new_n2928_), .A2(new_n2930_), .ZN(new_n2951_));
  NOR3_X1    g01947(.A1(new_n2950_), .A2(new_n2951_), .A3(new_n2916_), .ZN(new_n2952_));
  NOR3_X1    g01948(.A1(new_n2949_), .A2(new_n2952_), .A3(new_n2911_), .ZN(new_n2953_));
  INV_X1     g01949(.I(\A[453] ), .ZN(new_n2954_));
  NOR2_X1    g01950(.A1(new_n2954_), .A2(\A[452] ), .ZN(new_n2955_));
  INV_X1     g01951(.I(\A[452] ), .ZN(new_n2956_));
  NOR2_X1    g01952(.A1(new_n2956_), .A2(\A[453] ), .ZN(new_n2957_));
  OAI21_X1   g01953(.A1(new_n2955_), .A2(new_n2957_), .B(\A[451] ), .ZN(new_n2958_));
  INV_X1     g01954(.I(\A[451] ), .ZN(new_n2959_));
  NOR2_X1    g01955(.A1(\A[452] ), .A2(\A[453] ), .ZN(new_n2960_));
  NAND2_X1   g01956(.A1(\A[452] ), .A2(\A[453] ), .ZN(new_n2961_));
  INV_X1     g01957(.I(new_n2961_), .ZN(new_n2962_));
  OAI21_X1   g01958(.A1(new_n2962_), .A2(new_n2960_), .B(new_n2959_), .ZN(new_n2963_));
  NAND2_X1   g01959(.A1(new_n2958_), .A2(new_n2963_), .ZN(new_n2964_));
  INV_X1     g01960(.I(\A[454] ), .ZN(new_n2965_));
  INV_X1     g01961(.I(\A[455] ), .ZN(new_n2966_));
  NAND2_X1   g01962(.A1(new_n2966_), .A2(\A[456] ), .ZN(new_n2967_));
  INV_X1     g01963(.I(\A[456] ), .ZN(new_n2968_));
  NAND2_X1   g01964(.A1(new_n2968_), .A2(\A[455] ), .ZN(new_n2969_));
  AOI21_X1   g01965(.A1(new_n2967_), .A2(new_n2969_), .B(new_n2965_), .ZN(new_n2970_));
  NOR2_X1    g01966(.A1(\A[455] ), .A2(\A[456] ), .ZN(new_n2971_));
  INV_X1     g01967(.I(new_n2971_), .ZN(new_n2972_));
  NAND2_X1   g01968(.A1(\A[455] ), .A2(\A[456] ), .ZN(new_n2973_));
  AOI21_X1   g01969(.A1(new_n2972_), .A2(new_n2973_), .B(\A[454] ), .ZN(new_n2974_));
  NOR2_X1    g01970(.A1(new_n2974_), .A2(new_n2970_), .ZN(new_n2975_));
  NOR2_X1    g01971(.A1(new_n2975_), .A2(new_n2964_), .ZN(new_n2976_));
  NAND2_X1   g01972(.A1(new_n2956_), .A2(\A[453] ), .ZN(new_n2977_));
  NAND2_X1   g01973(.A1(new_n2954_), .A2(\A[452] ), .ZN(new_n2978_));
  AOI21_X1   g01974(.A1(new_n2977_), .A2(new_n2978_), .B(new_n2959_), .ZN(new_n2979_));
  INV_X1     g01975(.I(new_n2960_), .ZN(new_n2980_));
  AOI21_X1   g01976(.A1(new_n2980_), .A2(new_n2961_), .B(\A[451] ), .ZN(new_n2981_));
  NOR2_X1    g01977(.A1(new_n2981_), .A2(new_n2979_), .ZN(new_n2982_));
  NOR2_X1    g01978(.A1(new_n2968_), .A2(\A[455] ), .ZN(new_n2983_));
  NOR2_X1    g01979(.A1(new_n2966_), .A2(\A[456] ), .ZN(new_n2984_));
  OAI21_X1   g01980(.A1(new_n2983_), .A2(new_n2984_), .B(\A[454] ), .ZN(new_n2985_));
  INV_X1     g01981(.I(new_n2973_), .ZN(new_n2986_));
  OAI21_X1   g01982(.A1(new_n2986_), .A2(new_n2971_), .B(new_n2965_), .ZN(new_n2987_));
  NAND2_X1   g01983(.A1(new_n2985_), .A2(new_n2987_), .ZN(new_n2988_));
  NOR2_X1    g01984(.A1(new_n2982_), .A2(new_n2988_), .ZN(new_n2989_));
  NOR2_X1    g01985(.A1(new_n2945_), .A2(new_n2950_), .ZN(new_n2990_));
  NOR2_X1    g01986(.A1(new_n2939_), .A2(new_n2951_), .ZN(new_n2991_));
  OAI22_X1   g01987(.A1(new_n2976_), .A2(new_n2989_), .B1(new_n2990_), .B2(new_n2991_), .ZN(new_n2992_));
  NAND4_X1   g01988(.A1(new_n2958_), .A2(new_n2963_), .A3(new_n2985_), .A4(new_n2987_), .ZN(new_n2993_));
  AOI21_X1   g01989(.A1(new_n2965_), .A2(new_n2973_), .B(new_n2971_), .ZN(new_n2994_));
  AOI21_X1   g01990(.A1(new_n2959_), .A2(new_n2961_), .B(new_n2960_), .ZN(new_n2995_));
  NAND2_X1   g01991(.A1(new_n2994_), .A2(new_n2995_), .ZN(new_n2996_));
  NOR2_X1    g01992(.A1(new_n2993_), .A2(new_n2996_), .ZN(new_n2997_));
  NAND2_X1   g01993(.A1(new_n2911_), .A2(new_n2916_), .ZN(new_n2998_));
  INV_X1     g01994(.I(new_n2998_), .ZN(new_n2999_));
  OAI21_X1   g01995(.A1(new_n2939_), .A2(new_n2945_), .B(new_n2999_), .ZN(new_n3000_));
  NAND2_X1   g01996(.A1(new_n3000_), .A2(new_n2997_), .ZN(new_n3001_));
  NOR4_X1    g01997(.A1(new_n2947_), .A2(new_n2992_), .A3(new_n2953_), .A4(new_n3001_), .ZN(new_n3002_));
  NOR4_X1    g01998(.A1(new_n2979_), .A2(new_n2981_), .A3(new_n2974_), .A4(new_n2970_), .ZN(new_n3003_));
  INV_X1     g01999(.I(new_n2995_), .ZN(new_n3004_));
  NOR2_X1    g02000(.A1(new_n3003_), .A2(new_n3004_), .ZN(new_n3005_));
  NOR2_X1    g02001(.A1(new_n2993_), .A2(new_n2995_), .ZN(new_n3006_));
  OAI21_X1   g02002(.A1(new_n3005_), .A2(new_n3006_), .B(new_n2994_), .ZN(new_n3007_));
  INV_X1     g02003(.I(new_n2994_), .ZN(new_n3008_));
  NAND2_X1   g02004(.A1(new_n2993_), .A2(new_n2995_), .ZN(new_n3009_));
  NAND2_X1   g02005(.A1(new_n3003_), .A2(new_n3004_), .ZN(new_n3010_));
  NAND3_X1   g02006(.A1(new_n3010_), .A2(new_n3009_), .A3(new_n3008_), .ZN(new_n3011_));
  NAND2_X1   g02007(.A1(new_n3007_), .A2(new_n3011_), .ZN(new_n3012_));
  OAI21_X1   g02008(.A1(new_n2949_), .A2(new_n2952_), .B(new_n2911_), .ZN(new_n3013_));
  NAND3_X1   g02009(.A1(new_n2932_), .A2(new_n2946_), .A3(new_n2912_), .ZN(new_n3014_));
  NAND2_X1   g02010(.A1(new_n3013_), .A2(new_n3014_), .ZN(new_n3015_));
  NOR2_X1    g02011(.A1(new_n2976_), .A2(new_n2989_), .ZN(new_n3016_));
  NOR2_X1    g02012(.A1(new_n2990_), .A2(new_n2991_), .ZN(new_n3017_));
  INV_X1     g02013(.I(new_n2996_), .ZN(new_n3018_));
  NAND4_X1   g02014(.A1(new_n2948_), .A2(new_n3003_), .A3(new_n3018_), .A4(new_n2999_), .ZN(new_n3019_));
  NOR3_X1    g02015(.A1(new_n3016_), .A2(new_n3017_), .A3(new_n3019_), .ZN(new_n3020_));
  NOR2_X1    g02016(.A1(new_n3015_), .A2(new_n3020_), .ZN(new_n3021_));
  NOR3_X1    g02017(.A1(new_n3021_), .A2(new_n3002_), .A3(new_n3012_), .ZN(new_n3022_));
  NAND2_X1   g02018(.A1(new_n2982_), .A2(new_n2988_), .ZN(new_n3023_));
  NAND2_X1   g02019(.A1(new_n2975_), .A2(new_n2964_), .ZN(new_n3024_));
  NAND2_X1   g02020(.A1(new_n3023_), .A2(new_n3024_), .ZN(new_n3025_));
  NAND2_X1   g02021(.A1(new_n2939_), .A2(new_n2951_), .ZN(new_n3026_));
  NAND2_X1   g02022(.A1(new_n2945_), .A2(new_n2950_), .ZN(new_n3027_));
  NAND2_X1   g02023(.A1(new_n3026_), .A2(new_n3027_), .ZN(new_n3028_));
  NOR4_X1    g02024(.A1(new_n2931_), .A2(new_n2993_), .A3(new_n2996_), .A4(new_n2998_), .ZN(new_n3029_));
  NAND3_X1   g02025(.A1(new_n3025_), .A2(new_n3028_), .A3(new_n3029_), .ZN(new_n3030_));
  NAND2_X1   g02026(.A1(new_n3015_), .A2(new_n3030_), .ZN(new_n3031_));
  AOI22_X1   g02027(.A1(new_n3023_), .A2(new_n3024_), .B1(new_n3026_), .B2(new_n3027_), .ZN(new_n3032_));
  NAND4_X1   g02028(.A1(new_n3032_), .A2(new_n3013_), .A3(new_n3014_), .A4(new_n3029_), .ZN(new_n3033_));
  AOI21_X1   g02029(.A1(new_n3031_), .A2(new_n3033_), .B(new_n3012_), .ZN(new_n3034_));
  NOR2_X1    g02030(.A1(new_n3022_), .A2(new_n3034_), .ZN(new_n3035_));
  NAND2_X1   g02031(.A1(new_n3003_), .A2(new_n3018_), .ZN(new_n3036_));
  AOI21_X1   g02032(.A1(new_n2950_), .A2(new_n2951_), .B(new_n2998_), .ZN(new_n3037_));
  NOR2_X1    g02033(.A1(new_n3036_), .A2(new_n3037_), .ZN(new_n3038_));
  NAND4_X1   g02034(.A1(new_n3032_), .A2(new_n3013_), .A3(new_n3014_), .A4(new_n3038_), .ZN(new_n3039_));
  AOI21_X1   g02035(.A1(new_n3010_), .A2(new_n3009_), .B(new_n3008_), .ZN(new_n3040_));
  NOR3_X1    g02036(.A1(new_n3005_), .A2(new_n3006_), .A3(new_n2994_), .ZN(new_n3041_));
  NOR2_X1    g02037(.A1(new_n3040_), .A2(new_n3041_), .ZN(new_n3042_));
  NOR2_X1    g02038(.A1(new_n2953_), .A2(new_n2947_), .ZN(new_n3043_));
  NAND2_X1   g02039(.A1(new_n3043_), .A2(new_n3030_), .ZN(new_n3044_));
  NAND3_X1   g02040(.A1(new_n3044_), .A2(new_n3039_), .A3(new_n3042_), .ZN(new_n3045_));
  AOI22_X1   g02041(.A1(new_n3032_), .A2(new_n3029_), .B1(new_n3013_), .B2(new_n3014_), .ZN(new_n3046_));
  NOR4_X1    g02042(.A1(new_n2992_), .A2(new_n2953_), .A3(new_n2947_), .A4(new_n3019_), .ZN(new_n3047_));
  OAI21_X1   g02043(.A1(new_n3046_), .A2(new_n3047_), .B(new_n3042_), .ZN(new_n3048_));
  NOR2_X1    g02044(.A1(new_n2931_), .A2(new_n2998_), .ZN(new_n3049_));
  NAND2_X1   g02045(.A1(new_n3028_), .A2(new_n3049_), .ZN(new_n3050_));
  NOR2_X1    g02046(.A1(new_n3016_), .A2(new_n3036_), .ZN(new_n3051_));
  NAND2_X1   g02047(.A1(new_n3051_), .A2(new_n3050_), .ZN(new_n3052_));
  NOR3_X1    g02048(.A1(new_n3017_), .A2(new_n2931_), .A3(new_n2998_), .ZN(new_n3053_));
  NAND2_X1   g02049(.A1(new_n3025_), .A2(new_n2997_), .ZN(new_n3054_));
  NAND2_X1   g02050(.A1(new_n3053_), .A2(new_n3054_), .ZN(new_n3055_));
  INV_X1     g02051(.I(\A[450] ), .ZN(new_n3056_));
  NOR2_X1    g02052(.A1(new_n3056_), .A2(\A[449] ), .ZN(new_n3057_));
  INV_X1     g02053(.I(\A[449] ), .ZN(new_n3058_));
  NOR2_X1    g02054(.A1(new_n3058_), .A2(\A[450] ), .ZN(new_n3059_));
  OAI21_X1   g02055(.A1(new_n3057_), .A2(new_n3059_), .B(\A[448] ), .ZN(new_n3060_));
  INV_X1     g02056(.I(\A[448] ), .ZN(new_n3061_));
  NOR2_X1    g02057(.A1(\A[449] ), .A2(\A[450] ), .ZN(new_n3062_));
  NAND2_X1   g02058(.A1(\A[449] ), .A2(\A[450] ), .ZN(new_n3063_));
  INV_X1     g02059(.I(new_n3063_), .ZN(new_n3064_));
  OAI21_X1   g02060(.A1(new_n3064_), .A2(new_n3062_), .B(new_n3061_), .ZN(new_n3065_));
  NAND2_X1   g02061(.A1(new_n3060_), .A2(new_n3065_), .ZN(new_n3066_));
  AOI21_X1   g02062(.A1(new_n3061_), .A2(new_n3063_), .B(new_n3062_), .ZN(new_n3067_));
  NAND4_X1   g02063(.A1(new_n3067_), .A2(\A[445] ), .A3(\A[446] ), .A4(\A[447] ), .ZN(new_n3068_));
  NOR2_X1    g02064(.A1(new_n3066_), .A2(new_n3068_), .ZN(new_n3069_));
  INV_X1     g02065(.I(\A[445] ), .ZN(new_n3070_));
  INV_X1     g02066(.I(\A[446] ), .ZN(new_n3071_));
  NAND2_X1   g02067(.A1(new_n3071_), .A2(\A[447] ), .ZN(new_n3072_));
  INV_X1     g02068(.I(\A[447] ), .ZN(new_n3073_));
  NAND2_X1   g02069(.A1(new_n3073_), .A2(\A[446] ), .ZN(new_n3074_));
  AOI21_X1   g02070(.A1(new_n3072_), .A2(new_n3074_), .B(new_n3070_), .ZN(new_n3075_));
  NOR2_X1    g02071(.A1(\A[446] ), .A2(\A[447] ), .ZN(new_n3076_));
  INV_X1     g02072(.I(new_n3076_), .ZN(new_n3077_));
  NAND2_X1   g02073(.A1(\A[446] ), .A2(\A[447] ), .ZN(new_n3078_));
  AOI21_X1   g02074(.A1(new_n3077_), .A2(new_n3078_), .B(\A[445] ), .ZN(new_n3079_));
  NOR2_X1    g02075(.A1(new_n3079_), .A2(new_n3075_), .ZN(new_n3080_));
  NAND2_X1   g02076(.A1(new_n3080_), .A2(new_n3066_), .ZN(new_n3081_));
  NAND2_X1   g02077(.A1(new_n3058_), .A2(\A[450] ), .ZN(new_n3082_));
  NAND2_X1   g02078(.A1(new_n3056_), .A2(\A[449] ), .ZN(new_n3083_));
  AOI21_X1   g02079(.A1(new_n3082_), .A2(new_n3083_), .B(new_n3061_), .ZN(new_n3084_));
  INV_X1     g02080(.I(new_n3062_), .ZN(new_n3085_));
  AOI21_X1   g02081(.A1(new_n3085_), .A2(new_n3063_), .B(\A[448] ), .ZN(new_n3086_));
  NOR2_X1    g02082(.A1(new_n3086_), .A2(new_n3084_), .ZN(new_n3087_));
  NOR2_X1    g02083(.A1(new_n3073_), .A2(\A[446] ), .ZN(new_n3088_));
  NOR2_X1    g02084(.A1(new_n3071_), .A2(\A[447] ), .ZN(new_n3089_));
  OAI21_X1   g02085(.A1(new_n3088_), .A2(new_n3089_), .B(\A[445] ), .ZN(new_n3090_));
  INV_X1     g02086(.I(new_n3078_), .ZN(new_n3091_));
  OAI21_X1   g02087(.A1(new_n3091_), .A2(new_n3076_), .B(new_n3070_), .ZN(new_n3092_));
  NAND2_X1   g02088(.A1(new_n3090_), .A2(new_n3092_), .ZN(new_n3093_));
  NAND2_X1   g02089(.A1(new_n3087_), .A2(new_n3093_), .ZN(new_n3094_));
  NAND2_X1   g02090(.A1(new_n3081_), .A2(new_n3094_), .ZN(new_n3095_));
  INV_X1     g02091(.I(\A[439] ), .ZN(new_n3096_));
  INV_X1     g02092(.I(\A[440] ), .ZN(new_n3097_));
  NAND2_X1   g02093(.A1(new_n3097_), .A2(\A[441] ), .ZN(new_n3098_));
  INV_X1     g02094(.I(\A[441] ), .ZN(new_n3099_));
  NAND2_X1   g02095(.A1(new_n3099_), .A2(\A[440] ), .ZN(new_n3100_));
  AOI21_X1   g02096(.A1(new_n3098_), .A2(new_n3100_), .B(new_n3096_), .ZN(new_n3101_));
  NOR2_X1    g02097(.A1(\A[440] ), .A2(\A[441] ), .ZN(new_n3102_));
  INV_X1     g02098(.I(new_n3102_), .ZN(new_n3103_));
  NAND2_X1   g02099(.A1(\A[440] ), .A2(\A[441] ), .ZN(new_n3104_));
  AOI21_X1   g02100(.A1(new_n3103_), .A2(new_n3104_), .B(\A[439] ), .ZN(new_n3105_));
  NOR2_X1    g02101(.A1(new_n3105_), .A2(new_n3101_), .ZN(new_n3106_));
  INV_X1     g02102(.I(\A[442] ), .ZN(new_n3107_));
  INV_X1     g02103(.I(\A[443] ), .ZN(new_n3108_));
  NAND2_X1   g02104(.A1(new_n3108_), .A2(\A[444] ), .ZN(new_n3109_));
  INV_X1     g02105(.I(\A[444] ), .ZN(new_n3110_));
  NAND2_X1   g02106(.A1(new_n3110_), .A2(\A[443] ), .ZN(new_n3111_));
  AOI21_X1   g02107(.A1(new_n3109_), .A2(new_n3111_), .B(new_n3107_), .ZN(new_n3112_));
  NOR2_X1    g02108(.A1(\A[443] ), .A2(\A[444] ), .ZN(new_n3113_));
  INV_X1     g02109(.I(new_n3113_), .ZN(new_n3114_));
  NAND2_X1   g02110(.A1(\A[443] ), .A2(\A[444] ), .ZN(new_n3115_));
  AOI21_X1   g02111(.A1(new_n3114_), .A2(new_n3115_), .B(\A[442] ), .ZN(new_n3116_));
  NOR2_X1    g02112(.A1(new_n3116_), .A2(new_n3112_), .ZN(new_n3117_));
  AOI21_X1   g02113(.A1(new_n3107_), .A2(new_n3115_), .B(new_n3113_), .ZN(new_n3118_));
  AOI21_X1   g02114(.A1(new_n3096_), .A2(new_n3104_), .B(new_n3102_), .ZN(new_n3119_));
  NAND2_X1   g02115(.A1(new_n3118_), .A2(new_n3119_), .ZN(new_n3120_));
  NAND2_X1   g02116(.A1(new_n3095_), .A2(new_n3069_), .ZN(new_n3122_));
  AOI21_X1   g02117(.A1(new_n3055_), .A2(new_n3052_), .B(new_n3122_), .ZN(new_n3123_));
  AOI21_X1   g02118(.A1(new_n3045_), .A2(new_n3048_), .B(new_n3123_), .ZN(new_n3124_));
  NOR2_X1    g02119(.A1(new_n3053_), .A2(new_n3054_), .ZN(new_n3125_));
  NOR2_X1    g02120(.A1(new_n3051_), .A2(new_n3050_), .ZN(new_n3126_));
  INV_X1     g02121(.I(new_n3122_), .ZN(new_n3127_));
  OAI21_X1   g02122(.A1(new_n3125_), .A2(new_n3126_), .B(new_n3127_), .ZN(new_n3128_));
  NOR3_X1    g02123(.A1(new_n3022_), .A2(new_n3034_), .A3(new_n3128_), .ZN(new_n3129_));
  NOR4_X1    g02124(.A1(new_n3101_), .A2(new_n3105_), .A3(new_n3116_), .A4(new_n3112_), .ZN(new_n3130_));
  INV_X1     g02125(.I(new_n3119_), .ZN(new_n3131_));
  NOR2_X1    g02126(.A1(new_n3130_), .A2(new_n3131_), .ZN(new_n3132_));
  NOR2_X1    g02127(.A1(new_n3099_), .A2(\A[440] ), .ZN(new_n3133_));
  NOR2_X1    g02128(.A1(new_n3097_), .A2(\A[441] ), .ZN(new_n3134_));
  OAI21_X1   g02129(.A1(new_n3133_), .A2(new_n3134_), .B(\A[439] ), .ZN(new_n3135_));
  INV_X1     g02130(.I(new_n3104_), .ZN(new_n3136_));
  OAI21_X1   g02131(.A1(new_n3136_), .A2(new_n3102_), .B(new_n3096_), .ZN(new_n3137_));
  NAND2_X1   g02132(.A1(new_n3135_), .A2(new_n3137_), .ZN(new_n3138_));
  NOR2_X1    g02133(.A1(new_n3110_), .A2(\A[443] ), .ZN(new_n3139_));
  NOR2_X1    g02134(.A1(new_n3108_), .A2(\A[444] ), .ZN(new_n3140_));
  OAI21_X1   g02135(.A1(new_n3139_), .A2(new_n3140_), .B(\A[442] ), .ZN(new_n3141_));
  INV_X1     g02136(.I(new_n3115_), .ZN(new_n3142_));
  OAI21_X1   g02137(.A1(new_n3142_), .A2(new_n3113_), .B(new_n3107_), .ZN(new_n3143_));
  NAND2_X1   g02138(.A1(new_n3141_), .A2(new_n3143_), .ZN(new_n3144_));
  NOR3_X1    g02139(.A1(new_n3138_), .A2(new_n3144_), .A3(new_n3119_), .ZN(new_n3145_));
  OAI21_X1   g02140(.A1(new_n3132_), .A2(new_n3145_), .B(new_n3118_), .ZN(new_n3146_));
  INV_X1     g02141(.I(new_n3118_), .ZN(new_n3147_));
  OAI21_X1   g02142(.A1(new_n3138_), .A2(new_n3144_), .B(new_n3119_), .ZN(new_n3148_));
  NAND3_X1   g02143(.A1(new_n3106_), .A2(new_n3117_), .A3(new_n3131_), .ZN(new_n3149_));
  NAND3_X1   g02144(.A1(new_n3148_), .A2(new_n3149_), .A3(new_n3147_), .ZN(new_n3150_));
  NAND2_X1   g02145(.A1(new_n3146_), .A2(new_n3150_), .ZN(new_n3151_));
  NOR3_X1    g02146(.A1(new_n3138_), .A2(new_n3144_), .A3(new_n3120_), .ZN(new_n3152_));
  INV_X1     g02147(.I(new_n3152_), .ZN(new_n3153_));
  AOI21_X1   g02148(.A1(new_n3070_), .A2(new_n3078_), .B(new_n3076_), .ZN(new_n3154_));
  INV_X1     g02149(.I(new_n3154_), .ZN(new_n3155_));
  AOI21_X1   g02150(.A1(new_n3087_), .A2(new_n3080_), .B(new_n3155_), .ZN(new_n3156_));
  NOR3_X1    g02151(.A1(new_n3066_), .A2(new_n3093_), .A3(new_n3154_), .ZN(new_n3157_));
  OAI21_X1   g02152(.A1(new_n3156_), .A2(new_n3157_), .B(new_n3067_), .ZN(new_n3158_));
  INV_X1     g02153(.I(new_n3067_), .ZN(new_n3159_));
  OAI21_X1   g02154(.A1(new_n3066_), .A2(new_n3093_), .B(new_n3154_), .ZN(new_n3160_));
  NAND3_X1   g02155(.A1(new_n3087_), .A2(new_n3080_), .A3(new_n3155_), .ZN(new_n3161_));
  NAND3_X1   g02156(.A1(new_n3160_), .A2(new_n3161_), .A3(new_n3159_), .ZN(new_n3162_));
  NAND2_X1   g02157(.A1(new_n3158_), .A2(new_n3162_), .ZN(new_n3163_));
  NAND2_X1   g02158(.A1(new_n3106_), .A2(new_n3144_), .ZN(new_n3164_));
  NAND2_X1   g02159(.A1(new_n3117_), .A2(new_n3138_), .ZN(new_n3165_));
  NAND2_X1   g02160(.A1(new_n3164_), .A2(new_n3165_), .ZN(new_n3166_));
  NAND2_X1   g02161(.A1(new_n3095_), .A2(new_n3166_), .ZN(new_n3167_));
  NAND2_X1   g02162(.A1(new_n3067_), .A2(new_n3154_), .ZN(new_n3168_));
  AOI21_X1   g02163(.A1(new_n3066_), .A2(new_n3093_), .B(new_n3168_), .ZN(new_n3169_));
  NOR4_X1    g02164(.A1(new_n3163_), .A2(new_n3153_), .A3(new_n3167_), .A4(new_n3169_), .ZN(new_n3170_));
  XOR2_X1    g02165(.A1(new_n3087_), .A2(new_n3093_), .Z(new_n3171_));
  NOR2_X1    g02166(.A1(new_n3117_), .A2(new_n3138_), .ZN(new_n3172_));
  NOR2_X1    g02167(.A1(new_n3106_), .A2(new_n3144_), .ZN(new_n3173_));
  NOR2_X1    g02168(.A1(new_n3172_), .A2(new_n3173_), .ZN(new_n3174_));
  NAND2_X1   g02169(.A1(new_n3152_), .A2(new_n3069_), .ZN(new_n3175_));
  NOR3_X1    g02170(.A1(new_n3171_), .A2(new_n3174_), .A3(new_n3175_), .ZN(new_n3176_));
  NAND2_X1   g02171(.A1(new_n3176_), .A2(new_n3151_), .ZN(new_n3177_));
  AOI21_X1   g02172(.A1(new_n3160_), .A2(new_n3161_), .B(new_n3159_), .ZN(new_n3178_));
  NOR3_X1    g02173(.A1(new_n3156_), .A2(new_n3157_), .A3(new_n3067_), .ZN(new_n3179_));
  NOR2_X1    g02174(.A1(new_n3179_), .A2(new_n3178_), .ZN(new_n3180_));
  OAI21_X1   g02175(.A1(new_n3151_), .A2(new_n3176_), .B(new_n3180_), .ZN(new_n3181_));
  AOI21_X1   g02176(.A1(new_n3148_), .A2(new_n3149_), .B(new_n3147_), .ZN(new_n3182_));
  NOR3_X1    g02177(.A1(new_n3132_), .A2(new_n3145_), .A3(new_n3118_), .ZN(new_n3183_));
  NOR2_X1    g02178(.A1(new_n3183_), .A2(new_n3182_), .ZN(new_n3184_));
  NAND4_X1   g02179(.A1(new_n3095_), .A2(new_n3166_), .A3(new_n3069_), .A4(new_n3152_), .ZN(new_n3185_));
  NAND3_X1   g02180(.A1(new_n3184_), .A2(new_n3185_), .A3(new_n3163_), .ZN(new_n3186_));
  NAND2_X1   g02181(.A1(new_n3181_), .A2(new_n3186_), .ZN(new_n3187_));
  AOI22_X1   g02182(.A1(new_n3187_), .A2(new_n3177_), .B1(new_n3151_), .B2(new_n3170_), .ZN(new_n3188_));
  OAI22_X1   g02183(.A1(new_n3188_), .A2(new_n3035_), .B1(new_n3129_), .B2(new_n3124_), .ZN(new_n3189_));
  OAI21_X1   g02184(.A1(new_n2911_), .A2(new_n2916_), .B(new_n2948_), .ZN(new_n3190_));
  NAND2_X1   g02185(.A1(new_n3190_), .A2(new_n2998_), .ZN(new_n3191_));
  OAI21_X1   g02186(.A1(new_n2994_), .A2(new_n2995_), .B(new_n3003_), .ZN(new_n3192_));
  NAND2_X1   g02187(.A1(new_n3192_), .A2(new_n2996_), .ZN(new_n3193_));
  INV_X1     g02188(.I(new_n3193_), .ZN(new_n3194_));
  OAI21_X1   g02189(.A1(new_n3015_), .A2(new_n3020_), .B(new_n3012_), .ZN(new_n3195_));
  AOI21_X1   g02190(.A1(new_n3195_), .A2(new_n3039_), .B(new_n3194_), .ZN(new_n3196_));
  AOI21_X1   g02191(.A1(new_n3043_), .A2(new_n3030_), .B(new_n3042_), .ZN(new_n3197_));
  NOR3_X1    g02192(.A1(new_n3197_), .A2(new_n3002_), .A3(new_n3193_), .ZN(new_n3198_));
  OAI21_X1   g02193(.A1(new_n3198_), .A2(new_n3196_), .B(new_n3191_), .ZN(new_n3199_));
  INV_X1     g02194(.I(new_n3191_), .ZN(new_n3200_));
  OAI21_X1   g02195(.A1(new_n3197_), .A2(new_n3002_), .B(new_n3193_), .ZN(new_n3201_));
  NAND3_X1   g02196(.A1(new_n3195_), .A2(new_n3039_), .A3(new_n3194_), .ZN(new_n3202_));
  NAND3_X1   g02197(.A1(new_n3201_), .A2(new_n3202_), .A3(new_n3200_), .ZN(new_n3203_));
  NAND2_X1   g02198(.A1(new_n3199_), .A2(new_n3203_), .ZN(new_n3204_));
  NAND2_X1   g02199(.A1(new_n3159_), .A2(new_n3155_), .ZN(new_n3205_));
  NAND3_X1   g02200(.A1(new_n3205_), .A2(new_n3087_), .A3(new_n3080_), .ZN(new_n3206_));
  NAND2_X1   g02201(.A1(new_n3206_), .A2(new_n3168_), .ZN(new_n3207_));
  INV_X1     g02202(.I(new_n3207_), .ZN(new_n3208_));
  OAI21_X1   g02203(.A1(new_n3118_), .A2(new_n3119_), .B(new_n3130_), .ZN(new_n3209_));
  NAND2_X1   g02204(.A1(new_n3209_), .A2(new_n3120_), .ZN(new_n3210_));
  AOI21_X1   g02205(.A1(new_n3180_), .A2(new_n3185_), .B(new_n3184_), .ZN(new_n3211_));
  OAI21_X1   g02206(.A1(new_n3211_), .A2(new_n3170_), .B(new_n3210_), .ZN(new_n3212_));
  NOR2_X1    g02207(.A1(new_n3171_), .A2(new_n3174_), .ZN(new_n3213_));
  NOR2_X1    g02208(.A1(new_n3153_), .A2(new_n3169_), .ZN(new_n3214_));
  NAND3_X1   g02209(.A1(new_n3180_), .A2(new_n3213_), .A3(new_n3214_), .ZN(new_n3215_));
  INV_X1     g02210(.I(new_n3210_), .ZN(new_n3216_));
  OAI21_X1   g02211(.A1(new_n3163_), .A2(new_n3176_), .B(new_n3151_), .ZN(new_n3217_));
  NAND3_X1   g02212(.A1(new_n3217_), .A2(new_n3215_), .A3(new_n3216_), .ZN(new_n3218_));
  AOI21_X1   g02213(.A1(new_n3212_), .A2(new_n3218_), .B(new_n3208_), .ZN(new_n3219_));
  AOI21_X1   g02214(.A1(new_n3217_), .A2(new_n3215_), .B(new_n3216_), .ZN(new_n3220_));
  NOR3_X1    g02215(.A1(new_n3211_), .A2(new_n3170_), .A3(new_n3210_), .ZN(new_n3221_));
  NOR3_X1    g02216(.A1(new_n3221_), .A2(new_n3220_), .A3(new_n3207_), .ZN(new_n3222_));
  NOR2_X1    g02217(.A1(new_n3222_), .A2(new_n3219_), .ZN(new_n3223_));
  NAND2_X1   g02218(.A1(new_n3204_), .A2(new_n3223_), .ZN(new_n3224_));
  AOI21_X1   g02219(.A1(new_n3201_), .A2(new_n3202_), .B(new_n3200_), .ZN(new_n3225_));
  NOR3_X1    g02220(.A1(new_n3198_), .A2(new_n3196_), .A3(new_n3191_), .ZN(new_n3226_));
  NOR2_X1    g02221(.A1(new_n3226_), .A2(new_n3225_), .ZN(new_n3227_));
  OAI21_X1   g02222(.A1(new_n3221_), .A2(new_n3220_), .B(new_n3207_), .ZN(new_n3228_));
  NAND3_X1   g02223(.A1(new_n3212_), .A2(new_n3218_), .A3(new_n3208_), .ZN(new_n3229_));
  NAND2_X1   g02224(.A1(new_n3228_), .A2(new_n3229_), .ZN(new_n3230_));
  NAND2_X1   g02225(.A1(new_n3227_), .A2(new_n3230_), .ZN(new_n3231_));
  AOI21_X1   g02226(.A1(new_n3231_), .A2(new_n3224_), .B(new_n3189_), .ZN(new_n3232_));
  NAND2_X1   g02227(.A1(new_n3045_), .A2(new_n3048_), .ZN(new_n3233_));
  OAI21_X1   g02228(.A1(new_n3022_), .A2(new_n3034_), .B(new_n3128_), .ZN(new_n3234_));
  NAND3_X1   g02229(.A1(new_n3045_), .A2(new_n3123_), .A3(new_n3048_), .ZN(new_n3235_));
  NAND2_X1   g02230(.A1(new_n3170_), .A2(new_n3151_), .ZN(new_n3236_));
  AOI21_X1   g02231(.A1(new_n3184_), .A2(new_n3185_), .B(new_n3163_), .ZN(new_n3237_));
  NOR3_X1    g02232(.A1(new_n3180_), .A2(new_n3176_), .A3(new_n3151_), .ZN(new_n3238_));
  OAI21_X1   g02233(.A1(new_n3238_), .A2(new_n3237_), .B(new_n3177_), .ZN(new_n3239_));
  NAND2_X1   g02234(.A1(new_n3239_), .A2(new_n3236_), .ZN(new_n3240_));
  AOI22_X1   g02235(.A1(new_n3240_), .A2(new_n3233_), .B1(new_n3234_), .B2(new_n3235_), .ZN(new_n3241_));
  NAND4_X1   g02236(.A1(new_n3199_), .A2(new_n3203_), .A3(new_n3228_), .A4(new_n3229_), .ZN(new_n3242_));
  OAI22_X1   g02237(.A1(new_n3226_), .A2(new_n3225_), .B1(new_n3222_), .B2(new_n3219_), .ZN(new_n3243_));
  AOI21_X1   g02238(.A1(new_n3243_), .A2(new_n3242_), .B(new_n3241_), .ZN(new_n3244_));
  NOR3_X1    g02239(.A1(new_n3232_), .A2(new_n2907_), .A3(new_n3244_), .ZN(new_n3245_));
  NOR3_X1    g02240(.A1(new_n3240_), .A2(new_n3129_), .A3(new_n3124_), .ZN(new_n3246_));
  INV_X1     g02241(.I(new_n3246_), .ZN(new_n3247_));
  NOR2_X1    g02242(.A1(new_n3125_), .A2(new_n3126_), .ZN(new_n3248_));
  INV_X1     g02243(.I(new_n3069_), .ZN(new_n3249_));
  NOR2_X1    g02244(.A1(new_n3171_), .A2(new_n3249_), .ZN(new_n3250_));
  NOR2_X1    g02245(.A1(new_n3248_), .A2(new_n3250_), .ZN(new_n3251_));
  NAND2_X1   g02246(.A1(new_n3055_), .A2(new_n3052_), .ZN(new_n3252_));
  INV_X1     g02247(.I(new_n3250_), .ZN(new_n3253_));
  NOR2_X1    g02248(.A1(new_n3252_), .A2(new_n3253_), .ZN(new_n3254_));
  NOR2_X1    g02249(.A1(new_n2792_), .A2(new_n2793_), .ZN(new_n3255_));
  INV_X1     g02250(.I(new_n2848_), .ZN(new_n3256_));
  NOR2_X1    g02251(.A1(new_n3255_), .A2(new_n3256_), .ZN(new_n3257_));
  NAND2_X1   g02252(.A1(new_n2713_), .A2(new_n2709_), .ZN(new_n3258_));
  NOR2_X1    g02253(.A1(new_n3258_), .A2(new_n2848_), .ZN(new_n3259_));
  NOR4_X1    g02254(.A1(new_n3251_), .A2(new_n3254_), .A3(new_n3257_), .A4(new_n3259_), .ZN(new_n3260_));
  OR2_X2     g02255(.A1(new_n3246_), .A2(new_n3260_), .Z(new_n3261_));
  NAND2_X1   g02256(.A1(new_n3246_), .A2(new_n3260_), .ZN(new_n3262_));
  NAND3_X1   g02257(.A1(new_n2897_), .A2(new_n2842_), .A3(new_n2859_), .ZN(new_n3263_));
  NAND2_X1   g02258(.A1(new_n2860_), .A2(new_n2801_), .ZN(new_n3264_));
  NAND2_X1   g02259(.A1(new_n3264_), .A2(new_n3263_), .ZN(new_n3265_));
  AOI22_X1   g02260(.A1(new_n3261_), .A2(new_n3262_), .B1(new_n3247_), .B2(new_n3265_), .ZN(new_n3266_));
  OAI21_X1   g02261(.A1(new_n3232_), .A2(new_n3244_), .B(new_n2907_), .ZN(new_n3267_));
  AOI21_X1   g02262(.A1(new_n3267_), .A2(new_n3266_), .B(new_n3245_), .ZN(new_n3268_));
  NOR2_X1    g02263(.A1(new_n3200_), .A2(new_n3194_), .ZN(new_n3269_));
  NAND2_X1   g02264(.A1(new_n3195_), .A2(new_n3039_), .ZN(new_n3270_));
  AOI21_X1   g02265(.A1(new_n3200_), .A2(new_n3194_), .B(new_n3270_), .ZN(new_n3271_));
  NOR2_X1    g02266(.A1(new_n3271_), .A2(new_n3269_), .ZN(new_n3272_));
  AOI21_X1   g02267(.A1(new_n3227_), .A2(new_n3223_), .B(new_n3241_), .ZN(new_n3273_));
  NAND2_X1   g02268(.A1(new_n3217_), .A2(new_n3215_), .ZN(new_n3274_));
  XOR2_X1    g02269(.A1(new_n3193_), .A2(new_n3191_), .Z(new_n3275_));
  XOR2_X1    g02270(.A1(new_n3210_), .A2(new_n3207_), .Z(new_n3276_));
  NOR4_X1    g02271(.A1(new_n3270_), .A2(new_n3274_), .A3(new_n3276_), .A4(new_n3275_), .ZN(new_n3277_));
  INV_X1     g02272(.I(new_n3277_), .ZN(new_n3278_));
  NOR2_X1    g02273(.A1(new_n3216_), .A2(new_n3208_), .ZN(new_n3279_));
  AOI21_X1   g02274(.A1(new_n3208_), .A2(new_n3216_), .B(new_n3274_), .ZN(new_n3280_));
  NOR2_X1    g02275(.A1(new_n3280_), .A2(new_n3279_), .ZN(new_n3281_));
  INV_X1     g02276(.I(new_n3281_), .ZN(new_n3282_));
  OAI21_X1   g02277(.A1(new_n3273_), .A2(new_n3278_), .B(new_n3282_), .ZN(new_n3283_));
  NAND2_X1   g02278(.A1(new_n3242_), .A2(new_n3189_), .ZN(new_n3284_));
  NAND3_X1   g02279(.A1(new_n3284_), .A2(new_n3277_), .A3(new_n3281_), .ZN(new_n3285_));
  AOI21_X1   g02280(.A1(new_n3283_), .A2(new_n3285_), .B(new_n3272_), .ZN(new_n3286_));
  INV_X1     g02281(.I(new_n3272_), .ZN(new_n3287_));
  AOI21_X1   g02282(.A1(new_n3284_), .A2(new_n3277_), .B(new_n3281_), .ZN(new_n3288_));
  NOR3_X1    g02283(.A1(new_n3273_), .A2(new_n3278_), .A3(new_n3282_), .ZN(new_n3289_));
  NOR3_X1    g02284(.A1(new_n3289_), .A2(new_n3288_), .A3(new_n3287_), .ZN(new_n3290_));
  NAND2_X1   g02285(.A1(new_n2867_), .A2(new_n2865_), .ZN(new_n3291_));
  NOR2_X1    g02286(.A1(new_n2863_), .A2(new_n2862_), .ZN(new_n3292_));
  OAI21_X1   g02287(.A1(new_n2865_), .A2(new_n2867_), .B(new_n3292_), .ZN(new_n3293_));
  NAND2_X1   g02288(.A1(new_n3293_), .A2(new_n3291_), .ZN(new_n3294_));
  INV_X1     g02289(.I(new_n3294_), .ZN(new_n3295_));
  INV_X1     g02290(.I(new_n2881_), .ZN(new_n3296_));
  NAND3_X1   g02291(.A1(new_n2861_), .A2(new_n2869_), .A3(new_n3296_), .ZN(new_n3297_));
  OAI21_X1   g02292(.A1(new_n2872_), .A2(new_n2830_), .B(new_n2875_), .ZN(new_n3298_));
  NAND3_X1   g02293(.A1(new_n2879_), .A2(new_n2878_), .A3(new_n2876_), .ZN(new_n3299_));
  NAND2_X1   g02294(.A1(new_n2888_), .A2(new_n3299_), .ZN(new_n3300_));
  NAND2_X1   g02295(.A1(new_n3300_), .A2(new_n3298_), .ZN(new_n3301_));
  NAND2_X1   g02296(.A1(new_n3297_), .A2(new_n3301_), .ZN(new_n3302_));
  INV_X1     g02297(.I(new_n2904_), .ZN(new_n3303_));
  NAND3_X1   g02298(.A1(new_n3263_), .A2(new_n2802_), .A3(new_n2903_), .ZN(new_n3304_));
  INV_X1     g02299(.I(new_n3301_), .ZN(new_n3305_));
  NAND3_X1   g02300(.A1(new_n3304_), .A2(new_n3303_), .A3(new_n3305_), .ZN(new_n3306_));
  AOI21_X1   g02301(.A1(new_n3302_), .A2(new_n3306_), .B(new_n3295_), .ZN(new_n3307_));
  AOI21_X1   g02302(.A1(new_n3304_), .A2(new_n3303_), .B(new_n3305_), .ZN(new_n3308_));
  NOR4_X1    g02303(.A1(new_n2902_), .A2(new_n2886_), .A3(new_n2881_), .A4(new_n3301_), .ZN(new_n3309_));
  NOR3_X1    g02304(.A1(new_n3308_), .A2(new_n3309_), .A3(new_n3294_), .ZN(new_n3310_));
  NOR2_X1    g02305(.A1(new_n3307_), .A2(new_n3310_), .ZN(new_n3311_));
  OAI21_X1   g02306(.A1(new_n3286_), .A2(new_n3290_), .B(new_n3311_), .ZN(new_n3312_));
  OAI21_X1   g02307(.A1(new_n3289_), .A2(new_n3288_), .B(new_n3287_), .ZN(new_n3313_));
  NAND3_X1   g02308(.A1(new_n3283_), .A2(new_n3285_), .A3(new_n3272_), .ZN(new_n3314_));
  OAI21_X1   g02309(.A1(new_n3308_), .A2(new_n3309_), .B(new_n3294_), .ZN(new_n3315_));
  NAND3_X1   g02310(.A1(new_n3302_), .A2(new_n3306_), .A3(new_n3295_), .ZN(new_n3316_));
  NAND2_X1   g02311(.A1(new_n3316_), .A2(new_n3315_), .ZN(new_n3317_));
  NAND3_X1   g02312(.A1(new_n3317_), .A2(new_n3313_), .A3(new_n3314_), .ZN(new_n3318_));
  AOI21_X1   g02313(.A1(new_n3312_), .A2(new_n3318_), .B(new_n3268_), .ZN(new_n3319_));
  AND2_X2    g02314(.A1(new_n2882_), .A2(new_n2892_), .Z(new_n3320_));
  AND2_X2    g02315(.A1(new_n2903_), .A2(new_n2904_), .Z(new_n3321_));
  MUX2_X1    g02316(.I0(new_n3321_), .I1(new_n3320_), .S(new_n2861_), .Z(new_n3322_));
  NOR2_X1    g02317(.A1(new_n3227_), .A2(new_n3230_), .ZN(new_n3323_));
  NOR2_X1    g02318(.A1(new_n3204_), .A2(new_n3223_), .ZN(new_n3324_));
  OAI21_X1   g02319(.A1(new_n3323_), .A2(new_n3324_), .B(new_n3241_), .ZN(new_n3325_));
  INV_X1     g02320(.I(new_n3242_), .ZN(new_n3326_));
  AOI22_X1   g02321(.A1(new_n3199_), .A2(new_n3203_), .B1(new_n3228_), .B2(new_n3229_), .ZN(new_n3327_));
  OAI21_X1   g02322(.A1(new_n3326_), .A2(new_n3327_), .B(new_n3189_), .ZN(new_n3328_));
  NAND3_X1   g02323(.A1(new_n3322_), .A2(new_n3325_), .A3(new_n3328_), .ZN(new_n3329_));
  INV_X1     g02324(.I(new_n3266_), .ZN(new_n3330_));
  AOI21_X1   g02325(.A1(new_n3325_), .A2(new_n3328_), .B(new_n3322_), .ZN(new_n3331_));
  OAI21_X1   g02326(.A1(new_n3331_), .A2(new_n3330_), .B(new_n3329_), .ZN(new_n3332_));
  NAND4_X1   g02327(.A1(new_n3313_), .A2(new_n3314_), .A3(new_n3315_), .A4(new_n3316_), .ZN(new_n3333_));
  OAI21_X1   g02328(.A1(new_n3286_), .A2(new_n3290_), .B(new_n3317_), .ZN(new_n3334_));
  AOI21_X1   g02329(.A1(new_n3334_), .A2(new_n3333_), .B(new_n3332_), .ZN(new_n3335_));
  INV_X1     g02330(.I(\A[382] ), .ZN(new_n3336_));
  NOR2_X1    g02331(.A1(\A[383] ), .A2(\A[384] ), .ZN(new_n3337_));
  NAND2_X1   g02332(.A1(\A[383] ), .A2(\A[384] ), .ZN(new_n3338_));
  AOI21_X1   g02333(.A1(new_n3336_), .A2(new_n3338_), .B(new_n3337_), .ZN(new_n3339_));
  INV_X1     g02334(.I(new_n3339_), .ZN(new_n3340_));
  INV_X1     g02335(.I(\A[379] ), .ZN(new_n3341_));
  NOR2_X1    g02336(.A1(\A[380] ), .A2(\A[381] ), .ZN(new_n3342_));
  NAND2_X1   g02337(.A1(\A[380] ), .A2(\A[381] ), .ZN(new_n3343_));
  AOI21_X1   g02338(.A1(new_n3341_), .A2(new_n3343_), .B(new_n3342_), .ZN(new_n3344_));
  INV_X1     g02339(.I(\A[381] ), .ZN(new_n3345_));
  NOR2_X1    g02340(.A1(new_n3345_), .A2(\A[380] ), .ZN(new_n3346_));
  INV_X1     g02341(.I(\A[380] ), .ZN(new_n3347_));
  NOR2_X1    g02342(.A1(new_n3347_), .A2(\A[381] ), .ZN(new_n3348_));
  OAI21_X1   g02343(.A1(new_n3346_), .A2(new_n3348_), .B(\A[379] ), .ZN(new_n3349_));
  INV_X1     g02344(.I(new_n3343_), .ZN(new_n3350_));
  OAI21_X1   g02345(.A1(new_n3350_), .A2(new_n3342_), .B(new_n3341_), .ZN(new_n3351_));
  INV_X1     g02346(.I(\A[384] ), .ZN(new_n3352_));
  NOR2_X1    g02347(.A1(new_n3352_), .A2(\A[383] ), .ZN(new_n3353_));
  INV_X1     g02348(.I(\A[383] ), .ZN(new_n3354_));
  NOR2_X1    g02349(.A1(new_n3354_), .A2(\A[384] ), .ZN(new_n3355_));
  OAI21_X1   g02350(.A1(new_n3353_), .A2(new_n3355_), .B(\A[382] ), .ZN(new_n3356_));
  INV_X1     g02351(.I(new_n3338_), .ZN(new_n3357_));
  OAI21_X1   g02352(.A1(new_n3357_), .A2(new_n3337_), .B(new_n3336_), .ZN(new_n3358_));
  NAND4_X1   g02353(.A1(new_n3349_), .A2(new_n3351_), .A3(new_n3356_), .A4(new_n3358_), .ZN(new_n3359_));
  NAND2_X1   g02354(.A1(new_n3359_), .A2(new_n3344_), .ZN(new_n3360_));
  INV_X1     g02355(.I(new_n3344_), .ZN(new_n3361_));
  NAND2_X1   g02356(.A1(new_n3347_), .A2(\A[381] ), .ZN(new_n3362_));
  NAND2_X1   g02357(.A1(new_n3345_), .A2(\A[380] ), .ZN(new_n3363_));
  AOI21_X1   g02358(.A1(new_n3362_), .A2(new_n3363_), .B(new_n3341_), .ZN(new_n3364_));
  INV_X1     g02359(.I(new_n3342_), .ZN(new_n3365_));
  AOI21_X1   g02360(.A1(new_n3365_), .A2(new_n3343_), .B(\A[379] ), .ZN(new_n3366_));
  NAND2_X1   g02361(.A1(new_n3354_), .A2(\A[384] ), .ZN(new_n3367_));
  NAND2_X1   g02362(.A1(new_n3352_), .A2(\A[383] ), .ZN(new_n3368_));
  AOI21_X1   g02363(.A1(new_n3367_), .A2(new_n3368_), .B(new_n3336_), .ZN(new_n3369_));
  INV_X1     g02364(.I(new_n3337_), .ZN(new_n3370_));
  AOI21_X1   g02365(.A1(new_n3370_), .A2(new_n3338_), .B(\A[382] ), .ZN(new_n3371_));
  NOR4_X1    g02366(.A1(new_n3364_), .A2(new_n3366_), .A3(new_n3371_), .A4(new_n3369_), .ZN(new_n3372_));
  NAND2_X1   g02367(.A1(new_n3372_), .A2(new_n3361_), .ZN(new_n3373_));
  AOI21_X1   g02368(.A1(new_n3373_), .A2(new_n3360_), .B(new_n3340_), .ZN(new_n3374_));
  NOR2_X1    g02369(.A1(new_n3372_), .A2(new_n3361_), .ZN(new_n3375_));
  NOR2_X1    g02370(.A1(new_n3359_), .A2(new_n3344_), .ZN(new_n3376_));
  NOR3_X1    g02371(.A1(new_n3375_), .A2(new_n3376_), .A3(new_n3339_), .ZN(new_n3377_));
  NOR2_X1    g02372(.A1(new_n3374_), .A2(new_n3377_), .ZN(new_n3378_));
  INV_X1     g02373(.I(\A[388] ), .ZN(new_n3379_));
  NOR2_X1    g02374(.A1(\A[389] ), .A2(\A[390] ), .ZN(new_n3380_));
  NAND2_X1   g02375(.A1(\A[389] ), .A2(\A[390] ), .ZN(new_n3381_));
  AOI21_X1   g02376(.A1(new_n3379_), .A2(new_n3381_), .B(new_n3380_), .ZN(new_n3382_));
  INV_X1     g02377(.I(\A[385] ), .ZN(new_n3383_));
  NOR2_X1    g02378(.A1(\A[386] ), .A2(\A[387] ), .ZN(new_n3384_));
  NAND2_X1   g02379(.A1(\A[386] ), .A2(\A[387] ), .ZN(new_n3385_));
  AOI21_X1   g02380(.A1(new_n3383_), .A2(new_n3385_), .B(new_n3384_), .ZN(new_n3386_));
  NAND2_X1   g02381(.A1(new_n3382_), .A2(new_n3386_), .ZN(new_n3387_));
  INV_X1     g02382(.I(\A[386] ), .ZN(new_n3388_));
  NAND2_X1   g02383(.A1(new_n3388_), .A2(\A[387] ), .ZN(new_n3389_));
  INV_X1     g02384(.I(\A[387] ), .ZN(new_n3390_));
  NAND2_X1   g02385(.A1(new_n3390_), .A2(\A[386] ), .ZN(new_n3391_));
  AOI21_X1   g02386(.A1(new_n3389_), .A2(new_n3391_), .B(new_n3383_), .ZN(new_n3392_));
  INV_X1     g02387(.I(new_n3384_), .ZN(new_n3393_));
  AOI21_X1   g02388(.A1(new_n3393_), .A2(new_n3385_), .B(\A[385] ), .ZN(new_n3394_));
  NOR2_X1    g02389(.A1(new_n3394_), .A2(new_n3392_), .ZN(new_n3395_));
  INV_X1     g02390(.I(\A[390] ), .ZN(new_n3396_));
  NOR2_X1    g02391(.A1(new_n3396_), .A2(\A[389] ), .ZN(new_n3397_));
  INV_X1     g02392(.I(\A[389] ), .ZN(new_n3398_));
  NOR2_X1    g02393(.A1(new_n3398_), .A2(\A[390] ), .ZN(new_n3399_));
  OAI21_X1   g02394(.A1(new_n3397_), .A2(new_n3399_), .B(\A[388] ), .ZN(new_n3400_));
  AND2_X2    g02395(.A1(\A[389] ), .A2(\A[390] ), .Z(new_n3401_));
  OAI21_X1   g02396(.A1(new_n3401_), .A2(new_n3380_), .B(new_n3379_), .ZN(new_n3402_));
  NAND2_X1   g02397(.A1(new_n3400_), .A2(new_n3402_), .ZN(new_n3403_));
  NAND2_X1   g02398(.A1(new_n3395_), .A2(new_n3403_), .ZN(new_n3404_));
  NOR2_X1    g02399(.A1(new_n3390_), .A2(\A[386] ), .ZN(new_n3405_));
  NOR2_X1    g02400(.A1(new_n3388_), .A2(\A[387] ), .ZN(new_n3406_));
  OAI21_X1   g02401(.A1(new_n3405_), .A2(new_n3406_), .B(\A[385] ), .ZN(new_n3407_));
  INV_X1     g02402(.I(new_n3385_), .ZN(new_n3408_));
  OAI21_X1   g02403(.A1(new_n3408_), .A2(new_n3384_), .B(new_n3383_), .ZN(new_n3409_));
  NAND2_X1   g02404(.A1(new_n3407_), .A2(new_n3409_), .ZN(new_n3410_));
  NAND2_X1   g02405(.A1(new_n3398_), .A2(\A[390] ), .ZN(new_n3411_));
  NAND2_X1   g02406(.A1(new_n3396_), .A2(\A[389] ), .ZN(new_n3412_));
  AOI21_X1   g02407(.A1(new_n3411_), .A2(new_n3412_), .B(new_n3379_), .ZN(new_n3413_));
  INV_X1     g02408(.I(new_n3380_), .ZN(new_n3414_));
  AOI21_X1   g02409(.A1(new_n3414_), .A2(new_n3381_), .B(\A[388] ), .ZN(new_n3415_));
  NOR2_X1    g02410(.A1(new_n3415_), .A2(new_n3413_), .ZN(new_n3416_));
  NAND2_X1   g02411(.A1(new_n3416_), .A2(new_n3410_), .ZN(new_n3417_));
  AOI21_X1   g02412(.A1(new_n3417_), .A2(new_n3404_), .B(new_n3387_), .ZN(new_n3418_));
  INV_X1     g02413(.I(new_n3382_), .ZN(new_n3419_));
  NAND4_X1   g02414(.A1(new_n3407_), .A2(new_n3400_), .A3(new_n3409_), .A4(new_n3402_), .ZN(new_n3420_));
  NAND2_X1   g02415(.A1(new_n3420_), .A2(new_n3386_), .ZN(new_n3421_));
  INV_X1     g02416(.I(new_n3386_), .ZN(new_n3422_));
  NAND3_X1   g02417(.A1(new_n3395_), .A2(new_n3416_), .A3(new_n3422_), .ZN(new_n3423_));
  AOI21_X1   g02418(.A1(new_n3421_), .A2(new_n3423_), .B(new_n3419_), .ZN(new_n3424_));
  AOI21_X1   g02419(.A1(new_n3395_), .A2(new_n3416_), .B(new_n3422_), .ZN(new_n3425_));
  NOR3_X1    g02420(.A1(new_n3410_), .A2(new_n3403_), .A3(new_n3386_), .ZN(new_n3426_));
  NOR3_X1    g02421(.A1(new_n3425_), .A2(new_n3426_), .A3(new_n3382_), .ZN(new_n3427_));
  NOR2_X1    g02422(.A1(new_n3420_), .A2(new_n3387_), .ZN(new_n3428_));
  NOR4_X1    g02423(.A1(new_n3392_), .A2(new_n3394_), .A3(new_n3415_), .A4(new_n3413_), .ZN(new_n3429_));
  AOI22_X1   g02424(.A1(new_n3407_), .A2(new_n3409_), .B1(new_n3400_), .B2(new_n3402_), .ZN(new_n3430_));
  NOR2_X1    g02425(.A1(new_n3429_), .A2(new_n3430_), .ZN(new_n3431_));
  AOI22_X1   g02426(.A1(new_n3349_), .A2(new_n3351_), .B1(new_n3356_), .B2(new_n3358_), .ZN(new_n3432_));
  NOR2_X1    g02427(.A1(new_n3432_), .A2(new_n3372_), .ZN(new_n3433_));
  NAND2_X1   g02428(.A1(new_n3339_), .A2(new_n3344_), .ZN(new_n3434_));
  NOR2_X1    g02429(.A1(new_n3359_), .A2(new_n3434_), .ZN(new_n3435_));
  NAND4_X1   g02430(.A1(new_n3433_), .A2(new_n3431_), .A3(new_n3435_), .A4(new_n3428_), .ZN(new_n3436_));
  NOR4_X1    g02431(.A1(new_n3436_), .A2(new_n3418_), .A3(new_n3424_), .A4(new_n3427_), .ZN(new_n3437_));
  NOR3_X1    g02432(.A1(new_n3424_), .A2(new_n3427_), .A3(new_n3418_), .ZN(new_n3438_));
  INV_X1     g02433(.I(new_n3387_), .ZN(new_n3439_));
  NAND2_X1   g02434(.A1(new_n3429_), .A2(new_n3439_), .ZN(new_n3440_));
  NAND2_X1   g02435(.A1(new_n3410_), .A2(new_n3403_), .ZN(new_n3441_));
  NAND2_X1   g02436(.A1(new_n3441_), .A2(new_n3420_), .ZN(new_n3442_));
  OAI22_X1   g02437(.A1(new_n3364_), .A2(new_n3366_), .B1(new_n3371_), .B2(new_n3369_), .ZN(new_n3443_));
  NAND2_X1   g02438(.A1(new_n3443_), .A2(new_n3359_), .ZN(new_n3444_));
  NAND3_X1   g02439(.A1(new_n3372_), .A2(new_n3339_), .A3(new_n3344_), .ZN(new_n3445_));
  NOR4_X1    g02440(.A1(new_n3442_), .A2(new_n3445_), .A3(new_n3444_), .A4(new_n3440_), .ZN(new_n3446_));
  NOR2_X1    g02441(.A1(new_n3438_), .A2(new_n3446_), .ZN(new_n3447_));
  OAI21_X1   g02442(.A1(new_n3447_), .A2(new_n3437_), .B(new_n3378_), .ZN(new_n3448_));
  OAI21_X1   g02443(.A1(new_n3425_), .A2(new_n3426_), .B(new_n3382_), .ZN(new_n3449_));
  NAND3_X1   g02444(.A1(new_n3421_), .A2(new_n3423_), .A3(new_n3419_), .ZN(new_n3450_));
  NAND2_X1   g02445(.A1(new_n3450_), .A2(new_n3449_), .ZN(new_n3451_));
  OAI21_X1   g02446(.A1(new_n3451_), .A2(new_n3418_), .B(new_n3446_), .ZN(new_n3452_));
  NAND3_X1   g02447(.A1(new_n3433_), .A2(new_n3431_), .A3(new_n3428_), .ZN(new_n3453_));
  NOR2_X1    g02448(.A1(new_n3418_), .A2(new_n3445_), .ZN(new_n3454_));
  OAI21_X1   g02449(.A1(new_n3451_), .A2(new_n3453_), .B(new_n3454_), .ZN(new_n3455_));
  NAND3_X1   g02450(.A1(new_n3455_), .A2(new_n3452_), .A3(new_n3378_), .ZN(new_n3456_));
  NAND2_X1   g02451(.A1(new_n3456_), .A2(new_n3448_), .ZN(new_n3457_));
  OR2_X2     g02452(.A1(new_n3374_), .A2(new_n3377_), .Z(new_n3458_));
  NAND2_X1   g02453(.A1(new_n3438_), .A2(new_n3446_), .ZN(new_n3459_));
  OAI21_X1   g02454(.A1(new_n3451_), .A2(new_n3418_), .B(new_n3436_), .ZN(new_n3460_));
  AOI21_X1   g02455(.A1(new_n3460_), .A2(new_n3459_), .B(new_n3458_), .ZN(new_n3461_));
  NOR2_X1    g02456(.A1(new_n3438_), .A2(new_n3436_), .ZN(new_n3462_));
  NOR2_X1    g02457(.A1(new_n3424_), .A2(new_n3427_), .ZN(new_n3463_));
  NOR3_X1    g02458(.A1(new_n3442_), .A2(new_n3444_), .A3(new_n3440_), .ZN(new_n3464_));
  NOR2_X1    g02459(.A1(new_n3416_), .A2(new_n3410_), .ZN(new_n3465_));
  NOR2_X1    g02460(.A1(new_n3395_), .A2(new_n3403_), .ZN(new_n3466_));
  OAI21_X1   g02461(.A1(new_n3465_), .A2(new_n3466_), .B(new_n3439_), .ZN(new_n3467_));
  NAND2_X1   g02462(.A1(new_n3467_), .A2(new_n3435_), .ZN(new_n3468_));
  AOI21_X1   g02463(.A1(new_n3463_), .A2(new_n3464_), .B(new_n3468_), .ZN(new_n3469_));
  NOR3_X1    g02464(.A1(new_n3469_), .A2(new_n3462_), .A3(new_n3458_), .ZN(new_n3470_));
  NOR2_X1    g02465(.A1(new_n3442_), .A2(new_n3440_), .ZN(new_n3471_));
  NAND2_X1   g02466(.A1(new_n3433_), .A2(new_n3435_), .ZN(new_n3472_));
  NOR2_X1    g02467(.A1(new_n3471_), .A2(new_n3472_), .ZN(new_n3473_));
  NAND2_X1   g02468(.A1(new_n3431_), .A2(new_n3428_), .ZN(new_n3474_));
  NOR2_X1    g02469(.A1(new_n3445_), .A2(new_n3444_), .ZN(new_n3475_));
  NOR2_X1    g02470(.A1(new_n3475_), .A2(new_n3474_), .ZN(new_n3476_));
  INV_X1     g02471(.I(\A[375] ), .ZN(new_n3477_));
  NOR2_X1    g02472(.A1(new_n3477_), .A2(\A[374] ), .ZN(new_n3478_));
  INV_X1     g02473(.I(\A[374] ), .ZN(new_n3479_));
  NOR2_X1    g02474(.A1(new_n3479_), .A2(\A[375] ), .ZN(new_n3480_));
  OAI21_X1   g02475(.A1(new_n3478_), .A2(new_n3480_), .B(\A[373] ), .ZN(new_n3481_));
  INV_X1     g02476(.I(\A[373] ), .ZN(new_n3482_));
  NOR2_X1    g02477(.A1(\A[374] ), .A2(\A[375] ), .ZN(new_n3483_));
  NAND2_X1   g02478(.A1(\A[374] ), .A2(\A[375] ), .ZN(new_n3484_));
  INV_X1     g02479(.I(new_n3484_), .ZN(new_n3485_));
  OAI21_X1   g02480(.A1(new_n3485_), .A2(new_n3483_), .B(new_n3482_), .ZN(new_n3486_));
  NAND2_X1   g02481(.A1(new_n3481_), .A2(new_n3486_), .ZN(new_n3487_));
  INV_X1     g02482(.I(\A[378] ), .ZN(new_n3488_));
  NOR2_X1    g02483(.A1(new_n3488_), .A2(\A[377] ), .ZN(new_n3489_));
  INV_X1     g02484(.I(\A[377] ), .ZN(new_n3490_));
  NOR2_X1    g02485(.A1(new_n3490_), .A2(\A[378] ), .ZN(new_n3491_));
  OAI21_X1   g02486(.A1(new_n3489_), .A2(new_n3491_), .B(\A[376] ), .ZN(new_n3492_));
  INV_X1     g02487(.I(\A[376] ), .ZN(new_n3493_));
  NOR2_X1    g02488(.A1(\A[377] ), .A2(\A[378] ), .ZN(new_n3494_));
  AND2_X2    g02489(.A1(\A[377] ), .A2(\A[378] ), .Z(new_n3495_));
  OAI21_X1   g02490(.A1(new_n3495_), .A2(new_n3494_), .B(new_n3493_), .ZN(new_n3496_));
  NAND2_X1   g02491(.A1(new_n3492_), .A2(new_n3496_), .ZN(new_n3497_));
  NAND2_X1   g02492(.A1(\A[377] ), .A2(\A[378] ), .ZN(new_n3498_));
  AOI21_X1   g02493(.A1(new_n3493_), .A2(new_n3498_), .B(new_n3494_), .ZN(new_n3499_));
  AOI21_X1   g02494(.A1(new_n3482_), .A2(new_n3484_), .B(new_n3483_), .ZN(new_n3500_));
  NAND2_X1   g02495(.A1(new_n3499_), .A2(new_n3500_), .ZN(new_n3501_));
  NOR3_X1    g02496(.A1(new_n3487_), .A2(new_n3497_), .A3(new_n3501_), .ZN(new_n3502_));
  NOR2_X1    g02497(.A1(new_n3487_), .A2(new_n3497_), .ZN(new_n3503_));
  NAND2_X1   g02498(.A1(new_n3479_), .A2(\A[375] ), .ZN(new_n3504_));
  NAND2_X1   g02499(.A1(new_n3477_), .A2(\A[374] ), .ZN(new_n3505_));
  AOI21_X1   g02500(.A1(new_n3504_), .A2(new_n3505_), .B(new_n3482_), .ZN(new_n3506_));
  INV_X1     g02501(.I(new_n3483_), .ZN(new_n3507_));
  AOI21_X1   g02502(.A1(new_n3507_), .A2(new_n3484_), .B(\A[373] ), .ZN(new_n3508_));
  NOR2_X1    g02503(.A1(new_n3508_), .A2(new_n3506_), .ZN(new_n3509_));
  NAND2_X1   g02504(.A1(new_n3490_), .A2(\A[378] ), .ZN(new_n3510_));
  NAND2_X1   g02505(.A1(new_n3488_), .A2(\A[377] ), .ZN(new_n3511_));
  AOI21_X1   g02506(.A1(new_n3510_), .A2(new_n3511_), .B(new_n3493_), .ZN(new_n3512_));
  INV_X1     g02507(.I(new_n3494_), .ZN(new_n3513_));
  AOI21_X1   g02508(.A1(new_n3513_), .A2(new_n3498_), .B(\A[376] ), .ZN(new_n3514_));
  NOR2_X1    g02509(.A1(new_n3514_), .A2(new_n3512_), .ZN(new_n3515_));
  NOR2_X1    g02510(.A1(new_n3509_), .A2(new_n3515_), .ZN(new_n3516_));
  NOR2_X1    g02511(.A1(new_n3516_), .A2(new_n3503_), .ZN(new_n3517_));
  INV_X1     g02512(.I(\A[367] ), .ZN(new_n3518_));
  INV_X1     g02513(.I(\A[368] ), .ZN(new_n3519_));
  NAND2_X1   g02514(.A1(new_n3519_), .A2(\A[369] ), .ZN(new_n3520_));
  INV_X1     g02515(.I(\A[369] ), .ZN(new_n3521_));
  NAND2_X1   g02516(.A1(new_n3521_), .A2(\A[368] ), .ZN(new_n3522_));
  AOI21_X1   g02517(.A1(new_n3520_), .A2(new_n3522_), .B(new_n3518_), .ZN(new_n3523_));
  NOR2_X1    g02518(.A1(\A[368] ), .A2(\A[369] ), .ZN(new_n3524_));
  INV_X1     g02519(.I(new_n3524_), .ZN(new_n3525_));
  NAND2_X1   g02520(.A1(\A[368] ), .A2(\A[369] ), .ZN(new_n3526_));
  AOI21_X1   g02521(.A1(new_n3525_), .A2(new_n3526_), .B(\A[367] ), .ZN(new_n3527_));
  NOR2_X1    g02522(.A1(new_n3527_), .A2(new_n3523_), .ZN(new_n3528_));
  INV_X1     g02523(.I(\A[370] ), .ZN(new_n3529_));
  INV_X1     g02524(.I(\A[371] ), .ZN(new_n3530_));
  NAND2_X1   g02525(.A1(new_n3530_), .A2(\A[372] ), .ZN(new_n3531_));
  INV_X1     g02526(.I(\A[372] ), .ZN(new_n3532_));
  NAND2_X1   g02527(.A1(new_n3532_), .A2(\A[371] ), .ZN(new_n3533_));
  AOI21_X1   g02528(.A1(new_n3531_), .A2(new_n3533_), .B(new_n3529_), .ZN(new_n3534_));
  NOR2_X1    g02529(.A1(\A[371] ), .A2(\A[372] ), .ZN(new_n3535_));
  INV_X1     g02530(.I(new_n3535_), .ZN(new_n3536_));
  NAND2_X1   g02531(.A1(\A[371] ), .A2(\A[372] ), .ZN(new_n3537_));
  AOI21_X1   g02532(.A1(new_n3536_), .A2(new_n3537_), .B(\A[370] ), .ZN(new_n3538_));
  NOR2_X1    g02533(.A1(new_n3538_), .A2(new_n3534_), .ZN(new_n3539_));
  AOI21_X1   g02534(.A1(new_n3529_), .A2(new_n3537_), .B(new_n3535_), .ZN(new_n3540_));
  AOI21_X1   g02535(.A1(new_n3518_), .A2(new_n3526_), .B(new_n3524_), .ZN(new_n3541_));
  NAND2_X1   g02536(.A1(new_n3540_), .A2(new_n3541_), .ZN(new_n3542_));
  AND2_X2    g02537(.A1(new_n3517_), .A2(new_n3502_), .Z(new_n3544_));
  OR3_X2     g02538(.A1(new_n3473_), .A2(new_n3476_), .A3(new_n3544_), .Z(new_n3545_));
  OAI21_X1   g02539(.A1(new_n3461_), .A2(new_n3470_), .B(new_n3545_), .ZN(new_n3546_));
  NAND2_X1   g02540(.A1(new_n3475_), .A2(new_n3474_), .ZN(new_n3547_));
  NAND2_X1   g02541(.A1(new_n3471_), .A2(new_n3472_), .ZN(new_n3548_));
  NAND2_X1   g02542(.A1(new_n3548_), .A2(new_n3547_), .ZN(new_n3549_));
  NOR2_X1    g02543(.A1(new_n3549_), .A2(new_n3544_), .ZN(new_n3550_));
  NAND3_X1   g02544(.A1(new_n3456_), .A2(new_n3448_), .A3(new_n3550_), .ZN(new_n3551_));
  NAND2_X1   g02545(.A1(new_n3509_), .A2(new_n3515_), .ZN(new_n3552_));
  NAND2_X1   g02546(.A1(new_n3487_), .A2(new_n3497_), .ZN(new_n3553_));
  NAND3_X1   g02547(.A1(new_n3502_), .A2(new_n3552_), .A3(new_n3553_), .ZN(new_n3554_));
  NAND2_X1   g02548(.A1(new_n3528_), .A2(new_n3539_), .ZN(new_n3555_));
  NOR2_X1    g02549(.A1(new_n3521_), .A2(\A[368] ), .ZN(new_n3556_));
  NOR2_X1    g02550(.A1(new_n3519_), .A2(\A[369] ), .ZN(new_n3557_));
  OAI21_X1   g02551(.A1(new_n3556_), .A2(new_n3557_), .B(\A[367] ), .ZN(new_n3558_));
  INV_X1     g02552(.I(new_n3526_), .ZN(new_n3559_));
  OAI21_X1   g02553(.A1(new_n3559_), .A2(new_n3524_), .B(new_n3518_), .ZN(new_n3560_));
  NAND2_X1   g02554(.A1(new_n3558_), .A2(new_n3560_), .ZN(new_n3561_));
  NOR2_X1    g02555(.A1(new_n3532_), .A2(\A[371] ), .ZN(new_n3562_));
  NOR2_X1    g02556(.A1(new_n3530_), .A2(\A[372] ), .ZN(new_n3563_));
  OAI21_X1   g02557(.A1(new_n3562_), .A2(new_n3563_), .B(\A[370] ), .ZN(new_n3564_));
  INV_X1     g02558(.I(new_n3537_), .ZN(new_n3565_));
  OAI21_X1   g02559(.A1(new_n3565_), .A2(new_n3535_), .B(new_n3529_), .ZN(new_n3566_));
  NAND2_X1   g02560(.A1(new_n3564_), .A2(new_n3566_), .ZN(new_n3567_));
  NAND2_X1   g02561(.A1(new_n3561_), .A2(new_n3567_), .ZN(new_n3568_));
  NAND2_X1   g02562(.A1(new_n3555_), .A2(new_n3568_), .ZN(new_n3569_));
  INV_X1     g02563(.I(new_n3499_), .ZN(new_n3570_));
  OAI21_X1   g02564(.A1(new_n3487_), .A2(new_n3497_), .B(new_n3500_), .ZN(new_n3571_));
  INV_X1     g02565(.I(new_n3500_), .ZN(new_n3572_));
  NAND3_X1   g02566(.A1(new_n3509_), .A2(new_n3515_), .A3(new_n3572_), .ZN(new_n3573_));
  AOI21_X1   g02567(.A1(new_n3573_), .A2(new_n3571_), .B(new_n3570_), .ZN(new_n3574_));
  AOI21_X1   g02568(.A1(new_n3509_), .A2(new_n3515_), .B(new_n3572_), .ZN(new_n3575_));
  NOR3_X1    g02569(.A1(new_n3487_), .A2(new_n3497_), .A3(new_n3500_), .ZN(new_n3576_));
  NOR3_X1    g02570(.A1(new_n3575_), .A2(new_n3576_), .A3(new_n3499_), .ZN(new_n3577_));
  NOR4_X1    g02571(.A1(new_n3574_), .A2(new_n3577_), .A3(new_n3554_), .A4(new_n3569_), .ZN(new_n3578_));
  NOR3_X1    g02572(.A1(new_n3561_), .A2(new_n3567_), .A3(new_n3542_), .ZN(new_n3579_));
  INV_X1     g02573(.I(new_n3501_), .ZN(new_n3580_));
  NOR2_X1    g02574(.A1(new_n3515_), .A2(new_n3487_), .ZN(new_n3581_));
  NOR2_X1    g02575(.A1(new_n3509_), .A2(new_n3497_), .ZN(new_n3582_));
  OAI21_X1   g02576(.A1(new_n3581_), .A2(new_n3582_), .B(new_n3580_), .ZN(new_n3583_));
  NAND2_X1   g02577(.A1(new_n3583_), .A2(new_n3579_), .ZN(new_n3584_));
  INV_X1     g02578(.I(new_n3540_), .ZN(new_n3585_));
  OAI21_X1   g02579(.A1(new_n3561_), .A2(new_n3567_), .B(new_n3541_), .ZN(new_n3586_));
  INV_X1     g02580(.I(new_n3541_), .ZN(new_n3587_));
  NAND3_X1   g02581(.A1(new_n3528_), .A2(new_n3539_), .A3(new_n3587_), .ZN(new_n3588_));
  AOI21_X1   g02582(.A1(new_n3586_), .A2(new_n3588_), .B(new_n3585_), .ZN(new_n3589_));
  AOI21_X1   g02583(.A1(new_n3528_), .A2(new_n3539_), .B(new_n3587_), .ZN(new_n3590_));
  NOR3_X1    g02584(.A1(new_n3561_), .A2(new_n3567_), .A3(new_n3541_), .ZN(new_n3591_));
  NOR3_X1    g02585(.A1(new_n3590_), .A2(new_n3591_), .A3(new_n3540_), .ZN(new_n3592_));
  NOR2_X1    g02586(.A1(new_n3592_), .A2(new_n3589_), .ZN(new_n3593_));
  NOR3_X1    g02587(.A1(new_n3578_), .A2(new_n3593_), .A3(new_n3584_), .ZN(new_n3594_));
  INV_X1     g02588(.I(new_n3594_), .ZN(new_n3595_));
  OAI21_X1   g02589(.A1(new_n3590_), .A2(new_n3591_), .B(new_n3540_), .ZN(new_n3596_));
  NAND3_X1   g02590(.A1(new_n3586_), .A2(new_n3588_), .A3(new_n3585_), .ZN(new_n3597_));
  NAND2_X1   g02591(.A1(new_n3596_), .A2(new_n3597_), .ZN(new_n3598_));
  NOR4_X1    g02592(.A1(new_n3523_), .A2(new_n3527_), .A3(new_n3538_), .A4(new_n3534_), .ZN(new_n3599_));
  NOR2_X1    g02593(.A1(new_n3528_), .A2(new_n3539_), .ZN(new_n3600_));
  NOR2_X1    g02594(.A1(new_n3600_), .A2(new_n3599_), .ZN(new_n3601_));
  NAND4_X1   g02595(.A1(new_n3517_), .A2(new_n3601_), .A3(new_n3502_), .A4(new_n3579_), .ZN(new_n3602_));
  NAND2_X1   g02596(.A1(new_n3598_), .A2(new_n3602_), .ZN(new_n3603_));
  NAND2_X1   g02597(.A1(new_n3509_), .A2(new_n3497_), .ZN(new_n3604_));
  NAND2_X1   g02598(.A1(new_n3515_), .A2(new_n3487_), .ZN(new_n3605_));
  AOI21_X1   g02599(.A1(new_n3605_), .A2(new_n3604_), .B(new_n3501_), .ZN(new_n3606_));
  NOR3_X1    g02600(.A1(new_n3577_), .A2(new_n3574_), .A3(new_n3606_), .ZN(new_n3607_));
  NAND3_X1   g02601(.A1(new_n3579_), .A2(new_n3555_), .A3(new_n3568_), .ZN(new_n3608_));
  NOR4_X1    g02602(.A1(new_n3589_), .A2(new_n3592_), .A3(new_n3608_), .A4(new_n3554_), .ZN(new_n3609_));
  NOR2_X1    g02603(.A1(new_n3609_), .A2(new_n3607_), .ZN(new_n3610_));
  OAI21_X1   g02604(.A1(new_n3575_), .A2(new_n3576_), .B(new_n3499_), .ZN(new_n3611_));
  NAND3_X1   g02605(.A1(new_n3573_), .A2(new_n3571_), .A3(new_n3570_), .ZN(new_n3612_));
  NAND3_X1   g02606(.A1(new_n3611_), .A2(new_n3612_), .A3(new_n3583_), .ZN(new_n3613_));
  NOR3_X1    g02607(.A1(new_n3613_), .A2(new_n3598_), .A3(new_n3602_), .ZN(new_n3614_));
  OAI21_X1   g02608(.A1(new_n3610_), .A2(new_n3614_), .B(new_n3603_), .ZN(new_n3615_));
  NAND2_X1   g02609(.A1(new_n3615_), .A2(new_n3595_), .ZN(new_n3616_));
  AOI22_X1   g02610(.A1(new_n3546_), .A2(new_n3551_), .B1(new_n3616_), .B2(new_n3457_), .ZN(new_n3617_));
  NOR2_X1    g02611(.A1(new_n3462_), .A2(new_n3378_), .ZN(new_n3618_));
  NAND2_X1   g02612(.A1(new_n3422_), .A2(new_n3419_), .ZN(new_n3619_));
  AOI21_X1   g02613(.A1(new_n3429_), .A2(new_n3619_), .B(new_n3439_), .ZN(new_n3620_));
  NOR2_X1    g02614(.A1(new_n3339_), .A2(new_n3344_), .ZN(new_n3621_));
  OAI21_X1   g02615(.A1(new_n3359_), .A2(new_n3621_), .B(new_n3434_), .ZN(new_n3622_));
  XOR2_X1    g02616(.A1(new_n3620_), .A2(new_n3622_), .Z(new_n3623_));
  INV_X1     g02617(.I(new_n3623_), .ZN(new_n3624_));
  NOR3_X1    g02618(.A1(new_n3618_), .A2(new_n3624_), .A3(new_n3469_), .ZN(new_n3625_));
  NOR2_X1    g02619(.A1(new_n3578_), .A2(new_n3584_), .ZN(new_n3626_));
  INV_X1     g02620(.I(new_n3602_), .ZN(new_n3627_));
  AOI21_X1   g02621(.A1(new_n3627_), .A2(new_n3613_), .B(new_n3593_), .ZN(new_n3628_));
  NAND2_X1   g02622(.A1(new_n3572_), .A2(new_n3570_), .ZN(new_n3629_));
  AOI21_X1   g02623(.A1(new_n3503_), .A2(new_n3629_), .B(new_n3580_), .ZN(new_n3630_));
  NOR2_X1    g02624(.A1(new_n3540_), .A2(new_n3541_), .ZN(new_n3631_));
  OAI21_X1   g02625(.A1(new_n3555_), .A2(new_n3631_), .B(new_n3542_), .ZN(new_n3632_));
  XNOR2_X1   g02626(.A1(new_n3632_), .A2(new_n3630_), .ZN(new_n3633_));
  NOR3_X1    g02627(.A1(new_n3628_), .A2(new_n3626_), .A3(new_n3633_), .ZN(new_n3634_));
  XOR2_X1    g02628(.A1(new_n3625_), .A2(new_n3634_), .Z(new_n3635_));
  NAND2_X1   g02629(.A1(new_n3635_), .A2(new_n3617_), .ZN(new_n3636_));
  NOR2_X1    g02630(.A1(new_n3461_), .A2(new_n3470_), .ZN(new_n3637_));
  AOI21_X1   g02631(.A1(new_n3456_), .A2(new_n3448_), .B(new_n3550_), .ZN(new_n3638_));
  NOR3_X1    g02632(.A1(new_n3461_), .A2(new_n3470_), .A3(new_n3545_), .ZN(new_n3639_));
  OAI21_X1   g02633(.A1(new_n3598_), .A2(new_n3602_), .B(new_n3613_), .ZN(new_n3640_));
  NAND2_X1   g02634(.A1(new_n3609_), .A2(new_n3607_), .ZN(new_n3641_));
  NAND2_X1   g02635(.A1(new_n3640_), .A2(new_n3641_), .ZN(new_n3642_));
  AOI21_X1   g02636(.A1(new_n3642_), .A2(new_n3603_), .B(new_n3594_), .ZN(new_n3643_));
  OAI22_X1   g02637(.A1(new_n3638_), .A2(new_n3639_), .B1(new_n3643_), .B2(new_n3637_), .ZN(new_n3644_));
  NAND2_X1   g02638(.A1(new_n3452_), .A2(new_n3458_), .ZN(new_n3645_));
  NAND3_X1   g02639(.A1(new_n3645_), .A2(new_n3455_), .A3(new_n3623_), .ZN(new_n3646_));
  OR3_X2     g02640(.A1(new_n3628_), .A2(new_n3626_), .A3(new_n3633_), .Z(new_n3647_));
  NAND2_X1   g02641(.A1(new_n3647_), .A2(new_n3646_), .ZN(new_n3648_));
  NAND2_X1   g02642(.A1(new_n3625_), .A2(new_n3634_), .ZN(new_n3649_));
  NAND2_X1   g02643(.A1(new_n3648_), .A2(new_n3649_), .ZN(new_n3650_));
  NAND2_X1   g02644(.A1(new_n3650_), .A2(new_n3644_), .ZN(new_n3651_));
  NAND2_X1   g02645(.A1(new_n3636_), .A2(new_n3651_), .ZN(new_n3652_));
  INV_X1     g02646(.I(\A[412] ), .ZN(new_n3653_));
  NOR2_X1    g02647(.A1(\A[413] ), .A2(\A[414] ), .ZN(new_n3654_));
  NAND2_X1   g02648(.A1(\A[413] ), .A2(\A[414] ), .ZN(new_n3655_));
  AOI21_X1   g02649(.A1(new_n3653_), .A2(new_n3655_), .B(new_n3654_), .ZN(new_n3656_));
  INV_X1     g02650(.I(new_n3656_), .ZN(new_n3657_));
  INV_X1     g02651(.I(\A[409] ), .ZN(new_n3658_));
  NOR2_X1    g02652(.A1(\A[410] ), .A2(\A[411] ), .ZN(new_n3659_));
  NAND2_X1   g02653(.A1(\A[410] ), .A2(\A[411] ), .ZN(new_n3660_));
  AOI21_X1   g02654(.A1(new_n3658_), .A2(new_n3660_), .B(new_n3659_), .ZN(new_n3661_));
  INV_X1     g02655(.I(\A[411] ), .ZN(new_n3662_));
  NOR2_X1    g02656(.A1(new_n3662_), .A2(\A[410] ), .ZN(new_n3663_));
  INV_X1     g02657(.I(\A[410] ), .ZN(new_n3664_));
  NOR2_X1    g02658(.A1(new_n3664_), .A2(\A[411] ), .ZN(new_n3665_));
  OAI21_X1   g02659(.A1(new_n3663_), .A2(new_n3665_), .B(\A[409] ), .ZN(new_n3666_));
  INV_X1     g02660(.I(new_n3660_), .ZN(new_n3667_));
  OAI21_X1   g02661(.A1(new_n3667_), .A2(new_n3659_), .B(new_n3658_), .ZN(new_n3668_));
  INV_X1     g02662(.I(\A[414] ), .ZN(new_n3669_));
  NOR2_X1    g02663(.A1(new_n3669_), .A2(\A[413] ), .ZN(new_n3670_));
  INV_X1     g02664(.I(\A[413] ), .ZN(new_n3671_));
  NOR2_X1    g02665(.A1(new_n3671_), .A2(\A[414] ), .ZN(new_n3672_));
  OAI21_X1   g02666(.A1(new_n3670_), .A2(new_n3672_), .B(\A[412] ), .ZN(new_n3673_));
  INV_X1     g02667(.I(new_n3655_), .ZN(new_n3674_));
  OAI21_X1   g02668(.A1(new_n3674_), .A2(new_n3654_), .B(new_n3653_), .ZN(new_n3675_));
  NAND4_X1   g02669(.A1(new_n3666_), .A2(new_n3668_), .A3(new_n3673_), .A4(new_n3675_), .ZN(new_n3676_));
  NAND2_X1   g02670(.A1(new_n3676_), .A2(new_n3661_), .ZN(new_n3677_));
  INV_X1     g02671(.I(new_n3661_), .ZN(new_n3678_));
  NAND2_X1   g02672(.A1(new_n3671_), .A2(\A[414] ), .ZN(new_n3679_));
  NAND2_X1   g02673(.A1(new_n3669_), .A2(\A[413] ), .ZN(new_n3680_));
  AOI21_X1   g02674(.A1(new_n3679_), .A2(new_n3680_), .B(new_n3653_), .ZN(new_n3681_));
  INV_X1     g02675(.I(new_n3654_), .ZN(new_n3682_));
  AOI21_X1   g02676(.A1(new_n3682_), .A2(new_n3655_), .B(\A[412] ), .ZN(new_n3683_));
  NOR2_X1    g02677(.A1(new_n3683_), .A2(new_n3681_), .ZN(new_n3684_));
  NAND4_X1   g02678(.A1(new_n3684_), .A2(new_n3678_), .A3(new_n3666_), .A4(new_n3668_), .ZN(new_n3685_));
  AOI21_X1   g02679(.A1(new_n3677_), .A2(new_n3685_), .B(new_n3657_), .ZN(new_n3686_));
  NAND2_X1   g02680(.A1(new_n3664_), .A2(\A[411] ), .ZN(new_n3687_));
  NAND2_X1   g02681(.A1(new_n3662_), .A2(\A[410] ), .ZN(new_n3688_));
  AOI21_X1   g02682(.A1(new_n3687_), .A2(new_n3688_), .B(new_n3658_), .ZN(new_n3689_));
  INV_X1     g02683(.I(new_n3659_), .ZN(new_n3690_));
  AOI21_X1   g02684(.A1(new_n3690_), .A2(new_n3660_), .B(\A[409] ), .ZN(new_n3691_));
  NOR4_X1    g02685(.A1(new_n3689_), .A2(new_n3691_), .A3(new_n3683_), .A4(new_n3681_), .ZN(new_n3692_));
  NOR2_X1    g02686(.A1(new_n3692_), .A2(new_n3678_), .ZN(new_n3693_));
  NOR2_X1    g02687(.A1(new_n3676_), .A2(new_n3661_), .ZN(new_n3694_));
  NOR3_X1    g02688(.A1(new_n3693_), .A2(new_n3694_), .A3(new_n3656_), .ZN(new_n3695_));
  INV_X1     g02689(.I(\A[405] ), .ZN(new_n3696_));
  NOR2_X1    g02690(.A1(new_n3696_), .A2(\A[404] ), .ZN(new_n3697_));
  INV_X1     g02691(.I(\A[404] ), .ZN(new_n3698_));
  NOR2_X1    g02692(.A1(new_n3698_), .A2(\A[405] ), .ZN(new_n3699_));
  OAI21_X1   g02693(.A1(new_n3697_), .A2(new_n3699_), .B(\A[403] ), .ZN(new_n3700_));
  INV_X1     g02694(.I(\A[403] ), .ZN(new_n3701_));
  NOR2_X1    g02695(.A1(\A[404] ), .A2(\A[405] ), .ZN(new_n3702_));
  NAND2_X1   g02696(.A1(\A[404] ), .A2(\A[405] ), .ZN(new_n3703_));
  INV_X1     g02697(.I(new_n3703_), .ZN(new_n3704_));
  OAI21_X1   g02698(.A1(new_n3704_), .A2(new_n3702_), .B(new_n3701_), .ZN(new_n3705_));
  INV_X1     g02699(.I(\A[408] ), .ZN(new_n3706_));
  NOR2_X1    g02700(.A1(new_n3706_), .A2(\A[407] ), .ZN(new_n3707_));
  INV_X1     g02701(.I(\A[407] ), .ZN(new_n3708_));
  NOR2_X1    g02702(.A1(new_n3708_), .A2(\A[408] ), .ZN(new_n3709_));
  OAI21_X1   g02703(.A1(new_n3707_), .A2(new_n3709_), .B(\A[406] ), .ZN(new_n3710_));
  INV_X1     g02704(.I(\A[406] ), .ZN(new_n3711_));
  NOR2_X1    g02705(.A1(\A[407] ), .A2(\A[408] ), .ZN(new_n3712_));
  NAND2_X1   g02706(.A1(\A[407] ), .A2(\A[408] ), .ZN(new_n3713_));
  INV_X1     g02707(.I(new_n3713_), .ZN(new_n3714_));
  OAI21_X1   g02708(.A1(new_n3714_), .A2(new_n3712_), .B(new_n3711_), .ZN(new_n3715_));
  NAND4_X1   g02709(.A1(new_n3700_), .A2(new_n3705_), .A3(new_n3710_), .A4(new_n3715_), .ZN(new_n3716_));
  NAND2_X1   g02710(.A1(new_n3698_), .A2(\A[405] ), .ZN(new_n3717_));
  NAND2_X1   g02711(.A1(new_n3696_), .A2(\A[404] ), .ZN(new_n3718_));
  AOI21_X1   g02712(.A1(new_n3717_), .A2(new_n3718_), .B(new_n3701_), .ZN(new_n3719_));
  INV_X1     g02713(.I(new_n3702_), .ZN(new_n3720_));
  AOI21_X1   g02714(.A1(new_n3720_), .A2(new_n3703_), .B(\A[403] ), .ZN(new_n3721_));
  NAND2_X1   g02715(.A1(new_n3708_), .A2(\A[408] ), .ZN(new_n3722_));
  NAND2_X1   g02716(.A1(new_n3706_), .A2(\A[407] ), .ZN(new_n3723_));
  AOI21_X1   g02717(.A1(new_n3722_), .A2(new_n3723_), .B(new_n3711_), .ZN(new_n3724_));
  INV_X1     g02718(.I(new_n3712_), .ZN(new_n3725_));
  AOI21_X1   g02719(.A1(new_n3725_), .A2(new_n3713_), .B(\A[406] ), .ZN(new_n3726_));
  OAI22_X1   g02720(.A1(new_n3719_), .A2(new_n3721_), .B1(new_n3726_), .B2(new_n3724_), .ZN(new_n3727_));
  NAND2_X1   g02721(.A1(new_n3727_), .A2(new_n3716_), .ZN(new_n3728_));
  OAI22_X1   g02722(.A1(new_n3689_), .A2(new_n3691_), .B1(new_n3683_), .B2(new_n3681_), .ZN(new_n3729_));
  NAND2_X1   g02723(.A1(new_n3729_), .A2(new_n3676_), .ZN(new_n3730_));
  NAND2_X1   g02724(.A1(new_n3656_), .A2(new_n3661_), .ZN(new_n3731_));
  NOR2_X1    g02725(.A1(new_n3676_), .A2(new_n3731_), .ZN(new_n3732_));
  NOR2_X1    g02726(.A1(new_n3721_), .A2(new_n3719_), .ZN(new_n3733_));
  NOR2_X1    g02727(.A1(new_n3726_), .A2(new_n3724_), .ZN(new_n3734_));
  AOI21_X1   g02728(.A1(new_n3711_), .A2(new_n3713_), .B(new_n3712_), .ZN(new_n3735_));
  AOI21_X1   g02729(.A1(new_n3701_), .A2(new_n3703_), .B(new_n3702_), .ZN(new_n3736_));
  NAND4_X1   g02730(.A1(new_n3733_), .A2(new_n3734_), .A3(new_n3735_), .A4(new_n3736_), .ZN(new_n3737_));
  NOR4_X1    g02731(.A1(new_n3728_), .A2(new_n3730_), .A3(new_n3732_), .A4(new_n3737_), .ZN(new_n3738_));
  NOR3_X1    g02732(.A1(new_n3738_), .A2(new_n3686_), .A3(new_n3695_), .ZN(new_n3739_));
  NOR4_X1    g02733(.A1(new_n3719_), .A2(new_n3721_), .A3(new_n3726_), .A4(new_n3724_), .ZN(new_n3740_));
  INV_X1     g02734(.I(new_n3736_), .ZN(new_n3741_));
  NOR2_X1    g02735(.A1(new_n3740_), .A2(new_n3741_), .ZN(new_n3742_));
  NOR2_X1    g02736(.A1(new_n3716_), .A2(new_n3736_), .ZN(new_n3743_));
  OAI21_X1   g02737(.A1(new_n3742_), .A2(new_n3743_), .B(new_n3735_), .ZN(new_n3744_));
  INV_X1     g02738(.I(new_n3735_), .ZN(new_n3745_));
  NAND2_X1   g02739(.A1(new_n3716_), .A2(new_n3736_), .ZN(new_n3746_));
  NAND2_X1   g02740(.A1(new_n3740_), .A2(new_n3741_), .ZN(new_n3747_));
  NAND3_X1   g02741(.A1(new_n3747_), .A2(new_n3746_), .A3(new_n3745_), .ZN(new_n3748_));
  NAND2_X1   g02742(.A1(new_n3744_), .A2(new_n3748_), .ZN(new_n3749_));
  NAND4_X1   g02743(.A1(new_n3676_), .A2(new_n3727_), .A3(new_n3729_), .A4(new_n3716_), .ZN(new_n3750_));
  NAND2_X1   g02744(.A1(new_n3735_), .A2(new_n3736_), .ZN(new_n3751_));
  NOR2_X1    g02745(.A1(new_n3716_), .A2(new_n3751_), .ZN(new_n3752_));
  INV_X1     g02746(.I(new_n3731_), .ZN(new_n3753_));
  NAND2_X1   g02747(.A1(new_n3729_), .A2(new_n3753_), .ZN(new_n3754_));
  NAND2_X1   g02748(.A1(new_n3754_), .A2(new_n3752_), .ZN(new_n3755_));
  XNOR2_X1   g02749(.A1(new_n3656_), .A2(new_n3661_), .ZN(new_n3756_));
  NOR2_X1    g02750(.A1(new_n3756_), .A2(new_n3676_), .ZN(new_n3757_));
  NAND2_X1   g02751(.A1(new_n3657_), .A2(new_n3678_), .ZN(new_n3758_));
  AOI21_X1   g02752(.A1(new_n3731_), .A2(new_n3758_), .B(new_n3692_), .ZN(new_n3759_));
  NOR4_X1    g02753(.A1(new_n3755_), .A2(new_n3750_), .A3(new_n3757_), .A4(new_n3759_), .ZN(new_n3760_));
  NOR3_X1    g02754(.A1(new_n3739_), .A2(new_n3749_), .A3(new_n3760_), .ZN(new_n3761_));
  NAND2_X1   g02755(.A1(new_n3692_), .A2(new_n3753_), .ZN(new_n3762_));
  NAND2_X1   g02756(.A1(new_n3762_), .A2(new_n3752_), .ZN(new_n3763_));
  OAI22_X1   g02757(.A1(new_n3695_), .A2(new_n3686_), .B1(new_n3763_), .B2(new_n3750_), .ZN(new_n3764_));
  OAI21_X1   g02758(.A1(new_n3693_), .A2(new_n3694_), .B(new_n3656_), .ZN(new_n3765_));
  NAND3_X1   g02759(.A1(new_n3677_), .A2(new_n3685_), .A3(new_n3657_), .ZN(new_n3766_));
  AOI22_X1   g02760(.A1(new_n3700_), .A2(new_n3705_), .B1(new_n3710_), .B2(new_n3715_), .ZN(new_n3767_));
  AOI22_X1   g02761(.A1(new_n3666_), .A2(new_n3668_), .B1(new_n3673_), .B2(new_n3675_), .ZN(new_n3768_));
  NOR4_X1    g02762(.A1(new_n3692_), .A2(new_n3767_), .A3(new_n3768_), .A4(new_n3740_), .ZN(new_n3769_));
  NOR2_X1    g02763(.A1(new_n3732_), .A2(new_n3737_), .ZN(new_n3770_));
  NAND4_X1   g02764(.A1(new_n3765_), .A2(new_n3766_), .A3(new_n3770_), .A4(new_n3769_), .ZN(new_n3771_));
  AOI21_X1   g02765(.A1(new_n3764_), .A2(new_n3771_), .B(new_n3749_), .ZN(new_n3772_));
  NOR2_X1    g02766(.A1(new_n3761_), .A2(new_n3772_), .ZN(new_n3773_));
  NOR2_X1    g02767(.A1(new_n3767_), .A2(new_n3740_), .ZN(new_n3774_));
  NOR2_X1    g02768(.A1(new_n3768_), .A2(new_n3692_), .ZN(new_n3775_));
  NAND4_X1   g02769(.A1(new_n3774_), .A2(new_n3775_), .A3(new_n3762_), .A4(new_n3752_), .ZN(new_n3776_));
  NAND3_X1   g02770(.A1(new_n3776_), .A2(new_n3765_), .A3(new_n3766_), .ZN(new_n3777_));
  AOI21_X1   g02771(.A1(new_n3747_), .A2(new_n3746_), .B(new_n3745_), .ZN(new_n3778_));
  NOR3_X1    g02772(.A1(new_n3742_), .A2(new_n3743_), .A3(new_n3735_), .ZN(new_n3779_));
  NOR2_X1    g02773(.A1(new_n3778_), .A2(new_n3779_), .ZN(new_n3780_));
  AOI21_X1   g02774(.A1(new_n3729_), .A2(new_n3753_), .B(new_n3737_), .ZN(new_n3781_));
  NOR2_X1    g02775(.A1(new_n3757_), .A2(new_n3759_), .ZN(new_n3782_));
  NAND3_X1   g02776(.A1(new_n3782_), .A2(new_n3781_), .A3(new_n3769_), .ZN(new_n3783_));
  NAND3_X1   g02777(.A1(new_n3777_), .A2(new_n3783_), .A3(new_n3780_), .ZN(new_n3784_));
  AOI22_X1   g02778(.A1(new_n3765_), .A2(new_n3766_), .B1(new_n3770_), .B2(new_n3769_), .ZN(new_n3785_));
  NOR3_X1    g02779(.A1(new_n3776_), .A2(new_n3686_), .A3(new_n3695_), .ZN(new_n3786_));
  OAI21_X1   g02780(.A1(new_n3786_), .A2(new_n3785_), .B(new_n3780_), .ZN(new_n3787_));
  NOR2_X1    g02781(.A1(new_n3768_), .A2(new_n3692_), .ZN(new_n3788_));
  INV_X1     g02782(.I(new_n3788_), .ZN(new_n3789_));
  NAND3_X1   g02783(.A1(new_n3789_), .A2(new_n3774_), .A3(new_n3752_), .ZN(new_n3790_));
  NAND2_X1   g02784(.A1(new_n3774_), .A2(new_n3752_), .ZN(new_n3791_));
  NAND2_X1   g02785(.A1(new_n3791_), .A2(new_n3788_), .ZN(new_n3792_));
  INV_X1     g02786(.I(\A[400] ), .ZN(new_n3793_));
  NOR2_X1    g02787(.A1(\A[401] ), .A2(\A[402] ), .ZN(new_n3794_));
  NAND2_X1   g02788(.A1(\A[401] ), .A2(\A[402] ), .ZN(new_n3795_));
  AOI21_X1   g02789(.A1(new_n3793_), .A2(new_n3795_), .B(new_n3794_), .ZN(new_n3796_));
  INV_X1     g02790(.I(\A[397] ), .ZN(new_n3797_));
  NOR2_X1    g02791(.A1(\A[398] ), .A2(\A[399] ), .ZN(new_n3798_));
  NAND2_X1   g02792(.A1(\A[398] ), .A2(\A[399] ), .ZN(new_n3799_));
  AOI21_X1   g02793(.A1(new_n3797_), .A2(new_n3799_), .B(new_n3798_), .ZN(new_n3800_));
  NAND2_X1   g02794(.A1(new_n3796_), .A2(new_n3800_), .ZN(new_n3801_));
  INV_X1     g02795(.I(new_n3801_), .ZN(new_n3802_));
  INV_X1     g02796(.I(\A[399] ), .ZN(new_n3803_));
  NOR2_X1    g02797(.A1(new_n3803_), .A2(\A[398] ), .ZN(new_n3804_));
  INV_X1     g02798(.I(\A[398] ), .ZN(new_n3805_));
  NOR2_X1    g02799(.A1(new_n3805_), .A2(\A[399] ), .ZN(new_n3806_));
  OAI21_X1   g02800(.A1(new_n3804_), .A2(new_n3806_), .B(\A[397] ), .ZN(new_n3807_));
  INV_X1     g02801(.I(new_n3799_), .ZN(new_n3808_));
  OAI21_X1   g02802(.A1(new_n3808_), .A2(new_n3798_), .B(new_n3797_), .ZN(new_n3809_));
  NAND2_X1   g02803(.A1(new_n3807_), .A2(new_n3809_), .ZN(new_n3810_));
  INV_X1     g02804(.I(\A[402] ), .ZN(new_n3811_));
  NOR2_X1    g02805(.A1(new_n3811_), .A2(\A[401] ), .ZN(new_n3812_));
  INV_X1     g02806(.I(\A[401] ), .ZN(new_n3813_));
  NOR2_X1    g02807(.A1(new_n3813_), .A2(\A[402] ), .ZN(new_n3814_));
  OAI21_X1   g02808(.A1(new_n3812_), .A2(new_n3814_), .B(\A[400] ), .ZN(new_n3815_));
  AND2_X2    g02809(.A1(\A[401] ), .A2(\A[402] ), .Z(new_n3816_));
  OAI21_X1   g02810(.A1(new_n3816_), .A2(new_n3794_), .B(new_n3793_), .ZN(new_n3817_));
  NAND2_X1   g02811(.A1(new_n3815_), .A2(new_n3817_), .ZN(new_n3818_));
  NOR2_X1    g02812(.A1(new_n3810_), .A2(new_n3818_), .ZN(new_n3819_));
  NAND2_X1   g02813(.A1(new_n3819_), .A2(new_n3802_), .ZN(new_n3820_));
  NAND2_X1   g02814(.A1(new_n3805_), .A2(\A[399] ), .ZN(new_n3821_));
  NAND2_X1   g02815(.A1(new_n3803_), .A2(\A[398] ), .ZN(new_n3822_));
  AOI21_X1   g02816(.A1(new_n3821_), .A2(new_n3822_), .B(new_n3797_), .ZN(new_n3823_));
  INV_X1     g02817(.I(new_n3798_), .ZN(new_n3824_));
  AOI21_X1   g02818(.A1(new_n3824_), .A2(new_n3799_), .B(\A[397] ), .ZN(new_n3825_));
  NOR2_X1    g02819(.A1(new_n3825_), .A2(new_n3823_), .ZN(new_n3826_));
  NAND2_X1   g02820(.A1(new_n3813_), .A2(\A[402] ), .ZN(new_n3827_));
  NAND2_X1   g02821(.A1(new_n3811_), .A2(\A[401] ), .ZN(new_n3828_));
  AOI21_X1   g02822(.A1(new_n3827_), .A2(new_n3828_), .B(new_n3793_), .ZN(new_n3829_));
  INV_X1     g02823(.I(new_n3794_), .ZN(new_n3830_));
  AOI21_X1   g02824(.A1(new_n3830_), .A2(new_n3795_), .B(\A[400] ), .ZN(new_n3831_));
  NOR2_X1    g02825(.A1(new_n3831_), .A2(new_n3829_), .ZN(new_n3832_));
  NOR2_X1    g02826(.A1(new_n3826_), .A2(new_n3832_), .ZN(new_n3833_));
  NOR2_X1    g02827(.A1(new_n3833_), .A2(new_n3819_), .ZN(new_n3834_));
  INV_X1     g02828(.I(\A[391] ), .ZN(new_n3835_));
  INV_X1     g02829(.I(\A[392] ), .ZN(new_n3836_));
  NAND2_X1   g02830(.A1(new_n3836_), .A2(\A[393] ), .ZN(new_n3837_));
  INV_X1     g02831(.I(\A[393] ), .ZN(new_n3838_));
  NAND2_X1   g02832(.A1(new_n3838_), .A2(\A[392] ), .ZN(new_n3839_));
  AOI21_X1   g02833(.A1(new_n3837_), .A2(new_n3839_), .B(new_n3835_), .ZN(new_n3840_));
  NOR2_X1    g02834(.A1(\A[392] ), .A2(\A[393] ), .ZN(new_n3841_));
  INV_X1     g02835(.I(new_n3841_), .ZN(new_n3842_));
  NAND2_X1   g02836(.A1(\A[392] ), .A2(\A[393] ), .ZN(new_n3843_));
  AOI21_X1   g02837(.A1(new_n3842_), .A2(new_n3843_), .B(\A[391] ), .ZN(new_n3844_));
  NOR2_X1    g02838(.A1(new_n3844_), .A2(new_n3840_), .ZN(new_n3845_));
  INV_X1     g02839(.I(\A[394] ), .ZN(new_n3846_));
  INV_X1     g02840(.I(\A[395] ), .ZN(new_n3847_));
  NAND2_X1   g02841(.A1(new_n3847_), .A2(\A[396] ), .ZN(new_n3848_));
  INV_X1     g02842(.I(\A[396] ), .ZN(new_n3849_));
  NAND2_X1   g02843(.A1(new_n3849_), .A2(\A[395] ), .ZN(new_n3850_));
  AOI21_X1   g02844(.A1(new_n3848_), .A2(new_n3850_), .B(new_n3846_), .ZN(new_n3851_));
  NOR2_X1    g02845(.A1(\A[395] ), .A2(\A[396] ), .ZN(new_n3852_));
  INV_X1     g02846(.I(new_n3852_), .ZN(new_n3853_));
  NAND2_X1   g02847(.A1(\A[395] ), .A2(\A[396] ), .ZN(new_n3854_));
  AOI21_X1   g02848(.A1(new_n3853_), .A2(new_n3854_), .B(\A[394] ), .ZN(new_n3855_));
  NOR2_X1    g02849(.A1(new_n3855_), .A2(new_n3851_), .ZN(new_n3856_));
  AOI21_X1   g02850(.A1(new_n3846_), .A2(new_n3854_), .B(new_n3852_), .ZN(new_n3857_));
  AOI21_X1   g02851(.A1(new_n3835_), .A2(new_n3843_), .B(new_n3841_), .ZN(new_n3858_));
  NAND2_X1   g02852(.A1(new_n3857_), .A2(new_n3858_), .ZN(new_n3859_));
  INV_X1     g02853(.I(new_n3859_), .ZN(new_n3860_));
  NAND2_X1   g02854(.A1(new_n3834_), .A2(new_n3820_), .ZN(new_n3861_));
  AOI21_X1   g02855(.A1(new_n3792_), .A2(new_n3790_), .B(new_n3861_), .ZN(new_n3862_));
  AOI21_X1   g02856(.A1(new_n3787_), .A2(new_n3784_), .B(new_n3862_), .ZN(new_n3863_));
  NOR2_X1    g02857(.A1(new_n3791_), .A2(new_n3788_), .ZN(new_n3864_));
  AOI21_X1   g02858(.A1(new_n3774_), .A2(new_n3752_), .B(new_n3789_), .ZN(new_n3865_));
  INV_X1     g02859(.I(new_n3861_), .ZN(new_n3866_));
  OAI21_X1   g02860(.A1(new_n3865_), .A2(new_n3864_), .B(new_n3866_), .ZN(new_n3867_));
  NOR3_X1    g02861(.A1(new_n3761_), .A2(new_n3772_), .A3(new_n3867_), .ZN(new_n3868_));
  INV_X1     g02862(.I(new_n3857_), .ZN(new_n3869_));
  NOR2_X1    g02863(.A1(new_n3838_), .A2(\A[392] ), .ZN(new_n3870_));
  NOR2_X1    g02864(.A1(new_n3836_), .A2(\A[393] ), .ZN(new_n3871_));
  OAI21_X1   g02865(.A1(new_n3870_), .A2(new_n3871_), .B(\A[391] ), .ZN(new_n3872_));
  INV_X1     g02866(.I(new_n3843_), .ZN(new_n3873_));
  OAI21_X1   g02867(.A1(new_n3873_), .A2(new_n3841_), .B(new_n3835_), .ZN(new_n3874_));
  NAND2_X1   g02868(.A1(new_n3872_), .A2(new_n3874_), .ZN(new_n3875_));
  NOR2_X1    g02869(.A1(new_n3849_), .A2(\A[395] ), .ZN(new_n3876_));
  NOR2_X1    g02870(.A1(new_n3847_), .A2(\A[396] ), .ZN(new_n3877_));
  OAI21_X1   g02871(.A1(new_n3876_), .A2(new_n3877_), .B(\A[394] ), .ZN(new_n3878_));
  INV_X1     g02872(.I(new_n3854_), .ZN(new_n3879_));
  OAI21_X1   g02873(.A1(new_n3879_), .A2(new_n3852_), .B(new_n3846_), .ZN(new_n3880_));
  NAND2_X1   g02874(.A1(new_n3878_), .A2(new_n3880_), .ZN(new_n3881_));
  OAI21_X1   g02875(.A1(new_n3875_), .A2(new_n3881_), .B(new_n3858_), .ZN(new_n3882_));
  INV_X1     g02876(.I(new_n3858_), .ZN(new_n3883_));
  NAND3_X1   g02877(.A1(new_n3845_), .A2(new_n3856_), .A3(new_n3883_), .ZN(new_n3884_));
  AOI21_X1   g02878(.A1(new_n3882_), .A2(new_n3884_), .B(new_n3869_), .ZN(new_n3885_));
  NOR4_X1    g02879(.A1(new_n3840_), .A2(new_n3844_), .A3(new_n3855_), .A4(new_n3851_), .ZN(new_n3886_));
  NOR2_X1    g02880(.A1(new_n3886_), .A2(new_n3883_), .ZN(new_n3887_));
  NOR3_X1    g02881(.A1(new_n3875_), .A2(new_n3881_), .A3(new_n3858_), .ZN(new_n3888_));
  NOR3_X1    g02882(.A1(new_n3887_), .A2(new_n3888_), .A3(new_n3857_), .ZN(new_n3889_));
  NOR2_X1    g02883(.A1(new_n3889_), .A2(new_n3885_), .ZN(new_n3890_));
  NAND4_X1   g02884(.A1(new_n3807_), .A2(new_n3815_), .A3(new_n3809_), .A4(new_n3817_), .ZN(new_n3891_));
  NAND2_X1   g02885(.A1(new_n3810_), .A2(new_n3818_), .ZN(new_n3892_));
  NAND2_X1   g02886(.A1(new_n3892_), .A2(new_n3891_), .ZN(new_n3893_));
  NAND4_X1   g02887(.A1(new_n3872_), .A2(new_n3874_), .A3(new_n3878_), .A4(new_n3880_), .ZN(new_n3894_));
  OAI22_X1   g02888(.A1(new_n3840_), .A2(new_n3844_), .B1(new_n3855_), .B2(new_n3851_), .ZN(new_n3895_));
  NAND2_X1   g02889(.A1(new_n3895_), .A2(new_n3894_), .ZN(new_n3896_));
  NOR2_X1    g02890(.A1(new_n3893_), .A2(new_n3896_), .ZN(new_n3897_));
  NAND2_X1   g02891(.A1(new_n3886_), .A2(new_n3860_), .ZN(new_n3898_));
  AOI21_X1   g02892(.A1(new_n3802_), .A2(new_n3892_), .B(new_n3898_), .ZN(new_n3899_));
  XOR2_X1    g02893(.A1(new_n3796_), .A2(new_n3800_), .Z(new_n3900_));
  NAND2_X1   g02894(.A1(new_n3900_), .A2(new_n3819_), .ZN(new_n3901_));
  INV_X1     g02895(.I(new_n3796_), .ZN(new_n3902_));
  INV_X1     g02896(.I(new_n3800_), .ZN(new_n3903_));
  NAND2_X1   g02897(.A1(new_n3903_), .A2(new_n3902_), .ZN(new_n3904_));
  NAND2_X1   g02898(.A1(new_n3904_), .A2(new_n3801_), .ZN(new_n3905_));
  NAND2_X1   g02899(.A1(new_n3905_), .A2(new_n3891_), .ZN(new_n3906_));
  NAND4_X1   g02900(.A1(new_n3899_), .A2(new_n3897_), .A3(new_n3901_), .A4(new_n3906_), .ZN(new_n3907_));
  NOR2_X1    g02901(.A1(new_n3907_), .A2(new_n3890_), .ZN(new_n3908_));
  OAI21_X1   g02902(.A1(new_n3887_), .A2(new_n3888_), .B(new_n3857_), .ZN(new_n3909_));
  NAND3_X1   g02903(.A1(new_n3882_), .A2(new_n3884_), .A3(new_n3869_), .ZN(new_n3910_));
  NAND2_X1   g02904(.A1(new_n3909_), .A2(new_n3910_), .ZN(new_n3911_));
  NOR2_X1    g02905(.A1(new_n3891_), .A2(new_n3801_), .ZN(new_n3912_));
  NOR4_X1    g02906(.A1(new_n3893_), .A2(new_n3896_), .A3(new_n3898_), .A4(new_n3912_), .ZN(new_n3913_));
  NAND2_X1   g02907(.A1(new_n3911_), .A2(new_n3913_), .ZN(new_n3914_));
  NAND2_X1   g02908(.A1(new_n3891_), .A2(new_n3800_), .ZN(new_n3915_));
  NAND3_X1   g02909(.A1(new_n3826_), .A2(new_n3832_), .A3(new_n3903_), .ZN(new_n3916_));
  AOI21_X1   g02910(.A1(new_n3915_), .A2(new_n3916_), .B(new_n3902_), .ZN(new_n3917_));
  AOI21_X1   g02911(.A1(new_n3826_), .A2(new_n3832_), .B(new_n3903_), .ZN(new_n3918_));
  NOR3_X1    g02912(.A1(new_n3810_), .A2(new_n3818_), .A3(new_n3800_), .ZN(new_n3919_));
  NOR3_X1    g02913(.A1(new_n3918_), .A2(new_n3919_), .A3(new_n3796_), .ZN(new_n3920_));
  NOR2_X1    g02914(.A1(new_n3917_), .A2(new_n3920_), .ZN(new_n3921_));
  OAI21_X1   g02915(.A1(new_n3911_), .A2(new_n3913_), .B(new_n3921_), .ZN(new_n3922_));
  NOR2_X1    g02916(.A1(new_n3894_), .A2(new_n3859_), .ZN(new_n3923_));
  AOI22_X1   g02917(.A1(new_n3872_), .A2(new_n3874_), .B1(new_n3878_), .B2(new_n3880_), .ZN(new_n3924_));
  NOR2_X1    g02918(.A1(new_n3924_), .A2(new_n3886_), .ZN(new_n3925_));
  NAND4_X1   g02919(.A1(new_n3834_), .A2(new_n3820_), .A3(new_n3925_), .A4(new_n3923_), .ZN(new_n3926_));
  OAI21_X1   g02920(.A1(new_n3918_), .A2(new_n3919_), .B(new_n3796_), .ZN(new_n3927_));
  NAND3_X1   g02921(.A1(new_n3915_), .A2(new_n3916_), .A3(new_n3902_), .ZN(new_n3928_));
  NAND2_X1   g02922(.A1(new_n3928_), .A2(new_n3927_), .ZN(new_n3929_));
  NAND3_X1   g02923(.A1(new_n3890_), .A2(new_n3929_), .A3(new_n3926_), .ZN(new_n3930_));
  NAND2_X1   g02924(.A1(new_n3922_), .A2(new_n3930_), .ZN(new_n3931_));
  AOI21_X1   g02925(.A1(new_n3931_), .A2(new_n3914_), .B(new_n3908_), .ZN(new_n3932_));
  OAI22_X1   g02926(.A1(new_n3932_), .A2(new_n3773_), .B1(new_n3863_), .B2(new_n3868_), .ZN(new_n3933_));
  NAND2_X1   g02927(.A1(new_n3692_), .A2(new_n3758_), .ZN(new_n3934_));
  NAND2_X1   g02928(.A1(new_n3934_), .A2(new_n3731_), .ZN(new_n3935_));
  OAI21_X1   g02929(.A1(new_n3735_), .A2(new_n3736_), .B(new_n3740_), .ZN(new_n3936_));
  NAND2_X1   g02930(.A1(new_n3936_), .A2(new_n3751_), .ZN(new_n3937_));
  INV_X1     g02931(.I(new_n3937_), .ZN(new_n3938_));
  NAND2_X1   g02932(.A1(new_n3777_), .A2(new_n3749_), .ZN(new_n3939_));
  AOI21_X1   g02933(.A1(new_n3939_), .A2(new_n3783_), .B(new_n3938_), .ZN(new_n3940_));
  NOR2_X1    g02934(.A1(new_n3739_), .A2(new_n3780_), .ZN(new_n3941_));
  NOR3_X1    g02935(.A1(new_n3941_), .A2(new_n3760_), .A3(new_n3937_), .ZN(new_n3942_));
  OAI21_X1   g02936(.A1(new_n3942_), .A2(new_n3940_), .B(new_n3935_), .ZN(new_n3943_));
  INV_X1     g02937(.I(new_n3935_), .ZN(new_n3944_));
  OAI21_X1   g02938(.A1(new_n3941_), .A2(new_n3760_), .B(new_n3937_), .ZN(new_n3945_));
  NAND3_X1   g02939(.A1(new_n3939_), .A2(new_n3783_), .A3(new_n3938_), .ZN(new_n3946_));
  NAND3_X1   g02940(.A1(new_n3945_), .A2(new_n3946_), .A3(new_n3944_), .ZN(new_n3947_));
  NAND2_X1   g02941(.A1(new_n3943_), .A2(new_n3947_), .ZN(new_n3948_));
  AOI21_X1   g02942(.A1(new_n3819_), .A2(new_n3904_), .B(new_n3802_), .ZN(new_n3949_));
  INV_X1     g02943(.I(new_n3907_), .ZN(new_n3950_));
  OAI21_X1   g02944(.A1(new_n3857_), .A2(new_n3858_), .B(new_n3886_), .ZN(new_n3951_));
  NAND2_X1   g02945(.A1(new_n3951_), .A2(new_n3859_), .ZN(new_n3952_));
  AOI21_X1   g02946(.A1(new_n3926_), .A2(new_n3921_), .B(new_n3890_), .ZN(new_n3953_));
  OAI21_X1   g02947(.A1(new_n3953_), .A2(new_n3950_), .B(new_n3952_), .ZN(new_n3954_));
  INV_X1     g02948(.I(new_n3952_), .ZN(new_n3955_));
  OAI21_X1   g02949(.A1(new_n3913_), .A2(new_n3929_), .B(new_n3911_), .ZN(new_n3956_));
  NAND3_X1   g02950(.A1(new_n3956_), .A2(new_n3907_), .A3(new_n3955_), .ZN(new_n3957_));
  AOI21_X1   g02951(.A1(new_n3954_), .A2(new_n3957_), .B(new_n3949_), .ZN(new_n3958_));
  INV_X1     g02952(.I(new_n3949_), .ZN(new_n3959_));
  AOI21_X1   g02953(.A1(new_n3956_), .A2(new_n3907_), .B(new_n3955_), .ZN(new_n3960_));
  NOR3_X1    g02954(.A1(new_n3953_), .A2(new_n3950_), .A3(new_n3952_), .ZN(new_n3961_));
  NOR3_X1    g02955(.A1(new_n3961_), .A2(new_n3960_), .A3(new_n3959_), .ZN(new_n3962_));
  NOR2_X1    g02956(.A1(new_n3962_), .A2(new_n3958_), .ZN(new_n3963_));
  NAND2_X1   g02957(.A1(new_n3948_), .A2(new_n3963_), .ZN(new_n3964_));
  AOI21_X1   g02958(.A1(new_n3945_), .A2(new_n3946_), .B(new_n3944_), .ZN(new_n3965_));
  NOR3_X1    g02959(.A1(new_n3942_), .A2(new_n3940_), .A3(new_n3935_), .ZN(new_n3966_));
  NOR2_X1    g02960(.A1(new_n3966_), .A2(new_n3965_), .ZN(new_n3967_));
  OAI21_X1   g02961(.A1(new_n3961_), .A2(new_n3960_), .B(new_n3959_), .ZN(new_n3968_));
  NAND3_X1   g02962(.A1(new_n3954_), .A2(new_n3957_), .A3(new_n3949_), .ZN(new_n3969_));
  NAND2_X1   g02963(.A1(new_n3968_), .A2(new_n3969_), .ZN(new_n3970_));
  NAND2_X1   g02964(.A1(new_n3967_), .A2(new_n3970_), .ZN(new_n3971_));
  AOI21_X1   g02965(.A1(new_n3971_), .A2(new_n3964_), .B(new_n3933_), .ZN(new_n3972_));
  NAND2_X1   g02966(.A1(new_n3787_), .A2(new_n3784_), .ZN(new_n3973_));
  OAI21_X1   g02967(.A1(new_n3761_), .A2(new_n3772_), .B(new_n3867_), .ZN(new_n3974_));
  NAND3_X1   g02968(.A1(new_n3787_), .A2(new_n3784_), .A3(new_n3862_), .ZN(new_n3975_));
  INV_X1     g02969(.I(new_n3908_), .ZN(new_n3976_));
  AOI21_X1   g02970(.A1(new_n3890_), .A2(new_n3926_), .B(new_n3929_), .ZN(new_n3977_));
  NOR3_X1    g02971(.A1(new_n3911_), .A2(new_n3921_), .A3(new_n3913_), .ZN(new_n3978_));
  OAI21_X1   g02972(.A1(new_n3977_), .A2(new_n3978_), .B(new_n3914_), .ZN(new_n3979_));
  NAND2_X1   g02973(.A1(new_n3979_), .A2(new_n3976_), .ZN(new_n3980_));
  AOI22_X1   g02974(.A1(new_n3980_), .A2(new_n3973_), .B1(new_n3974_), .B2(new_n3975_), .ZN(new_n3981_));
  NAND2_X1   g02975(.A1(new_n3967_), .A2(new_n3963_), .ZN(new_n3982_));
  NAND2_X1   g02976(.A1(new_n3948_), .A2(new_n3970_), .ZN(new_n3983_));
  AOI21_X1   g02977(.A1(new_n3982_), .A2(new_n3983_), .B(new_n3981_), .ZN(new_n3984_));
  NOR3_X1    g02978(.A1(new_n3652_), .A2(new_n3972_), .A3(new_n3984_), .ZN(new_n3985_));
  INV_X1     g02979(.I(new_n3985_), .ZN(new_n3986_));
  INV_X1     g02980(.I(new_n3620_), .ZN(new_n3987_));
  NAND2_X1   g02981(.A1(new_n3987_), .A2(new_n3622_), .ZN(new_n3988_));
  NOR2_X1    g02982(.A1(new_n3618_), .A2(new_n3469_), .ZN(new_n3989_));
  OAI21_X1   g02983(.A1(new_n3987_), .A2(new_n3622_), .B(new_n3989_), .ZN(new_n3990_));
  NAND2_X1   g02984(.A1(new_n3990_), .A2(new_n3988_), .ZN(new_n3991_));
  AOI21_X1   g02985(.A1(new_n3644_), .A2(new_n3648_), .B(new_n3649_), .ZN(new_n3992_));
  INV_X1     g02986(.I(new_n3630_), .ZN(new_n3993_));
  NAND2_X1   g02987(.A1(new_n3993_), .A2(new_n3632_), .ZN(new_n3994_));
  NOR2_X1    g02988(.A1(new_n3993_), .A2(new_n3632_), .ZN(new_n3995_));
  OR3_X2     g02989(.A1(new_n3628_), .A2(new_n3626_), .A3(new_n3995_), .Z(new_n3996_));
  NAND2_X1   g02990(.A1(new_n3996_), .A2(new_n3994_), .ZN(new_n3997_));
  INV_X1     g02991(.I(new_n3997_), .ZN(new_n3998_));
  NOR2_X1    g02992(.A1(new_n3992_), .A2(new_n3998_), .ZN(new_n3999_));
  NOR4_X1    g02993(.A1(new_n3644_), .A2(new_n3646_), .A3(new_n3647_), .A4(new_n3997_), .ZN(new_n4000_));
  OAI21_X1   g02994(.A1(new_n3999_), .A2(new_n4000_), .B(new_n3991_), .ZN(new_n4001_));
  INV_X1     g02995(.I(new_n3991_), .ZN(new_n4002_));
  NAND3_X1   g02996(.A1(new_n3617_), .A2(new_n3625_), .A3(new_n3634_), .ZN(new_n4003_));
  NAND2_X1   g02997(.A1(new_n4003_), .A2(new_n3997_), .ZN(new_n4004_));
  NAND4_X1   g02998(.A1(new_n3998_), .A2(new_n3617_), .A3(new_n3625_), .A4(new_n3634_), .ZN(new_n4005_));
  NAND3_X1   g02999(.A1(new_n4004_), .A2(new_n4002_), .A3(new_n4005_), .ZN(new_n4006_));
  NAND2_X1   g03000(.A1(new_n4001_), .A2(new_n4006_), .ZN(new_n4007_));
  NAND2_X1   g03001(.A1(new_n3939_), .A2(new_n3783_), .ZN(new_n4008_));
  NAND2_X1   g03002(.A1(new_n3937_), .A2(new_n3935_), .ZN(new_n4009_));
  NOR2_X1    g03003(.A1(new_n3937_), .A2(new_n3935_), .ZN(new_n4010_));
  OAI21_X1   g03004(.A1(new_n4008_), .A2(new_n4010_), .B(new_n4009_), .ZN(new_n4011_));
  NAND2_X1   g03005(.A1(new_n3956_), .A2(new_n3907_), .ZN(new_n4012_));
  NOR2_X1    g03006(.A1(new_n3952_), .A2(new_n3959_), .ZN(new_n4013_));
  NOR2_X1    g03007(.A1(new_n4012_), .A2(new_n4013_), .ZN(new_n4014_));
  AOI21_X1   g03008(.A1(new_n3959_), .A2(new_n3952_), .B(new_n4014_), .ZN(new_n4015_));
  OAI21_X1   g03009(.A1(new_n3948_), .A2(new_n3970_), .B(new_n3933_), .ZN(new_n4016_));
  XOR2_X1    g03010(.A1(new_n3937_), .A2(new_n3935_), .Z(new_n4017_));
  XOR2_X1    g03011(.A1(new_n3952_), .A2(new_n3959_), .Z(new_n4018_));
  NOR4_X1    g03012(.A1(new_n4008_), .A2(new_n4012_), .A3(new_n4017_), .A4(new_n4018_), .ZN(new_n4019_));
  AOI21_X1   g03013(.A1(new_n4016_), .A2(new_n4019_), .B(new_n4015_), .ZN(new_n4020_));
  INV_X1     g03014(.I(new_n4015_), .ZN(new_n4021_));
  AOI21_X1   g03015(.A1(new_n3967_), .A2(new_n3963_), .B(new_n3981_), .ZN(new_n4022_));
  INV_X1     g03016(.I(new_n4019_), .ZN(new_n4023_));
  NOR3_X1    g03017(.A1(new_n4022_), .A2(new_n4021_), .A3(new_n4023_), .ZN(new_n4024_));
  OAI21_X1   g03018(.A1(new_n4024_), .A2(new_n4020_), .B(new_n4011_), .ZN(new_n4025_));
  INV_X1     g03019(.I(new_n4011_), .ZN(new_n4026_));
  OAI21_X1   g03020(.A1(new_n4022_), .A2(new_n4023_), .B(new_n4021_), .ZN(new_n4027_));
  NAND3_X1   g03021(.A1(new_n4016_), .A2(new_n4015_), .A3(new_n4019_), .ZN(new_n4028_));
  NAND3_X1   g03022(.A1(new_n4027_), .A2(new_n4028_), .A3(new_n4026_), .ZN(new_n4029_));
  NAND3_X1   g03023(.A1(new_n4007_), .A2(new_n4025_), .A3(new_n4029_), .ZN(new_n4030_));
  AOI21_X1   g03024(.A1(new_n4004_), .A2(new_n4005_), .B(new_n4002_), .ZN(new_n4031_));
  NOR3_X1    g03025(.A1(new_n3999_), .A2(new_n3991_), .A3(new_n4000_), .ZN(new_n4032_));
  NOR2_X1    g03026(.A1(new_n4032_), .A2(new_n4031_), .ZN(new_n4033_));
  NAND2_X1   g03027(.A1(new_n4025_), .A2(new_n4029_), .ZN(new_n4034_));
  NAND2_X1   g03028(.A1(new_n4034_), .A2(new_n4033_), .ZN(new_n4035_));
  AOI21_X1   g03029(.A1(new_n4035_), .A2(new_n4030_), .B(new_n3986_), .ZN(new_n4036_));
  NAND4_X1   g03030(.A1(new_n4025_), .A2(new_n4029_), .A3(new_n4001_), .A4(new_n4006_), .ZN(new_n4037_));
  AOI21_X1   g03031(.A1(new_n4027_), .A2(new_n4028_), .B(new_n4026_), .ZN(new_n4038_));
  NOR3_X1    g03032(.A1(new_n4024_), .A2(new_n4020_), .A3(new_n4011_), .ZN(new_n4039_));
  OAI22_X1   g03033(.A1(new_n4038_), .A2(new_n4039_), .B1(new_n4032_), .B2(new_n4031_), .ZN(new_n4040_));
  AOI21_X1   g03034(.A1(new_n4040_), .A2(new_n4037_), .B(new_n3985_), .ZN(new_n4041_));
  NOR4_X1    g03035(.A1(new_n4036_), .A2(new_n3319_), .A3(new_n3335_), .A4(new_n4041_), .ZN(new_n4042_));
  OAI21_X1   g03036(.A1(new_n3972_), .A2(new_n3984_), .B(new_n3652_), .ZN(new_n4043_));
  INV_X1     g03037(.I(new_n4043_), .ZN(new_n4044_));
  NOR2_X1    g03038(.A1(new_n4044_), .A2(new_n3985_), .ZN(new_n4045_));
  AOI21_X1   g03039(.A1(new_n3325_), .A2(new_n3328_), .B(new_n2907_), .ZN(new_n4046_));
  NOR3_X1    g03040(.A1(new_n3322_), .A2(new_n3232_), .A3(new_n3244_), .ZN(new_n4047_));
  OAI21_X1   g03041(.A1(new_n4047_), .A2(new_n4046_), .B(new_n3266_), .ZN(new_n4048_));
  AOI21_X1   g03042(.A1(new_n3329_), .A2(new_n3267_), .B(new_n3266_), .ZN(new_n4049_));
  INV_X1     g03043(.I(new_n4049_), .ZN(new_n4050_));
  NAND3_X1   g03044(.A1(new_n4045_), .A2(new_n4050_), .A3(new_n4048_), .ZN(new_n4051_));
  NAND2_X1   g03045(.A1(new_n3261_), .A2(new_n3262_), .ZN(new_n4052_));
  NOR2_X1    g03046(.A1(new_n4052_), .A2(new_n3265_), .ZN(new_n4053_));
  NOR2_X1    g03047(.A1(new_n3896_), .A2(new_n3898_), .ZN(new_n4054_));
  INV_X1     g03048(.I(new_n4054_), .ZN(new_n4055_));
  NAND2_X1   g03049(.A1(new_n3834_), .A2(new_n3820_), .ZN(new_n4056_));
  XOR2_X1    g03050(.A1(new_n4056_), .A2(new_n3789_), .Z(new_n4057_));
  NAND2_X1   g03051(.A1(new_n4057_), .A2(new_n4055_), .ZN(new_n4058_));
  XOR2_X1    g03052(.A1(new_n4056_), .A2(new_n3788_), .Z(new_n4059_));
  NAND2_X1   g03053(.A1(new_n4059_), .A2(new_n4054_), .ZN(new_n4060_));
  AOI22_X1   g03054(.A1(new_n4058_), .A2(new_n4060_), .B1(new_n3774_), .B2(new_n3752_), .ZN(new_n4061_));
  NOR2_X1    g03055(.A1(new_n4059_), .A2(new_n4054_), .ZN(new_n4062_));
  NOR2_X1    g03056(.A1(new_n4057_), .A2(new_n4055_), .ZN(new_n4063_));
  NOR3_X1    g03057(.A1(new_n4062_), .A2(new_n4063_), .A3(new_n3791_), .ZN(new_n4064_));
  NAND2_X1   g03058(.A1(new_n3549_), .A2(new_n3544_), .ZN(new_n4065_));
  NAND2_X1   g03059(.A1(new_n4065_), .A2(new_n3545_), .ZN(new_n4066_));
  NOR3_X1    g03060(.A1(new_n4061_), .A2(new_n4064_), .A3(new_n4066_), .ZN(new_n4067_));
  INV_X1     g03061(.I(new_n4067_), .ZN(new_n4068_));
  OAI21_X1   g03062(.A1(new_n4061_), .A2(new_n4064_), .B(new_n4066_), .ZN(new_n4069_));
  NOR2_X1    g03063(.A1(new_n3251_), .A2(new_n3254_), .ZN(new_n4070_));
  NOR2_X1    g03064(.A1(new_n3257_), .A2(new_n3259_), .ZN(new_n4071_));
  NOR2_X1    g03065(.A1(new_n4070_), .A2(new_n4071_), .ZN(new_n4072_));
  NOR2_X1    g03066(.A1(new_n4072_), .A2(new_n3260_), .ZN(new_n4073_));
  NAND3_X1   g03067(.A1(new_n4068_), .A2(new_n4073_), .A3(new_n4069_), .ZN(new_n4074_));
  INV_X1     g03068(.I(new_n4074_), .ZN(new_n4075_));
  NOR2_X1    g03069(.A1(new_n4053_), .A2(new_n4075_), .ZN(new_n4076_));
  NOR3_X1    g03070(.A1(new_n4052_), .A2(new_n4074_), .A3(new_n3265_), .ZN(new_n4077_));
  NOR2_X1    g03071(.A1(new_n3639_), .A2(new_n3638_), .ZN(new_n4078_));
  NOR2_X1    g03072(.A1(new_n4078_), .A2(new_n3616_), .ZN(new_n4079_));
  INV_X1     g03073(.I(new_n4079_), .ZN(new_n4080_));
  NOR3_X1    g03074(.A1(new_n3980_), .A2(new_n3863_), .A3(new_n3868_), .ZN(new_n4081_));
  INV_X1     g03075(.I(new_n4081_), .ZN(new_n4082_));
  NAND2_X1   g03076(.A1(new_n4078_), .A2(new_n3616_), .ZN(new_n4083_));
  NAND3_X1   g03077(.A1(new_n4080_), .A2(new_n4082_), .A3(new_n4083_), .ZN(new_n4084_));
  INV_X1     g03078(.I(new_n4083_), .ZN(new_n4085_));
  OAI21_X1   g03079(.A1(new_n4085_), .A2(new_n4079_), .B(new_n4081_), .ZN(new_n4086_));
  AOI21_X1   g03080(.A1(new_n4086_), .A2(new_n4084_), .B(new_n4067_), .ZN(new_n4087_));
  NOR3_X1    g03081(.A1(new_n4085_), .A2(new_n4079_), .A3(new_n4081_), .ZN(new_n4088_));
  AOI21_X1   g03082(.A1(new_n4080_), .A2(new_n4083_), .B(new_n4082_), .ZN(new_n4089_));
  NOR3_X1    g03083(.A1(new_n4089_), .A2(new_n4088_), .A3(new_n4068_), .ZN(new_n4090_));
  NOR2_X1    g03084(.A1(new_n4087_), .A2(new_n4090_), .ZN(new_n4091_));
  OAI22_X1   g03085(.A1(new_n4091_), .A2(new_n4053_), .B1(new_n4076_), .B2(new_n4077_), .ZN(new_n4092_));
  AOI21_X1   g03086(.A1(new_n4048_), .A2(new_n4050_), .B(new_n4045_), .ZN(new_n4093_));
  OAI21_X1   g03087(.A1(new_n4093_), .A2(new_n4092_), .B(new_n4051_), .ZN(new_n4094_));
  OAI22_X1   g03088(.A1(new_n4036_), .A2(new_n4041_), .B1(new_n3319_), .B2(new_n3335_), .ZN(new_n4095_));
  AOI21_X1   g03089(.A1(new_n4094_), .A2(new_n4095_), .B(new_n4042_), .ZN(new_n4096_));
  NOR3_X1    g03090(.A1(new_n3317_), .A2(new_n3290_), .A3(new_n3286_), .ZN(new_n4097_));
  NAND2_X1   g03091(.A1(new_n3284_), .A2(new_n3277_), .ZN(new_n4098_));
  XOR2_X1    g03092(.A1(new_n3294_), .A2(new_n3301_), .Z(new_n4099_));
  XOR2_X1    g03093(.A1(new_n3272_), .A2(new_n3281_), .Z(new_n4100_));
  NOR4_X1    g03094(.A1(new_n4098_), .A2(new_n4100_), .A3(new_n4099_), .A4(new_n3297_), .ZN(new_n4101_));
  OAI21_X1   g03095(.A1(new_n4097_), .A2(new_n3332_), .B(new_n4101_), .ZN(new_n4102_));
  NOR2_X1    g03096(.A1(new_n3287_), .A2(new_n3282_), .ZN(new_n4103_));
  INV_X1     g03097(.I(new_n4103_), .ZN(new_n4104_));
  NOR2_X1    g03098(.A1(new_n3272_), .A2(new_n3281_), .ZN(new_n4105_));
  OR3_X2     g03099(.A1(new_n3273_), .A2(new_n3278_), .A3(new_n4105_), .Z(new_n4106_));
  NAND2_X1   g03100(.A1(new_n3294_), .A2(new_n3301_), .ZN(new_n4107_));
  NAND4_X1   g03101(.A1(new_n3293_), .A2(new_n3291_), .A3(new_n3298_), .A4(new_n3300_), .ZN(new_n4108_));
  NAND3_X1   g03102(.A1(new_n3304_), .A2(new_n3303_), .A3(new_n4108_), .ZN(new_n4109_));
  NAND4_X1   g03103(.A1(new_n4106_), .A2(new_n4104_), .A3(new_n4107_), .A4(new_n4109_), .ZN(new_n4110_));
  NOR2_X1    g03104(.A1(new_n4098_), .A2(new_n4105_), .ZN(new_n4111_));
  NAND2_X1   g03105(.A1(new_n4109_), .A2(new_n4107_), .ZN(new_n4112_));
  OAI21_X1   g03106(.A1(new_n4111_), .A2(new_n4103_), .B(new_n4112_), .ZN(new_n4113_));
  AND2_X2    g03107(.A1(new_n4110_), .A2(new_n4113_), .Z(new_n4114_));
  NAND2_X1   g03108(.A1(new_n4102_), .A2(new_n4114_), .ZN(new_n4115_));
  NAND2_X1   g03109(.A1(new_n3333_), .A2(new_n3268_), .ZN(new_n4116_));
  NAND2_X1   g03110(.A1(new_n4110_), .A2(new_n4113_), .ZN(new_n4117_));
  NAND3_X1   g03111(.A1(new_n4116_), .A2(new_n4101_), .A3(new_n4117_), .ZN(new_n4118_));
  NAND2_X1   g03112(.A1(new_n4115_), .A2(new_n4118_), .ZN(new_n4119_));
  NAND2_X1   g03113(.A1(new_n4016_), .A2(new_n4019_), .ZN(new_n4120_));
  NAND2_X1   g03114(.A1(new_n4015_), .A2(new_n4026_), .ZN(new_n4121_));
  NOR2_X1    g03115(.A1(new_n4015_), .A2(new_n4026_), .ZN(new_n4122_));
  AOI21_X1   g03116(.A1(new_n4120_), .A2(new_n4121_), .B(new_n4122_), .ZN(new_n4123_));
  INV_X1     g03117(.I(new_n4123_), .ZN(new_n4124_));
  NOR2_X1    g03118(.A1(new_n3991_), .A2(new_n3997_), .ZN(new_n4125_));
  NAND2_X1   g03119(.A1(new_n3991_), .A2(new_n3997_), .ZN(new_n4126_));
  AOI21_X1   g03120(.A1(new_n3992_), .A2(new_n4126_), .B(new_n4125_), .ZN(new_n4127_));
  INV_X1     g03121(.I(new_n4127_), .ZN(new_n4128_));
  OAI21_X1   g03122(.A1(new_n4034_), .A2(new_n4007_), .B(new_n3986_), .ZN(new_n4129_));
  XOR2_X1    g03123(.A1(new_n3991_), .A2(new_n3997_), .Z(new_n4130_));
  XOR2_X1    g03124(.A1(new_n4015_), .A2(new_n4026_), .Z(new_n4131_));
  NOR4_X1    g03125(.A1(new_n4130_), .A2(new_n4003_), .A3(new_n4120_), .A4(new_n4131_), .ZN(new_n4132_));
  AOI21_X1   g03126(.A1(new_n4129_), .A2(new_n4132_), .B(new_n4128_), .ZN(new_n4133_));
  NOR2_X1    g03127(.A1(new_n4039_), .A2(new_n4038_), .ZN(new_n4134_));
  AOI21_X1   g03128(.A1(new_n4134_), .A2(new_n4033_), .B(new_n3985_), .ZN(new_n4135_));
  INV_X1     g03129(.I(new_n4132_), .ZN(new_n4136_));
  NOR3_X1    g03130(.A1(new_n4135_), .A2(new_n4127_), .A3(new_n4136_), .ZN(new_n4137_));
  OAI21_X1   g03131(.A1(new_n4137_), .A2(new_n4133_), .B(new_n4124_), .ZN(new_n4138_));
  OAI21_X1   g03132(.A1(new_n4135_), .A2(new_n4136_), .B(new_n4127_), .ZN(new_n4139_));
  NAND3_X1   g03133(.A1(new_n4129_), .A2(new_n4128_), .A3(new_n4132_), .ZN(new_n4140_));
  NAND3_X1   g03134(.A1(new_n4139_), .A2(new_n4140_), .A3(new_n4123_), .ZN(new_n4141_));
  NAND3_X1   g03135(.A1(new_n4119_), .A2(new_n4138_), .A3(new_n4141_), .ZN(new_n4142_));
  AOI21_X1   g03136(.A1(new_n4116_), .A2(new_n4101_), .B(new_n4117_), .ZN(new_n4143_));
  NOR2_X1    g03137(.A1(new_n4102_), .A2(new_n4114_), .ZN(new_n4144_));
  NOR2_X1    g03138(.A1(new_n4144_), .A2(new_n4143_), .ZN(new_n4145_));
  AOI21_X1   g03139(.A1(new_n4139_), .A2(new_n4140_), .B(new_n4123_), .ZN(new_n4146_));
  NOR3_X1    g03140(.A1(new_n4137_), .A2(new_n4133_), .A3(new_n4124_), .ZN(new_n4147_));
  OAI21_X1   g03141(.A1(new_n4146_), .A2(new_n4147_), .B(new_n4145_), .ZN(new_n4148_));
  AOI21_X1   g03142(.A1(new_n4148_), .A2(new_n4142_), .B(new_n4096_), .ZN(new_n4149_));
  AOI21_X1   g03143(.A1(new_n3313_), .A2(new_n3314_), .B(new_n3317_), .ZN(new_n4150_));
  NOR3_X1    g03144(.A1(new_n3311_), .A2(new_n3286_), .A3(new_n3290_), .ZN(new_n4151_));
  OAI21_X1   g03145(.A1(new_n4150_), .A2(new_n4151_), .B(new_n3332_), .ZN(new_n4152_));
  AOI22_X1   g03146(.A1(new_n3313_), .A2(new_n3314_), .B1(new_n3315_), .B2(new_n3316_), .ZN(new_n4153_));
  OAI21_X1   g03147(.A1(new_n4153_), .A2(new_n4097_), .B(new_n3268_), .ZN(new_n4154_));
  NOR2_X1    g03148(.A1(new_n4034_), .A2(new_n4033_), .ZN(new_n4155_));
  NOR2_X1    g03149(.A1(new_n4134_), .A2(new_n4007_), .ZN(new_n4156_));
  OAI21_X1   g03150(.A1(new_n4156_), .A2(new_n4155_), .B(new_n3985_), .ZN(new_n4157_));
  NOR4_X1    g03151(.A1(new_n4038_), .A2(new_n4039_), .A3(new_n4032_), .A4(new_n4031_), .ZN(new_n4158_));
  AOI22_X1   g03152(.A1(new_n4025_), .A2(new_n4029_), .B1(new_n4001_), .B2(new_n4006_), .ZN(new_n4159_));
  OAI21_X1   g03153(.A1(new_n4158_), .A2(new_n4159_), .B(new_n3986_), .ZN(new_n4160_));
  NAND4_X1   g03154(.A1(new_n4157_), .A2(new_n4152_), .A3(new_n4154_), .A4(new_n4160_), .ZN(new_n4161_));
  NAND2_X1   g03155(.A1(new_n3986_), .A2(new_n4043_), .ZN(new_n4162_));
  INV_X1     g03156(.I(new_n4048_), .ZN(new_n4163_));
  NOR3_X1    g03157(.A1(new_n4163_), .A2(new_n4162_), .A3(new_n4049_), .ZN(new_n4164_));
  NOR2_X1    g03158(.A1(new_n4076_), .A2(new_n4077_), .ZN(new_n4165_));
  NAND2_X1   g03159(.A1(new_n4053_), .A2(new_n4075_), .ZN(new_n4166_));
  OR2_X2     g03160(.A1(new_n4087_), .A2(new_n4090_), .Z(new_n4167_));
  OAI21_X1   g03161(.A1(new_n4167_), .A2(new_n4165_), .B(new_n4166_), .ZN(new_n4168_));
  OAI21_X1   g03162(.A1(new_n4163_), .A2(new_n4049_), .B(new_n4162_), .ZN(new_n4169_));
  AOI21_X1   g03163(.A1(new_n4168_), .A2(new_n4169_), .B(new_n4164_), .ZN(new_n4170_));
  AOI22_X1   g03164(.A1(new_n4157_), .A2(new_n4160_), .B1(new_n4152_), .B2(new_n4154_), .ZN(new_n4171_));
  OAI21_X1   g03165(.A1(new_n4170_), .A2(new_n4171_), .B(new_n4161_), .ZN(new_n4172_));
  NAND3_X1   g03166(.A1(new_n4145_), .A2(new_n4138_), .A3(new_n4141_), .ZN(new_n4173_));
  OAI21_X1   g03167(.A1(new_n4146_), .A2(new_n4147_), .B(new_n4119_), .ZN(new_n4174_));
  AOI21_X1   g03168(.A1(new_n4174_), .A2(new_n4173_), .B(new_n4172_), .ZN(new_n4175_));
  NOR4_X1    g03169(.A1(new_n4149_), .A2(new_n4175_), .A3(new_n2573_), .A4(new_n2596_), .ZN(new_n4176_));
  NAND2_X1   g03170(.A1(new_n4152_), .A2(new_n4154_), .ZN(new_n4177_));
  NOR2_X1    g03171(.A1(new_n4036_), .A2(new_n4041_), .ZN(new_n4178_));
  NOR2_X1    g03172(.A1(new_n4178_), .A2(new_n4177_), .ZN(new_n4179_));
  NOR2_X1    g03173(.A1(new_n3319_), .A2(new_n3335_), .ZN(new_n4180_));
  NAND2_X1   g03174(.A1(new_n4157_), .A2(new_n4160_), .ZN(new_n4181_));
  NOR2_X1    g03175(.A1(new_n4181_), .A2(new_n4180_), .ZN(new_n4182_));
  OAI21_X1   g03176(.A1(new_n4182_), .A2(new_n4179_), .B(new_n4094_), .ZN(new_n4183_));
  OAI21_X1   g03177(.A1(new_n4171_), .A2(new_n4042_), .B(new_n4170_), .ZN(new_n4184_));
  NAND2_X1   g03178(.A1(new_n2576_), .A2(new_n2578_), .ZN(new_n4185_));
  NOR2_X1    g03179(.A1(new_n2464_), .A2(new_n2485_), .ZN(new_n4186_));
  NOR2_X1    g03180(.A1(new_n4186_), .A2(new_n4185_), .ZN(new_n4187_));
  NOR2_X1    g03181(.A1(new_n1724_), .A2(new_n1742_), .ZN(new_n4188_));
  NAND2_X1   g03182(.A1(new_n2581_), .A2(new_n2584_), .ZN(new_n4189_));
  NOR2_X1    g03183(.A1(new_n4189_), .A2(new_n4188_), .ZN(new_n4190_));
  OAI21_X1   g03184(.A1(new_n4190_), .A2(new_n4187_), .B(new_n2517_), .ZN(new_n4191_));
  OAI21_X1   g03185(.A1(new_n2486_), .A2(new_n2592_), .B(new_n2591_), .ZN(new_n4192_));
  NAND4_X1   g03186(.A1(new_n4183_), .A2(new_n4191_), .A3(new_n4184_), .A4(new_n4192_), .ZN(new_n4193_));
  INV_X1     g03187(.I(new_n2586_), .ZN(new_n4194_));
  NAND2_X1   g03188(.A1(new_n4194_), .A2(new_n2587_), .ZN(new_n4195_));
  OAI21_X1   g03189(.A1(new_n1633_), .A2(new_n1647_), .B(new_n1729_), .ZN(new_n4196_));
  NAND3_X1   g03190(.A1(new_n1732_), .A2(new_n1735_), .A3(new_n1316_), .ZN(new_n4197_));
  AOI21_X1   g03191(.A1(new_n4196_), .A2(new_n4197_), .B(new_n1737_), .ZN(new_n4198_));
  AOI21_X1   g03192(.A1(new_n1736_), .A2(new_n1671_), .B(new_n1670_), .ZN(new_n4199_));
  NOR2_X1    g03193(.A1(new_n4198_), .A2(new_n4199_), .ZN(new_n4200_));
  NAND2_X1   g03194(.A1(new_n4200_), .A2(new_n2586_), .ZN(new_n4201_));
  AOI21_X1   g03195(.A1(new_n4195_), .A2(new_n4201_), .B(new_n2515_), .ZN(new_n4202_));
  AOI21_X1   g03196(.A1(new_n2497_), .A2(new_n2590_), .B(new_n2589_), .ZN(new_n4203_));
  OAI21_X1   g03197(.A1(new_n4163_), .A2(new_n4049_), .B(new_n4045_), .ZN(new_n4204_));
  NAND3_X1   g03198(.A1(new_n4050_), .A2(new_n4162_), .A3(new_n4048_), .ZN(new_n4205_));
  AOI21_X1   g03199(.A1(new_n4204_), .A2(new_n4205_), .B(new_n4092_), .ZN(new_n4206_));
  AOI21_X1   g03200(.A1(new_n4051_), .A2(new_n4169_), .B(new_n4168_), .ZN(new_n4207_));
  NOR4_X1    g03201(.A1(new_n4202_), .A2(new_n4203_), .A3(new_n4206_), .A4(new_n4207_), .ZN(new_n4208_));
  NAND2_X1   g03202(.A1(new_n4165_), .A2(new_n4091_), .ZN(new_n4209_));
  AOI21_X1   g03203(.A1(new_n4068_), .A2(new_n4069_), .B(new_n4073_), .ZN(new_n4210_));
  INV_X1     g03204(.I(new_n4210_), .ZN(new_n4211_));
  NAND2_X1   g03205(.A1(new_n4211_), .A2(new_n4074_), .ZN(new_n4212_));
  AOI21_X1   g03206(.A1(new_n2401_), .A2(new_n2506_), .B(new_n2503_), .ZN(new_n4213_));
  NOR2_X1    g03207(.A1(new_n4213_), .A2(new_n2510_), .ZN(new_n4214_));
  INV_X1     g03208(.I(new_n4214_), .ZN(new_n4215_));
  NOR2_X1    g03209(.A1(new_n4212_), .A2(new_n4215_), .ZN(new_n4216_));
  INV_X1     g03210(.I(new_n4216_), .ZN(new_n4217_));
  XOR2_X1    g03211(.A1(new_n4209_), .A2(new_n4217_), .Z(new_n4218_));
  XOR2_X1    g03212(.A1(new_n2514_), .A2(new_n2512_), .Z(new_n4219_));
  INV_X1     g03213(.I(new_n4219_), .ZN(new_n4220_));
  AOI21_X1   g03214(.A1(new_n4209_), .A2(new_n4220_), .B(new_n4218_), .ZN(new_n4221_));
  OAI22_X1   g03215(.A1(new_n4202_), .A2(new_n4203_), .B1(new_n4206_), .B2(new_n4207_), .ZN(new_n4222_));
  AOI21_X1   g03216(.A1(new_n4221_), .A2(new_n4222_), .B(new_n4208_), .ZN(new_n4223_));
  AOI22_X1   g03217(.A1(new_n4183_), .A2(new_n4184_), .B1(new_n4191_), .B2(new_n4192_), .ZN(new_n4224_));
  OAI21_X1   g03218(.A1(new_n4224_), .A2(new_n4223_), .B(new_n4193_), .ZN(new_n4225_));
  OAI22_X1   g03219(.A1(new_n4149_), .A2(new_n4175_), .B1(new_n2573_), .B2(new_n2596_), .ZN(new_n4226_));
  AOI21_X1   g03220(.A1(new_n4225_), .A2(new_n4226_), .B(new_n4176_), .ZN(new_n4227_));
  INV_X1     g03221(.I(new_n2525_), .ZN(new_n4228_));
  NAND2_X1   g03222(.A1(new_n2529_), .A2(new_n2527_), .ZN(new_n4229_));
  NAND2_X1   g03223(.A1(new_n1692_), .A2(new_n1687_), .ZN(new_n4230_));
  NAND2_X1   g03224(.A1(new_n2527_), .A2(new_n2521_), .ZN(new_n4231_));
  AND4_X2    g03225(.A1(new_n4230_), .A2(new_n4231_), .A3(new_n2530_), .A4(new_n2532_), .Z(new_n4232_));
  OAI22_X1   g03226(.A1(new_n4228_), .A2(new_n4232_), .B1(new_n4229_), .B2(new_n2534_), .ZN(new_n4233_));
  NAND2_X1   g03227(.A1(new_n2554_), .A2(new_n2557_), .ZN(new_n4234_));
  NAND2_X1   g03228(.A1(new_n2549_), .A2(new_n2428_), .ZN(new_n4235_));
  NAND2_X1   g03229(.A1(new_n2544_), .A2(new_n2438_), .ZN(new_n4236_));
  NAND4_X1   g03230(.A1(new_n4235_), .A2(new_n2545_), .A3(new_n2550_), .A4(new_n4236_), .ZN(new_n4237_));
  AOI22_X1   g03231(.A1(new_n4234_), .A2(new_n4237_), .B1(new_n2548_), .B2(new_n2552_), .ZN(new_n4238_));
  INV_X1     g03232(.I(new_n4238_), .ZN(new_n4239_));
  OAI21_X1   g03233(.A1(new_n4186_), .A2(new_n4188_), .B(new_n2517_), .ZN(new_n4240_));
  NAND3_X1   g03234(.A1(new_n2594_), .A2(new_n2585_), .A3(new_n4240_), .ZN(new_n4241_));
  XOR2_X1    g03235(.A1(new_n2552_), .A2(new_n2548_), .Z(new_n4242_));
  NOR4_X1    g03236(.A1(new_n4234_), .A2(new_n4242_), .A3(new_n2525_), .A4(new_n2538_), .ZN(new_n4243_));
  AOI21_X1   g03237(.A1(new_n4241_), .A2(new_n4243_), .B(new_n4239_), .ZN(new_n4244_));
  NOR3_X1    g03238(.A1(new_n2543_), .A2(new_n2571_), .A3(new_n2570_), .ZN(new_n4245_));
  OAI21_X1   g03239(.A1(new_n4245_), .A2(new_n2593_), .B(new_n4243_), .ZN(new_n4246_));
  NOR2_X1    g03240(.A1(new_n4246_), .A2(new_n4238_), .ZN(new_n4247_));
  OAI21_X1   g03241(.A1(new_n4247_), .A2(new_n4244_), .B(new_n4233_), .ZN(new_n4248_));
  INV_X1     g03242(.I(new_n4233_), .ZN(new_n4249_));
  NAND2_X1   g03243(.A1(new_n4246_), .A2(new_n4238_), .ZN(new_n4250_));
  NAND3_X1   g03244(.A1(new_n4241_), .A2(new_n4239_), .A3(new_n4243_), .ZN(new_n4251_));
  NAND3_X1   g03245(.A1(new_n4250_), .A2(new_n4251_), .A3(new_n4249_), .ZN(new_n4252_));
  NAND2_X1   g03246(.A1(new_n4248_), .A2(new_n4252_), .ZN(new_n4253_));
  NAND2_X1   g03247(.A1(new_n3287_), .A2(new_n3282_), .ZN(new_n4254_));
  NAND2_X1   g03248(.A1(new_n4104_), .A2(new_n4098_), .ZN(new_n4255_));
  NAND4_X1   g03249(.A1(new_n4255_), .A2(new_n4254_), .A3(new_n4107_), .A4(new_n4109_), .ZN(new_n4256_));
  NAND2_X1   g03250(.A1(new_n4102_), .A2(new_n4256_), .ZN(new_n4257_));
  NAND3_X1   g03251(.A1(new_n4106_), .A2(new_n4104_), .A3(new_n4112_), .ZN(new_n4258_));
  NAND2_X1   g03252(.A1(new_n4257_), .A2(new_n4258_), .ZN(new_n4259_));
  NAND2_X1   g03253(.A1(new_n4129_), .A2(new_n4132_), .ZN(new_n4260_));
  NAND4_X1   g03254(.A1(new_n4124_), .A2(new_n3991_), .A3(new_n3992_), .A4(new_n3997_), .ZN(new_n4261_));
  AOI22_X1   g03255(.A1(new_n4260_), .A2(new_n4261_), .B1(new_n4124_), .B2(new_n4127_), .ZN(new_n4262_));
  INV_X1     g03256(.I(new_n4262_), .ZN(new_n4263_));
  NAND2_X1   g03257(.A1(new_n4173_), .A2(new_n4096_), .ZN(new_n4264_));
  XNOR2_X1   g03258(.A1(new_n4123_), .A2(new_n4127_), .ZN(new_n4265_));
  NOR4_X1    g03259(.A1(new_n4260_), .A2(new_n4102_), .A3(new_n4265_), .A4(new_n4117_), .ZN(new_n4266_));
  AOI21_X1   g03260(.A1(new_n4264_), .A2(new_n4266_), .B(new_n4263_), .ZN(new_n4267_));
  NOR3_X1    g03261(.A1(new_n4146_), .A2(new_n4147_), .A3(new_n4119_), .ZN(new_n4268_));
  OAI21_X1   g03262(.A1(new_n4268_), .A2(new_n4172_), .B(new_n4266_), .ZN(new_n4269_));
  NOR2_X1    g03263(.A1(new_n4269_), .A2(new_n4262_), .ZN(new_n4270_));
  OAI21_X1   g03264(.A1(new_n4267_), .A2(new_n4270_), .B(new_n4259_), .ZN(new_n4271_));
  INV_X1     g03265(.I(new_n4259_), .ZN(new_n4272_));
  NAND2_X1   g03266(.A1(new_n4269_), .A2(new_n4262_), .ZN(new_n4273_));
  NAND3_X1   g03267(.A1(new_n4264_), .A2(new_n4263_), .A3(new_n4266_), .ZN(new_n4274_));
  NAND3_X1   g03268(.A1(new_n4274_), .A2(new_n4273_), .A3(new_n4272_), .ZN(new_n4275_));
  NAND3_X1   g03269(.A1(new_n4253_), .A2(new_n4271_), .A3(new_n4275_), .ZN(new_n4276_));
  AOI21_X1   g03270(.A1(new_n4250_), .A2(new_n4251_), .B(new_n4249_), .ZN(new_n4277_));
  NOR3_X1    g03271(.A1(new_n4247_), .A2(new_n4244_), .A3(new_n4233_), .ZN(new_n4278_));
  NOR2_X1    g03272(.A1(new_n4278_), .A2(new_n4277_), .ZN(new_n4279_));
  NAND2_X1   g03273(.A1(new_n4271_), .A2(new_n4275_), .ZN(new_n4280_));
  NAND2_X1   g03274(.A1(new_n4280_), .A2(new_n4279_), .ZN(new_n4281_));
  AOI21_X1   g03275(.A1(new_n4281_), .A2(new_n4276_), .B(new_n4227_), .ZN(new_n4282_));
  NOR3_X1    g03276(.A1(new_n2569_), .A2(new_n2571_), .A3(new_n2570_), .ZN(new_n4283_));
  AOI21_X1   g03277(.A1(new_n2562_), .A2(new_n2565_), .B(new_n2543_), .ZN(new_n4284_));
  OAI21_X1   g03278(.A1(new_n4284_), .A2(new_n4283_), .B(new_n2593_), .ZN(new_n4285_));
  AOI21_X1   g03279(.A1(new_n2562_), .A2(new_n2565_), .B(new_n2569_), .ZN(new_n4286_));
  OAI21_X1   g03280(.A1(new_n4286_), .A2(new_n4245_), .B(new_n2519_), .ZN(new_n4287_));
  NOR3_X1    g03281(.A1(new_n4145_), .A2(new_n4147_), .A3(new_n4146_), .ZN(new_n4288_));
  AOI21_X1   g03282(.A1(new_n4138_), .A2(new_n4141_), .B(new_n4119_), .ZN(new_n4289_));
  OAI21_X1   g03283(.A1(new_n4288_), .A2(new_n4289_), .B(new_n4172_), .ZN(new_n4290_));
  AOI21_X1   g03284(.A1(new_n4138_), .A2(new_n4141_), .B(new_n4145_), .ZN(new_n4291_));
  OAI21_X1   g03285(.A1(new_n4291_), .A2(new_n4268_), .B(new_n4096_), .ZN(new_n4292_));
  NAND4_X1   g03286(.A1(new_n4290_), .A2(new_n4292_), .A3(new_n4287_), .A4(new_n4285_), .ZN(new_n4293_));
  NAND2_X1   g03287(.A1(new_n4181_), .A2(new_n4180_), .ZN(new_n4294_));
  NAND2_X1   g03288(.A1(new_n4178_), .A2(new_n4177_), .ZN(new_n4295_));
  AOI21_X1   g03289(.A1(new_n4294_), .A2(new_n4295_), .B(new_n4170_), .ZN(new_n4296_));
  AOI21_X1   g03290(.A1(new_n4095_), .A2(new_n4161_), .B(new_n4094_), .ZN(new_n4297_));
  NAND2_X1   g03291(.A1(new_n4189_), .A2(new_n4188_), .ZN(new_n4298_));
  NAND2_X1   g03292(.A1(new_n4186_), .A2(new_n4185_), .ZN(new_n4299_));
  AOI21_X1   g03293(.A1(new_n4298_), .A2(new_n4299_), .B(new_n2591_), .ZN(new_n4300_));
  AOI21_X1   g03294(.A1(new_n2518_), .A2(new_n2585_), .B(new_n2517_), .ZN(new_n4301_));
  NOR4_X1    g03295(.A1(new_n4296_), .A2(new_n4300_), .A3(new_n4297_), .A4(new_n4301_), .ZN(new_n4302_));
  NOR2_X1    g03296(.A1(new_n4200_), .A2(new_n2586_), .ZN(new_n4303_));
  NOR2_X1    g03297(.A1(new_n4194_), .A2(new_n2587_), .ZN(new_n4304_));
  OAI21_X1   g03298(.A1(new_n4304_), .A2(new_n4303_), .B(new_n2589_), .ZN(new_n4305_));
  OAI21_X1   g03299(.A1(new_n2588_), .A2(new_n2516_), .B(new_n2515_), .ZN(new_n4306_));
  AOI21_X1   g03300(.A1(new_n4050_), .A2(new_n4048_), .B(new_n4162_), .ZN(new_n4307_));
  NOR3_X1    g03301(.A1(new_n4163_), .A2(new_n4045_), .A3(new_n4049_), .ZN(new_n4308_));
  OAI21_X1   g03302(.A1(new_n4308_), .A2(new_n4307_), .B(new_n4168_), .ZN(new_n4309_));
  OAI21_X1   g03303(.A1(new_n4093_), .A2(new_n4164_), .B(new_n4092_), .ZN(new_n4310_));
  NAND4_X1   g03304(.A1(new_n4305_), .A2(new_n4309_), .A3(new_n4310_), .A4(new_n4306_), .ZN(new_n4311_));
  XOR2_X1    g03305(.A1(new_n4209_), .A2(new_n4216_), .Z(new_n4312_));
  NOR2_X1    g03306(.A1(new_n4209_), .A2(new_n4217_), .ZN(new_n4313_));
  AOI21_X1   g03307(.A1(new_n4312_), .A2(new_n4219_), .B(new_n4313_), .ZN(new_n4314_));
  AOI22_X1   g03308(.A1(new_n4305_), .A2(new_n4306_), .B1(new_n4310_), .B2(new_n4309_), .ZN(new_n4315_));
  OAI21_X1   g03309(.A1(new_n4315_), .A2(new_n4314_), .B(new_n4311_), .ZN(new_n4316_));
  OAI22_X1   g03310(.A1(new_n4296_), .A2(new_n4297_), .B1(new_n4300_), .B2(new_n4301_), .ZN(new_n4317_));
  AOI21_X1   g03311(.A1(new_n4317_), .A2(new_n4316_), .B(new_n4302_), .ZN(new_n4318_));
  AOI22_X1   g03312(.A1(new_n4290_), .A2(new_n4292_), .B1(new_n4287_), .B2(new_n4285_), .ZN(new_n4319_));
  OAI21_X1   g03313(.A1(new_n4318_), .A2(new_n4319_), .B(new_n4293_), .ZN(new_n4320_));
  NAND4_X1   g03314(.A1(new_n4271_), .A2(new_n4275_), .A3(new_n4248_), .A4(new_n4252_), .ZN(new_n4321_));
  AOI21_X1   g03315(.A1(new_n4274_), .A2(new_n4273_), .B(new_n4272_), .ZN(new_n4322_));
  NOR3_X1    g03316(.A1(new_n4267_), .A2(new_n4270_), .A3(new_n4259_), .ZN(new_n4323_));
  OAI22_X1   g03317(.A1(new_n4322_), .A2(new_n4323_), .B1(new_n4277_), .B2(new_n4278_), .ZN(new_n4324_));
  AOI21_X1   g03318(.A1(new_n4324_), .A2(new_n4321_), .B(new_n4320_), .ZN(new_n4325_));
  INV_X1     g03319(.I(\A[142] ), .ZN(new_n4326_));
  NOR2_X1    g03320(.A1(\A[143] ), .A2(\A[144] ), .ZN(new_n4327_));
  NAND2_X1   g03321(.A1(\A[143] ), .A2(\A[144] ), .ZN(new_n4328_));
  AOI21_X1   g03322(.A1(new_n4326_), .A2(new_n4328_), .B(new_n4327_), .ZN(new_n4329_));
  INV_X1     g03323(.I(\A[139] ), .ZN(new_n4330_));
  NOR2_X1    g03324(.A1(\A[140] ), .A2(\A[141] ), .ZN(new_n4331_));
  NAND2_X1   g03325(.A1(\A[140] ), .A2(\A[141] ), .ZN(new_n4332_));
  AOI21_X1   g03326(.A1(new_n4330_), .A2(new_n4332_), .B(new_n4331_), .ZN(new_n4333_));
  INV_X1     g03327(.I(new_n4333_), .ZN(new_n4334_));
  INV_X1     g03328(.I(\A[140] ), .ZN(new_n4335_));
  NAND2_X1   g03329(.A1(new_n4335_), .A2(\A[141] ), .ZN(new_n4336_));
  INV_X1     g03330(.I(\A[141] ), .ZN(new_n4337_));
  NAND2_X1   g03331(.A1(new_n4337_), .A2(\A[140] ), .ZN(new_n4338_));
  AOI21_X1   g03332(.A1(new_n4336_), .A2(new_n4338_), .B(new_n4330_), .ZN(new_n4339_));
  INV_X1     g03333(.I(new_n4331_), .ZN(new_n4340_));
  AOI21_X1   g03334(.A1(new_n4340_), .A2(new_n4332_), .B(\A[139] ), .ZN(new_n4341_));
  INV_X1     g03335(.I(\A[143] ), .ZN(new_n4342_));
  NAND2_X1   g03336(.A1(new_n4342_), .A2(\A[144] ), .ZN(new_n4343_));
  INV_X1     g03337(.I(\A[144] ), .ZN(new_n4344_));
  NAND2_X1   g03338(.A1(new_n4344_), .A2(\A[143] ), .ZN(new_n4345_));
  AOI21_X1   g03339(.A1(new_n4343_), .A2(new_n4345_), .B(new_n4326_), .ZN(new_n4346_));
  INV_X1     g03340(.I(new_n4327_), .ZN(new_n4347_));
  AOI21_X1   g03341(.A1(new_n4347_), .A2(new_n4328_), .B(\A[142] ), .ZN(new_n4348_));
  NOR4_X1    g03342(.A1(new_n4339_), .A2(new_n4341_), .A3(new_n4348_), .A4(new_n4346_), .ZN(new_n4349_));
  NOR2_X1    g03343(.A1(new_n4349_), .A2(new_n4334_), .ZN(new_n4350_));
  INV_X1     g03344(.I(new_n4336_), .ZN(new_n4351_));
  NOR2_X1    g03345(.A1(new_n4335_), .A2(\A[141] ), .ZN(new_n4352_));
  OAI21_X1   g03346(.A1(new_n4351_), .A2(new_n4352_), .B(\A[139] ), .ZN(new_n4353_));
  INV_X1     g03347(.I(new_n4332_), .ZN(new_n4354_));
  OAI21_X1   g03348(.A1(new_n4354_), .A2(new_n4331_), .B(new_n4330_), .ZN(new_n4355_));
  NOR2_X1    g03349(.A1(new_n4344_), .A2(\A[143] ), .ZN(new_n4356_));
  NOR2_X1    g03350(.A1(new_n4342_), .A2(\A[144] ), .ZN(new_n4357_));
  OAI21_X1   g03351(.A1(new_n4356_), .A2(new_n4357_), .B(\A[142] ), .ZN(new_n4358_));
  INV_X1     g03352(.I(new_n4328_), .ZN(new_n4359_));
  OAI21_X1   g03353(.A1(new_n4359_), .A2(new_n4327_), .B(new_n4326_), .ZN(new_n4360_));
  NAND4_X1   g03354(.A1(new_n4353_), .A2(new_n4355_), .A3(new_n4360_), .A4(new_n4358_), .ZN(new_n4361_));
  NOR2_X1    g03355(.A1(new_n4361_), .A2(new_n4333_), .ZN(new_n4362_));
  OAI21_X1   g03356(.A1(new_n4362_), .A2(new_n4350_), .B(new_n4329_), .ZN(new_n4363_));
  INV_X1     g03357(.I(new_n4329_), .ZN(new_n4364_));
  NAND2_X1   g03358(.A1(new_n4361_), .A2(new_n4333_), .ZN(new_n4365_));
  NAND2_X1   g03359(.A1(new_n4349_), .A2(new_n4334_), .ZN(new_n4366_));
  NAND3_X1   g03360(.A1(new_n4365_), .A2(new_n4366_), .A3(new_n4364_), .ZN(new_n4367_));
  NAND2_X1   g03361(.A1(new_n4363_), .A2(new_n4367_), .ZN(new_n4368_));
  INV_X1     g03362(.I(\A[148] ), .ZN(new_n4369_));
  NOR2_X1    g03363(.A1(\A[149] ), .A2(\A[150] ), .ZN(new_n4370_));
  NAND2_X1   g03364(.A1(\A[149] ), .A2(\A[150] ), .ZN(new_n4371_));
  AOI21_X1   g03365(.A1(new_n4369_), .A2(new_n4371_), .B(new_n4370_), .ZN(new_n4372_));
  INV_X1     g03366(.I(\A[145] ), .ZN(new_n4373_));
  NOR2_X1    g03367(.A1(\A[146] ), .A2(\A[147] ), .ZN(new_n4374_));
  NAND2_X1   g03368(.A1(\A[146] ), .A2(\A[147] ), .ZN(new_n4375_));
  AOI21_X1   g03369(.A1(new_n4373_), .A2(new_n4375_), .B(new_n4374_), .ZN(new_n4376_));
  NAND2_X1   g03370(.A1(new_n4372_), .A2(new_n4376_), .ZN(new_n4377_));
  INV_X1     g03371(.I(\A[146] ), .ZN(new_n4378_));
  NAND2_X1   g03372(.A1(new_n4378_), .A2(\A[147] ), .ZN(new_n4379_));
  INV_X1     g03373(.I(\A[147] ), .ZN(new_n4380_));
  NAND2_X1   g03374(.A1(new_n4380_), .A2(\A[146] ), .ZN(new_n4381_));
  AOI21_X1   g03375(.A1(new_n4379_), .A2(new_n4381_), .B(new_n4373_), .ZN(new_n4382_));
  INV_X1     g03376(.I(new_n4374_), .ZN(new_n4383_));
  AOI21_X1   g03377(.A1(new_n4383_), .A2(new_n4375_), .B(\A[145] ), .ZN(new_n4384_));
  NOR2_X1    g03378(.A1(new_n4384_), .A2(new_n4382_), .ZN(new_n4385_));
  INV_X1     g03379(.I(\A[150] ), .ZN(new_n4386_));
  NOR2_X1    g03380(.A1(new_n4386_), .A2(\A[149] ), .ZN(new_n4387_));
  INV_X1     g03381(.I(\A[149] ), .ZN(new_n4388_));
  NOR2_X1    g03382(.A1(new_n4388_), .A2(\A[150] ), .ZN(new_n4389_));
  OAI21_X1   g03383(.A1(new_n4387_), .A2(new_n4389_), .B(\A[148] ), .ZN(new_n4390_));
  INV_X1     g03384(.I(new_n4371_), .ZN(new_n4391_));
  OAI21_X1   g03385(.A1(new_n4391_), .A2(new_n4370_), .B(new_n4369_), .ZN(new_n4392_));
  NAND2_X1   g03386(.A1(new_n4390_), .A2(new_n4392_), .ZN(new_n4393_));
  NAND2_X1   g03387(.A1(new_n4385_), .A2(new_n4393_), .ZN(new_n4394_));
  NOR2_X1    g03388(.A1(new_n4380_), .A2(\A[146] ), .ZN(new_n4395_));
  NOR2_X1    g03389(.A1(new_n4378_), .A2(\A[147] ), .ZN(new_n4396_));
  OAI21_X1   g03390(.A1(new_n4395_), .A2(new_n4396_), .B(\A[145] ), .ZN(new_n4397_));
  INV_X1     g03391(.I(new_n4375_), .ZN(new_n4398_));
  OAI21_X1   g03392(.A1(new_n4398_), .A2(new_n4374_), .B(new_n4373_), .ZN(new_n4399_));
  NAND2_X1   g03393(.A1(new_n4397_), .A2(new_n4399_), .ZN(new_n4400_));
  NAND2_X1   g03394(.A1(new_n4388_), .A2(\A[150] ), .ZN(new_n4401_));
  NAND2_X1   g03395(.A1(new_n4386_), .A2(\A[149] ), .ZN(new_n4402_));
  AOI21_X1   g03396(.A1(new_n4401_), .A2(new_n4402_), .B(new_n4369_), .ZN(new_n4403_));
  INV_X1     g03397(.I(new_n4370_), .ZN(new_n4404_));
  AOI21_X1   g03398(.A1(new_n4404_), .A2(new_n4371_), .B(\A[148] ), .ZN(new_n4405_));
  NOR2_X1    g03399(.A1(new_n4405_), .A2(new_n4403_), .ZN(new_n4406_));
  NAND2_X1   g03400(.A1(new_n4406_), .A2(new_n4400_), .ZN(new_n4407_));
  AOI21_X1   g03401(.A1(new_n4394_), .A2(new_n4407_), .B(new_n4377_), .ZN(new_n4408_));
  INV_X1     g03402(.I(new_n4372_), .ZN(new_n4409_));
  NAND4_X1   g03403(.A1(new_n4397_), .A2(new_n4399_), .A3(new_n4390_), .A4(new_n4392_), .ZN(new_n4410_));
  NAND2_X1   g03404(.A1(new_n4410_), .A2(new_n4376_), .ZN(new_n4411_));
  INV_X1     g03405(.I(new_n4376_), .ZN(new_n4412_));
  NAND3_X1   g03406(.A1(new_n4385_), .A2(new_n4406_), .A3(new_n4412_), .ZN(new_n4413_));
  AOI21_X1   g03407(.A1(new_n4411_), .A2(new_n4413_), .B(new_n4409_), .ZN(new_n4414_));
  NOR4_X1    g03408(.A1(new_n4382_), .A2(new_n4384_), .A3(new_n4405_), .A4(new_n4403_), .ZN(new_n4415_));
  NOR2_X1    g03409(.A1(new_n4415_), .A2(new_n4412_), .ZN(new_n4416_));
  NOR3_X1    g03410(.A1(new_n4400_), .A2(new_n4393_), .A3(new_n4376_), .ZN(new_n4417_));
  NOR3_X1    g03411(.A1(new_n4416_), .A2(new_n4417_), .A3(new_n4372_), .ZN(new_n4418_));
  NOR3_X1    g03412(.A1(new_n4418_), .A2(new_n4414_), .A3(new_n4408_), .ZN(new_n4419_));
  INV_X1     g03413(.I(new_n4377_), .ZN(new_n4420_));
  NAND2_X1   g03414(.A1(new_n4415_), .A2(new_n4420_), .ZN(new_n4421_));
  NAND2_X1   g03415(.A1(new_n4400_), .A2(new_n4393_), .ZN(new_n4422_));
  NAND2_X1   g03416(.A1(new_n4422_), .A2(new_n4410_), .ZN(new_n4423_));
  OAI22_X1   g03417(.A1(new_n4339_), .A2(new_n4341_), .B1(new_n4348_), .B2(new_n4346_), .ZN(new_n4424_));
  NAND2_X1   g03418(.A1(new_n4361_), .A2(new_n4424_), .ZN(new_n4425_));
  NAND3_X1   g03419(.A1(new_n4349_), .A2(new_n4329_), .A3(new_n4333_), .ZN(new_n4426_));
  NOR4_X1    g03420(.A1(new_n4423_), .A2(new_n4425_), .A3(new_n4426_), .A4(new_n4421_), .ZN(new_n4427_));
  NAND2_X1   g03421(.A1(new_n4419_), .A2(new_n4427_), .ZN(new_n4428_));
  NOR2_X1    g03422(.A1(new_n4406_), .A2(new_n4400_), .ZN(new_n4429_));
  NOR2_X1    g03423(.A1(new_n4385_), .A2(new_n4393_), .ZN(new_n4430_));
  OAI21_X1   g03424(.A1(new_n4429_), .A2(new_n4430_), .B(new_n4420_), .ZN(new_n4431_));
  OAI21_X1   g03425(.A1(new_n4416_), .A2(new_n4417_), .B(new_n4372_), .ZN(new_n4432_));
  NAND3_X1   g03426(.A1(new_n4411_), .A2(new_n4413_), .A3(new_n4409_), .ZN(new_n4433_));
  NAND3_X1   g03427(.A1(new_n4432_), .A2(new_n4433_), .A3(new_n4431_), .ZN(new_n4434_));
  NOR2_X1    g03428(.A1(new_n4410_), .A2(new_n4377_), .ZN(new_n4435_));
  NOR2_X1    g03429(.A1(new_n4385_), .A2(new_n4406_), .ZN(new_n4436_));
  NOR2_X1    g03430(.A1(new_n4436_), .A2(new_n4415_), .ZN(new_n4437_));
  AOI22_X1   g03431(.A1(new_n4353_), .A2(new_n4355_), .B1(new_n4360_), .B2(new_n4358_), .ZN(new_n4438_));
  NOR2_X1    g03432(.A1(new_n4438_), .A2(new_n4349_), .ZN(new_n4439_));
  NAND2_X1   g03433(.A1(new_n4329_), .A2(new_n4333_), .ZN(new_n4440_));
  NOR2_X1    g03434(.A1(new_n4361_), .A2(new_n4440_), .ZN(new_n4441_));
  NAND4_X1   g03435(.A1(new_n4437_), .A2(new_n4435_), .A3(new_n4439_), .A4(new_n4441_), .ZN(new_n4442_));
  NAND2_X1   g03436(.A1(new_n4434_), .A2(new_n4442_), .ZN(new_n4443_));
  AOI21_X1   g03437(.A1(new_n4428_), .A2(new_n4443_), .B(new_n4368_), .ZN(new_n4444_));
  NOR2_X1    g03438(.A1(new_n4419_), .A2(new_n4442_), .ZN(new_n4445_));
  NOR2_X1    g03439(.A1(new_n4418_), .A2(new_n4414_), .ZN(new_n4446_));
  NOR3_X1    g03440(.A1(new_n4423_), .A2(new_n4425_), .A3(new_n4421_), .ZN(new_n4447_));
  NAND2_X1   g03441(.A1(new_n4431_), .A2(new_n4441_), .ZN(new_n4448_));
  AOI21_X1   g03442(.A1(new_n4446_), .A2(new_n4447_), .B(new_n4448_), .ZN(new_n4449_));
  NOR3_X1    g03443(.A1(new_n4449_), .A2(new_n4445_), .A3(new_n4368_), .ZN(new_n4450_));
  NOR2_X1    g03444(.A1(new_n4450_), .A2(new_n4444_), .ZN(new_n4451_));
  AOI21_X1   g03445(.A1(new_n4365_), .A2(new_n4366_), .B(new_n4364_), .ZN(new_n4452_));
  NOR3_X1    g03446(.A1(new_n4362_), .A2(new_n4350_), .A3(new_n4329_), .ZN(new_n4453_));
  NOR2_X1    g03447(.A1(new_n4452_), .A2(new_n4453_), .ZN(new_n4454_));
  NOR2_X1    g03448(.A1(new_n4434_), .A2(new_n4442_), .ZN(new_n4455_));
  NOR2_X1    g03449(.A1(new_n4419_), .A2(new_n4427_), .ZN(new_n4456_));
  OAI21_X1   g03450(.A1(new_n4456_), .A2(new_n4455_), .B(new_n4454_), .ZN(new_n4457_));
  NAND2_X1   g03451(.A1(new_n4434_), .A2(new_n4427_), .ZN(new_n4458_));
  NAND2_X1   g03452(.A1(new_n4432_), .A2(new_n4433_), .ZN(new_n4459_));
  NAND3_X1   g03453(.A1(new_n4437_), .A2(new_n4435_), .A3(new_n4439_), .ZN(new_n4460_));
  NOR2_X1    g03454(.A1(new_n4408_), .A2(new_n4426_), .ZN(new_n4461_));
  OAI21_X1   g03455(.A1(new_n4459_), .A2(new_n4460_), .B(new_n4461_), .ZN(new_n4462_));
  NAND3_X1   g03456(.A1(new_n4462_), .A2(new_n4458_), .A3(new_n4454_), .ZN(new_n4463_));
  NOR2_X1    g03457(.A1(new_n4423_), .A2(new_n4421_), .ZN(new_n4464_));
  NAND2_X1   g03458(.A1(new_n4439_), .A2(new_n4441_), .ZN(new_n4465_));
  NOR2_X1    g03459(.A1(new_n4464_), .A2(new_n4465_), .ZN(new_n4466_));
  NAND2_X1   g03460(.A1(new_n4437_), .A2(new_n4435_), .ZN(new_n4467_));
  NOR2_X1    g03461(.A1(new_n4425_), .A2(new_n4426_), .ZN(new_n4468_));
  NOR2_X1    g03462(.A1(new_n4467_), .A2(new_n4468_), .ZN(new_n4469_));
  INV_X1     g03463(.I(\A[135] ), .ZN(new_n4470_));
  NOR2_X1    g03464(.A1(new_n4470_), .A2(\A[134] ), .ZN(new_n4471_));
  INV_X1     g03465(.I(\A[134] ), .ZN(new_n4472_));
  NOR2_X1    g03466(.A1(new_n4472_), .A2(\A[135] ), .ZN(new_n4473_));
  OAI21_X1   g03467(.A1(new_n4471_), .A2(new_n4473_), .B(\A[133] ), .ZN(new_n4474_));
  INV_X1     g03468(.I(\A[133] ), .ZN(new_n4475_));
  NOR2_X1    g03469(.A1(\A[134] ), .A2(\A[135] ), .ZN(new_n4476_));
  NAND2_X1   g03470(.A1(\A[134] ), .A2(\A[135] ), .ZN(new_n4477_));
  INV_X1     g03471(.I(new_n4477_), .ZN(new_n4478_));
  OAI21_X1   g03472(.A1(new_n4478_), .A2(new_n4476_), .B(new_n4475_), .ZN(new_n4479_));
  NAND2_X1   g03473(.A1(new_n4474_), .A2(new_n4479_), .ZN(new_n4480_));
  INV_X1     g03474(.I(\A[138] ), .ZN(new_n4481_));
  NOR2_X1    g03475(.A1(new_n4481_), .A2(\A[137] ), .ZN(new_n4482_));
  INV_X1     g03476(.I(\A[137] ), .ZN(new_n4483_));
  NOR2_X1    g03477(.A1(new_n4483_), .A2(\A[138] ), .ZN(new_n4484_));
  OAI21_X1   g03478(.A1(new_n4482_), .A2(new_n4484_), .B(\A[136] ), .ZN(new_n4485_));
  INV_X1     g03479(.I(\A[136] ), .ZN(new_n4486_));
  NOR2_X1    g03480(.A1(\A[137] ), .A2(\A[138] ), .ZN(new_n4487_));
  NAND2_X1   g03481(.A1(\A[137] ), .A2(\A[138] ), .ZN(new_n4488_));
  INV_X1     g03482(.I(new_n4488_), .ZN(new_n4489_));
  OAI21_X1   g03483(.A1(new_n4489_), .A2(new_n4487_), .B(new_n4486_), .ZN(new_n4490_));
  NAND2_X1   g03484(.A1(new_n4485_), .A2(new_n4490_), .ZN(new_n4491_));
  AOI21_X1   g03485(.A1(new_n4486_), .A2(new_n4488_), .B(new_n4487_), .ZN(new_n4492_));
  AOI21_X1   g03486(.A1(new_n4475_), .A2(new_n4477_), .B(new_n4476_), .ZN(new_n4493_));
  NAND2_X1   g03487(.A1(new_n4492_), .A2(new_n4493_), .ZN(new_n4494_));
  NOR3_X1    g03488(.A1(new_n4480_), .A2(new_n4491_), .A3(new_n4494_), .ZN(new_n4495_));
  NOR2_X1    g03489(.A1(new_n4480_), .A2(new_n4491_), .ZN(new_n4496_));
  NAND2_X1   g03490(.A1(new_n4472_), .A2(\A[135] ), .ZN(new_n4497_));
  NAND2_X1   g03491(.A1(new_n4470_), .A2(\A[134] ), .ZN(new_n4498_));
  AOI21_X1   g03492(.A1(new_n4497_), .A2(new_n4498_), .B(new_n4475_), .ZN(new_n4499_));
  INV_X1     g03493(.I(new_n4476_), .ZN(new_n4500_));
  AOI21_X1   g03494(.A1(new_n4500_), .A2(new_n4477_), .B(\A[133] ), .ZN(new_n4501_));
  NOR2_X1    g03495(.A1(new_n4501_), .A2(new_n4499_), .ZN(new_n4502_));
  NAND2_X1   g03496(.A1(new_n4483_), .A2(\A[138] ), .ZN(new_n4503_));
  NAND2_X1   g03497(.A1(new_n4481_), .A2(\A[137] ), .ZN(new_n4504_));
  AOI21_X1   g03498(.A1(new_n4503_), .A2(new_n4504_), .B(new_n4486_), .ZN(new_n4505_));
  INV_X1     g03499(.I(new_n4487_), .ZN(new_n4506_));
  AOI21_X1   g03500(.A1(new_n4506_), .A2(new_n4488_), .B(\A[136] ), .ZN(new_n4507_));
  NOR2_X1    g03501(.A1(new_n4507_), .A2(new_n4505_), .ZN(new_n4508_));
  NOR2_X1    g03502(.A1(new_n4502_), .A2(new_n4508_), .ZN(new_n4509_));
  NOR2_X1    g03503(.A1(new_n4509_), .A2(new_n4496_), .ZN(new_n4510_));
  INV_X1     g03504(.I(\A[127] ), .ZN(new_n4511_));
  INV_X1     g03505(.I(\A[128] ), .ZN(new_n4512_));
  NAND2_X1   g03506(.A1(new_n4512_), .A2(\A[129] ), .ZN(new_n4513_));
  INV_X1     g03507(.I(\A[129] ), .ZN(new_n4514_));
  NAND2_X1   g03508(.A1(new_n4514_), .A2(\A[128] ), .ZN(new_n4515_));
  AOI21_X1   g03509(.A1(new_n4513_), .A2(new_n4515_), .B(new_n4511_), .ZN(new_n4516_));
  NOR2_X1    g03510(.A1(\A[128] ), .A2(\A[129] ), .ZN(new_n4517_));
  INV_X1     g03511(.I(new_n4517_), .ZN(new_n4518_));
  NAND2_X1   g03512(.A1(\A[128] ), .A2(\A[129] ), .ZN(new_n4519_));
  AOI21_X1   g03513(.A1(new_n4518_), .A2(new_n4519_), .B(\A[127] ), .ZN(new_n4520_));
  NOR2_X1    g03514(.A1(new_n4520_), .A2(new_n4516_), .ZN(new_n4521_));
  INV_X1     g03515(.I(\A[130] ), .ZN(new_n4522_));
  INV_X1     g03516(.I(\A[131] ), .ZN(new_n4523_));
  NAND2_X1   g03517(.A1(new_n4523_), .A2(\A[132] ), .ZN(new_n4524_));
  INV_X1     g03518(.I(\A[132] ), .ZN(new_n4525_));
  NAND2_X1   g03519(.A1(new_n4525_), .A2(\A[131] ), .ZN(new_n4526_));
  AOI21_X1   g03520(.A1(new_n4524_), .A2(new_n4526_), .B(new_n4522_), .ZN(new_n4527_));
  NOR2_X1    g03521(.A1(\A[131] ), .A2(\A[132] ), .ZN(new_n4528_));
  INV_X1     g03522(.I(new_n4528_), .ZN(new_n4529_));
  NAND2_X1   g03523(.A1(\A[131] ), .A2(\A[132] ), .ZN(new_n4530_));
  AOI21_X1   g03524(.A1(new_n4529_), .A2(new_n4530_), .B(\A[130] ), .ZN(new_n4531_));
  NOR2_X1    g03525(.A1(new_n4531_), .A2(new_n4527_), .ZN(new_n4532_));
  AOI21_X1   g03526(.A1(new_n4522_), .A2(new_n4530_), .B(new_n4528_), .ZN(new_n4533_));
  AOI21_X1   g03527(.A1(new_n4511_), .A2(new_n4519_), .B(new_n4517_), .ZN(new_n4534_));
  NAND2_X1   g03528(.A1(new_n4533_), .A2(new_n4534_), .ZN(new_n4535_));
  NAND2_X1   g03529(.A1(new_n4510_), .A2(new_n4495_), .ZN(new_n4537_));
  INV_X1     g03530(.I(new_n4537_), .ZN(new_n4538_));
  NOR3_X1    g03531(.A1(new_n4469_), .A2(new_n4466_), .A3(new_n4538_), .ZN(new_n4539_));
  AOI21_X1   g03532(.A1(new_n4457_), .A2(new_n4463_), .B(new_n4539_), .ZN(new_n4540_));
  NOR2_X1    g03533(.A1(new_n4469_), .A2(new_n4466_), .ZN(new_n4541_));
  NAND2_X1   g03534(.A1(new_n4541_), .A2(new_n4537_), .ZN(new_n4542_));
  NOR3_X1    g03535(.A1(new_n4450_), .A2(new_n4444_), .A3(new_n4542_), .ZN(new_n4543_));
  INV_X1     g03536(.I(new_n4493_), .ZN(new_n4544_));
  AOI21_X1   g03537(.A1(new_n4502_), .A2(new_n4508_), .B(new_n4544_), .ZN(new_n4545_));
  NOR3_X1    g03538(.A1(new_n4480_), .A2(new_n4491_), .A3(new_n4493_), .ZN(new_n4546_));
  OAI21_X1   g03539(.A1(new_n4545_), .A2(new_n4546_), .B(new_n4492_), .ZN(new_n4547_));
  INV_X1     g03540(.I(new_n4492_), .ZN(new_n4548_));
  OAI21_X1   g03541(.A1(new_n4480_), .A2(new_n4491_), .B(new_n4493_), .ZN(new_n4549_));
  NAND3_X1   g03542(.A1(new_n4502_), .A2(new_n4508_), .A3(new_n4544_), .ZN(new_n4550_));
  NAND3_X1   g03543(.A1(new_n4549_), .A2(new_n4550_), .A3(new_n4548_), .ZN(new_n4551_));
  NAND2_X1   g03544(.A1(new_n4547_), .A2(new_n4551_), .ZN(new_n4552_));
  NOR4_X1    g03545(.A1(new_n4516_), .A2(new_n4520_), .A3(new_n4531_), .A4(new_n4527_), .ZN(new_n4553_));
  NOR2_X1    g03546(.A1(new_n4521_), .A2(new_n4532_), .ZN(new_n4554_));
  NOR2_X1    g03547(.A1(new_n4554_), .A2(new_n4553_), .ZN(new_n4555_));
  NAND3_X1   g03548(.A1(new_n4510_), .A2(new_n4555_), .A3(new_n4495_), .ZN(new_n4556_));
  NAND2_X1   g03549(.A1(new_n4521_), .A2(new_n4532_), .ZN(new_n4557_));
  NAND2_X1   g03550(.A1(new_n4502_), .A2(new_n4491_), .ZN(new_n4558_));
  NAND2_X1   g03551(.A1(new_n4508_), .A2(new_n4480_), .ZN(new_n4559_));
  AOI21_X1   g03552(.A1(new_n4558_), .A2(new_n4559_), .B(new_n4494_), .ZN(new_n4560_));
  NOR3_X1    g03553(.A1(new_n4560_), .A2(new_n4557_), .A3(new_n4535_), .ZN(new_n4561_));
  OAI21_X1   g03554(.A1(new_n4552_), .A2(new_n4556_), .B(new_n4561_), .ZN(new_n4562_));
  INV_X1     g03555(.I(new_n4533_), .ZN(new_n4563_));
  NOR2_X1    g03556(.A1(new_n4514_), .A2(\A[128] ), .ZN(new_n4564_));
  NOR2_X1    g03557(.A1(new_n4512_), .A2(\A[129] ), .ZN(new_n4565_));
  OAI21_X1   g03558(.A1(new_n4564_), .A2(new_n4565_), .B(\A[127] ), .ZN(new_n4566_));
  INV_X1     g03559(.I(new_n4519_), .ZN(new_n4567_));
  OAI21_X1   g03560(.A1(new_n4567_), .A2(new_n4517_), .B(new_n4511_), .ZN(new_n4568_));
  NAND2_X1   g03561(.A1(new_n4566_), .A2(new_n4568_), .ZN(new_n4569_));
  NOR2_X1    g03562(.A1(new_n4525_), .A2(\A[131] ), .ZN(new_n4570_));
  NOR2_X1    g03563(.A1(new_n4523_), .A2(\A[132] ), .ZN(new_n4571_));
  OAI21_X1   g03564(.A1(new_n4570_), .A2(new_n4571_), .B(\A[130] ), .ZN(new_n4572_));
  INV_X1     g03565(.I(new_n4530_), .ZN(new_n4573_));
  OAI21_X1   g03566(.A1(new_n4573_), .A2(new_n4528_), .B(new_n4522_), .ZN(new_n4574_));
  NAND2_X1   g03567(.A1(new_n4572_), .A2(new_n4574_), .ZN(new_n4575_));
  OAI21_X1   g03568(.A1(new_n4569_), .A2(new_n4575_), .B(new_n4534_), .ZN(new_n4576_));
  INV_X1     g03569(.I(new_n4534_), .ZN(new_n4577_));
  NAND3_X1   g03570(.A1(new_n4521_), .A2(new_n4532_), .A3(new_n4577_), .ZN(new_n4578_));
  AOI21_X1   g03571(.A1(new_n4576_), .A2(new_n4578_), .B(new_n4563_), .ZN(new_n4579_));
  NOR2_X1    g03572(.A1(new_n4553_), .A2(new_n4577_), .ZN(new_n4580_));
  NOR3_X1    g03573(.A1(new_n4569_), .A2(new_n4575_), .A3(new_n4534_), .ZN(new_n4581_));
  NOR3_X1    g03574(.A1(new_n4580_), .A2(new_n4581_), .A3(new_n4533_), .ZN(new_n4582_));
  NOR2_X1    g03575(.A1(new_n4582_), .A2(new_n4579_), .ZN(new_n4583_));
  NOR2_X1    g03576(.A1(new_n4562_), .A2(new_n4583_), .ZN(new_n4584_));
  OAI21_X1   g03577(.A1(new_n4580_), .A2(new_n4581_), .B(new_n4533_), .ZN(new_n4585_));
  NAND3_X1   g03578(.A1(new_n4576_), .A2(new_n4578_), .A3(new_n4563_), .ZN(new_n4586_));
  NAND2_X1   g03579(.A1(new_n4585_), .A2(new_n4586_), .ZN(new_n4587_));
  NOR3_X1    g03580(.A1(new_n4569_), .A2(new_n4575_), .A3(new_n4535_), .ZN(new_n4588_));
  NAND4_X1   g03581(.A1(new_n4510_), .A2(new_n4555_), .A3(new_n4495_), .A4(new_n4588_), .ZN(new_n4589_));
  NAND2_X1   g03582(.A1(new_n4587_), .A2(new_n4589_), .ZN(new_n4590_));
  INV_X1     g03583(.I(new_n4494_), .ZN(new_n4591_));
  NOR2_X1    g03584(.A1(new_n4508_), .A2(new_n4480_), .ZN(new_n4592_));
  NOR2_X1    g03585(.A1(new_n4502_), .A2(new_n4491_), .ZN(new_n4593_));
  OAI21_X1   g03586(.A1(new_n4592_), .A2(new_n4593_), .B(new_n4591_), .ZN(new_n4594_));
  NAND3_X1   g03587(.A1(new_n4547_), .A2(new_n4551_), .A3(new_n4594_), .ZN(new_n4595_));
  OAI21_X1   g03588(.A1(new_n4587_), .A2(new_n4589_), .B(new_n4595_), .ZN(new_n4596_));
  NAND2_X1   g03589(.A1(new_n4502_), .A2(new_n4508_), .ZN(new_n4597_));
  NAND2_X1   g03590(.A1(new_n4480_), .A2(new_n4491_), .ZN(new_n4598_));
  NAND3_X1   g03591(.A1(new_n4495_), .A2(new_n4597_), .A3(new_n4598_), .ZN(new_n4599_));
  NAND2_X1   g03592(.A1(new_n4569_), .A2(new_n4575_), .ZN(new_n4600_));
  NAND3_X1   g03593(.A1(new_n4588_), .A2(new_n4557_), .A3(new_n4600_), .ZN(new_n4601_));
  NOR2_X1    g03594(.A1(new_n4599_), .A2(new_n4601_), .ZN(new_n4602_));
  AOI21_X1   g03595(.A1(new_n4549_), .A2(new_n4550_), .B(new_n4548_), .ZN(new_n4603_));
  NOR3_X1    g03596(.A1(new_n4545_), .A2(new_n4546_), .A3(new_n4492_), .ZN(new_n4604_));
  NOR3_X1    g03597(.A1(new_n4604_), .A2(new_n4603_), .A3(new_n4560_), .ZN(new_n4605_));
  NAND3_X1   g03598(.A1(new_n4605_), .A2(new_n4583_), .A3(new_n4602_), .ZN(new_n4606_));
  NAND2_X1   g03599(.A1(new_n4596_), .A2(new_n4606_), .ZN(new_n4607_));
  AOI21_X1   g03600(.A1(new_n4607_), .A2(new_n4590_), .B(new_n4584_), .ZN(new_n4608_));
  OAI22_X1   g03601(.A1(new_n4540_), .A2(new_n4543_), .B1(new_n4608_), .B2(new_n4451_), .ZN(new_n4609_));
  OAI21_X1   g03602(.A1(new_n4419_), .A2(new_n4442_), .B(new_n4368_), .ZN(new_n4610_));
  NAND2_X1   g03603(.A1(new_n4409_), .A2(new_n4412_), .ZN(new_n4611_));
  AOI21_X1   g03604(.A1(new_n4415_), .A2(new_n4611_), .B(new_n4420_), .ZN(new_n4612_));
  NOR2_X1    g03605(.A1(new_n4329_), .A2(new_n4333_), .ZN(new_n4613_));
  OAI21_X1   g03606(.A1(new_n4361_), .A2(new_n4613_), .B(new_n4440_), .ZN(new_n4614_));
  XOR2_X1    g03607(.A1(new_n4614_), .A2(new_n4612_), .Z(new_n4615_));
  NAND3_X1   g03608(.A1(new_n4610_), .A2(new_n4462_), .A3(new_n4615_), .ZN(new_n4616_));
  NOR2_X1    g03609(.A1(new_n4604_), .A2(new_n4603_), .ZN(new_n4617_));
  NOR3_X1    g03610(.A1(new_n4599_), .A2(new_n4553_), .A3(new_n4554_), .ZN(new_n4618_));
  NAND2_X1   g03611(.A1(new_n4594_), .A2(new_n4588_), .ZN(new_n4619_));
  AOI21_X1   g03612(.A1(new_n4617_), .A2(new_n4618_), .B(new_n4619_), .ZN(new_n4620_));
  AOI21_X1   g03613(.A1(new_n4595_), .A2(new_n4602_), .B(new_n4583_), .ZN(new_n4621_));
  NOR2_X1    g03614(.A1(new_n4492_), .A2(new_n4493_), .ZN(new_n4622_));
  OAI21_X1   g03615(.A1(new_n4597_), .A2(new_n4622_), .B(new_n4494_), .ZN(new_n4623_));
  NOR2_X1    g03616(.A1(new_n4533_), .A2(new_n4534_), .ZN(new_n4624_));
  OAI21_X1   g03617(.A1(new_n4557_), .A2(new_n4624_), .B(new_n4535_), .ZN(new_n4625_));
  XOR2_X1    g03618(.A1(new_n4623_), .A2(new_n4625_), .Z(new_n4626_));
  NOR3_X1    g03619(.A1(new_n4621_), .A2(new_n4620_), .A3(new_n4626_), .ZN(new_n4627_));
  XOR2_X1    g03620(.A1(new_n4616_), .A2(new_n4627_), .Z(new_n4628_));
  NOR2_X1    g03621(.A1(new_n4609_), .A2(new_n4628_), .ZN(new_n4629_));
  NAND2_X1   g03622(.A1(new_n4457_), .A2(new_n4463_), .ZN(new_n4630_));
  OAI21_X1   g03623(.A1(new_n4450_), .A2(new_n4444_), .B(new_n4542_), .ZN(new_n4631_));
  NAND3_X1   g03624(.A1(new_n4457_), .A2(new_n4463_), .A3(new_n4539_), .ZN(new_n4632_));
  NAND2_X1   g03625(.A1(new_n4620_), .A2(new_n4587_), .ZN(new_n4633_));
  NOR4_X1    g03626(.A1(new_n4599_), .A2(new_n4582_), .A3(new_n4579_), .A4(new_n4601_), .ZN(new_n4634_));
  NOR2_X1    g03627(.A1(new_n4634_), .A2(new_n4605_), .ZN(new_n4635_));
  NOR3_X1    g03628(.A1(new_n4595_), .A2(new_n4587_), .A3(new_n4589_), .ZN(new_n4636_));
  OAI21_X1   g03629(.A1(new_n4635_), .A2(new_n4636_), .B(new_n4590_), .ZN(new_n4637_));
  NAND2_X1   g03630(.A1(new_n4637_), .A2(new_n4633_), .ZN(new_n4638_));
  AOI22_X1   g03631(.A1(new_n4631_), .A2(new_n4632_), .B1(new_n4638_), .B2(new_n4630_), .ZN(new_n4639_));
  AOI21_X1   g03632(.A1(new_n4434_), .A2(new_n4427_), .B(new_n4454_), .ZN(new_n4640_));
  INV_X1     g03633(.I(new_n4615_), .ZN(new_n4641_));
  NOR3_X1    g03634(.A1(new_n4640_), .A2(new_n4449_), .A3(new_n4641_), .ZN(new_n4642_));
  NOR2_X1    g03635(.A1(new_n4642_), .A2(new_n4627_), .ZN(new_n4643_));
  OAI21_X1   g03636(.A1(new_n4605_), .A2(new_n4589_), .B(new_n4587_), .ZN(new_n4644_));
  XNOR2_X1   g03637(.A1(new_n4623_), .A2(new_n4625_), .ZN(new_n4645_));
  NAND3_X1   g03638(.A1(new_n4562_), .A2(new_n4644_), .A3(new_n4645_), .ZN(new_n4646_));
  NOR2_X1    g03639(.A1(new_n4616_), .A2(new_n4646_), .ZN(new_n4647_));
  NOR2_X1    g03640(.A1(new_n4643_), .A2(new_n4647_), .ZN(new_n4648_));
  NOR2_X1    g03641(.A1(new_n4639_), .A2(new_n4648_), .ZN(new_n4649_));
  INV_X1     g03642(.I(\A[166] ), .ZN(new_n4650_));
  NOR2_X1    g03643(.A1(\A[167] ), .A2(\A[168] ), .ZN(new_n4651_));
  NAND2_X1   g03644(.A1(\A[167] ), .A2(\A[168] ), .ZN(new_n4652_));
  AOI21_X1   g03645(.A1(new_n4650_), .A2(new_n4652_), .B(new_n4651_), .ZN(new_n4653_));
  INV_X1     g03646(.I(\A[163] ), .ZN(new_n4654_));
  NOR2_X1    g03647(.A1(\A[164] ), .A2(\A[165] ), .ZN(new_n4655_));
  NAND2_X1   g03648(.A1(\A[164] ), .A2(\A[165] ), .ZN(new_n4656_));
  AOI21_X1   g03649(.A1(new_n4654_), .A2(new_n4656_), .B(new_n4655_), .ZN(new_n4657_));
  INV_X1     g03650(.I(new_n4657_), .ZN(new_n4658_));
  INV_X1     g03651(.I(\A[164] ), .ZN(new_n4659_));
  NAND2_X1   g03652(.A1(new_n4659_), .A2(\A[165] ), .ZN(new_n4660_));
  INV_X1     g03653(.I(\A[165] ), .ZN(new_n4661_));
  NAND2_X1   g03654(.A1(new_n4661_), .A2(\A[164] ), .ZN(new_n4662_));
  AOI21_X1   g03655(.A1(new_n4660_), .A2(new_n4662_), .B(new_n4654_), .ZN(new_n4663_));
  INV_X1     g03656(.I(new_n4655_), .ZN(new_n4664_));
  AOI21_X1   g03657(.A1(new_n4664_), .A2(new_n4656_), .B(\A[163] ), .ZN(new_n4665_));
  INV_X1     g03658(.I(\A[167] ), .ZN(new_n4666_));
  NAND2_X1   g03659(.A1(new_n4666_), .A2(\A[168] ), .ZN(new_n4667_));
  INV_X1     g03660(.I(\A[168] ), .ZN(new_n4668_));
  NAND2_X1   g03661(.A1(new_n4668_), .A2(\A[167] ), .ZN(new_n4669_));
  AOI21_X1   g03662(.A1(new_n4667_), .A2(new_n4669_), .B(new_n4650_), .ZN(new_n4670_));
  INV_X1     g03663(.I(new_n4651_), .ZN(new_n4671_));
  AOI21_X1   g03664(.A1(new_n4671_), .A2(new_n4652_), .B(\A[166] ), .ZN(new_n4672_));
  NOR4_X1    g03665(.A1(new_n4663_), .A2(new_n4665_), .A3(new_n4672_), .A4(new_n4670_), .ZN(new_n4673_));
  NOR2_X1    g03666(.A1(new_n4673_), .A2(new_n4658_), .ZN(new_n4674_));
  NOR2_X1    g03667(.A1(new_n4661_), .A2(\A[164] ), .ZN(new_n4675_));
  NOR2_X1    g03668(.A1(new_n4659_), .A2(\A[165] ), .ZN(new_n4676_));
  OAI21_X1   g03669(.A1(new_n4675_), .A2(new_n4676_), .B(\A[163] ), .ZN(new_n4677_));
  INV_X1     g03670(.I(new_n4656_), .ZN(new_n4678_));
  OAI21_X1   g03671(.A1(new_n4678_), .A2(new_n4655_), .B(new_n4654_), .ZN(new_n4679_));
  NOR2_X1    g03672(.A1(new_n4668_), .A2(\A[167] ), .ZN(new_n4680_));
  NOR2_X1    g03673(.A1(new_n4666_), .A2(\A[168] ), .ZN(new_n4681_));
  OAI21_X1   g03674(.A1(new_n4680_), .A2(new_n4681_), .B(\A[166] ), .ZN(new_n4682_));
  INV_X1     g03675(.I(new_n4652_), .ZN(new_n4683_));
  OAI21_X1   g03676(.A1(new_n4683_), .A2(new_n4651_), .B(new_n4650_), .ZN(new_n4684_));
  NAND4_X1   g03677(.A1(new_n4677_), .A2(new_n4679_), .A3(new_n4682_), .A4(new_n4684_), .ZN(new_n4685_));
  NOR2_X1    g03678(.A1(new_n4685_), .A2(new_n4657_), .ZN(new_n4686_));
  OAI21_X1   g03679(.A1(new_n4674_), .A2(new_n4686_), .B(new_n4653_), .ZN(new_n4687_));
  INV_X1     g03680(.I(new_n4653_), .ZN(new_n4688_));
  NAND2_X1   g03681(.A1(new_n4685_), .A2(new_n4657_), .ZN(new_n4689_));
  NAND2_X1   g03682(.A1(new_n4673_), .A2(new_n4658_), .ZN(new_n4690_));
  NAND3_X1   g03683(.A1(new_n4690_), .A2(new_n4689_), .A3(new_n4688_), .ZN(new_n4691_));
  NAND2_X1   g03684(.A1(new_n4687_), .A2(new_n4691_), .ZN(new_n4692_));
  INV_X1     g03685(.I(\A[172] ), .ZN(new_n4693_));
  NOR2_X1    g03686(.A1(\A[173] ), .A2(\A[174] ), .ZN(new_n4694_));
  NAND2_X1   g03687(.A1(\A[173] ), .A2(\A[174] ), .ZN(new_n4695_));
  AOI21_X1   g03688(.A1(new_n4693_), .A2(new_n4695_), .B(new_n4694_), .ZN(new_n4696_));
  INV_X1     g03689(.I(\A[169] ), .ZN(new_n4697_));
  NOR2_X1    g03690(.A1(\A[170] ), .A2(\A[171] ), .ZN(new_n4698_));
  NAND2_X1   g03691(.A1(\A[170] ), .A2(\A[171] ), .ZN(new_n4699_));
  AOI21_X1   g03692(.A1(new_n4697_), .A2(new_n4699_), .B(new_n4698_), .ZN(new_n4700_));
  NAND2_X1   g03693(.A1(new_n4696_), .A2(new_n4700_), .ZN(new_n4701_));
  INV_X1     g03694(.I(\A[170] ), .ZN(new_n4702_));
  NAND2_X1   g03695(.A1(new_n4702_), .A2(\A[171] ), .ZN(new_n4703_));
  INV_X1     g03696(.I(\A[171] ), .ZN(new_n4704_));
  NAND2_X1   g03697(.A1(new_n4704_), .A2(\A[170] ), .ZN(new_n4705_));
  AOI21_X1   g03698(.A1(new_n4703_), .A2(new_n4705_), .B(new_n4697_), .ZN(new_n4706_));
  INV_X1     g03699(.I(new_n4698_), .ZN(new_n4707_));
  AOI21_X1   g03700(.A1(new_n4707_), .A2(new_n4699_), .B(\A[169] ), .ZN(new_n4708_));
  NOR2_X1    g03701(.A1(new_n4708_), .A2(new_n4706_), .ZN(new_n4709_));
  INV_X1     g03702(.I(\A[174] ), .ZN(new_n4710_));
  NOR2_X1    g03703(.A1(new_n4710_), .A2(\A[173] ), .ZN(new_n4711_));
  INV_X1     g03704(.I(\A[173] ), .ZN(new_n4712_));
  NOR2_X1    g03705(.A1(new_n4712_), .A2(\A[174] ), .ZN(new_n4713_));
  OAI21_X1   g03706(.A1(new_n4711_), .A2(new_n4713_), .B(\A[172] ), .ZN(new_n4714_));
  AND2_X2    g03707(.A1(\A[173] ), .A2(\A[174] ), .Z(new_n4715_));
  OAI21_X1   g03708(.A1(new_n4715_), .A2(new_n4694_), .B(new_n4693_), .ZN(new_n4716_));
  NAND2_X1   g03709(.A1(new_n4714_), .A2(new_n4716_), .ZN(new_n4717_));
  NAND2_X1   g03710(.A1(new_n4709_), .A2(new_n4717_), .ZN(new_n4718_));
  NOR2_X1    g03711(.A1(new_n4704_), .A2(\A[170] ), .ZN(new_n4719_));
  NOR2_X1    g03712(.A1(new_n4702_), .A2(\A[171] ), .ZN(new_n4720_));
  OAI21_X1   g03713(.A1(new_n4719_), .A2(new_n4720_), .B(\A[169] ), .ZN(new_n4721_));
  AND2_X2    g03714(.A1(\A[170] ), .A2(\A[171] ), .Z(new_n4722_));
  OAI21_X1   g03715(.A1(new_n4722_), .A2(new_n4698_), .B(new_n4697_), .ZN(new_n4723_));
  NAND2_X1   g03716(.A1(new_n4721_), .A2(new_n4723_), .ZN(new_n4724_));
  NAND2_X1   g03717(.A1(new_n4712_), .A2(\A[174] ), .ZN(new_n4725_));
  NAND2_X1   g03718(.A1(new_n4710_), .A2(\A[173] ), .ZN(new_n4726_));
  AOI21_X1   g03719(.A1(new_n4725_), .A2(new_n4726_), .B(new_n4693_), .ZN(new_n4727_));
  INV_X1     g03720(.I(new_n4694_), .ZN(new_n4728_));
  AOI21_X1   g03721(.A1(new_n4728_), .A2(new_n4695_), .B(\A[172] ), .ZN(new_n4729_));
  NOR2_X1    g03722(.A1(new_n4729_), .A2(new_n4727_), .ZN(new_n4730_));
  NAND2_X1   g03723(.A1(new_n4730_), .A2(new_n4724_), .ZN(new_n4731_));
  AOI21_X1   g03724(.A1(new_n4718_), .A2(new_n4731_), .B(new_n4701_), .ZN(new_n4732_));
  INV_X1     g03725(.I(new_n4696_), .ZN(new_n4733_));
  NAND4_X1   g03726(.A1(new_n4721_), .A2(new_n4714_), .A3(new_n4723_), .A4(new_n4716_), .ZN(new_n4734_));
  NAND2_X1   g03727(.A1(new_n4734_), .A2(new_n4700_), .ZN(new_n4735_));
  INV_X1     g03728(.I(new_n4700_), .ZN(new_n4736_));
  NAND3_X1   g03729(.A1(new_n4709_), .A2(new_n4730_), .A3(new_n4736_), .ZN(new_n4737_));
  AOI21_X1   g03730(.A1(new_n4735_), .A2(new_n4737_), .B(new_n4733_), .ZN(new_n4738_));
  AOI21_X1   g03731(.A1(new_n4709_), .A2(new_n4730_), .B(new_n4736_), .ZN(new_n4739_));
  NOR3_X1    g03732(.A1(new_n4724_), .A2(new_n4717_), .A3(new_n4700_), .ZN(new_n4740_));
  NOR3_X1    g03733(.A1(new_n4739_), .A2(new_n4740_), .A3(new_n4696_), .ZN(new_n4741_));
  NOR3_X1    g03734(.A1(new_n4738_), .A2(new_n4741_), .A3(new_n4732_), .ZN(new_n4742_));
  INV_X1     g03735(.I(new_n4701_), .ZN(new_n4743_));
  NOR4_X1    g03736(.A1(new_n4706_), .A2(new_n4708_), .A3(new_n4729_), .A4(new_n4727_), .ZN(new_n4744_));
  NAND2_X1   g03737(.A1(new_n4744_), .A2(new_n4743_), .ZN(new_n4745_));
  NAND2_X1   g03738(.A1(new_n4724_), .A2(new_n4717_), .ZN(new_n4746_));
  NAND2_X1   g03739(.A1(new_n4746_), .A2(new_n4734_), .ZN(new_n4747_));
  OAI22_X1   g03740(.A1(new_n4663_), .A2(new_n4665_), .B1(new_n4672_), .B2(new_n4670_), .ZN(new_n4748_));
  NAND2_X1   g03741(.A1(new_n4748_), .A2(new_n4685_), .ZN(new_n4749_));
  NAND2_X1   g03742(.A1(new_n4653_), .A2(new_n4657_), .ZN(new_n4750_));
  INV_X1     g03743(.I(new_n4750_), .ZN(new_n4751_));
  NAND2_X1   g03744(.A1(new_n4673_), .A2(new_n4751_), .ZN(new_n4752_));
  NOR4_X1    g03745(.A1(new_n4747_), .A2(new_n4749_), .A3(new_n4745_), .A4(new_n4752_), .ZN(new_n4753_));
  NAND2_X1   g03746(.A1(new_n4742_), .A2(new_n4753_), .ZN(new_n4754_));
  NOR2_X1    g03747(.A1(new_n4730_), .A2(new_n4724_), .ZN(new_n4755_));
  NOR2_X1    g03748(.A1(new_n4709_), .A2(new_n4717_), .ZN(new_n4756_));
  OAI21_X1   g03749(.A1(new_n4755_), .A2(new_n4756_), .B(new_n4743_), .ZN(new_n4757_));
  OAI21_X1   g03750(.A1(new_n4739_), .A2(new_n4740_), .B(new_n4696_), .ZN(new_n4758_));
  NAND3_X1   g03751(.A1(new_n4735_), .A2(new_n4737_), .A3(new_n4733_), .ZN(new_n4759_));
  NAND3_X1   g03752(.A1(new_n4759_), .A2(new_n4758_), .A3(new_n4757_), .ZN(new_n4760_));
  NOR2_X1    g03753(.A1(new_n4734_), .A2(new_n4701_), .ZN(new_n4761_));
  AOI22_X1   g03754(.A1(new_n4721_), .A2(new_n4723_), .B1(new_n4714_), .B2(new_n4716_), .ZN(new_n4762_));
  NOR2_X1    g03755(.A1(new_n4744_), .A2(new_n4762_), .ZN(new_n4763_));
  AOI22_X1   g03756(.A1(new_n4677_), .A2(new_n4679_), .B1(new_n4682_), .B2(new_n4684_), .ZN(new_n4764_));
  NOR2_X1    g03757(.A1(new_n4764_), .A2(new_n4673_), .ZN(new_n4765_));
  NOR2_X1    g03758(.A1(new_n4685_), .A2(new_n4750_), .ZN(new_n4766_));
  NAND4_X1   g03759(.A1(new_n4765_), .A2(new_n4763_), .A3(new_n4766_), .A4(new_n4761_), .ZN(new_n4767_));
  NAND2_X1   g03760(.A1(new_n4760_), .A2(new_n4767_), .ZN(new_n4768_));
  AOI21_X1   g03761(.A1(new_n4754_), .A2(new_n4768_), .B(new_n4692_), .ZN(new_n4769_));
  NOR2_X1    g03762(.A1(new_n4742_), .A2(new_n4767_), .ZN(new_n4770_));
  NOR2_X1    g03763(.A1(new_n4738_), .A2(new_n4741_), .ZN(new_n4771_));
  NAND3_X1   g03764(.A1(new_n4765_), .A2(new_n4763_), .A3(new_n4761_), .ZN(new_n4772_));
  INV_X1     g03765(.I(new_n4772_), .ZN(new_n4773_));
  NAND2_X1   g03766(.A1(new_n4757_), .A2(new_n4766_), .ZN(new_n4774_));
  AOI21_X1   g03767(.A1(new_n4773_), .A2(new_n4771_), .B(new_n4774_), .ZN(new_n4775_));
  NOR3_X1    g03768(.A1(new_n4775_), .A2(new_n4770_), .A3(new_n4692_), .ZN(new_n4776_));
  NOR2_X1    g03769(.A1(new_n4776_), .A2(new_n4769_), .ZN(new_n4777_));
  AOI21_X1   g03770(.A1(new_n4690_), .A2(new_n4689_), .B(new_n4688_), .ZN(new_n4778_));
  NOR3_X1    g03771(.A1(new_n4674_), .A2(new_n4686_), .A3(new_n4653_), .ZN(new_n4779_));
  NOR2_X1    g03772(.A1(new_n4778_), .A2(new_n4779_), .ZN(new_n4780_));
  NOR4_X1    g03773(.A1(new_n4767_), .A2(new_n4732_), .A3(new_n4738_), .A4(new_n4741_), .ZN(new_n4781_));
  NOR2_X1    g03774(.A1(new_n4742_), .A2(new_n4753_), .ZN(new_n4782_));
  OAI21_X1   g03775(.A1(new_n4782_), .A2(new_n4781_), .B(new_n4780_), .ZN(new_n4783_));
  NAND2_X1   g03776(.A1(new_n4760_), .A2(new_n4753_), .ZN(new_n4784_));
  NAND2_X1   g03777(.A1(new_n4759_), .A2(new_n4758_), .ZN(new_n4785_));
  NOR2_X1    g03778(.A1(new_n4732_), .A2(new_n4752_), .ZN(new_n4786_));
  OAI21_X1   g03779(.A1(new_n4785_), .A2(new_n4772_), .B(new_n4786_), .ZN(new_n4787_));
  NAND3_X1   g03780(.A1(new_n4787_), .A2(new_n4784_), .A3(new_n4780_), .ZN(new_n4788_));
  NOR2_X1    g03781(.A1(new_n4747_), .A2(new_n4745_), .ZN(new_n4789_));
  NAND2_X1   g03782(.A1(new_n4765_), .A2(new_n4766_), .ZN(new_n4790_));
  NOR2_X1    g03783(.A1(new_n4789_), .A2(new_n4790_), .ZN(new_n4791_));
  NAND2_X1   g03784(.A1(new_n4789_), .A2(new_n4790_), .ZN(new_n4792_));
  INV_X1     g03785(.I(new_n4792_), .ZN(new_n4793_));
  INV_X1     g03786(.I(\A[159] ), .ZN(new_n4794_));
  NOR2_X1    g03787(.A1(new_n4794_), .A2(\A[158] ), .ZN(new_n4795_));
  INV_X1     g03788(.I(\A[158] ), .ZN(new_n4796_));
  NOR2_X1    g03789(.A1(new_n4796_), .A2(\A[159] ), .ZN(new_n4797_));
  OAI21_X1   g03790(.A1(new_n4795_), .A2(new_n4797_), .B(\A[157] ), .ZN(new_n4798_));
  INV_X1     g03791(.I(\A[157] ), .ZN(new_n4799_));
  NOR2_X1    g03792(.A1(\A[158] ), .A2(\A[159] ), .ZN(new_n4800_));
  NAND2_X1   g03793(.A1(\A[158] ), .A2(\A[159] ), .ZN(new_n4801_));
  INV_X1     g03794(.I(new_n4801_), .ZN(new_n4802_));
  OAI21_X1   g03795(.A1(new_n4802_), .A2(new_n4800_), .B(new_n4799_), .ZN(new_n4803_));
  NAND2_X1   g03796(.A1(new_n4798_), .A2(new_n4803_), .ZN(new_n4804_));
  INV_X1     g03797(.I(\A[162] ), .ZN(new_n4805_));
  NOR2_X1    g03798(.A1(new_n4805_), .A2(\A[161] ), .ZN(new_n4806_));
  INV_X1     g03799(.I(\A[161] ), .ZN(new_n4807_));
  NOR2_X1    g03800(.A1(new_n4807_), .A2(\A[162] ), .ZN(new_n4808_));
  OAI21_X1   g03801(.A1(new_n4806_), .A2(new_n4808_), .B(\A[160] ), .ZN(new_n4809_));
  INV_X1     g03802(.I(\A[160] ), .ZN(new_n4810_));
  NOR2_X1    g03803(.A1(\A[161] ), .A2(\A[162] ), .ZN(new_n4811_));
  AND2_X2    g03804(.A1(\A[161] ), .A2(\A[162] ), .Z(new_n4812_));
  OAI21_X1   g03805(.A1(new_n4812_), .A2(new_n4811_), .B(new_n4810_), .ZN(new_n4813_));
  NAND2_X1   g03806(.A1(new_n4809_), .A2(new_n4813_), .ZN(new_n4814_));
  NAND2_X1   g03807(.A1(\A[161] ), .A2(\A[162] ), .ZN(new_n4815_));
  AOI21_X1   g03808(.A1(new_n4810_), .A2(new_n4815_), .B(new_n4811_), .ZN(new_n4816_));
  AOI21_X1   g03809(.A1(new_n4799_), .A2(new_n4801_), .B(new_n4800_), .ZN(new_n4817_));
  NAND2_X1   g03810(.A1(new_n4816_), .A2(new_n4817_), .ZN(new_n4818_));
  NOR3_X1    g03811(.A1(new_n4804_), .A2(new_n4814_), .A3(new_n4818_), .ZN(new_n4819_));
  NOR2_X1    g03812(.A1(new_n4804_), .A2(new_n4814_), .ZN(new_n4820_));
  NAND2_X1   g03813(.A1(new_n4796_), .A2(\A[159] ), .ZN(new_n4821_));
  NAND2_X1   g03814(.A1(new_n4794_), .A2(\A[158] ), .ZN(new_n4822_));
  AOI21_X1   g03815(.A1(new_n4821_), .A2(new_n4822_), .B(new_n4799_), .ZN(new_n4823_));
  INV_X1     g03816(.I(new_n4800_), .ZN(new_n4824_));
  AOI21_X1   g03817(.A1(new_n4824_), .A2(new_n4801_), .B(\A[157] ), .ZN(new_n4825_));
  NOR2_X1    g03818(.A1(new_n4825_), .A2(new_n4823_), .ZN(new_n4826_));
  NAND2_X1   g03819(.A1(new_n4807_), .A2(\A[162] ), .ZN(new_n4827_));
  NAND2_X1   g03820(.A1(new_n4805_), .A2(\A[161] ), .ZN(new_n4828_));
  AOI21_X1   g03821(.A1(new_n4827_), .A2(new_n4828_), .B(new_n4810_), .ZN(new_n4829_));
  INV_X1     g03822(.I(new_n4811_), .ZN(new_n4830_));
  AOI21_X1   g03823(.A1(new_n4830_), .A2(new_n4815_), .B(\A[160] ), .ZN(new_n4831_));
  NOR2_X1    g03824(.A1(new_n4831_), .A2(new_n4829_), .ZN(new_n4832_));
  NOR2_X1    g03825(.A1(new_n4826_), .A2(new_n4832_), .ZN(new_n4833_));
  NOR2_X1    g03826(.A1(new_n4833_), .A2(new_n4820_), .ZN(new_n4834_));
  INV_X1     g03827(.I(\A[151] ), .ZN(new_n4835_));
  INV_X1     g03828(.I(\A[152] ), .ZN(new_n4836_));
  NAND2_X1   g03829(.A1(new_n4836_), .A2(\A[153] ), .ZN(new_n4837_));
  INV_X1     g03830(.I(\A[153] ), .ZN(new_n4838_));
  NAND2_X1   g03831(.A1(new_n4838_), .A2(\A[152] ), .ZN(new_n4839_));
  AOI21_X1   g03832(.A1(new_n4837_), .A2(new_n4839_), .B(new_n4835_), .ZN(new_n4840_));
  NOR2_X1    g03833(.A1(\A[152] ), .A2(\A[153] ), .ZN(new_n4841_));
  INV_X1     g03834(.I(new_n4841_), .ZN(new_n4842_));
  NAND2_X1   g03835(.A1(\A[152] ), .A2(\A[153] ), .ZN(new_n4843_));
  AOI21_X1   g03836(.A1(new_n4842_), .A2(new_n4843_), .B(\A[151] ), .ZN(new_n4844_));
  NOR2_X1    g03837(.A1(new_n4844_), .A2(new_n4840_), .ZN(new_n4845_));
  INV_X1     g03838(.I(\A[154] ), .ZN(new_n4846_));
  INV_X1     g03839(.I(\A[155] ), .ZN(new_n4847_));
  NAND2_X1   g03840(.A1(new_n4847_), .A2(\A[156] ), .ZN(new_n4848_));
  INV_X1     g03841(.I(\A[156] ), .ZN(new_n4849_));
  NAND2_X1   g03842(.A1(new_n4849_), .A2(\A[155] ), .ZN(new_n4850_));
  AOI21_X1   g03843(.A1(new_n4848_), .A2(new_n4850_), .B(new_n4846_), .ZN(new_n4851_));
  OR2_X2     g03844(.A1(\A[155] ), .A2(\A[156] ), .Z(new_n4852_));
  NAND2_X1   g03845(.A1(\A[155] ), .A2(\A[156] ), .ZN(new_n4853_));
  AOI21_X1   g03846(.A1(new_n4852_), .A2(new_n4853_), .B(\A[154] ), .ZN(new_n4854_));
  NOR2_X1    g03847(.A1(new_n4851_), .A2(new_n4854_), .ZN(new_n4855_));
  NOR2_X1    g03848(.A1(\A[155] ), .A2(\A[156] ), .ZN(new_n4856_));
  AOI21_X1   g03849(.A1(new_n4846_), .A2(new_n4853_), .B(new_n4856_), .ZN(new_n4857_));
  AOI21_X1   g03850(.A1(new_n4835_), .A2(new_n4843_), .B(new_n4841_), .ZN(new_n4858_));
  NAND2_X1   g03851(.A1(new_n4857_), .A2(new_n4858_), .ZN(new_n4859_));
  NAND2_X1   g03852(.A1(new_n4834_), .A2(new_n4819_), .ZN(new_n4861_));
  INV_X1     g03853(.I(new_n4861_), .ZN(new_n4862_));
  NOR3_X1    g03854(.A1(new_n4793_), .A2(new_n4791_), .A3(new_n4862_), .ZN(new_n4863_));
  AOI21_X1   g03855(.A1(new_n4788_), .A2(new_n4783_), .B(new_n4863_), .ZN(new_n4864_));
  INV_X1     g03856(.I(new_n4791_), .ZN(new_n4865_));
  NAND3_X1   g03857(.A1(new_n4865_), .A2(new_n4792_), .A3(new_n4861_), .ZN(new_n4866_));
  NOR3_X1    g03858(.A1(new_n4776_), .A2(new_n4769_), .A3(new_n4866_), .ZN(new_n4867_));
  INV_X1     g03859(.I(new_n4817_), .ZN(new_n4868_));
  AOI21_X1   g03860(.A1(new_n4826_), .A2(new_n4832_), .B(new_n4868_), .ZN(new_n4869_));
  NOR3_X1    g03861(.A1(new_n4804_), .A2(new_n4814_), .A3(new_n4817_), .ZN(new_n4870_));
  OAI21_X1   g03862(.A1(new_n4869_), .A2(new_n4870_), .B(new_n4816_), .ZN(new_n4871_));
  INV_X1     g03863(.I(new_n4816_), .ZN(new_n4872_));
  OAI21_X1   g03864(.A1(new_n4804_), .A2(new_n4814_), .B(new_n4817_), .ZN(new_n4873_));
  NAND3_X1   g03865(.A1(new_n4826_), .A2(new_n4832_), .A3(new_n4868_), .ZN(new_n4874_));
  NAND3_X1   g03866(.A1(new_n4874_), .A2(new_n4873_), .A3(new_n4872_), .ZN(new_n4875_));
  NAND2_X1   g03867(.A1(new_n4871_), .A2(new_n4875_), .ZN(new_n4876_));
  NOR4_X1    g03868(.A1(new_n4840_), .A2(new_n4844_), .A3(new_n4851_), .A4(new_n4854_), .ZN(new_n4877_));
  NOR2_X1    g03869(.A1(new_n4845_), .A2(new_n4855_), .ZN(new_n4878_));
  NOR2_X1    g03870(.A1(new_n4878_), .A2(new_n4877_), .ZN(new_n4879_));
  NAND3_X1   g03871(.A1(new_n4834_), .A2(new_n4879_), .A3(new_n4819_), .ZN(new_n4880_));
  NAND2_X1   g03872(.A1(new_n4845_), .A2(new_n4855_), .ZN(new_n4881_));
  NAND2_X1   g03873(.A1(new_n4826_), .A2(new_n4814_), .ZN(new_n4882_));
  NAND2_X1   g03874(.A1(new_n4832_), .A2(new_n4804_), .ZN(new_n4883_));
  AOI21_X1   g03875(.A1(new_n4883_), .A2(new_n4882_), .B(new_n4818_), .ZN(new_n4884_));
  NOR3_X1    g03876(.A1(new_n4884_), .A2(new_n4881_), .A3(new_n4859_), .ZN(new_n4885_));
  OAI21_X1   g03877(.A1(new_n4876_), .A2(new_n4880_), .B(new_n4885_), .ZN(new_n4886_));
  INV_X1     g03878(.I(new_n4857_), .ZN(new_n4887_));
  NOR2_X1    g03879(.A1(new_n4838_), .A2(\A[152] ), .ZN(new_n4888_));
  NOR2_X1    g03880(.A1(new_n4836_), .A2(\A[153] ), .ZN(new_n4889_));
  OAI21_X1   g03881(.A1(new_n4888_), .A2(new_n4889_), .B(\A[151] ), .ZN(new_n4890_));
  INV_X1     g03882(.I(new_n4843_), .ZN(new_n4891_));
  OAI21_X1   g03883(.A1(new_n4891_), .A2(new_n4841_), .B(new_n4835_), .ZN(new_n4892_));
  NAND2_X1   g03884(.A1(new_n4890_), .A2(new_n4892_), .ZN(new_n4893_));
  NOR2_X1    g03885(.A1(new_n4849_), .A2(\A[155] ), .ZN(new_n4894_));
  NOR2_X1    g03886(.A1(new_n4847_), .A2(\A[156] ), .ZN(new_n4895_));
  OAI21_X1   g03887(.A1(new_n4894_), .A2(new_n4895_), .B(\A[154] ), .ZN(new_n4896_));
  AND2_X2    g03888(.A1(\A[155] ), .A2(\A[156] ), .Z(new_n4897_));
  OAI21_X1   g03889(.A1(new_n4897_), .A2(new_n4856_), .B(new_n4846_), .ZN(new_n4898_));
  NAND2_X1   g03890(.A1(new_n4896_), .A2(new_n4898_), .ZN(new_n4899_));
  OAI21_X1   g03891(.A1(new_n4893_), .A2(new_n4899_), .B(new_n4858_), .ZN(new_n4900_));
  INV_X1     g03892(.I(new_n4858_), .ZN(new_n4901_));
  NAND3_X1   g03893(.A1(new_n4845_), .A2(new_n4855_), .A3(new_n4901_), .ZN(new_n4902_));
  AOI21_X1   g03894(.A1(new_n4900_), .A2(new_n4902_), .B(new_n4887_), .ZN(new_n4903_));
  NOR2_X1    g03895(.A1(new_n4877_), .A2(new_n4901_), .ZN(new_n4904_));
  NOR3_X1    g03896(.A1(new_n4893_), .A2(new_n4899_), .A3(new_n4858_), .ZN(new_n4905_));
  NOR3_X1    g03897(.A1(new_n4904_), .A2(new_n4857_), .A3(new_n4905_), .ZN(new_n4906_));
  NOR2_X1    g03898(.A1(new_n4906_), .A2(new_n4903_), .ZN(new_n4907_));
  NOR2_X1    g03899(.A1(new_n4886_), .A2(new_n4907_), .ZN(new_n4908_));
  OAI21_X1   g03900(.A1(new_n4904_), .A2(new_n4905_), .B(new_n4857_), .ZN(new_n4909_));
  NAND3_X1   g03901(.A1(new_n4900_), .A2(new_n4902_), .A3(new_n4887_), .ZN(new_n4910_));
  NAND2_X1   g03902(.A1(new_n4909_), .A2(new_n4910_), .ZN(new_n4911_));
  NOR3_X1    g03903(.A1(new_n4893_), .A2(new_n4899_), .A3(new_n4859_), .ZN(new_n4912_));
  NAND4_X1   g03904(.A1(new_n4834_), .A2(new_n4879_), .A3(new_n4819_), .A4(new_n4912_), .ZN(new_n4913_));
  NAND2_X1   g03905(.A1(new_n4911_), .A2(new_n4913_), .ZN(new_n4914_));
  INV_X1     g03906(.I(new_n4818_), .ZN(new_n4915_));
  NOR2_X1    g03907(.A1(new_n4832_), .A2(new_n4804_), .ZN(new_n4916_));
  NOR2_X1    g03908(.A1(new_n4826_), .A2(new_n4814_), .ZN(new_n4917_));
  OAI21_X1   g03909(.A1(new_n4916_), .A2(new_n4917_), .B(new_n4915_), .ZN(new_n4918_));
  NAND3_X1   g03910(.A1(new_n4871_), .A2(new_n4875_), .A3(new_n4918_), .ZN(new_n4919_));
  OAI21_X1   g03911(.A1(new_n4911_), .A2(new_n4913_), .B(new_n4919_), .ZN(new_n4920_));
  NAND2_X1   g03912(.A1(new_n4826_), .A2(new_n4832_), .ZN(new_n4921_));
  NAND2_X1   g03913(.A1(new_n4804_), .A2(new_n4814_), .ZN(new_n4922_));
  NAND3_X1   g03914(.A1(new_n4819_), .A2(new_n4921_), .A3(new_n4922_), .ZN(new_n4923_));
  NAND2_X1   g03915(.A1(new_n4893_), .A2(new_n4899_), .ZN(new_n4924_));
  NAND3_X1   g03916(.A1(new_n4912_), .A2(new_n4881_), .A3(new_n4924_), .ZN(new_n4925_));
  NOR2_X1    g03917(.A1(new_n4923_), .A2(new_n4925_), .ZN(new_n4926_));
  AOI21_X1   g03918(.A1(new_n4874_), .A2(new_n4873_), .B(new_n4872_), .ZN(new_n4927_));
  NOR3_X1    g03919(.A1(new_n4869_), .A2(new_n4870_), .A3(new_n4816_), .ZN(new_n4928_));
  NOR3_X1    g03920(.A1(new_n4928_), .A2(new_n4927_), .A3(new_n4884_), .ZN(new_n4929_));
  NAND3_X1   g03921(.A1(new_n4929_), .A2(new_n4907_), .A3(new_n4926_), .ZN(new_n4930_));
  NAND2_X1   g03922(.A1(new_n4920_), .A2(new_n4930_), .ZN(new_n4931_));
  AOI21_X1   g03923(.A1(new_n4931_), .A2(new_n4914_), .B(new_n4908_), .ZN(new_n4932_));
  OAI22_X1   g03924(.A1(new_n4864_), .A2(new_n4867_), .B1(new_n4932_), .B2(new_n4777_), .ZN(new_n4933_));
  OAI21_X1   g03925(.A1(new_n4742_), .A2(new_n4767_), .B(new_n4692_), .ZN(new_n4934_));
  NOR2_X1    g03926(.A1(new_n4696_), .A2(new_n4700_), .ZN(new_n4935_));
  OAI21_X1   g03927(.A1(new_n4734_), .A2(new_n4935_), .B(new_n4701_), .ZN(new_n4936_));
  NAND2_X1   g03928(.A1(new_n4688_), .A2(new_n4658_), .ZN(new_n4937_));
  AOI21_X1   g03929(.A1(new_n4673_), .A2(new_n4937_), .B(new_n4751_), .ZN(new_n4938_));
  XOR2_X1    g03930(.A1(new_n4938_), .A2(new_n4936_), .Z(new_n4939_));
  NAND3_X1   g03931(.A1(new_n4934_), .A2(new_n4787_), .A3(new_n4939_), .ZN(new_n4940_));
  NOR2_X1    g03932(.A1(new_n4928_), .A2(new_n4927_), .ZN(new_n4941_));
  NOR3_X1    g03933(.A1(new_n4923_), .A2(new_n4877_), .A3(new_n4878_), .ZN(new_n4942_));
  NAND2_X1   g03934(.A1(new_n4918_), .A2(new_n4912_), .ZN(new_n4943_));
  AOI21_X1   g03935(.A1(new_n4941_), .A2(new_n4942_), .B(new_n4943_), .ZN(new_n4944_));
  AOI21_X1   g03936(.A1(new_n4919_), .A2(new_n4926_), .B(new_n4907_), .ZN(new_n4945_));
  NOR2_X1    g03937(.A1(new_n4816_), .A2(new_n4817_), .ZN(new_n4946_));
  OAI21_X1   g03938(.A1(new_n4921_), .A2(new_n4946_), .B(new_n4818_), .ZN(new_n4947_));
  NOR2_X1    g03939(.A1(new_n4857_), .A2(new_n4858_), .ZN(new_n4948_));
  OAI21_X1   g03940(.A1(new_n4881_), .A2(new_n4948_), .B(new_n4859_), .ZN(new_n4949_));
  XOR2_X1    g03941(.A1(new_n4947_), .A2(new_n4949_), .Z(new_n4950_));
  NOR3_X1    g03942(.A1(new_n4945_), .A2(new_n4944_), .A3(new_n4950_), .ZN(new_n4951_));
  XOR2_X1    g03943(.A1(new_n4940_), .A2(new_n4951_), .Z(new_n4952_));
  NOR2_X1    g03944(.A1(new_n4933_), .A2(new_n4952_), .ZN(new_n4953_));
  NAND2_X1   g03945(.A1(new_n4788_), .A2(new_n4783_), .ZN(new_n4954_));
  OAI21_X1   g03946(.A1(new_n4776_), .A2(new_n4769_), .B(new_n4866_), .ZN(new_n4955_));
  NAND3_X1   g03947(.A1(new_n4788_), .A2(new_n4783_), .A3(new_n4863_), .ZN(new_n4956_));
  NAND2_X1   g03948(.A1(new_n4944_), .A2(new_n4911_), .ZN(new_n4957_));
  NOR4_X1    g03949(.A1(new_n4923_), .A2(new_n4906_), .A3(new_n4903_), .A4(new_n4925_), .ZN(new_n4958_));
  NOR2_X1    g03950(.A1(new_n4958_), .A2(new_n4929_), .ZN(new_n4959_));
  NOR3_X1    g03951(.A1(new_n4919_), .A2(new_n4911_), .A3(new_n4913_), .ZN(new_n4960_));
  OAI21_X1   g03952(.A1(new_n4959_), .A2(new_n4960_), .B(new_n4914_), .ZN(new_n4961_));
  NAND2_X1   g03953(.A1(new_n4961_), .A2(new_n4957_), .ZN(new_n4962_));
  AOI22_X1   g03954(.A1(new_n4955_), .A2(new_n4956_), .B1(new_n4962_), .B2(new_n4954_), .ZN(new_n4963_));
  AOI21_X1   g03955(.A1(new_n4760_), .A2(new_n4753_), .B(new_n4780_), .ZN(new_n4964_));
  INV_X1     g03956(.I(new_n4939_), .ZN(new_n4965_));
  NOR3_X1    g03957(.A1(new_n4964_), .A2(new_n4775_), .A3(new_n4965_), .ZN(new_n4966_));
  NOR2_X1    g03958(.A1(new_n4966_), .A2(new_n4951_), .ZN(new_n4967_));
  OAI21_X1   g03959(.A1(new_n4929_), .A2(new_n4913_), .B(new_n4911_), .ZN(new_n4968_));
  XNOR2_X1   g03960(.A1(new_n4947_), .A2(new_n4949_), .ZN(new_n4969_));
  NAND3_X1   g03961(.A1(new_n4886_), .A2(new_n4968_), .A3(new_n4969_), .ZN(new_n4970_));
  NOR2_X1    g03962(.A1(new_n4940_), .A2(new_n4970_), .ZN(new_n4971_));
  NOR2_X1    g03963(.A1(new_n4967_), .A2(new_n4971_), .ZN(new_n4972_));
  NOR2_X1    g03964(.A1(new_n4963_), .A2(new_n4972_), .ZN(new_n4973_));
  NOR4_X1    g03965(.A1(new_n4629_), .A2(new_n4953_), .A3(new_n4649_), .A4(new_n4973_), .ZN(new_n4974_));
  NOR2_X1    g03966(.A1(new_n4867_), .A2(new_n4864_), .ZN(new_n4975_));
  NAND2_X1   g03967(.A1(new_n4975_), .A2(new_n4932_), .ZN(new_n4976_));
  AOI21_X1   g03968(.A1(new_n4865_), .A2(new_n4792_), .B(new_n4861_), .ZN(new_n4977_));
  NOR2_X1    g03969(.A1(new_n4977_), .A2(new_n4863_), .ZN(new_n4978_));
  OAI21_X1   g03970(.A1(new_n4466_), .A2(new_n4469_), .B(new_n4538_), .ZN(new_n4979_));
  NAND3_X1   g03971(.A1(new_n4978_), .A2(new_n4542_), .A3(new_n4979_), .ZN(new_n4980_));
  NAND2_X1   g03972(.A1(new_n4976_), .A2(new_n4980_), .ZN(new_n4981_));
  INV_X1     g03973(.I(new_n4980_), .ZN(new_n4982_));
  NAND3_X1   g03974(.A1(new_n4982_), .A2(new_n4975_), .A3(new_n4932_), .ZN(new_n4983_));
  OAI21_X1   g03975(.A1(new_n4543_), .A2(new_n4540_), .B(new_n4608_), .ZN(new_n4984_));
  NAND3_X1   g03976(.A1(new_n4631_), .A2(new_n4638_), .A3(new_n4632_), .ZN(new_n4985_));
  NAND2_X1   g03977(.A1(new_n4984_), .A2(new_n4985_), .ZN(new_n4986_));
  AOI22_X1   g03978(.A1(new_n4981_), .A2(new_n4983_), .B1(new_n4986_), .B2(new_n4976_), .ZN(new_n4987_));
  OAI22_X1   g03979(.A1(new_n4629_), .A2(new_n4649_), .B1(new_n4953_), .B2(new_n4973_), .ZN(new_n4988_));
  AOI21_X1   g03980(.A1(new_n4987_), .A2(new_n4988_), .B(new_n4974_), .ZN(new_n4989_));
  INV_X1     g03981(.I(new_n4612_), .ZN(new_n4990_));
  NAND2_X1   g03982(.A1(new_n4990_), .A2(new_n4614_), .ZN(new_n4991_));
  NOR2_X1    g03983(.A1(new_n4640_), .A2(new_n4449_), .ZN(new_n4992_));
  OAI21_X1   g03984(.A1(new_n4990_), .A2(new_n4614_), .B(new_n4992_), .ZN(new_n4993_));
  NAND2_X1   g03985(.A1(new_n4993_), .A2(new_n4991_), .ZN(new_n4994_));
  INV_X1     g03986(.I(new_n4623_), .ZN(new_n4995_));
  INV_X1     g03987(.I(new_n4625_), .ZN(new_n4996_));
  NOR2_X1    g03988(.A1(new_n4996_), .A2(new_n4995_), .ZN(new_n4997_));
  NAND2_X1   g03989(.A1(new_n4644_), .A2(new_n4562_), .ZN(new_n4998_));
  AOI21_X1   g03990(.A1(new_n4995_), .A2(new_n4996_), .B(new_n4998_), .ZN(new_n4999_));
  NOR2_X1    g03991(.A1(new_n4999_), .A2(new_n4997_), .ZN(new_n5000_));
  NAND2_X1   g03992(.A1(new_n4616_), .A2(new_n4646_), .ZN(new_n5001_));
  NAND2_X1   g03993(.A1(new_n4642_), .A2(new_n4627_), .ZN(new_n5002_));
  AOI21_X1   g03994(.A1(new_n4609_), .A2(new_n5001_), .B(new_n5002_), .ZN(new_n5003_));
  NOR2_X1    g03995(.A1(new_n5003_), .A2(new_n5000_), .ZN(new_n5004_));
  NAND4_X1   g03996(.A1(new_n4639_), .A2(new_n5000_), .A3(new_n4642_), .A4(new_n4627_), .ZN(new_n5005_));
  INV_X1     g03997(.I(new_n5005_), .ZN(new_n5006_));
  OAI21_X1   g03998(.A1(new_n5004_), .A2(new_n5006_), .B(new_n4994_), .ZN(new_n5007_));
  INV_X1     g03999(.I(new_n4994_), .ZN(new_n5008_));
  INV_X1     g04000(.I(new_n5000_), .ZN(new_n5009_));
  NAND3_X1   g04001(.A1(new_n4639_), .A2(new_n4642_), .A3(new_n4627_), .ZN(new_n5010_));
  NAND2_X1   g04002(.A1(new_n5010_), .A2(new_n5009_), .ZN(new_n5011_));
  NAND3_X1   g04003(.A1(new_n5011_), .A2(new_n5008_), .A3(new_n5005_), .ZN(new_n5012_));
  NAND2_X1   g04004(.A1(new_n5007_), .A2(new_n5012_), .ZN(new_n5013_));
  INV_X1     g04005(.I(new_n4938_), .ZN(new_n5014_));
  NAND2_X1   g04006(.A1(new_n5014_), .A2(new_n4936_), .ZN(new_n5015_));
  NOR2_X1    g04007(.A1(new_n4964_), .A2(new_n4775_), .ZN(new_n5016_));
  OAI21_X1   g04008(.A1(new_n4936_), .A2(new_n5014_), .B(new_n5016_), .ZN(new_n5017_));
  NAND2_X1   g04009(.A1(new_n5017_), .A2(new_n5015_), .ZN(new_n5018_));
  INV_X1     g04010(.I(new_n5018_), .ZN(new_n5019_));
  NAND3_X1   g04011(.A1(new_n4963_), .A2(new_n4966_), .A3(new_n4951_), .ZN(new_n5020_));
  NAND2_X1   g04012(.A1(new_n4947_), .A2(new_n4949_), .ZN(new_n5021_));
  NOR2_X1    g04013(.A1(new_n4945_), .A2(new_n4944_), .ZN(new_n5022_));
  OAI21_X1   g04014(.A1(new_n4947_), .A2(new_n4949_), .B(new_n5022_), .ZN(new_n5023_));
  NAND2_X1   g04015(.A1(new_n5023_), .A2(new_n5021_), .ZN(new_n5024_));
  NAND2_X1   g04016(.A1(new_n5020_), .A2(new_n5024_), .ZN(new_n5025_));
  INV_X1     g04017(.I(new_n5024_), .ZN(new_n5026_));
  NAND4_X1   g04018(.A1(new_n5026_), .A2(new_n4963_), .A3(new_n4966_), .A4(new_n4951_), .ZN(new_n5027_));
  AOI21_X1   g04019(.A1(new_n5025_), .A2(new_n5027_), .B(new_n5019_), .ZN(new_n5028_));
  NAND2_X1   g04020(.A1(new_n4940_), .A2(new_n4970_), .ZN(new_n5029_));
  NAND2_X1   g04021(.A1(new_n4933_), .A2(new_n5029_), .ZN(new_n5030_));
  AOI21_X1   g04022(.A1(new_n5030_), .A2(new_n4971_), .B(new_n5026_), .ZN(new_n5031_));
  NOR4_X1    g04023(.A1(new_n4933_), .A2(new_n4940_), .A3(new_n4970_), .A4(new_n5024_), .ZN(new_n5032_));
  NOR3_X1    g04024(.A1(new_n5031_), .A2(new_n5018_), .A3(new_n5032_), .ZN(new_n5033_));
  NOR2_X1    g04025(.A1(new_n5033_), .A2(new_n5028_), .ZN(new_n5034_));
  NAND2_X1   g04026(.A1(new_n5013_), .A2(new_n5034_), .ZN(new_n5035_));
  AOI21_X1   g04027(.A1(new_n5011_), .A2(new_n5005_), .B(new_n5008_), .ZN(new_n5036_));
  NOR3_X1    g04028(.A1(new_n5004_), .A2(new_n5006_), .A3(new_n4994_), .ZN(new_n5037_));
  NOR2_X1    g04029(.A1(new_n5037_), .A2(new_n5036_), .ZN(new_n5038_));
  OAI21_X1   g04030(.A1(new_n5031_), .A2(new_n5032_), .B(new_n5018_), .ZN(new_n5039_));
  NAND3_X1   g04031(.A1(new_n5025_), .A2(new_n5019_), .A3(new_n5027_), .ZN(new_n5040_));
  NAND2_X1   g04032(.A1(new_n5039_), .A2(new_n5040_), .ZN(new_n5041_));
  NAND2_X1   g04033(.A1(new_n5038_), .A2(new_n5041_), .ZN(new_n5042_));
  AOI21_X1   g04034(.A1(new_n5035_), .A2(new_n5042_), .B(new_n4989_), .ZN(new_n5043_));
  XOR2_X1    g04035(.A1(new_n4616_), .A2(new_n4646_), .Z(new_n5044_));
  NAND2_X1   g04036(.A1(new_n5044_), .A2(new_n4639_), .ZN(new_n5045_));
  NAND2_X1   g04037(.A1(new_n5002_), .A2(new_n5001_), .ZN(new_n5046_));
  NAND2_X1   g04038(.A1(new_n4609_), .A2(new_n5046_), .ZN(new_n5047_));
  XOR2_X1    g04039(.A1(new_n4940_), .A2(new_n4970_), .Z(new_n5048_));
  NAND2_X1   g04040(.A1(new_n5048_), .A2(new_n4963_), .ZN(new_n5049_));
  NAND2_X1   g04041(.A1(new_n4966_), .A2(new_n4951_), .ZN(new_n5050_));
  NAND2_X1   g04042(.A1(new_n5050_), .A2(new_n5029_), .ZN(new_n5051_));
  NAND2_X1   g04043(.A1(new_n4933_), .A2(new_n5051_), .ZN(new_n5052_));
  NAND4_X1   g04044(.A1(new_n5045_), .A2(new_n5047_), .A3(new_n5049_), .A4(new_n5052_), .ZN(new_n5053_));
  NAND2_X1   g04045(.A1(new_n4955_), .A2(new_n4956_), .ZN(new_n5054_));
  NOR2_X1    g04046(.A1(new_n5054_), .A2(new_n4962_), .ZN(new_n5055_));
  NOR2_X1    g04047(.A1(new_n5055_), .A2(new_n4982_), .ZN(new_n5056_));
  NOR2_X1    g04048(.A1(new_n4976_), .A2(new_n4980_), .ZN(new_n5057_));
  AOI21_X1   g04049(.A1(new_n4631_), .A2(new_n4632_), .B(new_n4638_), .ZN(new_n5058_));
  NOR3_X1    g04050(.A1(new_n4543_), .A2(new_n4608_), .A3(new_n4540_), .ZN(new_n5059_));
  NOR2_X1    g04051(.A1(new_n5059_), .A2(new_n5058_), .ZN(new_n5060_));
  OAI22_X1   g04052(.A1(new_n5057_), .A2(new_n5056_), .B1(new_n5055_), .B2(new_n5060_), .ZN(new_n5061_));
  AOI22_X1   g04053(.A1(new_n5045_), .A2(new_n5047_), .B1(new_n5049_), .B2(new_n5052_), .ZN(new_n5062_));
  OAI21_X1   g04054(.A1(new_n5061_), .A2(new_n5062_), .B(new_n5053_), .ZN(new_n5063_));
  NAND2_X1   g04055(.A1(new_n5038_), .A2(new_n5034_), .ZN(new_n5064_));
  NAND2_X1   g04056(.A1(new_n5013_), .A2(new_n5041_), .ZN(new_n5065_));
  AOI21_X1   g04057(.A1(new_n5064_), .A2(new_n5065_), .B(new_n5063_), .ZN(new_n5066_));
  INV_X1     g04058(.I(\A[94] ), .ZN(new_n5067_));
  NOR2_X1    g04059(.A1(\A[95] ), .A2(\A[96] ), .ZN(new_n5068_));
  NAND2_X1   g04060(.A1(\A[95] ), .A2(\A[96] ), .ZN(new_n5069_));
  AOI21_X1   g04061(.A1(new_n5067_), .A2(new_n5069_), .B(new_n5068_), .ZN(new_n5070_));
  INV_X1     g04062(.I(\A[91] ), .ZN(new_n5071_));
  NOR2_X1    g04063(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n5072_));
  NAND2_X1   g04064(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n5073_));
  AOI21_X1   g04065(.A1(new_n5071_), .A2(new_n5073_), .B(new_n5072_), .ZN(new_n5074_));
  INV_X1     g04066(.I(new_n5074_), .ZN(new_n5075_));
  INV_X1     g04067(.I(\A[92] ), .ZN(new_n5076_));
  NAND2_X1   g04068(.A1(new_n5076_), .A2(\A[93] ), .ZN(new_n5077_));
  INV_X1     g04069(.I(\A[93] ), .ZN(new_n5078_));
  NAND2_X1   g04070(.A1(new_n5078_), .A2(\A[92] ), .ZN(new_n5079_));
  AOI21_X1   g04071(.A1(new_n5077_), .A2(new_n5079_), .B(new_n5071_), .ZN(new_n5080_));
  INV_X1     g04072(.I(new_n5072_), .ZN(new_n5081_));
  AOI21_X1   g04073(.A1(new_n5081_), .A2(new_n5073_), .B(\A[91] ), .ZN(new_n5082_));
  INV_X1     g04074(.I(\A[95] ), .ZN(new_n5083_));
  NAND2_X1   g04075(.A1(new_n5083_), .A2(\A[96] ), .ZN(new_n5084_));
  INV_X1     g04076(.I(\A[96] ), .ZN(new_n5085_));
  NAND2_X1   g04077(.A1(new_n5085_), .A2(\A[95] ), .ZN(new_n5086_));
  AOI21_X1   g04078(.A1(new_n5084_), .A2(new_n5086_), .B(new_n5067_), .ZN(new_n5087_));
  INV_X1     g04079(.I(new_n5068_), .ZN(new_n5088_));
  AOI21_X1   g04080(.A1(new_n5088_), .A2(new_n5069_), .B(\A[94] ), .ZN(new_n5089_));
  NOR4_X1    g04081(.A1(new_n5080_), .A2(new_n5082_), .A3(new_n5089_), .A4(new_n5087_), .ZN(new_n5090_));
  NOR2_X1    g04082(.A1(new_n5090_), .A2(new_n5075_), .ZN(new_n5091_));
  NOR2_X1    g04083(.A1(new_n5078_), .A2(\A[92] ), .ZN(new_n5092_));
  NOR2_X1    g04084(.A1(new_n5076_), .A2(\A[93] ), .ZN(new_n5093_));
  OAI21_X1   g04085(.A1(new_n5092_), .A2(new_n5093_), .B(\A[91] ), .ZN(new_n5094_));
  INV_X1     g04086(.I(new_n5073_), .ZN(new_n5095_));
  OAI21_X1   g04087(.A1(new_n5095_), .A2(new_n5072_), .B(new_n5071_), .ZN(new_n5096_));
  NOR2_X1    g04088(.A1(new_n5085_), .A2(\A[95] ), .ZN(new_n5097_));
  NOR2_X1    g04089(.A1(new_n5083_), .A2(\A[96] ), .ZN(new_n5098_));
  OAI21_X1   g04090(.A1(new_n5097_), .A2(new_n5098_), .B(\A[94] ), .ZN(new_n5099_));
  INV_X1     g04091(.I(new_n5069_), .ZN(new_n5100_));
  OAI21_X1   g04092(.A1(new_n5100_), .A2(new_n5068_), .B(new_n5067_), .ZN(new_n5101_));
  NAND4_X1   g04093(.A1(new_n5094_), .A2(new_n5096_), .A3(new_n5099_), .A4(new_n5101_), .ZN(new_n5102_));
  NOR2_X1    g04094(.A1(new_n5102_), .A2(new_n5074_), .ZN(new_n5103_));
  OAI21_X1   g04095(.A1(new_n5091_), .A2(new_n5103_), .B(new_n5070_), .ZN(new_n5104_));
  INV_X1     g04096(.I(new_n5070_), .ZN(new_n5105_));
  NAND2_X1   g04097(.A1(new_n5102_), .A2(new_n5074_), .ZN(new_n5106_));
  NAND2_X1   g04098(.A1(new_n5090_), .A2(new_n5075_), .ZN(new_n5107_));
  NAND3_X1   g04099(.A1(new_n5107_), .A2(new_n5106_), .A3(new_n5105_), .ZN(new_n5108_));
  NAND2_X1   g04100(.A1(new_n5104_), .A2(new_n5108_), .ZN(new_n5109_));
  INV_X1     g04101(.I(\A[100] ), .ZN(new_n5110_));
  NOR2_X1    g04102(.A1(\A[101] ), .A2(\A[102] ), .ZN(new_n5111_));
  NAND2_X1   g04103(.A1(\A[101] ), .A2(\A[102] ), .ZN(new_n5112_));
  AOI21_X1   g04104(.A1(new_n5110_), .A2(new_n5112_), .B(new_n5111_), .ZN(new_n5113_));
  INV_X1     g04105(.I(\A[97] ), .ZN(new_n5114_));
  NOR2_X1    g04106(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n5115_));
  NAND2_X1   g04107(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n5116_));
  AOI21_X1   g04108(.A1(new_n5114_), .A2(new_n5116_), .B(new_n5115_), .ZN(new_n5117_));
  NAND2_X1   g04109(.A1(new_n5113_), .A2(new_n5117_), .ZN(new_n5118_));
  INV_X1     g04110(.I(\A[98] ), .ZN(new_n5119_));
  NAND2_X1   g04111(.A1(new_n5119_), .A2(\A[99] ), .ZN(new_n5120_));
  INV_X1     g04112(.I(\A[99] ), .ZN(new_n5121_));
  NAND2_X1   g04113(.A1(new_n5121_), .A2(\A[98] ), .ZN(new_n5122_));
  AOI21_X1   g04114(.A1(new_n5120_), .A2(new_n5122_), .B(new_n5114_), .ZN(new_n5123_));
  INV_X1     g04115(.I(new_n5115_), .ZN(new_n5124_));
  AOI21_X1   g04116(.A1(new_n5124_), .A2(new_n5116_), .B(\A[97] ), .ZN(new_n5125_));
  NOR2_X1    g04117(.A1(new_n5125_), .A2(new_n5123_), .ZN(new_n5126_));
  INV_X1     g04118(.I(\A[102] ), .ZN(new_n5127_));
  NOR2_X1    g04119(.A1(new_n5127_), .A2(\A[101] ), .ZN(new_n5128_));
  INV_X1     g04120(.I(\A[101] ), .ZN(new_n5129_));
  NOR2_X1    g04121(.A1(new_n5129_), .A2(\A[102] ), .ZN(new_n5130_));
  OAI21_X1   g04122(.A1(new_n5128_), .A2(new_n5130_), .B(\A[100] ), .ZN(new_n5131_));
  INV_X1     g04123(.I(new_n5112_), .ZN(new_n5132_));
  OAI21_X1   g04124(.A1(new_n5132_), .A2(new_n5111_), .B(new_n5110_), .ZN(new_n5133_));
  NAND2_X1   g04125(.A1(new_n5131_), .A2(new_n5133_), .ZN(new_n5134_));
  NAND2_X1   g04126(.A1(new_n5126_), .A2(new_n5134_), .ZN(new_n5135_));
  NOR2_X1    g04127(.A1(new_n5121_), .A2(\A[98] ), .ZN(new_n5136_));
  NOR2_X1    g04128(.A1(new_n5119_), .A2(\A[99] ), .ZN(new_n5137_));
  OAI21_X1   g04129(.A1(new_n5136_), .A2(new_n5137_), .B(\A[97] ), .ZN(new_n5138_));
  INV_X1     g04130(.I(new_n5116_), .ZN(new_n5139_));
  OAI21_X1   g04131(.A1(new_n5139_), .A2(new_n5115_), .B(new_n5114_), .ZN(new_n5140_));
  NAND2_X1   g04132(.A1(new_n5138_), .A2(new_n5140_), .ZN(new_n5141_));
  NAND2_X1   g04133(.A1(new_n5129_), .A2(\A[102] ), .ZN(new_n5142_));
  NAND2_X1   g04134(.A1(new_n5127_), .A2(\A[101] ), .ZN(new_n5143_));
  AOI21_X1   g04135(.A1(new_n5142_), .A2(new_n5143_), .B(new_n5110_), .ZN(new_n5144_));
  INV_X1     g04136(.I(new_n5111_), .ZN(new_n5145_));
  AOI21_X1   g04137(.A1(new_n5145_), .A2(new_n5112_), .B(\A[100] ), .ZN(new_n5146_));
  NOR2_X1    g04138(.A1(new_n5146_), .A2(new_n5144_), .ZN(new_n5147_));
  NAND2_X1   g04139(.A1(new_n5147_), .A2(new_n5141_), .ZN(new_n5148_));
  AOI21_X1   g04140(.A1(new_n5135_), .A2(new_n5148_), .B(new_n5118_), .ZN(new_n5149_));
  INV_X1     g04141(.I(new_n5113_), .ZN(new_n5150_));
  NAND4_X1   g04142(.A1(new_n5138_), .A2(new_n5140_), .A3(new_n5131_), .A4(new_n5133_), .ZN(new_n5151_));
  NAND2_X1   g04143(.A1(new_n5151_), .A2(new_n5117_), .ZN(new_n5152_));
  INV_X1     g04144(.I(new_n5117_), .ZN(new_n5153_));
  NAND3_X1   g04145(.A1(new_n5126_), .A2(new_n5147_), .A3(new_n5153_), .ZN(new_n5154_));
  AOI21_X1   g04146(.A1(new_n5152_), .A2(new_n5154_), .B(new_n5150_), .ZN(new_n5155_));
  AOI21_X1   g04147(.A1(new_n5126_), .A2(new_n5147_), .B(new_n5153_), .ZN(new_n5156_));
  NOR3_X1    g04148(.A1(new_n5141_), .A2(new_n5134_), .A3(new_n5117_), .ZN(new_n5157_));
  NOR3_X1    g04149(.A1(new_n5156_), .A2(new_n5157_), .A3(new_n5113_), .ZN(new_n5158_));
  NOR3_X1    g04150(.A1(new_n5155_), .A2(new_n5158_), .A3(new_n5149_), .ZN(new_n5159_));
  INV_X1     g04151(.I(new_n5118_), .ZN(new_n5160_));
  NOR4_X1    g04152(.A1(new_n5123_), .A2(new_n5125_), .A3(new_n5146_), .A4(new_n5144_), .ZN(new_n5161_));
  NAND2_X1   g04153(.A1(new_n5161_), .A2(new_n5160_), .ZN(new_n5162_));
  NAND2_X1   g04154(.A1(new_n5141_), .A2(new_n5134_), .ZN(new_n5163_));
  NAND2_X1   g04155(.A1(new_n5163_), .A2(new_n5151_), .ZN(new_n5164_));
  OAI22_X1   g04156(.A1(new_n5080_), .A2(new_n5082_), .B1(new_n5089_), .B2(new_n5087_), .ZN(new_n5165_));
  NAND2_X1   g04157(.A1(new_n5165_), .A2(new_n5102_), .ZN(new_n5166_));
  NAND3_X1   g04158(.A1(new_n5090_), .A2(new_n5070_), .A3(new_n5074_), .ZN(new_n5167_));
  NOR4_X1    g04159(.A1(new_n5164_), .A2(new_n5162_), .A3(new_n5167_), .A4(new_n5166_), .ZN(new_n5168_));
  NAND2_X1   g04160(.A1(new_n5159_), .A2(new_n5168_), .ZN(new_n5169_));
  OAI21_X1   g04161(.A1(new_n5156_), .A2(new_n5157_), .B(new_n5113_), .ZN(new_n5170_));
  NAND3_X1   g04162(.A1(new_n5152_), .A2(new_n5154_), .A3(new_n5150_), .ZN(new_n5171_));
  NAND2_X1   g04163(.A1(new_n5170_), .A2(new_n5171_), .ZN(new_n5172_));
  NOR2_X1    g04164(.A1(new_n5151_), .A2(new_n5118_), .ZN(new_n5173_));
  NOR2_X1    g04165(.A1(new_n5126_), .A2(new_n5147_), .ZN(new_n5174_));
  NOR2_X1    g04166(.A1(new_n5174_), .A2(new_n5161_), .ZN(new_n5175_));
  AOI22_X1   g04167(.A1(new_n5094_), .A2(new_n5096_), .B1(new_n5099_), .B2(new_n5101_), .ZN(new_n5176_));
  NOR2_X1    g04168(.A1(new_n5176_), .A2(new_n5090_), .ZN(new_n5177_));
  NAND2_X1   g04169(.A1(new_n5070_), .A2(new_n5074_), .ZN(new_n5178_));
  NOR2_X1    g04170(.A1(new_n5102_), .A2(new_n5178_), .ZN(new_n5179_));
  NAND4_X1   g04171(.A1(new_n5175_), .A2(new_n5177_), .A3(new_n5173_), .A4(new_n5179_), .ZN(new_n5180_));
  OAI21_X1   g04172(.A1(new_n5172_), .A2(new_n5149_), .B(new_n5180_), .ZN(new_n5181_));
  AOI21_X1   g04173(.A1(new_n5181_), .A2(new_n5169_), .B(new_n5109_), .ZN(new_n5182_));
  NOR2_X1    g04174(.A1(new_n5159_), .A2(new_n5180_), .ZN(new_n5183_));
  NOR2_X1    g04175(.A1(new_n5155_), .A2(new_n5158_), .ZN(new_n5184_));
  NOR3_X1    g04176(.A1(new_n5164_), .A2(new_n5166_), .A3(new_n5162_), .ZN(new_n5185_));
  NOR2_X1    g04177(.A1(new_n5147_), .A2(new_n5141_), .ZN(new_n5186_));
  NOR2_X1    g04178(.A1(new_n5126_), .A2(new_n5134_), .ZN(new_n5187_));
  OAI21_X1   g04179(.A1(new_n5186_), .A2(new_n5187_), .B(new_n5160_), .ZN(new_n5188_));
  NAND2_X1   g04180(.A1(new_n5188_), .A2(new_n5179_), .ZN(new_n5189_));
  AOI21_X1   g04181(.A1(new_n5184_), .A2(new_n5185_), .B(new_n5189_), .ZN(new_n5190_));
  NOR3_X1    g04182(.A1(new_n5190_), .A2(new_n5183_), .A3(new_n5109_), .ZN(new_n5191_));
  NOR2_X1    g04183(.A1(new_n5182_), .A2(new_n5191_), .ZN(new_n5192_));
  INV_X1     g04184(.I(new_n5109_), .ZN(new_n5193_));
  NOR4_X1    g04185(.A1(new_n5180_), .A2(new_n5149_), .A3(new_n5155_), .A4(new_n5158_), .ZN(new_n5194_));
  NOR2_X1    g04186(.A1(new_n5159_), .A2(new_n5168_), .ZN(new_n5195_));
  OAI21_X1   g04187(.A1(new_n5195_), .A2(new_n5194_), .B(new_n5193_), .ZN(new_n5196_));
  OAI21_X1   g04188(.A1(new_n5172_), .A2(new_n5149_), .B(new_n5168_), .ZN(new_n5197_));
  NOR4_X1    g04189(.A1(new_n5090_), .A2(new_n5176_), .A3(new_n5151_), .A4(new_n5118_), .ZN(new_n5198_));
  NAND4_X1   g04190(.A1(new_n5170_), .A2(new_n5171_), .A3(new_n5175_), .A4(new_n5198_), .ZN(new_n5199_));
  NAND3_X1   g04191(.A1(new_n5199_), .A2(new_n5188_), .A3(new_n5179_), .ZN(new_n5200_));
  NAND3_X1   g04192(.A1(new_n5200_), .A2(new_n5197_), .A3(new_n5193_), .ZN(new_n5201_));
  NAND2_X1   g04193(.A1(new_n5175_), .A2(new_n5173_), .ZN(new_n5202_));
  NOR2_X1    g04194(.A1(new_n5167_), .A2(new_n5166_), .ZN(new_n5203_));
  NAND2_X1   g04195(.A1(new_n5202_), .A2(new_n5203_), .ZN(new_n5204_));
  NOR2_X1    g04196(.A1(new_n5164_), .A2(new_n5162_), .ZN(new_n5205_));
  NAND2_X1   g04197(.A1(new_n5177_), .A2(new_n5179_), .ZN(new_n5206_));
  NAND2_X1   g04198(.A1(new_n5205_), .A2(new_n5206_), .ZN(new_n5207_));
  NAND2_X1   g04199(.A1(new_n5204_), .A2(new_n5207_), .ZN(new_n5208_));
  INV_X1     g04200(.I(\A[87] ), .ZN(new_n5209_));
  NOR2_X1    g04201(.A1(new_n5209_), .A2(\A[86] ), .ZN(new_n5210_));
  INV_X1     g04202(.I(\A[86] ), .ZN(new_n5211_));
  NOR2_X1    g04203(.A1(new_n5211_), .A2(\A[87] ), .ZN(new_n5212_));
  OAI21_X1   g04204(.A1(new_n5210_), .A2(new_n5212_), .B(\A[85] ), .ZN(new_n5213_));
  INV_X1     g04205(.I(\A[85] ), .ZN(new_n5214_));
  NOR2_X1    g04206(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n5215_));
  NAND2_X1   g04207(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n5216_));
  INV_X1     g04208(.I(new_n5216_), .ZN(new_n5217_));
  OAI21_X1   g04209(.A1(new_n5217_), .A2(new_n5215_), .B(new_n5214_), .ZN(new_n5218_));
  NAND2_X1   g04210(.A1(new_n5213_), .A2(new_n5218_), .ZN(new_n5219_));
  INV_X1     g04211(.I(\A[90] ), .ZN(new_n5220_));
  NOR2_X1    g04212(.A1(new_n5220_), .A2(\A[89] ), .ZN(new_n5221_));
  INV_X1     g04213(.I(\A[89] ), .ZN(new_n5222_));
  NOR2_X1    g04214(.A1(new_n5222_), .A2(\A[90] ), .ZN(new_n5223_));
  OAI21_X1   g04215(.A1(new_n5221_), .A2(new_n5223_), .B(\A[88] ), .ZN(new_n5224_));
  INV_X1     g04216(.I(\A[88] ), .ZN(new_n5225_));
  NOR2_X1    g04217(.A1(\A[89] ), .A2(\A[90] ), .ZN(new_n5226_));
  NAND2_X1   g04218(.A1(\A[89] ), .A2(\A[90] ), .ZN(new_n5227_));
  INV_X1     g04219(.I(new_n5227_), .ZN(new_n5228_));
  OAI21_X1   g04220(.A1(new_n5228_), .A2(new_n5226_), .B(new_n5225_), .ZN(new_n5229_));
  NAND2_X1   g04221(.A1(new_n5224_), .A2(new_n5229_), .ZN(new_n5230_));
  AOI21_X1   g04222(.A1(new_n5225_), .A2(new_n5227_), .B(new_n5226_), .ZN(new_n5231_));
  AOI21_X1   g04223(.A1(new_n5214_), .A2(new_n5216_), .B(new_n5215_), .ZN(new_n5232_));
  NAND2_X1   g04224(.A1(new_n5231_), .A2(new_n5232_), .ZN(new_n5233_));
  NOR3_X1    g04225(.A1(new_n5219_), .A2(new_n5230_), .A3(new_n5233_), .ZN(new_n5234_));
  NOR2_X1    g04226(.A1(new_n5219_), .A2(new_n5230_), .ZN(new_n5235_));
  NAND2_X1   g04227(.A1(new_n5211_), .A2(\A[87] ), .ZN(new_n5236_));
  NAND2_X1   g04228(.A1(new_n5209_), .A2(\A[86] ), .ZN(new_n5237_));
  AOI21_X1   g04229(.A1(new_n5236_), .A2(new_n5237_), .B(new_n5214_), .ZN(new_n5238_));
  INV_X1     g04230(.I(new_n5215_), .ZN(new_n5239_));
  AOI21_X1   g04231(.A1(new_n5239_), .A2(new_n5216_), .B(\A[85] ), .ZN(new_n5240_));
  NOR2_X1    g04232(.A1(new_n5240_), .A2(new_n5238_), .ZN(new_n5241_));
  NAND2_X1   g04233(.A1(new_n5222_), .A2(\A[90] ), .ZN(new_n5242_));
  NAND2_X1   g04234(.A1(new_n5220_), .A2(\A[89] ), .ZN(new_n5243_));
  AOI21_X1   g04235(.A1(new_n5242_), .A2(new_n5243_), .B(new_n5225_), .ZN(new_n5244_));
  INV_X1     g04236(.I(new_n5226_), .ZN(new_n5245_));
  AOI21_X1   g04237(.A1(new_n5245_), .A2(new_n5227_), .B(\A[88] ), .ZN(new_n5246_));
  NOR2_X1    g04238(.A1(new_n5246_), .A2(new_n5244_), .ZN(new_n5247_));
  NOR2_X1    g04239(.A1(new_n5241_), .A2(new_n5247_), .ZN(new_n5248_));
  NOR2_X1    g04240(.A1(new_n5248_), .A2(new_n5235_), .ZN(new_n5249_));
  INV_X1     g04241(.I(\A[79] ), .ZN(new_n5250_));
  INV_X1     g04242(.I(\A[80] ), .ZN(new_n5251_));
  NAND2_X1   g04243(.A1(new_n5251_), .A2(\A[81] ), .ZN(new_n5252_));
  INV_X1     g04244(.I(\A[81] ), .ZN(new_n5253_));
  NAND2_X1   g04245(.A1(new_n5253_), .A2(\A[80] ), .ZN(new_n5254_));
  AOI21_X1   g04246(.A1(new_n5252_), .A2(new_n5254_), .B(new_n5250_), .ZN(new_n5255_));
  NOR2_X1    g04247(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n5256_));
  INV_X1     g04248(.I(new_n5256_), .ZN(new_n5257_));
  NAND2_X1   g04249(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n5258_));
  AOI21_X1   g04250(.A1(new_n5257_), .A2(new_n5258_), .B(\A[79] ), .ZN(new_n5259_));
  NOR2_X1    g04251(.A1(new_n5259_), .A2(new_n5255_), .ZN(new_n5260_));
  INV_X1     g04252(.I(\A[82] ), .ZN(new_n5261_));
  INV_X1     g04253(.I(\A[83] ), .ZN(new_n5262_));
  NAND2_X1   g04254(.A1(new_n5262_), .A2(\A[84] ), .ZN(new_n5263_));
  INV_X1     g04255(.I(\A[84] ), .ZN(new_n5264_));
  NAND2_X1   g04256(.A1(new_n5264_), .A2(\A[83] ), .ZN(new_n5265_));
  AOI21_X1   g04257(.A1(new_n5263_), .A2(new_n5265_), .B(new_n5261_), .ZN(new_n5266_));
  NOR2_X1    g04258(.A1(\A[83] ), .A2(\A[84] ), .ZN(new_n5267_));
  INV_X1     g04259(.I(new_n5267_), .ZN(new_n5268_));
  NAND2_X1   g04260(.A1(\A[83] ), .A2(\A[84] ), .ZN(new_n5269_));
  AOI21_X1   g04261(.A1(new_n5268_), .A2(new_n5269_), .B(\A[82] ), .ZN(new_n5270_));
  NOR2_X1    g04262(.A1(new_n5270_), .A2(new_n5266_), .ZN(new_n5271_));
  AOI21_X1   g04263(.A1(new_n5261_), .A2(new_n5269_), .B(new_n5267_), .ZN(new_n5272_));
  AOI21_X1   g04264(.A1(new_n5250_), .A2(new_n5258_), .B(new_n5256_), .ZN(new_n5273_));
  NAND2_X1   g04265(.A1(new_n5272_), .A2(new_n5273_), .ZN(new_n5274_));
  NAND2_X1   g04266(.A1(new_n5249_), .A2(new_n5234_), .ZN(new_n5276_));
  INV_X1     g04267(.I(new_n5276_), .ZN(new_n5277_));
  NOR2_X1    g04268(.A1(new_n5208_), .A2(new_n5277_), .ZN(new_n5278_));
  AOI21_X1   g04269(.A1(new_n5201_), .A2(new_n5196_), .B(new_n5278_), .ZN(new_n5279_));
  NOR2_X1    g04270(.A1(new_n5205_), .A2(new_n5206_), .ZN(new_n5280_));
  NOR2_X1    g04271(.A1(new_n5202_), .A2(new_n5203_), .ZN(new_n5281_));
  NOR2_X1    g04272(.A1(new_n5281_), .A2(new_n5280_), .ZN(new_n5282_));
  NAND2_X1   g04273(.A1(new_n5282_), .A2(new_n5276_), .ZN(new_n5283_));
  NOR3_X1    g04274(.A1(new_n5182_), .A2(new_n5191_), .A3(new_n5283_), .ZN(new_n5284_));
  INV_X1     g04275(.I(new_n5232_), .ZN(new_n5285_));
  AOI21_X1   g04276(.A1(new_n5241_), .A2(new_n5247_), .B(new_n5285_), .ZN(new_n5286_));
  NOR3_X1    g04277(.A1(new_n5219_), .A2(new_n5230_), .A3(new_n5232_), .ZN(new_n5287_));
  OAI21_X1   g04278(.A1(new_n5286_), .A2(new_n5287_), .B(new_n5231_), .ZN(new_n5288_));
  INV_X1     g04279(.I(new_n5231_), .ZN(new_n5289_));
  OAI21_X1   g04280(.A1(new_n5219_), .A2(new_n5230_), .B(new_n5232_), .ZN(new_n5290_));
  NAND3_X1   g04281(.A1(new_n5241_), .A2(new_n5247_), .A3(new_n5285_), .ZN(new_n5291_));
  NAND3_X1   g04282(.A1(new_n5290_), .A2(new_n5291_), .A3(new_n5289_), .ZN(new_n5292_));
  NAND2_X1   g04283(.A1(new_n5288_), .A2(new_n5292_), .ZN(new_n5293_));
  INV_X1     g04284(.I(new_n5233_), .ZN(new_n5294_));
  NAND3_X1   g04285(.A1(new_n5294_), .A2(new_n5241_), .A3(new_n5247_), .ZN(new_n5295_));
  NOR3_X1    g04286(.A1(new_n5295_), .A2(new_n5248_), .A3(new_n5235_), .ZN(new_n5296_));
  NOR4_X1    g04287(.A1(new_n5255_), .A2(new_n5259_), .A3(new_n5270_), .A4(new_n5266_), .ZN(new_n5297_));
  NOR2_X1    g04288(.A1(new_n5260_), .A2(new_n5271_), .ZN(new_n5298_));
  NOR2_X1    g04289(.A1(new_n5298_), .A2(new_n5297_), .ZN(new_n5299_));
  NAND2_X1   g04290(.A1(new_n5296_), .A2(new_n5299_), .ZN(new_n5300_));
  NAND2_X1   g04291(.A1(new_n5260_), .A2(new_n5271_), .ZN(new_n5301_));
  NAND2_X1   g04292(.A1(new_n5241_), .A2(new_n5230_), .ZN(new_n5302_));
  NAND2_X1   g04293(.A1(new_n5247_), .A2(new_n5219_), .ZN(new_n5303_));
  AOI21_X1   g04294(.A1(new_n5302_), .A2(new_n5303_), .B(new_n5233_), .ZN(new_n5304_));
  NOR3_X1    g04295(.A1(new_n5304_), .A2(new_n5301_), .A3(new_n5274_), .ZN(new_n5305_));
  OAI21_X1   g04296(.A1(new_n5293_), .A2(new_n5300_), .B(new_n5305_), .ZN(new_n5306_));
  INV_X1     g04297(.I(new_n5273_), .ZN(new_n5307_));
  NOR2_X1    g04298(.A1(new_n5297_), .A2(new_n5307_), .ZN(new_n5308_));
  NOR2_X1    g04299(.A1(new_n5253_), .A2(\A[80] ), .ZN(new_n5309_));
  NOR2_X1    g04300(.A1(new_n5251_), .A2(\A[81] ), .ZN(new_n5310_));
  OAI21_X1   g04301(.A1(new_n5309_), .A2(new_n5310_), .B(\A[79] ), .ZN(new_n5311_));
  INV_X1     g04302(.I(new_n5258_), .ZN(new_n5312_));
  OAI21_X1   g04303(.A1(new_n5312_), .A2(new_n5256_), .B(new_n5250_), .ZN(new_n5313_));
  NAND2_X1   g04304(.A1(new_n5311_), .A2(new_n5313_), .ZN(new_n5314_));
  NOR2_X1    g04305(.A1(new_n5264_), .A2(\A[83] ), .ZN(new_n5315_));
  NOR2_X1    g04306(.A1(new_n5262_), .A2(\A[84] ), .ZN(new_n5316_));
  OAI21_X1   g04307(.A1(new_n5315_), .A2(new_n5316_), .B(\A[82] ), .ZN(new_n5317_));
  INV_X1     g04308(.I(new_n5269_), .ZN(new_n5318_));
  OAI21_X1   g04309(.A1(new_n5318_), .A2(new_n5267_), .B(new_n5261_), .ZN(new_n5319_));
  NAND2_X1   g04310(.A1(new_n5317_), .A2(new_n5319_), .ZN(new_n5320_));
  NOR3_X1    g04311(.A1(new_n5314_), .A2(new_n5320_), .A3(new_n5273_), .ZN(new_n5321_));
  OAI21_X1   g04312(.A1(new_n5308_), .A2(new_n5321_), .B(new_n5272_), .ZN(new_n5322_));
  INV_X1     g04313(.I(new_n5272_), .ZN(new_n5323_));
  OAI21_X1   g04314(.A1(new_n5314_), .A2(new_n5320_), .B(new_n5273_), .ZN(new_n5324_));
  NAND3_X1   g04315(.A1(new_n5260_), .A2(new_n5271_), .A3(new_n5307_), .ZN(new_n5325_));
  NAND3_X1   g04316(.A1(new_n5324_), .A2(new_n5325_), .A3(new_n5323_), .ZN(new_n5326_));
  NAND2_X1   g04317(.A1(new_n5322_), .A2(new_n5326_), .ZN(new_n5327_));
  INV_X1     g04318(.I(new_n5327_), .ZN(new_n5328_));
  NOR2_X1    g04319(.A1(new_n5306_), .A2(new_n5328_), .ZN(new_n5329_));
  NOR3_X1    g04320(.A1(new_n5314_), .A2(new_n5320_), .A3(new_n5274_), .ZN(new_n5330_));
  NAND3_X1   g04321(.A1(new_n5296_), .A2(new_n5330_), .A3(new_n5299_), .ZN(new_n5331_));
  NAND2_X1   g04322(.A1(new_n5331_), .A2(new_n5327_), .ZN(new_n5332_));
  NOR2_X1    g04323(.A1(new_n5247_), .A2(new_n5219_), .ZN(new_n5333_));
  NOR2_X1    g04324(.A1(new_n5241_), .A2(new_n5230_), .ZN(new_n5334_));
  OAI21_X1   g04325(.A1(new_n5333_), .A2(new_n5334_), .B(new_n5294_), .ZN(new_n5335_));
  NAND3_X1   g04326(.A1(new_n5288_), .A2(new_n5292_), .A3(new_n5335_), .ZN(new_n5336_));
  OAI21_X1   g04327(.A1(new_n5327_), .A2(new_n5331_), .B(new_n5336_), .ZN(new_n5337_));
  AOI21_X1   g04328(.A1(new_n5290_), .A2(new_n5291_), .B(new_n5289_), .ZN(new_n5338_));
  NOR3_X1    g04329(.A1(new_n5286_), .A2(new_n5287_), .A3(new_n5231_), .ZN(new_n5339_));
  NOR3_X1    g04330(.A1(new_n5339_), .A2(new_n5338_), .A3(new_n5304_), .ZN(new_n5340_));
  NAND2_X1   g04331(.A1(new_n5241_), .A2(new_n5247_), .ZN(new_n5341_));
  NAND2_X1   g04332(.A1(new_n5219_), .A2(new_n5230_), .ZN(new_n5342_));
  NAND3_X1   g04333(.A1(new_n5234_), .A2(new_n5341_), .A3(new_n5342_), .ZN(new_n5343_));
  NAND2_X1   g04334(.A1(new_n5314_), .A2(new_n5320_), .ZN(new_n5344_));
  NAND3_X1   g04335(.A1(new_n5330_), .A2(new_n5301_), .A3(new_n5344_), .ZN(new_n5345_));
  AOI21_X1   g04336(.A1(new_n5324_), .A2(new_n5325_), .B(new_n5323_), .ZN(new_n5346_));
  NOR3_X1    g04337(.A1(new_n5308_), .A2(new_n5321_), .A3(new_n5272_), .ZN(new_n5347_));
  NOR4_X1    g04338(.A1(new_n5347_), .A2(new_n5346_), .A3(new_n5343_), .A4(new_n5345_), .ZN(new_n5348_));
  NAND2_X1   g04339(.A1(new_n5348_), .A2(new_n5340_), .ZN(new_n5349_));
  NAND2_X1   g04340(.A1(new_n5337_), .A2(new_n5349_), .ZN(new_n5350_));
  AOI21_X1   g04341(.A1(new_n5350_), .A2(new_n5332_), .B(new_n5329_), .ZN(new_n5351_));
  OAI22_X1   g04342(.A1(new_n5279_), .A2(new_n5284_), .B1(new_n5351_), .B2(new_n5192_), .ZN(new_n5352_));
  OAI21_X1   g04343(.A1(new_n5159_), .A2(new_n5180_), .B(new_n5109_), .ZN(new_n5353_));
  NAND2_X1   g04344(.A1(new_n5150_), .A2(new_n5153_), .ZN(new_n5354_));
  AOI21_X1   g04345(.A1(new_n5161_), .A2(new_n5354_), .B(new_n5160_), .ZN(new_n5355_));
  NOR2_X1    g04346(.A1(new_n5070_), .A2(new_n5074_), .ZN(new_n5356_));
  OAI21_X1   g04347(.A1(new_n5102_), .A2(new_n5356_), .B(new_n5178_), .ZN(new_n5357_));
  XOR2_X1    g04348(.A1(new_n5355_), .A2(new_n5357_), .Z(new_n5358_));
  NAND3_X1   g04349(.A1(new_n5353_), .A2(new_n5200_), .A3(new_n5358_), .ZN(new_n5359_));
  OAI21_X1   g04350(.A1(new_n5340_), .A2(new_n5331_), .B(new_n5327_), .ZN(new_n5360_));
  NOR2_X1    g04351(.A1(new_n5231_), .A2(new_n5232_), .ZN(new_n5361_));
  OAI21_X1   g04352(.A1(new_n5341_), .A2(new_n5361_), .B(new_n5233_), .ZN(new_n5362_));
  NOR2_X1    g04353(.A1(new_n5272_), .A2(new_n5273_), .ZN(new_n5363_));
  OAI21_X1   g04354(.A1(new_n5301_), .A2(new_n5363_), .B(new_n5274_), .ZN(new_n5364_));
  XNOR2_X1   g04355(.A1(new_n5362_), .A2(new_n5364_), .ZN(new_n5365_));
  NAND3_X1   g04356(.A1(new_n5306_), .A2(new_n5360_), .A3(new_n5365_), .ZN(new_n5366_));
  XNOR2_X1   g04357(.A1(new_n5359_), .A2(new_n5366_), .ZN(new_n5367_));
  NOR2_X1    g04358(.A1(new_n5352_), .A2(new_n5367_), .ZN(new_n5368_));
  NAND2_X1   g04359(.A1(new_n5201_), .A2(new_n5196_), .ZN(new_n5369_));
  OAI21_X1   g04360(.A1(new_n5182_), .A2(new_n5191_), .B(new_n5283_), .ZN(new_n5370_));
  NAND3_X1   g04361(.A1(new_n5201_), .A2(new_n5196_), .A3(new_n5278_), .ZN(new_n5371_));
  NOR2_X1    g04362(.A1(new_n5339_), .A2(new_n5338_), .ZN(new_n5372_));
  NOR3_X1    g04363(.A1(new_n5343_), .A2(new_n5297_), .A3(new_n5298_), .ZN(new_n5373_));
  NAND2_X1   g04364(.A1(new_n5335_), .A2(new_n5330_), .ZN(new_n5374_));
  AOI21_X1   g04365(.A1(new_n5372_), .A2(new_n5373_), .B(new_n5374_), .ZN(new_n5375_));
  NAND2_X1   g04366(.A1(new_n5375_), .A2(new_n5327_), .ZN(new_n5376_));
  NOR2_X1    g04367(.A1(new_n5348_), .A2(new_n5340_), .ZN(new_n5377_));
  NOR3_X1    g04368(.A1(new_n5336_), .A2(new_n5331_), .A3(new_n5327_), .ZN(new_n5378_));
  OAI21_X1   g04369(.A1(new_n5377_), .A2(new_n5378_), .B(new_n5332_), .ZN(new_n5379_));
  NAND2_X1   g04370(.A1(new_n5379_), .A2(new_n5376_), .ZN(new_n5380_));
  AOI22_X1   g04371(.A1(new_n5370_), .A2(new_n5371_), .B1(new_n5380_), .B2(new_n5369_), .ZN(new_n5381_));
  INV_X1     g04372(.I(new_n5359_), .ZN(new_n5382_));
  AND3_X2    g04373(.A1(new_n5360_), .A2(new_n5306_), .A3(new_n5365_), .Z(new_n5383_));
  NOR2_X1    g04374(.A1(new_n5382_), .A2(new_n5383_), .ZN(new_n5384_));
  NOR2_X1    g04375(.A1(new_n5359_), .A2(new_n5366_), .ZN(new_n5385_));
  NOR2_X1    g04376(.A1(new_n5384_), .A2(new_n5385_), .ZN(new_n5386_));
  NOR2_X1    g04377(.A1(new_n5386_), .A2(new_n5381_), .ZN(new_n5387_));
  INV_X1     g04378(.I(\A[118] ), .ZN(new_n5388_));
  NOR2_X1    g04379(.A1(\A[119] ), .A2(\A[120] ), .ZN(new_n5389_));
  NAND2_X1   g04380(.A1(\A[119] ), .A2(\A[120] ), .ZN(new_n5390_));
  AOI21_X1   g04381(.A1(new_n5388_), .A2(new_n5390_), .B(new_n5389_), .ZN(new_n5391_));
  INV_X1     g04382(.I(\A[115] ), .ZN(new_n5392_));
  NOR2_X1    g04383(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n5393_));
  NAND2_X1   g04384(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n5394_));
  AOI21_X1   g04385(.A1(new_n5392_), .A2(new_n5394_), .B(new_n5393_), .ZN(new_n5395_));
  INV_X1     g04386(.I(new_n5395_), .ZN(new_n5396_));
  INV_X1     g04387(.I(\A[116] ), .ZN(new_n5397_));
  NAND2_X1   g04388(.A1(new_n5397_), .A2(\A[117] ), .ZN(new_n5398_));
  INV_X1     g04389(.I(\A[117] ), .ZN(new_n5399_));
  NAND2_X1   g04390(.A1(new_n5399_), .A2(\A[116] ), .ZN(new_n5400_));
  AOI21_X1   g04391(.A1(new_n5398_), .A2(new_n5400_), .B(new_n5392_), .ZN(new_n5401_));
  INV_X1     g04392(.I(new_n5393_), .ZN(new_n5402_));
  AOI21_X1   g04393(.A1(new_n5402_), .A2(new_n5394_), .B(\A[115] ), .ZN(new_n5403_));
  INV_X1     g04394(.I(\A[119] ), .ZN(new_n5404_));
  NAND2_X1   g04395(.A1(new_n5404_), .A2(\A[120] ), .ZN(new_n5405_));
  INV_X1     g04396(.I(\A[120] ), .ZN(new_n5406_));
  NAND2_X1   g04397(.A1(new_n5406_), .A2(\A[119] ), .ZN(new_n5407_));
  AOI21_X1   g04398(.A1(new_n5405_), .A2(new_n5407_), .B(new_n5388_), .ZN(new_n5408_));
  INV_X1     g04399(.I(new_n5389_), .ZN(new_n5409_));
  AOI21_X1   g04400(.A1(new_n5409_), .A2(new_n5390_), .B(\A[118] ), .ZN(new_n5410_));
  NOR4_X1    g04401(.A1(new_n5401_), .A2(new_n5403_), .A3(new_n5410_), .A4(new_n5408_), .ZN(new_n5411_));
  NOR2_X1    g04402(.A1(new_n5411_), .A2(new_n5396_), .ZN(new_n5412_));
  NOR2_X1    g04403(.A1(new_n5399_), .A2(\A[116] ), .ZN(new_n5413_));
  NOR2_X1    g04404(.A1(new_n5397_), .A2(\A[117] ), .ZN(new_n5414_));
  OAI21_X1   g04405(.A1(new_n5413_), .A2(new_n5414_), .B(\A[115] ), .ZN(new_n5415_));
  INV_X1     g04406(.I(new_n5394_), .ZN(new_n5416_));
  OAI21_X1   g04407(.A1(new_n5416_), .A2(new_n5393_), .B(new_n5392_), .ZN(new_n5417_));
  NOR2_X1    g04408(.A1(new_n5406_), .A2(\A[119] ), .ZN(new_n5418_));
  NOR2_X1    g04409(.A1(new_n5404_), .A2(\A[120] ), .ZN(new_n5419_));
  OAI21_X1   g04410(.A1(new_n5418_), .A2(new_n5419_), .B(\A[118] ), .ZN(new_n5420_));
  INV_X1     g04411(.I(new_n5390_), .ZN(new_n5421_));
  OAI21_X1   g04412(.A1(new_n5421_), .A2(new_n5389_), .B(new_n5388_), .ZN(new_n5422_));
  NAND4_X1   g04413(.A1(new_n5415_), .A2(new_n5417_), .A3(new_n5420_), .A4(new_n5422_), .ZN(new_n5423_));
  NOR2_X1    g04414(.A1(new_n5423_), .A2(new_n5395_), .ZN(new_n5424_));
  OAI21_X1   g04415(.A1(new_n5412_), .A2(new_n5424_), .B(new_n5391_), .ZN(new_n5425_));
  INV_X1     g04416(.I(new_n5391_), .ZN(new_n5426_));
  NAND2_X1   g04417(.A1(new_n5423_), .A2(new_n5395_), .ZN(new_n5427_));
  NOR2_X1    g04418(.A1(new_n5410_), .A2(new_n5408_), .ZN(new_n5428_));
  NAND4_X1   g04419(.A1(new_n5428_), .A2(new_n5396_), .A3(new_n5415_), .A4(new_n5417_), .ZN(new_n5429_));
  NAND3_X1   g04420(.A1(new_n5427_), .A2(new_n5429_), .A3(new_n5426_), .ZN(new_n5430_));
  NAND2_X1   g04421(.A1(new_n5425_), .A2(new_n5430_), .ZN(new_n5431_));
  INV_X1     g04422(.I(\A[124] ), .ZN(new_n5432_));
  NOR2_X1    g04423(.A1(\A[125] ), .A2(\A[126] ), .ZN(new_n5433_));
  NAND2_X1   g04424(.A1(\A[125] ), .A2(\A[126] ), .ZN(new_n5434_));
  AOI21_X1   g04425(.A1(new_n5432_), .A2(new_n5434_), .B(new_n5433_), .ZN(new_n5435_));
  INV_X1     g04426(.I(\A[121] ), .ZN(new_n5436_));
  NOR2_X1    g04427(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n5437_));
  NAND2_X1   g04428(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n5438_));
  AOI21_X1   g04429(.A1(new_n5436_), .A2(new_n5438_), .B(new_n5437_), .ZN(new_n5439_));
  NAND2_X1   g04430(.A1(new_n5435_), .A2(new_n5439_), .ZN(new_n5440_));
  INV_X1     g04431(.I(\A[122] ), .ZN(new_n5441_));
  NAND2_X1   g04432(.A1(new_n5441_), .A2(\A[123] ), .ZN(new_n5442_));
  INV_X1     g04433(.I(\A[123] ), .ZN(new_n5443_));
  NAND2_X1   g04434(.A1(new_n5443_), .A2(\A[122] ), .ZN(new_n5444_));
  AOI21_X1   g04435(.A1(new_n5442_), .A2(new_n5444_), .B(new_n5436_), .ZN(new_n5445_));
  INV_X1     g04436(.I(new_n5437_), .ZN(new_n5446_));
  AOI21_X1   g04437(.A1(new_n5446_), .A2(new_n5438_), .B(\A[121] ), .ZN(new_n5447_));
  NOR2_X1    g04438(.A1(new_n5447_), .A2(new_n5445_), .ZN(new_n5448_));
  INV_X1     g04439(.I(\A[126] ), .ZN(new_n5449_));
  NOR2_X1    g04440(.A1(new_n5449_), .A2(\A[125] ), .ZN(new_n5450_));
  INV_X1     g04441(.I(\A[125] ), .ZN(new_n5451_));
  NOR2_X1    g04442(.A1(new_n5451_), .A2(\A[126] ), .ZN(new_n5452_));
  OAI21_X1   g04443(.A1(new_n5450_), .A2(new_n5452_), .B(\A[124] ), .ZN(new_n5453_));
  AND2_X2    g04444(.A1(\A[125] ), .A2(\A[126] ), .Z(new_n5454_));
  OAI21_X1   g04445(.A1(new_n5454_), .A2(new_n5433_), .B(new_n5432_), .ZN(new_n5455_));
  NAND2_X1   g04446(.A1(new_n5453_), .A2(new_n5455_), .ZN(new_n5456_));
  NAND2_X1   g04447(.A1(new_n5448_), .A2(new_n5456_), .ZN(new_n5457_));
  NOR2_X1    g04448(.A1(new_n5443_), .A2(\A[122] ), .ZN(new_n5458_));
  NOR2_X1    g04449(.A1(new_n5441_), .A2(\A[123] ), .ZN(new_n5459_));
  OAI21_X1   g04450(.A1(new_n5458_), .A2(new_n5459_), .B(\A[121] ), .ZN(new_n5460_));
  INV_X1     g04451(.I(new_n5438_), .ZN(new_n5461_));
  OAI21_X1   g04452(.A1(new_n5461_), .A2(new_n5437_), .B(new_n5436_), .ZN(new_n5462_));
  NAND2_X1   g04453(.A1(new_n5460_), .A2(new_n5462_), .ZN(new_n5463_));
  NAND2_X1   g04454(.A1(new_n5451_), .A2(\A[126] ), .ZN(new_n5464_));
  NAND2_X1   g04455(.A1(new_n5449_), .A2(\A[125] ), .ZN(new_n5465_));
  AOI21_X1   g04456(.A1(new_n5464_), .A2(new_n5465_), .B(new_n5432_), .ZN(new_n5466_));
  INV_X1     g04457(.I(new_n5433_), .ZN(new_n5467_));
  AOI21_X1   g04458(.A1(new_n5467_), .A2(new_n5434_), .B(\A[124] ), .ZN(new_n5468_));
  NOR2_X1    g04459(.A1(new_n5468_), .A2(new_n5466_), .ZN(new_n5469_));
  NAND2_X1   g04460(.A1(new_n5469_), .A2(new_n5463_), .ZN(new_n5470_));
  AOI21_X1   g04461(.A1(new_n5470_), .A2(new_n5457_), .B(new_n5440_), .ZN(new_n5471_));
  INV_X1     g04462(.I(new_n5435_), .ZN(new_n5472_));
  NAND4_X1   g04463(.A1(new_n5460_), .A2(new_n5453_), .A3(new_n5462_), .A4(new_n5455_), .ZN(new_n5473_));
  NAND2_X1   g04464(.A1(new_n5473_), .A2(new_n5439_), .ZN(new_n5474_));
  INV_X1     g04465(.I(new_n5439_), .ZN(new_n5475_));
  NAND3_X1   g04466(.A1(new_n5448_), .A2(new_n5469_), .A3(new_n5475_), .ZN(new_n5476_));
  AOI21_X1   g04467(.A1(new_n5474_), .A2(new_n5476_), .B(new_n5472_), .ZN(new_n5477_));
  AOI21_X1   g04468(.A1(new_n5448_), .A2(new_n5469_), .B(new_n5475_), .ZN(new_n5478_));
  NOR3_X1    g04469(.A1(new_n5463_), .A2(new_n5456_), .A3(new_n5439_), .ZN(new_n5479_));
  NOR3_X1    g04470(.A1(new_n5478_), .A2(new_n5479_), .A3(new_n5435_), .ZN(new_n5480_));
  NOR3_X1    g04471(.A1(new_n5477_), .A2(new_n5480_), .A3(new_n5471_), .ZN(new_n5481_));
  INV_X1     g04472(.I(new_n5440_), .ZN(new_n5482_));
  NOR4_X1    g04473(.A1(new_n5445_), .A2(new_n5447_), .A3(new_n5468_), .A4(new_n5466_), .ZN(new_n5483_));
  NAND2_X1   g04474(.A1(new_n5483_), .A2(new_n5482_), .ZN(new_n5484_));
  NAND2_X1   g04475(.A1(new_n5463_), .A2(new_n5456_), .ZN(new_n5485_));
  NAND2_X1   g04476(.A1(new_n5485_), .A2(new_n5473_), .ZN(new_n5486_));
  OAI22_X1   g04477(.A1(new_n5401_), .A2(new_n5403_), .B1(new_n5410_), .B2(new_n5408_), .ZN(new_n5487_));
  NAND2_X1   g04478(.A1(new_n5487_), .A2(new_n5423_), .ZN(new_n5488_));
  NAND2_X1   g04479(.A1(new_n5391_), .A2(new_n5395_), .ZN(new_n5489_));
  INV_X1     g04480(.I(new_n5489_), .ZN(new_n5490_));
  NAND2_X1   g04481(.A1(new_n5411_), .A2(new_n5490_), .ZN(new_n5491_));
  NOR4_X1    g04482(.A1(new_n5486_), .A2(new_n5488_), .A3(new_n5484_), .A4(new_n5491_), .ZN(new_n5492_));
  NAND2_X1   g04483(.A1(new_n5481_), .A2(new_n5492_), .ZN(new_n5493_));
  NOR2_X1    g04484(.A1(new_n5469_), .A2(new_n5463_), .ZN(new_n5494_));
  NOR2_X1    g04485(.A1(new_n5448_), .A2(new_n5456_), .ZN(new_n5495_));
  OAI21_X1   g04486(.A1(new_n5494_), .A2(new_n5495_), .B(new_n5482_), .ZN(new_n5496_));
  OAI21_X1   g04487(.A1(new_n5478_), .A2(new_n5479_), .B(new_n5435_), .ZN(new_n5497_));
  NAND3_X1   g04488(.A1(new_n5474_), .A2(new_n5476_), .A3(new_n5472_), .ZN(new_n5498_));
  NAND3_X1   g04489(.A1(new_n5498_), .A2(new_n5497_), .A3(new_n5496_), .ZN(new_n5499_));
  NOR2_X1    g04490(.A1(new_n5473_), .A2(new_n5440_), .ZN(new_n5500_));
  AOI22_X1   g04491(.A1(new_n5460_), .A2(new_n5462_), .B1(new_n5453_), .B2(new_n5455_), .ZN(new_n5501_));
  NOR2_X1    g04492(.A1(new_n5483_), .A2(new_n5501_), .ZN(new_n5502_));
  AOI22_X1   g04493(.A1(new_n5415_), .A2(new_n5417_), .B1(new_n5420_), .B2(new_n5422_), .ZN(new_n5503_));
  NOR2_X1    g04494(.A1(new_n5503_), .A2(new_n5411_), .ZN(new_n5504_));
  NOR2_X1    g04495(.A1(new_n5423_), .A2(new_n5489_), .ZN(new_n5505_));
  NAND4_X1   g04496(.A1(new_n5504_), .A2(new_n5502_), .A3(new_n5505_), .A4(new_n5500_), .ZN(new_n5506_));
  NAND2_X1   g04497(.A1(new_n5499_), .A2(new_n5506_), .ZN(new_n5507_));
  AOI21_X1   g04498(.A1(new_n5493_), .A2(new_n5507_), .B(new_n5431_), .ZN(new_n5508_));
  NOR2_X1    g04499(.A1(new_n5481_), .A2(new_n5506_), .ZN(new_n5509_));
  NOR2_X1    g04500(.A1(new_n5477_), .A2(new_n5480_), .ZN(new_n5510_));
  NAND3_X1   g04501(.A1(new_n5504_), .A2(new_n5502_), .A3(new_n5500_), .ZN(new_n5511_));
  INV_X1     g04502(.I(new_n5511_), .ZN(new_n5512_));
  NAND2_X1   g04503(.A1(new_n5496_), .A2(new_n5505_), .ZN(new_n5513_));
  AOI21_X1   g04504(.A1(new_n5512_), .A2(new_n5510_), .B(new_n5513_), .ZN(new_n5514_));
  NOR3_X1    g04505(.A1(new_n5514_), .A2(new_n5509_), .A3(new_n5431_), .ZN(new_n5515_));
  NOR2_X1    g04506(.A1(new_n5515_), .A2(new_n5508_), .ZN(new_n5516_));
  AOI21_X1   g04507(.A1(new_n5427_), .A2(new_n5429_), .B(new_n5426_), .ZN(new_n5517_));
  NOR3_X1    g04508(.A1(new_n5412_), .A2(new_n5424_), .A3(new_n5391_), .ZN(new_n5518_));
  NOR2_X1    g04509(.A1(new_n5518_), .A2(new_n5517_), .ZN(new_n5519_));
  NOR4_X1    g04510(.A1(new_n5506_), .A2(new_n5471_), .A3(new_n5477_), .A4(new_n5480_), .ZN(new_n5520_));
  NOR2_X1    g04511(.A1(new_n5481_), .A2(new_n5492_), .ZN(new_n5521_));
  OAI21_X1   g04512(.A1(new_n5521_), .A2(new_n5520_), .B(new_n5519_), .ZN(new_n5522_));
  NAND2_X1   g04513(.A1(new_n5499_), .A2(new_n5492_), .ZN(new_n5523_));
  NAND2_X1   g04514(.A1(new_n5498_), .A2(new_n5497_), .ZN(new_n5524_));
  NOR2_X1    g04515(.A1(new_n5471_), .A2(new_n5491_), .ZN(new_n5525_));
  OAI21_X1   g04516(.A1(new_n5524_), .A2(new_n5511_), .B(new_n5525_), .ZN(new_n5526_));
  NAND3_X1   g04517(.A1(new_n5526_), .A2(new_n5523_), .A3(new_n5519_), .ZN(new_n5527_));
  NOR2_X1    g04518(.A1(new_n5486_), .A2(new_n5484_), .ZN(new_n5528_));
  NAND2_X1   g04519(.A1(new_n5504_), .A2(new_n5505_), .ZN(new_n5529_));
  NOR2_X1    g04520(.A1(new_n5528_), .A2(new_n5529_), .ZN(new_n5530_));
  NAND2_X1   g04521(.A1(new_n5528_), .A2(new_n5529_), .ZN(new_n5531_));
  INV_X1     g04522(.I(new_n5531_), .ZN(new_n5532_));
  INV_X1     g04523(.I(\A[111] ), .ZN(new_n5533_));
  NOR2_X1    g04524(.A1(new_n5533_), .A2(\A[110] ), .ZN(new_n5534_));
  INV_X1     g04525(.I(\A[110] ), .ZN(new_n5535_));
  NOR2_X1    g04526(.A1(new_n5535_), .A2(\A[111] ), .ZN(new_n5536_));
  OAI21_X1   g04527(.A1(new_n5534_), .A2(new_n5536_), .B(\A[109] ), .ZN(new_n5537_));
  INV_X1     g04528(.I(\A[109] ), .ZN(new_n5538_));
  NOR2_X1    g04529(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n5539_));
  NAND2_X1   g04530(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n5540_));
  INV_X1     g04531(.I(new_n5540_), .ZN(new_n5541_));
  OAI21_X1   g04532(.A1(new_n5541_), .A2(new_n5539_), .B(new_n5538_), .ZN(new_n5542_));
  NAND2_X1   g04533(.A1(new_n5537_), .A2(new_n5542_), .ZN(new_n5543_));
  INV_X1     g04534(.I(\A[114] ), .ZN(new_n5544_));
  NOR2_X1    g04535(.A1(new_n5544_), .A2(\A[113] ), .ZN(new_n5545_));
  INV_X1     g04536(.I(\A[113] ), .ZN(new_n5546_));
  NOR2_X1    g04537(.A1(new_n5546_), .A2(\A[114] ), .ZN(new_n5547_));
  OAI21_X1   g04538(.A1(new_n5545_), .A2(new_n5547_), .B(\A[112] ), .ZN(new_n5548_));
  INV_X1     g04539(.I(\A[112] ), .ZN(new_n5549_));
  NOR2_X1    g04540(.A1(\A[113] ), .A2(\A[114] ), .ZN(new_n5550_));
  AND2_X2    g04541(.A1(\A[113] ), .A2(\A[114] ), .Z(new_n5551_));
  OAI21_X1   g04542(.A1(new_n5551_), .A2(new_n5550_), .B(new_n5549_), .ZN(new_n5552_));
  NAND2_X1   g04543(.A1(new_n5548_), .A2(new_n5552_), .ZN(new_n5553_));
  NAND2_X1   g04544(.A1(\A[113] ), .A2(\A[114] ), .ZN(new_n5554_));
  AOI21_X1   g04545(.A1(new_n5549_), .A2(new_n5554_), .B(new_n5550_), .ZN(new_n5555_));
  AOI21_X1   g04546(.A1(new_n5538_), .A2(new_n5540_), .B(new_n5539_), .ZN(new_n5556_));
  NAND2_X1   g04547(.A1(new_n5555_), .A2(new_n5556_), .ZN(new_n5557_));
  NOR3_X1    g04548(.A1(new_n5543_), .A2(new_n5553_), .A3(new_n5557_), .ZN(new_n5558_));
  NOR2_X1    g04549(.A1(new_n5543_), .A2(new_n5553_), .ZN(new_n5559_));
  NAND2_X1   g04550(.A1(new_n5535_), .A2(\A[111] ), .ZN(new_n5560_));
  NAND2_X1   g04551(.A1(new_n5533_), .A2(\A[110] ), .ZN(new_n5561_));
  AOI21_X1   g04552(.A1(new_n5560_), .A2(new_n5561_), .B(new_n5538_), .ZN(new_n5562_));
  INV_X1     g04553(.I(new_n5539_), .ZN(new_n5563_));
  AOI21_X1   g04554(.A1(new_n5563_), .A2(new_n5540_), .B(\A[109] ), .ZN(new_n5564_));
  NOR2_X1    g04555(.A1(new_n5564_), .A2(new_n5562_), .ZN(new_n5565_));
  NAND2_X1   g04556(.A1(new_n5546_), .A2(\A[114] ), .ZN(new_n5566_));
  NAND2_X1   g04557(.A1(new_n5544_), .A2(\A[113] ), .ZN(new_n5567_));
  AOI21_X1   g04558(.A1(new_n5566_), .A2(new_n5567_), .B(new_n5549_), .ZN(new_n5568_));
  INV_X1     g04559(.I(new_n5550_), .ZN(new_n5569_));
  AOI21_X1   g04560(.A1(new_n5569_), .A2(new_n5554_), .B(\A[112] ), .ZN(new_n5570_));
  NOR2_X1    g04561(.A1(new_n5570_), .A2(new_n5568_), .ZN(new_n5571_));
  NOR2_X1    g04562(.A1(new_n5565_), .A2(new_n5571_), .ZN(new_n5572_));
  NOR2_X1    g04563(.A1(new_n5572_), .A2(new_n5559_), .ZN(new_n5573_));
  INV_X1     g04564(.I(\A[103] ), .ZN(new_n5574_));
  INV_X1     g04565(.I(\A[104] ), .ZN(new_n5575_));
  NAND2_X1   g04566(.A1(new_n5575_), .A2(\A[105] ), .ZN(new_n5576_));
  INV_X1     g04567(.I(\A[105] ), .ZN(new_n5577_));
  NAND2_X1   g04568(.A1(new_n5577_), .A2(\A[104] ), .ZN(new_n5578_));
  AOI21_X1   g04569(.A1(new_n5576_), .A2(new_n5578_), .B(new_n5574_), .ZN(new_n5579_));
  NOR2_X1    g04570(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n5580_));
  INV_X1     g04571(.I(new_n5580_), .ZN(new_n5581_));
  NAND2_X1   g04572(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n5582_));
  AOI21_X1   g04573(.A1(new_n5581_), .A2(new_n5582_), .B(\A[103] ), .ZN(new_n5583_));
  NOR2_X1    g04574(.A1(new_n5583_), .A2(new_n5579_), .ZN(new_n5584_));
  INV_X1     g04575(.I(\A[106] ), .ZN(new_n5585_));
  INV_X1     g04576(.I(\A[107] ), .ZN(new_n5586_));
  NAND2_X1   g04577(.A1(new_n5586_), .A2(\A[108] ), .ZN(new_n5587_));
  INV_X1     g04578(.I(\A[108] ), .ZN(new_n5588_));
  NAND2_X1   g04579(.A1(new_n5588_), .A2(\A[107] ), .ZN(new_n5589_));
  AOI21_X1   g04580(.A1(new_n5587_), .A2(new_n5589_), .B(new_n5585_), .ZN(new_n5590_));
  NOR2_X1    g04581(.A1(\A[107] ), .A2(\A[108] ), .ZN(new_n5591_));
  INV_X1     g04582(.I(new_n5591_), .ZN(new_n5592_));
  NAND2_X1   g04583(.A1(\A[107] ), .A2(\A[108] ), .ZN(new_n5593_));
  AOI21_X1   g04584(.A1(new_n5592_), .A2(new_n5593_), .B(\A[106] ), .ZN(new_n5594_));
  NOR2_X1    g04585(.A1(new_n5594_), .A2(new_n5590_), .ZN(new_n5595_));
  AOI21_X1   g04586(.A1(new_n5585_), .A2(new_n5593_), .B(new_n5591_), .ZN(new_n5596_));
  AOI21_X1   g04587(.A1(new_n5574_), .A2(new_n5582_), .B(new_n5580_), .ZN(new_n5597_));
  NAND2_X1   g04588(.A1(new_n5596_), .A2(new_n5597_), .ZN(new_n5598_));
  INV_X1     g04589(.I(new_n5598_), .ZN(new_n5599_));
  NAND2_X1   g04590(.A1(new_n5573_), .A2(new_n5558_), .ZN(new_n5600_));
  INV_X1     g04591(.I(new_n5600_), .ZN(new_n5601_));
  NOR3_X1    g04592(.A1(new_n5532_), .A2(new_n5530_), .A3(new_n5601_), .ZN(new_n5602_));
  AOI21_X1   g04593(.A1(new_n5527_), .A2(new_n5522_), .B(new_n5602_), .ZN(new_n5603_));
  INV_X1     g04594(.I(new_n5530_), .ZN(new_n5604_));
  NAND3_X1   g04595(.A1(new_n5604_), .A2(new_n5531_), .A3(new_n5600_), .ZN(new_n5605_));
  NOR3_X1    g04596(.A1(new_n5515_), .A2(new_n5508_), .A3(new_n5605_), .ZN(new_n5606_));
  INV_X1     g04597(.I(new_n5556_), .ZN(new_n5607_));
  AOI21_X1   g04598(.A1(new_n5565_), .A2(new_n5571_), .B(new_n5607_), .ZN(new_n5608_));
  NOR3_X1    g04599(.A1(new_n5543_), .A2(new_n5553_), .A3(new_n5556_), .ZN(new_n5609_));
  OAI21_X1   g04600(.A1(new_n5608_), .A2(new_n5609_), .B(new_n5555_), .ZN(new_n5610_));
  INV_X1     g04601(.I(new_n5555_), .ZN(new_n5611_));
  OAI21_X1   g04602(.A1(new_n5543_), .A2(new_n5553_), .B(new_n5556_), .ZN(new_n5612_));
  NAND3_X1   g04603(.A1(new_n5565_), .A2(new_n5571_), .A3(new_n5607_), .ZN(new_n5613_));
  NAND3_X1   g04604(.A1(new_n5613_), .A2(new_n5612_), .A3(new_n5611_), .ZN(new_n5614_));
  NAND2_X1   g04605(.A1(new_n5610_), .A2(new_n5614_), .ZN(new_n5615_));
  NOR4_X1    g04606(.A1(new_n5579_), .A2(new_n5583_), .A3(new_n5594_), .A4(new_n5590_), .ZN(new_n5616_));
  NOR2_X1    g04607(.A1(new_n5584_), .A2(new_n5595_), .ZN(new_n5617_));
  NOR2_X1    g04608(.A1(new_n5617_), .A2(new_n5616_), .ZN(new_n5618_));
  NAND3_X1   g04609(.A1(new_n5573_), .A2(new_n5618_), .A3(new_n5558_), .ZN(new_n5619_));
  NAND2_X1   g04610(.A1(new_n5584_), .A2(new_n5595_), .ZN(new_n5620_));
  NAND2_X1   g04611(.A1(new_n5565_), .A2(new_n5553_), .ZN(new_n5621_));
  NAND2_X1   g04612(.A1(new_n5571_), .A2(new_n5543_), .ZN(new_n5622_));
  AOI21_X1   g04613(.A1(new_n5622_), .A2(new_n5621_), .B(new_n5557_), .ZN(new_n5623_));
  NOR3_X1    g04614(.A1(new_n5623_), .A2(new_n5620_), .A3(new_n5598_), .ZN(new_n5624_));
  OAI21_X1   g04615(.A1(new_n5619_), .A2(new_n5615_), .B(new_n5624_), .ZN(new_n5625_));
  INV_X1     g04616(.I(new_n5596_), .ZN(new_n5626_));
  NOR2_X1    g04617(.A1(new_n5577_), .A2(\A[104] ), .ZN(new_n5627_));
  NOR2_X1    g04618(.A1(new_n5575_), .A2(\A[105] ), .ZN(new_n5628_));
  OAI21_X1   g04619(.A1(new_n5627_), .A2(new_n5628_), .B(\A[103] ), .ZN(new_n5629_));
  INV_X1     g04620(.I(new_n5582_), .ZN(new_n5630_));
  OAI21_X1   g04621(.A1(new_n5630_), .A2(new_n5580_), .B(new_n5574_), .ZN(new_n5631_));
  NAND2_X1   g04622(.A1(new_n5629_), .A2(new_n5631_), .ZN(new_n5632_));
  NOR2_X1    g04623(.A1(new_n5588_), .A2(\A[107] ), .ZN(new_n5633_));
  NOR2_X1    g04624(.A1(new_n5586_), .A2(\A[108] ), .ZN(new_n5634_));
  OAI21_X1   g04625(.A1(new_n5633_), .A2(new_n5634_), .B(\A[106] ), .ZN(new_n5635_));
  INV_X1     g04626(.I(new_n5593_), .ZN(new_n5636_));
  OAI21_X1   g04627(.A1(new_n5636_), .A2(new_n5591_), .B(new_n5585_), .ZN(new_n5637_));
  NAND2_X1   g04628(.A1(new_n5635_), .A2(new_n5637_), .ZN(new_n5638_));
  OAI21_X1   g04629(.A1(new_n5632_), .A2(new_n5638_), .B(new_n5597_), .ZN(new_n5639_));
  INV_X1     g04630(.I(new_n5597_), .ZN(new_n5640_));
  NAND3_X1   g04631(.A1(new_n5584_), .A2(new_n5595_), .A3(new_n5640_), .ZN(new_n5641_));
  AOI21_X1   g04632(.A1(new_n5639_), .A2(new_n5641_), .B(new_n5626_), .ZN(new_n5642_));
  AOI21_X1   g04633(.A1(new_n5584_), .A2(new_n5595_), .B(new_n5640_), .ZN(new_n5643_));
  NOR3_X1    g04634(.A1(new_n5632_), .A2(new_n5638_), .A3(new_n5597_), .ZN(new_n5644_));
  NOR3_X1    g04635(.A1(new_n5643_), .A2(new_n5644_), .A3(new_n5596_), .ZN(new_n5645_));
  NOR2_X1    g04636(.A1(new_n5645_), .A2(new_n5642_), .ZN(new_n5646_));
  NOR2_X1    g04637(.A1(new_n5625_), .A2(new_n5646_), .ZN(new_n5647_));
  OAI21_X1   g04638(.A1(new_n5643_), .A2(new_n5644_), .B(new_n5596_), .ZN(new_n5648_));
  NAND3_X1   g04639(.A1(new_n5639_), .A2(new_n5641_), .A3(new_n5626_), .ZN(new_n5649_));
  NAND2_X1   g04640(.A1(new_n5648_), .A2(new_n5649_), .ZN(new_n5650_));
  NOR3_X1    g04641(.A1(new_n5632_), .A2(new_n5638_), .A3(new_n5598_), .ZN(new_n5651_));
  NAND4_X1   g04642(.A1(new_n5573_), .A2(new_n5618_), .A3(new_n5558_), .A4(new_n5651_), .ZN(new_n5652_));
  NAND2_X1   g04643(.A1(new_n5650_), .A2(new_n5652_), .ZN(new_n5653_));
  INV_X1     g04644(.I(new_n5557_), .ZN(new_n5654_));
  NOR2_X1    g04645(.A1(new_n5571_), .A2(new_n5543_), .ZN(new_n5655_));
  NOR2_X1    g04646(.A1(new_n5565_), .A2(new_n5553_), .ZN(new_n5656_));
  OAI21_X1   g04647(.A1(new_n5655_), .A2(new_n5656_), .B(new_n5654_), .ZN(new_n5657_));
  NAND3_X1   g04648(.A1(new_n5610_), .A2(new_n5614_), .A3(new_n5657_), .ZN(new_n5658_));
  OAI21_X1   g04649(.A1(new_n5650_), .A2(new_n5652_), .B(new_n5658_), .ZN(new_n5659_));
  AOI21_X1   g04650(.A1(new_n5613_), .A2(new_n5612_), .B(new_n5611_), .ZN(new_n5660_));
  NOR3_X1    g04651(.A1(new_n5608_), .A2(new_n5609_), .A3(new_n5555_), .ZN(new_n5661_));
  NOR3_X1    g04652(.A1(new_n5661_), .A2(new_n5660_), .A3(new_n5623_), .ZN(new_n5662_));
  NAND2_X1   g04653(.A1(new_n5565_), .A2(new_n5571_), .ZN(new_n5663_));
  NAND2_X1   g04654(.A1(new_n5543_), .A2(new_n5553_), .ZN(new_n5664_));
  NAND3_X1   g04655(.A1(new_n5558_), .A2(new_n5663_), .A3(new_n5664_), .ZN(new_n5665_));
  NAND2_X1   g04656(.A1(new_n5632_), .A2(new_n5638_), .ZN(new_n5666_));
  NAND3_X1   g04657(.A1(new_n5651_), .A2(new_n5620_), .A3(new_n5666_), .ZN(new_n5667_));
  NOR4_X1    g04658(.A1(new_n5642_), .A2(new_n5645_), .A3(new_n5667_), .A4(new_n5665_), .ZN(new_n5668_));
  NAND2_X1   g04659(.A1(new_n5668_), .A2(new_n5662_), .ZN(new_n5669_));
  NAND2_X1   g04660(.A1(new_n5659_), .A2(new_n5669_), .ZN(new_n5670_));
  AOI21_X1   g04661(.A1(new_n5670_), .A2(new_n5653_), .B(new_n5647_), .ZN(new_n5671_));
  OAI22_X1   g04662(.A1(new_n5603_), .A2(new_n5606_), .B1(new_n5671_), .B2(new_n5516_), .ZN(new_n5672_));
  AOI21_X1   g04663(.A1(new_n5499_), .A2(new_n5492_), .B(new_n5519_), .ZN(new_n5673_));
  NAND2_X1   g04664(.A1(new_n5475_), .A2(new_n5472_), .ZN(new_n5674_));
  AOI21_X1   g04665(.A1(new_n5483_), .A2(new_n5674_), .B(new_n5482_), .ZN(new_n5675_));
  NAND2_X1   g04666(.A1(new_n5426_), .A2(new_n5396_), .ZN(new_n5676_));
  AOI21_X1   g04667(.A1(new_n5411_), .A2(new_n5676_), .B(new_n5490_), .ZN(new_n5677_));
  XOR2_X1    g04668(.A1(new_n5675_), .A2(new_n5677_), .Z(new_n5678_));
  NOR3_X1    g04669(.A1(new_n5673_), .A2(new_n5514_), .A3(new_n5678_), .ZN(new_n5679_));
  OAI21_X1   g04670(.A1(new_n5662_), .A2(new_n5652_), .B(new_n5650_), .ZN(new_n5680_));
  NOR2_X1    g04671(.A1(new_n5555_), .A2(new_n5556_), .ZN(new_n5681_));
  OAI21_X1   g04672(.A1(new_n5663_), .A2(new_n5681_), .B(new_n5557_), .ZN(new_n5682_));
  NAND2_X1   g04673(.A1(new_n5626_), .A2(new_n5640_), .ZN(new_n5683_));
  AOI21_X1   g04674(.A1(new_n5616_), .A2(new_n5683_), .B(new_n5599_), .ZN(new_n5684_));
  XOR2_X1    g04675(.A1(new_n5682_), .A2(new_n5684_), .Z(new_n5685_));
  NAND3_X1   g04676(.A1(new_n5680_), .A2(new_n5625_), .A3(new_n5685_), .ZN(new_n5686_));
  XOR2_X1    g04677(.A1(new_n5679_), .A2(new_n5686_), .Z(new_n5687_));
  NOR2_X1    g04678(.A1(new_n5672_), .A2(new_n5687_), .ZN(new_n5688_));
  NAND2_X1   g04679(.A1(new_n5527_), .A2(new_n5522_), .ZN(new_n5689_));
  OAI21_X1   g04680(.A1(new_n5515_), .A2(new_n5508_), .B(new_n5605_), .ZN(new_n5690_));
  NAND3_X1   g04681(.A1(new_n5527_), .A2(new_n5522_), .A3(new_n5602_), .ZN(new_n5691_));
  NOR2_X1    g04682(.A1(new_n5661_), .A2(new_n5660_), .ZN(new_n5692_));
  NOR3_X1    g04683(.A1(new_n5665_), .A2(new_n5616_), .A3(new_n5617_), .ZN(new_n5693_));
  NAND2_X1   g04684(.A1(new_n5657_), .A2(new_n5651_), .ZN(new_n5694_));
  AOI21_X1   g04685(.A1(new_n5692_), .A2(new_n5693_), .B(new_n5694_), .ZN(new_n5695_));
  NAND2_X1   g04686(.A1(new_n5695_), .A2(new_n5650_), .ZN(new_n5696_));
  NOR2_X1    g04687(.A1(new_n5668_), .A2(new_n5662_), .ZN(new_n5697_));
  NOR3_X1    g04688(.A1(new_n5658_), .A2(new_n5650_), .A3(new_n5652_), .ZN(new_n5698_));
  OAI21_X1   g04689(.A1(new_n5697_), .A2(new_n5698_), .B(new_n5653_), .ZN(new_n5699_));
  NAND2_X1   g04690(.A1(new_n5699_), .A2(new_n5696_), .ZN(new_n5700_));
  AOI22_X1   g04691(.A1(new_n5690_), .A2(new_n5691_), .B1(new_n5700_), .B2(new_n5689_), .ZN(new_n5701_));
  INV_X1     g04692(.I(new_n5652_), .ZN(new_n5702_));
  AOI21_X1   g04693(.A1(new_n5702_), .A2(new_n5658_), .B(new_n5646_), .ZN(new_n5703_));
  XNOR2_X1   g04694(.A1(new_n5682_), .A2(new_n5684_), .ZN(new_n5704_));
  NOR3_X1    g04695(.A1(new_n5703_), .A2(new_n5695_), .A3(new_n5704_), .ZN(new_n5705_));
  NOR2_X1    g04696(.A1(new_n5705_), .A2(new_n5679_), .ZN(new_n5706_));
  OAI21_X1   g04697(.A1(new_n5481_), .A2(new_n5506_), .B(new_n5431_), .ZN(new_n5707_));
  INV_X1     g04698(.I(new_n5678_), .ZN(new_n5708_));
  NAND3_X1   g04699(.A1(new_n5707_), .A2(new_n5708_), .A3(new_n5526_), .ZN(new_n5709_));
  NOR2_X1    g04700(.A1(new_n5709_), .A2(new_n5686_), .ZN(new_n5710_));
  NOR2_X1    g04701(.A1(new_n5706_), .A2(new_n5710_), .ZN(new_n5711_));
  NOR2_X1    g04702(.A1(new_n5701_), .A2(new_n5711_), .ZN(new_n5712_));
  NOR4_X1    g04703(.A1(new_n5368_), .A2(new_n5387_), .A3(new_n5688_), .A4(new_n5712_), .ZN(new_n5713_));
  NOR3_X1    g04704(.A1(new_n5603_), .A2(new_n5606_), .A3(new_n5700_), .ZN(new_n5714_));
  INV_X1     g04705(.I(new_n5714_), .ZN(new_n5715_));
  OAI21_X1   g04706(.A1(new_n5532_), .A2(new_n5530_), .B(new_n5601_), .ZN(new_n5716_));
  NOR2_X1    g04707(.A1(new_n5282_), .A2(new_n5276_), .ZN(new_n5717_));
  NOR2_X1    g04708(.A1(new_n5717_), .A2(new_n5278_), .ZN(new_n5718_));
  NAND3_X1   g04709(.A1(new_n5718_), .A2(new_n5605_), .A3(new_n5716_), .ZN(new_n5719_));
  NAND2_X1   g04710(.A1(new_n5715_), .A2(new_n5719_), .ZN(new_n5720_));
  INV_X1     g04711(.I(new_n5719_), .ZN(new_n5721_));
  NAND2_X1   g04712(.A1(new_n5721_), .A2(new_n5714_), .ZN(new_n5722_));
  OAI21_X1   g04713(.A1(new_n5284_), .A2(new_n5279_), .B(new_n5351_), .ZN(new_n5723_));
  NAND3_X1   g04714(.A1(new_n5370_), .A2(new_n5371_), .A3(new_n5380_), .ZN(new_n5724_));
  NAND2_X1   g04715(.A1(new_n5723_), .A2(new_n5724_), .ZN(new_n5725_));
  AOI22_X1   g04716(.A1(new_n5720_), .A2(new_n5722_), .B1(new_n5715_), .B2(new_n5725_), .ZN(new_n5726_));
  OAI22_X1   g04717(.A1(new_n5368_), .A2(new_n5387_), .B1(new_n5688_), .B2(new_n5712_), .ZN(new_n5727_));
  AOI21_X1   g04718(.A1(new_n5726_), .A2(new_n5727_), .B(new_n5713_), .ZN(new_n5728_));
  INV_X1     g04719(.I(new_n5355_), .ZN(new_n5729_));
  NAND2_X1   g04720(.A1(new_n5729_), .A2(new_n5357_), .ZN(new_n5730_));
  AOI21_X1   g04721(.A1(new_n5109_), .A2(new_n5197_), .B(new_n5190_), .ZN(new_n5731_));
  OAI21_X1   g04722(.A1(new_n5729_), .A2(new_n5357_), .B(new_n5731_), .ZN(new_n5732_));
  NAND2_X1   g04723(.A1(new_n5732_), .A2(new_n5730_), .ZN(new_n5733_));
  AND2_X2    g04724(.A1(new_n5360_), .A2(new_n5306_), .Z(new_n5734_));
  INV_X1     g04725(.I(new_n5362_), .ZN(new_n5735_));
  INV_X1     g04726(.I(new_n5364_), .ZN(new_n5736_));
  NOR2_X1    g04727(.A1(new_n5736_), .A2(new_n5735_), .ZN(new_n5737_));
  NAND2_X1   g04728(.A1(new_n5736_), .A2(new_n5735_), .ZN(new_n5738_));
  AOI21_X1   g04729(.A1(new_n5734_), .A2(new_n5738_), .B(new_n5737_), .ZN(new_n5739_));
  NAND2_X1   g04730(.A1(new_n5359_), .A2(new_n5366_), .ZN(new_n5740_));
  INV_X1     g04731(.I(new_n5385_), .ZN(new_n5741_));
  AOI21_X1   g04732(.A1(new_n5352_), .A2(new_n5740_), .B(new_n5741_), .ZN(new_n5742_));
  NOR2_X1    g04733(.A1(new_n5742_), .A2(new_n5739_), .ZN(new_n5743_));
  NAND4_X1   g04734(.A1(new_n5381_), .A2(new_n5382_), .A3(new_n5383_), .A4(new_n5739_), .ZN(new_n5744_));
  INV_X1     g04735(.I(new_n5744_), .ZN(new_n5745_));
  OAI21_X1   g04736(.A1(new_n5743_), .A2(new_n5745_), .B(new_n5733_), .ZN(new_n5746_));
  INV_X1     g04737(.I(new_n5733_), .ZN(new_n5747_));
  INV_X1     g04738(.I(new_n5739_), .ZN(new_n5748_));
  NAND3_X1   g04739(.A1(new_n5381_), .A2(new_n5382_), .A3(new_n5383_), .ZN(new_n5749_));
  NAND2_X1   g04740(.A1(new_n5749_), .A2(new_n5748_), .ZN(new_n5750_));
  NAND3_X1   g04741(.A1(new_n5750_), .A2(new_n5747_), .A3(new_n5744_), .ZN(new_n5751_));
  NAND2_X1   g04742(.A1(new_n5746_), .A2(new_n5751_), .ZN(new_n5752_));
  OR2_X2     g04743(.A1(new_n5675_), .A2(new_n5677_), .Z(new_n5753_));
  NAND2_X1   g04744(.A1(new_n5675_), .A2(new_n5677_), .ZN(new_n5754_));
  NAND3_X1   g04745(.A1(new_n5707_), .A2(new_n5526_), .A3(new_n5754_), .ZN(new_n5755_));
  NAND2_X1   g04746(.A1(new_n5755_), .A2(new_n5753_), .ZN(new_n5756_));
  INV_X1     g04747(.I(new_n5756_), .ZN(new_n5757_));
  NAND3_X1   g04748(.A1(new_n5701_), .A2(new_n5679_), .A3(new_n5705_), .ZN(new_n5758_));
  INV_X1     g04749(.I(new_n5684_), .ZN(new_n5759_));
  NAND2_X1   g04750(.A1(new_n5759_), .A2(new_n5682_), .ZN(new_n5760_));
  OR2_X2     g04751(.A1(new_n5759_), .A2(new_n5682_), .Z(new_n5761_));
  NAND3_X1   g04752(.A1(new_n5680_), .A2(new_n5625_), .A3(new_n5761_), .ZN(new_n5762_));
  NAND2_X1   g04753(.A1(new_n5762_), .A2(new_n5760_), .ZN(new_n5763_));
  NAND2_X1   g04754(.A1(new_n5758_), .A2(new_n5763_), .ZN(new_n5764_));
  INV_X1     g04755(.I(new_n5763_), .ZN(new_n5765_));
  NAND4_X1   g04756(.A1(new_n5701_), .A2(new_n5765_), .A3(new_n5679_), .A4(new_n5705_), .ZN(new_n5766_));
  AOI21_X1   g04757(.A1(new_n5764_), .A2(new_n5766_), .B(new_n5757_), .ZN(new_n5767_));
  NAND2_X1   g04758(.A1(new_n5709_), .A2(new_n5686_), .ZN(new_n5768_));
  NAND2_X1   g04759(.A1(new_n5672_), .A2(new_n5768_), .ZN(new_n5769_));
  AOI21_X1   g04760(.A1(new_n5769_), .A2(new_n5710_), .B(new_n5765_), .ZN(new_n5770_));
  INV_X1     g04761(.I(new_n5766_), .ZN(new_n5771_));
  NOR3_X1    g04762(.A1(new_n5770_), .A2(new_n5771_), .A3(new_n5756_), .ZN(new_n5772_));
  NOR2_X1    g04763(.A1(new_n5772_), .A2(new_n5767_), .ZN(new_n5773_));
  NAND2_X1   g04764(.A1(new_n5752_), .A2(new_n5773_), .ZN(new_n5774_));
  AOI21_X1   g04765(.A1(new_n5750_), .A2(new_n5744_), .B(new_n5747_), .ZN(new_n5775_));
  NOR3_X1    g04766(.A1(new_n5743_), .A2(new_n5745_), .A3(new_n5733_), .ZN(new_n5776_));
  NOR2_X1    g04767(.A1(new_n5776_), .A2(new_n5775_), .ZN(new_n5777_));
  OAI21_X1   g04768(.A1(new_n5770_), .A2(new_n5771_), .B(new_n5756_), .ZN(new_n5778_));
  NAND3_X1   g04769(.A1(new_n5764_), .A2(new_n5757_), .A3(new_n5766_), .ZN(new_n5779_));
  NAND2_X1   g04770(.A1(new_n5778_), .A2(new_n5779_), .ZN(new_n5780_));
  NAND2_X1   g04771(.A1(new_n5777_), .A2(new_n5780_), .ZN(new_n5781_));
  AOI21_X1   g04772(.A1(new_n5774_), .A2(new_n5781_), .B(new_n5728_), .ZN(new_n5782_));
  XOR2_X1    g04773(.A1(new_n5359_), .A2(new_n5366_), .Z(new_n5783_));
  NAND2_X1   g04774(.A1(new_n5381_), .A2(new_n5783_), .ZN(new_n5784_));
  NAND2_X1   g04775(.A1(new_n5741_), .A2(new_n5740_), .ZN(new_n5785_));
  NAND2_X1   g04776(.A1(new_n5785_), .A2(new_n5352_), .ZN(new_n5786_));
  XOR2_X1    g04777(.A1(new_n5709_), .A2(new_n5686_), .Z(new_n5787_));
  NAND2_X1   g04778(.A1(new_n5701_), .A2(new_n5787_), .ZN(new_n5788_));
  INV_X1     g04779(.I(new_n5710_), .ZN(new_n5789_));
  NAND2_X1   g04780(.A1(new_n5789_), .A2(new_n5768_), .ZN(new_n5790_));
  NAND2_X1   g04781(.A1(new_n5790_), .A2(new_n5672_), .ZN(new_n5791_));
  NAND4_X1   g04782(.A1(new_n5786_), .A2(new_n5791_), .A3(new_n5784_), .A4(new_n5788_), .ZN(new_n5792_));
  NOR2_X1    g04783(.A1(new_n5721_), .A2(new_n5714_), .ZN(new_n5793_));
  NOR2_X1    g04784(.A1(new_n5715_), .A2(new_n5719_), .ZN(new_n5794_));
  AOI21_X1   g04785(.A1(new_n5370_), .A2(new_n5371_), .B(new_n5380_), .ZN(new_n5795_));
  NOR3_X1    g04786(.A1(new_n5279_), .A2(new_n5284_), .A3(new_n5351_), .ZN(new_n5796_));
  NOR2_X1    g04787(.A1(new_n5796_), .A2(new_n5795_), .ZN(new_n5797_));
  OAI22_X1   g04788(.A1(new_n5794_), .A2(new_n5793_), .B1(new_n5797_), .B2(new_n5714_), .ZN(new_n5798_));
  AOI22_X1   g04789(.A1(new_n5786_), .A2(new_n5784_), .B1(new_n5791_), .B2(new_n5788_), .ZN(new_n5799_));
  OAI21_X1   g04790(.A1(new_n5798_), .A2(new_n5799_), .B(new_n5792_), .ZN(new_n5800_));
  NAND4_X1   g04791(.A1(new_n5746_), .A2(new_n5778_), .A3(new_n5751_), .A4(new_n5779_), .ZN(new_n5801_));
  NAND2_X1   g04792(.A1(new_n5752_), .A2(new_n5780_), .ZN(new_n5802_));
  AOI21_X1   g04793(.A1(new_n5802_), .A2(new_n5801_), .B(new_n5800_), .ZN(new_n5803_));
  NOR4_X1    g04794(.A1(new_n5782_), .A2(new_n5043_), .A3(new_n5066_), .A4(new_n5803_), .ZN(new_n5804_));
  NAND2_X1   g04795(.A1(new_n5786_), .A2(new_n5784_), .ZN(new_n5805_));
  NOR2_X1    g04796(.A1(new_n5688_), .A2(new_n5712_), .ZN(new_n5806_));
  NOR2_X1    g04797(.A1(new_n5805_), .A2(new_n5806_), .ZN(new_n5807_));
  NOR2_X1    g04798(.A1(new_n5368_), .A2(new_n5387_), .ZN(new_n5808_));
  NAND2_X1   g04799(.A1(new_n5791_), .A2(new_n5788_), .ZN(new_n5809_));
  NOR2_X1    g04800(.A1(new_n5808_), .A2(new_n5809_), .ZN(new_n5810_));
  OAI21_X1   g04801(.A1(new_n5810_), .A2(new_n5807_), .B(new_n5726_), .ZN(new_n5811_));
  AOI21_X1   g04802(.A1(new_n5792_), .A2(new_n5727_), .B(new_n5726_), .ZN(new_n5812_));
  INV_X1     g04803(.I(new_n5812_), .ZN(new_n5813_));
  NAND2_X1   g04804(.A1(new_n5045_), .A2(new_n5047_), .ZN(new_n5814_));
  NOR2_X1    g04805(.A1(new_n4953_), .A2(new_n4973_), .ZN(new_n5815_));
  NOR2_X1    g04806(.A1(new_n5814_), .A2(new_n5815_), .ZN(new_n5816_));
  NOR2_X1    g04807(.A1(new_n4629_), .A2(new_n4649_), .ZN(new_n5817_));
  NAND2_X1   g04808(.A1(new_n5049_), .A2(new_n5052_), .ZN(new_n5818_));
  NOR2_X1    g04809(.A1(new_n5817_), .A2(new_n5818_), .ZN(new_n5819_));
  OAI21_X1   g04810(.A1(new_n5819_), .A2(new_n5816_), .B(new_n4987_), .ZN(new_n5820_));
  AOI21_X1   g04811(.A1(new_n4988_), .A2(new_n5053_), .B(new_n4987_), .ZN(new_n5821_));
  INV_X1     g04812(.I(new_n5821_), .ZN(new_n5822_));
  NAND4_X1   g04813(.A1(new_n5813_), .A2(new_n5822_), .A3(new_n5811_), .A4(new_n5820_), .ZN(new_n5823_));
  NAND3_X1   g04814(.A1(new_n4981_), .A2(new_n5060_), .A3(new_n4983_), .ZN(new_n5824_));
  NAND2_X1   g04815(.A1(new_n4542_), .A2(new_n4979_), .ZN(new_n5825_));
  OAI21_X1   g04816(.A1(new_n4863_), .A2(new_n4977_), .B(new_n5825_), .ZN(new_n5826_));
  NAND2_X1   g04817(.A1(new_n5826_), .A2(new_n4980_), .ZN(new_n5827_));
  NAND2_X1   g04818(.A1(new_n5716_), .A2(new_n5605_), .ZN(new_n5828_));
  OAI21_X1   g04819(.A1(new_n5278_), .A2(new_n5717_), .B(new_n5828_), .ZN(new_n5829_));
  NAND2_X1   g04820(.A1(new_n5719_), .A2(new_n5829_), .ZN(new_n5830_));
  NOR2_X1    g04821(.A1(new_n5827_), .A2(new_n5830_), .ZN(new_n5831_));
  INV_X1     g04822(.I(new_n5831_), .ZN(new_n5832_));
  NAND2_X1   g04823(.A1(new_n5824_), .A2(new_n5832_), .ZN(new_n5833_));
  NAND4_X1   g04824(.A1(new_n5831_), .A2(new_n4981_), .A3(new_n4983_), .A4(new_n5060_), .ZN(new_n5834_));
  NAND2_X1   g04825(.A1(new_n5720_), .A2(new_n5722_), .ZN(new_n5835_));
  XOR2_X1    g04826(.A1(new_n5835_), .A2(new_n5725_), .Z(new_n5836_));
  AOI22_X1   g04827(.A1(new_n5836_), .A2(new_n5824_), .B1(new_n5833_), .B2(new_n5834_), .ZN(new_n5837_));
  INV_X1     g04828(.I(new_n5837_), .ZN(new_n5838_));
  AOI22_X1   g04829(.A1(new_n5813_), .A2(new_n5811_), .B1(new_n5822_), .B2(new_n5820_), .ZN(new_n5839_));
  OAI21_X1   g04830(.A1(new_n5838_), .A2(new_n5839_), .B(new_n5823_), .ZN(new_n5840_));
  OAI22_X1   g04831(.A1(new_n5043_), .A2(new_n5066_), .B1(new_n5782_), .B2(new_n5803_), .ZN(new_n5841_));
  AOI21_X1   g04832(.A1(new_n5841_), .A2(new_n5840_), .B(new_n5804_), .ZN(new_n5842_));
  NAND2_X1   g04833(.A1(new_n5019_), .A2(new_n5026_), .ZN(new_n5843_));
  INV_X1     g04834(.I(new_n5020_), .ZN(new_n5844_));
  OAI21_X1   g04835(.A1(new_n5019_), .A2(new_n5026_), .B(new_n5844_), .ZN(new_n5845_));
  NAND2_X1   g04836(.A1(new_n5845_), .A2(new_n5843_), .ZN(new_n5846_));
  INV_X1     g04837(.I(new_n5846_), .ZN(new_n5847_));
  OAI21_X1   g04838(.A1(new_n5013_), .A2(new_n5041_), .B(new_n4989_), .ZN(new_n5848_));
  XNOR2_X1   g04839(.A1(new_n4994_), .A2(new_n5000_), .ZN(new_n5849_));
  XOR2_X1    g04840(.A1(new_n5018_), .A2(new_n5024_), .Z(new_n5850_));
  NOR4_X1    g04841(.A1(new_n5849_), .A2(new_n5850_), .A3(new_n5010_), .A4(new_n5020_), .ZN(new_n5851_));
  NAND2_X1   g04842(.A1(new_n5008_), .A2(new_n5000_), .ZN(new_n5852_));
  NAND2_X1   g04843(.A1(new_n5009_), .A2(new_n4994_), .ZN(new_n5853_));
  NAND2_X1   g04844(.A1(new_n5853_), .A2(new_n5003_), .ZN(new_n5854_));
  NAND2_X1   g04845(.A1(new_n5854_), .A2(new_n5852_), .ZN(new_n5855_));
  AOI21_X1   g04846(.A1(new_n5848_), .A2(new_n5851_), .B(new_n5855_), .ZN(new_n5856_));
  AOI21_X1   g04847(.A1(new_n5038_), .A2(new_n5034_), .B(new_n5063_), .ZN(new_n5857_));
  INV_X1     g04848(.I(new_n5851_), .ZN(new_n5858_));
  INV_X1     g04849(.I(new_n5855_), .ZN(new_n5859_));
  NOR3_X1    g04850(.A1(new_n5857_), .A2(new_n5858_), .A3(new_n5859_), .ZN(new_n5860_));
  OAI21_X1   g04851(.A1(new_n5860_), .A2(new_n5856_), .B(new_n5847_), .ZN(new_n5861_));
  OAI21_X1   g04852(.A1(new_n5857_), .A2(new_n5858_), .B(new_n5859_), .ZN(new_n5862_));
  NAND3_X1   g04853(.A1(new_n5848_), .A2(new_n5851_), .A3(new_n5855_), .ZN(new_n5863_));
  NAND3_X1   g04854(.A1(new_n5862_), .A2(new_n5863_), .A3(new_n5846_), .ZN(new_n5864_));
  NAND2_X1   g04855(.A1(new_n5861_), .A2(new_n5864_), .ZN(new_n5865_));
  NAND2_X1   g04856(.A1(new_n5757_), .A2(new_n5765_), .ZN(new_n5866_));
  INV_X1     g04857(.I(new_n5758_), .ZN(new_n5867_));
  OAI21_X1   g04858(.A1(new_n5757_), .A2(new_n5765_), .B(new_n5867_), .ZN(new_n5868_));
  NAND2_X1   g04859(.A1(new_n5868_), .A2(new_n5866_), .ZN(new_n5869_));
  AOI21_X1   g04860(.A1(new_n5777_), .A2(new_n5773_), .B(new_n5800_), .ZN(new_n5870_));
  XOR2_X1    g04861(.A1(new_n5733_), .A2(new_n5739_), .Z(new_n5871_));
  INV_X1     g04862(.I(new_n5871_), .ZN(new_n5872_));
  XOR2_X1    g04863(.A1(new_n5756_), .A2(new_n5763_), .Z(new_n5873_));
  NOR4_X1    g04864(.A1(new_n5872_), .A2(new_n5873_), .A3(new_n5749_), .A4(new_n5758_), .ZN(new_n5874_));
  INV_X1     g04865(.I(new_n5874_), .ZN(new_n5875_));
  NAND2_X1   g04866(.A1(new_n5747_), .A2(new_n5739_), .ZN(new_n5876_));
  NAND2_X1   g04867(.A1(new_n5733_), .A2(new_n5748_), .ZN(new_n5877_));
  NAND2_X1   g04868(.A1(new_n5742_), .A2(new_n5877_), .ZN(new_n5878_));
  NAND2_X1   g04869(.A1(new_n5878_), .A2(new_n5876_), .ZN(new_n5879_));
  INV_X1     g04870(.I(new_n5879_), .ZN(new_n5880_));
  OAI21_X1   g04871(.A1(new_n5870_), .A2(new_n5875_), .B(new_n5880_), .ZN(new_n5881_));
  OAI21_X1   g04872(.A1(new_n5752_), .A2(new_n5780_), .B(new_n5728_), .ZN(new_n5882_));
  NAND3_X1   g04873(.A1(new_n5882_), .A2(new_n5874_), .A3(new_n5879_), .ZN(new_n5883_));
  AOI21_X1   g04874(.A1(new_n5881_), .A2(new_n5883_), .B(new_n5869_), .ZN(new_n5884_));
  INV_X1     g04875(.I(new_n5869_), .ZN(new_n5885_));
  AOI21_X1   g04876(.A1(new_n5882_), .A2(new_n5874_), .B(new_n5879_), .ZN(new_n5886_));
  NOR3_X1    g04877(.A1(new_n5870_), .A2(new_n5875_), .A3(new_n5880_), .ZN(new_n5887_));
  NOR3_X1    g04878(.A1(new_n5887_), .A2(new_n5886_), .A3(new_n5885_), .ZN(new_n5888_));
  NOR2_X1    g04879(.A1(new_n5888_), .A2(new_n5884_), .ZN(new_n5889_));
  NAND2_X1   g04880(.A1(new_n5889_), .A2(new_n5865_), .ZN(new_n5890_));
  AOI21_X1   g04881(.A1(new_n5862_), .A2(new_n5863_), .B(new_n5846_), .ZN(new_n5891_));
  NOR3_X1    g04882(.A1(new_n5860_), .A2(new_n5856_), .A3(new_n5847_), .ZN(new_n5892_));
  NOR2_X1    g04883(.A1(new_n5892_), .A2(new_n5891_), .ZN(new_n5893_));
  OAI21_X1   g04884(.A1(new_n5887_), .A2(new_n5886_), .B(new_n5885_), .ZN(new_n5894_));
  NAND3_X1   g04885(.A1(new_n5881_), .A2(new_n5883_), .A3(new_n5869_), .ZN(new_n5895_));
  NAND2_X1   g04886(.A1(new_n5894_), .A2(new_n5895_), .ZN(new_n5896_));
  NAND2_X1   g04887(.A1(new_n5893_), .A2(new_n5896_), .ZN(new_n5897_));
  AOI21_X1   g04888(.A1(new_n5897_), .A2(new_n5890_), .B(new_n5842_), .ZN(new_n5898_));
  NOR2_X1    g04889(.A1(new_n5038_), .A2(new_n5041_), .ZN(new_n5899_));
  NOR2_X1    g04890(.A1(new_n5013_), .A2(new_n5034_), .ZN(new_n5900_));
  OAI21_X1   g04891(.A1(new_n5900_), .A2(new_n5899_), .B(new_n5063_), .ZN(new_n5901_));
  NOR2_X1    g04892(.A1(new_n5013_), .A2(new_n5041_), .ZN(new_n5902_));
  AOI22_X1   g04893(.A1(new_n5007_), .A2(new_n5012_), .B1(new_n5039_), .B2(new_n5040_), .ZN(new_n5903_));
  OAI21_X1   g04894(.A1(new_n5902_), .A2(new_n5903_), .B(new_n4989_), .ZN(new_n5904_));
  NOR2_X1    g04895(.A1(new_n5777_), .A2(new_n5780_), .ZN(new_n5905_));
  NOR2_X1    g04896(.A1(new_n5752_), .A2(new_n5773_), .ZN(new_n5906_));
  OAI21_X1   g04897(.A1(new_n5906_), .A2(new_n5905_), .B(new_n5800_), .ZN(new_n5907_));
  INV_X1     g04898(.I(new_n5801_), .ZN(new_n5908_));
  NOR2_X1    g04899(.A1(new_n5777_), .A2(new_n5773_), .ZN(new_n5909_));
  OAI21_X1   g04900(.A1(new_n5908_), .A2(new_n5909_), .B(new_n5728_), .ZN(new_n5910_));
  NAND4_X1   g04901(.A1(new_n5907_), .A2(new_n5910_), .A3(new_n5901_), .A4(new_n5904_), .ZN(new_n5911_));
  INV_X1     g04902(.I(new_n5811_), .ZN(new_n5912_));
  INV_X1     g04903(.I(new_n5820_), .ZN(new_n5913_));
  NOR4_X1    g04904(.A1(new_n5912_), .A2(new_n5913_), .A3(new_n5812_), .A4(new_n5821_), .ZN(new_n5914_));
  NAND2_X1   g04905(.A1(new_n5813_), .A2(new_n5811_), .ZN(new_n5915_));
  NAND2_X1   g04906(.A1(new_n5822_), .A2(new_n5820_), .ZN(new_n5916_));
  NAND2_X1   g04907(.A1(new_n5915_), .A2(new_n5916_), .ZN(new_n5917_));
  AOI21_X1   g04908(.A1(new_n5917_), .A2(new_n5837_), .B(new_n5914_), .ZN(new_n5918_));
  AOI22_X1   g04909(.A1(new_n5910_), .A2(new_n5907_), .B1(new_n5901_), .B2(new_n5904_), .ZN(new_n5919_));
  OAI21_X1   g04910(.A1(new_n5919_), .A2(new_n5918_), .B(new_n5911_), .ZN(new_n5920_));
  NAND4_X1   g04911(.A1(new_n5861_), .A2(new_n5894_), .A3(new_n5895_), .A4(new_n5864_), .ZN(new_n5921_));
  NAND2_X1   g04912(.A1(new_n5896_), .A2(new_n5865_), .ZN(new_n5922_));
  AOI21_X1   g04913(.A1(new_n5922_), .A2(new_n5921_), .B(new_n5920_), .ZN(new_n5923_));
  INV_X1     g04914(.I(\A[238] ), .ZN(new_n5924_));
  NOR2_X1    g04915(.A1(\A[239] ), .A2(\A[240] ), .ZN(new_n5925_));
  NAND2_X1   g04916(.A1(\A[239] ), .A2(\A[240] ), .ZN(new_n5926_));
  AOI21_X1   g04917(.A1(new_n5924_), .A2(new_n5926_), .B(new_n5925_), .ZN(new_n5927_));
  INV_X1     g04918(.I(\A[235] ), .ZN(new_n5928_));
  NOR2_X1    g04919(.A1(\A[236] ), .A2(\A[237] ), .ZN(new_n5929_));
  NAND2_X1   g04920(.A1(\A[236] ), .A2(\A[237] ), .ZN(new_n5930_));
  AOI21_X1   g04921(.A1(new_n5928_), .A2(new_n5930_), .B(new_n5929_), .ZN(new_n5931_));
  INV_X1     g04922(.I(new_n5931_), .ZN(new_n5932_));
  INV_X1     g04923(.I(\A[236] ), .ZN(new_n5933_));
  NAND2_X1   g04924(.A1(new_n5933_), .A2(\A[237] ), .ZN(new_n5934_));
  INV_X1     g04925(.I(\A[237] ), .ZN(new_n5935_));
  NAND2_X1   g04926(.A1(new_n5935_), .A2(\A[236] ), .ZN(new_n5936_));
  AOI21_X1   g04927(.A1(new_n5934_), .A2(new_n5936_), .B(new_n5928_), .ZN(new_n5937_));
  INV_X1     g04928(.I(new_n5929_), .ZN(new_n5938_));
  AOI21_X1   g04929(.A1(new_n5938_), .A2(new_n5930_), .B(\A[235] ), .ZN(new_n5939_));
  NOR2_X1    g04930(.A1(new_n5939_), .A2(new_n5937_), .ZN(new_n5940_));
  INV_X1     g04931(.I(\A[239] ), .ZN(new_n5941_));
  NAND2_X1   g04932(.A1(new_n5941_), .A2(\A[240] ), .ZN(new_n5942_));
  INV_X1     g04933(.I(\A[240] ), .ZN(new_n5943_));
  NAND2_X1   g04934(.A1(new_n5943_), .A2(\A[239] ), .ZN(new_n5944_));
  AOI21_X1   g04935(.A1(new_n5942_), .A2(new_n5944_), .B(new_n5924_), .ZN(new_n5945_));
  OR2_X2     g04936(.A1(\A[239] ), .A2(\A[240] ), .Z(new_n5946_));
  AOI21_X1   g04937(.A1(new_n5946_), .A2(new_n5926_), .B(\A[238] ), .ZN(new_n5947_));
  NOR2_X1    g04938(.A1(new_n5945_), .A2(new_n5947_), .ZN(new_n5948_));
  AOI21_X1   g04939(.A1(new_n5940_), .A2(new_n5948_), .B(new_n5932_), .ZN(new_n5949_));
  NOR2_X1    g04940(.A1(new_n5935_), .A2(\A[236] ), .ZN(new_n5950_));
  NOR2_X1    g04941(.A1(new_n5933_), .A2(\A[237] ), .ZN(new_n5951_));
  OAI21_X1   g04942(.A1(new_n5950_), .A2(new_n5951_), .B(\A[235] ), .ZN(new_n5952_));
  INV_X1     g04943(.I(new_n5930_), .ZN(new_n5953_));
  OAI21_X1   g04944(.A1(new_n5953_), .A2(new_n5929_), .B(new_n5928_), .ZN(new_n5954_));
  NAND2_X1   g04945(.A1(new_n5952_), .A2(new_n5954_), .ZN(new_n5955_));
  NOR2_X1    g04946(.A1(new_n5943_), .A2(\A[239] ), .ZN(new_n5956_));
  NOR2_X1    g04947(.A1(new_n5941_), .A2(\A[240] ), .ZN(new_n5957_));
  OAI21_X1   g04948(.A1(new_n5956_), .A2(new_n5957_), .B(\A[238] ), .ZN(new_n5958_));
  INV_X1     g04949(.I(new_n5926_), .ZN(new_n5959_));
  OAI21_X1   g04950(.A1(new_n5959_), .A2(new_n5925_), .B(new_n5924_), .ZN(new_n5960_));
  NAND2_X1   g04951(.A1(new_n5958_), .A2(new_n5960_), .ZN(new_n5961_));
  NOR3_X1    g04952(.A1(new_n5955_), .A2(new_n5961_), .A3(new_n5931_), .ZN(new_n5962_));
  OAI21_X1   g04953(.A1(new_n5962_), .A2(new_n5949_), .B(new_n5927_), .ZN(new_n5963_));
  INV_X1     g04954(.I(new_n5927_), .ZN(new_n5964_));
  OAI21_X1   g04955(.A1(new_n5955_), .A2(new_n5961_), .B(new_n5931_), .ZN(new_n5965_));
  NAND3_X1   g04956(.A1(new_n5940_), .A2(new_n5948_), .A3(new_n5932_), .ZN(new_n5966_));
  NAND3_X1   g04957(.A1(new_n5965_), .A2(new_n5966_), .A3(new_n5964_), .ZN(new_n5967_));
  NAND2_X1   g04958(.A1(new_n5963_), .A2(new_n5967_), .ZN(new_n5968_));
  INV_X1     g04959(.I(\A[244] ), .ZN(new_n5969_));
  NOR2_X1    g04960(.A1(\A[245] ), .A2(\A[246] ), .ZN(new_n5970_));
  NAND2_X1   g04961(.A1(\A[245] ), .A2(\A[246] ), .ZN(new_n5971_));
  AOI21_X1   g04962(.A1(new_n5969_), .A2(new_n5971_), .B(new_n5970_), .ZN(new_n5972_));
  INV_X1     g04963(.I(new_n5972_), .ZN(new_n5973_));
  INV_X1     g04964(.I(\A[241] ), .ZN(new_n5974_));
  NOR2_X1    g04965(.A1(\A[242] ), .A2(\A[243] ), .ZN(new_n5975_));
  NAND2_X1   g04966(.A1(\A[242] ), .A2(\A[243] ), .ZN(new_n5976_));
  AOI21_X1   g04967(.A1(new_n5974_), .A2(new_n5976_), .B(new_n5975_), .ZN(new_n5977_));
  INV_X1     g04968(.I(\A[246] ), .ZN(new_n5978_));
  NOR2_X1    g04969(.A1(new_n5978_), .A2(\A[245] ), .ZN(new_n5979_));
  INV_X1     g04970(.I(\A[245] ), .ZN(new_n5980_));
  NOR2_X1    g04971(.A1(new_n5980_), .A2(\A[246] ), .ZN(new_n5981_));
  OAI21_X1   g04972(.A1(new_n5979_), .A2(new_n5981_), .B(\A[244] ), .ZN(new_n5982_));
  INV_X1     g04973(.I(new_n5971_), .ZN(new_n5983_));
  OAI21_X1   g04974(.A1(new_n5983_), .A2(new_n5970_), .B(new_n5969_), .ZN(new_n5984_));
  INV_X1     g04975(.I(\A[243] ), .ZN(new_n5985_));
  NOR2_X1    g04976(.A1(new_n5985_), .A2(\A[242] ), .ZN(new_n5986_));
  INV_X1     g04977(.I(\A[242] ), .ZN(new_n5987_));
  NOR2_X1    g04978(.A1(new_n5987_), .A2(\A[243] ), .ZN(new_n5988_));
  OAI21_X1   g04979(.A1(new_n5986_), .A2(new_n5988_), .B(\A[241] ), .ZN(new_n5989_));
  AND2_X2    g04980(.A1(\A[242] ), .A2(\A[243] ), .Z(new_n5990_));
  OAI21_X1   g04981(.A1(new_n5990_), .A2(new_n5975_), .B(new_n5974_), .ZN(new_n5991_));
  NAND4_X1   g04982(.A1(new_n5982_), .A2(new_n5989_), .A3(new_n5984_), .A4(new_n5991_), .ZN(new_n5992_));
  NAND2_X1   g04983(.A1(new_n5992_), .A2(new_n5977_), .ZN(new_n5993_));
  INV_X1     g04984(.I(new_n5977_), .ZN(new_n5994_));
  NAND2_X1   g04985(.A1(new_n5980_), .A2(\A[246] ), .ZN(new_n5995_));
  NAND2_X1   g04986(.A1(new_n5978_), .A2(\A[245] ), .ZN(new_n5996_));
  AOI21_X1   g04987(.A1(new_n5995_), .A2(new_n5996_), .B(new_n5969_), .ZN(new_n5997_));
  INV_X1     g04988(.I(new_n5970_), .ZN(new_n5998_));
  AOI21_X1   g04989(.A1(new_n5998_), .A2(new_n5971_), .B(\A[244] ), .ZN(new_n5999_));
  NOR2_X1    g04990(.A1(new_n5999_), .A2(new_n5997_), .ZN(new_n6000_));
  NAND2_X1   g04991(.A1(new_n5987_), .A2(\A[243] ), .ZN(new_n6001_));
  NAND2_X1   g04992(.A1(new_n5985_), .A2(\A[242] ), .ZN(new_n6002_));
  AOI21_X1   g04993(.A1(new_n6001_), .A2(new_n6002_), .B(new_n5974_), .ZN(new_n6003_));
  INV_X1     g04994(.I(new_n5975_), .ZN(new_n6004_));
  AOI21_X1   g04995(.A1(new_n6004_), .A2(new_n5976_), .B(\A[241] ), .ZN(new_n6005_));
  NOR2_X1    g04996(.A1(new_n6005_), .A2(new_n6003_), .ZN(new_n6006_));
  NAND3_X1   g04997(.A1(new_n6000_), .A2(new_n6006_), .A3(new_n5994_), .ZN(new_n6007_));
  AOI21_X1   g04998(.A1(new_n5993_), .A2(new_n6007_), .B(new_n5973_), .ZN(new_n6008_));
  AOI21_X1   g04999(.A1(new_n6000_), .A2(new_n6006_), .B(new_n5994_), .ZN(new_n6009_));
  NOR2_X1    g05000(.A1(new_n5992_), .A2(new_n5977_), .ZN(new_n6010_));
  NOR3_X1    g05001(.A1(new_n6010_), .A2(new_n6009_), .A3(new_n5972_), .ZN(new_n6011_));
  NOR2_X1    g05002(.A1(new_n6011_), .A2(new_n6008_), .ZN(new_n6012_));
  NAND2_X1   g05003(.A1(new_n5927_), .A2(new_n5931_), .ZN(new_n6013_));
  NOR3_X1    g05004(.A1(new_n5955_), .A2(new_n5961_), .A3(new_n6013_), .ZN(new_n6014_));
  NAND2_X1   g05005(.A1(new_n5982_), .A2(new_n5984_), .ZN(new_n6015_));
  NAND2_X1   g05006(.A1(new_n5989_), .A2(new_n5991_), .ZN(new_n6016_));
  NAND2_X1   g05007(.A1(new_n6015_), .A2(new_n6016_), .ZN(new_n6017_));
  NAND3_X1   g05008(.A1(new_n6014_), .A2(new_n5992_), .A3(new_n6017_), .ZN(new_n6018_));
  NAND2_X1   g05009(.A1(new_n5940_), .A2(new_n5948_), .ZN(new_n6019_));
  NAND2_X1   g05010(.A1(new_n5955_), .A2(new_n5961_), .ZN(new_n6020_));
  NAND2_X1   g05011(.A1(new_n6020_), .A2(new_n6019_), .ZN(new_n6021_));
  NAND4_X1   g05012(.A1(new_n6000_), .A2(new_n6006_), .A3(new_n5972_), .A4(new_n5977_), .ZN(new_n6022_));
  NOR3_X1    g05013(.A1(new_n6018_), .A2(new_n6021_), .A3(new_n6022_), .ZN(new_n6023_));
  NOR2_X1    g05014(.A1(new_n6000_), .A2(new_n6006_), .ZN(new_n6024_));
  NAND2_X1   g05015(.A1(new_n5972_), .A2(new_n5977_), .ZN(new_n6025_));
  NOR2_X1    g05016(.A1(new_n6024_), .A2(new_n6025_), .ZN(new_n6026_));
  NOR3_X1    g05017(.A1(new_n6018_), .A2(new_n6021_), .A3(new_n6026_), .ZN(new_n6027_));
  AOI21_X1   g05018(.A1(new_n6012_), .A2(new_n6023_), .B(new_n5968_), .ZN(new_n6028_));
  INV_X1     g05019(.I(new_n5992_), .ZN(new_n6029_));
  NOR3_X1    g05020(.A1(new_n6022_), .A2(new_n6029_), .A3(new_n6024_), .ZN(new_n6030_));
  NAND3_X1   g05021(.A1(new_n6014_), .A2(new_n6020_), .A3(new_n6019_), .ZN(new_n6031_));
  NOR2_X1    g05022(.A1(new_n6030_), .A2(new_n6031_), .ZN(new_n6032_));
  NOR3_X1    g05023(.A1(new_n6015_), .A2(new_n6016_), .A3(new_n6025_), .ZN(new_n6033_));
  NAND3_X1   g05024(.A1(new_n6033_), .A2(new_n6017_), .A3(new_n5992_), .ZN(new_n6034_));
  NOR2_X1    g05025(.A1(new_n5955_), .A2(new_n5961_), .ZN(new_n6035_));
  NAND4_X1   g05026(.A1(new_n5940_), .A2(new_n5948_), .A3(new_n5927_), .A4(new_n5931_), .ZN(new_n6036_));
  NOR2_X1    g05027(.A1(new_n5940_), .A2(new_n5948_), .ZN(new_n6037_));
  NOR3_X1    g05028(.A1(new_n6036_), .A2(new_n6035_), .A3(new_n6037_), .ZN(new_n6038_));
  NOR2_X1    g05029(.A1(new_n6038_), .A2(new_n6034_), .ZN(new_n6039_));
  INV_X1     g05030(.I(\A[231] ), .ZN(new_n6040_));
  NOR2_X1    g05031(.A1(new_n6040_), .A2(\A[230] ), .ZN(new_n6041_));
  INV_X1     g05032(.I(\A[230] ), .ZN(new_n6042_));
  NOR2_X1    g05033(.A1(new_n6042_), .A2(\A[231] ), .ZN(new_n6043_));
  OAI21_X1   g05034(.A1(new_n6041_), .A2(new_n6043_), .B(\A[229] ), .ZN(new_n6044_));
  INV_X1     g05035(.I(\A[229] ), .ZN(new_n6045_));
  NAND2_X1   g05036(.A1(\A[230] ), .A2(\A[231] ), .ZN(new_n6046_));
  INV_X1     g05037(.I(new_n6046_), .ZN(new_n6047_));
  NOR2_X1    g05038(.A1(\A[230] ), .A2(\A[231] ), .ZN(new_n6048_));
  OAI21_X1   g05039(.A1(new_n6047_), .A2(new_n6048_), .B(new_n6045_), .ZN(new_n6049_));
  NAND2_X1   g05040(.A1(new_n6044_), .A2(new_n6049_), .ZN(new_n6050_));
  INV_X1     g05041(.I(\A[234] ), .ZN(new_n6051_));
  NOR2_X1    g05042(.A1(new_n6051_), .A2(\A[233] ), .ZN(new_n6052_));
  INV_X1     g05043(.I(\A[233] ), .ZN(new_n6053_));
  NOR2_X1    g05044(.A1(new_n6053_), .A2(\A[234] ), .ZN(new_n6054_));
  OAI21_X1   g05045(.A1(new_n6052_), .A2(new_n6054_), .B(\A[232] ), .ZN(new_n6055_));
  INV_X1     g05046(.I(\A[232] ), .ZN(new_n6056_));
  NAND2_X1   g05047(.A1(\A[233] ), .A2(\A[234] ), .ZN(new_n6057_));
  INV_X1     g05048(.I(new_n6057_), .ZN(new_n6058_));
  NOR2_X1    g05049(.A1(\A[233] ), .A2(\A[234] ), .ZN(new_n6059_));
  OAI21_X1   g05050(.A1(new_n6058_), .A2(new_n6059_), .B(new_n6056_), .ZN(new_n6060_));
  NAND2_X1   g05051(.A1(new_n6055_), .A2(new_n6060_), .ZN(new_n6061_));
  NAND2_X1   g05052(.A1(new_n6050_), .A2(new_n6061_), .ZN(new_n6062_));
  NAND2_X1   g05053(.A1(new_n6042_), .A2(\A[231] ), .ZN(new_n6063_));
  NAND2_X1   g05054(.A1(new_n6040_), .A2(\A[230] ), .ZN(new_n6064_));
  AOI21_X1   g05055(.A1(new_n6063_), .A2(new_n6064_), .B(new_n6045_), .ZN(new_n6065_));
  INV_X1     g05056(.I(new_n6048_), .ZN(new_n6066_));
  AOI21_X1   g05057(.A1(new_n6066_), .A2(new_n6046_), .B(\A[229] ), .ZN(new_n6067_));
  NOR2_X1    g05058(.A1(new_n6067_), .A2(new_n6065_), .ZN(new_n6068_));
  NAND2_X1   g05059(.A1(new_n6053_), .A2(\A[234] ), .ZN(new_n6069_));
  NAND2_X1   g05060(.A1(new_n6051_), .A2(\A[233] ), .ZN(new_n6070_));
  AOI21_X1   g05061(.A1(new_n6069_), .A2(new_n6070_), .B(new_n6056_), .ZN(new_n6071_));
  INV_X1     g05062(.I(new_n6059_), .ZN(new_n6072_));
  AOI21_X1   g05063(.A1(new_n6072_), .A2(new_n6057_), .B(\A[232] ), .ZN(new_n6073_));
  NOR2_X1    g05064(.A1(new_n6073_), .A2(new_n6071_), .ZN(new_n6074_));
  NAND2_X1   g05065(.A1(new_n6068_), .A2(new_n6074_), .ZN(new_n6075_));
  NAND2_X1   g05066(.A1(new_n6075_), .A2(new_n6062_), .ZN(new_n6076_));
  AOI21_X1   g05067(.A1(new_n6056_), .A2(new_n6057_), .B(new_n6059_), .ZN(new_n6077_));
  AOI21_X1   g05068(.A1(new_n6045_), .A2(new_n6046_), .B(new_n6048_), .ZN(new_n6078_));
  NAND2_X1   g05069(.A1(new_n6077_), .A2(new_n6078_), .ZN(new_n6079_));
  NOR3_X1    g05070(.A1(new_n6050_), .A2(new_n6061_), .A3(new_n6079_), .ZN(new_n6080_));
  INV_X1     g05071(.I(new_n6080_), .ZN(new_n6081_));
  INV_X1     g05072(.I(\A[225] ), .ZN(new_n6082_));
  NOR2_X1    g05073(.A1(new_n6082_), .A2(\A[224] ), .ZN(new_n6083_));
  INV_X1     g05074(.I(\A[224] ), .ZN(new_n6084_));
  NOR2_X1    g05075(.A1(new_n6084_), .A2(\A[225] ), .ZN(new_n6085_));
  OAI21_X1   g05076(.A1(new_n6083_), .A2(new_n6085_), .B(\A[223] ), .ZN(new_n6086_));
  INV_X1     g05077(.I(\A[223] ), .ZN(new_n6087_));
  NOR2_X1    g05078(.A1(\A[224] ), .A2(\A[225] ), .ZN(new_n6088_));
  NAND2_X1   g05079(.A1(\A[224] ), .A2(\A[225] ), .ZN(new_n6089_));
  INV_X1     g05080(.I(new_n6089_), .ZN(new_n6090_));
  OAI21_X1   g05081(.A1(new_n6090_), .A2(new_n6088_), .B(new_n6087_), .ZN(new_n6091_));
  NAND2_X1   g05082(.A1(new_n6086_), .A2(new_n6091_), .ZN(new_n6092_));
  INV_X1     g05083(.I(\A[228] ), .ZN(new_n6094_));
  NOR2_X1    g05084(.A1(new_n6094_), .A2(\A[227] ), .ZN(new_n6095_));
  INV_X1     g05085(.I(\A[227] ), .ZN(new_n6096_));
  NOR2_X1    g05086(.A1(new_n6096_), .A2(\A[228] ), .ZN(new_n6097_));
  OAI21_X1   g05087(.A1(new_n6095_), .A2(new_n6097_), .B(\A[226] ), .ZN(new_n6098_));
  INV_X1     g05088(.I(\A[226] ), .ZN(new_n6099_));
  NOR2_X1    g05089(.A1(\A[227] ), .A2(\A[228] ), .ZN(new_n6100_));
  NAND2_X1   g05090(.A1(\A[227] ), .A2(\A[228] ), .ZN(new_n6101_));
  INV_X1     g05091(.I(new_n6101_), .ZN(new_n6102_));
  OAI21_X1   g05092(.A1(new_n6102_), .A2(new_n6100_), .B(new_n6099_), .ZN(new_n6103_));
  NAND2_X1   g05093(.A1(new_n6098_), .A2(new_n6103_), .ZN(new_n6104_));
  AOI21_X1   g05094(.A1(new_n6099_), .A2(new_n6101_), .B(new_n6100_), .ZN(new_n6106_));
  AOI21_X1   g05095(.A1(new_n6087_), .A2(new_n6089_), .B(new_n6088_), .ZN(new_n6107_));
  NAND2_X1   g05096(.A1(new_n6106_), .A2(new_n6107_), .ZN(new_n6108_));
  NOR2_X1    g05097(.A1(new_n6076_), .A2(new_n6081_), .ZN(new_n6110_));
  OAI21_X1   g05098(.A1(new_n6032_), .A2(new_n6039_), .B(new_n6110_), .ZN(new_n6111_));
  NOR2_X1    g05099(.A1(new_n6028_), .A2(new_n6111_), .ZN(new_n6112_));
  AOI21_X1   g05100(.A1(new_n5965_), .A2(new_n5966_), .B(new_n5964_), .ZN(new_n6113_));
  NOR3_X1    g05101(.A1(new_n5962_), .A2(new_n5949_), .A3(new_n5927_), .ZN(new_n6114_));
  NOR2_X1    g05102(.A1(new_n6114_), .A2(new_n6113_), .ZN(new_n6115_));
  OAI21_X1   g05103(.A1(new_n6010_), .A2(new_n6009_), .B(new_n5972_), .ZN(new_n6116_));
  NAND3_X1   g05104(.A1(new_n5993_), .A2(new_n6007_), .A3(new_n5973_), .ZN(new_n6117_));
  NAND2_X1   g05105(.A1(new_n6116_), .A2(new_n6117_), .ZN(new_n6118_));
  NOR3_X1    g05106(.A1(new_n6036_), .A2(new_n6029_), .A3(new_n6024_), .ZN(new_n6119_));
  NAND4_X1   g05107(.A1(new_n6119_), .A2(new_n6019_), .A3(new_n6020_), .A4(new_n6033_), .ZN(new_n6120_));
  OAI21_X1   g05108(.A1(new_n6120_), .A2(new_n6118_), .B(new_n6115_), .ZN(new_n6121_));
  NAND2_X1   g05109(.A1(new_n6038_), .A2(new_n6034_), .ZN(new_n6122_));
  NAND2_X1   g05110(.A1(new_n6030_), .A2(new_n6031_), .ZN(new_n6123_));
  NOR2_X1    g05111(.A1(new_n6068_), .A2(new_n6074_), .ZN(new_n6124_));
  NOR4_X1    g05112(.A1(new_n6065_), .A2(new_n6067_), .A3(new_n6073_), .A4(new_n6071_), .ZN(new_n6125_));
  NOR2_X1    g05113(.A1(new_n6124_), .A2(new_n6125_), .ZN(new_n6126_));
  NAND2_X1   g05114(.A1(new_n6126_), .A2(new_n6080_), .ZN(new_n6127_));
  AOI21_X1   g05115(.A1(new_n6123_), .A2(new_n6122_), .B(new_n6127_), .ZN(new_n6128_));
  NOR2_X1    g05116(.A1(new_n6121_), .A2(new_n6128_), .ZN(new_n6129_));
  NOR2_X1    g05117(.A1(new_n6028_), .A2(new_n6111_), .ZN(new_n6130_));
  NOR2_X1    g05118(.A1(new_n6129_), .A2(new_n6130_), .ZN(new_n6131_));
  INV_X1     g05119(.I(new_n6077_), .ZN(new_n6132_));
  OAI21_X1   g05120(.A1(new_n6050_), .A2(new_n6061_), .B(new_n6078_), .ZN(new_n6133_));
  INV_X1     g05121(.I(new_n6078_), .ZN(new_n6134_));
  NAND2_X1   g05122(.A1(new_n6125_), .A2(new_n6134_), .ZN(new_n6135_));
  AOI21_X1   g05123(.A1(new_n6135_), .A2(new_n6133_), .B(new_n6132_), .ZN(new_n6136_));
  NOR2_X1    g05124(.A1(new_n6125_), .A2(new_n6134_), .ZN(new_n6137_));
  NOR3_X1    g05125(.A1(new_n6050_), .A2(new_n6061_), .A3(new_n6078_), .ZN(new_n6138_));
  NOR3_X1    g05126(.A1(new_n6137_), .A2(new_n6138_), .A3(new_n6077_), .ZN(new_n6139_));
  NOR3_X1    g05127(.A1(new_n6092_), .A2(new_n6104_), .A3(new_n6108_), .ZN(new_n6140_));
  NAND2_X1   g05128(.A1(new_n6084_), .A2(\A[225] ), .ZN(new_n6141_));
  NAND2_X1   g05129(.A1(new_n6082_), .A2(\A[224] ), .ZN(new_n6142_));
  AOI21_X1   g05130(.A1(new_n6141_), .A2(new_n6142_), .B(new_n6087_), .ZN(new_n6143_));
  INV_X1     g05131(.I(new_n6088_), .ZN(new_n6144_));
  AOI21_X1   g05132(.A1(new_n6144_), .A2(new_n6089_), .B(\A[223] ), .ZN(new_n6145_));
  NAND2_X1   g05133(.A1(new_n6096_), .A2(\A[228] ), .ZN(new_n6146_));
  NAND2_X1   g05134(.A1(new_n6094_), .A2(\A[227] ), .ZN(new_n6147_));
  AOI21_X1   g05135(.A1(new_n6146_), .A2(new_n6147_), .B(new_n6099_), .ZN(new_n6148_));
  INV_X1     g05136(.I(new_n6100_), .ZN(new_n6149_));
  AOI21_X1   g05137(.A1(new_n6149_), .A2(new_n6101_), .B(\A[226] ), .ZN(new_n6150_));
  NOR4_X1    g05138(.A1(new_n6143_), .A2(new_n6145_), .A3(new_n6150_), .A4(new_n6148_), .ZN(new_n6151_));
  AOI22_X1   g05139(.A1(new_n6086_), .A2(new_n6091_), .B1(new_n6098_), .B2(new_n6103_), .ZN(new_n6152_));
  NOR2_X1    g05140(.A1(new_n6152_), .A2(new_n6151_), .ZN(new_n6153_));
  INV_X1     g05141(.I(new_n6079_), .ZN(new_n6154_));
  NAND2_X1   g05142(.A1(new_n6132_), .A2(new_n6134_), .ZN(new_n6155_));
  AOI21_X1   g05143(.A1(new_n6125_), .A2(new_n6155_), .B(new_n6154_), .ZN(new_n6156_));
  NAND4_X1   g05144(.A1(new_n6126_), .A2(new_n6153_), .A3(new_n6156_), .A4(new_n6140_), .ZN(new_n6157_));
  NOR3_X1    g05145(.A1(new_n6157_), .A2(new_n6136_), .A3(new_n6139_), .ZN(new_n6158_));
  INV_X1     g05146(.I(new_n6107_), .ZN(new_n6159_));
  NOR2_X1    g05147(.A1(new_n6151_), .A2(new_n6159_), .ZN(new_n6160_));
  NOR3_X1    g05148(.A1(new_n6092_), .A2(new_n6104_), .A3(new_n6107_), .ZN(new_n6161_));
  OAI21_X1   g05149(.A1(new_n6160_), .A2(new_n6161_), .B(new_n6106_), .ZN(new_n6162_));
  INV_X1     g05150(.I(new_n6106_), .ZN(new_n6163_));
  OAI21_X1   g05151(.A1(new_n6092_), .A2(new_n6104_), .B(new_n6107_), .ZN(new_n6164_));
  NAND2_X1   g05152(.A1(new_n6151_), .A2(new_n6159_), .ZN(new_n6165_));
  NAND3_X1   g05153(.A1(new_n6165_), .A2(new_n6164_), .A3(new_n6163_), .ZN(new_n6166_));
  NAND2_X1   g05154(.A1(new_n6162_), .A2(new_n6166_), .ZN(new_n6167_));
  NAND2_X1   g05155(.A1(new_n6158_), .A2(new_n6167_), .ZN(new_n6168_));
  NAND4_X1   g05156(.A1(new_n6126_), .A2(new_n6080_), .A3(new_n6153_), .A4(new_n6140_), .ZN(new_n6169_));
  NAND2_X1   g05157(.A1(new_n6167_), .A2(new_n6169_), .ZN(new_n6170_));
  NOR4_X1    g05158(.A1(new_n6124_), .A2(new_n6125_), .A3(new_n6132_), .A4(new_n6134_), .ZN(new_n6171_));
  NOR3_X1    g05159(.A1(new_n6139_), .A2(new_n6136_), .A3(new_n6171_), .ZN(new_n6172_));
  NAND3_X1   g05160(.A1(new_n6080_), .A2(new_n6075_), .A3(new_n6062_), .ZN(new_n6173_));
  NAND2_X1   g05161(.A1(new_n6153_), .A2(new_n6140_), .ZN(new_n6174_));
  AOI21_X1   g05162(.A1(new_n6165_), .A2(new_n6164_), .B(new_n6163_), .ZN(new_n6175_));
  NOR3_X1    g05163(.A1(new_n6160_), .A2(new_n6161_), .A3(new_n6106_), .ZN(new_n6176_));
  NOR4_X1    g05164(.A1(new_n6175_), .A2(new_n6176_), .A3(new_n6174_), .A4(new_n6173_), .ZN(new_n6177_));
  NOR2_X1    g05165(.A1(new_n6177_), .A2(new_n6172_), .ZN(new_n6178_));
  OAI21_X1   g05166(.A1(new_n6137_), .A2(new_n6138_), .B(new_n6077_), .ZN(new_n6179_));
  NAND3_X1   g05167(.A1(new_n6135_), .A2(new_n6133_), .A3(new_n6132_), .ZN(new_n6180_));
  NAND4_X1   g05168(.A1(new_n6075_), .A2(new_n6062_), .A3(new_n6077_), .A4(new_n6078_), .ZN(new_n6181_));
  NAND3_X1   g05169(.A1(new_n6179_), .A2(new_n6180_), .A3(new_n6181_), .ZN(new_n6182_));
  NOR3_X1    g05170(.A1(new_n6182_), .A2(new_n6167_), .A3(new_n6169_), .ZN(new_n6183_));
  OAI21_X1   g05171(.A1(new_n6178_), .A2(new_n6183_), .B(new_n6170_), .ZN(new_n6184_));
  NAND2_X1   g05172(.A1(new_n6184_), .A2(new_n6168_), .ZN(new_n6185_));
  NOR2_X1    g05173(.A1(new_n6185_), .A2(new_n6131_), .ZN(new_n6186_));
  NAND2_X1   g05174(.A1(new_n6012_), .A2(new_n6027_), .ZN(new_n6187_));
  OAI21_X1   g05175(.A1(new_n6120_), .A2(new_n6118_), .B(new_n5968_), .ZN(new_n6188_));
  NOR2_X1    g05176(.A1(new_n5972_), .A2(new_n5977_), .ZN(new_n6189_));
  OAI21_X1   g05177(.A1(new_n5992_), .A2(new_n6189_), .B(new_n6025_), .ZN(new_n6190_));
  NOR2_X1    g05178(.A1(new_n5927_), .A2(new_n5931_), .ZN(new_n6191_));
  OAI21_X1   g05179(.A1(new_n6019_), .A2(new_n6191_), .B(new_n6013_), .ZN(new_n6192_));
  XNOR2_X1   g05180(.A1(new_n6192_), .A2(new_n6190_), .ZN(new_n6193_));
  NAND3_X1   g05181(.A1(new_n6188_), .A2(new_n6193_), .A3(new_n6187_), .ZN(new_n6194_));
  INV_X1     g05182(.I(new_n6173_), .ZN(new_n6195_));
  NAND4_X1   g05183(.A1(new_n6182_), .A2(new_n6195_), .A3(new_n6140_), .A4(new_n6153_), .ZN(new_n6196_));
  AOI21_X1   g05184(.A1(new_n6196_), .A2(new_n6167_), .B(new_n6158_), .ZN(new_n6197_));
  INV_X1     g05185(.I(new_n6156_), .ZN(new_n6198_));
  NAND3_X1   g05186(.A1(new_n6179_), .A2(new_n6180_), .A3(new_n6126_), .ZN(new_n6199_));
  INV_X1     g05187(.I(new_n6151_), .ZN(new_n6200_));
  NOR2_X1    g05188(.A1(new_n6106_), .A2(new_n6107_), .ZN(new_n6201_));
  OAI21_X1   g05189(.A1(new_n6200_), .A2(new_n6201_), .B(new_n6108_), .ZN(new_n6202_));
  AOI21_X1   g05190(.A1(new_n6199_), .A2(new_n6198_), .B(new_n6202_), .ZN(new_n6203_));
  NOR3_X1    g05191(.A1(new_n6139_), .A2(new_n6136_), .A3(new_n6076_), .ZN(new_n6204_));
  INV_X1     g05192(.I(new_n6202_), .ZN(new_n6205_));
  NOR3_X1    g05193(.A1(new_n6204_), .A2(new_n6156_), .A3(new_n6205_), .ZN(new_n6206_));
  NOR2_X1    g05194(.A1(new_n6206_), .A2(new_n6203_), .ZN(new_n6207_));
  AOI21_X1   g05195(.A1(new_n6197_), .A2(new_n6207_), .B(new_n6194_), .ZN(new_n6208_));
  INV_X1     g05196(.I(new_n6194_), .ZN(new_n6209_));
  OR3_X2     g05197(.A1(new_n6157_), .A2(new_n6136_), .A3(new_n6139_), .Z(new_n6210_));
  OAI21_X1   g05198(.A1(new_n6172_), .A2(new_n6169_), .B(new_n6167_), .ZN(new_n6211_));
  OAI21_X1   g05199(.A1(new_n6204_), .A2(new_n6156_), .B(new_n6205_), .ZN(new_n6212_));
  NAND3_X1   g05200(.A1(new_n6199_), .A2(new_n6198_), .A3(new_n6202_), .ZN(new_n6213_));
  NAND4_X1   g05201(.A1(new_n6210_), .A2(new_n6211_), .A3(new_n6212_), .A4(new_n6213_), .ZN(new_n6214_));
  NOR2_X1    g05202(.A1(new_n6209_), .A2(new_n6214_), .ZN(new_n6215_));
  OAI22_X1   g05203(.A1(new_n6186_), .A2(new_n6112_), .B1(new_n6208_), .B2(new_n6215_), .ZN(new_n6216_));
  NAND2_X1   g05204(.A1(new_n6028_), .A2(new_n6111_), .ZN(new_n6217_));
  NAND2_X1   g05205(.A1(new_n6121_), .A2(new_n6128_), .ZN(new_n6218_));
  NAND2_X1   g05206(.A1(new_n6218_), .A2(new_n6217_), .ZN(new_n6219_));
  INV_X1     g05207(.I(new_n6168_), .ZN(new_n6220_));
  OAI21_X1   g05208(.A1(new_n6167_), .A2(new_n6169_), .B(new_n6182_), .ZN(new_n6221_));
  NAND2_X1   g05209(.A1(new_n6177_), .A2(new_n6172_), .ZN(new_n6222_));
  NAND2_X1   g05210(.A1(new_n6221_), .A2(new_n6222_), .ZN(new_n6223_));
  AOI21_X1   g05211(.A1(new_n6223_), .A2(new_n6170_), .B(new_n6220_), .ZN(new_n6224_));
  OAI21_X1   g05212(.A1(new_n6224_), .A2(new_n6121_), .B(new_n6219_), .ZN(new_n6225_));
  NAND2_X1   g05213(.A1(new_n6214_), .A2(new_n6194_), .ZN(new_n6226_));
  NAND3_X1   g05214(.A1(new_n6209_), .A2(new_n6207_), .A3(new_n6197_), .ZN(new_n6227_));
  NAND2_X1   g05215(.A1(new_n6227_), .A2(new_n6226_), .ZN(new_n6228_));
  NAND2_X1   g05216(.A1(new_n6228_), .A2(new_n6225_), .ZN(new_n6229_));
  NAND2_X1   g05217(.A1(new_n6229_), .A2(new_n6216_), .ZN(new_n6230_));
  INV_X1     g05218(.I(\A[268] ), .ZN(new_n6231_));
  NOR2_X1    g05219(.A1(\A[269] ), .A2(\A[270] ), .ZN(new_n6232_));
  NAND2_X1   g05220(.A1(\A[269] ), .A2(\A[270] ), .ZN(new_n6233_));
  AOI21_X1   g05221(.A1(new_n6231_), .A2(new_n6233_), .B(new_n6232_), .ZN(new_n6234_));
  INV_X1     g05222(.I(new_n6234_), .ZN(new_n6235_));
  INV_X1     g05223(.I(\A[265] ), .ZN(new_n6236_));
  NOR2_X1    g05224(.A1(\A[266] ), .A2(\A[267] ), .ZN(new_n6237_));
  NAND2_X1   g05225(.A1(\A[266] ), .A2(\A[267] ), .ZN(new_n6238_));
  AOI21_X1   g05226(.A1(new_n6236_), .A2(new_n6238_), .B(new_n6237_), .ZN(new_n6239_));
  INV_X1     g05227(.I(\A[267] ), .ZN(new_n6240_));
  NOR2_X1    g05228(.A1(new_n6240_), .A2(\A[266] ), .ZN(new_n6241_));
  INV_X1     g05229(.I(\A[266] ), .ZN(new_n6242_));
  NOR2_X1    g05230(.A1(new_n6242_), .A2(\A[267] ), .ZN(new_n6243_));
  OAI21_X1   g05231(.A1(new_n6241_), .A2(new_n6243_), .B(\A[265] ), .ZN(new_n6244_));
  INV_X1     g05232(.I(new_n6238_), .ZN(new_n6245_));
  OAI21_X1   g05233(.A1(new_n6245_), .A2(new_n6237_), .B(new_n6236_), .ZN(new_n6246_));
  NAND2_X1   g05234(.A1(new_n6244_), .A2(new_n6246_), .ZN(new_n6247_));
  INV_X1     g05235(.I(\A[270] ), .ZN(new_n6248_));
  NOR2_X1    g05236(.A1(new_n6248_), .A2(\A[269] ), .ZN(new_n6249_));
  INV_X1     g05237(.I(\A[269] ), .ZN(new_n6250_));
  NOR2_X1    g05238(.A1(new_n6250_), .A2(\A[270] ), .ZN(new_n6251_));
  OAI21_X1   g05239(.A1(new_n6249_), .A2(new_n6251_), .B(\A[268] ), .ZN(new_n6252_));
  INV_X1     g05240(.I(new_n6233_), .ZN(new_n6253_));
  OAI21_X1   g05241(.A1(new_n6253_), .A2(new_n6232_), .B(new_n6231_), .ZN(new_n6254_));
  NAND2_X1   g05242(.A1(new_n6252_), .A2(new_n6254_), .ZN(new_n6255_));
  OAI21_X1   g05243(.A1(new_n6247_), .A2(new_n6255_), .B(new_n6239_), .ZN(new_n6256_));
  INV_X1     g05244(.I(new_n6239_), .ZN(new_n6257_));
  NAND2_X1   g05245(.A1(new_n6242_), .A2(\A[267] ), .ZN(new_n6258_));
  NAND2_X1   g05246(.A1(new_n6240_), .A2(\A[266] ), .ZN(new_n6259_));
  AOI21_X1   g05247(.A1(new_n6258_), .A2(new_n6259_), .B(new_n6236_), .ZN(new_n6260_));
  INV_X1     g05248(.I(new_n6237_), .ZN(new_n6261_));
  AOI21_X1   g05249(.A1(new_n6261_), .A2(new_n6238_), .B(\A[265] ), .ZN(new_n6262_));
  NOR2_X1    g05250(.A1(new_n6262_), .A2(new_n6260_), .ZN(new_n6263_));
  NAND2_X1   g05251(.A1(new_n6250_), .A2(\A[270] ), .ZN(new_n6264_));
  NAND2_X1   g05252(.A1(new_n6248_), .A2(\A[269] ), .ZN(new_n6265_));
  AOI21_X1   g05253(.A1(new_n6264_), .A2(new_n6265_), .B(new_n6231_), .ZN(new_n6266_));
  INV_X1     g05254(.I(new_n6232_), .ZN(new_n6267_));
  AOI21_X1   g05255(.A1(new_n6267_), .A2(new_n6233_), .B(\A[268] ), .ZN(new_n6268_));
  NOR2_X1    g05256(.A1(new_n6268_), .A2(new_n6266_), .ZN(new_n6269_));
  NAND3_X1   g05257(.A1(new_n6263_), .A2(new_n6269_), .A3(new_n6257_), .ZN(new_n6270_));
  AOI21_X1   g05258(.A1(new_n6256_), .A2(new_n6270_), .B(new_n6235_), .ZN(new_n6271_));
  NOR4_X1    g05259(.A1(new_n6260_), .A2(new_n6262_), .A3(new_n6268_), .A4(new_n6266_), .ZN(new_n6272_));
  NOR2_X1    g05260(.A1(new_n6272_), .A2(new_n6257_), .ZN(new_n6273_));
  NOR3_X1    g05261(.A1(new_n6247_), .A2(new_n6255_), .A3(new_n6239_), .ZN(new_n6274_));
  NOR3_X1    g05262(.A1(new_n6273_), .A2(new_n6274_), .A3(new_n6234_), .ZN(new_n6275_));
  INV_X1     g05263(.I(\A[261] ), .ZN(new_n6276_));
  NOR2_X1    g05264(.A1(new_n6276_), .A2(\A[260] ), .ZN(new_n6277_));
  INV_X1     g05265(.I(\A[260] ), .ZN(new_n6278_));
  NOR2_X1    g05266(.A1(new_n6278_), .A2(\A[261] ), .ZN(new_n6279_));
  OAI21_X1   g05267(.A1(new_n6277_), .A2(new_n6279_), .B(\A[259] ), .ZN(new_n6280_));
  INV_X1     g05268(.I(\A[259] ), .ZN(new_n6281_));
  NOR2_X1    g05269(.A1(\A[260] ), .A2(\A[261] ), .ZN(new_n6282_));
  NAND2_X1   g05270(.A1(\A[260] ), .A2(\A[261] ), .ZN(new_n6283_));
  INV_X1     g05271(.I(new_n6283_), .ZN(new_n6284_));
  OAI21_X1   g05272(.A1(new_n6284_), .A2(new_n6282_), .B(new_n6281_), .ZN(new_n6285_));
  NAND2_X1   g05273(.A1(new_n6280_), .A2(new_n6285_), .ZN(new_n6286_));
  INV_X1     g05274(.I(\A[262] ), .ZN(new_n6287_));
  INV_X1     g05275(.I(\A[263] ), .ZN(new_n6288_));
  NAND2_X1   g05276(.A1(new_n6288_), .A2(\A[264] ), .ZN(new_n6289_));
  INV_X1     g05277(.I(\A[264] ), .ZN(new_n6290_));
  NAND2_X1   g05278(.A1(new_n6290_), .A2(\A[263] ), .ZN(new_n6291_));
  AOI21_X1   g05279(.A1(new_n6289_), .A2(new_n6291_), .B(new_n6287_), .ZN(new_n6292_));
  NOR2_X1    g05280(.A1(\A[263] ), .A2(\A[264] ), .ZN(new_n6293_));
  INV_X1     g05281(.I(new_n6293_), .ZN(new_n6294_));
  NAND2_X1   g05282(.A1(\A[263] ), .A2(\A[264] ), .ZN(new_n6295_));
  AOI21_X1   g05283(.A1(new_n6294_), .A2(new_n6295_), .B(\A[262] ), .ZN(new_n6296_));
  NOR2_X1    g05284(.A1(new_n6296_), .A2(new_n6292_), .ZN(new_n6297_));
  NOR2_X1    g05285(.A1(new_n6297_), .A2(new_n6286_), .ZN(new_n6298_));
  NAND2_X1   g05286(.A1(new_n6278_), .A2(\A[261] ), .ZN(new_n6299_));
  NAND2_X1   g05287(.A1(new_n6276_), .A2(\A[260] ), .ZN(new_n6300_));
  AOI21_X1   g05288(.A1(new_n6299_), .A2(new_n6300_), .B(new_n6281_), .ZN(new_n6301_));
  INV_X1     g05289(.I(new_n6282_), .ZN(new_n6302_));
  AOI21_X1   g05290(.A1(new_n6302_), .A2(new_n6283_), .B(\A[259] ), .ZN(new_n6303_));
  NOR2_X1    g05291(.A1(new_n6303_), .A2(new_n6301_), .ZN(new_n6304_));
  NOR2_X1    g05292(.A1(new_n6290_), .A2(\A[263] ), .ZN(new_n6305_));
  NOR2_X1    g05293(.A1(new_n6288_), .A2(\A[264] ), .ZN(new_n6306_));
  OAI21_X1   g05294(.A1(new_n6305_), .A2(new_n6306_), .B(\A[262] ), .ZN(new_n6307_));
  INV_X1     g05295(.I(new_n6295_), .ZN(new_n6308_));
  OAI21_X1   g05296(.A1(new_n6308_), .A2(new_n6293_), .B(new_n6287_), .ZN(new_n6309_));
  NAND2_X1   g05297(.A1(new_n6307_), .A2(new_n6309_), .ZN(new_n6310_));
  NOR2_X1    g05298(.A1(new_n6304_), .A2(new_n6310_), .ZN(new_n6311_));
  NOR2_X1    g05299(.A1(new_n6269_), .A2(new_n6247_), .ZN(new_n6312_));
  NOR2_X1    g05300(.A1(new_n6263_), .A2(new_n6255_), .ZN(new_n6313_));
  OAI22_X1   g05301(.A1(new_n6298_), .A2(new_n6311_), .B1(new_n6312_), .B2(new_n6313_), .ZN(new_n6314_));
  NAND4_X1   g05302(.A1(new_n6280_), .A2(new_n6285_), .A3(new_n6307_), .A4(new_n6309_), .ZN(new_n6315_));
  AOI21_X1   g05303(.A1(new_n6287_), .A2(new_n6295_), .B(new_n6293_), .ZN(new_n6316_));
  AOI21_X1   g05304(.A1(new_n6281_), .A2(new_n6283_), .B(new_n6282_), .ZN(new_n6317_));
  NAND2_X1   g05305(.A1(new_n6316_), .A2(new_n6317_), .ZN(new_n6318_));
  NOR2_X1    g05306(.A1(new_n6315_), .A2(new_n6318_), .ZN(new_n6319_));
  NAND2_X1   g05307(.A1(new_n6234_), .A2(new_n6239_), .ZN(new_n6320_));
  AOI21_X1   g05308(.A1(new_n6247_), .A2(new_n6255_), .B(new_n6320_), .ZN(new_n6321_));
  INV_X1     g05309(.I(new_n6321_), .ZN(new_n6322_));
  NAND2_X1   g05310(.A1(new_n6322_), .A2(new_n6319_), .ZN(new_n6323_));
  NOR4_X1    g05311(.A1(new_n6323_), .A2(new_n6314_), .A3(new_n6275_), .A4(new_n6271_), .ZN(new_n6324_));
  NOR4_X1    g05312(.A1(new_n6301_), .A2(new_n6303_), .A3(new_n6296_), .A4(new_n6292_), .ZN(new_n6325_));
  INV_X1     g05313(.I(new_n6317_), .ZN(new_n6326_));
  NOR2_X1    g05314(.A1(new_n6325_), .A2(new_n6326_), .ZN(new_n6327_));
  NOR2_X1    g05315(.A1(new_n6315_), .A2(new_n6317_), .ZN(new_n6328_));
  OAI21_X1   g05316(.A1(new_n6327_), .A2(new_n6328_), .B(new_n6316_), .ZN(new_n6329_));
  INV_X1     g05317(.I(new_n6316_), .ZN(new_n6330_));
  NAND2_X1   g05318(.A1(new_n6315_), .A2(new_n6317_), .ZN(new_n6331_));
  NAND3_X1   g05319(.A1(new_n6304_), .A2(new_n6297_), .A3(new_n6326_), .ZN(new_n6332_));
  NAND3_X1   g05320(.A1(new_n6331_), .A2(new_n6332_), .A3(new_n6330_), .ZN(new_n6333_));
  NAND2_X1   g05321(.A1(new_n6329_), .A2(new_n6333_), .ZN(new_n6334_));
  OAI21_X1   g05322(.A1(new_n6273_), .A2(new_n6274_), .B(new_n6234_), .ZN(new_n6335_));
  NAND3_X1   g05323(.A1(new_n6256_), .A2(new_n6270_), .A3(new_n6235_), .ZN(new_n6336_));
  NAND2_X1   g05324(.A1(new_n6335_), .A2(new_n6336_), .ZN(new_n6337_));
  NOR2_X1    g05325(.A1(new_n6298_), .A2(new_n6311_), .ZN(new_n6338_));
  NOR2_X1    g05326(.A1(new_n6312_), .A2(new_n6313_), .ZN(new_n6339_));
  INV_X1     g05327(.I(new_n6318_), .ZN(new_n6340_));
  INV_X1     g05328(.I(new_n6320_), .ZN(new_n6341_));
  NAND4_X1   g05329(.A1(new_n6272_), .A2(new_n6325_), .A3(new_n6340_), .A4(new_n6341_), .ZN(new_n6342_));
  NOR3_X1    g05330(.A1(new_n6338_), .A2(new_n6339_), .A3(new_n6342_), .ZN(new_n6343_));
  NOR2_X1    g05331(.A1(new_n6337_), .A2(new_n6343_), .ZN(new_n6344_));
  NOR3_X1    g05332(.A1(new_n6344_), .A2(new_n6324_), .A3(new_n6334_), .ZN(new_n6345_));
  OAI22_X1   g05333(.A1(new_n6314_), .A2(new_n6342_), .B1(new_n6275_), .B2(new_n6271_), .ZN(new_n6346_));
  NAND2_X1   g05334(.A1(new_n6304_), .A2(new_n6310_), .ZN(new_n6347_));
  NAND2_X1   g05335(.A1(new_n6297_), .A2(new_n6286_), .ZN(new_n6348_));
  NAND2_X1   g05336(.A1(new_n6263_), .A2(new_n6255_), .ZN(new_n6349_));
  NAND2_X1   g05337(.A1(new_n6269_), .A2(new_n6247_), .ZN(new_n6350_));
  AOI22_X1   g05338(.A1(new_n6347_), .A2(new_n6348_), .B1(new_n6349_), .B2(new_n6350_), .ZN(new_n6351_));
  INV_X1     g05339(.I(new_n6342_), .ZN(new_n6352_));
  NAND4_X1   g05340(.A1(new_n6351_), .A2(new_n6352_), .A3(new_n6335_), .A4(new_n6336_), .ZN(new_n6353_));
  AOI21_X1   g05341(.A1(new_n6346_), .A2(new_n6353_), .B(new_n6334_), .ZN(new_n6354_));
  NOR2_X1    g05342(.A1(new_n6345_), .A2(new_n6354_), .ZN(new_n6355_));
  NAND2_X1   g05343(.A1(new_n6325_), .A2(new_n6340_), .ZN(new_n6356_));
  NOR2_X1    g05344(.A1(new_n6356_), .A2(new_n6321_), .ZN(new_n6357_));
  NAND4_X1   g05345(.A1(new_n6351_), .A2(new_n6335_), .A3(new_n6336_), .A4(new_n6357_), .ZN(new_n6358_));
  AOI21_X1   g05346(.A1(new_n6331_), .A2(new_n6332_), .B(new_n6330_), .ZN(new_n6359_));
  NOR3_X1    g05347(.A1(new_n6327_), .A2(new_n6328_), .A3(new_n6316_), .ZN(new_n6360_));
  NOR2_X1    g05348(.A1(new_n6360_), .A2(new_n6359_), .ZN(new_n6361_));
  NOR2_X1    g05349(.A1(new_n6275_), .A2(new_n6271_), .ZN(new_n6362_));
  NAND2_X1   g05350(.A1(new_n6347_), .A2(new_n6348_), .ZN(new_n6363_));
  NAND2_X1   g05351(.A1(new_n6349_), .A2(new_n6350_), .ZN(new_n6364_));
  NOR3_X1    g05352(.A1(new_n6247_), .A2(new_n6255_), .A3(new_n6320_), .ZN(new_n6365_));
  NAND4_X1   g05353(.A1(new_n6363_), .A2(new_n6364_), .A3(new_n6319_), .A4(new_n6365_), .ZN(new_n6366_));
  NAND2_X1   g05354(.A1(new_n6362_), .A2(new_n6366_), .ZN(new_n6367_));
  NAND3_X1   g05355(.A1(new_n6367_), .A2(new_n6358_), .A3(new_n6361_), .ZN(new_n6368_));
  AOI22_X1   g05356(.A1(new_n6351_), .A2(new_n6352_), .B1(new_n6335_), .B2(new_n6336_), .ZN(new_n6369_));
  NOR4_X1    g05357(.A1(new_n6314_), .A2(new_n6275_), .A3(new_n6271_), .A4(new_n6342_), .ZN(new_n6370_));
  OAI21_X1   g05358(.A1(new_n6369_), .A2(new_n6370_), .B(new_n6361_), .ZN(new_n6371_));
  NAND2_X1   g05359(.A1(new_n6364_), .A2(new_n6365_), .ZN(new_n6372_));
  NOR2_X1    g05360(.A1(new_n6338_), .A2(new_n6356_), .ZN(new_n6373_));
  NAND2_X1   g05361(.A1(new_n6373_), .A2(new_n6372_), .ZN(new_n6374_));
  NAND2_X1   g05362(.A1(new_n6272_), .A2(new_n6341_), .ZN(new_n6375_));
  NOR2_X1    g05363(.A1(new_n6339_), .A2(new_n6375_), .ZN(new_n6376_));
  NAND2_X1   g05364(.A1(new_n6363_), .A2(new_n6319_), .ZN(new_n6377_));
  NAND2_X1   g05365(.A1(new_n6376_), .A2(new_n6377_), .ZN(new_n6378_));
  INV_X1     g05366(.I(\A[258] ), .ZN(new_n6379_));
  NOR2_X1    g05367(.A1(new_n6379_), .A2(\A[257] ), .ZN(new_n6380_));
  INV_X1     g05368(.I(\A[257] ), .ZN(new_n6381_));
  NOR2_X1    g05369(.A1(new_n6381_), .A2(\A[258] ), .ZN(new_n6382_));
  OAI21_X1   g05370(.A1(new_n6380_), .A2(new_n6382_), .B(\A[256] ), .ZN(new_n6383_));
  INV_X1     g05371(.I(\A[256] ), .ZN(new_n6384_));
  NOR2_X1    g05372(.A1(\A[257] ), .A2(\A[258] ), .ZN(new_n6385_));
  NAND2_X1   g05373(.A1(\A[257] ), .A2(\A[258] ), .ZN(new_n6386_));
  INV_X1     g05374(.I(new_n6386_), .ZN(new_n6387_));
  OAI21_X1   g05375(.A1(new_n6387_), .A2(new_n6385_), .B(new_n6384_), .ZN(new_n6388_));
  NAND2_X1   g05376(.A1(new_n6383_), .A2(new_n6388_), .ZN(new_n6389_));
  AOI21_X1   g05377(.A1(new_n6384_), .A2(new_n6386_), .B(new_n6385_), .ZN(new_n6390_));
  NAND4_X1   g05378(.A1(new_n6390_), .A2(\A[253] ), .A3(\A[254] ), .A4(\A[255] ), .ZN(new_n6391_));
  NOR2_X1    g05379(.A1(new_n6389_), .A2(new_n6391_), .ZN(new_n6392_));
  INV_X1     g05380(.I(\A[255] ), .ZN(new_n6393_));
  NOR2_X1    g05381(.A1(new_n6393_), .A2(\A[254] ), .ZN(new_n6394_));
  INV_X1     g05382(.I(\A[254] ), .ZN(new_n6395_));
  NOR2_X1    g05383(.A1(new_n6395_), .A2(\A[255] ), .ZN(new_n6396_));
  OAI21_X1   g05384(.A1(new_n6394_), .A2(new_n6396_), .B(\A[253] ), .ZN(new_n6397_));
  INV_X1     g05385(.I(\A[253] ), .ZN(new_n6398_));
  NOR2_X1    g05386(.A1(\A[254] ), .A2(\A[255] ), .ZN(new_n6399_));
  NAND2_X1   g05387(.A1(\A[254] ), .A2(\A[255] ), .ZN(new_n6400_));
  INV_X1     g05388(.I(new_n6400_), .ZN(new_n6401_));
  OAI21_X1   g05389(.A1(new_n6401_), .A2(new_n6399_), .B(new_n6398_), .ZN(new_n6402_));
  NAND2_X1   g05390(.A1(new_n6397_), .A2(new_n6402_), .ZN(new_n6403_));
  XOR2_X1    g05391(.A1(new_n6389_), .A2(new_n6403_), .Z(new_n6404_));
  INV_X1     g05392(.I(\A[247] ), .ZN(new_n6405_));
  INV_X1     g05393(.I(\A[248] ), .ZN(new_n6406_));
  NAND2_X1   g05394(.A1(new_n6406_), .A2(\A[249] ), .ZN(new_n6407_));
  INV_X1     g05395(.I(\A[249] ), .ZN(new_n6408_));
  NAND2_X1   g05396(.A1(new_n6408_), .A2(\A[248] ), .ZN(new_n6409_));
  AOI21_X1   g05397(.A1(new_n6407_), .A2(new_n6409_), .B(new_n6405_), .ZN(new_n6410_));
  NOR2_X1    g05398(.A1(\A[248] ), .A2(\A[249] ), .ZN(new_n6411_));
  INV_X1     g05399(.I(new_n6411_), .ZN(new_n6412_));
  NAND2_X1   g05400(.A1(\A[248] ), .A2(\A[249] ), .ZN(new_n6413_));
  AOI21_X1   g05401(.A1(new_n6412_), .A2(new_n6413_), .B(\A[247] ), .ZN(new_n6414_));
  NOR2_X1    g05402(.A1(new_n6414_), .A2(new_n6410_), .ZN(new_n6415_));
  INV_X1     g05403(.I(\A[250] ), .ZN(new_n6416_));
  INV_X1     g05404(.I(\A[251] ), .ZN(new_n6417_));
  NAND2_X1   g05405(.A1(new_n6417_), .A2(\A[252] ), .ZN(new_n6418_));
  INV_X1     g05406(.I(\A[252] ), .ZN(new_n6419_));
  NAND2_X1   g05407(.A1(new_n6419_), .A2(\A[251] ), .ZN(new_n6420_));
  AOI21_X1   g05408(.A1(new_n6418_), .A2(new_n6420_), .B(new_n6416_), .ZN(new_n6421_));
  NOR2_X1    g05409(.A1(\A[251] ), .A2(\A[252] ), .ZN(new_n6422_));
  INV_X1     g05410(.I(new_n6422_), .ZN(new_n6423_));
  NAND2_X1   g05411(.A1(\A[251] ), .A2(\A[252] ), .ZN(new_n6424_));
  AOI21_X1   g05412(.A1(new_n6423_), .A2(new_n6424_), .B(\A[250] ), .ZN(new_n6425_));
  NOR2_X1    g05413(.A1(new_n6425_), .A2(new_n6421_), .ZN(new_n6426_));
  AOI21_X1   g05414(.A1(new_n6416_), .A2(new_n6424_), .B(new_n6422_), .ZN(new_n6427_));
  AOI21_X1   g05415(.A1(new_n6405_), .A2(new_n6413_), .B(new_n6411_), .ZN(new_n6428_));
  NAND2_X1   g05416(.A1(new_n6427_), .A2(new_n6428_), .ZN(new_n6429_));
  INV_X1     g05417(.I(new_n6429_), .ZN(new_n6430_));
  NAND2_X1   g05418(.A1(new_n6404_), .A2(new_n6392_), .ZN(new_n6431_));
  AOI21_X1   g05419(.A1(new_n6374_), .A2(new_n6378_), .B(new_n6431_), .ZN(new_n6432_));
  AOI21_X1   g05420(.A1(new_n6368_), .A2(new_n6371_), .B(new_n6432_), .ZN(new_n6433_));
  NOR2_X1    g05421(.A1(new_n6376_), .A2(new_n6377_), .ZN(new_n6434_));
  NOR2_X1    g05422(.A1(new_n6373_), .A2(new_n6372_), .ZN(new_n6435_));
  INV_X1     g05423(.I(new_n6431_), .ZN(new_n6436_));
  OAI21_X1   g05424(.A1(new_n6435_), .A2(new_n6434_), .B(new_n6436_), .ZN(new_n6437_));
  NOR3_X1    g05425(.A1(new_n6345_), .A2(new_n6437_), .A3(new_n6354_), .ZN(new_n6438_));
  NOR4_X1    g05426(.A1(new_n6410_), .A2(new_n6414_), .A3(new_n6425_), .A4(new_n6421_), .ZN(new_n6439_));
  INV_X1     g05427(.I(new_n6428_), .ZN(new_n6440_));
  NOR2_X1    g05428(.A1(new_n6439_), .A2(new_n6440_), .ZN(new_n6441_));
  NOR2_X1    g05429(.A1(new_n6408_), .A2(\A[248] ), .ZN(new_n6442_));
  NOR2_X1    g05430(.A1(new_n6406_), .A2(\A[249] ), .ZN(new_n6443_));
  OAI21_X1   g05431(.A1(new_n6442_), .A2(new_n6443_), .B(\A[247] ), .ZN(new_n6444_));
  INV_X1     g05432(.I(new_n6413_), .ZN(new_n6445_));
  OAI21_X1   g05433(.A1(new_n6445_), .A2(new_n6411_), .B(new_n6405_), .ZN(new_n6446_));
  NAND2_X1   g05434(.A1(new_n6444_), .A2(new_n6446_), .ZN(new_n6447_));
  NOR2_X1    g05435(.A1(new_n6419_), .A2(\A[251] ), .ZN(new_n6448_));
  NOR2_X1    g05436(.A1(new_n6417_), .A2(\A[252] ), .ZN(new_n6449_));
  OAI21_X1   g05437(.A1(new_n6448_), .A2(new_n6449_), .B(\A[250] ), .ZN(new_n6450_));
  INV_X1     g05438(.I(new_n6424_), .ZN(new_n6451_));
  OAI21_X1   g05439(.A1(new_n6451_), .A2(new_n6422_), .B(new_n6416_), .ZN(new_n6452_));
  NAND2_X1   g05440(.A1(new_n6450_), .A2(new_n6452_), .ZN(new_n6453_));
  NOR3_X1    g05441(.A1(new_n6447_), .A2(new_n6453_), .A3(new_n6428_), .ZN(new_n6454_));
  OAI21_X1   g05442(.A1(new_n6441_), .A2(new_n6454_), .B(new_n6427_), .ZN(new_n6455_));
  INV_X1     g05443(.I(new_n6427_), .ZN(new_n6456_));
  NAND4_X1   g05444(.A1(new_n6444_), .A2(new_n6446_), .A3(new_n6450_), .A4(new_n6452_), .ZN(new_n6457_));
  NAND2_X1   g05445(.A1(new_n6457_), .A2(new_n6428_), .ZN(new_n6458_));
  NAND3_X1   g05446(.A1(new_n6415_), .A2(new_n6426_), .A3(new_n6440_), .ZN(new_n6459_));
  NAND3_X1   g05447(.A1(new_n6458_), .A2(new_n6459_), .A3(new_n6456_), .ZN(new_n6460_));
  NAND2_X1   g05448(.A1(new_n6455_), .A2(new_n6460_), .ZN(new_n6461_));
  NAND2_X1   g05449(.A1(new_n6439_), .A2(new_n6430_), .ZN(new_n6462_));
  NAND2_X1   g05450(.A1(new_n6381_), .A2(\A[258] ), .ZN(new_n6463_));
  NAND2_X1   g05451(.A1(new_n6379_), .A2(\A[257] ), .ZN(new_n6464_));
  AOI21_X1   g05452(.A1(new_n6463_), .A2(new_n6464_), .B(new_n6384_), .ZN(new_n6465_));
  INV_X1     g05453(.I(new_n6385_), .ZN(new_n6466_));
  AOI21_X1   g05454(.A1(new_n6466_), .A2(new_n6386_), .B(\A[256] ), .ZN(new_n6467_));
  NOR2_X1    g05455(.A1(new_n6467_), .A2(new_n6465_), .ZN(new_n6468_));
  NAND2_X1   g05456(.A1(new_n6395_), .A2(\A[255] ), .ZN(new_n6469_));
  NAND2_X1   g05457(.A1(new_n6393_), .A2(\A[254] ), .ZN(new_n6470_));
  AOI21_X1   g05458(.A1(new_n6469_), .A2(new_n6470_), .B(new_n6398_), .ZN(new_n6471_));
  INV_X1     g05459(.I(new_n6399_), .ZN(new_n6472_));
  AOI21_X1   g05460(.A1(new_n6472_), .A2(new_n6400_), .B(\A[253] ), .ZN(new_n6473_));
  NOR2_X1    g05461(.A1(new_n6473_), .A2(new_n6471_), .ZN(new_n6474_));
  AOI21_X1   g05462(.A1(new_n6398_), .A2(new_n6400_), .B(new_n6399_), .ZN(new_n6475_));
  INV_X1     g05463(.I(new_n6475_), .ZN(new_n6476_));
  AOI21_X1   g05464(.A1(new_n6468_), .A2(new_n6474_), .B(new_n6476_), .ZN(new_n6477_));
  NOR3_X1    g05465(.A1(new_n6389_), .A2(new_n6403_), .A3(new_n6475_), .ZN(new_n6478_));
  OAI21_X1   g05466(.A1(new_n6477_), .A2(new_n6478_), .B(new_n6390_), .ZN(new_n6479_));
  INV_X1     g05467(.I(new_n6390_), .ZN(new_n6480_));
  OAI21_X1   g05468(.A1(new_n6389_), .A2(new_n6403_), .B(new_n6475_), .ZN(new_n6481_));
  NAND3_X1   g05469(.A1(new_n6468_), .A2(new_n6474_), .A3(new_n6476_), .ZN(new_n6482_));
  NAND3_X1   g05470(.A1(new_n6481_), .A2(new_n6482_), .A3(new_n6480_), .ZN(new_n6483_));
  NAND2_X1   g05471(.A1(new_n6479_), .A2(new_n6483_), .ZN(new_n6484_));
  NAND2_X1   g05472(.A1(new_n6415_), .A2(new_n6453_), .ZN(new_n6485_));
  NAND2_X1   g05473(.A1(new_n6426_), .A2(new_n6447_), .ZN(new_n6486_));
  NAND2_X1   g05474(.A1(new_n6485_), .A2(new_n6486_), .ZN(new_n6487_));
  NAND2_X1   g05475(.A1(new_n6404_), .A2(new_n6487_), .ZN(new_n6488_));
  NAND2_X1   g05476(.A1(new_n6390_), .A2(new_n6475_), .ZN(new_n6489_));
  AOI21_X1   g05477(.A1(new_n6389_), .A2(new_n6403_), .B(new_n6489_), .ZN(new_n6490_));
  NOR4_X1    g05478(.A1(new_n6484_), .A2(new_n6488_), .A3(new_n6462_), .A4(new_n6490_), .ZN(new_n6491_));
  XOR2_X1    g05479(.A1(new_n6468_), .A2(new_n6403_), .Z(new_n6492_));
  NOR2_X1    g05480(.A1(new_n6426_), .A2(new_n6447_), .ZN(new_n6493_));
  NOR2_X1    g05481(.A1(new_n6415_), .A2(new_n6453_), .ZN(new_n6494_));
  NOR2_X1    g05482(.A1(new_n6493_), .A2(new_n6494_), .ZN(new_n6495_));
  NAND3_X1   g05483(.A1(new_n6392_), .A2(new_n6439_), .A3(new_n6430_), .ZN(new_n6496_));
  NOR3_X1    g05484(.A1(new_n6492_), .A2(new_n6495_), .A3(new_n6496_), .ZN(new_n6497_));
  NAND2_X1   g05485(.A1(new_n6497_), .A2(new_n6461_), .ZN(new_n6498_));
  AOI21_X1   g05486(.A1(new_n6481_), .A2(new_n6482_), .B(new_n6480_), .ZN(new_n6499_));
  NOR3_X1    g05487(.A1(new_n6477_), .A2(new_n6478_), .A3(new_n6390_), .ZN(new_n6500_));
  NOR2_X1    g05488(.A1(new_n6500_), .A2(new_n6499_), .ZN(new_n6501_));
  OAI21_X1   g05489(.A1(new_n6461_), .A2(new_n6497_), .B(new_n6501_), .ZN(new_n6502_));
  AOI21_X1   g05490(.A1(new_n6458_), .A2(new_n6459_), .B(new_n6456_), .ZN(new_n6503_));
  NOR3_X1    g05491(.A1(new_n6441_), .A2(new_n6454_), .A3(new_n6427_), .ZN(new_n6504_));
  NOR2_X1    g05492(.A1(new_n6504_), .A2(new_n6503_), .ZN(new_n6505_));
  NOR2_X1    g05493(.A1(new_n6457_), .A2(new_n6429_), .ZN(new_n6506_));
  NAND4_X1   g05494(.A1(new_n6404_), .A2(new_n6392_), .A3(new_n6487_), .A4(new_n6506_), .ZN(new_n6507_));
  NAND3_X1   g05495(.A1(new_n6507_), .A2(new_n6505_), .A3(new_n6484_), .ZN(new_n6508_));
  NAND2_X1   g05496(.A1(new_n6502_), .A2(new_n6508_), .ZN(new_n6509_));
  AOI22_X1   g05497(.A1(new_n6509_), .A2(new_n6498_), .B1(new_n6461_), .B2(new_n6491_), .ZN(new_n6510_));
  OAI22_X1   g05498(.A1(new_n6510_), .A2(new_n6355_), .B1(new_n6433_), .B2(new_n6438_), .ZN(new_n6511_));
  OAI21_X1   g05499(.A1(new_n6234_), .A2(new_n6239_), .B(new_n6272_), .ZN(new_n6512_));
  NAND2_X1   g05500(.A1(new_n6512_), .A2(new_n6320_), .ZN(new_n6513_));
  OAI21_X1   g05501(.A1(new_n6316_), .A2(new_n6317_), .B(new_n6325_), .ZN(new_n6514_));
  NAND2_X1   g05502(.A1(new_n6514_), .A2(new_n6318_), .ZN(new_n6515_));
  INV_X1     g05503(.I(new_n6515_), .ZN(new_n6516_));
  OAI21_X1   g05504(.A1(new_n6337_), .A2(new_n6343_), .B(new_n6334_), .ZN(new_n6517_));
  AOI21_X1   g05505(.A1(new_n6517_), .A2(new_n6358_), .B(new_n6516_), .ZN(new_n6518_));
  AOI21_X1   g05506(.A1(new_n6362_), .A2(new_n6366_), .B(new_n6361_), .ZN(new_n6519_));
  NOR3_X1    g05507(.A1(new_n6519_), .A2(new_n6324_), .A3(new_n6515_), .ZN(new_n6520_));
  OAI21_X1   g05508(.A1(new_n6520_), .A2(new_n6518_), .B(new_n6513_), .ZN(new_n6521_));
  INV_X1     g05509(.I(new_n6513_), .ZN(new_n6522_));
  OAI21_X1   g05510(.A1(new_n6519_), .A2(new_n6324_), .B(new_n6515_), .ZN(new_n6523_));
  NAND3_X1   g05511(.A1(new_n6517_), .A2(new_n6358_), .A3(new_n6516_), .ZN(new_n6524_));
  NAND3_X1   g05512(.A1(new_n6523_), .A2(new_n6524_), .A3(new_n6522_), .ZN(new_n6525_));
  NAND2_X1   g05513(.A1(new_n6521_), .A2(new_n6525_), .ZN(new_n6526_));
  NAND2_X1   g05514(.A1(new_n6480_), .A2(new_n6476_), .ZN(new_n6527_));
  NAND3_X1   g05515(.A1(new_n6527_), .A2(new_n6468_), .A3(new_n6474_), .ZN(new_n6528_));
  NAND2_X1   g05516(.A1(new_n6528_), .A2(new_n6489_), .ZN(new_n6529_));
  INV_X1     g05517(.I(new_n6529_), .ZN(new_n6530_));
  OAI21_X1   g05518(.A1(new_n6427_), .A2(new_n6428_), .B(new_n6439_), .ZN(new_n6531_));
  NAND2_X1   g05519(.A1(new_n6531_), .A2(new_n6429_), .ZN(new_n6532_));
  AOI21_X1   g05520(.A1(new_n6501_), .A2(new_n6507_), .B(new_n6505_), .ZN(new_n6533_));
  OAI21_X1   g05521(.A1(new_n6533_), .A2(new_n6491_), .B(new_n6532_), .ZN(new_n6534_));
  NOR2_X1    g05522(.A1(new_n6492_), .A2(new_n6495_), .ZN(new_n6535_));
  NOR2_X1    g05523(.A1(new_n6462_), .A2(new_n6490_), .ZN(new_n6536_));
  NAND3_X1   g05524(.A1(new_n6501_), .A2(new_n6535_), .A3(new_n6536_), .ZN(new_n6537_));
  INV_X1     g05525(.I(new_n6532_), .ZN(new_n6538_));
  OAI21_X1   g05526(.A1(new_n6484_), .A2(new_n6497_), .B(new_n6461_), .ZN(new_n6539_));
  NAND3_X1   g05527(.A1(new_n6539_), .A2(new_n6537_), .A3(new_n6538_), .ZN(new_n6540_));
  AOI21_X1   g05528(.A1(new_n6534_), .A2(new_n6540_), .B(new_n6530_), .ZN(new_n6541_));
  AOI21_X1   g05529(.A1(new_n6539_), .A2(new_n6537_), .B(new_n6538_), .ZN(new_n6542_));
  NOR3_X1    g05530(.A1(new_n6533_), .A2(new_n6491_), .A3(new_n6532_), .ZN(new_n6543_));
  NOR3_X1    g05531(.A1(new_n6543_), .A2(new_n6542_), .A3(new_n6529_), .ZN(new_n6544_));
  NOR2_X1    g05532(.A1(new_n6544_), .A2(new_n6541_), .ZN(new_n6545_));
  NAND2_X1   g05533(.A1(new_n6545_), .A2(new_n6526_), .ZN(new_n6546_));
  AOI21_X1   g05534(.A1(new_n6523_), .A2(new_n6524_), .B(new_n6522_), .ZN(new_n6547_));
  NOR3_X1    g05535(.A1(new_n6520_), .A2(new_n6518_), .A3(new_n6513_), .ZN(new_n6548_));
  NOR2_X1    g05536(.A1(new_n6548_), .A2(new_n6547_), .ZN(new_n6549_));
  OAI21_X1   g05537(.A1(new_n6543_), .A2(new_n6542_), .B(new_n6529_), .ZN(new_n6550_));
  NAND3_X1   g05538(.A1(new_n6534_), .A2(new_n6540_), .A3(new_n6530_), .ZN(new_n6551_));
  NAND2_X1   g05539(.A1(new_n6550_), .A2(new_n6551_), .ZN(new_n6552_));
  NAND2_X1   g05540(.A1(new_n6549_), .A2(new_n6552_), .ZN(new_n6553_));
  AOI21_X1   g05541(.A1(new_n6546_), .A2(new_n6553_), .B(new_n6511_), .ZN(new_n6554_));
  NAND2_X1   g05542(.A1(new_n6368_), .A2(new_n6371_), .ZN(new_n6555_));
  OAI21_X1   g05543(.A1(new_n6345_), .A2(new_n6354_), .B(new_n6437_), .ZN(new_n6556_));
  NAND3_X1   g05544(.A1(new_n6368_), .A2(new_n6432_), .A3(new_n6371_), .ZN(new_n6557_));
  NAND2_X1   g05545(.A1(new_n6491_), .A2(new_n6461_), .ZN(new_n6558_));
  AOI21_X1   g05546(.A1(new_n6507_), .A2(new_n6505_), .B(new_n6484_), .ZN(new_n6559_));
  NOR3_X1    g05547(.A1(new_n6501_), .A2(new_n6497_), .A3(new_n6461_), .ZN(new_n6560_));
  OAI21_X1   g05548(.A1(new_n6560_), .A2(new_n6559_), .B(new_n6498_), .ZN(new_n6561_));
  NAND2_X1   g05549(.A1(new_n6561_), .A2(new_n6558_), .ZN(new_n6562_));
  AOI22_X1   g05550(.A1(new_n6562_), .A2(new_n6555_), .B1(new_n6556_), .B2(new_n6557_), .ZN(new_n6563_));
  NAND4_X1   g05551(.A1(new_n6521_), .A2(new_n6525_), .A3(new_n6550_), .A4(new_n6551_), .ZN(new_n6564_));
  OAI22_X1   g05552(.A1(new_n6547_), .A2(new_n6548_), .B1(new_n6544_), .B2(new_n6541_), .ZN(new_n6565_));
  AOI21_X1   g05553(.A1(new_n6565_), .A2(new_n6564_), .B(new_n6563_), .ZN(new_n6566_));
  NOR3_X1    g05554(.A1(new_n6554_), .A2(new_n6230_), .A3(new_n6566_), .ZN(new_n6567_));
  NOR3_X1    g05555(.A1(new_n6562_), .A2(new_n6433_), .A3(new_n6438_), .ZN(new_n6568_));
  INV_X1     g05556(.I(new_n6568_), .ZN(new_n6569_));
  NAND2_X1   g05557(.A1(new_n6374_), .A2(new_n6378_), .ZN(new_n6570_));
  INV_X1     g05558(.I(new_n6392_), .ZN(new_n6571_));
  NOR2_X1    g05559(.A1(new_n6492_), .A2(new_n6571_), .ZN(new_n6572_));
  INV_X1     g05560(.I(new_n6572_), .ZN(new_n6573_));
  AND2_X2    g05561(.A1(new_n6570_), .A2(new_n6573_), .Z(new_n6574_));
  NOR2_X1    g05562(.A1(new_n6570_), .A2(new_n6573_), .ZN(new_n6575_));
  NOR2_X1    g05563(.A1(new_n6032_), .A2(new_n6039_), .ZN(new_n6576_));
  NOR2_X1    g05564(.A1(new_n6576_), .A2(new_n6195_), .ZN(new_n6577_));
  AND2_X2    g05565(.A1(new_n6576_), .A2(new_n6195_), .Z(new_n6578_));
  NOR4_X1    g05566(.A1(new_n6574_), .A2(new_n6575_), .A3(new_n6578_), .A4(new_n6577_), .ZN(new_n6579_));
  NOR2_X1    g05567(.A1(new_n6568_), .A2(new_n6579_), .ZN(new_n6580_));
  INV_X1     g05568(.I(new_n6580_), .ZN(new_n6581_));
  NAND2_X1   g05569(.A1(new_n6568_), .A2(new_n6579_), .ZN(new_n6582_));
  NAND3_X1   g05570(.A1(new_n6219_), .A2(new_n6168_), .A3(new_n6184_), .ZN(new_n6583_));
  NAND2_X1   g05571(.A1(new_n6185_), .A2(new_n6131_), .ZN(new_n6584_));
  NAND2_X1   g05572(.A1(new_n6584_), .A2(new_n6583_), .ZN(new_n6585_));
  AOI22_X1   g05573(.A1(new_n6581_), .A2(new_n6582_), .B1(new_n6569_), .B2(new_n6585_), .ZN(new_n6586_));
  OAI21_X1   g05574(.A1(new_n6554_), .A2(new_n6566_), .B(new_n6230_), .ZN(new_n6587_));
  AOI21_X1   g05575(.A1(new_n6587_), .A2(new_n6586_), .B(new_n6567_), .ZN(new_n6588_));
  NOR2_X1    g05576(.A1(new_n6522_), .A2(new_n6516_), .ZN(new_n6589_));
  NAND2_X1   g05577(.A1(new_n6517_), .A2(new_n6358_), .ZN(new_n6590_));
  AOI21_X1   g05578(.A1(new_n6522_), .A2(new_n6516_), .B(new_n6590_), .ZN(new_n6591_));
  NOR2_X1    g05579(.A1(new_n6591_), .A2(new_n6589_), .ZN(new_n6592_));
  AOI21_X1   g05580(.A1(new_n6549_), .A2(new_n6545_), .B(new_n6563_), .ZN(new_n6593_));
  NAND2_X1   g05581(.A1(new_n6539_), .A2(new_n6537_), .ZN(new_n6594_));
  XOR2_X1    g05582(.A1(new_n6515_), .A2(new_n6513_), .Z(new_n6595_));
  XOR2_X1    g05583(.A1(new_n6532_), .A2(new_n6529_), .Z(new_n6596_));
  NOR4_X1    g05584(.A1(new_n6590_), .A2(new_n6594_), .A3(new_n6596_), .A4(new_n6595_), .ZN(new_n6597_));
  INV_X1     g05585(.I(new_n6597_), .ZN(new_n6598_));
  NOR2_X1    g05586(.A1(new_n6538_), .A2(new_n6530_), .ZN(new_n6599_));
  AOI21_X1   g05587(.A1(new_n6530_), .A2(new_n6538_), .B(new_n6594_), .ZN(new_n6600_));
  NOR2_X1    g05588(.A1(new_n6600_), .A2(new_n6599_), .ZN(new_n6601_));
  INV_X1     g05589(.I(new_n6601_), .ZN(new_n6602_));
  OAI21_X1   g05590(.A1(new_n6593_), .A2(new_n6598_), .B(new_n6602_), .ZN(new_n6603_));
  NAND2_X1   g05591(.A1(new_n6564_), .A2(new_n6511_), .ZN(new_n6604_));
  NAND3_X1   g05592(.A1(new_n6604_), .A2(new_n6597_), .A3(new_n6601_), .ZN(new_n6605_));
  AOI21_X1   g05593(.A1(new_n6603_), .A2(new_n6605_), .B(new_n6592_), .ZN(new_n6606_));
  INV_X1     g05594(.I(new_n6592_), .ZN(new_n6607_));
  AOI21_X1   g05595(.A1(new_n6604_), .A2(new_n6597_), .B(new_n6601_), .ZN(new_n6608_));
  NOR3_X1    g05596(.A1(new_n6593_), .A2(new_n6598_), .A3(new_n6602_), .ZN(new_n6609_));
  NOR3_X1    g05597(.A1(new_n6609_), .A2(new_n6608_), .A3(new_n6607_), .ZN(new_n6610_));
  NAND2_X1   g05598(.A1(new_n6192_), .A2(new_n6190_), .ZN(new_n6611_));
  OR2_X2     g05599(.A1(new_n6192_), .A2(new_n6190_), .Z(new_n6612_));
  NAND3_X1   g05600(.A1(new_n6188_), .A2(new_n6187_), .A3(new_n6612_), .ZN(new_n6613_));
  NAND2_X1   g05601(.A1(new_n6613_), .A2(new_n6611_), .ZN(new_n6614_));
  INV_X1     g05602(.I(new_n6614_), .ZN(new_n6615_));
  NAND2_X1   g05603(.A1(new_n6121_), .A2(new_n6128_), .ZN(new_n6616_));
  OAI21_X1   g05604(.A1(new_n6185_), .A2(new_n6131_), .B(new_n6616_), .ZN(new_n6617_));
  INV_X1     g05605(.I(new_n6214_), .ZN(new_n6618_));
  NAND3_X1   g05606(.A1(new_n6617_), .A2(new_n6209_), .A3(new_n6618_), .ZN(new_n6619_));
  OAI21_X1   g05607(.A1(new_n6204_), .A2(new_n6156_), .B(new_n6202_), .ZN(new_n6620_));
  NAND3_X1   g05608(.A1(new_n6199_), .A2(new_n6198_), .A3(new_n6205_), .ZN(new_n6621_));
  NAND2_X1   g05609(.A1(new_n6197_), .A2(new_n6621_), .ZN(new_n6622_));
  NAND2_X1   g05610(.A1(new_n6622_), .A2(new_n6620_), .ZN(new_n6623_));
  NAND2_X1   g05611(.A1(new_n6619_), .A2(new_n6623_), .ZN(new_n6624_));
  INV_X1     g05612(.I(new_n6227_), .ZN(new_n6625_));
  NAND3_X1   g05613(.A1(new_n6583_), .A2(new_n6616_), .A3(new_n6226_), .ZN(new_n6626_));
  INV_X1     g05614(.I(new_n6623_), .ZN(new_n6627_));
  NAND3_X1   g05615(.A1(new_n6626_), .A2(new_n6627_), .A3(new_n6625_), .ZN(new_n6628_));
  AOI21_X1   g05616(.A1(new_n6624_), .A2(new_n6628_), .B(new_n6615_), .ZN(new_n6629_));
  AOI21_X1   g05617(.A1(new_n6626_), .A2(new_n6625_), .B(new_n6627_), .ZN(new_n6630_));
  NOR4_X1    g05618(.A1(new_n6225_), .A2(new_n6194_), .A3(new_n6214_), .A4(new_n6623_), .ZN(new_n6631_));
  NOR3_X1    g05619(.A1(new_n6630_), .A2(new_n6631_), .A3(new_n6614_), .ZN(new_n6632_));
  NOR2_X1    g05620(.A1(new_n6629_), .A2(new_n6632_), .ZN(new_n6633_));
  OAI21_X1   g05621(.A1(new_n6606_), .A2(new_n6610_), .B(new_n6633_), .ZN(new_n6634_));
  OAI21_X1   g05622(.A1(new_n6609_), .A2(new_n6608_), .B(new_n6607_), .ZN(new_n6635_));
  NAND3_X1   g05623(.A1(new_n6603_), .A2(new_n6605_), .A3(new_n6592_), .ZN(new_n6636_));
  OAI21_X1   g05624(.A1(new_n6630_), .A2(new_n6631_), .B(new_n6614_), .ZN(new_n6637_));
  NAND3_X1   g05625(.A1(new_n6624_), .A2(new_n6628_), .A3(new_n6615_), .ZN(new_n6638_));
  NAND2_X1   g05626(.A1(new_n6638_), .A2(new_n6637_), .ZN(new_n6639_));
  NAND3_X1   g05627(.A1(new_n6639_), .A2(new_n6635_), .A3(new_n6636_), .ZN(new_n6640_));
  AOI21_X1   g05628(.A1(new_n6634_), .A2(new_n6640_), .B(new_n6588_), .ZN(new_n6641_));
  NOR2_X1    g05629(.A1(new_n6215_), .A2(new_n6208_), .ZN(new_n6642_));
  NOR2_X1    g05630(.A1(new_n6225_), .A2(new_n6642_), .ZN(new_n6643_));
  AOI21_X1   g05631(.A1(new_n6226_), .A2(new_n6227_), .B(new_n6617_), .ZN(new_n6644_));
  NOR2_X1    g05632(.A1(new_n6643_), .A2(new_n6644_), .ZN(new_n6645_));
  NOR2_X1    g05633(.A1(new_n6549_), .A2(new_n6552_), .ZN(new_n6646_));
  NOR2_X1    g05634(.A1(new_n6545_), .A2(new_n6526_), .ZN(new_n6647_));
  OAI21_X1   g05635(.A1(new_n6647_), .A2(new_n6646_), .B(new_n6563_), .ZN(new_n6648_));
  NOR2_X1    g05636(.A1(new_n6526_), .A2(new_n6552_), .ZN(new_n6649_));
  AOI22_X1   g05637(.A1(new_n6521_), .A2(new_n6525_), .B1(new_n6550_), .B2(new_n6551_), .ZN(new_n6650_));
  OAI21_X1   g05638(.A1(new_n6649_), .A2(new_n6650_), .B(new_n6511_), .ZN(new_n6651_));
  NAND3_X1   g05639(.A1(new_n6648_), .A2(new_n6645_), .A3(new_n6651_), .ZN(new_n6652_));
  INV_X1     g05640(.I(new_n6586_), .ZN(new_n6653_));
  AOI21_X1   g05641(.A1(new_n6648_), .A2(new_n6651_), .B(new_n6645_), .ZN(new_n6654_));
  OAI21_X1   g05642(.A1(new_n6654_), .A2(new_n6653_), .B(new_n6652_), .ZN(new_n6655_));
  NAND3_X1   g05643(.A1(new_n6633_), .A2(new_n6635_), .A3(new_n6636_), .ZN(new_n6656_));
  OAI21_X1   g05644(.A1(new_n6606_), .A2(new_n6610_), .B(new_n6639_), .ZN(new_n6657_));
  AOI21_X1   g05645(.A1(new_n6657_), .A2(new_n6656_), .B(new_n6655_), .ZN(new_n6658_));
  INV_X1     g05646(.I(\A[190] ), .ZN(new_n6659_));
  NOR2_X1    g05647(.A1(\A[191] ), .A2(\A[192] ), .ZN(new_n6660_));
  NAND2_X1   g05648(.A1(\A[191] ), .A2(\A[192] ), .ZN(new_n6661_));
  AOI21_X1   g05649(.A1(new_n6659_), .A2(new_n6661_), .B(new_n6660_), .ZN(new_n6662_));
  INV_X1     g05650(.I(\A[187] ), .ZN(new_n6663_));
  NOR2_X1    g05651(.A1(\A[188] ), .A2(\A[189] ), .ZN(new_n6664_));
  NAND2_X1   g05652(.A1(\A[188] ), .A2(\A[189] ), .ZN(new_n6665_));
  AOI21_X1   g05653(.A1(new_n6663_), .A2(new_n6665_), .B(new_n6664_), .ZN(new_n6666_));
  INV_X1     g05654(.I(new_n6666_), .ZN(new_n6667_));
  INV_X1     g05655(.I(\A[188] ), .ZN(new_n6668_));
  NAND2_X1   g05656(.A1(new_n6668_), .A2(\A[189] ), .ZN(new_n6669_));
  INV_X1     g05657(.I(\A[189] ), .ZN(new_n6670_));
  NAND2_X1   g05658(.A1(new_n6670_), .A2(\A[188] ), .ZN(new_n6671_));
  AOI21_X1   g05659(.A1(new_n6669_), .A2(new_n6671_), .B(new_n6663_), .ZN(new_n6672_));
  INV_X1     g05660(.I(new_n6664_), .ZN(new_n6673_));
  AOI21_X1   g05661(.A1(new_n6673_), .A2(new_n6665_), .B(\A[187] ), .ZN(new_n6674_));
  INV_X1     g05662(.I(\A[191] ), .ZN(new_n6675_));
  NAND2_X1   g05663(.A1(new_n6675_), .A2(\A[192] ), .ZN(new_n6676_));
  INV_X1     g05664(.I(\A[192] ), .ZN(new_n6677_));
  NAND2_X1   g05665(.A1(new_n6677_), .A2(\A[191] ), .ZN(new_n6678_));
  AOI21_X1   g05666(.A1(new_n6676_), .A2(new_n6678_), .B(new_n6659_), .ZN(new_n6679_));
  INV_X1     g05667(.I(new_n6660_), .ZN(new_n6680_));
  AOI21_X1   g05668(.A1(new_n6680_), .A2(new_n6661_), .B(\A[190] ), .ZN(new_n6681_));
  NOR4_X1    g05669(.A1(new_n6672_), .A2(new_n6674_), .A3(new_n6681_), .A4(new_n6679_), .ZN(new_n6682_));
  NOR2_X1    g05670(.A1(new_n6682_), .A2(new_n6667_), .ZN(new_n6683_));
  NOR2_X1    g05671(.A1(new_n6670_), .A2(\A[188] ), .ZN(new_n6684_));
  NOR2_X1    g05672(.A1(new_n6668_), .A2(\A[189] ), .ZN(new_n6685_));
  OAI21_X1   g05673(.A1(new_n6684_), .A2(new_n6685_), .B(\A[187] ), .ZN(new_n6686_));
  INV_X1     g05674(.I(new_n6665_), .ZN(new_n6687_));
  OAI21_X1   g05675(.A1(new_n6687_), .A2(new_n6664_), .B(new_n6663_), .ZN(new_n6688_));
  NOR2_X1    g05676(.A1(new_n6677_), .A2(\A[191] ), .ZN(new_n6689_));
  NOR2_X1    g05677(.A1(new_n6675_), .A2(\A[192] ), .ZN(new_n6690_));
  OAI21_X1   g05678(.A1(new_n6689_), .A2(new_n6690_), .B(\A[190] ), .ZN(new_n6691_));
  INV_X1     g05679(.I(new_n6661_), .ZN(new_n6692_));
  OAI21_X1   g05680(.A1(new_n6692_), .A2(new_n6660_), .B(new_n6659_), .ZN(new_n6693_));
  NAND4_X1   g05681(.A1(new_n6686_), .A2(new_n6688_), .A3(new_n6691_), .A4(new_n6693_), .ZN(new_n6694_));
  NOR2_X1    g05682(.A1(new_n6694_), .A2(new_n6666_), .ZN(new_n6695_));
  OAI21_X1   g05683(.A1(new_n6683_), .A2(new_n6695_), .B(new_n6662_), .ZN(new_n6696_));
  INV_X1     g05684(.I(new_n6662_), .ZN(new_n6697_));
  NAND2_X1   g05685(.A1(new_n6694_), .A2(new_n6666_), .ZN(new_n6698_));
  NOR2_X1    g05686(.A1(new_n6681_), .A2(new_n6679_), .ZN(new_n6699_));
  NAND4_X1   g05687(.A1(new_n6699_), .A2(new_n6667_), .A3(new_n6686_), .A4(new_n6688_), .ZN(new_n6700_));
  NAND3_X1   g05688(.A1(new_n6698_), .A2(new_n6700_), .A3(new_n6697_), .ZN(new_n6701_));
  NAND2_X1   g05689(.A1(new_n6696_), .A2(new_n6701_), .ZN(new_n6702_));
  INV_X1     g05690(.I(new_n6702_), .ZN(new_n6703_));
  INV_X1     g05691(.I(\A[196] ), .ZN(new_n6704_));
  NOR2_X1    g05692(.A1(\A[197] ), .A2(\A[198] ), .ZN(new_n6705_));
  NAND2_X1   g05693(.A1(\A[197] ), .A2(\A[198] ), .ZN(new_n6706_));
  AOI21_X1   g05694(.A1(new_n6704_), .A2(new_n6706_), .B(new_n6705_), .ZN(new_n6707_));
  INV_X1     g05695(.I(\A[193] ), .ZN(new_n6708_));
  NOR2_X1    g05696(.A1(\A[194] ), .A2(\A[195] ), .ZN(new_n6709_));
  NAND2_X1   g05697(.A1(\A[194] ), .A2(\A[195] ), .ZN(new_n6710_));
  AOI21_X1   g05698(.A1(new_n6708_), .A2(new_n6710_), .B(new_n6709_), .ZN(new_n6711_));
  NAND2_X1   g05699(.A1(new_n6707_), .A2(new_n6711_), .ZN(new_n6712_));
  INV_X1     g05700(.I(\A[194] ), .ZN(new_n6713_));
  NAND2_X1   g05701(.A1(new_n6713_), .A2(\A[195] ), .ZN(new_n6714_));
  INV_X1     g05702(.I(\A[195] ), .ZN(new_n6715_));
  NAND2_X1   g05703(.A1(new_n6715_), .A2(\A[194] ), .ZN(new_n6716_));
  AOI21_X1   g05704(.A1(new_n6714_), .A2(new_n6716_), .B(new_n6708_), .ZN(new_n6717_));
  INV_X1     g05705(.I(new_n6709_), .ZN(new_n6718_));
  AOI21_X1   g05706(.A1(new_n6718_), .A2(new_n6710_), .B(\A[193] ), .ZN(new_n6719_));
  NOR2_X1    g05707(.A1(new_n6719_), .A2(new_n6717_), .ZN(new_n6720_));
  INV_X1     g05708(.I(\A[198] ), .ZN(new_n6721_));
  NOR2_X1    g05709(.A1(new_n6721_), .A2(\A[197] ), .ZN(new_n6722_));
  INV_X1     g05710(.I(\A[197] ), .ZN(new_n6723_));
  NOR2_X1    g05711(.A1(new_n6723_), .A2(\A[198] ), .ZN(new_n6724_));
  OAI21_X1   g05712(.A1(new_n6722_), .A2(new_n6724_), .B(\A[196] ), .ZN(new_n6725_));
  INV_X1     g05713(.I(new_n6706_), .ZN(new_n6726_));
  OAI21_X1   g05714(.A1(new_n6726_), .A2(new_n6705_), .B(new_n6704_), .ZN(new_n6727_));
  NAND2_X1   g05715(.A1(new_n6725_), .A2(new_n6727_), .ZN(new_n6728_));
  NAND2_X1   g05716(.A1(new_n6720_), .A2(new_n6728_), .ZN(new_n6729_));
  NOR2_X1    g05717(.A1(new_n6715_), .A2(\A[194] ), .ZN(new_n6730_));
  NOR2_X1    g05718(.A1(new_n6713_), .A2(\A[195] ), .ZN(new_n6731_));
  OAI21_X1   g05719(.A1(new_n6730_), .A2(new_n6731_), .B(\A[193] ), .ZN(new_n6732_));
  INV_X1     g05720(.I(new_n6710_), .ZN(new_n6733_));
  OAI21_X1   g05721(.A1(new_n6733_), .A2(new_n6709_), .B(new_n6708_), .ZN(new_n6734_));
  NAND2_X1   g05722(.A1(new_n6732_), .A2(new_n6734_), .ZN(new_n6735_));
  NAND2_X1   g05723(.A1(new_n6723_), .A2(\A[198] ), .ZN(new_n6736_));
  NAND2_X1   g05724(.A1(new_n6721_), .A2(\A[197] ), .ZN(new_n6737_));
  AOI21_X1   g05725(.A1(new_n6736_), .A2(new_n6737_), .B(new_n6704_), .ZN(new_n6738_));
  INV_X1     g05726(.I(new_n6705_), .ZN(new_n6739_));
  AOI21_X1   g05727(.A1(new_n6739_), .A2(new_n6706_), .B(\A[196] ), .ZN(new_n6740_));
  NOR2_X1    g05728(.A1(new_n6740_), .A2(new_n6738_), .ZN(new_n6741_));
  NAND2_X1   g05729(.A1(new_n6741_), .A2(new_n6735_), .ZN(new_n6742_));
  AOI21_X1   g05730(.A1(new_n6729_), .A2(new_n6742_), .B(new_n6712_), .ZN(new_n6743_));
  INV_X1     g05731(.I(new_n6707_), .ZN(new_n6744_));
  NAND4_X1   g05732(.A1(new_n6732_), .A2(new_n6734_), .A3(new_n6725_), .A4(new_n6727_), .ZN(new_n6745_));
  NAND2_X1   g05733(.A1(new_n6745_), .A2(new_n6711_), .ZN(new_n6746_));
  INV_X1     g05734(.I(new_n6711_), .ZN(new_n6747_));
  NAND3_X1   g05735(.A1(new_n6720_), .A2(new_n6741_), .A3(new_n6747_), .ZN(new_n6748_));
  AOI21_X1   g05736(.A1(new_n6746_), .A2(new_n6748_), .B(new_n6744_), .ZN(new_n6749_));
  AOI21_X1   g05737(.A1(new_n6720_), .A2(new_n6741_), .B(new_n6747_), .ZN(new_n6750_));
  NOR3_X1    g05738(.A1(new_n6735_), .A2(new_n6728_), .A3(new_n6711_), .ZN(new_n6751_));
  NOR3_X1    g05739(.A1(new_n6750_), .A2(new_n6751_), .A3(new_n6707_), .ZN(new_n6752_));
  NOR2_X1    g05740(.A1(new_n6745_), .A2(new_n6712_), .ZN(new_n6753_));
  NOR4_X1    g05741(.A1(new_n6717_), .A2(new_n6719_), .A3(new_n6740_), .A4(new_n6738_), .ZN(new_n6754_));
  AOI22_X1   g05742(.A1(new_n6732_), .A2(new_n6734_), .B1(new_n6725_), .B2(new_n6727_), .ZN(new_n6755_));
  NOR2_X1    g05743(.A1(new_n6755_), .A2(new_n6754_), .ZN(new_n6756_));
  AOI22_X1   g05744(.A1(new_n6686_), .A2(new_n6688_), .B1(new_n6691_), .B2(new_n6693_), .ZN(new_n6757_));
  NOR2_X1    g05745(.A1(new_n6757_), .A2(new_n6682_), .ZN(new_n6758_));
  NAND2_X1   g05746(.A1(new_n6662_), .A2(new_n6666_), .ZN(new_n6759_));
  NOR2_X1    g05747(.A1(new_n6694_), .A2(new_n6759_), .ZN(new_n6760_));
  NAND4_X1   g05748(.A1(new_n6756_), .A2(new_n6758_), .A3(new_n6753_), .A4(new_n6760_), .ZN(new_n6761_));
  NOR4_X1    g05749(.A1(new_n6761_), .A2(new_n6743_), .A3(new_n6749_), .A4(new_n6752_), .ZN(new_n6762_));
  NOR3_X1    g05750(.A1(new_n6749_), .A2(new_n6752_), .A3(new_n6743_), .ZN(new_n6763_));
  INV_X1     g05751(.I(new_n6712_), .ZN(new_n6764_));
  NAND2_X1   g05752(.A1(new_n6754_), .A2(new_n6764_), .ZN(new_n6765_));
  OR2_X2     g05753(.A1(new_n6755_), .A2(new_n6754_), .Z(new_n6766_));
  OAI22_X1   g05754(.A1(new_n6672_), .A2(new_n6674_), .B1(new_n6681_), .B2(new_n6679_), .ZN(new_n6767_));
  NAND2_X1   g05755(.A1(new_n6767_), .A2(new_n6694_), .ZN(new_n6768_));
  NAND3_X1   g05756(.A1(new_n6682_), .A2(new_n6662_), .A3(new_n6666_), .ZN(new_n6769_));
  NOR4_X1    g05757(.A1(new_n6766_), .A2(new_n6768_), .A3(new_n6765_), .A4(new_n6769_), .ZN(new_n6770_));
  NOR2_X1    g05758(.A1(new_n6763_), .A2(new_n6770_), .ZN(new_n6771_));
  OAI21_X1   g05759(.A1(new_n6771_), .A2(new_n6762_), .B(new_n6703_), .ZN(new_n6772_));
  OAI21_X1   g05760(.A1(new_n6750_), .A2(new_n6751_), .B(new_n6707_), .ZN(new_n6773_));
  NAND3_X1   g05761(.A1(new_n6746_), .A2(new_n6748_), .A3(new_n6744_), .ZN(new_n6774_));
  NAND2_X1   g05762(.A1(new_n6773_), .A2(new_n6774_), .ZN(new_n6775_));
  OAI21_X1   g05763(.A1(new_n6775_), .A2(new_n6743_), .B(new_n6770_), .ZN(new_n6776_));
  NOR4_X1    g05764(.A1(new_n6682_), .A2(new_n6757_), .A3(new_n6745_), .A4(new_n6712_), .ZN(new_n6777_));
  NAND2_X1   g05765(.A1(new_n6777_), .A2(new_n6756_), .ZN(new_n6778_));
  NOR2_X1    g05766(.A1(new_n6743_), .A2(new_n6769_), .ZN(new_n6779_));
  OAI21_X1   g05767(.A1(new_n6775_), .A2(new_n6778_), .B(new_n6779_), .ZN(new_n6780_));
  NAND3_X1   g05768(.A1(new_n6776_), .A2(new_n6780_), .A3(new_n6703_), .ZN(new_n6781_));
  NAND2_X1   g05769(.A1(new_n6781_), .A2(new_n6772_), .ZN(new_n6782_));
  NAND2_X1   g05770(.A1(new_n6763_), .A2(new_n6770_), .ZN(new_n6783_));
  OAI21_X1   g05771(.A1(new_n6775_), .A2(new_n6743_), .B(new_n6761_), .ZN(new_n6784_));
  AOI21_X1   g05772(.A1(new_n6784_), .A2(new_n6783_), .B(new_n6702_), .ZN(new_n6785_));
  NOR2_X1    g05773(.A1(new_n6763_), .A2(new_n6761_), .ZN(new_n6786_));
  NOR2_X1    g05774(.A1(new_n6749_), .A2(new_n6752_), .ZN(new_n6787_));
  NOR3_X1    g05775(.A1(new_n6766_), .A2(new_n6768_), .A3(new_n6765_), .ZN(new_n6788_));
  NOR2_X1    g05776(.A1(new_n6741_), .A2(new_n6735_), .ZN(new_n6789_));
  NOR2_X1    g05777(.A1(new_n6720_), .A2(new_n6728_), .ZN(new_n6790_));
  OAI21_X1   g05778(.A1(new_n6789_), .A2(new_n6790_), .B(new_n6764_), .ZN(new_n6791_));
  NAND2_X1   g05779(.A1(new_n6791_), .A2(new_n6760_), .ZN(new_n6792_));
  AOI21_X1   g05780(.A1(new_n6787_), .A2(new_n6788_), .B(new_n6792_), .ZN(new_n6793_));
  NOR3_X1    g05781(.A1(new_n6793_), .A2(new_n6786_), .A3(new_n6702_), .ZN(new_n6794_));
  NOR2_X1    g05782(.A1(new_n6766_), .A2(new_n6765_), .ZN(new_n6795_));
  NAND2_X1   g05783(.A1(new_n6758_), .A2(new_n6760_), .ZN(new_n6796_));
  NOR2_X1    g05784(.A1(new_n6795_), .A2(new_n6796_), .ZN(new_n6797_));
  NOR2_X1    g05785(.A1(new_n6769_), .A2(new_n6768_), .ZN(new_n6798_));
  NOR3_X1    g05786(.A1(new_n6798_), .A2(new_n6765_), .A3(new_n6766_), .ZN(new_n6799_));
  INV_X1     g05787(.I(\A[183] ), .ZN(new_n6800_));
  NOR2_X1    g05788(.A1(new_n6800_), .A2(\A[182] ), .ZN(new_n6801_));
  INV_X1     g05789(.I(\A[182] ), .ZN(new_n6802_));
  NOR2_X1    g05790(.A1(new_n6802_), .A2(\A[183] ), .ZN(new_n6803_));
  OAI21_X1   g05791(.A1(new_n6801_), .A2(new_n6803_), .B(\A[181] ), .ZN(new_n6804_));
  INV_X1     g05792(.I(\A[181] ), .ZN(new_n6805_));
  NOR2_X1    g05793(.A1(\A[182] ), .A2(\A[183] ), .ZN(new_n6806_));
  NAND2_X1   g05794(.A1(\A[182] ), .A2(\A[183] ), .ZN(new_n6807_));
  INV_X1     g05795(.I(new_n6807_), .ZN(new_n6808_));
  OAI21_X1   g05796(.A1(new_n6808_), .A2(new_n6806_), .B(new_n6805_), .ZN(new_n6809_));
  NAND2_X1   g05797(.A1(new_n6804_), .A2(new_n6809_), .ZN(new_n6810_));
  INV_X1     g05798(.I(\A[186] ), .ZN(new_n6811_));
  NOR2_X1    g05799(.A1(new_n6811_), .A2(\A[185] ), .ZN(new_n6812_));
  INV_X1     g05800(.I(\A[185] ), .ZN(new_n6813_));
  NOR2_X1    g05801(.A1(new_n6813_), .A2(\A[186] ), .ZN(new_n6814_));
  OAI21_X1   g05802(.A1(new_n6812_), .A2(new_n6814_), .B(\A[184] ), .ZN(new_n6815_));
  INV_X1     g05803(.I(\A[184] ), .ZN(new_n6816_));
  NOR2_X1    g05804(.A1(\A[185] ), .A2(\A[186] ), .ZN(new_n6817_));
  AND2_X2    g05805(.A1(\A[185] ), .A2(\A[186] ), .Z(new_n6818_));
  OAI21_X1   g05806(.A1(new_n6818_), .A2(new_n6817_), .B(new_n6816_), .ZN(new_n6819_));
  NAND2_X1   g05807(.A1(new_n6815_), .A2(new_n6819_), .ZN(new_n6820_));
  NAND2_X1   g05808(.A1(\A[185] ), .A2(\A[186] ), .ZN(new_n6821_));
  AOI21_X1   g05809(.A1(new_n6816_), .A2(new_n6821_), .B(new_n6817_), .ZN(new_n6822_));
  AOI21_X1   g05810(.A1(new_n6805_), .A2(new_n6807_), .B(new_n6806_), .ZN(new_n6823_));
  NAND2_X1   g05811(.A1(new_n6822_), .A2(new_n6823_), .ZN(new_n6824_));
  NOR3_X1    g05812(.A1(new_n6810_), .A2(new_n6820_), .A3(new_n6824_), .ZN(new_n6825_));
  NOR2_X1    g05813(.A1(new_n6810_), .A2(new_n6820_), .ZN(new_n6826_));
  NAND2_X1   g05814(.A1(new_n6802_), .A2(\A[183] ), .ZN(new_n6827_));
  NAND2_X1   g05815(.A1(new_n6800_), .A2(\A[182] ), .ZN(new_n6828_));
  AOI21_X1   g05816(.A1(new_n6827_), .A2(new_n6828_), .B(new_n6805_), .ZN(new_n6829_));
  INV_X1     g05817(.I(new_n6806_), .ZN(new_n6830_));
  AOI21_X1   g05818(.A1(new_n6830_), .A2(new_n6807_), .B(\A[181] ), .ZN(new_n6831_));
  NOR2_X1    g05819(.A1(new_n6831_), .A2(new_n6829_), .ZN(new_n6832_));
  NAND2_X1   g05820(.A1(new_n6813_), .A2(\A[186] ), .ZN(new_n6833_));
  NAND2_X1   g05821(.A1(new_n6811_), .A2(\A[185] ), .ZN(new_n6834_));
  AOI21_X1   g05822(.A1(new_n6833_), .A2(new_n6834_), .B(new_n6816_), .ZN(new_n6835_));
  INV_X1     g05823(.I(new_n6817_), .ZN(new_n6836_));
  AOI21_X1   g05824(.A1(new_n6836_), .A2(new_n6821_), .B(\A[184] ), .ZN(new_n6837_));
  NOR2_X1    g05825(.A1(new_n6837_), .A2(new_n6835_), .ZN(new_n6838_));
  NOR2_X1    g05826(.A1(new_n6832_), .A2(new_n6838_), .ZN(new_n6839_));
  NOR2_X1    g05827(.A1(new_n6839_), .A2(new_n6826_), .ZN(new_n6840_));
  INV_X1     g05828(.I(\A[175] ), .ZN(new_n6841_));
  INV_X1     g05829(.I(\A[176] ), .ZN(new_n6842_));
  NAND2_X1   g05830(.A1(new_n6842_), .A2(\A[177] ), .ZN(new_n6843_));
  INV_X1     g05831(.I(\A[177] ), .ZN(new_n6844_));
  NAND2_X1   g05832(.A1(new_n6844_), .A2(\A[176] ), .ZN(new_n6845_));
  AOI21_X1   g05833(.A1(new_n6843_), .A2(new_n6845_), .B(new_n6841_), .ZN(new_n6846_));
  NOR2_X1    g05834(.A1(\A[176] ), .A2(\A[177] ), .ZN(new_n6847_));
  INV_X1     g05835(.I(new_n6847_), .ZN(new_n6848_));
  NAND2_X1   g05836(.A1(\A[176] ), .A2(\A[177] ), .ZN(new_n6849_));
  AOI21_X1   g05837(.A1(new_n6848_), .A2(new_n6849_), .B(\A[175] ), .ZN(new_n6850_));
  NOR2_X1    g05838(.A1(new_n6850_), .A2(new_n6846_), .ZN(new_n6851_));
  INV_X1     g05839(.I(\A[178] ), .ZN(new_n6852_));
  INV_X1     g05840(.I(\A[179] ), .ZN(new_n6853_));
  NAND2_X1   g05841(.A1(new_n6853_), .A2(\A[180] ), .ZN(new_n6854_));
  INV_X1     g05842(.I(\A[180] ), .ZN(new_n6855_));
  NAND2_X1   g05843(.A1(new_n6855_), .A2(\A[179] ), .ZN(new_n6856_));
  AOI21_X1   g05844(.A1(new_n6854_), .A2(new_n6856_), .B(new_n6852_), .ZN(new_n6857_));
  NOR2_X1    g05845(.A1(\A[179] ), .A2(\A[180] ), .ZN(new_n6858_));
  INV_X1     g05846(.I(new_n6858_), .ZN(new_n6859_));
  NAND2_X1   g05847(.A1(\A[179] ), .A2(\A[180] ), .ZN(new_n6860_));
  AOI21_X1   g05848(.A1(new_n6859_), .A2(new_n6860_), .B(\A[178] ), .ZN(new_n6861_));
  NOR2_X1    g05849(.A1(new_n6861_), .A2(new_n6857_), .ZN(new_n6862_));
  AOI21_X1   g05850(.A1(new_n6852_), .A2(new_n6860_), .B(new_n6858_), .ZN(new_n6863_));
  AOI21_X1   g05851(.A1(new_n6841_), .A2(new_n6849_), .B(new_n6847_), .ZN(new_n6864_));
  NAND2_X1   g05852(.A1(new_n6863_), .A2(new_n6864_), .ZN(new_n6865_));
  AND2_X2    g05853(.A1(new_n6840_), .A2(new_n6825_), .Z(new_n6867_));
  OR3_X2     g05854(.A1(new_n6797_), .A2(new_n6799_), .A3(new_n6867_), .Z(new_n6868_));
  OAI21_X1   g05855(.A1(new_n6785_), .A2(new_n6794_), .B(new_n6868_), .ZN(new_n6869_));
  NOR3_X1    g05856(.A1(new_n6797_), .A2(new_n6799_), .A3(new_n6867_), .ZN(new_n6870_));
  NAND3_X1   g05857(.A1(new_n6781_), .A2(new_n6772_), .A3(new_n6870_), .ZN(new_n6871_));
  NAND2_X1   g05858(.A1(new_n6832_), .A2(new_n6838_), .ZN(new_n6872_));
  NAND2_X1   g05859(.A1(new_n6810_), .A2(new_n6820_), .ZN(new_n6873_));
  NAND3_X1   g05860(.A1(new_n6825_), .A2(new_n6872_), .A3(new_n6873_), .ZN(new_n6874_));
  NOR4_X1    g05861(.A1(new_n6846_), .A2(new_n6850_), .A3(new_n6861_), .A4(new_n6857_), .ZN(new_n6875_));
  INV_X1     g05862(.I(new_n6875_), .ZN(new_n6876_));
  NOR2_X1    g05863(.A1(new_n6844_), .A2(\A[176] ), .ZN(new_n6877_));
  NOR2_X1    g05864(.A1(new_n6842_), .A2(\A[177] ), .ZN(new_n6878_));
  OAI21_X1   g05865(.A1(new_n6877_), .A2(new_n6878_), .B(\A[175] ), .ZN(new_n6879_));
  INV_X1     g05866(.I(new_n6849_), .ZN(new_n6880_));
  OAI21_X1   g05867(.A1(new_n6880_), .A2(new_n6847_), .B(new_n6841_), .ZN(new_n6881_));
  NAND2_X1   g05868(.A1(new_n6879_), .A2(new_n6881_), .ZN(new_n6882_));
  NOR2_X1    g05869(.A1(new_n6855_), .A2(\A[179] ), .ZN(new_n6883_));
  NOR2_X1    g05870(.A1(new_n6853_), .A2(\A[180] ), .ZN(new_n6884_));
  OAI21_X1   g05871(.A1(new_n6883_), .A2(new_n6884_), .B(\A[178] ), .ZN(new_n6885_));
  INV_X1     g05872(.I(new_n6860_), .ZN(new_n6886_));
  OAI21_X1   g05873(.A1(new_n6886_), .A2(new_n6858_), .B(new_n6852_), .ZN(new_n6887_));
  NAND2_X1   g05874(.A1(new_n6885_), .A2(new_n6887_), .ZN(new_n6888_));
  NAND2_X1   g05875(.A1(new_n6882_), .A2(new_n6888_), .ZN(new_n6889_));
  NAND2_X1   g05876(.A1(new_n6876_), .A2(new_n6889_), .ZN(new_n6890_));
  INV_X1     g05877(.I(new_n6822_), .ZN(new_n6891_));
  OAI21_X1   g05878(.A1(new_n6810_), .A2(new_n6820_), .B(new_n6823_), .ZN(new_n6892_));
  INV_X1     g05879(.I(new_n6823_), .ZN(new_n6893_));
  NAND3_X1   g05880(.A1(new_n6832_), .A2(new_n6838_), .A3(new_n6893_), .ZN(new_n6894_));
  AOI21_X1   g05881(.A1(new_n6894_), .A2(new_n6892_), .B(new_n6891_), .ZN(new_n6895_));
  AOI21_X1   g05882(.A1(new_n6832_), .A2(new_n6838_), .B(new_n6893_), .ZN(new_n6896_));
  NOR3_X1    g05883(.A1(new_n6810_), .A2(new_n6820_), .A3(new_n6823_), .ZN(new_n6897_));
  NOR3_X1    g05884(.A1(new_n6896_), .A2(new_n6897_), .A3(new_n6822_), .ZN(new_n6898_));
  NOR4_X1    g05885(.A1(new_n6895_), .A2(new_n6898_), .A3(new_n6874_), .A4(new_n6890_), .ZN(new_n6899_));
  NOR3_X1    g05886(.A1(new_n6882_), .A2(new_n6888_), .A3(new_n6865_), .ZN(new_n6900_));
  INV_X1     g05887(.I(new_n6824_), .ZN(new_n6901_));
  NOR2_X1    g05888(.A1(new_n6838_), .A2(new_n6810_), .ZN(new_n6902_));
  NOR2_X1    g05889(.A1(new_n6832_), .A2(new_n6820_), .ZN(new_n6903_));
  OAI21_X1   g05890(.A1(new_n6902_), .A2(new_n6903_), .B(new_n6901_), .ZN(new_n6904_));
  NAND2_X1   g05891(.A1(new_n6904_), .A2(new_n6900_), .ZN(new_n6905_));
  INV_X1     g05892(.I(new_n6863_), .ZN(new_n6906_));
  OAI21_X1   g05893(.A1(new_n6882_), .A2(new_n6888_), .B(new_n6864_), .ZN(new_n6907_));
  INV_X1     g05894(.I(new_n6864_), .ZN(new_n6908_));
  NAND3_X1   g05895(.A1(new_n6851_), .A2(new_n6862_), .A3(new_n6908_), .ZN(new_n6909_));
  AOI21_X1   g05896(.A1(new_n6907_), .A2(new_n6909_), .B(new_n6906_), .ZN(new_n6910_));
  NOR2_X1    g05897(.A1(new_n6875_), .A2(new_n6908_), .ZN(new_n6911_));
  NOR3_X1    g05898(.A1(new_n6882_), .A2(new_n6888_), .A3(new_n6864_), .ZN(new_n6912_));
  NOR3_X1    g05899(.A1(new_n6911_), .A2(new_n6912_), .A3(new_n6863_), .ZN(new_n6913_));
  NOR2_X1    g05900(.A1(new_n6913_), .A2(new_n6910_), .ZN(new_n6914_));
  NOR3_X1    g05901(.A1(new_n6899_), .A2(new_n6905_), .A3(new_n6914_), .ZN(new_n6915_));
  INV_X1     g05902(.I(new_n6915_), .ZN(new_n6916_));
  OAI21_X1   g05903(.A1(new_n6911_), .A2(new_n6912_), .B(new_n6863_), .ZN(new_n6917_));
  NAND3_X1   g05904(.A1(new_n6907_), .A2(new_n6909_), .A3(new_n6906_), .ZN(new_n6918_));
  NAND2_X1   g05905(.A1(new_n6917_), .A2(new_n6918_), .ZN(new_n6919_));
  NOR2_X1    g05906(.A1(new_n6851_), .A2(new_n6862_), .ZN(new_n6920_));
  NOR2_X1    g05907(.A1(new_n6920_), .A2(new_n6875_), .ZN(new_n6921_));
  NAND4_X1   g05908(.A1(new_n6840_), .A2(new_n6921_), .A3(new_n6825_), .A4(new_n6900_), .ZN(new_n6922_));
  NAND2_X1   g05909(.A1(new_n6919_), .A2(new_n6922_), .ZN(new_n6923_));
  NAND2_X1   g05910(.A1(new_n6832_), .A2(new_n6820_), .ZN(new_n6924_));
  NAND2_X1   g05911(.A1(new_n6838_), .A2(new_n6810_), .ZN(new_n6925_));
  AOI21_X1   g05912(.A1(new_n6925_), .A2(new_n6924_), .B(new_n6824_), .ZN(new_n6926_));
  NOR3_X1    g05913(.A1(new_n6898_), .A2(new_n6895_), .A3(new_n6926_), .ZN(new_n6927_));
  NAND3_X1   g05914(.A1(new_n6876_), .A2(new_n6900_), .A3(new_n6889_), .ZN(new_n6928_));
  NOR4_X1    g05915(.A1(new_n6913_), .A2(new_n6910_), .A3(new_n6928_), .A4(new_n6874_), .ZN(new_n6929_));
  NOR2_X1    g05916(.A1(new_n6929_), .A2(new_n6927_), .ZN(new_n6930_));
  OAI21_X1   g05917(.A1(new_n6896_), .A2(new_n6897_), .B(new_n6822_), .ZN(new_n6931_));
  NAND3_X1   g05918(.A1(new_n6894_), .A2(new_n6892_), .A3(new_n6891_), .ZN(new_n6932_));
  NAND3_X1   g05919(.A1(new_n6931_), .A2(new_n6932_), .A3(new_n6904_), .ZN(new_n6933_));
  NOR3_X1    g05920(.A1(new_n6933_), .A2(new_n6919_), .A3(new_n6922_), .ZN(new_n6934_));
  OAI21_X1   g05921(.A1(new_n6930_), .A2(new_n6934_), .B(new_n6923_), .ZN(new_n6935_));
  NAND2_X1   g05922(.A1(new_n6935_), .A2(new_n6916_), .ZN(new_n6936_));
  AOI22_X1   g05923(.A1(new_n6869_), .A2(new_n6871_), .B1(new_n6936_), .B2(new_n6782_), .ZN(new_n6937_));
  OAI21_X1   g05924(.A1(new_n6763_), .A2(new_n6761_), .B(new_n6702_), .ZN(new_n6938_));
  NAND2_X1   g05925(.A1(new_n6744_), .A2(new_n6747_), .ZN(new_n6939_));
  AOI21_X1   g05926(.A1(new_n6754_), .A2(new_n6939_), .B(new_n6764_), .ZN(new_n6940_));
  NOR2_X1    g05927(.A1(new_n6662_), .A2(new_n6666_), .ZN(new_n6941_));
  OAI21_X1   g05928(.A1(new_n6694_), .A2(new_n6941_), .B(new_n6759_), .ZN(new_n6942_));
  XOR2_X1    g05929(.A1(new_n6940_), .A2(new_n6942_), .Z(new_n6943_));
  NAND3_X1   g05930(.A1(new_n6938_), .A2(new_n6780_), .A3(new_n6943_), .ZN(new_n6944_));
  NOR2_X1    g05931(.A1(new_n6874_), .A2(new_n6890_), .ZN(new_n6945_));
  NAND3_X1   g05932(.A1(new_n6945_), .A2(new_n6931_), .A3(new_n6932_), .ZN(new_n6946_));
  INV_X1     g05933(.I(new_n6905_), .ZN(new_n6947_));
  NAND2_X1   g05934(.A1(new_n6946_), .A2(new_n6947_), .ZN(new_n6948_));
  OAI21_X1   g05935(.A1(new_n6927_), .A2(new_n6922_), .B(new_n6919_), .ZN(new_n6949_));
  NOR2_X1    g05936(.A1(new_n6822_), .A2(new_n6823_), .ZN(new_n6950_));
  OAI21_X1   g05937(.A1(new_n6872_), .A2(new_n6950_), .B(new_n6824_), .ZN(new_n6951_));
  NOR2_X1    g05938(.A1(new_n6863_), .A2(new_n6864_), .ZN(new_n6952_));
  OAI21_X1   g05939(.A1(new_n6876_), .A2(new_n6952_), .B(new_n6865_), .ZN(new_n6953_));
  XNOR2_X1   g05940(.A1(new_n6953_), .A2(new_n6951_), .ZN(new_n6954_));
  NAND3_X1   g05941(.A1(new_n6948_), .A2(new_n6949_), .A3(new_n6954_), .ZN(new_n6955_));
  XOR2_X1    g05942(.A1(new_n6955_), .A2(new_n6944_), .Z(new_n6956_));
  NAND2_X1   g05943(.A1(new_n6956_), .A2(new_n6937_), .ZN(new_n6957_));
  NAND3_X1   g05944(.A1(new_n6781_), .A2(new_n6772_), .A3(new_n6870_), .ZN(new_n6958_));
  AOI21_X1   g05945(.A1(new_n6781_), .A2(new_n6772_), .B(new_n6870_), .ZN(new_n6959_));
  NOR3_X1    g05946(.A1(new_n6785_), .A2(new_n6794_), .A3(new_n6868_), .ZN(new_n6960_));
  OAI21_X1   g05947(.A1(new_n6919_), .A2(new_n6922_), .B(new_n6933_), .ZN(new_n6961_));
  NAND2_X1   g05948(.A1(new_n6929_), .A2(new_n6927_), .ZN(new_n6962_));
  NAND2_X1   g05949(.A1(new_n6961_), .A2(new_n6962_), .ZN(new_n6963_));
  AOI21_X1   g05950(.A1(new_n6963_), .A2(new_n6923_), .B(new_n6915_), .ZN(new_n6964_));
  OAI21_X1   g05951(.A1(new_n6960_), .A2(new_n6959_), .B(new_n6964_), .ZN(new_n6965_));
  NAND2_X1   g05952(.A1(new_n6955_), .A2(new_n6944_), .ZN(new_n6966_));
  INV_X1     g05953(.I(new_n6944_), .ZN(new_n6967_));
  NOR2_X1    g05954(.A1(new_n6899_), .A2(new_n6905_), .ZN(new_n6968_));
  INV_X1     g05955(.I(new_n6922_), .ZN(new_n6969_));
  AOI21_X1   g05956(.A1(new_n6969_), .A2(new_n6933_), .B(new_n6914_), .ZN(new_n6970_));
  XOR2_X1    g05957(.A1(new_n6953_), .A2(new_n6951_), .Z(new_n6971_));
  NOR3_X1    g05958(.A1(new_n6970_), .A2(new_n6968_), .A3(new_n6971_), .ZN(new_n6972_));
  NAND2_X1   g05959(.A1(new_n6967_), .A2(new_n6972_), .ZN(new_n6973_));
  NAND2_X1   g05960(.A1(new_n6973_), .A2(new_n6966_), .ZN(new_n6974_));
  NAND3_X1   g05961(.A1(new_n6974_), .A2(new_n6965_), .A3(new_n6958_), .ZN(new_n6975_));
  AND2_X2    g05962(.A1(new_n6975_), .A2(new_n6957_), .Z(new_n6976_));
  INV_X1     g05963(.I(\A[220] ), .ZN(new_n6977_));
  NOR2_X1    g05964(.A1(\A[221] ), .A2(\A[222] ), .ZN(new_n6978_));
  NAND2_X1   g05965(.A1(\A[221] ), .A2(\A[222] ), .ZN(new_n6979_));
  AOI21_X1   g05966(.A1(new_n6977_), .A2(new_n6979_), .B(new_n6978_), .ZN(new_n6980_));
  INV_X1     g05967(.I(new_n6980_), .ZN(new_n6981_));
  INV_X1     g05968(.I(\A[217] ), .ZN(new_n6982_));
  NOR2_X1    g05969(.A1(\A[218] ), .A2(\A[219] ), .ZN(new_n6983_));
  NAND2_X1   g05970(.A1(\A[218] ), .A2(\A[219] ), .ZN(new_n6984_));
  AOI21_X1   g05971(.A1(new_n6982_), .A2(new_n6984_), .B(new_n6983_), .ZN(new_n6985_));
  INV_X1     g05972(.I(\A[219] ), .ZN(new_n6986_));
  NOR2_X1    g05973(.A1(new_n6986_), .A2(\A[218] ), .ZN(new_n6987_));
  INV_X1     g05974(.I(\A[218] ), .ZN(new_n6988_));
  NOR2_X1    g05975(.A1(new_n6988_), .A2(\A[219] ), .ZN(new_n6989_));
  OAI21_X1   g05976(.A1(new_n6987_), .A2(new_n6989_), .B(\A[217] ), .ZN(new_n6990_));
  INV_X1     g05977(.I(new_n6984_), .ZN(new_n6991_));
  OAI21_X1   g05978(.A1(new_n6991_), .A2(new_n6983_), .B(new_n6982_), .ZN(new_n6992_));
  INV_X1     g05979(.I(\A[222] ), .ZN(new_n6993_));
  NOR2_X1    g05980(.A1(new_n6993_), .A2(\A[221] ), .ZN(new_n6994_));
  INV_X1     g05981(.I(\A[221] ), .ZN(new_n6995_));
  NOR2_X1    g05982(.A1(new_n6995_), .A2(\A[222] ), .ZN(new_n6996_));
  OAI21_X1   g05983(.A1(new_n6994_), .A2(new_n6996_), .B(\A[220] ), .ZN(new_n6997_));
  INV_X1     g05984(.I(new_n6979_), .ZN(new_n6998_));
  OAI21_X1   g05985(.A1(new_n6998_), .A2(new_n6978_), .B(new_n6977_), .ZN(new_n6999_));
  NAND4_X1   g05986(.A1(new_n6990_), .A2(new_n6992_), .A3(new_n6997_), .A4(new_n6999_), .ZN(new_n7000_));
  NAND2_X1   g05987(.A1(new_n7000_), .A2(new_n6985_), .ZN(new_n7001_));
  INV_X1     g05988(.I(new_n6985_), .ZN(new_n7002_));
  NAND2_X1   g05989(.A1(new_n6988_), .A2(\A[219] ), .ZN(new_n7003_));
  NAND2_X1   g05990(.A1(new_n6986_), .A2(\A[218] ), .ZN(new_n7004_));
  AOI21_X1   g05991(.A1(new_n7003_), .A2(new_n7004_), .B(new_n6982_), .ZN(new_n7005_));
  INV_X1     g05992(.I(new_n6983_), .ZN(new_n7006_));
  AOI21_X1   g05993(.A1(new_n7006_), .A2(new_n6984_), .B(\A[217] ), .ZN(new_n7007_));
  NAND2_X1   g05994(.A1(new_n6995_), .A2(\A[222] ), .ZN(new_n7008_));
  NAND2_X1   g05995(.A1(new_n6993_), .A2(\A[221] ), .ZN(new_n7009_));
  AOI21_X1   g05996(.A1(new_n7008_), .A2(new_n7009_), .B(new_n6977_), .ZN(new_n7010_));
  INV_X1     g05997(.I(new_n6978_), .ZN(new_n7011_));
  AOI21_X1   g05998(.A1(new_n7011_), .A2(new_n6979_), .B(\A[220] ), .ZN(new_n7012_));
  NOR4_X1    g05999(.A1(new_n7005_), .A2(new_n7007_), .A3(new_n7012_), .A4(new_n7010_), .ZN(new_n7013_));
  NAND2_X1   g06000(.A1(new_n7013_), .A2(new_n7002_), .ZN(new_n7014_));
  AOI21_X1   g06001(.A1(new_n7014_), .A2(new_n7001_), .B(new_n6981_), .ZN(new_n7015_));
  NOR2_X1    g06002(.A1(new_n7013_), .A2(new_n7002_), .ZN(new_n7016_));
  NOR2_X1    g06003(.A1(new_n7000_), .A2(new_n6985_), .ZN(new_n7017_));
  NOR3_X1    g06004(.A1(new_n7016_), .A2(new_n7017_), .A3(new_n6980_), .ZN(new_n7018_));
  INV_X1     g06005(.I(\A[213] ), .ZN(new_n7019_));
  NOR2_X1    g06006(.A1(new_n7019_), .A2(\A[212] ), .ZN(new_n7020_));
  INV_X1     g06007(.I(\A[212] ), .ZN(new_n7021_));
  NOR2_X1    g06008(.A1(new_n7021_), .A2(\A[213] ), .ZN(new_n7022_));
  OAI21_X1   g06009(.A1(new_n7020_), .A2(new_n7022_), .B(\A[211] ), .ZN(new_n7023_));
  INV_X1     g06010(.I(\A[211] ), .ZN(new_n7024_));
  NOR2_X1    g06011(.A1(\A[212] ), .A2(\A[213] ), .ZN(new_n7025_));
  NAND2_X1   g06012(.A1(\A[212] ), .A2(\A[213] ), .ZN(new_n7026_));
  INV_X1     g06013(.I(new_n7026_), .ZN(new_n7027_));
  OAI21_X1   g06014(.A1(new_n7027_), .A2(new_n7025_), .B(new_n7024_), .ZN(new_n7028_));
  INV_X1     g06015(.I(\A[216] ), .ZN(new_n7029_));
  NOR2_X1    g06016(.A1(new_n7029_), .A2(\A[215] ), .ZN(new_n7030_));
  INV_X1     g06017(.I(\A[215] ), .ZN(new_n7031_));
  NOR2_X1    g06018(.A1(new_n7031_), .A2(\A[216] ), .ZN(new_n7032_));
  OAI21_X1   g06019(.A1(new_n7030_), .A2(new_n7032_), .B(\A[214] ), .ZN(new_n7033_));
  INV_X1     g06020(.I(\A[214] ), .ZN(new_n7034_));
  NOR2_X1    g06021(.A1(\A[215] ), .A2(\A[216] ), .ZN(new_n7035_));
  NAND2_X1   g06022(.A1(\A[215] ), .A2(\A[216] ), .ZN(new_n7036_));
  INV_X1     g06023(.I(new_n7036_), .ZN(new_n7037_));
  OAI21_X1   g06024(.A1(new_n7037_), .A2(new_n7035_), .B(new_n7034_), .ZN(new_n7038_));
  NAND4_X1   g06025(.A1(new_n7023_), .A2(new_n7028_), .A3(new_n7033_), .A4(new_n7038_), .ZN(new_n7039_));
  NAND2_X1   g06026(.A1(new_n7021_), .A2(\A[213] ), .ZN(new_n7040_));
  NAND2_X1   g06027(.A1(new_n7019_), .A2(\A[212] ), .ZN(new_n7041_));
  AOI21_X1   g06028(.A1(new_n7040_), .A2(new_n7041_), .B(new_n7024_), .ZN(new_n7042_));
  INV_X1     g06029(.I(new_n7025_), .ZN(new_n7043_));
  AOI21_X1   g06030(.A1(new_n7043_), .A2(new_n7026_), .B(\A[211] ), .ZN(new_n7044_));
  NAND2_X1   g06031(.A1(new_n7031_), .A2(\A[216] ), .ZN(new_n7045_));
  NAND2_X1   g06032(.A1(new_n7029_), .A2(\A[215] ), .ZN(new_n7046_));
  AOI21_X1   g06033(.A1(new_n7045_), .A2(new_n7046_), .B(new_n7034_), .ZN(new_n7047_));
  INV_X1     g06034(.I(new_n7035_), .ZN(new_n7048_));
  AOI21_X1   g06035(.A1(new_n7048_), .A2(new_n7036_), .B(\A[214] ), .ZN(new_n7049_));
  OAI22_X1   g06036(.A1(new_n7042_), .A2(new_n7044_), .B1(new_n7049_), .B2(new_n7047_), .ZN(new_n7050_));
  NAND2_X1   g06037(.A1(new_n7050_), .A2(new_n7039_), .ZN(new_n7051_));
  OAI22_X1   g06038(.A1(new_n7005_), .A2(new_n7007_), .B1(new_n7012_), .B2(new_n7010_), .ZN(new_n7052_));
  NAND2_X1   g06039(.A1(new_n7052_), .A2(new_n7000_), .ZN(new_n7053_));
  NAND2_X1   g06040(.A1(new_n6980_), .A2(new_n6985_), .ZN(new_n7054_));
  NOR2_X1    g06041(.A1(new_n7000_), .A2(new_n7054_), .ZN(new_n7055_));
  NOR4_X1    g06042(.A1(new_n7042_), .A2(new_n7044_), .A3(new_n7049_), .A4(new_n7047_), .ZN(new_n7056_));
  AOI21_X1   g06043(.A1(new_n7034_), .A2(new_n7036_), .B(new_n7035_), .ZN(new_n7057_));
  AOI21_X1   g06044(.A1(new_n7024_), .A2(new_n7026_), .B(new_n7025_), .ZN(new_n7058_));
  NAND3_X1   g06045(.A1(new_n7056_), .A2(new_n7057_), .A3(new_n7058_), .ZN(new_n7059_));
  NOR4_X1    g06046(.A1(new_n7051_), .A2(new_n7059_), .A3(new_n7053_), .A4(new_n7055_), .ZN(new_n7060_));
  NOR3_X1    g06047(.A1(new_n7060_), .A2(new_n7015_), .A3(new_n7018_), .ZN(new_n7061_));
  INV_X1     g06048(.I(new_n7058_), .ZN(new_n7062_));
  NOR2_X1    g06049(.A1(new_n7056_), .A2(new_n7062_), .ZN(new_n7063_));
  NOR2_X1    g06050(.A1(new_n7039_), .A2(new_n7058_), .ZN(new_n7064_));
  OAI21_X1   g06051(.A1(new_n7063_), .A2(new_n7064_), .B(new_n7057_), .ZN(new_n7065_));
  INV_X1     g06052(.I(new_n7057_), .ZN(new_n7066_));
  NAND2_X1   g06053(.A1(new_n7039_), .A2(new_n7058_), .ZN(new_n7067_));
  NAND2_X1   g06054(.A1(new_n7056_), .A2(new_n7062_), .ZN(new_n7068_));
  NAND3_X1   g06055(.A1(new_n7068_), .A2(new_n7067_), .A3(new_n7066_), .ZN(new_n7069_));
  NAND2_X1   g06056(.A1(new_n7065_), .A2(new_n7069_), .ZN(new_n7070_));
  NAND4_X1   g06057(.A1(new_n7000_), .A2(new_n7050_), .A3(new_n7052_), .A4(new_n7039_), .ZN(new_n7071_));
  AOI22_X1   g06058(.A1(new_n6990_), .A2(new_n6992_), .B1(new_n6997_), .B2(new_n6999_), .ZN(new_n7072_));
  NAND2_X1   g06059(.A1(new_n7057_), .A2(new_n7058_), .ZN(new_n7073_));
  NOR2_X1    g06060(.A1(new_n7039_), .A2(new_n7073_), .ZN(new_n7074_));
  OAI21_X1   g06061(.A1(new_n7072_), .A2(new_n7054_), .B(new_n7074_), .ZN(new_n7075_));
  XOR2_X1    g06062(.A1(new_n6980_), .A2(new_n6985_), .Z(new_n7076_));
  NAND2_X1   g06063(.A1(new_n7076_), .A2(new_n7013_), .ZN(new_n7077_));
  NAND2_X1   g06064(.A1(new_n6981_), .A2(new_n7002_), .ZN(new_n7078_));
  NAND2_X1   g06065(.A1(new_n7078_), .A2(new_n7054_), .ZN(new_n7079_));
  NAND2_X1   g06066(.A1(new_n7079_), .A2(new_n7000_), .ZN(new_n7080_));
  NAND2_X1   g06067(.A1(new_n7080_), .A2(new_n7077_), .ZN(new_n7081_));
  NOR3_X1    g06068(.A1(new_n7081_), .A2(new_n7075_), .A3(new_n7071_), .ZN(new_n7082_));
  NOR3_X1    g06069(.A1(new_n7061_), .A2(new_n7082_), .A3(new_n7070_), .ZN(new_n7083_));
  INV_X1     g06070(.I(new_n7054_), .ZN(new_n7084_));
  NAND2_X1   g06071(.A1(new_n7013_), .A2(new_n7084_), .ZN(new_n7085_));
  NAND2_X1   g06072(.A1(new_n7085_), .A2(new_n7074_), .ZN(new_n7086_));
  OAI22_X1   g06073(.A1(new_n7015_), .A2(new_n7018_), .B1(new_n7086_), .B2(new_n7071_), .ZN(new_n7087_));
  OAI21_X1   g06074(.A1(new_n7016_), .A2(new_n7017_), .B(new_n6980_), .ZN(new_n7088_));
  NAND3_X1   g06075(.A1(new_n7014_), .A2(new_n7001_), .A3(new_n6981_), .ZN(new_n7089_));
  AOI22_X1   g06076(.A1(new_n7023_), .A2(new_n7028_), .B1(new_n7033_), .B2(new_n7038_), .ZN(new_n7090_));
  NOR4_X1    g06077(.A1(new_n7013_), .A2(new_n7090_), .A3(new_n7072_), .A4(new_n7056_), .ZN(new_n7091_));
  NOR2_X1    g06078(.A1(new_n7059_), .A2(new_n7055_), .ZN(new_n7092_));
  NAND4_X1   g06079(.A1(new_n7088_), .A2(new_n7089_), .A3(new_n7092_), .A4(new_n7091_), .ZN(new_n7093_));
  AOI21_X1   g06080(.A1(new_n7087_), .A2(new_n7093_), .B(new_n7070_), .ZN(new_n7094_));
  NOR2_X1    g06081(.A1(new_n7083_), .A2(new_n7094_), .ZN(new_n7095_));
  NOR2_X1    g06082(.A1(new_n7090_), .A2(new_n7056_), .ZN(new_n7096_));
  NOR2_X1    g06083(.A1(new_n7072_), .A2(new_n7013_), .ZN(new_n7097_));
  NAND4_X1   g06084(.A1(new_n7096_), .A2(new_n7097_), .A3(new_n7085_), .A4(new_n7074_), .ZN(new_n7098_));
  NAND3_X1   g06085(.A1(new_n7098_), .A2(new_n7088_), .A3(new_n7089_), .ZN(new_n7099_));
  AOI21_X1   g06086(.A1(new_n7068_), .A2(new_n7067_), .B(new_n7066_), .ZN(new_n7100_));
  NOR3_X1    g06087(.A1(new_n7063_), .A2(new_n7064_), .A3(new_n7057_), .ZN(new_n7101_));
  NOR2_X1    g06088(.A1(new_n7100_), .A2(new_n7101_), .ZN(new_n7102_));
  NOR2_X1    g06089(.A1(new_n7072_), .A2(new_n7054_), .ZN(new_n7103_));
  NOR2_X1    g06090(.A1(new_n7059_), .A2(new_n7103_), .ZN(new_n7104_));
  NAND4_X1   g06091(.A1(new_n7104_), .A2(new_n7091_), .A3(new_n7077_), .A4(new_n7080_), .ZN(new_n7105_));
  NAND3_X1   g06092(.A1(new_n7099_), .A2(new_n7102_), .A3(new_n7105_), .ZN(new_n7106_));
  AOI22_X1   g06093(.A1(new_n7088_), .A2(new_n7089_), .B1(new_n7092_), .B2(new_n7091_), .ZN(new_n7107_));
  NOR3_X1    g06094(.A1(new_n7098_), .A2(new_n7015_), .A3(new_n7018_), .ZN(new_n7108_));
  OAI21_X1   g06095(.A1(new_n7108_), .A2(new_n7107_), .B(new_n7102_), .ZN(new_n7109_));
  NOR2_X1    g06096(.A1(new_n7072_), .A2(new_n7013_), .ZN(new_n7110_));
  INV_X1     g06097(.I(new_n7110_), .ZN(new_n7111_));
  NAND2_X1   g06098(.A1(new_n7096_), .A2(new_n7074_), .ZN(new_n7112_));
  INV_X1     g06099(.I(new_n7112_), .ZN(new_n7113_));
  NAND2_X1   g06100(.A1(new_n7113_), .A2(new_n7111_), .ZN(new_n7114_));
  NAND2_X1   g06101(.A1(new_n7112_), .A2(new_n7110_), .ZN(new_n7115_));
  INV_X1     g06102(.I(\A[208] ), .ZN(new_n7116_));
  NOR2_X1    g06103(.A1(\A[209] ), .A2(\A[210] ), .ZN(new_n7117_));
  NAND2_X1   g06104(.A1(\A[209] ), .A2(\A[210] ), .ZN(new_n7118_));
  AOI21_X1   g06105(.A1(new_n7116_), .A2(new_n7118_), .B(new_n7117_), .ZN(new_n7119_));
  INV_X1     g06106(.I(\A[205] ), .ZN(new_n7120_));
  NOR2_X1    g06107(.A1(\A[206] ), .A2(\A[207] ), .ZN(new_n7121_));
  NAND2_X1   g06108(.A1(\A[206] ), .A2(\A[207] ), .ZN(new_n7122_));
  AOI21_X1   g06109(.A1(new_n7120_), .A2(new_n7122_), .B(new_n7121_), .ZN(new_n7123_));
  NAND2_X1   g06110(.A1(new_n7119_), .A2(new_n7123_), .ZN(new_n7124_));
  INV_X1     g06111(.I(new_n7124_), .ZN(new_n7125_));
  INV_X1     g06112(.I(\A[207] ), .ZN(new_n7126_));
  NOR2_X1    g06113(.A1(new_n7126_), .A2(\A[206] ), .ZN(new_n7127_));
  INV_X1     g06114(.I(\A[206] ), .ZN(new_n7128_));
  NOR2_X1    g06115(.A1(new_n7128_), .A2(\A[207] ), .ZN(new_n7129_));
  OAI21_X1   g06116(.A1(new_n7127_), .A2(new_n7129_), .B(\A[205] ), .ZN(new_n7130_));
  INV_X1     g06117(.I(new_n7122_), .ZN(new_n7131_));
  OAI21_X1   g06118(.A1(new_n7131_), .A2(new_n7121_), .B(new_n7120_), .ZN(new_n7132_));
  NAND2_X1   g06119(.A1(new_n7130_), .A2(new_n7132_), .ZN(new_n7133_));
  INV_X1     g06120(.I(\A[210] ), .ZN(new_n7134_));
  NOR2_X1    g06121(.A1(new_n7134_), .A2(\A[209] ), .ZN(new_n7135_));
  INV_X1     g06122(.I(\A[209] ), .ZN(new_n7136_));
  NOR2_X1    g06123(.A1(new_n7136_), .A2(\A[210] ), .ZN(new_n7137_));
  OAI21_X1   g06124(.A1(new_n7135_), .A2(new_n7137_), .B(\A[208] ), .ZN(new_n7138_));
  AND2_X2    g06125(.A1(\A[209] ), .A2(\A[210] ), .Z(new_n7139_));
  OAI21_X1   g06126(.A1(new_n7139_), .A2(new_n7117_), .B(new_n7116_), .ZN(new_n7140_));
  NAND2_X1   g06127(.A1(new_n7138_), .A2(new_n7140_), .ZN(new_n7141_));
  NOR2_X1    g06128(.A1(new_n7133_), .A2(new_n7141_), .ZN(new_n7142_));
  NAND2_X1   g06129(.A1(new_n7142_), .A2(new_n7125_), .ZN(new_n7143_));
  NAND2_X1   g06130(.A1(new_n7128_), .A2(\A[207] ), .ZN(new_n7144_));
  NAND2_X1   g06131(.A1(new_n7126_), .A2(\A[206] ), .ZN(new_n7145_));
  AOI21_X1   g06132(.A1(new_n7144_), .A2(new_n7145_), .B(new_n7120_), .ZN(new_n7146_));
  INV_X1     g06133(.I(new_n7121_), .ZN(new_n7147_));
  AOI21_X1   g06134(.A1(new_n7147_), .A2(new_n7122_), .B(\A[205] ), .ZN(new_n7148_));
  NOR2_X1    g06135(.A1(new_n7148_), .A2(new_n7146_), .ZN(new_n7149_));
  NAND2_X1   g06136(.A1(new_n7136_), .A2(\A[210] ), .ZN(new_n7150_));
  NAND2_X1   g06137(.A1(new_n7134_), .A2(\A[209] ), .ZN(new_n7151_));
  AOI21_X1   g06138(.A1(new_n7150_), .A2(new_n7151_), .B(new_n7116_), .ZN(new_n7152_));
  INV_X1     g06139(.I(new_n7117_), .ZN(new_n7153_));
  AOI21_X1   g06140(.A1(new_n7153_), .A2(new_n7118_), .B(\A[208] ), .ZN(new_n7154_));
  NOR2_X1    g06141(.A1(new_n7154_), .A2(new_n7152_), .ZN(new_n7155_));
  NOR2_X1    g06142(.A1(new_n7149_), .A2(new_n7155_), .ZN(new_n7156_));
  NOR2_X1    g06143(.A1(new_n7156_), .A2(new_n7142_), .ZN(new_n7157_));
  INV_X1     g06144(.I(\A[199] ), .ZN(new_n7158_));
  INV_X1     g06145(.I(\A[200] ), .ZN(new_n7159_));
  NAND2_X1   g06146(.A1(new_n7159_), .A2(\A[201] ), .ZN(new_n7160_));
  INV_X1     g06147(.I(\A[201] ), .ZN(new_n7161_));
  NAND2_X1   g06148(.A1(new_n7161_), .A2(\A[200] ), .ZN(new_n7162_));
  AOI21_X1   g06149(.A1(new_n7160_), .A2(new_n7162_), .B(new_n7158_), .ZN(new_n7163_));
  NOR2_X1    g06150(.A1(\A[200] ), .A2(\A[201] ), .ZN(new_n7164_));
  INV_X1     g06151(.I(new_n7164_), .ZN(new_n7165_));
  NAND2_X1   g06152(.A1(\A[200] ), .A2(\A[201] ), .ZN(new_n7166_));
  AOI21_X1   g06153(.A1(new_n7165_), .A2(new_n7166_), .B(\A[199] ), .ZN(new_n7167_));
  NOR2_X1    g06154(.A1(new_n7167_), .A2(new_n7163_), .ZN(new_n7168_));
  INV_X1     g06155(.I(\A[202] ), .ZN(new_n7169_));
  INV_X1     g06156(.I(\A[203] ), .ZN(new_n7170_));
  NAND2_X1   g06157(.A1(new_n7170_), .A2(\A[204] ), .ZN(new_n7171_));
  INV_X1     g06158(.I(\A[204] ), .ZN(new_n7172_));
  NAND2_X1   g06159(.A1(new_n7172_), .A2(\A[203] ), .ZN(new_n7173_));
  AOI21_X1   g06160(.A1(new_n7171_), .A2(new_n7173_), .B(new_n7169_), .ZN(new_n7174_));
  NOR2_X1    g06161(.A1(\A[203] ), .A2(\A[204] ), .ZN(new_n7175_));
  INV_X1     g06162(.I(new_n7175_), .ZN(new_n7176_));
  NAND2_X1   g06163(.A1(\A[203] ), .A2(\A[204] ), .ZN(new_n7177_));
  AOI21_X1   g06164(.A1(new_n7176_), .A2(new_n7177_), .B(\A[202] ), .ZN(new_n7178_));
  NOR2_X1    g06165(.A1(new_n7178_), .A2(new_n7174_), .ZN(new_n7179_));
  AOI21_X1   g06166(.A1(new_n7169_), .A2(new_n7177_), .B(new_n7175_), .ZN(new_n7180_));
  AOI21_X1   g06167(.A1(new_n7158_), .A2(new_n7166_), .B(new_n7164_), .ZN(new_n7181_));
  NAND2_X1   g06168(.A1(new_n7180_), .A2(new_n7181_), .ZN(new_n7182_));
  INV_X1     g06169(.I(new_n7182_), .ZN(new_n7183_));
  NAND2_X1   g06170(.A1(new_n7157_), .A2(new_n7143_), .ZN(new_n7184_));
  AOI21_X1   g06171(.A1(new_n7114_), .A2(new_n7115_), .B(new_n7184_), .ZN(new_n7185_));
  AOI21_X1   g06172(.A1(new_n7109_), .A2(new_n7106_), .B(new_n7185_), .ZN(new_n7186_));
  NOR2_X1    g06173(.A1(new_n7112_), .A2(new_n7110_), .ZN(new_n7187_));
  AOI21_X1   g06174(.A1(new_n7096_), .A2(new_n7074_), .B(new_n7111_), .ZN(new_n7188_));
  INV_X1     g06175(.I(new_n7184_), .ZN(new_n7189_));
  OAI21_X1   g06176(.A1(new_n7188_), .A2(new_n7187_), .B(new_n7189_), .ZN(new_n7190_));
  NOR3_X1    g06177(.A1(new_n7083_), .A2(new_n7094_), .A3(new_n7190_), .ZN(new_n7191_));
  INV_X1     g06178(.I(new_n7180_), .ZN(new_n7192_));
  NOR2_X1    g06179(.A1(new_n7161_), .A2(\A[200] ), .ZN(new_n7193_));
  NOR2_X1    g06180(.A1(new_n7159_), .A2(\A[201] ), .ZN(new_n7194_));
  OAI21_X1   g06181(.A1(new_n7193_), .A2(new_n7194_), .B(\A[199] ), .ZN(new_n7195_));
  INV_X1     g06182(.I(new_n7166_), .ZN(new_n7196_));
  OAI21_X1   g06183(.A1(new_n7196_), .A2(new_n7164_), .B(new_n7158_), .ZN(new_n7197_));
  NOR2_X1    g06184(.A1(new_n7172_), .A2(\A[203] ), .ZN(new_n7198_));
  NOR2_X1    g06185(.A1(new_n7170_), .A2(\A[204] ), .ZN(new_n7199_));
  OAI21_X1   g06186(.A1(new_n7198_), .A2(new_n7199_), .B(\A[202] ), .ZN(new_n7200_));
  INV_X1     g06187(.I(new_n7177_), .ZN(new_n7201_));
  OAI21_X1   g06188(.A1(new_n7201_), .A2(new_n7175_), .B(new_n7169_), .ZN(new_n7202_));
  NAND4_X1   g06189(.A1(new_n7195_), .A2(new_n7197_), .A3(new_n7200_), .A4(new_n7202_), .ZN(new_n7203_));
  NAND2_X1   g06190(.A1(new_n7203_), .A2(new_n7181_), .ZN(new_n7204_));
  INV_X1     g06191(.I(new_n7181_), .ZN(new_n7205_));
  NAND3_X1   g06192(.A1(new_n7168_), .A2(new_n7179_), .A3(new_n7205_), .ZN(new_n7206_));
  AOI21_X1   g06193(.A1(new_n7204_), .A2(new_n7206_), .B(new_n7192_), .ZN(new_n7207_));
  NOR4_X1    g06194(.A1(new_n7163_), .A2(new_n7167_), .A3(new_n7178_), .A4(new_n7174_), .ZN(new_n7208_));
  NOR2_X1    g06195(.A1(new_n7208_), .A2(new_n7205_), .ZN(new_n7209_));
  NOR2_X1    g06196(.A1(new_n7203_), .A2(new_n7181_), .ZN(new_n7210_));
  NOR3_X1    g06197(.A1(new_n7209_), .A2(new_n7210_), .A3(new_n7180_), .ZN(new_n7211_));
  NOR2_X1    g06198(.A1(new_n7211_), .A2(new_n7207_), .ZN(new_n7212_));
  NOR2_X1    g06199(.A1(new_n7168_), .A2(new_n7179_), .ZN(new_n7213_));
  NOR2_X1    g06200(.A1(new_n7213_), .A2(new_n7208_), .ZN(new_n7214_));
  NAND2_X1   g06201(.A1(new_n7133_), .A2(new_n7141_), .ZN(new_n7215_));
  NAND2_X1   g06202(.A1(new_n7208_), .A2(new_n7183_), .ZN(new_n7216_));
  AOI21_X1   g06203(.A1(new_n7125_), .A2(new_n7215_), .B(new_n7216_), .ZN(new_n7217_));
  NAND4_X1   g06204(.A1(new_n7130_), .A2(new_n7138_), .A3(new_n7132_), .A4(new_n7140_), .ZN(new_n7218_));
  XNOR2_X1   g06205(.A1(new_n7119_), .A2(new_n7123_), .ZN(new_n7219_));
  NOR2_X1    g06206(.A1(new_n7219_), .A2(new_n7218_), .ZN(new_n7220_));
  INV_X1     g06207(.I(new_n7119_), .ZN(new_n7221_));
  INV_X1     g06208(.I(new_n7123_), .ZN(new_n7222_));
  NAND2_X1   g06209(.A1(new_n7222_), .A2(new_n7221_), .ZN(new_n7223_));
  AOI21_X1   g06210(.A1(new_n7124_), .A2(new_n7223_), .B(new_n7142_), .ZN(new_n7224_));
  NOR2_X1    g06211(.A1(new_n7224_), .A2(new_n7220_), .ZN(new_n7225_));
  NAND4_X1   g06212(.A1(new_n7225_), .A2(new_n7157_), .A3(new_n7214_), .A4(new_n7217_), .ZN(new_n7226_));
  NOR2_X1    g06213(.A1(new_n7226_), .A2(new_n7212_), .ZN(new_n7227_));
  OAI21_X1   g06214(.A1(new_n7209_), .A2(new_n7210_), .B(new_n7180_), .ZN(new_n7228_));
  NAND3_X1   g06215(.A1(new_n7204_), .A2(new_n7206_), .A3(new_n7192_), .ZN(new_n7229_));
  NAND2_X1   g06216(.A1(new_n7228_), .A2(new_n7229_), .ZN(new_n7230_));
  NOR2_X1    g06217(.A1(new_n7218_), .A2(new_n7124_), .ZN(new_n7231_));
  NAND2_X1   g06218(.A1(new_n7215_), .A2(new_n7218_), .ZN(new_n7232_));
  NAND2_X1   g06219(.A1(new_n7195_), .A2(new_n7197_), .ZN(new_n7233_));
  NAND2_X1   g06220(.A1(new_n7200_), .A2(new_n7202_), .ZN(new_n7234_));
  NAND2_X1   g06221(.A1(new_n7233_), .A2(new_n7234_), .ZN(new_n7235_));
  NAND2_X1   g06222(.A1(new_n7235_), .A2(new_n7203_), .ZN(new_n7236_));
  NOR4_X1    g06223(.A1(new_n7236_), .A2(new_n7232_), .A3(new_n7231_), .A4(new_n7216_), .ZN(new_n7237_));
  NAND2_X1   g06224(.A1(new_n7230_), .A2(new_n7237_), .ZN(new_n7238_));
  NAND2_X1   g06225(.A1(new_n7218_), .A2(new_n7123_), .ZN(new_n7239_));
  NAND3_X1   g06226(.A1(new_n7149_), .A2(new_n7155_), .A3(new_n7222_), .ZN(new_n7240_));
  AOI21_X1   g06227(.A1(new_n7239_), .A2(new_n7240_), .B(new_n7221_), .ZN(new_n7241_));
  AOI21_X1   g06228(.A1(new_n7149_), .A2(new_n7155_), .B(new_n7222_), .ZN(new_n7242_));
  NOR3_X1    g06229(.A1(new_n7133_), .A2(new_n7141_), .A3(new_n7123_), .ZN(new_n7243_));
  NOR3_X1    g06230(.A1(new_n7242_), .A2(new_n7243_), .A3(new_n7119_), .ZN(new_n7244_));
  NOR2_X1    g06231(.A1(new_n7241_), .A2(new_n7244_), .ZN(new_n7245_));
  OAI21_X1   g06232(.A1(new_n7230_), .A2(new_n7237_), .B(new_n7245_), .ZN(new_n7246_));
  NOR2_X1    g06233(.A1(new_n7203_), .A2(new_n7182_), .ZN(new_n7247_));
  NAND4_X1   g06234(.A1(new_n7157_), .A2(new_n7214_), .A3(new_n7143_), .A4(new_n7247_), .ZN(new_n7248_));
  OAI21_X1   g06235(.A1(new_n7242_), .A2(new_n7243_), .B(new_n7119_), .ZN(new_n7249_));
  NAND3_X1   g06236(.A1(new_n7239_), .A2(new_n7240_), .A3(new_n7221_), .ZN(new_n7250_));
  NAND2_X1   g06237(.A1(new_n7250_), .A2(new_n7249_), .ZN(new_n7251_));
  NAND3_X1   g06238(.A1(new_n7212_), .A2(new_n7251_), .A3(new_n7248_), .ZN(new_n7252_));
  NAND2_X1   g06239(.A1(new_n7246_), .A2(new_n7252_), .ZN(new_n7253_));
  AOI21_X1   g06240(.A1(new_n7253_), .A2(new_n7238_), .B(new_n7227_), .ZN(new_n7254_));
  OAI22_X1   g06241(.A1(new_n7254_), .A2(new_n7095_), .B1(new_n7186_), .B2(new_n7191_), .ZN(new_n7255_));
  NAND2_X1   g06242(.A1(new_n7013_), .A2(new_n7078_), .ZN(new_n7256_));
  NAND2_X1   g06243(.A1(new_n7256_), .A2(new_n7054_), .ZN(new_n7257_));
  OAI21_X1   g06244(.A1(new_n7057_), .A2(new_n7058_), .B(new_n7056_), .ZN(new_n7258_));
  NAND2_X1   g06245(.A1(new_n7258_), .A2(new_n7073_), .ZN(new_n7259_));
  INV_X1     g06246(.I(new_n7259_), .ZN(new_n7260_));
  NAND2_X1   g06247(.A1(new_n7099_), .A2(new_n7070_), .ZN(new_n7261_));
  AOI21_X1   g06248(.A1(new_n7261_), .A2(new_n7105_), .B(new_n7260_), .ZN(new_n7262_));
  NOR2_X1    g06249(.A1(new_n7061_), .A2(new_n7102_), .ZN(new_n7263_));
  NOR3_X1    g06250(.A1(new_n7263_), .A2(new_n7082_), .A3(new_n7259_), .ZN(new_n7264_));
  OAI21_X1   g06251(.A1(new_n7264_), .A2(new_n7262_), .B(new_n7257_), .ZN(new_n7265_));
  INV_X1     g06252(.I(new_n7257_), .ZN(new_n7266_));
  OAI21_X1   g06253(.A1(new_n7263_), .A2(new_n7082_), .B(new_n7259_), .ZN(new_n7267_));
  NAND3_X1   g06254(.A1(new_n7261_), .A2(new_n7105_), .A3(new_n7260_), .ZN(new_n7268_));
  NAND3_X1   g06255(.A1(new_n7267_), .A2(new_n7268_), .A3(new_n7266_), .ZN(new_n7269_));
  NAND2_X1   g06256(.A1(new_n7265_), .A2(new_n7269_), .ZN(new_n7270_));
  AOI21_X1   g06257(.A1(new_n7142_), .A2(new_n7223_), .B(new_n7125_), .ZN(new_n7271_));
  NAND2_X1   g06258(.A1(new_n7157_), .A2(new_n7214_), .ZN(new_n7272_));
  OAI21_X1   g06259(.A1(new_n7124_), .A2(new_n7156_), .B(new_n7247_), .ZN(new_n7273_));
  NOR4_X1    g06260(.A1(new_n7272_), .A2(new_n7273_), .A3(new_n7220_), .A4(new_n7224_), .ZN(new_n7274_));
  OAI21_X1   g06261(.A1(new_n7180_), .A2(new_n7181_), .B(new_n7208_), .ZN(new_n7275_));
  NAND2_X1   g06262(.A1(new_n7275_), .A2(new_n7182_), .ZN(new_n7276_));
  AOI21_X1   g06263(.A1(new_n7248_), .A2(new_n7245_), .B(new_n7212_), .ZN(new_n7277_));
  OAI21_X1   g06264(.A1(new_n7277_), .A2(new_n7274_), .B(new_n7276_), .ZN(new_n7278_));
  INV_X1     g06265(.I(new_n7276_), .ZN(new_n7279_));
  OAI21_X1   g06266(.A1(new_n7237_), .A2(new_n7251_), .B(new_n7230_), .ZN(new_n7280_));
  NAND3_X1   g06267(.A1(new_n7280_), .A2(new_n7226_), .A3(new_n7279_), .ZN(new_n7281_));
  AOI21_X1   g06268(.A1(new_n7278_), .A2(new_n7281_), .B(new_n7271_), .ZN(new_n7282_));
  INV_X1     g06269(.I(new_n7271_), .ZN(new_n7283_));
  AOI21_X1   g06270(.A1(new_n7280_), .A2(new_n7226_), .B(new_n7279_), .ZN(new_n7284_));
  NOR3_X1    g06271(.A1(new_n7277_), .A2(new_n7274_), .A3(new_n7276_), .ZN(new_n7285_));
  NOR3_X1    g06272(.A1(new_n7285_), .A2(new_n7284_), .A3(new_n7283_), .ZN(new_n7286_));
  NOR2_X1    g06273(.A1(new_n7286_), .A2(new_n7282_), .ZN(new_n7287_));
  NAND2_X1   g06274(.A1(new_n7270_), .A2(new_n7287_), .ZN(new_n7288_));
  AOI21_X1   g06275(.A1(new_n7267_), .A2(new_n7268_), .B(new_n7266_), .ZN(new_n7289_));
  NOR3_X1    g06276(.A1(new_n7264_), .A2(new_n7262_), .A3(new_n7257_), .ZN(new_n7290_));
  NOR2_X1    g06277(.A1(new_n7290_), .A2(new_n7289_), .ZN(new_n7291_));
  OAI21_X1   g06278(.A1(new_n7285_), .A2(new_n7284_), .B(new_n7283_), .ZN(new_n7292_));
  NAND3_X1   g06279(.A1(new_n7278_), .A2(new_n7281_), .A3(new_n7271_), .ZN(new_n7293_));
  NAND2_X1   g06280(.A1(new_n7292_), .A2(new_n7293_), .ZN(new_n7294_));
  NAND2_X1   g06281(.A1(new_n7291_), .A2(new_n7294_), .ZN(new_n7295_));
  AOI21_X1   g06282(.A1(new_n7288_), .A2(new_n7295_), .B(new_n7255_), .ZN(new_n7296_));
  INV_X1     g06283(.I(new_n7296_), .ZN(new_n7297_));
  NAND2_X1   g06284(.A1(new_n7109_), .A2(new_n7106_), .ZN(new_n7298_));
  OAI21_X1   g06285(.A1(new_n7083_), .A2(new_n7094_), .B(new_n7190_), .ZN(new_n7299_));
  NAND3_X1   g06286(.A1(new_n7109_), .A2(new_n7185_), .A3(new_n7106_), .ZN(new_n7300_));
  NAND2_X1   g06287(.A1(new_n7274_), .A2(new_n7230_), .ZN(new_n7301_));
  AOI21_X1   g06288(.A1(new_n7212_), .A2(new_n7248_), .B(new_n7251_), .ZN(new_n7302_));
  NOR3_X1    g06289(.A1(new_n7230_), .A2(new_n7245_), .A3(new_n7237_), .ZN(new_n7303_));
  OAI21_X1   g06290(.A1(new_n7302_), .A2(new_n7303_), .B(new_n7238_), .ZN(new_n7304_));
  NAND2_X1   g06291(.A1(new_n7304_), .A2(new_n7301_), .ZN(new_n7305_));
  AOI22_X1   g06292(.A1(new_n7305_), .A2(new_n7298_), .B1(new_n7299_), .B2(new_n7300_), .ZN(new_n7306_));
  NAND2_X1   g06293(.A1(new_n7291_), .A2(new_n7287_), .ZN(new_n7307_));
  NAND2_X1   g06294(.A1(new_n7270_), .A2(new_n7294_), .ZN(new_n7308_));
  AOI21_X1   g06295(.A1(new_n7307_), .A2(new_n7308_), .B(new_n7306_), .ZN(new_n7309_));
  INV_X1     g06296(.I(new_n7309_), .ZN(new_n7310_));
  NAND3_X1   g06297(.A1(new_n7297_), .A2(new_n7310_), .A3(new_n6976_), .ZN(new_n7311_));
  INV_X1     g06298(.I(new_n6940_), .ZN(new_n7312_));
  NAND2_X1   g06299(.A1(new_n7312_), .A2(new_n6942_), .ZN(new_n7313_));
  AOI21_X1   g06300(.A1(new_n6776_), .A2(new_n6702_), .B(new_n6793_), .ZN(new_n7314_));
  OAI21_X1   g06301(.A1(new_n7312_), .A2(new_n6942_), .B(new_n7314_), .ZN(new_n7315_));
  NAND2_X1   g06302(.A1(new_n7315_), .A2(new_n7313_), .ZN(new_n7316_));
  INV_X1     g06303(.I(new_n6973_), .ZN(new_n7317_));
  NAND3_X1   g06304(.A1(new_n6965_), .A2(new_n6958_), .A3(new_n6966_), .ZN(new_n7318_));
  NOR2_X1    g06305(.A1(new_n6970_), .A2(new_n6968_), .ZN(new_n7319_));
  INV_X1     g06306(.I(new_n6951_), .ZN(new_n7320_));
  INV_X1     g06307(.I(new_n6953_), .ZN(new_n7321_));
  NOR2_X1    g06308(.A1(new_n7321_), .A2(new_n7320_), .ZN(new_n7322_));
  NAND2_X1   g06309(.A1(new_n7321_), .A2(new_n7320_), .ZN(new_n7323_));
  AOI21_X1   g06310(.A1(new_n7319_), .A2(new_n7323_), .B(new_n7322_), .ZN(new_n7324_));
  AOI21_X1   g06311(.A1(new_n7318_), .A2(new_n7317_), .B(new_n7324_), .ZN(new_n7325_));
  AND4_X2    g06312(.A1(new_n6937_), .A2(new_n6967_), .A3(new_n6972_), .A4(new_n7324_), .Z(new_n7326_));
  OAI21_X1   g06313(.A1(new_n7325_), .A2(new_n7326_), .B(new_n7316_), .ZN(new_n7327_));
  INV_X1     g06314(.I(new_n7316_), .ZN(new_n7328_));
  NAND3_X1   g06315(.A1(new_n6937_), .A2(new_n6967_), .A3(new_n6972_), .ZN(new_n7329_));
  INV_X1     g06316(.I(new_n7324_), .ZN(new_n7330_));
  NAND2_X1   g06317(.A1(new_n7329_), .A2(new_n7330_), .ZN(new_n7331_));
  NAND4_X1   g06318(.A1(new_n6937_), .A2(new_n6967_), .A3(new_n6972_), .A4(new_n7324_), .ZN(new_n7332_));
  NAND3_X1   g06319(.A1(new_n7331_), .A2(new_n7328_), .A3(new_n7332_), .ZN(new_n7333_));
  NAND2_X1   g06320(.A1(new_n7327_), .A2(new_n7333_), .ZN(new_n7334_));
  NAND2_X1   g06321(.A1(new_n7261_), .A2(new_n7105_), .ZN(new_n7335_));
  NAND2_X1   g06322(.A1(new_n7259_), .A2(new_n7257_), .ZN(new_n7336_));
  NOR2_X1    g06323(.A1(new_n7259_), .A2(new_n7257_), .ZN(new_n7337_));
  OAI21_X1   g06324(.A1(new_n7335_), .A2(new_n7337_), .B(new_n7336_), .ZN(new_n7338_));
  NOR2_X1    g06325(.A1(new_n7279_), .A2(new_n7271_), .ZN(new_n7339_));
  NAND2_X1   g06326(.A1(new_n7280_), .A2(new_n7226_), .ZN(new_n7340_));
  NOR2_X1    g06327(.A1(new_n7276_), .A2(new_n7283_), .ZN(new_n7341_));
  NOR2_X1    g06328(.A1(new_n7340_), .A2(new_n7341_), .ZN(new_n7342_));
  NOR2_X1    g06329(.A1(new_n7342_), .A2(new_n7339_), .ZN(new_n7343_));
  OAI21_X1   g06330(.A1(new_n7270_), .A2(new_n7294_), .B(new_n7255_), .ZN(new_n7344_));
  XOR2_X1    g06331(.A1(new_n7259_), .A2(new_n7257_), .Z(new_n7345_));
  XOR2_X1    g06332(.A1(new_n7276_), .A2(new_n7283_), .Z(new_n7346_));
  NOR4_X1    g06333(.A1(new_n7335_), .A2(new_n7340_), .A3(new_n7345_), .A4(new_n7346_), .ZN(new_n7347_));
  AOI21_X1   g06334(.A1(new_n7344_), .A2(new_n7347_), .B(new_n7343_), .ZN(new_n7348_));
  INV_X1     g06335(.I(new_n7343_), .ZN(new_n7349_));
  AOI21_X1   g06336(.A1(new_n7291_), .A2(new_n7287_), .B(new_n7306_), .ZN(new_n7350_));
  INV_X1     g06337(.I(new_n7347_), .ZN(new_n7351_));
  NOR3_X1    g06338(.A1(new_n7350_), .A2(new_n7349_), .A3(new_n7351_), .ZN(new_n7352_));
  OAI21_X1   g06339(.A1(new_n7352_), .A2(new_n7348_), .B(new_n7338_), .ZN(new_n7353_));
  INV_X1     g06340(.I(new_n7338_), .ZN(new_n7354_));
  OAI21_X1   g06341(.A1(new_n7350_), .A2(new_n7351_), .B(new_n7349_), .ZN(new_n7355_));
  NAND3_X1   g06342(.A1(new_n7344_), .A2(new_n7343_), .A3(new_n7347_), .ZN(new_n7356_));
  NAND3_X1   g06343(.A1(new_n7355_), .A2(new_n7356_), .A3(new_n7354_), .ZN(new_n7357_));
  NAND3_X1   g06344(.A1(new_n7334_), .A2(new_n7353_), .A3(new_n7357_), .ZN(new_n7358_));
  AOI21_X1   g06345(.A1(new_n7331_), .A2(new_n7332_), .B(new_n7328_), .ZN(new_n7359_));
  NOR3_X1    g06346(.A1(new_n7325_), .A2(new_n7326_), .A3(new_n7316_), .ZN(new_n7360_));
  NOR2_X1    g06347(.A1(new_n7360_), .A2(new_n7359_), .ZN(new_n7361_));
  NAND2_X1   g06348(.A1(new_n7353_), .A2(new_n7357_), .ZN(new_n7362_));
  NAND2_X1   g06349(.A1(new_n7362_), .A2(new_n7361_), .ZN(new_n7363_));
  AOI21_X1   g06350(.A1(new_n7363_), .A2(new_n7358_), .B(new_n7311_), .ZN(new_n7364_));
  NAND2_X1   g06351(.A1(new_n6975_), .A2(new_n6957_), .ZN(new_n7365_));
  NOR3_X1    g06352(.A1(new_n7365_), .A2(new_n7296_), .A3(new_n7309_), .ZN(new_n7366_));
  NAND4_X1   g06353(.A1(new_n7353_), .A2(new_n7357_), .A3(new_n7327_), .A4(new_n7333_), .ZN(new_n7367_));
  AOI21_X1   g06354(.A1(new_n7355_), .A2(new_n7356_), .B(new_n7354_), .ZN(new_n7368_));
  NOR3_X1    g06355(.A1(new_n7352_), .A2(new_n7348_), .A3(new_n7338_), .ZN(new_n7369_));
  OAI22_X1   g06356(.A1(new_n7369_), .A2(new_n7368_), .B1(new_n7359_), .B2(new_n7360_), .ZN(new_n7370_));
  AOI21_X1   g06357(.A1(new_n7370_), .A2(new_n7367_), .B(new_n7366_), .ZN(new_n7371_));
  NOR4_X1    g06358(.A1(new_n7364_), .A2(new_n6641_), .A3(new_n6658_), .A4(new_n7371_), .ZN(new_n7372_));
  OAI21_X1   g06359(.A1(new_n7296_), .A2(new_n7309_), .B(new_n7365_), .ZN(new_n7373_));
  INV_X1     g06360(.I(new_n7373_), .ZN(new_n7374_));
  NOR2_X1    g06361(.A1(new_n7374_), .A2(new_n7366_), .ZN(new_n7375_));
  OAI21_X1   g06362(.A1(new_n6554_), .A2(new_n6566_), .B(new_n6645_), .ZN(new_n7376_));
  NAND3_X1   g06363(.A1(new_n6648_), .A2(new_n6230_), .A3(new_n6651_), .ZN(new_n7377_));
  AOI21_X1   g06364(.A1(new_n7376_), .A2(new_n7377_), .B(new_n6653_), .ZN(new_n7378_));
  INV_X1     g06365(.I(new_n7378_), .ZN(new_n7379_));
  AOI21_X1   g06366(.A1(new_n6652_), .A2(new_n6587_), .B(new_n6586_), .ZN(new_n7380_));
  INV_X1     g06367(.I(new_n7380_), .ZN(new_n7381_));
  NAND3_X1   g06368(.A1(new_n7379_), .A2(new_n7381_), .A3(new_n7375_), .ZN(new_n7382_));
  NAND4_X1   g06369(.A1(new_n6581_), .A2(new_n6582_), .A3(new_n6583_), .A4(new_n6584_), .ZN(new_n7383_));
  NAND2_X1   g06370(.A1(new_n7157_), .A2(new_n7143_), .ZN(new_n7384_));
  XOR2_X1    g06371(.A1(new_n7384_), .A2(new_n7110_), .Z(new_n7385_));
  NOR2_X1    g06372(.A1(new_n7385_), .A2(new_n7113_), .ZN(new_n7386_));
  NAND2_X1   g06373(.A1(new_n7385_), .A2(new_n7113_), .ZN(new_n7387_));
  INV_X1     g06374(.I(new_n7387_), .ZN(new_n7388_));
  NOR2_X1    g06375(.A1(new_n7388_), .A2(new_n7386_), .ZN(new_n7389_));
  INV_X1     g06376(.I(new_n7389_), .ZN(new_n7390_));
  OAI21_X1   g06377(.A1(new_n6797_), .A2(new_n6799_), .B(new_n6867_), .ZN(new_n7391_));
  NAND2_X1   g06378(.A1(new_n6868_), .A2(new_n7391_), .ZN(new_n7392_));
  NOR2_X1    g06379(.A1(new_n7390_), .A2(new_n7392_), .ZN(new_n7393_));
  INV_X1     g06380(.I(new_n7393_), .ZN(new_n7394_));
  NAND2_X1   g06381(.A1(new_n7390_), .A2(new_n7392_), .ZN(new_n7395_));
  NOR2_X1    g06382(.A1(new_n6574_), .A2(new_n6575_), .ZN(new_n7396_));
  NOR2_X1    g06383(.A1(new_n6578_), .A2(new_n6577_), .ZN(new_n7397_));
  NOR2_X1    g06384(.A1(new_n7396_), .A2(new_n7397_), .ZN(new_n7398_));
  NOR2_X1    g06385(.A1(new_n7398_), .A2(new_n6579_), .ZN(new_n7399_));
  NAND3_X1   g06386(.A1(new_n7394_), .A2(new_n7395_), .A3(new_n7399_), .ZN(new_n7400_));
  XNOR2_X1   g06387(.A1(new_n7400_), .A2(new_n7383_), .ZN(new_n7401_));
  NOR2_X1    g06388(.A1(new_n7400_), .A2(new_n7383_), .ZN(new_n7402_));
  NOR3_X1    g06389(.A1(new_n7305_), .A2(new_n7186_), .A3(new_n7191_), .ZN(new_n7403_));
  INV_X1     g06390(.I(new_n7403_), .ZN(new_n7404_));
  NOR3_X1    g06391(.A1(new_n6960_), .A2(new_n6964_), .A3(new_n6959_), .ZN(new_n7405_));
  INV_X1     g06392(.I(new_n7405_), .ZN(new_n7406_));
  AND3_X2    g06393(.A1(new_n7406_), .A2(new_n6965_), .A3(new_n7404_), .Z(new_n7407_));
  AOI21_X1   g06394(.A1(new_n7406_), .A2(new_n6965_), .B(new_n7404_), .ZN(new_n7408_));
  NOR2_X1    g06395(.A1(new_n7407_), .A2(new_n7408_), .ZN(new_n7409_));
  NOR2_X1    g06396(.A1(new_n7409_), .A2(new_n7393_), .ZN(new_n7410_));
  NOR3_X1    g06397(.A1(new_n7407_), .A2(new_n7394_), .A3(new_n7408_), .ZN(new_n7411_));
  NOR2_X1    g06398(.A1(new_n7410_), .A2(new_n7411_), .ZN(new_n7412_));
  AOI21_X1   g06399(.A1(new_n7401_), .A2(new_n7412_), .B(new_n7402_), .ZN(new_n7413_));
  AOI21_X1   g06400(.A1(new_n7379_), .A2(new_n7381_), .B(new_n7375_), .ZN(new_n7414_));
  OAI21_X1   g06401(.A1(new_n7413_), .A2(new_n7414_), .B(new_n7382_), .ZN(new_n7415_));
  OAI22_X1   g06402(.A1(new_n7364_), .A2(new_n7371_), .B1(new_n6641_), .B2(new_n6658_), .ZN(new_n7416_));
  AOI21_X1   g06403(.A1(new_n7415_), .A2(new_n7416_), .B(new_n7372_), .ZN(new_n7417_));
  NOR3_X1    g06404(.A1(new_n6639_), .A2(new_n6610_), .A3(new_n6606_), .ZN(new_n7418_));
  NAND2_X1   g06405(.A1(new_n6604_), .A2(new_n6597_), .ZN(new_n7419_));
  XOR2_X1    g06406(.A1(new_n6623_), .A2(new_n6614_), .Z(new_n7420_));
  XOR2_X1    g06407(.A1(new_n6592_), .A2(new_n6601_), .Z(new_n7421_));
  NOR4_X1    g06408(.A1(new_n7419_), .A2(new_n7421_), .A3(new_n6619_), .A4(new_n7420_), .ZN(new_n7422_));
  OAI21_X1   g06409(.A1(new_n7418_), .A2(new_n6655_), .B(new_n7422_), .ZN(new_n7423_));
  NOR2_X1    g06410(.A1(new_n6607_), .A2(new_n6602_), .ZN(new_n7424_));
  INV_X1     g06411(.I(new_n7424_), .ZN(new_n7425_));
  NOR2_X1    g06412(.A1(new_n6592_), .A2(new_n6601_), .ZN(new_n7426_));
  OR3_X2     g06413(.A1(new_n6593_), .A2(new_n6598_), .A3(new_n7426_), .Z(new_n7427_));
  NAND2_X1   g06414(.A1(new_n6623_), .A2(new_n6614_), .ZN(new_n7428_));
  NAND3_X1   g06415(.A1(new_n6615_), .A2(new_n6620_), .A3(new_n6622_), .ZN(new_n7429_));
  NAND3_X1   g06416(.A1(new_n6626_), .A2(new_n6625_), .A3(new_n7429_), .ZN(new_n7430_));
  NAND4_X1   g06417(.A1(new_n7427_), .A2(new_n7425_), .A3(new_n7428_), .A4(new_n7430_), .ZN(new_n7431_));
  NOR2_X1    g06418(.A1(new_n7419_), .A2(new_n7426_), .ZN(new_n7432_));
  NAND2_X1   g06419(.A1(new_n7430_), .A2(new_n7428_), .ZN(new_n7433_));
  OAI21_X1   g06420(.A1(new_n7432_), .A2(new_n7424_), .B(new_n7433_), .ZN(new_n7434_));
  AND2_X2    g06421(.A1(new_n7431_), .A2(new_n7434_), .Z(new_n7435_));
  NAND2_X1   g06422(.A1(new_n7423_), .A2(new_n7435_), .ZN(new_n7436_));
  NAND2_X1   g06423(.A1(new_n6656_), .A2(new_n6588_), .ZN(new_n7437_));
  NAND2_X1   g06424(.A1(new_n7431_), .A2(new_n7434_), .ZN(new_n7438_));
  NAND3_X1   g06425(.A1(new_n7437_), .A2(new_n7422_), .A3(new_n7438_), .ZN(new_n7439_));
  NAND2_X1   g06426(.A1(new_n7436_), .A2(new_n7439_), .ZN(new_n7440_));
  NAND2_X1   g06427(.A1(new_n7344_), .A2(new_n7347_), .ZN(new_n7441_));
  NAND2_X1   g06428(.A1(new_n7354_), .A2(new_n7343_), .ZN(new_n7442_));
  NOR2_X1    g06429(.A1(new_n7354_), .A2(new_n7343_), .ZN(new_n7443_));
  AOI21_X1   g06430(.A1(new_n7441_), .A2(new_n7442_), .B(new_n7443_), .ZN(new_n7444_));
  INV_X1     g06431(.I(new_n7444_), .ZN(new_n7445_));
  NOR2_X1    g06432(.A1(new_n7316_), .A2(new_n7330_), .ZN(new_n7446_));
  NOR2_X1    g06433(.A1(new_n7328_), .A2(new_n7324_), .ZN(new_n7447_));
  NOR2_X1    g06434(.A1(new_n7447_), .A2(new_n7329_), .ZN(new_n7448_));
  NOR2_X1    g06435(.A1(new_n7448_), .A2(new_n7446_), .ZN(new_n7449_));
  INV_X1     g06436(.I(new_n7449_), .ZN(new_n7450_));
  OAI21_X1   g06437(.A1(new_n7362_), .A2(new_n7334_), .B(new_n7311_), .ZN(new_n7451_));
  XOR2_X1    g06438(.A1(new_n7316_), .A2(new_n7330_), .Z(new_n7452_));
  XNOR2_X1   g06439(.A1(new_n7343_), .A2(new_n7338_), .ZN(new_n7453_));
  NOR4_X1    g06440(.A1(new_n7452_), .A2(new_n7441_), .A3(new_n7329_), .A4(new_n7453_), .ZN(new_n7454_));
  AOI21_X1   g06441(.A1(new_n7451_), .A2(new_n7454_), .B(new_n7450_), .ZN(new_n7455_));
  NOR2_X1    g06442(.A1(new_n7369_), .A2(new_n7368_), .ZN(new_n7456_));
  AOI21_X1   g06443(.A1(new_n7456_), .A2(new_n7361_), .B(new_n7366_), .ZN(new_n7457_));
  INV_X1     g06444(.I(new_n7454_), .ZN(new_n7458_));
  NOR3_X1    g06445(.A1(new_n7457_), .A2(new_n7449_), .A3(new_n7458_), .ZN(new_n7459_));
  OAI21_X1   g06446(.A1(new_n7459_), .A2(new_n7455_), .B(new_n7445_), .ZN(new_n7460_));
  OAI21_X1   g06447(.A1(new_n7457_), .A2(new_n7458_), .B(new_n7449_), .ZN(new_n7461_));
  NAND3_X1   g06448(.A1(new_n7451_), .A2(new_n7450_), .A3(new_n7454_), .ZN(new_n7462_));
  NAND3_X1   g06449(.A1(new_n7461_), .A2(new_n7462_), .A3(new_n7444_), .ZN(new_n7463_));
  NAND3_X1   g06450(.A1(new_n7440_), .A2(new_n7460_), .A3(new_n7463_), .ZN(new_n7464_));
  AOI21_X1   g06451(.A1(new_n7437_), .A2(new_n7422_), .B(new_n7438_), .ZN(new_n7465_));
  NOR2_X1    g06452(.A1(new_n7423_), .A2(new_n7435_), .ZN(new_n7466_));
  NOR2_X1    g06453(.A1(new_n7466_), .A2(new_n7465_), .ZN(new_n7467_));
  AOI21_X1   g06454(.A1(new_n7461_), .A2(new_n7462_), .B(new_n7444_), .ZN(new_n7468_));
  NOR3_X1    g06455(.A1(new_n7459_), .A2(new_n7455_), .A3(new_n7445_), .ZN(new_n7469_));
  OAI21_X1   g06456(.A1(new_n7468_), .A2(new_n7469_), .B(new_n7467_), .ZN(new_n7470_));
  AOI21_X1   g06457(.A1(new_n7470_), .A2(new_n7464_), .B(new_n7417_), .ZN(new_n7471_));
  AOI21_X1   g06458(.A1(new_n6635_), .A2(new_n6636_), .B(new_n6639_), .ZN(new_n7472_));
  NOR3_X1    g06459(.A1(new_n6633_), .A2(new_n6610_), .A3(new_n6606_), .ZN(new_n7473_));
  OAI21_X1   g06460(.A1(new_n7472_), .A2(new_n7473_), .B(new_n6655_), .ZN(new_n7474_));
  AOI21_X1   g06461(.A1(new_n6635_), .A2(new_n6636_), .B(new_n6633_), .ZN(new_n7475_));
  OAI21_X1   g06462(.A1(new_n7475_), .A2(new_n7418_), .B(new_n6588_), .ZN(new_n7476_));
  NOR2_X1    g06463(.A1(new_n7362_), .A2(new_n7361_), .ZN(new_n7477_));
  NOR2_X1    g06464(.A1(new_n7456_), .A2(new_n7334_), .ZN(new_n7478_));
  OAI21_X1   g06465(.A1(new_n7478_), .A2(new_n7477_), .B(new_n7366_), .ZN(new_n7479_));
  NOR3_X1    g06466(.A1(new_n7334_), .A2(new_n7368_), .A3(new_n7369_), .ZN(new_n7480_));
  AOI22_X1   g06467(.A1(new_n7353_), .A2(new_n7357_), .B1(new_n7327_), .B2(new_n7333_), .ZN(new_n7481_));
  OAI21_X1   g06468(.A1(new_n7480_), .A2(new_n7481_), .B(new_n7311_), .ZN(new_n7482_));
  NAND4_X1   g06469(.A1(new_n7479_), .A2(new_n7474_), .A3(new_n7482_), .A4(new_n7476_), .ZN(new_n7483_));
  NAND2_X1   g06470(.A1(new_n7311_), .A2(new_n7373_), .ZN(new_n7484_));
  NOR3_X1    g06471(.A1(new_n7484_), .A2(new_n7378_), .A3(new_n7380_), .ZN(new_n7485_));
  XOR2_X1    g06472(.A1(new_n7400_), .A2(new_n7383_), .Z(new_n7486_));
  OR2_X2     g06473(.A1(new_n7410_), .A2(new_n7411_), .Z(new_n7487_));
  AOI21_X1   g06474(.A1(new_n7487_), .A2(new_n7383_), .B(new_n7486_), .ZN(new_n7488_));
  OAI21_X1   g06475(.A1(new_n7378_), .A2(new_n7380_), .B(new_n7484_), .ZN(new_n7489_));
  AOI21_X1   g06476(.A1(new_n7488_), .A2(new_n7489_), .B(new_n7485_), .ZN(new_n7490_));
  AOI22_X1   g06477(.A1(new_n7479_), .A2(new_n7482_), .B1(new_n7474_), .B2(new_n7476_), .ZN(new_n7491_));
  OAI21_X1   g06478(.A1(new_n7490_), .A2(new_n7491_), .B(new_n7483_), .ZN(new_n7492_));
  NAND3_X1   g06479(.A1(new_n7467_), .A2(new_n7460_), .A3(new_n7463_), .ZN(new_n7493_));
  OAI21_X1   g06480(.A1(new_n7468_), .A2(new_n7469_), .B(new_n7440_), .ZN(new_n7494_));
  AOI21_X1   g06481(.A1(new_n7493_), .A2(new_n7494_), .B(new_n7492_), .ZN(new_n7495_));
  NOR4_X1    g06482(.A1(new_n5898_), .A2(new_n5923_), .A3(new_n7471_), .A4(new_n7495_), .ZN(new_n7496_));
  NAND2_X1   g06483(.A1(new_n7476_), .A2(new_n7474_), .ZN(new_n7497_));
  NOR2_X1    g06484(.A1(new_n7364_), .A2(new_n7371_), .ZN(new_n7498_));
  NOR2_X1    g06485(.A1(new_n7498_), .A2(new_n7497_), .ZN(new_n7499_));
  NOR2_X1    g06486(.A1(new_n6641_), .A2(new_n6658_), .ZN(new_n7500_));
  NOR3_X1    g06487(.A1(new_n7500_), .A2(new_n7364_), .A3(new_n7371_), .ZN(new_n7501_));
  OAI21_X1   g06488(.A1(new_n7499_), .A2(new_n7501_), .B(new_n7415_), .ZN(new_n7502_));
  OAI21_X1   g06489(.A1(new_n7372_), .A2(new_n7491_), .B(new_n7490_), .ZN(new_n7503_));
  NAND2_X1   g06490(.A1(new_n5901_), .A2(new_n5904_), .ZN(new_n7504_));
  NOR2_X1    g06491(.A1(new_n5782_), .A2(new_n5803_), .ZN(new_n7505_));
  NOR2_X1    g06492(.A1(new_n7505_), .A2(new_n7504_), .ZN(new_n7506_));
  NOR2_X1    g06493(.A1(new_n5043_), .A2(new_n5066_), .ZN(new_n7507_));
  NAND2_X1   g06494(.A1(new_n5910_), .A2(new_n5907_), .ZN(new_n7508_));
  NOR2_X1    g06495(.A1(new_n7508_), .A2(new_n7507_), .ZN(new_n7509_));
  OAI21_X1   g06496(.A1(new_n7509_), .A2(new_n7506_), .B(new_n5840_), .ZN(new_n7510_));
  OAI21_X1   g06497(.A1(new_n5919_), .A2(new_n5804_), .B(new_n5918_), .ZN(new_n7511_));
  NAND4_X1   g06498(.A1(new_n7510_), .A2(new_n7502_), .A3(new_n7503_), .A4(new_n7511_), .ZN(new_n7512_));
  NAND3_X1   g06499(.A1(new_n5916_), .A2(new_n5811_), .A3(new_n5813_), .ZN(new_n7513_));
  NAND3_X1   g06500(.A1(new_n5915_), .A2(new_n5820_), .A3(new_n5822_), .ZN(new_n7514_));
  AOI21_X1   g06501(.A1(new_n7514_), .A2(new_n7513_), .B(new_n5838_), .ZN(new_n7515_));
  AOI21_X1   g06502(.A1(new_n5917_), .A2(new_n5823_), .B(new_n5837_), .ZN(new_n7516_));
  OAI21_X1   g06503(.A1(new_n7378_), .A2(new_n7380_), .B(new_n7375_), .ZN(new_n7517_));
  NAND3_X1   g06504(.A1(new_n7379_), .A2(new_n7381_), .A3(new_n7484_), .ZN(new_n7518_));
  AOI21_X1   g06505(.A1(new_n7518_), .A2(new_n7517_), .B(new_n7413_), .ZN(new_n7519_));
  OAI21_X1   g06506(.A1(new_n7414_), .A2(new_n7485_), .B(new_n7413_), .ZN(new_n7520_));
  INV_X1     g06507(.I(new_n7520_), .ZN(new_n7521_));
  NOR4_X1    g06508(.A1(new_n7521_), .A2(new_n7515_), .A3(new_n7516_), .A4(new_n7519_), .ZN(new_n7522_));
  INV_X1     g06509(.I(new_n7522_), .ZN(new_n7523_));
  AOI22_X1   g06510(.A1(new_n7510_), .A2(new_n7511_), .B1(new_n7502_), .B2(new_n7503_), .ZN(new_n7524_));
  OAI21_X1   g06511(.A1(new_n7524_), .A2(new_n7523_), .B(new_n7512_), .ZN(new_n7525_));
  OAI22_X1   g06512(.A1(new_n5898_), .A2(new_n5923_), .B1(new_n7471_), .B2(new_n7495_), .ZN(new_n7526_));
  AOI21_X1   g06513(.A1(new_n7525_), .A2(new_n7526_), .B(new_n7496_), .ZN(new_n7527_));
  NAND2_X1   g06514(.A1(new_n5848_), .A2(new_n5851_), .ZN(new_n7528_));
  NOR3_X1    g06515(.A1(new_n5020_), .A2(new_n5019_), .A3(new_n5024_), .ZN(new_n7529_));
  AOI21_X1   g06516(.A1(new_n5020_), .A2(new_n5024_), .B(new_n5018_), .ZN(new_n7530_));
  NOR2_X1    g06517(.A1(new_n7529_), .A2(new_n7530_), .ZN(new_n7531_));
  NAND2_X1   g06518(.A1(new_n5852_), .A2(new_n5010_), .ZN(new_n7532_));
  NAND2_X1   g06519(.A1(new_n7532_), .A2(new_n5853_), .ZN(new_n7533_));
  OAI21_X1   g06520(.A1(new_n7531_), .A2(new_n7533_), .B(new_n7528_), .ZN(new_n7534_));
  NAND2_X1   g06521(.A1(new_n5847_), .A2(new_n5859_), .ZN(new_n7535_));
  NAND2_X1   g06522(.A1(new_n7534_), .A2(new_n7535_), .ZN(new_n7536_));
  NAND2_X1   g06523(.A1(new_n5882_), .A2(new_n5874_), .ZN(new_n7537_));
  NOR3_X1    g06524(.A1(new_n5758_), .A2(new_n5757_), .A3(new_n5763_), .ZN(new_n7538_));
  AOI21_X1   g06525(.A1(new_n5758_), .A2(new_n5763_), .B(new_n5756_), .ZN(new_n7539_));
  NOR2_X1    g06526(.A1(new_n7538_), .A2(new_n7539_), .ZN(new_n7540_));
  NAND2_X1   g06527(.A1(new_n5876_), .A2(new_n5749_), .ZN(new_n7541_));
  NAND2_X1   g06528(.A1(new_n7541_), .A2(new_n5877_), .ZN(new_n7542_));
  OAI21_X1   g06529(.A1(new_n7540_), .A2(new_n7542_), .B(new_n7537_), .ZN(new_n7543_));
  NAND2_X1   g06530(.A1(new_n5885_), .A2(new_n5880_), .ZN(new_n7544_));
  NAND2_X1   g06531(.A1(new_n7543_), .A2(new_n7544_), .ZN(new_n7545_));
  INV_X1     g06532(.I(new_n7545_), .ZN(new_n7546_));
  NAND2_X1   g06533(.A1(new_n5842_), .A2(new_n5921_), .ZN(new_n7547_));
  XOR2_X1    g06534(.A1(new_n5846_), .A2(new_n5855_), .Z(new_n7548_));
  XOR2_X1    g06535(.A1(new_n5869_), .A2(new_n5879_), .Z(new_n7549_));
  NOR4_X1    g06536(.A1(new_n7537_), .A2(new_n7549_), .A3(new_n7548_), .A4(new_n7528_), .ZN(new_n7550_));
  AOI21_X1   g06537(.A1(new_n7547_), .A2(new_n7550_), .B(new_n7546_), .ZN(new_n7551_));
  NOR4_X1    g06538(.A1(new_n5892_), .A2(new_n5884_), .A3(new_n5888_), .A4(new_n5891_), .ZN(new_n7552_));
  OAI21_X1   g06539(.A1(new_n7552_), .A2(new_n5920_), .B(new_n7550_), .ZN(new_n7553_));
  NOR2_X1    g06540(.A1(new_n7553_), .A2(new_n7545_), .ZN(new_n7554_));
  OAI21_X1   g06541(.A1(new_n7554_), .A2(new_n7551_), .B(new_n7536_), .ZN(new_n7555_));
  INV_X1     g06542(.I(new_n7536_), .ZN(new_n7556_));
  NAND2_X1   g06543(.A1(new_n7553_), .A2(new_n7545_), .ZN(new_n7557_));
  NAND3_X1   g06544(.A1(new_n7547_), .A2(new_n7546_), .A3(new_n7550_), .ZN(new_n7558_));
  NAND3_X1   g06545(.A1(new_n7557_), .A2(new_n7558_), .A3(new_n7556_), .ZN(new_n7559_));
  NAND2_X1   g06546(.A1(new_n7555_), .A2(new_n7559_), .ZN(new_n7560_));
  NAND2_X1   g06547(.A1(new_n6607_), .A2(new_n6602_), .ZN(new_n7561_));
  NAND2_X1   g06548(.A1(new_n7425_), .A2(new_n7419_), .ZN(new_n7562_));
  NAND4_X1   g06549(.A1(new_n7562_), .A2(new_n7561_), .A3(new_n7428_), .A4(new_n7430_), .ZN(new_n7563_));
  NAND2_X1   g06550(.A1(new_n7423_), .A2(new_n7563_), .ZN(new_n7564_));
  NAND3_X1   g06551(.A1(new_n7427_), .A2(new_n7425_), .A3(new_n7433_), .ZN(new_n7565_));
  NAND2_X1   g06552(.A1(new_n7564_), .A2(new_n7565_), .ZN(new_n7566_));
  INV_X1     g06553(.I(new_n7566_), .ZN(new_n7567_));
  NAND2_X1   g06554(.A1(new_n7451_), .A2(new_n7454_), .ZN(new_n7568_));
  OR4_X2     g06555(.A1(new_n7328_), .A2(new_n7444_), .A3(new_n7329_), .A4(new_n7324_), .Z(new_n7569_));
  AOI22_X1   g06556(.A1(new_n7568_), .A2(new_n7569_), .B1(new_n7445_), .B2(new_n7449_), .ZN(new_n7570_));
  NOR3_X1    g06557(.A1(new_n7468_), .A2(new_n7469_), .A3(new_n7440_), .ZN(new_n7571_));
  XNOR2_X1   g06558(.A1(new_n7449_), .A2(new_n7444_), .ZN(new_n7572_));
  NOR4_X1    g06559(.A1(new_n7568_), .A2(new_n7423_), .A3(new_n7438_), .A4(new_n7572_), .ZN(new_n7573_));
  OAI21_X1   g06560(.A1(new_n7571_), .A2(new_n7492_), .B(new_n7573_), .ZN(new_n7574_));
  NAND2_X1   g06561(.A1(new_n7574_), .A2(new_n7570_), .ZN(new_n7575_));
  INV_X1     g06562(.I(new_n7570_), .ZN(new_n7576_));
  NAND2_X1   g06563(.A1(new_n7417_), .A2(new_n7493_), .ZN(new_n7577_));
  NAND3_X1   g06564(.A1(new_n7577_), .A2(new_n7576_), .A3(new_n7573_), .ZN(new_n7578_));
  AOI21_X1   g06565(.A1(new_n7575_), .A2(new_n7578_), .B(new_n7567_), .ZN(new_n7579_));
  AOI21_X1   g06566(.A1(new_n7577_), .A2(new_n7573_), .B(new_n7576_), .ZN(new_n7580_));
  NOR2_X1    g06567(.A1(new_n7574_), .A2(new_n7570_), .ZN(new_n7581_));
  NOR3_X1    g06568(.A1(new_n7581_), .A2(new_n7580_), .A3(new_n7566_), .ZN(new_n7582_));
  NOR2_X1    g06569(.A1(new_n7582_), .A2(new_n7579_), .ZN(new_n7583_));
  NAND2_X1   g06570(.A1(new_n7583_), .A2(new_n7560_), .ZN(new_n7584_));
  AOI21_X1   g06571(.A1(new_n7557_), .A2(new_n7558_), .B(new_n7556_), .ZN(new_n7585_));
  NOR3_X1    g06572(.A1(new_n7554_), .A2(new_n7551_), .A3(new_n7536_), .ZN(new_n7586_));
  NOR2_X1    g06573(.A1(new_n7586_), .A2(new_n7585_), .ZN(new_n7587_));
  OAI21_X1   g06574(.A1(new_n7581_), .A2(new_n7580_), .B(new_n7566_), .ZN(new_n7588_));
  NAND3_X1   g06575(.A1(new_n7575_), .A2(new_n7578_), .A3(new_n7567_), .ZN(new_n7589_));
  NAND2_X1   g06576(.A1(new_n7588_), .A2(new_n7589_), .ZN(new_n7590_));
  NAND2_X1   g06577(.A1(new_n7587_), .A2(new_n7590_), .ZN(new_n7591_));
  AOI21_X1   g06578(.A1(new_n7584_), .A2(new_n7591_), .B(new_n7527_), .ZN(new_n7592_));
  NOR2_X1    g06579(.A1(new_n5893_), .A2(new_n5896_), .ZN(new_n7593_));
  NOR2_X1    g06580(.A1(new_n5889_), .A2(new_n5865_), .ZN(new_n7594_));
  OAI21_X1   g06581(.A1(new_n7593_), .A2(new_n7594_), .B(new_n5920_), .ZN(new_n7595_));
  AOI22_X1   g06582(.A1(new_n5894_), .A2(new_n5895_), .B1(new_n5861_), .B2(new_n5864_), .ZN(new_n7596_));
  OAI21_X1   g06583(.A1(new_n7552_), .A2(new_n7596_), .B(new_n5842_), .ZN(new_n7597_));
  NOR3_X1    g06584(.A1(new_n7467_), .A2(new_n7469_), .A3(new_n7468_), .ZN(new_n7598_));
  AOI21_X1   g06585(.A1(new_n7460_), .A2(new_n7463_), .B(new_n7440_), .ZN(new_n7599_));
  OAI21_X1   g06586(.A1(new_n7598_), .A2(new_n7599_), .B(new_n7492_), .ZN(new_n7600_));
  AOI21_X1   g06587(.A1(new_n7460_), .A2(new_n7463_), .B(new_n7467_), .ZN(new_n7601_));
  OAI21_X1   g06588(.A1(new_n7601_), .A2(new_n7571_), .B(new_n7417_), .ZN(new_n7602_));
  NAND4_X1   g06589(.A1(new_n7595_), .A2(new_n7597_), .A3(new_n7600_), .A4(new_n7602_), .ZN(new_n7603_));
  OAI21_X1   g06590(.A1(new_n7364_), .A2(new_n7371_), .B(new_n7500_), .ZN(new_n7604_));
  NAND2_X1   g06591(.A1(new_n7498_), .A2(new_n7497_), .ZN(new_n7605_));
  AOI21_X1   g06592(.A1(new_n7604_), .A2(new_n7605_), .B(new_n7490_), .ZN(new_n7606_));
  AOI21_X1   g06593(.A1(new_n7483_), .A2(new_n7416_), .B(new_n7415_), .ZN(new_n7607_));
  NAND2_X1   g06594(.A1(new_n7508_), .A2(new_n7507_), .ZN(new_n7608_));
  NAND2_X1   g06595(.A1(new_n7505_), .A2(new_n7504_), .ZN(new_n7609_));
  AOI21_X1   g06596(.A1(new_n7608_), .A2(new_n7609_), .B(new_n5918_), .ZN(new_n7610_));
  AOI21_X1   g06597(.A1(new_n5841_), .A2(new_n5911_), .B(new_n5840_), .ZN(new_n7611_));
  NOR4_X1    g06598(.A1(new_n7606_), .A2(new_n7610_), .A3(new_n7607_), .A4(new_n7611_), .ZN(new_n7612_));
  OAI22_X1   g06599(.A1(new_n7606_), .A2(new_n7607_), .B1(new_n7610_), .B2(new_n7611_), .ZN(new_n7613_));
  AOI21_X1   g06600(.A1(new_n7613_), .A2(new_n7522_), .B(new_n7612_), .ZN(new_n7614_));
  AOI22_X1   g06601(.A1(new_n7595_), .A2(new_n7597_), .B1(new_n7600_), .B2(new_n7602_), .ZN(new_n7615_));
  OAI21_X1   g06602(.A1(new_n7614_), .A2(new_n7615_), .B(new_n7603_), .ZN(new_n7616_));
  NAND4_X1   g06603(.A1(new_n7555_), .A2(new_n7559_), .A3(new_n7588_), .A4(new_n7589_), .ZN(new_n7617_));
  OAI22_X1   g06604(.A1(new_n7585_), .A2(new_n7586_), .B1(new_n7582_), .B2(new_n7579_), .ZN(new_n7618_));
  AOI21_X1   g06605(.A1(new_n7618_), .A2(new_n7617_), .B(new_n7616_), .ZN(new_n7619_));
  NOR4_X1    g06606(.A1(new_n7592_), .A2(new_n4282_), .A3(new_n4325_), .A4(new_n7619_), .ZN(new_n7620_));
  NAND2_X1   g06607(.A1(new_n7600_), .A2(new_n7602_), .ZN(new_n7621_));
  NAND3_X1   g06608(.A1(new_n7621_), .A2(new_n7595_), .A3(new_n7597_), .ZN(new_n7622_));
  NAND2_X1   g06609(.A1(new_n7595_), .A2(new_n7597_), .ZN(new_n7623_));
  NOR2_X1    g06610(.A1(new_n7495_), .A2(new_n7471_), .ZN(new_n7624_));
  NAND2_X1   g06611(.A1(new_n7623_), .A2(new_n7624_), .ZN(new_n7625_));
  AOI21_X1   g06612(.A1(new_n7625_), .A2(new_n7622_), .B(new_n7614_), .ZN(new_n7626_));
  AOI21_X1   g06613(.A1(new_n7603_), .A2(new_n7526_), .B(new_n7525_), .ZN(new_n7627_));
  NOR2_X1    g06614(.A1(new_n7626_), .A2(new_n7627_), .ZN(new_n7628_));
  NOR2_X1    g06615(.A1(new_n2573_), .A2(new_n2596_), .ZN(new_n7629_));
  NAND2_X1   g06616(.A1(new_n4292_), .A2(new_n4290_), .ZN(new_n7630_));
  NAND2_X1   g06617(.A1(new_n7630_), .A2(new_n7629_), .ZN(new_n7631_));
  NAND2_X1   g06618(.A1(new_n4287_), .A2(new_n4285_), .ZN(new_n7632_));
  NOR2_X1    g06619(.A1(new_n4149_), .A2(new_n4175_), .ZN(new_n7633_));
  NAND2_X1   g06620(.A1(new_n7633_), .A2(new_n7632_), .ZN(new_n7634_));
  AOI21_X1   g06621(.A1(new_n7631_), .A2(new_n7634_), .B(new_n4318_), .ZN(new_n7635_));
  AOI21_X1   g06622(.A1(new_n4293_), .A2(new_n4226_), .B(new_n4225_), .ZN(new_n7636_));
  NOR2_X1    g06623(.A1(new_n7635_), .A2(new_n7636_), .ZN(new_n7637_));
  NAND2_X1   g06624(.A1(new_n7628_), .A2(new_n7637_), .ZN(new_n7638_));
  NOR2_X1    g06625(.A1(new_n4296_), .A2(new_n4297_), .ZN(new_n7639_));
  NAND2_X1   g06626(.A1(new_n4191_), .A2(new_n4192_), .ZN(new_n7640_));
  NAND2_X1   g06627(.A1(new_n7639_), .A2(new_n7640_), .ZN(new_n7641_));
  NAND2_X1   g06628(.A1(new_n4183_), .A2(new_n4184_), .ZN(new_n7642_));
  NOR2_X1    g06629(.A1(new_n4300_), .A2(new_n4301_), .ZN(new_n7643_));
  NAND2_X1   g06630(.A1(new_n7642_), .A2(new_n7643_), .ZN(new_n7644_));
  AOI21_X1   g06631(.A1(new_n7644_), .A2(new_n7641_), .B(new_n4223_), .ZN(new_n7645_));
  AOI21_X1   g06632(.A1(new_n4317_), .A2(new_n4193_), .B(new_n4316_), .ZN(new_n7646_));
  NOR2_X1    g06633(.A1(new_n7606_), .A2(new_n7607_), .ZN(new_n7647_));
  NAND2_X1   g06634(.A1(new_n7510_), .A2(new_n7511_), .ZN(new_n7648_));
  NAND2_X1   g06635(.A1(new_n7647_), .A2(new_n7648_), .ZN(new_n7649_));
  NAND2_X1   g06636(.A1(new_n7502_), .A2(new_n7503_), .ZN(new_n7650_));
  NOR2_X1    g06637(.A1(new_n7610_), .A2(new_n7611_), .ZN(new_n7651_));
  NAND2_X1   g06638(.A1(new_n7651_), .A2(new_n7650_), .ZN(new_n7652_));
  AOI21_X1   g06639(.A1(new_n7649_), .A2(new_n7652_), .B(new_n7523_), .ZN(new_n7653_));
  AOI21_X1   g06640(.A1(new_n7613_), .A2(new_n7512_), .B(new_n7522_), .ZN(new_n7654_));
  NOR4_X1    g06641(.A1(new_n7653_), .A2(new_n7645_), .A3(new_n7646_), .A4(new_n7654_), .ZN(new_n7655_));
  OAI22_X1   g06642(.A1(new_n7521_), .A2(new_n7519_), .B1(new_n7515_), .B2(new_n7516_), .ZN(new_n7656_));
  INV_X1     g06643(.I(new_n7656_), .ZN(new_n7657_));
  NOR2_X1    g06644(.A1(new_n7657_), .A2(new_n7522_), .ZN(new_n7658_));
  NOR2_X1    g06645(.A1(new_n4206_), .A2(new_n4207_), .ZN(new_n7659_));
  NOR3_X1    g06646(.A1(new_n7659_), .A2(new_n4202_), .A3(new_n4203_), .ZN(new_n7660_));
  NOR2_X1    g06647(.A1(new_n4202_), .A2(new_n4203_), .ZN(new_n7661_));
  NAND2_X1   g06648(.A1(new_n4310_), .A2(new_n4309_), .ZN(new_n7662_));
  NOR2_X1    g06649(.A1(new_n7661_), .A2(new_n7662_), .ZN(new_n7663_));
  OAI21_X1   g06650(.A1(new_n7663_), .A2(new_n7660_), .B(new_n4221_), .ZN(new_n7664_));
  OAI21_X1   g06651(.A1(new_n4315_), .A2(new_n4208_), .B(new_n4314_), .ZN(new_n7665_));
  NAND3_X1   g06652(.A1(new_n7658_), .A2(new_n7665_), .A3(new_n7664_), .ZN(new_n7666_));
  NAND2_X1   g06653(.A1(new_n4218_), .A2(new_n4219_), .ZN(new_n7667_));
  INV_X1     g06654(.I(new_n7667_), .ZN(new_n7668_));
  NAND2_X1   g06655(.A1(new_n4212_), .A2(new_n4215_), .ZN(new_n7669_));
  NAND2_X1   g06656(.A1(new_n4217_), .A2(new_n7669_), .ZN(new_n7670_));
  NAND2_X1   g06657(.A1(new_n7394_), .A2(new_n7395_), .ZN(new_n7671_));
  XNOR2_X1   g06658(.A1(new_n7671_), .A2(new_n7399_), .ZN(new_n7672_));
  NAND2_X1   g06659(.A1(new_n5827_), .A2(new_n5830_), .ZN(new_n7673_));
  NAND2_X1   g06660(.A1(new_n5832_), .A2(new_n7673_), .ZN(new_n7674_));
  INV_X1     g06661(.I(new_n7674_), .ZN(new_n7675_));
  NAND2_X1   g06662(.A1(new_n7672_), .A2(new_n7675_), .ZN(new_n7676_));
  OR2_X2     g06663(.A1(new_n7672_), .A2(new_n7675_), .Z(new_n7677_));
  NAND2_X1   g06664(.A1(new_n7677_), .A2(new_n7676_), .ZN(new_n7678_));
  NOR2_X1    g06665(.A1(new_n7678_), .A2(new_n7670_), .ZN(new_n7679_));
  INV_X1     g06666(.I(new_n7679_), .ZN(new_n7680_));
  NAND2_X1   g06667(.A1(new_n7680_), .A2(new_n7667_), .ZN(new_n7681_));
  NAND2_X1   g06668(.A1(new_n7668_), .A2(new_n7679_), .ZN(new_n7682_));
  NAND2_X1   g06669(.A1(new_n7682_), .A2(new_n7681_), .ZN(new_n7683_));
  NAND2_X1   g06670(.A1(new_n7412_), .A2(new_n7486_), .ZN(new_n7684_));
  NAND2_X1   g06671(.A1(new_n5833_), .A2(new_n5834_), .ZN(new_n7685_));
  XNOR2_X1   g06672(.A1(new_n5836_), .A2(new_n7685_), .ZN(new_n7686_));
  NAND2_X1   g06673(.A1(new_n7686_), .A2(new_n7684_), .ZN(new_n7687_));
  INV_X1     g06674(.I(new_n7684_), .ZN(new_n7688_));
  XOR2_X1    g06675(.A1(new_n5836_), .A2(new_n7685_), .Z(new_n7689_));
  NAND2_X1   g06676(.A1(new_n7689_), .A2(new_n7688_), .ZN(new_n7690_));
  AOI22_X1   g06677(.A1(new_n7687_), .A2(new_n7690_), .B1(new_n7672_), .B2(new_n7675_), .ZN(new_n7691_));
  NOR2_X1    g06678(.A1(new_n7689_), .A2(new_n7688_), .ZN(new_n7692_));
  NOR2_X1    g06679(.A1(new_n7686_), .A2(new_n7684_), .ZN(new_n7693_));
  NOR3_X1    g06680(.A1(new_n7692_), .A2(new_n7693_), .A3(new_n7676_), .ZN(new_n7694_));
  NOR2_X1    g06681(.A1(new_n7691_), .A2(new_n7694_), .ZN(new_n7695_));
  OAI21_X1   g06682(.A1(new_n7695_), .A2(new_n7668_), .B(new_n7683_), .ZN(new_n7696_));
  AOI21_X1   g06683(.A1(new_n7664_), .A2(new_n7665_), .B(new_n7658_), .ZN(new_n7697_));
  OAI21_X1   g06684(.A1(new_n7696_), .A2(new_n7697_), .B(new_n7666_), .ZN(new_n7698_));
  OAI22_X1   g06685(.A1(new_n7653_), .A2(new_n7654_), .B1(new_n7645_), .B2(new_n7646_), .ZN(new_n7699_));
  AOI21_X1   g06686(.A1(new_n7699_), .A2(new_n7698_), .B(new_n7655_), .ZN(new_n7700_));
  NOR2_X1    g06687(.A1(new_n7623_), .A2(new_n7624_), .ZN(new_n7701_));
  AOI21_X1   g06688(.A1(new_n7595_), .A2(new_n7597_), .B(new_n7621_), .ZN(new_n7702_));
  OAI21_X1   g06689(.A1(new_n7702_), .A2(new_n7701_), .B(new_n7525_), .ZN(new_n7703_));
  OAI21_X1   g06690(.A1(new_n7496_), .A2(new_n7615_), .B(new_n7614_), .ZN(new_n7704_));
  NOR2_X1    g06691(.A1(new_n7633_), .A2(new_n7632_), .ZN(new_n7705_));
  NOR2_X1    g06692(.A1(new_n7630_), .A2(new_n7629_), .ZN(new_n7706_));
  OAI21_X1   g06693(.A1(new_n7706_), .A2(new_n7705_), .B(new_n4225_), .ZN(new_n7707_));
  OAI21_X1   g06694(.A1(new_n4176_), .A2(new_n4319_), .B(new_n4318_), .ZN(new_n7708_));
  AOI22_X1   g06695(.A1(new_n7703_), .A2(new_n7704_), .B1(new_n7707_), .B2(new_n7708_), .ZN(new_n7709_));
  OAI21_X1   g06696(.A1(new_n7700_), .A2(new_n7709_), .B(new_n7638_), .ZN(new_n7710_));
  NOR2_X1    g06697(.A1(new_n4280_), .A2(new_n4279_), .ZN(new_n7711_));
  NOR2_X1    g06698(.A1(new_n4322_), .A2(new_n4323_), .ZN(new_n7712_));
  NOR2_X1    g06699(.A1(new_n7712_), .A2(new_n4253_), .ZN(new_n7713_));
  OAI21_X1   g06700(.A1(new_n7713_), .A2(new_n7711_), .B(new_n4320_), .ZN(new_n7714_));
  NOR2_X1    g06701(.A1(new_n4280_), .A2(new_n4253_), .ZN(new_n7715_));
  AOI22_X1   g06702(.A1(new_n4271_), .A2(new_n4275_), .B1(new_n4248_), .B2(new_n4252_), .ZN(new_n7716_));
  OAI21_X1   g06703(.A1(new_n7715_), .A2(new_n7716_), .B(new_n4227_), .ZN(new_n7717_));
  NAND2_X1   g06704(.A1(new_n7714_), .A2(new_n7717_), .ZN(new_n7718_));
  NOR2_X1    g06705(.A1(new_n7587_), .A2(new_n7590_), .ZN(new_n7719_));
  NOR2_X1    g06706(.A1(new_n7583_), .A2(new_n7560_), .ZN(new_n7720_));
  OAI21_X1   g06707(.A1(new_n7720_), .A2(new_n7719_), .B(new_n7616_), .ZN(new_n7721_));
  NOR2_X1    g06708(.A1(new_n7560_), .A2(new_n7590_), .ZN(new_n7722_));
  AOI22_X1   g06709(.A1(new_n7555_), .A2(new_n7559_), .B1(new_n7588_), .B2(new_n7589_), .ZN(new_n7723_));
  OAI21_X1   g06710(.A1(new_n7722_), .A2(new_n7723_), .B(new_n7527_), .ZN(new_n7724_));
  NAND2_X1   g06711(.A1(new_n7721_), .A2(new_n7724_), .ZN(new_n7725_));
  NAND2_X1   g06712(.A1(new_n7725_), .A2(new_n7718_), .ZN(new_n7726_));
  AOI21_X1   g06713(.A1(new_n7726_), .A2(new_n7710_), .B(new_n7620_), .ZN(new_n7727_));
  OAI21_X1   g06714(.A1(new_n4259_), .A2(new_n4263_), .B(new_n4269_), .ZN(new_n7728_));
  NAND2_X1   g06715(.A1(new_n4259_), .A2(new_n4262_), .ZN(new_n7729_));
  NAND2_X1   g06716(.A1(new_n7728_), .A2(new_n7729_), .ZN(new_n7730_));
  NAND2_X1   g06717(.A1(new_n4321_), .A2(new_n4227_), .ZN(new_n7731_));
  NAND2_X1   g06718(.A1(new_n4239_), .A2(new_n4233_), .ZN(new_n7732_));
  NAND2_X1   g06719(.A1(new_n4249_), .A2(new_n4238_), .ZN(new_n7733_));
  NAND2_X1   g06720(.A1(new_n7733_), .A2(new_n7732_), .ZN(new_n7734_));
  XOR2_X1    g06721(.A1(new_n4259_), .A2(new_n4262_), .Z(new_n7735_));
  NOR4_X1    g06722(.A1(new_n7734_), .A2(new_n4269_), .A3(new_n7735_), .A4(new_n4246_), .ZN(new_n7736_));
  NOR2_X1    g06723(.A1(new_n4249_), .A2(new_n4239_), .ZN(new_n7737_));
  AOI21_X1   g06724(.A1(new_n4246_), .A2(new_n7733_), .B(new_n7737_), .ZN(new_n7738_));
  AOI21_X1   g06725(.A1(new_n7731_), .A2(new_n7736_), .B(new_n7738_), .ZN(new_n7739_));
  AOI21_X1   g06726(.A1(new_n7712_), .A2(new_n4279_), .B(new_n4320_), .ZN(new_n7740_));
  INV_X1     g06727(.I(new_n7736_), .ZN(new_n7741_));
  INV_X1     g06728(.I(new_n7738_), .ZN(new_n7742_));
  NOR3_X1    g06729(.A1(new_n7740_), .A2(new_n7741_), .A3(new_n7742_), .ZN(new_n7743_));
  OAI21_X1   g06730(.A1(new_n7743_), .A2(new_n7739_), .B(new_n7730_), .ZN(new_n7744_));
  INV_X1     g06731(.I(new_n7730_), .ZN(new_n7745_));
  OAI21_X1   g06732(.A1(new_n7740_), .A2(new_n7741_), .B(new_n7742_), .ZN(new_n7746_));
  NAND3_X1   g06733(.A1(new_n7731_), .A2(new_n7736_), .A3(new_n7738_), .ZN(new_n7747_));
  NAND3_X1   g06734(.A1(new_n7746_), .A2(new_n7747_), .A3(new_n7745_), .ZN(new_n7748_));
  OAI21_X1   g06735(.A1(new_n7566_), .A2(new_n7576_), .B(new_n7574_), .ZN(new_n7749_));
  NAND2_X1   g06736(.A1(new_n7566_), .A2(new_n7570_), .ZN(new_n7750_));
  NAND2_X1   g06737(.A1(new_n7749_), .A2(new_n7750_), .ZN(new_n7751_));
  NAND2_X1   g06738(.A1(new_n7617_), .A2(new_n7527_), .ZN(new_n7752_));
  INV_X1     g06739(.I(new_n7553_), .ZN(new_n7753_));
  INV_X1     g06740(.I(new_n7574_), .ZN(new_n7754_));
  XNOR2_X1   g06741(.A1(new_n7545_), .A2(new_n7536_), .ZN(new_n7755_));
  XNOR2_X1   g06742(.A1(new_n7566_), .A2(new_n7570_), .ZN(new_n7756_));
  NAND4_X1   g06743(.A1(new_n7753_), .A2(new_n7754_), .A3(new_n7755_), .A4(new_n7756_), .ZN(new_n7757_));
  INV_X1     g06744(.I(new_n7757_), .ZN(new_n7758_));
  NOR2_X1    g06745(.A1(new_n7545_), .A2(new_n7536_), .ZN(new_n7759_));
  NOR2_X1    g06746(.A1(new_n7546_), .A2(new_n7556_), .ZN(new_n7760_));
  AOI21_X1   g06747(.A1(new_n7553_), .A2(new_n7759_), .B(new_n7760_), .ZN(new_n7761_));
  AOI21_X1   g06748(.A1(new_n7752_), .A2(new_n7758_), .B(new_n7761_), .ZN(new_n7762_));
  AOI21_X1   g06749(.A1(new_n7587_), .A2(new_n7583_), .B(new_n7616_), .ZN(new_n7763_));
  INV_X1     g06750(.I(new_n7761_), .ZN(new_n7764_));
  NOR3_X1    g06751(.A1(new_n7763_), .A2(new_n7757_), .A3(new_n7764_), .ZN(new_n7765_));
  OAI21_X1   g06752(.A1(new_n7762_), .A2(new_n7765_), .B(new_n7751_), .ZN(new_n7766_));
  INV_X1     g06753(.I(new_n7751_), .ZN(new_n7767_));
  OAI21_X1   g06754(.A1(new_n7763_), .A2(new_n7757_), .B(new_n7764_), .ZN(new_n7768_));
  NAND3_X1   g06755(.A1(new_n7752_), .A2(new_n7758_), .A3(new_n7761_), .ZN(new_n7769_));
  NAND3_X1   g06756(.A1(new_n7769_), .A2(new_n7768_), .A3(new_n7767_), .ZN(new_n7770_));
  NAND4_X1   g06757(.A1(new_n7766_), .A2(new_n7770_), .A3(new_n7744_), .A4(new_n7748_), .ZN(new_n7771_));
  NAND2_X1   g06758(.A1(new_n7727_), .A2(new_n7771_), .ZN(new_n7772_));
  NAND2_X1   g06759(.A1(new_n7731_), .A2(new_n7736_), .ZN(new_n7773_));
  NAND2_X1   g06760(.A1(new_n7752_), .A2(new_n7758_), .ZN(new_n7774_));
  XOR2_X1    g06761(.A1(new_n7730_), .A2(new_n7742_), .Z(new_n7775_));
  XOR2_X1    g06762(.A1(new_n7751_), .A2(new_n7764_), .Z(new_n7776_));
  NOR4_X1    g06763(.A1(new_n7774_), .A2(new_n7773_), .A3(new_n7775_), .A4(new_n7776_), .ZN(new_n7777_));
  NAND2_X1   g06764(.A1(new_n7772_), .A2(new_n7777_), .ZN(new_n7778_));
  INV_X1     g06765(.I(new_n7778_), .ZN(new_n7779_));
  NAND3_X1   g06766(.A1(new_n7773_), .A2(new_n7745_), .A3(new_n7738_), .ZN(new_n7780_));
  NAND2_X1   g06767(.A1(new_n7730_), .A2(new_n7742_), .ZN(new_n7781_));
  NAND2_X1   g06768(.A1(new_n7780_), .A2(new_n7781_), .ZN(new_n7782_));
  NAND3_X1   g06769(.A1(new_n7774_), .A2(new_n7767_), .A3(new_n7761_), .ZN(new_n7783_));
  NAND2_X1   g06770(.A1(new_n7751_), .A2(new_n7764_), .ZN(new_n7784_));
  NAND2_X1   g06771(.A1(new_n7783_), .A2(new_n7784_), .ZN(new_n7785_));
  NOR3_X1    g06772(.A1(new_n7779_), .A2(new_n7782_), .A3(new_n7785_), .ZN(new_n7786_));
  INV_X1     g06773(.I(new_n7786_), .ZN(new_n7787_));
  INV_X1     g06774(.I(new_n7782_), .ZN(new_n7788_));
  INV_X1     g06775(.I(new_n7785_), .ZN(new_n7789_));
  NOR2_X1    g06776(.A1(new_n7789_), .A2(new_n7788_), .ZN(new_n7790_));
  INV_X1     g06777(.I(new_n7790_), .ZN(new_n7791_));
  INV_X1     g06778(.I(\A[910] ), .ZN(new_n7792_));
  NOR2_X1    g06779(.A1(\A[911] ), .A2(\A[912] ), .ZN(new_n7793_));
  NAND2_X1   g06780(.A1(\A[911] ), .A2(\A[912] ), .ZN(new_n7794_));
  AOI21_X1   g06781(.A1(new_n7792_), .A2(new_n7794_), .B(new_n7793_), .ZN(new_n7795_));
  INV_X1     g06782(.I(new_n7795_), .ZN(new_n7796_));
  INV_X1     g06783(.I(\A[907] ), .ZN(new_n7797_));
  NOR2_X1    g06784(.A1(\A[908] ), .A2(\A[909] ), .ZN(new_n7798_));
  NAND2_X1   g06785(.A1(\A[908] ), .A2(\A[909] ), .ZN(new_n7799_));
  AOI21_X1   g06786(.A1(new_n7797_), .A2(new_n7799_), .B(new_n7798_), .ZN(new_n7800_));
  INV_X1     g06787(.I(\A[909] ), .ZN(new_n7801_));
  NOR2_X1    g06788(.A1(new_n7801_), .A2(\A[908] ), .ZN(new_n7802_));
  INV_X1     g06789(.I(\A[908] ), .ZN(new_n7803_));
  NOR2_X1    g06790(.A1(new_n7803_), .A2(\A[909] ), .ZN(new_n7804_));
  OAI21_X1   g06791(.A1(new_n7802_), .A2(new_n7804_), .B(\A[907] ), .ZN(new_n7805_));
  INV_X1     g06792(.I(new_n7799_), .ZN(new_n7806_));
  OAI21_X1   g06793(.A1(new_n7806_), .A2(new_n7798_), .B(new_n7797_), .ZN(new_n7807_));
  INV_X1     g06794(.I(\A[912] ), .ZN(new_n7808_));
  NOR2_X1    g06795(.A1(new_n7808_), .A2(\A[911] ), .ZN(new_n7809_));
  INV_X1     g06796(.I(\A[911] ), .ZN(new_n7810_));
  NOR2_X1    g06797(.A1(new_n7810_), .A2(\A[912] ), .ZN(new_n7811_));
  OAI21_X1   g06798(.A1(new_n7809_), .A2(new_n7811_), .B(\A[910] ), .ZN(new_n7812_));
  INV_X1     g06799(.I(new_n7794_), .ZN(new_n7813_));
  OAI21_X1   g06800(.A1(new_n7813_), .A2(new_n7793_), .B(new_n7792_), .ZN(new_n7814_));
  NAND4_X1   g06801(.A1(new_n7805_), .A2(new_n7807_), .A3(new_n7812_), .A4(new_n7814_), .ZN(new_n7815_));
  NAND2_X1   g06802(.A1(new_n7815_), .A2(new_n7800_), .ZN(new_n7816_));
  INV_X1     g06803(.I(new_n7800_), .ZN(new_n7817_));
  NAND2_X1   g06804(.A1(new_n7803_), .A2(\A[909] ), .ZN(new_n7818_));
  NAND2_X1   g06805(.A1(new_n7801_), .A2(\A[908] ), .ZN(new_n7819_));
  AOI21_X1   g06806(.A1(new_n7818_), .A2(new_n7819_), .B(new_n7797_), .ZN(new_n7820_));
  INV_X1     g06807(.I(new_n7798_), .ZN(new_n7821_));
  AOI21_X1   g06808(.A1(new_n7821_), .A2(new_n7799_), .B(\A[907] ), .ZN(new_n7822_));
  NAND2_X1   g06809(.A1(new_n7810_), .A2(\A[912] ), .ZN(new_n7823_));
  NAND2_X1   g06810(.A1(new_n7808_), .A2(\A[911] ), .ZN(new_n7824_));
  AOI21_X1   g06811(.A1(new_n7823_), .A2(new_n7824_), .B(new_n7792_), .ZN(new_n7825_));
  INV_X1     g06812(.I(new_n7793_), .ZN(new_n7826_));
  AOI21_X1   g06813(.A1(new_n7826_), .A2(new_n7794_), .B(\A[910] ), .ZN(new_n7827_));
  NOR4_X1    g06814(.A1(new_n7820_), .A2(new_n7822_), .A3(new_n7827_), .A4(new_n7825_), .ZN(new_n7828_));
  NAND2_X1   g06815(.A1(new_n7828_), .A2(new_n7817_), .ZN(new_n7829_));
  AOI21_X1   g06816(.A1(new_n7829_), .A2(new_n7816_), .B(new_n7796_), .ZN(new_n7830_));
  NOR2_X1    g06817(.A1(new_n7828_), .A2(new_n7817_), .ZN(new_n7831_));
  NOR2_X1    g06818(.A1(new_n7815_), .A2(new_n7800_), .ZN(new_n7832_));
  NOR3_X1    g06819(.A1(new_n7831_), .A2(new_n7832_), .A3(new_n7795_), .ZN(new_n7833_));
  NOR2_X1    g06820(.A1(new_n7830_), .A2(new_n7833_), .ZN(new_n7834_));
  INV_X1     g06821(.I(\A[916] ), .ZN(new_n7835_));
  NOR2_X1    g06822(.A1(\A[917] ), .A2(\A[918] ), .ZN(new_n7836_));
  NAND2_X1   g06823(.A1(\A[917] ), .A2(\A[918] ), .ZN(new_n7837_));
  AOI21_X1   g06824(.A1(new_n7835_), .A2(new_n7837_), .B(new_n7836_), .ZN(new_n7838_));
  INV_X1     g06825(.I(\A[913] ), .ZN(new_n7839_));
  NOR2_X1    g06826(.A1(\A[914] ), .A2(\A[915] ), .ZN(new_n7840_));
  NAND2_X1   g06827(.A1(\A[914] ), .A2(\A[915] ), .ZN(new_n7841_));
  AOI21_X1   g06828(.A1(new_n7839_), .A2(new_n7841_), .B(new_n7840_), .ZN(new_n7842_));
  NAND2_X1   g06829(.A1(new_n7838_), .A2(new_n7842_), .ZN(new_n7843_));
  INV_X1     g06830(.I(\A[914] ), .ZN(new_n7844_));
  NAND2_X1   g06831(.A1(new_n7844_), .A2(\A[915] ), .ZN(new_n7845_));
  INV_X1     g06832(.I(\A[915] ), .ZN(new_n7846_));
  NAND2_X1   g06833(.A1(new_n7846_), .A2(\A[914] ), .ZN(new_n7847_));
  AOI21_X1   g06834(.A1(new_n7845_), .A2(new_n7847_), .B(new_n7839_), .ZN(new_n7848_));
  INV_X1     g06835(.I(new_n7840_), .ZN(new_n7849_));
  AOI21_X1   g06836(.A1(new_n7849_), .A2(new_n7841_), .B(\A[913] ), .ZN(new_n7850_));
  NOR2_X1    g06837(.A1(new_n7850_), .A2(new_n7848_), .ZN(new_n7851_));
  INV_X1     g06838(.I(\A[918] ), .ZN(new_n7852_));
  NOR2_X1    g06839(.A1(new_n7852_), .A2(\A[917] ), .ZN(new_n7853_));
  INV_X1     g06840(.I(\A[917] ), .ZN(new_n7854_));
  NOR2_X1    g06841(.A1(new_n7854_), .A2(\A[918] ), .ZN(new_n7855_));
  OAI21_X1   g06842(.A1(new_n7853_), .A2(new_n7855_), .B(\A[916] ), .ZN(new_n7856_));
  INV_X1     g06843(.I(new_n7837_), .ZN(new_n7857_));
  OAI21_X1   g06844(.A1(new_n7857_), .A2(new_n7836_), .B(new_n7835_), .ZN(new_n7858_));
  NAND2_X1   g06845(.A1(new_n7856_), .A2(new_n7858_), .ZN(new_n7859_));
  NAND2_X1   g06846(.A1(new_n7851_), .A2(new_n7859_), .ZN(new_n7860_));
  NOR2_X1    g06847(.A1(new_n7846_), .A2(\A[914] ), .ZN(new_n7861_));
  NOR2_X1    g06848(.A1(new_n7844_), .A2(\A[915] ), .ZN(new_n7862_));
  OAI21_X1   g06849(.A1(new_n7861_), .A2(new_n7862_), .B(\A[913] ), .ZN(new_n7863_));
  INV_X1     g06850(.I(new_n7841_), .ZN(new_n7864_));
  OAI21_X1   g06851(.A1(new_n7864_), .A2(new_n7840_), .B(new_n7839_), .ZN(new_n7865_));
  NAND2_X1   g06852(.A1(new_n7863_), .A2(new_n7865_), .ZN(new_n7866_));
  NAND2_X1   g06853(.A1(new_n7854_), .A2(\A[918] ), .ZN(new_n7867_));
  NAND2_X1   g06854(.A1(new_n7852_), .A2(\A[917] ), .ZN(new_n7868_));
  AOI21_X1   g06855(.A1(new_n7867_), .A2(new_n7868_), .B(new_n7835_), .ZN(new_n7869_));
  INV_X1     g06856(.I(new_n7836_), .ZN(new_n7870_));
  AOI21_X1   g06857(.A1(new_n7870_), .A2(new_n7837_), .B(\A[916] ), .ZN(new_n7871_));
  NOR2_X1    g06858(.A1(new_n7871_), .A2(new_n7869_), .ZN(new_n7872_));
  NAND2_X1   g06859(.A1(new_n7872_), .A2(new_n7866_), .ZN(new_n7873_));
  AOI21_X1   g06860(.A1(new_n7860_), .A2(new_n7873_), .B(new_n7843_), .ZN(new_n7874_));
  INV_X1     g06861(.I(new_n7838_), .ZN(new_n7875_));
  NAND4_X1   g06862(.A1(new_n7863_), .A2(new_n7865_), .A3(new_n7856_), .A4(new_n7858_), .ZN(new_n7876_));
  NAND2_X1   g06863(.A1(new_n7876_), .A2(new_n7842_), .ZN(new_n7877_));
  INV_X1     g06864(.I(new_n7842_), .ZN(new_n7878_));
  NAND3_X1   g06865(.A1(new_n7851_), .A2(new_n7872_), .A3(new_n7878_), .ZN(new_n7879_));
  AOI21_X1   g06866(.A1(new_n7877_), .A2(new_n7879_), .B(new_n7875_), .ZN(new_n7880_));
  AOI21_X1   g06867(.A1(new_n7851_), .A2(new_n7872_), .B(new_n7878_), .ZN(new_n7881_));
  NOR3_X1    g06868(.A1(new_n7866_), .A2(new_n7859_), .A3(new_n7842_), .ZN(new_n7882_));
  NOR3_X1    g06869(.A1(new_n7881_), .A2(new_n7882_), .A3(new_n7838_), .ZN(new_n7883_));
  NOR2_X1    g06870(.A1(new_n7876_), .A2(new_n7843_), .ZN(new_n7884_));
  NOR4_X1    g06871(.A1(new_n7848_), .A2(new_n7850_), .A3(new_n7871_), .A4(new_n7869_), .ZN(new_n7885_));
  NOR2_X1    g06872(.A1(new_n7851_), .A2(new_n7872_), .ZN(new_n7886_));
  NOR2_X1    g06873(.A1(new_n7886_), .A2(new_n7885_), .ZN(new_n7887_));
  AOI22_X1   g06874(.A1(new_n7805_), .A2(new_n7807_), .B1(new_n7812_), .B2(new_n7814_), .ZN(new_n7888_));
  NOR2_X1    g06875(.A1(new_n7888_), .A2(new_n7828_), .ZN(new_n7889_));
  NAND2_X1   g06876(.A1(new_n7795_), .A2(new_n7800_), .ZN(new_n7890_));
  NOR2_X1    g06877(.A1(new_n7815_), .A2(new_n7890_), .ZN(new_n7891_));
  NAND4_X1   g06878(.A1(new_n7887_), .A2(new_n7889_), .A3(new_n7884_), .A4(new_n7891_), .ZN(new_n7892_));
  NOR4_X1    g06879(.A1(new_n7892_), .A2(new_n7874_), .A3(new_n7880_), .A4(new_n7883_), .ZN(new_n7893_));
  NOR3_X1    g06880(.A1(new_n7880_), .A2(new_n7883_), .A3(new_n7874_), .ZN(new_n7894_));
  INV_X1     g06881(.I(new_n7843_), .ZN(new_n7895_));
  NAND2_X1   g06882(.A1(new_n7885_), .A2(new_n7895_), .ZN(new_n7896_));
  NAND2_X1   g06883(.A1(new_n7866_), .A2(new_n7859_), .ZN(new_n7897_));
  NAND2_X1   g06884(.A1(new_n7897_), .A2(new_n7876_), .ZN(new_n7898_));
  OAI22_X1   g06885(.A1(new_n7820_), .A2(new_n7822_), .B1(new_n7827_), .B2(new_n7825_), .ZN(new_n7899_));
  NAND2_X1   g06886(.A1(new_n7899_), .A2(new_n7815_), .ZN(new_n7900_));
  NAND3_X1   g06887(.A1(new_n7828_), .A2(new_n7795_), .A3(new_n7800_), .ZN(new_n7901_));
  NOR4_X1    g06888(.A1(new_n7898_), .A2(new_n7896_), .A3(new_n7901_), .A4(new_n7900_), .ZN(new_n7902_));
  NOR2_X1    g06889(.A1(new_n7894_), .A2(new_n7902_), .ZN(new_n7903_));
  OAI21_X1   g06890(.A1(new_n7903_), .A2(new_n7893_), .B(new_n7834_), .ZN(new_n7904_));
  OAI21_X1   g06891(.A1(new_n7881_), .A2(new_n7882_), .B(new_n7838_), .ZN(new_n7905_));
  NAND3_X1   g06892(.A1(new_n7877_), .A2(new_n7879_), .A3(new_n7875_), .ZN(new_n7906_));
  NAND2_X1   g06893(.A1(new_n7905_), .A2(new_n7906_), .ZN(new_n7907_));
  OAI21_X1   g06894(.A1(new_n7907_), .A2(new_n7874_), .B(new_n7902_), .ZN(new_n7908_));
  NAND3_X1   g06895(.A1(new_n7887_), .A2(new_n7884_), .A3(new_n7889_), .ZN(new_n7909_));
  NOR2_X1    g06896(.A1(new_n7874_), .A2(new_n7901_), .ZN(new_n7910_));
  OAI21_X1   g06897(.A1(new_n7907_), .A2(new_n7909_), .B(new_n7910_), .ZN(new_n7911_));
  NAND3_X1   g06898(.A1(new_n7911_), .A2(new_n7908_), .A3(new_n7834_), .ZN(new_n7912_));
  NAND2_X1   g06899(.A1(new_n7912_), .A2(new_n7904_), .ZN(new_n7913_));
  INV_X1     g06900(.I(new_n7834_), .ZN(new_n7914_));
  NAND2_X1   g06901(.A1(new_n7894_), .A2(new_n7902_), .ZN(new_n7915_));
  OAI21_X1   g06902(.A1(new_n7907_), .A2(new_n7874_), .B(new_n7892_), .ZN(new_n7916_));
  AOI21_X1   g06903(.A1(new_n7916_), .A2(new_n7915_), .B(new_n7914_), .ZN(new_n7917_));
  NOR2_X1    g06904(.A1(new_n7894_), .A2(new_n7892_), .ZN(new_n7918_));
  NOR2_X1    g06905(.A1(new_n7880_), .A2(new_n7883_), .ZN(new_n7919_));
  NOR3_X1    g06906(.A1(new_n7898_), .A2(new_n7900_), .A3(new_n7896_), .ZN(new_n7920_));
  NOR2_X1    g06907(.A1(new_n7872_), .A2(new_n7866_), .ZN(new_n7921_));
  NOR2_X1    g06908(.A1(new_n7851_), .A2(new_n7859_), .ZN(new_n7922_));
  OAI21_X1   g06909(.A1(new_n7921_), .A2(new_n7922_), .B(new_n7895_), .ZN(new_n7923_));
  NAND2_X1   g06910(.A1(new_n7923_), .A2(new_n7891_), .ZN(new_n7924_));
  AOI21_X1   g06911(.A1(new_n7919_), .A2(new_n7920_), .B(new_n7924_), .ZN(new_n7925_));
  NOR3_X1    g06912(.A1(new_n7925_), .A2(new_n7918_), .A3(new_n7914_), .ZN(new_n7926_));
  NOR2_X1    g06913(.A1(new_n7898_), .A2(new_n7896_), .ZN(new_n7927_));
  NAND2_X1   g06914(.A1(new_n7889_), .A2(new_n7891_), .ZN(new_n7928_));
  NOR2_X1    g06915(.A1(new_n7927_), .A2(new_n7928_), .ZN(new_n7929_));
  NAND2_X1   g06916(.A1(new_n7887_), .A2(new_n7884_), .ZN(new_n7930_));
  NOR2_X1    g06917(.A1(new_n7901_), .A2(new_n7900_), .ZN(new_n7931_));
  NOR2_X1    g06918(.A1(new_n7930_), .A2(new_n7931_), .ZN(new_n7932_));
  NOR2_X1    g06919(.A1(new_n7932_), .A2(new_n7929_), .ZN(new_n7933_));
  INV_X1     g06920(.I(\A[903] ), .ZN(new_n7934_));
  NOR2_X1    g06921(.A1(new_n7934_), .A2(\A[902] ), .ZN(new_n7935_));
  INV_X1     g06922(.I(\A[902] ), .ZN(new_n7936_));
  NOR2_X1    g06923(.A1(new_n7936_), .A2(\A[903] ), .ZN(new_n7937_));
  OAI21_X1   g06924(.A1(new_n7935_), .A2(new_n7937_), .B(\A[901] ), .ZN(new_n7938_));
  INV_X1     g06925(.I(\A[901] ), .ZN(new_n7939_));
  NOR2_X1    g06926(.A1(\A[902] ), .A2(\A[903] ), .ZN(new_n7940_));
  NAND2_X1   g06927(.A1(\A[902] ), .A2(\A[903] ), .ZN(new_n7941_));
  INV_X1     g06928(.I(new_n7941_), .ZN(new_n7942_));
  OAI21_X1   g06929(.A1(new_n7942_), .A2(new_n7940_), .B(new_n7939_), .ZN(new_n7943_));
  NAND2_X1   g06930(.A1(new_n7938_), .A2(new_n7943_), .ZN(new_n7944_));
  INV_X1     g06931(.I(\A[906] ), .ZN(new_n7945_));
  NOR2_X1    g06932(.A1(new_n7945_), .A2(\A[905] ), .ZN(new_n7946_));
  INV_X1     g06933(.I(\A[905] ), .ZN(new_n7947_));
  NOR2_X1    g06934(.A1(new_n7947_), .A2(\A[906] ), .ZN(new_n7948_));
  OAI21_X1   g06935(.A1(new_n7946_), .A2(new_n7948_), .B(\A[904] ), .ZN(new_n7949_));
  INV_X1     g06936(.I(\A[904] ), .ZN(new_n7950_));
  NOR2_X1    g06937(.A1(\A[905] ), .A2(\A[906] ), .ZN(new_n7951_));
  NAND2_X1   g06938(.A1(\A[905] ), .A2(\A[906] ), .ZN(new_n7952_));
  INV_X1     g06939(.I(new_n7952_), .ZN(new_n7953_));
  OAI21_X1   g06940(.A1(new_n7953_), .A2(new_n7951_), .B(new_n7950_), .ZN(new_n7954_));
  NAND2_X1   g06941(.A1(new_n7949_), .A2(new_n7954_), .ZN(new_n7955_));
  AOI21_X1   g06942(.A1(new_n7950_), .A2(new_n7952_), .B(new_n7951_), .ZN(new_n7956_));
  AOI21_X1   g06943(.A1(new_n7939_), .A2(new_n7941_), .B(new_n7940_), .ZN(new_n7957_));
  NAND2_X1   g06944(.A1(new_n7956_), .A2(new_n7957_), .ZN(new_n7958_));
  NOR3_X1    g06945(.A1(new_n7944_), .A2(new_n7955_), .A3(new_n7958_), .ZN(new_n7959_));
  NOR2_X1    g06946(.A1(new_n7944_), .A2(new_n7955_), .ZN(new_n7960_));
  NAND2_X1   g06947(.A1(new_n7936_), .A2(\A[903] ), .ZN(new_n7961_));
  NAND2_X1   g06948(.A1(new_n7934_), .A2(\A[902] ), .ZN(new_n7962_));
  AOI21_X1   g06949(.A1(new_n7961_), .A2(new_n7962_), .B(new_n7939_), .ZN(new_n7963_));
  INV_X1     g06950(.I(new_n7940_), .ZN(new_n7964_));
  AOI21_X1   g06951(.A1(new_n7964_), .A2(new_n7941_), .B(\A[901] ), .ZN(new_n7965_));
  NOR2_X1    g06952(.A1(new_n7965_), .A2(new_n7963_), .ZN(new_n7966_));
  NAND2_X1   g06953(.A1(new_n7947_), .A2(\A[906] ), .ZN(new_n7967_));
  NAND2_X1   g06954(.A1(new_n7945_), .A2(\A[905] ), .ZN(new_n7968_));
  AOI21_X1   g06955(.A1(new_n7967_), .A2(new_n7968_), .B(new_n7950_), .ZN(new_n7969_));
  INV_X1     g06956(.I(new_n7951_), .ZN(new_n7970_));
  AOI21_X1   g06957(.A1(new_n7970_), .A2(new_n7952_), .B(\A[904] ), .ZN(new_n7971_));
  NOR2_X1    g06958(.A1(new_n7971_), .A2(new_n7969_), .ZN(new_n7972_));
  NOR2_X1    g06959(.A1(new_n7966_), .A2(new_n7972_), .ZN(new_n7973_));
  NOR2_X1    g06960(.A1(new_n7973_), .A2(new_n7960_), .ZN(new_n7974_));
  INV_X1     g06961(.I(\A[895] ), .ZN(new_n7975_));
  INV_X1     g06962(.I(\A[896] ), .ZN(new_n7976_));
  NAND2_X1   g06963(.A1(new_n7976_), .A2(\A[897] ), .ZN(new_n7977_));
  INV_X1     g06964(.I(\A[897] ), .ZN(new_n7978_));
  NAND2_X1   g06965(.A1(new_n7978_), .A2(\A[896] ), .ZN(new_n7979_));
  AOI21_X1   g06966(.A1(new_n7977_), .A2(new_n7979_), .B(new_n7975_), .ZN(new_n7980_));
  NOR2_X1    g06967(.A1(\A[896] ), .A2(\A[897] ), .ZN(new_n7981_));
  INV_X1     g06968(.I(new_n7981_), .ZN(new_n7982_));
  NAND2_X1   g06969(.A1(\A[896] ), .A2(\A[897] ), .ZN(new_n7983_));
  AOI21_X1   g06970(.A1(new_n7982_), .A2(new_n7983_), .B(\A[895] ), .ZN(new_n7984_));
  NOR2_X1    g06971(.A1(new_n7984_), .A2(new_n7980_), .ZN(new_n7985_));
  INV_X1     g06972(.I(\A[898] ), .ZN(new_n7986_));
  INV_X1     g06973(.I(\A[899] ), .ZN(new_n7987_));
  NAND2_X1   g06974(.A1(new_n7987_), .A2(\A[900] ), .ZN(new_n7988_));
  INV_X1     g06975(.I(\A[900] ), .ZN(new_n7989_));
  NAND2_X1   g06976(.A1(new_n7989_), .A2(\A[899] ), .ZN(new_n7990_));
  AOI21_X1   g06977(.A1(new_n7988_), .A2(new_n7990_), .B(new_n7986_), .ZN(new_n7991_));
  NOR2_X1    g06978(.A1(\A[899] ), .A2(\A[900] ), .ZN(new_n7992_));
  INV_X1     g06979(.I(new_n7992_), .ZN(new_n7993_));
  NAND2_X1   g06980(.A1(\A[899] ), .A2(\A[900] ), .ZN(new_n7994_));
  AOI21_X1   g06981(.A1(new_n7993_), .A2(new_n7994_), .B(\A[898] ), .ZN(new_n7995_));
  NOR2_X1    g06982(.A1(new_n7995_), .A2(new_n7991_), .ZN(new_n7996_));
  AOI21_X1   g06983(.A1(new_n7986_), .A2(new_n7994_), .B(new_n7992_), .ZN(new_n7997_));
  AOI21_X1   g06984(.A1(new_n7975_), .A2(new_n7983_), .B(new_n7981_), .ZN(new_n7998_));
  NAND2_X1   g06985(.A1(new_n7997_), .A2(new_n7998_), .ZN(new_n7999_));
  NAND2_X1   g06986(.A1(new_n7974_), .A2(new_n7959_), .ZN(new_n8001_));
  NAND2_X1   g06987(.A1(new_n7933_), .A2(new_n8001_), .ZN(new_n8002_));
  OAI21_X1   g06988(.A1(new_n7917_), .A2(new_n7926_), .B(new_n8002_), .ZN(new_n8003_));
  AND2_X2    g06989(.A1(new_n7974_), .A2(new_n7959_), .Z(new_n8004_));
  NOR3_X1    g06990(.A1(new_n7929_), .A2(new_n7932_), .A3(new_n8004_), .ZN(new_n8005_));
  NAND3_X1   g06991(.A1(new_n7912_), .A2(new_n7904_), .A3(new_n8005_), .ZN(new_n8006_));
  NAND2_X1   g06992(.A1(new_n7966_), .A2(new_n7972_), .ZN(new_n8007_));
  NAND2_X1   g06993(.A1(new_n7944_), .A2(new_n7955_), .ZN(new_n8008_));
  NAND3_X1   g06994(.A1(new_n7959_), .A2(new_n8007_), .A3(new_n8008_), .ZN(new_n8009_));
  NAND2_X1   g06995(.A1(new_n7985_), .A2(new_n7996_), .ZN(new_n8010_));
  NOR2_X1    g06996(.A1(new_n7978_), .A2(\A[896] ), .ZN(new_n8011_));
  NOR2_X1    g06997(.A1(new_n7976_), .A2(\A[897] ), .ZN(new_n8012_));
  OAI21_X1   g06998(.A1(new_n8011_), .A2(new_n8012_), .B(\A[895] ), .ZN(new_n8013_));
  INV_X1     g06999(.I(new_n7983_), .ZN(new_n8014_));
  OAI21_X1   g07000(.A1(new_n8014_), .A2(new_n7981_), .B(new_n7975_), .ZN(new_n8015_));
  NAND2_X1   g07001(.A1(new_n8013_), .A2(new_n8015_), .ZN(new_n8016_));
  NOR2_X1    g07002(.A1(new_n7989_), .A2(\A[899] ), .ZN(new_n8017_));
  NOR2_X1    g07003(.A1(new_n7987_), .A2(\A[900] ), .ZN(new_n8018_));
  OAI21_X1   g07004(.A1(new_n8017_), .A2(new_n8018_), .B(\A[898] ), .ZN(new_n8019_));
  INV_X1     g07005(.I(new_n7994_), .ZN(new_n8020_));
  OAI21_X1   g07006(.A1(new_n8020_), .A2(new_n7992_), .B(new_n7986_), .ZN(new_n8021_));
  NAND2_X1   g07007(.A1(new_n8019_), .A2(new_n8021_), .ZN(new_n8022_));
  NAND2_X1   g07008(.A1(new_n8016_), .A2(new_n8022_), .ZN(new_n8023_));
  NAND2_X1   g07009(.A1(new_n8010_), .A2(new_n8023_), .ZN(new_n8024_));
  INV_X1     g07010(.I(new_n7956_), .ZN(new_n8025_));
  OAI21_X1   g07011(.A1(new_n7944_), .A2(new_n7955_), .B(new_n7957_), .ZN(new_n8026_));
  INV_X1     g07012(.I(new_n7957_), .ZN(new_n8027_));
  NAND3_X1   g07013(.A1(new_n7966_), .A2(new_n7972_), .A3(new_n8027_), .ZN(new_n8028_));
  AOI21_X1   g07014(.A1(new_n8026_), .A2(new_n8028_), .B(new_n8025_), .ZN(new_n8029_));
  AOI21_X1   g07015(.A1(new_n7966_), .A2(new_n7972_), .B(new_n8027_), .ZN(new_n8030_));
  NOR3_X1    g07016(.A1(new_n7944_), .A2(new_n7955_), .A3(new_n7957_), .ZN(new_n8031_));
  NOR3_X1    g07017(.A1(new_n8030_), .A2(new_n8031_), .A3(new_n7956_), .ZN(new_n8032_));
  NOR4_X1    g07018(.A1(new_n8029_), .A2(new_n8032_), .A3(new_n8009_), .A4(new_n8024_), .ZN(new_n8033_));
  NOR3_X1    g07019(.A1(new_n8016_), .A2(new_n8022_), .A3(new_n7999_), .ZN(new_n8034_));
  INV_X1     g07020(.I(new_n7958_), .ZN(new_n8035_));
  NOR2_X1    g07021(.A1(new_n7972_), .A2(new_n7944_), .ZN(new_n8036_));
  NOR2_X1    g07022(.A1(new_n7966_), .A2(new_n7955_), .ZN(new_n8037_));
  OAI21_X1   g07023(.A1(new_n8036_), .A2(new_n8037_), .B(new_n8035_), .ZN(new_n8038_));
  NAND2_X1   g07024(.A1(new_n8038_), .A2(new_n8034_), .ZN(new_n8039_));
  NOR2_X1    g07025(.A1(new_n8033_), .A2(new_n8039_), .ZN(new_n8040_));
  NOR4_X1    g07026(.A1(new_n7980_), .A2(new_n7984_), .A3(new_n7995_), .A4(new_n7991_), .ZN(new_n8041_));
  INV_X1     g07027(.I(new_n7998_), .ZN(new_n8042_));
  NOR2_X1    g07028(.A1(new_n8041_), .A2(new_n8042_), .ZN(new_n8043_));
  NOR3_X1    g07029(.A1(new_n8016_), .A2(new_n8022_), .A3(new_n7998_), .ZN(new_n8044_));
  OAI21_X1   g07030(.A1(new_n8043_), .A2(new_n8044_), .B(new_n7997_), .ZN(new_n8045_));
  INV_X1     g07031(.I(new_n7997_), .ZN(new_n8046_));
  OAI21_X1   g07032(.A1(new_n8016_), .A2(new_n8022_), .B(new_n7998_), .ZN(new_n8047_));
  NAND3_X1   g07033(.A1(new_n7985_), .A2(new_n7996_), .A3(new_n8042_), .ZN(new_n8048_));
  NAND3_X1   g07034(.A1(new_n8047_), .A2(new_n8048_), .A3(new_n8046_), .ZN(new_n8049_));
  NAND2_X1   g07035(.A1(new_n8045_), .A2(new_n8049_), .ZN(new_n8050_));
  NAND2_X1   g07036(.A1(new_n8040_), .A2(new_n8050_), .ZN(new_n8051_));
  NOR2_X1    g07037(.A1(new_n7985_), .A2(new_n7996_), .ZN(new_n8052_));
  NOR2_X1    g07038(.A1(new_n8052_), .A2(new_n8041_), .ZN(new_n8053_));
  NAND4_X1   g07039(.A1(new_n7974_), .A2(new_n8053_), .A3(new_n7959_), .A4(new_n8034_), .ZN(new_n8054_));
  NAND2_X1   g07040(.A1(new_n8050_), .A2(new_n8054_), .ZN(new_n8055_));
  AOI21_X1   g07041(.A1(new_n8047_), .A2(new_n8048_), .B(new_n8046_), .ZN(new_n8056_));
  NOR3_X1    g07042(.A1(new_n8043_), .A2(new_n8044_), .A3(new_n7997_), .ZN(new_n8057_));
  NOR2_X1    g07043(.A1(new_n8057_), .A2(new_n8056_), .ZN(new_n8058_));
  NAND3_X1   g07044(.A1(new_n8034_), .A2(new_n8010_), .A3(new_n8023_), .ZN(new_n8059_));
  NOR2_X1    g07045(.A1(new_n8009_), .A2(new_n8059_), .ZN(new_n8060_));
  NAND2_X1   g07046(.A1(new_n7966_), .A2(new_n7955_), .ZN(new_n8061_));
  NAND2_X1   g07047(.A1(new_n7972_), .A2(new_n7944_), .ZN(new_n8062_));
  AOI21_X1   g07048(.A1(new_n8061_), .A2(new_n8062_), .B(new_n7958_), .ZN(new_n8063_));
  NOR3_X1    g07049(.A1(new_n8032_), .A2(new_n8029_), .A3(new_n8063_), .ZN(new_n8064_));
  AOI21_X1   g07050(.A1(new_n8058_), .A2(new_n8060_), .B(new_n8064_), .ZN(new_n8065_));
  OAI21_X1   g07051(.A1(new_n8030_), .A2(new_n8031_), .B(new_n7956_), .ZN(new_n8066_));
  NAND3_X1   g07052(.A1(new_n8026_), .A2(new_n8028_), .A3(new_n8025_), .ZN(new_n8067_));
  NAND3_X1   g07053(.A1(new_n8066_), .A2(new_n8067_), .A3(new_n8038_), .ZN(new_n8068_));
  NOR3_X1    g07054(.A1(new_n8068_), .A2(new_n8050_), .A3(new_n8054_), .ZN(new_n8069_));
  OAI21_X1   g07055(.A1(new_n8065_), .A2(new_n8069_), .B(new_n8055_), .ZN(new_n8070_));
  NAND2_X1   g07056(.A1(new_n8070_), .A2(new_n8051_), .ZN(new_n8071_));
  AOI22_X1   g07057(.A1(new_n8003_), .A2(new_n8006_), .B1(new_n8071_), .B2(new_n7913_), .ZN(new_n8072_));
  NOR2_X1    g07058(.A1(new_n7918_), .A2(new_n7834_), .ZN(new_n8073_));
  NOR2_X1    g07059(.A1(new_n7838_), .A2(new_n7842_), .ZN(new_n8074_));
  OAI21_X1   g07060(.A1(new_n7876_), .A2(new_n8074_), .B(new_n7843_), .ZN(new_n8075_));
  NOR2_X1    g07061(.A1(new_n7795_), .A2(new_n7800_), .ZN(new_n8076_));
  OAI21_X1   g07062(.A1(new_n7815_), .A2(new_n8076_), .B(new_n7890_), .ZN(new_n8077_));
  XNOR2_X1   g07063(.A1(new_n8075_), .A2(new_n8077_), .ZN(new_n8078_));
  INV_X1     g07064(.I(new_n8078_), .ZN(new_n8079_));
  NOR3_X1    g07065(.A1(new_n8073_), .A2(new_n7925_), .A3(new_n8079_), .ZN(new_n8080_));
  AOI21_X1   g07066(.A1(new_n8068_), .A2(new_n8060_), .B(new_n8058_), .ZN(new_n8081_));
  NAND2_X1   g07067(.A1(new_n8025_), .A2(new_n8027_), .ZN(new_n8082_));
  AOI21_X1   g07068(.A1(new_n7960_), .A2(new_n8082_), .B(new_n8035_), .ZN(new_n8083_));
  NOR2_X1    g07069(.A1(new_n7997_), .A2(new_n7998_), .ZN(new_n8084_));
  OAI21_X1   g07070(.A1(new_n8010_), .A2(new_n8084_), .B(new_n7999_), .ZN(new_n8085_));
  XNOR2_X1   g07071(.A1(new_n8083_), .A2(new_n8085_), .ZN(new_n8086_));
  NOR3_X1    g07072(.A1(new_n8081_), .A2(new_n8040_), .A3(new_n8086_), .ZN(new_n8087_));
  XOR2_X1    g07073(.A1(new_n8080_), .A2(new_n8087_), .Z(new_n8088_));
  NAND2_X1   g07074(.A1(new_n8088_), .A2(new_n8072_), .ZN(new_n8089_));
  NOR2_X1    g07075(.A1(new_n7917_), .A2(new_n7926_), .ZN(new_n8090_));
  AOI21_X1   g07076(.A1(new_n7912_), .A2(new_n7904_), .B(new_n8005_), .ZN(new_n8091_));
  NOR3_X1    g07077(.A1(new_n7917_), .A2(new_n7926_), .A3(new_n8002_), .ZN(new_n8092_));
  OAI21_X1   g07078(.A1(new_n8050_), .A2(new_n8054_), .B(new_n8068_), .ZN(new_n8093_));
  NAND3_X1   g07079(.A1(new_n8064_), .A2(new_n8058_), .A3(new_n8060_), .ZN(new_n8094_));
  NAND2_X1   g07080(.A1(new_n8093_), .A2(new_n8094_), .ZN(new_n8095_));
  AOI22_X1   g07081(.A1(new_n8095_), .A2(new_n8055_), .B1(new_n8040_), .B2(new_n8050_), .ZN(new_n8096_));
  OAI22_X1   g07082(.A1(new_n8090_), .A2(new_n8096_), .B1(new_n8092_), .B2(new_n8091_), .ZN(new_n8097_));
  NAND2_X1   g07083(.A1(new_n7908_), .A2(new_n7914_), .ZN(new_n8098_));
  NAND3_X1   g07084(.A1(new_n8098_), .A2(new_n8078_), .A3(new_n7911_), .ZN(new_n8099_));
  INV_X1     g07085(.I(new_n8087_), .ZN(new_n8100_));
  NAND2_X1   g07086(.A1(new_n8100_), .A2(new_n8099_), .ZN(new_n8101_));
  NAND2_X1   g07087(.A1(new_n8080_), .A2(new_n8087_), .ZN(new_n8102_));
  NAND2_X1   g07088(.A1(new_n8101_), .A2(new_n8102_), .ZN(new_n8103_));
  NAND2_X1   g07089(.A1(new_n8097_), .A2(new_n8103_), .ZN(new_n8104_));
  NAND2_X1   g07090(.A1(new_n8089_), .A2(new_n8104_), .ZN(new_n8105_));
  INV_X1     g07091(.I(\A[934] ), .ZN(new_n8106_));
  NOR2_X1    g07092(.A1(\A[935] ), .A2(\A[936] ), .ZN(new_n8107_));
  NAND2_X1   g07093(.A1(\A[935] ), .A2(\A[936] ), .ZN(new_n8108_));
  AOI21_X1   g07094(.A1(new_n8106_), .A2(new_n8108_), .B(new_n8107_), .ZN(new_n8109_));
  INV_X1     g07095(.I(new_n8109_), .ZN(new_n8110_));
  INV_X1     g07096(.I(\A[931] ), .ZN(new_n8111_));
  NOR2_X1    g07097(.A1(\A[932] ), .A2(\A[933] ), .ZN(new_n8112_));
  NAND2_X1   g07098(.A1(\A[932] ), .A2(\A[933] ), .ZN(new_n8113_));
  AOI21_X1   g07099(.A1(new_n8111_), .A2(new_n8113_), .B(new_n8112_), .ZN(new_n8114_));
  INV_X1     g07100(.I(\A[933] ), .ZN(new_n8115_));
  NOR2_X1    g07101(.A1(new_n8115_), .A2(\A[932] ), .ZN(new_n8116_));
  INV_X1     g07102(.I(\A[932] ), .ZN(new_n8117_));
  NOR2_X1    g07103(.A1(new_n8117_), .A2(\A[933] ), .ZN(new_n8118_));
  OAI21_X1   g07104(.A1(new_n8116_), .A2(new_n8118_), .B(\A[931] ), .ZN(new_n8119_));
  INV_X1     g07105(.I(new_n8113_), .ZN(new_n8120_));
  OAI21_X1   g07106(.A1(new_n8120_), .A2(new_n8112_), .B(new_n8111_), .ZN(new_n8121_));
  INV_X1     g07107(.I(\A[936] ), .ZN(new_n8122_));
  NOR2_X1    g07108(.A1(new_n8122_), .A2(\A[935] ), .ZN(new_n8123_));
  INV_X1     g07109(.I(\A[935] ), .ZN(new_n8124_));
  NOR2_X1    g07110(.A1(new_n8124_), .A2(\A[936] ), .ZN(new_n8125_));
  OAI21_X1   g07111(.A1(new_n8123_), .A2(new_n8125_), .B(\A[934] ), .ZN(new_n8126_));
  INV_X1     g07112(.I(new_n8108_), .ZN(new_n8127_));
  OAI21_X1   g07113(.A1(new_n8127_), .A2(new_n8107_), .B(new_n8106_), .ZN(new_n8128_));
  NAND4_X1   g07114(.A1(new_n8119_), .A2(new_n8121_), .A3(new_n8126_), .A4(new_n8128_), .ZN(new_n8129_));
  NAND2_X1   g07115(.A1(new_n8129_), .A2(new_n8114_), .ZN(new_n8130_));
  INV_X1     g07116(.I(new_n8114_), .ZN(new_n8131_));
  INV_X1     g07117(.I(new_n8116_), .ZN(new_n8132_));
  NAND2_X1   g07118(.A1(new_n8115_), .A2(\A[932] ), .ZN(new_n8133_));
  AOI21_X1   g07119(.A1(new_n8132_), .A2(new_n8133_), .B(new_n8111_), .ZN(new_n8134_));
  INV_X1     g07120(.I(new_n8112_), .ZN(new_n8135_));
  AOI21_X1   g07121(.A1(new_n8135_), .A2(new_n8113_), .B(\A[931] ), .ZN(new_n8136_));
  NAND2_X1   g07122(.A1(new_n8124_), .A2(\A[936] ), .ZN(new_n8137_));
  NAND2_X1   g07123(.A1(new_n8122_), .A2(\A[935] ), .ZN(new_n8138_));
  AOI21_X1   g07124(.A1(new_n8137_), .A2(new_n8138_), .B(new_n8106_), .ZN(new_n8139_));
  INV_X1     g07125(.I(new_n8107_), .ZN(new_n8140_));
  AOI21_X1   g07126(.A1(new_n8140_), .A2(new_n8108_), .B(\A[934] ), .ZN(new_n8141_));
  NOR4_X1    g07127(.A1(new_n8134_), .A2(new_n8136_), .A3(new_n8141_), .A4(new_n8139_), .ZN(new_n8142_));
  NAND2_X1   g07128(.A1(new_n8142_), .A2(new_n8131_), .ZN(new_n8143_));
  AOI21_X1   g07129(.A1(new_n8143_), .A2(new_n8130_), .B(new_n8110_), .ZN(new_n8144_));
  NOR2_X1    g07130(.A1(new_n8142_), .A2(new_n8131_), .ZN(new_n8145_));
  NOR2_X1    g07131(.A1(new_n8129_), .A2(new_n8114_), .ZN(new_n8146_));
  NOR3_X1    g07132(.A1(new_n8145_), .A2(new_n8146_), .A3(new_n8109_), .ZN(new_n8147_));
  NOR2_X1    g07133(.A1(new_n8147_), .A2(new_n8144_), .ZN(new_n8148_));
  INV_X1     g07134(.I(\A[940] ), .ZN(new_n8149_));
  NOR2_X1    g07135(.A1(\A[941] ), .A2(\A[942] ), .ZN(new_n8150_));
  NAND2_X1   g07136(.A1(\A[941] ), .A2(\A[942] ), .ZN(new_n8151_));
  AOI21_X1   g07137(.A1(new_n8149_), .A2(new_n8151_), .B(new_n8150_), .ZN(new_n8152_));
  INV_X1     g07138(.I(\A[937] ), .ZN(new_n8153_));
  NOR2_X1    g07139(.A1(\A[938] ), .A2(\A[939] ), .ZN(new_n8154_));
  NAND2_X1   g07140(.A1(\A[938] ), .A2(\A[939] ), .ZN(new_n8155_));
  AOI21_X1   g07141(.A1(new_n8153_), .A2(new_n8155_), .B(new_n8154_), .ZN(new_n8156_));
  NAND2_X1   g07142(.A1(new_n8152_), .A2(new_n8156_), .ZN(new_n8157_));
  INV_X1     g07143(.I(\A[938] ), .ZN(new_n8158_));
  NAND2_X1   g07144(.A1(new_n8158_), .A2(\A[939] ), .ZN(new_n8159_));
  INV_X1     g07145(.I(\A[939] ), .ZN(new_n8160_));
  NAND2_X1   g07146(.A1(new_n8160_), .A2(\A[938] ), .ZN(new_n8161_));
  AOI21_X1   g07147(.A1(new_n8159_), .A2(new_n8161_), .B(new_n8153_), .ZN(new_n8162_));
  INV_X1     g07148(.I(new_n8154_), .ZN(new_n8163_));
  AOI21_X1   g07149(.A1(new_n8163_), .A2(new_n8155_), .B(\A[937] ), .ZN(new_n8164_));
  NOR2_X1    g07150(.A1(new_n8164_), .A2(new_n8162_), .ZN(new_n8165_));
  INV_X1     g07151(.I(\A[942] ), .ZN(new_n8166_));
  NOR2_X1    g07152(.A1(new_n8166_), .A2(\A[941] ), .ZN(new_n8167_));
  INV_X1     g07153(.I(\A[941] ), .ZN(new_n8168_));
  NOR2_X1    g07154(.A1(new_n8168_), .A2(\A[942] ), .ZN(new_n8169_));
  OAI21_X1   g07155(.A1(new_n8167_), .A2(new_n8169_), .B(\A[940] ), .ZN(new_n8170_));
  AND2_X2    g07156(.A1(\A[941] ), .A2(\A[942] ), .Z(new_n8171_));
  OAI21_X1   g07157(.A1(new_n8171_), .A2(new_n8150_), .B(new_n8149_), .ZN(new_n8172_));
  NAND2_X1   g07158(.A1(new_n8170_), .A2(new_n8172_), .ZN(new_n8173_));
  NAND2_X1   g07159(.A1(new_n8165_), .A2(new_n8173_), .ZN(new_n8174_));
  NOR2_X1    g07160(.A1(new_n8160_), .A2(\A[938] ), .ZN(new_n8175_));
  NOR2_X1    g07161(.A1(new_n8158_), .A2(\A[939] ), .ZN(new_n8176_));
  OAI21_X1   g07162(.A1(new_n8175_), .A2(new_n8176_), .B(\A[937] ), .ZN(new_n8177_));
  INV_X1     g07163(.I(new_n8155_), .ZN(new_n8178_));
  OAI21_X1   g07164(.A1(new_n8178_), .A2(new_n8154_), .B(new_n8153_), .ZN(new_n8179_));
  NAND2_X1   g07165(.A1(new_n8177_), .A2(new_n8179_), .ZN(new_n8180_));
  NAND2_X1   g07166(.A1(new_n8168_), .A2(\A[942] ), .ZN(new_n8181_));
  NAND2_X1   g07167(.A1(new_n8166_), .A2(\A[941] ), .ZN(new_n8182_));
  AOI21_X1   g07168(.A1(new_n8181_), .A2(new_n8182_), .B(new_n8149_), .ZN(new_n8183_));
  INV_X1     g07169(.I(new_n8150_), .ZN(new_n8184_));
  AOI21_X1   g07170(.A1(new_n8184_), .A2(new_n8151_), .B(\A[940] ), .ZN(new_n8185_));
  NOR2_X1    g07171(.A1(new_n8185_), .A2(new_n8183_), .ZN(new_n8186_));
  NAND2_X1   g07172(.A1(new_n8186_), .A2(new_n8180_), .ZN(new_n8187_));
  AOI21_X1   g07173(.A1(new_n8187_), .A2(new_n8174_), .B(new_n8157_), .ZN(new_n8188_));
  INV_X1     g07174(.I(new_n8152_), .ZN(new_n8189_));
  NAND4_X1   g07175(.A1(new_n8177_), .A2(new_n8170_), .A3(new_n8179_), .A4(new_n8172_), .ZN(new_n8190_));
  NAND2_X1   g07176(.A1(new_n8190_), .A2(new_n8156_), .ZN(new_n8191_));
  INV_X1     g07177(.I(new_n8156_), .ZN(new_n8192_));
  NAND3_X1   g07178(.A1(new_n8165_), .A2(new_n8186_), .A3(new_n8192_), .ZN(new_n8193_));
  AOI21_X1   g07179(.A1(new_n8191_), .A2(new_n8193_), .B(new_n8189_), .ZN(new_n8194_));
  AOI21_X1   g07180(.A1(new_n8165_), .A2(new_n8186_), .B(new_n8192_), .ZN(new_n8195_));
  NOR3_X1    g07181(.A1(new_n8180_), .A2(new_n8173_), .A3(new_n8156_), .ZN(new_n8196_));
  NOR3_X1    g07182(.A1(new_n8195_), .A2(new_n8196_), .A3(new_n8152_), .ZN(new_n8197_));
  NOR2_X1    g07183(.A1(new_n8190_), .A2(new_n8157_), .ZN(new_n8198_));
  NOR2_X1    g07184(.A1(new_n8180_), .A2(new_n8173_), .ZN(new_n8199_));
  AOI22_X1   g07185(.A1(new_n8177_), .A2(new_n8179_), .B1(new_n8170_), .B2(new_n8172_), .ZN(new_n8200_));
  NOR2_X1    g07186(.A1(new_n8199_), .A2(new_n8200_), .ZN(new_n8201_));
  AOI22_X1   g07187(.A1(new_n8119_), .A2(new_n8121_), .B1(new_n8126_), .B2(new_n8128_), .ZN(new_n8202_));
  NOR2_X1    g07188(.A1(new_n8142_), .A2(new_n8202_), .ZN(new_n8203_));
  NAND2_X1   g07189(.A1(new_n8109_), .A2(new_n8114_), .ZN(new_n8204_));
  NOR2_X1    g07190(.A1(new_n8129_), .A2(new_n8204_), .ZN(new_n8205_));
  NAND4_X1   g07191(.A1(new_n8201_), .A2(new_n8203_), .A3(new_n8198_), .A4(new_n8205_), .ZN(new_n8206_));
  NOR4_X1    g07192(.A1(new_n8206_), .A2(new_n8188_), .A3(new_n8194_), .A4(new_n8197_), .ZN(new_n8207_));
  NOR3_X1    g07193(.A1(new_n8194_), .A2(new_n8197_), .A3(new_n8188_), .ZN(new_n8208_));
  INV_X1     g07194(.I(new_n8198_), .ZN(new_n8209_));
  NAND2_X1   g07195(.A1(new_n8180_), .A2(new_n8173_), .ZN(new_n8210_));
  NAND2_X1   g07196(.A1(new_n8210_), .A2(new_n8190_), .ZN(new_n8211_));
  OAI22_X1   g07197(.A1(new_n8134_), .A2(new_n8136_), .B1(new_n8141_), .B2(new_n8139_), .ZN(new_n8212_));
  NAND2_X1   g07198(.A1(new_n8212_), .A2(new_n8129_), .ZN(new_n8213_));
  NAND3_X1   g07199(.A1(new_n8142_), .A2(new_n8109_), .A3(new_n8114_), .ZN(new_n8214_));
  NOR4_X1    g07200(.A1(new_n8209_), .A2(new_n8214_), .A3(new_n8211_), .A4(new_n8213_), .ZN(new_n8215_));
  NOR2_X1    g07201(.A1(new_n8208_), .A2(new_n8215_), .ZN(new_n8216_));
  OAI21_X1   g07202(.A1(new_n8216_), .A2(new_n8207_), .B(new_n8148_), .ZN(new_n8217_));
  OAI21_X1   g07203(.A1(new_n8195_), .A2(new_n8196_), .B(new_n8152_), .ZN(new_n8218_));
  NAND3_X1   g07204(.A1(new_n8191_), .A2(new_n8193_), .A3(new_n8189_), .ZN(new_n8219_));
  NAND2_X1   g07205(.A1(new_n8219_), .A2(new_n8218_), .ZN(new_n8220_));
  OAI21_X1   g07206(.A1(new_n8220_), .A2(new_n8188_), .B(new_n8215_), .ZN(new_n8221_));
  NAND3_X1   g07207(.A1(new_n8201_), .A2(new_n8203_), .A3(new_n8198_), .ZN(new_n8222_));
  NOR2_X1    g07208(.A1(new_n8188_), .A2(new_n8214_), .ZN(new_n8223_));
  OAI21_X1   g07209(.A1(new_n8220_), .A2(new_n8222_), .B(new_n8223_), .ZN(new_n8224_));
  NAND3_X1   g07210(.A1(new_n8221_), .A2(new_n8224_), .A3(new_n8148_), .ZN(new_n8225_));
  NAND2_X1   g07211(.A1(new_n8225_), .A2(new_n8217_), .ZN(new_n8226_));
  OR2_X2     g07212(.A1(new_n8147_), .A2(new_n8144_), .Z(new_n8227_));
  NAND2_X1   g07213(.A1(new_n8208_), .A2(new_n8215_), .ZN(new_n8228_));
  OAI21_X1   g07214(.A1(new_n8220_), .A2(new_n8188_), .B(new_n8206_), .ZN(new_n8229_));
  AOI21_X1   g07215(.A1(new_n8229_), .A2(new_n8228_), .B(new_n8227_), .ZN(new_n8230_));
  NOR2_X1    g07216(.A1(new_n8208_), .A2(new_n8206_), .ZN(new_n8231_));
  NOR2_X1    g07217(.A1(new_n8194_), .A2(new_n8197_), .ZN(new_n8232_));
  NOR3_X1    g07218(.A1(new_n8209_), .A2(new_n8211_), .A3(new_n8213_), .ZN(new_n8233_));
  NOR2_X1    g07219(.A1(new_n8186_), .A2(new_n8180_), .ZN(new_n8234_));
  NOR2_X1    g07220(.A1(new_n8165_), .A2(new_n8173_), .ZN(new_n8235_));
  NOR2_X1    g07221(.A1(new_n8234_), .A2(new_n8235_), .ZN(new_n8236_));
  OAI21_X1   g07222(.A1(new_n8236_), .A2(new_n8157_), .B(new_n8205_), .ZN(new_n8237_));
  AOI21_X1   g07223(.A1(new_n8232_), .A2(new_n8233_), .B(new_n8237_), .ZN(new_n8238_));
  NOR3_X1    g07224(.A1(new_n8238_), .A2(new_n8231_), .A3(new_n8227_), .ZN(new_n8239_));
  NOR2_X1    g07225(.A1(new_n8209_), .A2(new_n8211_), .ZN(new_n8240_));
  NAND2_X1   g07226(.A1(new_n8203_), .A2(new_n8205_), .ZN(new_n8241_));
  NOR2_X1    g07227(.A1(new_n8240_), .A2(new_n8241_), .ZN(new_n8242_));
  NAND2_X1   g07228(.A1(new_n8201_), .A2(new_n8198_), .ZN(new_n8243_));
  NOR2_X1    g07229(.A1(new_n8214_), .A2(new_n8213_), .ZN(new_n8244_));
  NOR2_X1    g07230(.A1(new_n8244_), .A2(new_n8243_), .ZN(new_n8245_));
  INV_X1     g07231(.I(\A[927] ), .ZN(new_n8246_));
  NOR2_X1    g07232(.A1(new_n8246_), .A2(\A[926] ), .ZN(new_n8247_));
  INV_X1     g07233(.I(\A[926] ), .ZN(new_n8248_));
  NOR2_X1    g07234(.A1(new_n8248_), .A2(\A[927] ), .ZN(new_n8249_));
  OAI21_X1   g07235(.A1(new_n8247_), .A2(new_n8249_), .B(\A[925] ), .ZN(new_n8250_));
  INV_X1     g07236(.I(\A[925] ), .ZN(new_n8251_));
  NOR2_X1    g07237(.A1(\A[926] ), .A2(\A[927] ), .ZN(new_n8252_));
  NAND2_X1   g07238(.A1(\A[926] ), .A2(\A[927] ), .ZN(new_n8253_));
  INV_X1     g07239(.I(new_n8253_), .ZN(new_n8254_));
  OAI21_X1   g07240(.A1(new_n8254_), .A2(new_n8252_), .B(new_n8251_), .ZN(new_n8255_));
  NAND2_X1   g07241(.A1(new_n8250_), .A2(new_n8255_), .ZN(new_n8256_));
  INV_X1     g07242(.I(\A[930] ), .ZN(new_n8257_));
  NOR2_X1    g07243(.A1(new_n8257_), .A2(\A[929] ), .ZN(new_n8258_));
  INV_X1     g07244(.I(\A[929] ), .ZN(new_n8259_));
  NOR2_X1    g07245(.A1(new_n8259_), .A2(\A[930] ), .ZN(new_n8260_));
  OAI21_X1   g07246(.A1(new_n8258_), .A2(new_n8260_), .B(\A[928] ), .ZN(new_n8261_));
  INV_X1     g07247(.I(\A[928] ), .ZN(new_n8262_));
  NOR2_X1    g07248(.A1(\A[929] ), .A2(\A[930] ), .ZN(new_n8263_));
  AND2_X2    g07249(.A1(\A[929] ), .A2(\A[930] ), .Z(new_n8264_));
  OAI21_X1   g07250(.A1(new_n8264_), .A2(new_n8263_), .B(new_n8262_), .ZN(new_n8265_));
  NAND2_X1   g07251(.A1(new_n8261_), .A2(new_n8265_), .ZN(new_n8266_));
  NAND2_X1   g07252(.A1(\A[929] ), .A2(\A[930] ), .ZN(new_n8267_));
  AOI21_X1   g07253(.A1(new_n8262_), .A2(new_n8267_), .B(new_n8263_), .ZN(new_n8268_));
  AOI21_X1   g07254(.A1(new_n8251_), .A2(new_n8253_), .B(new_n8252_), .ZN(new_n8269_));
  NAND2_X1   g07255(.A1(new_n8268_), .A2(new_n8269_), .ZN(new_n8270_));
  NOR3_X1    g07256(.A1(new_n8256_), .A2(new_n8266_), .A3(new_n8270_), .ZN(new_n8271_));
  NOR2_X1    g07257(.A1(new_n8256_), .A2(new_n8266_), .ZN(new_n8272_));
  NAND2_X1   g07258(.A1(new_n8248_), .A2(\A[927] ), .ZN(new_n8273_));
  NAND2_X1   g07259(.A1(new_n8246_), .A2(\A[926] ), .ZN(new_n8274_));
  AOI21_X1   g07260(.A1(new_n8273_), .A2(new_n8274_), .B(new_n8251_), .ZN(new_n8275_));
  INV_X1     g07261(.I(new_n8252_), .ZN(new_n8276_));
  AOI21_X1   g07262(.A1(new_n8276_), .A2(new_n8253_), .B(\A[925] ), .ZN(new_n8277_));
  NOR2_X1    g07263(.A1(new_n8277_), .A2(new_n8275_), .ZN(new_n8278_));
  NAND2_X1   g07264(.A1(new_n8259_), .A2(\A[930] ), .ZN(new_n8279_));
  NAND2_X1   g07265(.A1(new_n8257_), .A2(\A[929] ), .ZN(new_n8280_));
  AOI21_X1   g07266(.A1(new_n8279_), .A2(new_n8280_), .B(new_n8262_), .ZN(new_n8281_));
  INV_X1     g07267(.I(new_n8263_), .ZN(new_n8282_));
  AOI21_X1   g07268(.A1(new_n8282_), .A2(new_n8267_), .B(\A[928] ), .ZN(new_n8283_));
  NOR2_X1    g07269(.A1(new_n8283_), .A2(new_n8281_), .ZN(new_n8284_));
  NOR2_X1    g07270(.A1(new_n8278_), .A2(new_n8284_), .ZN(new_n8285_));
  NOR2_X1    g07271(.A1(new_n8285_), .A2(new_n8272_), .ZN(new_n8286_));
  INV_X1     g07272(.I(\A[919] ), .ZN(new_n8287_));
  INV_X1     g07273(.I(\A[920] ), .ZN(new_n8288_));
  NAND2_X1   g07274(.A1(new_n8288_), .A2(\A[921] ), .ZN(new_n8289_));
  INV_X1     g07275(.I(\A[921] ), .ZN(new_n8290_));
  NAND2_X1   g07276(.A1(new_n8290_), .A2(\A[920] ), .ZN(new_n8291_));
  AOI21_X1   g07277(.A1(new_n8289_), .A2(new_n8291_), .B(new_n8287_), .ZN(new_n8292_));
  NOR2_X1    g07278(.A1(\A[920] ), .A2(\A[921] ), .ZN(new_n8293_));
  INV_X1     g07279(.I(new_n8293_), .ZN(new_n8294_));
  NAND2_X1   g07280(.A1(\A[920] ), .A2(\A[921] ), .ZN(new_n8295_));
  AOI21_X1   g07281(.A1(new_n8294_), .A2(new_n8295_), .B(\A[919] ), .ZN(new_n8296_));
  NOR2_X1    g07282(.A1(new_n8296_), .A2(new_n8292_), .ZN(new_n8297_));
  INV_X1     g07283(.I(\A[922] ), .ZN(new_n8298_));
  INV_X1     g07284(.I(\A[923] ), .ZN(new_n8299_));
  NAND2_X1   g07285(.A1(new_n8299_), .A2(\A[924] ), .ZN(new_n8300_));
  INV_X1     g07286(.I(\A[924] ), .ZN(new_n8301_));
  NAND2_X1   g07287(.A1(new_n8301_), .A2(\A[923] ), .ZN(new_n8302_));
  AOI21_X1   g07288(.A1(new_n8300_), .A2(new_n8302_), .B(new_n8298_), .ZN(new_n8303_));
  NOR2_X1    g07289(.A1(\A[923] ), .A2(\A[924] ), .ZN(new_n8304_));
  INV_X1     g07290(.I(new_n8304_), .ZN(new_n8305_));
  NAND2_X1   g07291(.A1(\A[923] ), .A2(\A[924] ), .ZN(new_n8306_));
  AOI21_X1   g07292(.A1(new_n8305_), .A2(new_n8306_), .B(\A[922] ), .ZN(new_n8307_));
  NOR2_X1    g07293(.A1(new_n8307_), .A2(new_n8303_), .ZN(new_n8308_));
  AOI21_X1   g07294(.A1(new_n8298_), .A2(new_n8306_), .B(new_n8304_), .ZN(new_n8309_));
  AOI21_X1   g07295(.A1(new_n8287_), .A2(new_n8295_), .B(new_n8293_), .ZN(new_n8310_));
  NAND2_X1   g07296(.A1(new_n8309_), .A2(new_n8310_), .ZN(new_n8311_));
  AND2_X2    g07297(.A1(new_n8286_), .A2(new_n8271_), .Z(new_n8313_));
  NOR3_X1    g07298(.A1(new_n8242_), .A2(new_n8245_), .A3(new_n8313_), .ZN(new_n8314_));
  INV_X1     g07299(.I(new_n8314_), .ZN(new_n8315_));
  OAI21_X1   g07300(.A1(new_n8230_), .A2(new_n8239_), .B(new_n8315_), .ZN(new_n8316_));
  NAND3_X1   g07301(.A1(new_n8225_), .A2(new_n8217_), .A3(new_n8314_), .ZN(new_n8317_));
  NAND2_X1   g07302(.A1(new_n8278_), .A2(new_n8284_), .ZN(new_n8318_));
  NAND2_X1   g07303(.A1(new_n8256_), .A2(new_n8266_), .ZN(new_n8319_));
  NAND3_X1   g07304(.A1(new_n8271_), .A2(new_n8318_), .A3(new_n8319_), .ZN(new_n8320_));
  NOR4_X1    g07305(.A1(new_n8292_), .A2(new_n8296_), .A3(new_n8307_), .A4(new_n8303_), .ZN(new_n8321_));
  INV_X1     g07306(.I(new_n8321_), .ZN(new_n8322_));
  NOR2_X1    g07307(.A1(new_n8290_), .A2(\A[920] ), .ZN(new_n8323_));
  NOR2_X1    g07308(.A1(new_n8288_), .A2(\A[921] ), .ZN(new_n8324_));
  OAI21_X1   g07309(.A1(new_n8323_), .A2(new_n8324_), .B(\A[919] ), .ZN(new_n8325_));
  INV_X1     g07310(.I(new_n8295_), .ZN(new_n8326_));
  OAI21_X1   g07311(.A1(new_n8326_), .A2(new_n8293_), .B(new_n8287_), .ZN(new_n8327_));
  NAND2_X1   g07312(.A1(new_n8325_), .A2(new_n8327_), .ZN(new_n8328_));
  NOR2_X1    g07313(.A1(new_n8301_), .A2(\A[923] ), .ZN(new_n8329_));
  NOR2_X1    g07314(.A1(new_n8299_), .A2(\A[924] ), .ZN(new_n8330_));
  OAI21_X1   g07315(.A1(new_n8329_), .A2(new_n8330_), .B(\A[922] ), .ZN(new_n8331_));
  INV_X1     g07316(.I(new_n8306_), .ZN(new_n8332_));
  OAI21_X1   g07317(.A1(new_n8332_), .A2(new_n8304_), .B(new_n8298_), .ZN(new_n8333_));
  NAND2_X1   g07318(.A1(new_n8331_), .A2(new_n8333_), .ZN(new_n8334_));
  NAND2_X1   g07319(.A1(new_n8328_), .A2(new_n8334_), .ZN(new_n8335_));
  NAND2_X1   g07320(.A1(new_n8322_), .A2(new_n8335_), .ZN(new_n8336_));
  INV_X1     g07321(.I(new_n8268_), .ZN(new_n8337_));
  OAI21_X1   g07322(.A1(new_n8256_), .A2(new_n8266_), .B(new_n8269_), .ZN(new_n8338_));
  INV_X1     g07323(.I(new_n8269_), .ZN(new_n8339_));
  NAND3_X1   g07324(.A1(new_n8278_), .A2(new_n8284_), .A3(new_n8339_), .ZN(new_n8340_));
  AOI21_X1   g07325(.A1(new_n8340_), .A2(new_n8338_), .B(new_n8337_), .ZN(new_n8341_));
  AOI21_X1   g07326(.A1(new_n8278_), .A2(new_n8284_), .B(new_n8339_), .ZN(new_n8342_));
  NOR3_X1    g07327(.A1(new_n8256_), .A2(new_n8266_), .A3(new_n8269_), .ZN(new_n8343_));
  NOR3_X1    g07328(.A1(new_n8342_), .A2(new_n8343_), .A3(new_n8268_), .ZN(new_n8344_));
  NOR4_X1    g07329(.A1(new_n8341_), .A2(new_n8344_), .A3(new_n8320_), .A4(new_n8336_), .ZN(new_n8345_));
  NOR3_X1    g07330(.A1(new_n8328_), .A2(new_n8334_), .A3(new_n8311_), .ZN(new_n8346_));
  INV_X1     g07331(.I(new_n8270_), .ZN(new_n8347_));
  NOR2_X1    g07332(.A1(new_n8284_), .A2(new_n8256_), .ZN(new_n8348_));
  NOR2_X1    g07333(.A1(new_n8278_), .A2(new_n8266_), .ZN(new_n8349_));
  OAI21_X1   g07334(.A1(new_n8348_), .A2(new_n8349_), .B(new_n8347_), .ZN(new_n8350_));
  NAND2_X1   g07335(.A1(new_n8350_), .A2(new_n8346_), .ZN(new_n8351_));
  INV_X1     g07336(.I(new_n8309_), .ZN(new_n8352_));
  OAI21_X1   g07337(.A1(new_n8328_), .A2(new_n8334_), .B(new_n8310_), .ZN(new_n8353_));
  INV_X1     g07338(.I(new_n8310_), .ZN(new_n8354_));
  NAND3_X1   g07339(.A1(new_n8297_), .A2(new_n8308_), .A3(new_n8354_), .ZN(new_n8355_));
  AOI21_X1   g07340(.A1(new_n8353_), .A2(new_n8355_), .B(new_n8352_), .ZN(new_n8356_));
  NOR2_X1    g07341(.A1(new_n8321_), .A2(new_n8354_), .ZN(new_n8357_));
  NOR3_X1    g07342(.A1(new_n8328_), .A2(new_n8334_), .A3(new_n8310_), .ZN(new_n8358_));
  NOR3_X1    g07343(.A1(new_n8357_), .A2(new_n8358_), .A3(new_n8309_), .ZN(new_n8359_));
  NOR2_X1    g07344(.A1(new_n8359_), .A2(new_n8356_), .ZN(new_n8360_));
  NOR3_X1    g07345(.A1(new_n8345_), .A2(new_n8360_), .A3(new_n8351_), .ZN(new_n8361_));
  INV_X1     g07346(.I(new_n8361_), .ZN(new_n8362_));
  OAI21_X1   g07347(.A1(new_n8357_), .A2(new_n8358_), .B(new_n8309_), .ZN(new_n8363_));
  NAND3_X1   g07348(.A1(new_n8353_), .A2(new_n8355_), .A3(new_n8352_), .ZN(new_n8364_));
  NAND2_X1   g07349(.A1(new_n8363_), .A2(new_n8364_), .ZN(new_n8365_));
  NOR2_X1    g07350(.A1(new_n8297_), .A2(new_n8308_), .ZN(new_n8366_));
  NOR2_X1    g07351(.A1(new_n8366_), .A2(new_n8321_), .ZN(new_n8367_));
  NAND4_X1   g07352(.A1(new_n8286_), .A2(new_n8367_), .A3(new_n8271_), .A4(new_n8346_), .ZN(new_n8368_));
  NAND2_X1   g07353(.A1(new_n8365_), .A2(new_n8368_), .ZN(new_n8369_));
  NAND3_X1   g07354(.A1(new_n8322_), .A2(new_n8346_), .A3(new_n8335_), .ZN(new_n8370_));
  NOR2_X1    g07355(.A1(new_n8370_), .A2(new_n8320_), .ZN(new_n8371_));
  NAND2_X1   g07356(.A1(new_n8278_), .A2(new_n8266_), .ZN(new_n8372_));
  NAND2_X1   g07357(.A1(new_n8284_), .A2(new_n8256_), .ZN(new_n8373_));
  AOI21_X1   g07358(.A1(new_n8373_), .A2(new_n8372_), .B(new_n8270_), .ZN(new_n8374_));
  NOR3_X1    g07359(.A1(new_n8344_), .A2(new_n8341_), .A3(new_n8374_), .ZN(new_n8375_));
  AOI21_X1   g07360(.A1(new_n8360_), .A2(new_n8371_), .B(new_n8375_), .ZN(new_n8376_));
  OAI21_X1   g07361(.A1(new_n8342_), .A2(new_n8343_), .B(new_n8268_), .ZN(new_n8377_));
  NAND3_X1   g07362(.A1(new_n8340_), .A2(new_n8338_), .A3(new_n8337_), .ZN(new_n8378_));
  NAND3_X1   g07363(.A1(new_n8377_), .A2(new_n8378_), .A3(new_n8350_), .ZN(new_n8379_));
  NOR3_X1    g07364(.A1(new_n8379_), .A2(new_n8365_), .A3(new_n8368_), .ZN(new_n8380_));
  OAI21_X1   g07365(.A1(new_n8376_), .A2(new_n8380_), .B(new_n8369_), .ZN(new_n8381_));
  NAND2_X1   g07366(.A1(new_n8381_), .A2(new_n8362_), .ZN(new_n8382_));
  AOI22_X1   g07367(.A1(new_n8316_), .A2(new_n8317_), .B1(new_n8382_), .B2(new_n8226_), .ZN(new_n8383_));
  NOR2_X1    g07368(.A1(new_n8231_), .A2(new_n8148_), .ZN(new_n8384_));
  NOR2_X1    g07369(.A1(new_n8152_), .A2(new_n8156_), .ZN(new_n8385_));
  OAI21_X1   g07370(.A1(new_n8190_), .A2(new_n8385_), .B(new_n8157_), .ZN(new_n8386_));
  NOR2_X1    g07371(.A1(new_n8109_), .A2(new_n8114_), .ZN(new_n8387_));
  OAI21_X1   g07372(.A1(new_n8129_), .A2(new_n8387_), .B(new_n8204_), .ZN(new_n8388_));
  XNOR2_X1   g07373(.A1(new_n8388_), .A2(new_n8386_), .ZN(new_n8389_));
  INV_X1     g07374(.I(new_n8389_), .ZN(new_n8390_));
  NOR3_X1    g07375(.A1(new_n8384_), .A2(new_n8390_), .A3(new_n8238_), .ZN(new_n8391_));
  NOR2_X1    g07376(.A1(new_n8345_), .A2(new_n8351_), .ZN(new_n8392_));
  AOI21_X1   g07377(.A1(new_n8371_), .A2(new_n8379_), .B(new_n8360_), .ZN(new_n8393_));
  NAND2_X1   g07378(.A1(new_n8339_), .A2(new_n8337_), .ZN(new_n8394_));
  AOI21_X1   g07379(.A1(new_n8272_), .A2(new_n8394_), .B(new_n8347_), .ZN(new_n8395_));
  NOR2_X1    g07380(.A1(new_n8309_), .A2(new_n8310_), .ZN(new_n8396_));
  OAI21_X1   g07381(.A1(new_n8322_), .A2(new_n8396_), .B(new_n8311_), .ZN(new_n8397_));
  XNOR2_X1   g07382(.A1(new_n8397_), .A2(new_n8395_), .ZN(new_n8398_));
  NOR3_X1    g07383(.A1(new_n8393_), .A2(new_n8398_), .A3(new_n8392_), .ZN(new_n8399_));
  XOR2_X1    g07384(.A1(new_n8391_), .A2(new_n8399_), .Z(new_n8400_));
  NAND2_X1   g07385(.A1(new_n8400_), .A2(new_n8383_), .ZN(new_n8401_));
  NOR2_X1    g07386(.A1(new_n8239_), .A2(new_n8230_), .ZN(new_n8402_));
  AOI21_X1   g07387(.A1(new_n8225_), .A2(new_n8217_), .B(new_n8314_), .ZN(new_n8403_));
  NOR3_X1    g07388(.A1(new_n8239_), .A2(new_n8315_), .A3(new_n8230_), .ZN(new_n8404_));
  OAI21_X1   g07389(.A1(new_n8365_), .A2(new_n8368_), .B(new_n8379_), .ZN(new_n8405_));
  NAND3_X1   g07390(.A1(new_n8375_), .A2(new_n8360_), .A3(new_n8371_), .ZN(new_n8406_));
  NAND2_X1   g07391(.A1(new_n8405_), .A2(new_n8406_), .ZN(new_n8407_));
  AOI21_X1   g07392(.A1(new_n8407_), .A2(new_n8369_), .B(new_n8361_), .ZN(new_n8408_));
  OAI22_X1   g07393(.A1(new_n8404_), .A2(new_n8403_), .B1(new_n8408_), .B2(new_n8402_), .ZN(new_n8409_));
  NOR2_X1    g07394(.A1(new_n8391_), .A2(new_n8399_), .ZN(new_n8410_));
  NAND2_X1   g07395(.A1(new_n8221_), .A2(new_n8227_), .ZN(new_n8411_));
  NAND3_X1   g07396(.A1(new_n8411_), .A2(new_n8389_), .A3(new_n8224_), .ZN(new_n8412_));
  INV_X1     g07397(.I(new_n8399_), .ZN(new_n8413_));
  NOR2_X1    g07398(.A1(new_n8413_), .A2(new_n8412_), .ZN(new_n8414_));
  OAI21_X1   g07399(.A1(new_n8410_), .A2(new_n8414_), .B(new_n8409_), .ZN(new_n8415_));
  NAND2_X1   g07400(.A1(new_n8415_), .A2(new_n8401_), .ZN(new_n8416_));
  NOR2_X1    g07401(.A1(new_n8416_), .A2(new_n8105_), .ZN(new_n8417_));
  NOR3_X1    g07402(.A1(new_n8404_), .A2(new_n8382_), .A3(new_n8403_), .ZN(new_n8418_));
  INV_X1     g07403(.I(new_n8418_), .ZN(new_n8419_));
  OAI21_X1   g07404(.A1(new_n8242_), .A2(new_n8245_), .B(new_n8313_), .ZN(new_n8420_));
  NOR2_X1    g07405(.A1(new_n7933_), .A2(new_n8001_), .ZN(new_n8421_));
  NOR2_X1    g07406(.A1(new_n8421_), .A2(new_n8005_), .ZN(new_n8422_));
  NAND3_X1   g07407(.A1(new_n8422_), .A2(new_n8315_), .A3(new_n8420_), .ZN(new_n8423_));
  INV_X1     g07408(.I(new_n8423_), .ZN(new_n8424_));
  NOR2_X1    g07409(.A1(new_n8424_), .A2(new_n8418_), .ZN(new_n8425_));
  INV_X1     g07410(.I(new_n8425_), .ZN(new_n8426_));
  NAND2_X1   g07411(.A1(new_n8424_), .A2(new_n8418_), .ZN(new_n8427_));
  OAI21_X1   g07412(.A1(new_n8092_), .A2(new_n8091_), .B(new_n8096_), .ZN(new_n8428_));
  NAND3_X1   g07413(.A1(new_n8003_), .A2(new_n8071_), .A3(new_n8006_), .ZN(new_n8429_));
  NAND2_X1   g07414(.A1(new_n8428_), .A2(new_n8429_), .ZN(new_n8430_));
  AOI22_X1   g07415(.A1(new_n8426_), .A2(new_n8427_), .B1(new_n8419_), .B2(new_n8430_), .ZN(new_n8431_));
  AOI22_X1   g07416(.A1(new_n8401_), .A2(new_n8415_), .B1(new_n8089_), .B2(new_n8104_), .ZN(new_n8432_));
  INV_X1     g07417(.I(new_n8432_), .ZN(new_n8433_));
  AOI21_X1   g07418(.A1(new_n8433_), .A2(new_n8431_), .B(new_n8417_), .ZN(new_n8434_));
  NAND2_X1   g07419(.A1(new_n8075_), .A2(new_n8077_), .ZN(new_n8435_));
  NOR2_X1    g07420(.A1(new_n8073_), .A2(new_n7925_), .ZN(new_n8436_));
  OAI21_X1   g07421(.A1(new_n8075_), .A2(new_n8077_), .B(new_n8436_), .ZN(new_n8437_));
  NAND2_X1   g07422(.A1(new_n8437_), .A2(new_n8435_), .ZN(new_n8438_));
  INV_X1     g07423(.I(new_n8083_), .ZN(new_n8439_));
  NAND2_X1   g07424(.A1(new_n8439_), .A2(new_n8085_), .ZN(new_n8440_));
  NOR2_X1    g07425(.A1(new_n8081_), .A2(new_n8040_), .ZN(new_n8441_));
  OAI21_X1   g07426(.A1(new_n8439_), .A2(new_n8085_), .B(new_n8441_), .ZN(new_n8442_));
  NAND2_X1   g07427(.A1(new_n8442_), .A2(new_n8440_), .ZN(new_n8443_));
  INV_X1     g07428(.I(new_n8443_), .ZN(new_n8444_));
  AOI21_X1   g07429(.A1(new_n8097_), .A2(new_n8101_), .B(new_n8102_), .ZN(new_n8445_));
  NOR2_X1    g07430(.A1(new_n8445_), .A2(new_n8444_), .ZN(new_n8446_));
  NAND3_X1   g07431(.A1(new_n8072_), .A2(new_n8080_), .A3(new_n8087_), .ZN(new_n8447_));
  NOR2_X1    g07432(.A1(new_n8447_), .A2(new_n8443_), .ZN(new_n8448_));
  OAI21_X1   g07433(.A1(new_n8446_), .A2(new_n8448_), .B(new_n8438_), .ZN(new_n8449_));
  INV_X1     g07434(.I(new_n8438_), .ZN(new_n8450_));
  NAND2_X1   g07435(.A1(new_n8447_), .A2(new_n8443_), .ZN(new_n8451_));
  NAND4_X1   g07436(.A1(new_n8444_), .A2(new_n8072_), .A3(new_n8080_), .A4(new_n8087_), .ZN(new_n8452_));
  NAND3_X1   g07437(.A1(new_n8451_), .A2(new_n8450_), .A3(new_n8452_), .ZN(new_n8453_));
  NAND2_X1   g07438(.A1(new_n8449_), .A2(new_n8453_), .ZN(new_n8454_));
  NAND2_X1   g07439(.A1(new_n8388_), .A2(new_n8386_), .ZN(new_n8455_));
  NOR2_X1    g07440(.A1(new_n8384_), .A2(new_n8238_), .ZN(new_n8456_));
  OAI21_X1   g07441(.A1(new_n8386_), .A2(new_n8388_), .B(new_n8456_), .ZN(new_n8457_));
  NAND2_X1   g07442(.A1(new_n8457_), .A2(new_n8455_), .ZN(new_n8458_));
  INV_X1     g07443(.I(new_n8458_), .ZN(new_n8459_));
  INV_X1     g07444(.I(new_n8395_), .ZN(new_n8460_));
  NAND2_X1   g07445(.A1(new_n8460_), .A2(new_n8397_), .ZN(new_n8461_));
  NOR2_X1    g07446(.A1(new_n8393_), .A2(new_n8392_), .ZN(new_n8462_));
  OAI21_X1   g07447(.A1(new_n8460_), .A2(new_n8397_), .B(new_n8462_), .ZN(new_n8463_));
  NAND2_X1   g07448(.A1(new_n8463_), .A2(new_n8461_), .ZN(new_n8464_));
  NAND3_X1   g07449(.A1(new_n8383_), .A2(new_n8391_), .A3(new_n8399_), .ZN(new_n8465_));
  NAND2_X1   g07450(.A1(new_n8465_), .A2(new_n8464_), .ZN(new_n8466_));
  INV_X1     g07451(.I(new_n8464_), .ZN(new_n8467_));
  NAND4_X1   g07452(.A1(new_n8467_), .A2(new_n8383_), .A3(new_n8391_), .A4(new_n8399_), .ZN(new_n8468_));
  AOI21_X1   g07453(.A1(new_n8466_), .A2(new_n8468_), .B(new_n8459_), .ZN(new_n8469_));
  INV_X1     g07454(.I(new_n8410_), .ZN(new_n8470_));
  NAND2_X1   g07455(.A1(new_n8409_), .A2(new_n8470_), .ZN(new_n8471_));
  AOI21_X1   g07456(.A1(new_n8471_), .A2(new_n8414_), .B(new_n8467_), .ZN(new_n8472_));
  NOR4_X1    g07457(.A1(new_n8409_), .A2(new_n8412_), .A3(new_n8413_), .A4(new_n8464_), .ZN(new_n8473_));
  NOR3_X1    g07458(.A1(new_n8472_), .A2(new_n8458_), .A3(new_n8473_), .ZN(new_n8474_));
  NOR2_X1    g07459(.A1(new_n8474_), .A2(new_n8469_), .ZN(new_n8475_));
  NAND2_X1   g07460(.A1(new_n8454_), .A2(new_n8475_), .ZN(new_n8476_));
  AOI21_X1   g07461(.A1(new_n8451_), .A2(new_n8452_), .B(new_n8450_), .ZN(new_n8477_));
  NOR3_X1    g07462(.A1(new_n8446_), .A2(new_n8448_), .A3(new_n8438_), .ZN(new_n8478_));
  NOR2_X1    g07463(.A1(new_n8478_), .A2(new_n8477_), .ZN(new_n8479_));
  OAI21_X1   g07464(.A1(new_n8472_), .A2(new_n8473_), .B(new_n8458_), .ZN(new_n8480_));
  NAND3_X1   g07465(.A1(new_n8466_), .A2(new_n8459_), .A3(new_n8468_), .ZN(new_n8481_));
  NAND2_X1   g07466(.A1(new_n8480_), .A2(new_n8481_), .ZN(new_n8482_));
  NAND2_X1   g07467(.A1(new_n8479_), .A2(new_n8482_), .ZN(new_n8483_));
  AOI21_X1   g07468(.A1(new_n8476_), .A2(new_n8483_), .B(new_n8434_), .ZN(new_n8484_));
  NAND4_X1   g07469(.A1(new_n8089_), .A2(new_n8415_), .A3(new_n8401_), .A4(new_n8104_), .ZN(new_n8485_));
  INV_X1     g07470(.I(new_n8427_), .ZN(new_n8486_));
  INV_X1     g07471(.I(new_n8430_), .ZN(new_n8487_));
  OAI22_X1   g07472(.A1(new_n8487_), .A2(new_n8418_), .B1(new_n8486_), .B2(new_n8425_), .ZN(new_n8488_));
  OAI21_X1   g07473(.A1(new_n8488_), .A2(new_n8432_), .B(new_n8485_), .ZN(new_n8489_));
  NAND4_X1   g07474(.A1(new_n8449_), .A2(new_n8453_), .A3(new_n8480_), .A4(new_n8481_), .ZN(new_n8490_));
  NAND2_X1   g07475(.A1(new_n8454_), .A2(new_n8482_), .ZN(new_n8491_));
  AOI21_X1   g07476(.A1(new_n8491_), .A2(new_n8490_), .B(new_n8489_), .ZN(new_n8492_));
  INV_X1     g07477(.I(\A[862] ), .ZN(new_n8493_));
  NOR2_X1    g07478(.A1(\A[863] ), .A2(\A[864] ), .ZN(new_n8494_));
  NAND2_X1   g07479(.A1(\A[863] ), .A2(\A[864] ), .ZN(new_n8495_));
  AOI21_X1   g07480(.A1(new_n8493_), .A2(new_n8495_), .B(new_n8494_), .ZN(new_n8496_));
  INV_X1     g07481(.I(\A[859] ), .ZN(new_n8497_));
  NOR2_X1    g07482(.A1(\A[860] ), .A2(\A[861] ), .ZN(new_n8498_));
  NAND2_X1   g07483(.A1(\A[860] ), .A2(\A[861] ), .ZN(new_n8499_));
  AOI21_X1   g07484(.A1(new_n8497_), .A2(new_n8499_), .B(new_n8498_), .ZN(new_n8500_));
  INV_X1     g07485(.I(new_n8500_), .ZN(new_n8501_));
  INV_X1     g07486(.I(\A[860] ), .ZN(new_n8502_));
  NAND2_X1   g07487(.A1(new_n8502_), .A2(\A[861] ), .ZN(new_n8503_));
  INV_X1     g07488(.I(\A[861] ), .ZN(new_n8504_));
  NAND2_X1   g07489(.A1(new_n8504_), .A2(\A[860] ), .ZN(new_n8505_));
  AOI21_X1   g07490(.A1(new_n8503_), .A2(new_n8505_), .B(new_n8497_), .ZN(new_n8506_));
  INV_X1     g07491(.I(new_n8498_), .ZN(new_n8507_));
  AOI21_X1   g07492(.A1(new_n8507_), .A2(new_n8499_), .B(\A[859] ), .ZN(new_n8508_));
  INV_X1     g07493(.I(\A[863] ), .ZN(new_n8509_));
  NAND2_X1   g07494(.A1(new_n8509_), .A2(\A[864] ), .ZN(new_n8510_));
  INV_X1     g07495(.I(\A[864] ), .ZN(new_n8511_));
  NAND2_X1   g07496(.A1(new_n8511_), .A2(\A[863] ), .ZN(new_n8512_));
  AOI21_X1   g07497(.A1(new_n8510_), .A2(new_n8512_), .B(new_n8493_), .ZN(new_n8513_));
  INV_X1     g07498(.I(new_n8494_), .ZN(new_n8514_));
  AOI21_X1   g07499(.A1(new_n8514_), .A2(new_n8495_), .B(\A[862] ), .ZN(new_n8515_));
  NOR4_X1    g07500(.A1(new_n8506_), .A2(new_n8508_), .A3(new_n8515_), .A4(new_n8513_), .ZN(new_n8516_));
  NOR2_X1    g07501(.A1(new_n8516_), .A2(new_n8501_), .ZN(new_n8517_));
  NOR2_X1    g07502(.A1(new_n8504_), .A2(\A[860] ), .ZN(new_n8518_));
  NOR2_X1    g07503(.A1(new_n8502_), .A2(\A[861] ), .ZN(new_n8519_));
  OAI21_X1   g07504(.A1(new_n8518_), .A2(new_n8519_), .B(\A[859] ), .ZN(new_n8520_));
  INV_X1     g07505(.I(new_n8499_), .ZN(new_n8521_));
  OAI21_X1   g07506(.A1(new_n8521_), .A2(new_n8498_), .B(new_n8497_), .ZN(new_n8522_));
  NOR2_X1    g07507(.A1(new_n8511_), .A2(\A[863] ), .ZN(new_n8523_));
  NOR2_X1    g07508(.A1(new_n8509_), .A2(\A[864] ), .ZN(new_n8524_));
  OAI21_X1   g07509(.A1(new_n8523_), .A2(new_n8524_), .B(\A[862] ), .ZN(new_n8525_));
  INV_X1     g07510(.I(new_n8495_), .ZN(new_n8526_));
  OAI21_X1   g07511(.A1(new_n8526_), .A2(new_n8494_), .B(new_n8493_), .ZN(new_n8527_));
  NAND4_X1   g07512(.A1(new_n8520_), .A2(new_n8522_), .A3(new_n8525_), .A4(new_n8527_), .ZN(new_n8528_));
  NOR2_X1    g07513(.A1(new_n8528_), .A2(new_n8500_), .ZN(new_n8529_));
  OAI21_X1   g07514(.A1(new_n8517_), .A2(new_n8529_), .B(new_n8496_), .ZN(new_n8530_));
  INV_X1     g07515(.I(new_n8496_), .ZN(new_n8531_));
  NAND2_X1   g07516(.A1(new_n8528_), .A2(new_n8500_), .ZN(new_n8532_));
  NAND2_X1   g07517(.A1(new_n8516_), .A2(new_n8501_), .ZN(new_n8533_));
  NAND3_X1   g07518(.A1(new_n8533_), .A2(new_n8532_), .A3(new_n8531_), .ZN(new_n8534_));
  NAND2_X1   g07519(.A1(new_n8530_), .A2(new_n8534_), .ZN(new_n8535_));
  INV_X1     g07520(.I(new_n8535_), .ZN(new_n8536_));
  INV_X1     g07521(.I(\A[868] ), .ZN(new_n8537_));
  NOR2_X1    g07522(.A1(\A[869] ), .A2(\A[870] ), .ZN(new_n8538_));
  NAND2_X1   g07523(.A1(\A[869] ), .A2(\A[870] ), .ZN(new_n8539_));
  AOI21_X1   g07524(.A1(new_n8537_), .A2(new_n8539_), .B(new_n8538_), .ZN(new_n8540_));
  INV_X1     g07525(.I(\A[865] ), .ZN(new_n8541_));
  NOR2_X1    g07526(.A1(\A[866] ), .A2(\A[867] ), .ZN(new_n8542_));
  NAND2_X1   g07527(.A1(\A[866] ), .A2(\A[867] ), .ZN(new_n8543_));
  AOI21_X1   g07528(.A1(new_n8541_), .A2(new_n8543_), .B(new_n8542_), .ZN(new_n8544_));
  NAND2_X1   g07529(.A1(new_n8540_), .A2(new_n8544_), .ZN(new_n8545_));
  INV_X1     g07530(.I(\A[866] ), .ZN(new_n8546_));
  NAND2_X1   g07531(.A1(new_n8546_), .A2(\A[867] ), .ZN(new_n8547_));
  INV_X1     g07532(.I(\A[867] ), .ZN(new_n8548_));
  NAND2_X1   g07533(.A1(new_n8548_), .A2(\A[866] ), .ZN(new_n8549_));
  AOI21_X1   g07534(.A1(new_n8547_), .A2(new_n8549_), .B(new_n8541_), .ZN(new_n8550_));
  INV_X1     g07535(.I(new_n8542_), .ZN(new_n8551_));
  AOI21_X1   g07536(.A1(new_n8551_), .A2(new_n8543_), .B(\A[865] ), .ZN(new_n8552_));
  NOR2_X1    g07537(.A1(new_n8552_), .A2(new_n8550_), .ZN(new_n8553_));
  INV_X1     g07538(.I(\A[870] ), .ZN(new_n8554_));
  NOR2_X1    g07539(.A1(new_n8554_), .A2(\A[869] ), .ZN(new_n8555_));
  INV_X1     g07540(.I(\A[869] ), .ZN(new_n8556_));
  NOR2_X1    g07541(.A1(new_n8556_), .A2(\A[870] ), .ZN(new_n8557_));
  OAI21_X1   g07542(.A1(new_n8555_), .A2(new_n8557_), .B(\A[868] ), .ZN(new_n8558_));
  INV_X1     g07543(.I(new_n8539_), .ZN(new_n8559_));
  OAI21_X1   g07544(.A1(new_n8559_), .A2(new_n8538_), .B(new_n8537_), .ZN(new_n8560_));
  NAND2_X1   g07545(.A1(new_n8558_), .A2(new_n8560_), .ZN(new_n8561_));
  NAND2_X1   g07546(.A1(new_n8553_), .A2(new_n8561_), .ZN(new_n8562_));
  NOR2_X1    g07547(.A1(new_n8548_), .A2(\A[866] ), .ZN(new_n8563_));
  NOR2_X1    g07548(.A1(new_n8546_), .A2(\A[867] ), .ZN(new_n8564_));
  OAI21_X1   g07549(.A1(new_n8563_), .A2(new_n8564_), .B(\A[865] ), .ZN(new_n8565_));
  INV_X1     g07550(.I(new_n8543_), .ZN(new_n8566_));
  OAI21_X1   g07551(.A1(new_n8566_), .A2(new_n8542_), .B(new_n8541_), .ZN(new_n8567_));
  NAND2_X1   g07552(.A1(new_n8565_), .A2(new_n8567_), .ZN(new_n8568_));
  NAND2_X1   g07553(.A1(new_n8556_), .A2(\A[870] ), .ZN(new_n8569_));
  NAND2_X1   g07554(.A1(new_n8554_), .A2(\A[869] ), .ZN(new_n8570_));
  AOI21_X1   g07555(.A1(new_n8569_), .A2(new_n8570_), .B(new_n8537_), .ZN(new_n8571_));
  INV_X1     g07556(.I(new_n8538_), .ZN(new_n8572_));
  AOI21_X1   g07557(.A1(new_n8572_), .A2(new_n8539_), .B(\A[868] ), .ZN(new_n8573_));
  NOR2_X1    g07558(.A1(new_n8573_), .A2(new_n8571_), .ZN(new_n8574_));
  NAND2_X1   g07559(.A1(new_n8574_), .A2(new_n8568_), .ZN(new_n8575_));
  AOI21_X1   g07560(.A1(new_n8562_), .A2(new_n8575_), .B(new_n8545_), .ZN(new_n8576_));
  INV_X1     g07561(.I(new_n8540_), .ZN(new_n8577_));
  NAND4_X1   g07562(.A1(new_n8565_), .A2(new_n8567_), .A3(new_n8558_), .A4(new_n8560_), .ZN(new_n8578_));
  NAND2_X1   g07563(.A1(new_n8578_), .A2(new_n8544_), .ZN(new_n8579_));
  INV_X1     g07564(.I(new_n8544_), .ZN(new_n8580_));
  NAND3_X1   g07565(.A1(new_n8553_), .A2(new_n8574_), .A3(new_n8580_), .ZN(new_n8581_));
  AOI21_X1   g07566(.A1(new_n8579_), .A2(new_n8581_), .B(new_n8577_), .ZN(new_n8582_));
  AOI21_X1   g07567(.A1(new_n8553_), .A2(new_n8574_), .B(new_n8580_), .ZN(new_n8583_));
  NOR3_X1    g07568(.A1(new_n8568_), .A2(new_n8561_), .A3(new_n8544_), .ZN(new_n8584_));
  NOR3_X1    g07569(.A1(new_n8583_), .A2(new_n8584_), .A3(new_n8540_), .ZN(new_n8585_));
  NOR2_X1    g07570(.A1(new_n8578_), .A2(new_n8545_), .ZN(new_n8586_));
  NOR4_X1    g07571(.A1(new_n8550_), .A2(new_n8552_), .A3(new_n8573_), .A4(new_n8571_), .ZN(new_n8587_));
  NOR2_X1    g07572(.A1(new_n8553_), .A2(new_n8574_), .ZN(new_n8588_));
  NOR2_X1    g07573(.A1(new_n8588_), .A2(new_n8587_), .ZN(new_n8589_));
  AOI22_X1   g07574(.A1(new_n8520_), .A2(new_n8522_), .B1(new_n8525_), .B2(new_n8527_), .ZN(new_n8590_));
  NOR2_X1    g07575(.A1(new_n8590_), .A2(new_n8516_), .ZN(new_n8591_));
  NAND2_X1   g07576(.A1(new_n8496_), .A2(new_n8500_), .ZN(new_n8592_));
  NOR2_X1    g07577(.A1(new_n8528_), .A2(new_n8592_), .ZN(new_n8593_));
  NAND4_X1   g07578(.A1(new_n8589_), .A2(new_n8591_), .A3(new_n8586_), .A4(new_n8593_), .ZN(new_n8594_));
  NOR4_X1    g07579(.A1(new_n8594_), .A2(new_n8576_), .A3(new_n8582_), .A4(new_n8585_), .ZN(new_n8595_));
  NOR3_X1    g07580(.A1(new_n8582_), .A2(new_n8585_), .A3(new_n8576_), .ZN(new_n8596_));
  INV_X1     g07581(.I(new_n8545_), .ZN(new_n8597_));
  NAND2_X1   g07582(.A1(new_n8587_), .A2(new_n8597_), .ZN(new_n8598_));
  NAND2_X1   g07583(.A1(new_n8568_), .A2(new_n8561_), .ZN(new_n8599_));
  NAND2_X1   g07584(.A1(new_n8599_), .A2(new_n8578_), .ZN(new_n8600_));
  OAI22_X1   g07585(.A1(new_n8506_), .A2(new_n8508_), .B1(new_n8515_), .B2(new_n8513_), .ZN(new_n8601_));
  NAND2_X1   g07586(.A1(new_n8601_), .A2(new_n8528_), .ZN(new_n8602_));
  NAND3_X1   g07587(.A1(new_n8516_), .A2(new_n8496_), .A3(new_n8500_), .ZN(new_n8603_));
  NOR4_X1    g07588(.A1(new_n8600_), .A2(new_n8598_), .A3(new_n8603_), .A4(new_n8602_), .ZN(new_n8604_));
  NOR2_X1    g07589(.A1(new_n8596_), .A2(new_n8604_), .ZN(new_n8605_));
  OAI21_X1   g07590(.A1(new_n8605_), .A2(new_n8595_), .B(new_n8536_), .ZN(new_n8606_));
  OAI21_X1   g07591(.A1(new_n8583_), .A2(new_n8584_), .B(new_n8540_), .ZN(new_n8607_));
  NAND3_X1   g07592(.A1(new_n8579_), .A2(new_n8581_), .A3(new_n8577_), .ZN(new_n8608_));
  NAND2_X1   g07593(.A1(new_n8607_), .A2(new_n8608_), .ZN(new_n8609_));
  OAI21_X1   g07594(.A1(new_n8609_), .A2(new_n8576_), .B(new_n8604_), .ZN(new_n8610_));
  NOR2_X1    g07595(.A1(new_n8574_), .A2(new_n8568_), .ZN(new_n8611_));
  NOR2_X1    g07596(.A1(new_n8553_), .A2(new_n8561_), .ZN(new_n8612_));
  OAI21_X1   g07597(.A1(new_n8611_), .A2(new_n8612_), .B(new_n8597_), .ZN(new_n8613_));
  NOR4_X1    g07598(.A1(new_n8516_), .A2(new_n8590_), .A3(new_n8578_), .A4(new_n8545_), .ZN(new_n8614_));
  NAND4_X1   g07599(.A1(new_n8607_), .A2(new_n8608_), .A3(new_n8589_), .A4(new_n8614_), .ZN(new_n8615_));
  NAND3_X1   g07600(.A1(new_n8615_), .A2(new_n8613_), .A3(new_n8593_), .ZN(new_n8616_));
  NAND3_X1   g07601(.A1(new_n8616_), .A2(new_n8610_), .A3(new_n8536_), .ZN(new_n8617_));
  NAND2_X1   g07602(.A1(new_n8617_), .A2(new_n8606_), .ZN(new_n8618_));
  NAND2_X1   g07603(.A1(new_n8596_), .A2(new_n8604_), .ZN(new_n8619_));
  OAI21_X1   g07604(.A1(new_n8609_), .A2(new_n8576_), .B(new_n8594_), .ZN(new_n8620_));
  AOI21_X1   g07605(.A1(new_n8620_), .A2(new_n8619_), .B(new_n8535_), .ZN(new_n8621_));
  NOR2_X1    g07606(.A1(new_n8596_), .A2(new_n8594_), .ZN(new_n8622_));
  NOR2_X1    g07607(.A1(new_n8582_), .A2(new_n8585_), .ZN(new_n8623_));
  NOR3_X1    g07608(.A1(new_n8600_), .A2(new_n8602_), .A3(new_n8598_), .ZN(new_n8624_));
  NAND2_X1   g07609(.A1(new_n8613_), .A2(new_n8593_), .ZN(new_n8625_));
  AOI21_X1   g07610(.A1(new_n8623_), .A2(new_n8624_), .B(new_n8625_), .ZN(new_n8626_));
  NOR3_X1    g07611(.A1(new_n8626_), .A2(new_n8622_), .A3(new_n8535_), .ZN(new_n8627_));
  NOR2_X1    g07612(.A1(new_n8600_), .A2(new_n8598_), .ZN(new_n8628_));
  NAND2_X1   g07613(.A1(new_n8591_), .A2(new_n8593_), .ZN(new_n8629_));
  NOR2_X1    g07614(.A1(new_n8628_), .A2(new_n8629_), .ZN(new_n8630_));
  NAND2_X1   g07615(.A1(new_n8589_), .A2(new_n8586_), .ZN(new_n8631_));
  NOR2_X1    g07616(.A1(new_n8603_), .A2(new_n8602_), .ZN(new_n8632_));
  NOR2_X1    g07617(.A1(new_n8631_), .A2(new_n8632_), .ZN(new_n8633_));
  NOR2_X1    g07618(.A1(new_n8633_), .A2(new_n8630_), .ZN(new_n8634_));
  INV_X1     g07619(.I(\A[855] ), .ZN(new_n8635_));
  NOR2_X1    g07620(.A1(new_n8635_), .A2(\A[854] ), .ZN(new_n8636_));
  INV_X1     g07621(.I(\A[854] ), .ZN(new_n8637_));
  NOR2_X1    g07622(.A1(new_n8637_), .A2(\A[855] ), .ZN(new_n8638_));
  OAI21_X1   g07623(.A1(new_n8636_), .A2(new_n8638_), .B(\A[853] ), .ZN(new_n8639_));
  INV_X1     g07624(.I(\A[853] ), .ZN(new_n8640_));
  NOR2_X1    g07625(.A1(\A[854] ), .A2(\A[855] ), .ZN(new_n8641_));
  NAND2_X1   g07626(.A1(\A[854] ), .A2(\A[855] ), .ZN(new_n8642_));
  INV_X1     g07627(.I(new_n8642_), .ZN(new_n8643_));
  OAI21_X1   g07628(.A1(new_n8643_), .A2(new_n8641_), .B(new_n8640_), .ZN(new_n8644_));
  NAND2_X1   g07629(.A1(new_n8639_), .A2(new_n8644_), .ZN(new_n8645_));
  INV_X1     g07630(.I(\A[858] ), .ZN(new_n8646_));
  NOR2_X1    g07631(.A1(new_n8646_), .A2(\A[857] ), .ZN(new_n8647_));
  INV_X1     g07632(.I(\A[857] ), .ZN(new_n8648_));
  NOR2_X1    g07633(.A1(new_n8648_), .A2(\A[858] ), .ZN(new_n8649_));
  OAI21_X1   g07634(.A1(new_n8647_), .A2(new_n8649_), .B(\A[856] ), .ZN(new_n8650_));
  INV_X1     g07635(.I(\A[856] ), .ZN(new_n8651_));
  NOR2_X1    g07636(.A1(\A[857] ), .A2(\A[858] ), .ZN(new_n8652_));
  NAND2_X1   g07637(.A1(\A[857] ), .A2(\A[858] ), .ZN(new_n8653_));
  INV_X1     g07638(.I(new_n8653_), .ZN(new_n8654_));
  OAI21_X1   g07639(.A1(new_n8654_), .A2(new_n8652_), .B(new_n8651_), .ZN(new_n8655_));
  NAND2_X1   g07640(.A1(new_n8650_), .A2(new_n8655_), .ZN(new_n8656_));
  AOI21_X1   g07641(.A1(new_n8651_), .A2(new_n8653_), .B(new_n8652_), .ZN(new_n8657_));
  AOI21_X1   g07642(.A1(new_n8640_), .A2(new_n8642_), .B(new_n8641_), .ZN(new_n8658_));
  NAND2_X1   g07643(.A1(new_n8657_), .A2(new_n8658_), .ZN(new_n8659_));
  NOR3_X1    g07644(.A1(new_n8645_), .A2(new_n8656_), .A3(new_n8659_), .ZN(new_n8660_));
  NOR2_X1    g07645(.A1(new_n8645_), .A2(new_n8656_), .ZN(new_n8661_));
  NAND2_X1   g07646(.A1(new_n8637_), .A2(\A[855] ), .ZN(new_n8662_));
  NAND2_X1   g07647(.A1(new_n8635_), .A2(\A[854] ), .ZN(new_n8663_));
  AOI21_X1   g07648(.A1(new_n8662_), .A2(new_n8663_), .B(new_n8640_), .ZN(new_n8664_));
  INV_X1     g07649(.I(new_n8641_), .ZN(new_n8665_));
  AOI21_X1   g07650(.A1(new_n8665_), .A2(new_n8642_), .B(\A[853] ), .ZN(new_n8666_));
  NOR2_X1    g07651(.A1(new_n8666_), .A2(new_n8664_), .ZN(new_n8667_));
  NAND2_X1   g07652(.A1(new_n8648_), .A2(\A[858] ), .ZN(new_n8668_));
  NAND2_X1   g07653(.A1(new_n8646_), .A2(\A[857] ), .ZN(new_n8669_));
  AOI21_X1   g07654(.A1(new_n8668_), .A2(new_n8669_), .B(new_n8651_), .ZN(new_n8670_));
  INV_X1     g07655(.I(new_n8652_), .ZN(new_n8671_));
  AOI21_X1   g07656(.A1(new_n8671_), .A2(new_n8653_), .B(\A[856] ), .ZN(new_n8672_));
  NOR2_X1    g07657(.A1(new_n8672_), .A2(new_n8670_), .ZN(new_n8673_));
  NOR2_X1    g07658(.A1(new_n8667_), .A2(new_n8673_), .ZN(new_n8674_));
  NOR2_X1    g07659(.A1(new_n8674_), .A2(new_n8661_), .ZN(new_n8675_));
  INV_X1     g07660(.I(\A[847] ), .ZN(new_n8676_));
  INV_X1     g07661(.I(\A[848] ), .ZN(new_n8677_));
  NAND2_X1   g07662(.A1(new_n8677_), .A2(\A[849] ), .ZN(new_n8678_));
  INV_X1     g07663(.I(\A[849] ), .ZN(new_n8679_));
  NAND2_X1   g07664(.A1(new_n8679_), .A2(\A[848] ), .ZN(new_n8680_));
  AOI21_X1   g07665(.A1(new_n8678_), .A2(new_n8680_), .B(new_n8676_), .ZN(new_n8681_));
  NOR2_X1    g07666(.A1(\A[848] ), .A2(\A[849] ), .ZN(new_n8682_));
  INV_X1     g07667(.I(new_n8682_), .ZN(new_n8683_));
  NAND2_X1   g07668(.A1(\A[848] ), .A2(\A[849] ), .ZN(new_n8684_));
  AOI21_X1   g07669(.A1(new_n8683_), .A2(new_n8684_), .B(\A[847] ), .ZN(new_n8685_));
  NOR2_X1    g07670(.A1(new_n8685_), .A2(new_n8681_), .ZN(new_n8686_));
  INV_X1     g07671(.I(\A[850] ), .ZN(new_n8687_));
  INV_X1     g07672(.I(\A[851] ), .ZN(new_n8688_));
  NAND2_X1   g07673(.A1(new_n8688_), .A2(\A[852] ), .ZN(new_n8689_));
  INV_X1     g07674(.I(\A[852] ), .ZN(new_n8690_));
  NAND2_X1   g07675(.A1(new_n8690_), .A2(\A[851] ), .ZN(new_n8691_));
  AOI21_X1   g07676(.A1(new_n8689_), .A2(new_n8691_), .B(new_n8687_), .ZN(new_n8692_));
  NOR2_X1    g07677(.A1(\A[851] ), .A2(\A[852] ), .ZN(new_n8693_));
  INV_X1     g07678(.I(new_n8693_), .ZN(new_n8694_));
  NAND2_X1   g07679(.A1(\A[851] ), .A2(\A[852] ), .ZN(new_n8695_));
  AOI21_X1   g07680(.A1(new_n8694_), .A2(new_n8695_), .B(\A[850] ), .ZN(new_n8696_));
  NOR2_X1    g07681(.A1(new_n8696_), .A2(new_n8692_), .ZN(new_n8697_));
  AOI21_X1   g07682(.A1(new_n8687_), .A2(new_n8695_), .B(new_n8693_), .ZN(new_n8698_));
  AOI21_X1   g07683(.A1(new_n8676_), .A2(new_n8684_), .B(new_n8682_), .ZN(new_n8699_));
  NAND2_X1   g07684(.A1(new_n8698_), .A2(new_n8699_), .ZN(new_n8700_));
  NAND2_X1   g07685(.A1(new_n8675_), .A2(new_n8660_), .ZN(new_n8702_));
  NAND2_X1   g07686(.A1(new_n8634_), .A2(new_n8702_), .ZN(new_n8703_));
  OAI21_X1   g07687(.A1(new_n8621_), .A2(new_n8627_), .B(new_n8703_), .ZN(new_n8704_));
  AND2_X2    g07688(.A1(new_n8675_), .A2(new_n8660_), .Z(new_n8705_));
  NOR3_X1    g07689(.A1(new_n8630_), .A2(new_n8633_), .A3(new_n8705_), .ZN(new_n8706_));
  NAND3_X1   g07690(.A1(new_n8617_), .A2(new_n8606_), .A3(new_n8706_), .ZN(new_n8707_));
  INV_X1     g07691(.I(new_n8659_), .ZN(new_n8708_));
  NAND3_X1   g07692(.A1(new_n8708_), .A2(new_n8667_), .A3(new_n8673_), .ZN(new_n8709_));
  NOR3_X1    g07693(.A1(new_n8709_), .A2(new_n8674_), .A3(new_n8661_), .ZN(new_n8710_));
  NOR4_X1    g07694(.A1(new_n8681_), .A2(new_n8685_), .A3(new_n8696_), .A4(new_n8692_), .ZN(new_n8711_));
  NOR2_X1    g07695(.A1(new_n8686_), .A2(new_n8697_), .ZN(new_n8712_));
  NOR2_X1    g07696(.A1(new_n8712_), .A2(new_n8711_), .ZN(new_n8713_));
  INV_X1     g07697(.I(new_n8658_), .ZN(new_n8714_));
  AOI21_X1   g07698(.A1(new_n8667_), .A2(new_n8673_), .B(new_n8714_), .ZN(new_n8715_));
  NOR3_X1    g07699(.A1(new_n8645_), .A2(new_n8656_), .A3(new_n8658_), .ZN(new_n8716_));
  OAI21_X1   g07700(.A1(new_n8715_), .A2(new_n8716_), .B(new_n8657_), .ZN(new_n8717_));
  INV_X1     g07701(.I(new_n8657_), .ZN(new_n8718_));
  OAI21_X1   g07702(.A1(new_n8645_), .A2(new_n8656_), .B(new_n8658_), .ZN(new_n8719_));
  NAND3_X1   g07703(.A1(new_n8667_), .A2(new_n8673_), .A3(new_n8714_), .ZN(new_n8720_));
  NAND3_X1   g07704(.A1(new_n8719_), .A2(new_n8720_), .A3(new_n8718_), .ZN(new_n8721_));
  NAND4_X1   g07705(.A1(new_n8710_), .A2(new_n8717_), .A3(new_n8721_), .A4(new_n8713_), .ZN(new_n8722_));
  NAND2_X1   g07706(.A1(new_n8686_), .A2(new_n8697_), .ZN(new_n8723_));
  NAND2_X1   g07707(.A1(new_n8667_), .A2(new_n8656_), .ZN(new_n8724_));
  NAND2_X1   g07708(.A1(new_n8673_), .A2(new_n8645_), .ZN(new_n8725_));
  AOI21_X1   g07709(.A1(new_n8724_), .A2(new_n8725_), .B(new_n8659_), .ZN(new_n8726_));
  NOR3_X1    g07710(.A1(new_n8726_), .A2(new_n8723_), .A3(new_n8700_), .ZN(new_n8727_));
  INV_X1     g07711(.I(new_n8699_), .ZN(new_n8728_));
  NOR2_X1    g07712(.A1(new_n8711_), .A2(new_n8728_), .ZN(new_n8729_));
  NOR2_X1    g07713(.A1(new_n8679_), .A2(\A[848] ), .ZN(new_n8730_));
  NOR2_X1    g07714(.A1(new_n8677_), .A2(\A[849] ), .ZN(new_n8731_));
  OAI21_X1   g07715(.A1(new_n8730_), .A2(new_n8731_), .B(\A[847] ), .ZN(new_n8732_));
  INV_X1     g07716(.I(new_n8684_), .ZN(new_n8733_));
  OAI21_X1   g07717(.A1(new_n8733_), .A2(new_n8682_), .B(new_n8676_), .ZN(new_n8734_));
  NAND2_X1   g07718(.A1(new_n8732_), .A2(new_n8734_), .ZN(new_n8735_));
  NOR2_X1    g07719(.A1(new_n8690_), .A2(\A[851] ), .ZN(new_n8736_));
  NOR2_X1    g07720(.A1(new_n8688_), .A2(\A[852] ), .ZN(new_n8737_));
  OAI21_X1   g07721(.A1(new_n8736_), .A2(new_n8737_), .B(\A[850] ), .ZN(new_n8738_));
  INV_X1     g07722(.I(new_n8695_), .ZN(new_n8739_));
  OAI21_X1   g07723(.A1(new_n8739_), .A2(new_n8693_), .B(new_n8687_), .ZN(new_n8740_));
  NAND2_X1   g07724(.A1(new_n8738_), .A2(new_n8740_), .ZN(new_n8741_));
  NOR3_X1    g07725(.A1(new_n8735_), .A2(new_n8741_), .A3(new_n8699_), .ZN(new_n8742_));
  OAI21_X1   g07726(.A1(new_n8729_), .A2(new_n8742_), .B(new_n8698_), .ZN(new_n8743_));
  INV_X1     g07727(.I(new_n8698_), .ZN(new_n8744_));
  OAI21_X1   g07728(.A1(new_n8735_), .A2(new_n8741_), .B(new_n8699_), .ZN(new_n8745_));
  NAND3_X1   g07729(.A1(new_n8686_), .A2(new_n8697_), .A3(new_n8728_), .ZN(new_n8746_));
  NAND3_X1   g07730(.A1(new_n8745_), .A2(new_n8746_), .A3(new_n8744_), .ZN(new_n8747_));
  NAND2_X1   g07731(.A1(new_n8743_), .A2(new_n8747_), .ZN(new_n8748_));
  NAND3_X1   g07732(.A1(new_n8722_), .A2(new_n8727_), .A3(new_n8748_), .ZN(new_n8749_));
  NOR3_X1    g07733(.A1(new_n8735_), .A2(new_n8741_), .A3(new_n8700_), .ZN(new_n8750_));
  NAND3_X1   g07734(.A1(new_n8710_), .A2(new_n8750_), .A3(new_n8713_), .ZN(new_n8751_));
  NAND2_X1   g07735(.A1(new_n8751_), .A2(new_n8748_), .ZN(new_n8752_));
  AOI21_X1   g07736(.A1(new_n8719_), .A2(new_n8720_), .B(new_n8718_), .ZN(new_n8753_));
  NOR3_X1    g07737(.A1(new_n8715_), .A2(new_n8716_), .A3(new_n8657_), .ZN(new_n8754_));
  NOR3_X1    g07738(.A1(new_n8754_), .A2(new_n8753_), .A3(new_n8726_), .ZN(new_n8755_));
  NAND2_X1   g07739(.A1(new_n8667_), .A2(new_n8673_), .ZN(new_n8756_));
  NAND2_X1   g07740(.A1(new_n8645_), .A2(new_n8656_), .ZN(new_n8757_));
  NAND3_X1   g07741(.A1(new_n8660_), .A2(new_n8756_), .A3(new_n8757_), .ZN(new_n8758_));
  NAND2_X1   g07742(.A1(new_n8735_), .A2(new_n8741_), .ZN(new_n8759_));
  NAND3_X1   g07743(.A1(new_n8750_), .A2(new_n8723_), .A3(new_n8759_), .ZN(new_n8760_));
  AOI21_X1   g07744(.A1(new_n8745_), .A2(new_n8746_), .B(new_n8744_), .ZN(new_n8761_));
  NOR3_X1    g07745(.A1(new_n8729_), .A2(new_n8742_), .A3(new_n8698_), .ZN(new_n8762_));
  NOR4_X1    g07746(.A1(new_n8762_), .A2(new_n8761_), .A3(new_n8758_), .A4(new_n8760_), .ZN(new_n8763_));
  NOR2_X1    g07747(.A1(new_n8763_), .A2(new_n8755_), .ZN(new_n8764_));
  NOR2_X1    g07748(.A1(new_n8673_), .A2(new_n8645_), .ZN(new_n8765_));
  NOR2_X1    g07749(.A1(new_n8667_), .A2(new_n8656_), .ZN(new_n8766_));
  OAI21_X1   g07750(.A1(new_n8765_), .A2(new_n8766_), .B(new_n8708_), .ZN(new_n8767_));
  NAND3_X1   g07751(.A1(new_n8717_), .A2(new_n8721_), .A3(new_n8767_), .ZN(new_n8768_));
  NOR3_X1    g07752(.A1(new_n8768_), .A2(new_n8751_), .A3(new_n8748_), .ZN(new_n8769_));
  OAI21_X1   g07753(.A1(new_n8764_), .A2(new_n8769_), .B(new_n8752_), .ZN(new_n8770_));
  NAND2_X1   g07754(.A1(new_n8770_), .A2(new_n8749_), .ZN(new_n8771_));
  AOI22_X1   g07755(.A1(new_n8704_), .A2(new_n8707_), .B1(new_n8771_), .B2(new_n8618_), .ZN(new_n8772_));
  NAND2_X1   g07756(.A1(new_n8610_), .A2(new_n8535_), .ZN(new_n8773_));
  NOR2_X1    g07757(.A1(new_n8540_), .A2(new_n8544_), .ZN(new_n8774_));
  OAI21_X1   g07758(.A1(new_n8578_), .A2(new_n8774_), .B(new_n8545_), .ZN(new_n8775_));
  NOR2_X1    g07759(.A1(new_n8496_), .A2(new_n8500_), .ZN(new_n8776_));
  OAI21_X1   g07760(.A1(new_n8528_), .A2(new_n8776_), .B(new_n8592_), .ZN(new_n8777_));
  XNOR2_X1   g07761(.A1(new_n8775_), .A2(new_n8777_), .ZN(new_n8778_));
  NAND3_X1   g07762(.A1(new_n8773_), .A2(new_n8778_), .A3(new_n8616_), .ZN(new_n8779_));
  NAND2_X1   g07763(.A1(new_n8722_), .A2(new_n8727_), .ZN(new_n8780_));
  OAI21_X1   g07764(.A1(new_n8755_), .A2(new_n8751_), .B(new_n8748_), .ZN(new_n8781_));
  NAND2_X1   g07765(.A1(new_n8718_), .A2(new_n8714_), .ZN(new_n8782_));
  AOI21_X1   g07766(.A1(new_n8661_), .A2(new_n8782_), .B(new_n8708_), .ZN(new_n8783_));
  NOR2_X1    g07767(.A1(new_n8698_), .A2(new_n8699_), .ZN(new_n8784_));
  OAI21_X1   g07768(.A1(new_n8723_), .A2(new_n8784_), .B(new_n8700_), .ZN(new_n8785_));
  XOR2_X1    g07769(.A1(new_n8783_), .A2(new_n8785_), .Z(new_n8786_));
  NAND3_X1   g07770(.A1(new_n8781_), .A2(new_n8780_), .A3(new_n8786_), .ZN(new_n8787_));
  XOR2_X1    g07771(.A1(new_n8779_), .A2(new_n8787_), .Z(new_n8788_));
  NAND2_X1   g07772(.A1(new_n8788_), .A2(new_n8772_), .ZN(new_n8789_));
  NOR2_X1    g07773(.A1(new_n8621_), .A2(new_n8627_), .ZN(new_n8790_));
  AOI21_X1   g07774(.A1(new_n8617_), .A2(new_n8606_), .B(new_n8706_), .ZN(new_n8791_));
  NOR3_X1    g07775(.A1(new_n8621_), .A2(new_n8627_), .A3(new_n8703_), .ZN(new_n8792_));
  INV_X1     g07776(.I(new_n8749_), .ZN(new_n8793_));
  OAI21_X1   g07777(.A1(new_n8748_), .A2(new_n8751_), .B(new_n8768_), .ZN(new_n8794_));
  NOR2_X1    g07778(.A1(new_n8762_), .A2(new_n8761_), .ZN(new_n8795_));
  NOR2_X1    g07779(.A1(new_n8758_), .A2(new_n8760_), .ZN(new_n8796_));
  NAND3_X1   g07780(.A1(new_n8755_), .A2(new_n8795_), .A3(new_n8796_), .ZN(new_n8797_));
  NAND2_X1   g07781(.A1(new_n8794_), .A2(new_n8797_), .ZN(new_n8798_));
  AOI21_X1   g07782(.A1(new_n8798_), .A2(new_n8752_), .B(new_n8793_), .ZN(new_n8799_));
  OAI22_X1   g07783(.A1(new_n8791_), .A2(new_n8792_), .B1(new_n8799_), .B2(new_n8790_), .ZN(new_n8800_));
  NAND2_X1   g07784(.A1(new_n8779_), .A2(new_n8787_), .ZN(new_n8801_));
  NOR2_X1    g07785(.A1(new_n8622_), .A2(new_n8536_), .ZN(new_n8802_));
  INV_X1     g07786(.I(new_n8778_), .ZN(new_n8803_));
  NOR3_X1    g07787(.A1(new_n8802_), .A2(new_n8626_), .A3(new_n8803_), .ZN(new_n8804_));
  INV_X1     g07788(.I(new_n8787_), .ZN(new_n8805_));
  NAND2_X1   g07789(.A1(new_n8805_), .A2(new_n8804_), .ZN(new_n8806_));
  NAND2_X1   g07790(.A1(new_n8806_), .A2(new_n8801_), .ZN(new_n8807_));
  NAND2_X1   g07791(.A1(new_n8807_), .A2(new_n8800_), .ZN(new_n8808_));
  NAND2_X1   g07792(.A1(new_n8789_), .A2(new_n8808_), .ZN(new_n8809_));
  INV_X1     g07793(.I(\A[886] ), .ZN(new_n8810_));
  NOR2_X1    g07794(.A1(\A[887] ), .A2(\A[888] ), .ZN(new_n8811_));
  NAND2_X1   g07795(.A1(\A[887] ), .A2(\A[888] ), .ZN(new_n8812_));
  AOI21_X1   g07796(.A1(new_n8810_), .A2(new_n8812_), .B(new_n8811_), .ZN(new_n8813_));
  INV_X1     g07797(.I(new_n8813_), .ZN(new_n8814_));
  INV_X1     g07798(.I(\A[883] ), .ZN(new_n8815_));
  NOR2_X1    g07799(.A1(\A[884] ), .A2(\A[885] ), .ZN(new_n8816_));
  NAND2_X1   g07800(.A1(\A[884] ), .A2(\A[885] ), .ZN(new_n8817_));
  AOI21_X1   g07801(.A1(new_n8815_), .A2(new_n8817_), .B(new_n8816_), .ZN(new_n8818_));
  INV_X1     g07802(.I(\A[885] ), .ZN(new_n8819_));
  NOR2_X1    g07803(.A1(new_n8819_), .A2(\A[884] ), .ZN(new_n8820_));
  INV_X1     g07804(.I(\A[884] ), .ZN(new_n8821_));
  NOR2_X1    g07805(.A1(new_n8821_), .A2(\A[885] ), .ZN(new_n8822_));
  OAI21_X1   g07806(.A1(new_n8820_), .A2(new_n8822_), .B(\A[883] ), .ZN(new_n8823_));
  INV_X1     g07807(.I(new_n8817_), .ZN(new_n8824_));
  OAI21_X1   g07808(.A1(new_n8824_), .A2(new_n8816_), .B(new_n8815_), .ZN(new_n8825_));
  INV_X1     g07809(.I(\A[888] ), .ZN(new_n8826_));
  NOR2_X1    g07810(.A1(new_n8826_), .A2(\A[887] ), .ZN(new_n8827_));
  INV_X1     g07811(.I(\A[887] ), .ZN(new_n8828_));
  NOR2_X1    g07812(.A1(new_n8828_), .A2(\A[888] ), .ZN(new_n8829_));
  OAI21_X1   g07813(.A1(new_n8827_), .A2(new_n8829_), .B(\A[886] ), .ZN(new_n8830_));
  INV_X1     g07814(.I(new_n8812_), .ZN(new_n8831_));
  OAI21_X1   g07815(.A1(new_n8831_), .A2(new_n8811_), .B(new_n8810_), .ZN(new_n8832_));
  NAND4_X1   g07816(.A1(new_n8823_), .A2(new_n8825_), .A3(new_n8830_), .A4(new_n8832_), .ZN(new_n8833_));
  NAND2_X1   g07817(.A1(new_n8833_), .A2(new_n8818_), .ZN(new_n8834_));
  INV_X1     g07818(.I(new_n8818_), .ZN(new_n8835_));
  NAND2_X1   g07819(.A1(new_n8821_), .A2(\A[885] ), .ZN(new_n8836_));
  NAND2_X1   g07820(.A1(new_n8819_), .A2(\A[884] ), .ZN(new_n8837_));
  AOI21_X1   g07821(.A1(new_n8836_), .A2(new_n8837_), .B(new_n8815_), .ZN(new_n8838_));
  INV_X1     g07822(.I(new_n8816_), .ZN(new_n8839_));
  AOI21_X1   g07823(.A1(new_n8839_), .A2(new_n8817_), .B(\A[883] ), .ZN(new_n8840_));
  NAND2_X1   g07824(.A1(new_n8828_), .A2(\A[888] ), .ZN(new_n8841_));
  NAND2_X1   g07825(.A1(new_n8826_), .A2(\A[887] ), .ZN(new_n8842_));
  AOI21_X1   g07826(.A1(new_n8841_), .A2(new_n8842_), .B(new_n8810_), .ZN(new_n8843_));
  INV_X1     g07827(.I(new_n8811_), .ZN(new_n8844_));
  AOI21_X1   g07828(.A1(new_n8844_), .A2(new_n8812_), .B(\A[886] ), .ZN(new_n8845_));
  NOR4_X1    g07829(.A1(new_n8838_), .A2(new_n8840_), .A3(new_n8845_), .A4(new_n8843_), .ZN(new_n8846_));
  NAND2_X1   g07830(.A1(new_n8846_), .A2(new_n8835_), .ZN(new_n8847_));
  AOI21_X1   g07831(.A1(new_n8847_), .A2(new_n8834_), .B(new_n8814_), .ZN(new_n8848_));
  NOR2_X1    g07832(.A1(new_n8846_), .A2(new_n8835_), .ZN(new_n8849_));
  NOR2_X1    g07833(.A1(new_n8833_), .A2(new_n8818_), .ZN(new_n8850_));
  NOR3_X1    g07834(.A1(new_n8849_), .A2(new_n8850_), .A3(new_n8813_), .ZN(new_n8851_));
  NOR2_X1    g07835(.A1(new_n8848_), .A2(new_n8851_), .ZN(new_n8852_));
  INV_X1     g07836(.I(\A[892] ), .ZN(new_n8853_));
  NOR2_X1    g07837(.A1(\A[893] ), .A2(\A[894] ), .ZN(new_n8854_));
  NAND2_X1   g07838(.A1(\A[893] ), .A2(\A[894] ), .ZN(new_n8855_));
  AOI21_X1   g07839(.A1(new_n8853_), .A2(new_n8855_), .B(new_n8854_), .ZN(new_n8856_));
  INV_X1     g07840(.I(\A[889] ), .ZN(new_n8857_));
  NOR2_X1    g07841(.A1(\A[890] ), .A2(\A[891] ), .ZN(new_n8858_));
  NAND2_X1   g07842(.A1(\A[890] ), .A2(\A[891] ), .ZN(new_n8859_));
  AOI21_X1   g07843(.A1(new_n8857_), .A2(new_n8859_), .B(new_n8858_), .ZN(new_n8860_));
  NAND2_X1   g07844(.A1(new_n8856_), .A2(new_n8860_), .ZN(new_n8861_));
  INV_X1     g07845(.I(\A[890] ), .ZN(new_n8862_));
  NAND2_X1   g07846(.A1(new_n8862_), .A2(\A[891] ), .ZN(new_n8863_));
  INV_X1     g07847(.I(\A[891] ), .ZN(new_n8864_));
  NAND2_X1   g07848(.A1(new_n8864_), .A2(\A[890] ), .ZN(new_n8865_));
  AOI21_X1   g07849(.A1(new_n8863_), .A2(new_n8865_), .B(new_n8857_), .ZN(new_n8866_));
  INV_X1     g07850(.I(new_n8858_), .ZN(new_n8867_));
  AOI21_X1   g07851(.A1(new_n8867_), .A2(new_n8859_), .B(\A[889] ), .ZN(new_n8868_));
  NOR2_X1    g07852(.A1(new_n8868_), .A2(new_n8866_), .ZN(new_n8869_));
  INV_X1     g07853(.I(\A[894] ), .ZN(new_n8870_));
  NOR2_X1    g07854(.A1(new_n8870_), .A2(\A[893] ), .ZN(new_n8871_));
  INV_X1     g07855(.I(\A[893] ), .ZN(new_n8872_));
  NOR2_X1    g07856(.A1(new_n8872_), .A2(\A[894] ), .ZN(new_n8873_));
  OAI21_X1   g07857(.A1(new_n8871_), .A2(new_n8873_), .B(\A[892] ), .ZN(new_n8874_));
  AND2_X2    g07858(.A1(\A[893] ), .A2(\A[894] ), .Z(new_n8875_));
  OAI21_X1   g07859(.A1(new_n8875_), .A2(new_n8854_), .B(new_n8853_), .ZN(new_n8876_));
  NAND2_X1   g07860(.A1(new_n8874_), .A2(new_n8876_), .ZN(new_n8877_));
  NAND2_X1   g07861(.A1(new_n8869_), .A2(new_n8877_), .ZN(new_n8878_));
  NOR2_X1    g07862(.A1(new_n8864_), .A2(\A[890] ), .ZN(new_n8879_));
  NOR2_X1    g07863(.A1(new_n8862_), .A2(\A[891] ), .ZN(new_n8880_));
  OAI21_X1   g07864(.A1(new_n8879_), .A2(new_n8880_), .B(\A[889] ), .ZN(new_n8881_));
  AND2_X2    g07865(.A1(\A[890] ), .A2(\A[891] ), .Z(new_n8882_));
  OAI21_X1   g07866(.A1(new_n8882_), .A2(new_n8858_), .B(new_n8857_), .ZN(new_n8883_));
  NAND2_X1   g07867(.A1(new_n8881_), .A2(new_n8883_), .ZN(new_n8884_));
  NAND2_X1   g07868(.A1(new_n8872_), .A2(\A[894] ), .ZN(new_n8885_));
  NAND2_X1   g07869(.A1(new_n8870_), .A2(\A[893] ), .ZN(new_n8886_));
  AOI21_X1   g07870(.A1(new_n8885_), .A2(new_n8886_), .B(new_n8853_), .ZN(new_n8887_));
  OR2_X2     g07871(.A1(\A[893] ), .A2(\A[894] ), .Z(new_n8888_));
  AOI21_X1   g07872(.A1(new_n8888_), .A2(new_n8855_), .B(\A[892] ), .ZN(new_n8889_));
  NOR2_X1    g07873(.A1(new_n8887_), .A2(new_n8889_), .ZN(new_n8890_));
  NAND2_X1   g07874(.A1(new_n8890_), .A2(new_n8884_), .ZN(new_n8891_));
  AOI21_X1   g07875(.A1(new_n8878_), .A2(new_n8891_), .B(new_n8861_), .ZN(new_n8892_));
  INV_X1     g07876(.I(new_n8856_), .ZN(new_n8893_));
  NAND4_X1   g07877(.A1(new_n8881_), .A2(new_n8874_), .A3(new_n8883_), .A4(new_n8876_), .ZN(new_n8894_));
  NAND2_X1   g07878(.A1(new_n8894_), .A2(new_n8860_), .ZN(new_n8895_));
  INV_X1     g07879(.I(new_n8860_), .ZN(new_n8896_));
  NAND3_X1   g07880(.A1(new_n8869_), .A2(new_n8890_), .A3(new_n8896_), .ZN(new_n8897_));
  AOI21_X1   g07881(.A1(new_n8895_), .A2(new_n8897_), .B(new_n8893_), .ZN(new_n8898_));
  AOI21_X1   g07882(.A1(new_n8869_), .A2(new_n8890_), .B(new_n8896_), .ZN(new_n8899_));
  NOR3_X1    g07883(.A1(new_n8884_), .A2(new_n8877_), .A3(new_n8860_), .ZN(new_n8900_));
  NOR3_X1    g07884(.A1(new_n8899_), .A2(new_n8900_), .A3(new_n8856_), .ZN(new_n8901_));
  NOR2_X1    g07885(.A1(new_n8894_), .A2(new_n8861_), .ZN(new_n8902_));
  NOR4_X1    g07886(.A1(new_n8866_), .A2(new_n8868_), .A3(new_n8887_), .A4(new_n8889_), .ZN(new_n8903_));
  AOI22_X1   g07887(.A1(new_n8881_), .A2(new_n8883_), .B1(new_n8874_), .B2(new_n8876_), .ZN(new_n8904_));
  NOR2_X1    g07888(.A1(new_n8904_), .A2(new_n8903_), .ZN(new_n8905_));
  AOI22_X1   g07889(.A1(new_n8823_), .A2(new_n8825_), .B1(new_n8830_), .B2(new_n8832_), .ZN(new_n8906_));
  NOR2_X1    g07890(.A1(new_n8906_), .A2(new_n8846_), .ZN(new_n8907_));
  NAND2_X1   g07891(.A1(new_n8813_), .A2(new_n8818_), .ZN(new_n8908_));
  NOR2_X1    g07892(.A1(new_n8833_), .A2(new_n8908_), .ZN(new_n8909_));
  NAND4_X1   g07893(.A1(new_n8907_), .A2(new_n8905_), .A3(new_n8909_), .A4(new_n8902_), .ZN(new_n8910_));
  NOR4_X1    g07894(.A1(new_n8910_), .A2(new_n8892_), .A3(new_n8898_), .A4(new_n8901_), .ZN(new_n8911_));
  NOR3_X1    g07895(.A1(new_n8898_), .A2(new_n8901_), .A3(new_n8892_), .ZN(new_n8912_));
  INV_X1     g07896(.I(new_n8861_), .ZN(new_n8913_));
  NAND2_X1   g07897(.A1(new_n8903_), .A2(new_n8913_), .ZN(new_n8914_));
  NAND2_X1   g07898(.A1(new_n8884_), .A2(new_n8877_), .ZN(new_n8915_));
  NAND2_X1   g07899(.A1(new_n8915_), .A2(new_n8894_), .ZN(new_n8916_));
  OAI22_X1   g07900(.A1(new_n8838_), .A2(new_n8840_), .B1(new_n8845_), .B2(new_n8843_), .ZN(new_n8917_));
  NAND2_X1   g07901(.A1(new_n8917_), .A2(new_n8833_), .ZN(new_n8918_));
  NAND3_X1   g07902(.A1(new_n8846_), .A2(new_n8813_), .A3(new_n8818_), .ZN(new_n8919_));
  NOR4_X1    g07903(.A1(new_n8916_), .A2(new_n8919_), .A3(new_n8918_), .A4(new_n8914_), .ZN(new_n8920_));
  NOR2_X1    g07904(.A1(new_n8912_), .A2(new_n8920_), .ZN(new_n8921_));
  OAI21_X1   g07905(.A1(new_n8921_), .A2(new_n8911_), .B(new_n8852_), .ZN(new_n8922_));
  OAI21_X1   g07906(.A1(new_n8899_), .A2(new_n8900_), .B(new_n8856_), .ZN(new_n8923_));
  NAND3_X1   g07907(.A1(new_n8895_), .A2(new_n8897_), .A3(new_n8893_), .ZN(new_n8924_));
  NAND2_X1   g07908(.A1(new_n8923_), .A2(new_n8924_), .ZN(new_n8925_));
  OAI21_X1   g07909(.A1(new_n8925_), .A2(new_n8892_), .B(new_n8920_), .ZN(new_n8926_));
  NAND3_X1   g07910(.A1(new_n8907_), .A2(new_n8905_), .A3(new_n8902_), .ZN(new_n8927_));
  NOR2_X1    g07911(.A1(new_n8892_), .A2(new_n8919_), .ZN(new_n8928_));
  OAI21_X1   g07912(.A1(new_n8925_), .A2(new_n8927_), .B(new_n8928_), .ZN(new_n8929_));
  NAND3_X1   g07913(.A1(new_n8926_), .A2(new_n8929_), .A3(new_n8852_), .ZN(new_n8930_));
  NAND2_X1   g07914(.A1(new_n8930_), .A2(new_n8922_), .ZN(new_n8931_));
  OR2_X2     g07915(.A1(new_n8848_), .A2(new_n8851_), .Z(new_n8932_));
  NAND2_X1   g07916(.A1(new_n8912_), .A2(new_n8920_), .ZN(new_n8933_));
  OAI21_X1   g07917(.A1(new_n8925_), .A2(new_n8892_), .B(new_n8910_), .ZN(new_n8934_));
  AOI21_X1   g07918(.A1(new_n8934_), .A2(new_n8933_), .B(new_n8932_), .ZN(new_n8935_));
  NOR2_X1    g07919(.A1(new_n8912_), .A2(new_n8910_), .ZN(new_n8936_));
  NOR2_X1    g07920(.A1(new_n8898_), .A2(new_n8901_), .ZN(new_n8937_));
  NOR3_X1    g07921(.A1(new_n8916_), .A2(new_n8918_), .A3(new_n8914_), .ZN(new_n8938_));
  NOR2_X1    g07922(.A1(new_n8890_), .A2(new_n8884_), .ZN(new_n8939_));
  NOR2_X1    g07923(.A1(new_n8869_), .A2(new_n8877_), .ZN(new_n8940_));
  OAI21_X1   g07924(.A1(new_n8939_), .A2(new_n8940_), .B(new_n8913_), .ZN(new_n8941_));
  NAND2_X1   g07925(.A1(new_n8941_), .A2(new_n8909_), .ZN(new_n8942_));
  AOI21_X1   g07926(.A1(new_n8937_), .A2(new_n8938_), .B(new_n8942_), .ZN(new_n8943_));
  NOR3_X1    g07927(.A1(new_n8943_), .A2(new_n8936_), .A3(new_n8932_), .ZN(new_n8944_));
  NOR2_X1    g07928(.A1(new_n8916_), .A2(new_n8914_), .ZN(new_n8945_));
  NAND2_X1   g07929(.A1(new_n8907_), .A2(new_n8909_), .ZN(new_n8946_));
  NOR2_X1    g07930(.A1(new_n8945_), .A2(new_n8946_), .ZN(new_n8947_));
  NAND2_X1   g07931(.A1(new_n8905_), .A2(new_n8902_), .ZN(new_n8948_));
  NOR2_X1    g07932(.A1(new_n8919_), .A2(new_n8918_), .ZN(new_n8949_));
  NOR2_X1    g07933(.A1(new_n8949_), .A2(new_n8948_), .ZN(new_n8950_));
  INV_X1     g07934(.I(\A[879] ), .ZN(new_n8951_));
  NOR2_X1    g07935(.A1(new_n8951_), .A2(\A[878] ), .ZN(new_n8952_));
  INV_X1     g07936(.I(\A[878] ), .ZN(new_n8953_));
  NOR2_X1    g07937(.A1(new_n8953_), .A2(\A[879] ), .ZN(new_n8954_));
  OAI21_X1   g07938(.A1(new_n8952_), .A2(new_n8954_), .B(\A[877] ), .ZN(new_n8955_));
  INV_X1     g07939(.I(\A[877] ), .ZN(new_n8956_));
  NOR2_X1    g07940(.A1(\A[878] ), .A2(\A[879] ), .ZN(new_n8957_));
  NAND2_X1   g07941(.A1(\A[878] ), .A2(\A[879] ), .ZN(new_n8958_));
  INV_X1     g07942(.I(new_n8958_), .ZN(new_n8959_));
  OAI21_X1   g07943(.A1(new_n8959_), .A2(new_n8957_), .B(new_n8956_), .ZN(new_n8960_));
  NAND2_X1   g07944(.A1(new_n8955_), .A2(new_n8960_), .ZN(new_n8961_));
  INV_X1     g07945(.I(\A[882] ), .ZN(new_n8962_));
  NOR2_X1    g07946(.A1(new_n8962_), .A2(\A[881] ), .ZN(new_n8963_));
  INV_X1     g07947(.I(\A[881] ), .ZN(new_n8964_));
  NOR2_X1    g07948(.A1(new_n8964_), .A2(\A[882] ), .ZN(new_n8965_));
  OAI21_X1   g07949(.A1(new_n8963_), .A2(new_n8965_), .B(\A[880] ), .ZN(new_n8966_));
  INV_X1     g07950(.I(\A[880] ), .ZN(new_n8967_));
  NOR2_X1    g07951(.A1(\A[881] ), .A2(\A[882] ), .ZN(new_n8968_));
  AND2_X2    g07952(.A1(\A[881] ), .A2(\A[882] ), .Z(new_n8969_));
  OAI21_X1   g07953(.A1(new_n8969_), .A2(new_n8968_), .B(new_n8967_), .ZN(new_n8970_));
  NAND2_X1   g07954(.A1(new_n8966_), .A2(new_n8970_), .ZN(new_n8971_));
  NAND2_X1   g07955(.A1(\A[881] ), .A2(\A[882] ), .ZN(new_n8972_));
  AOI21_X1   g07956(.A1(new_n8967_), .A2(new_n8972_), .B(new_n8968_), .ZN(new_n8973_));
  AOI21_X1   g07957(.A1(new_n8956_), .A2(new_n8958_), .B(new_n8957_), .ZN(new_n8974_));
  NAND2_X1   g07958(.A1(new_n8973_), .A2(new_n8974_), .ZN(new_n8975_));
  NOR3_X1    g07959(.A1(new_n8961_), .A2(new_n8971_), .A3(new_n8975_), .ZN(new_n8976_));
  NOR2_X1    g07960(.A1(new_n8961_), .A2(new_n8971_), .ZN(new_n8977_));
  NAND2_X1   g07961(.A1(new_n8953_), .A2(\A[879] ), .ZN(new_n8978_));
  NAND2_X1   g07962(.A1(new_n8951_), .A2(\A[878] ), .ZN(new_n8979_));
  AOI21_X1   g07963(.A1(new_n8978_), .A2(new_n8979_), .B(new_n8956_), .ZN(new_n8980_));
  INV_X1     g07964(.I(new_n8957_), .ZN(new_n8981_));
  AOI21_X1   g07965(.A1(new_n8981_), .A2(new_n8958_), .B(\A[877] ), .ZN(new_n8982_));
  NOR2_X1    g07966(.A1(new_n8982_), .A2(new_n8980_), .ZN(new_n8983_));
  NAND2_X1   g07967(.A1(new_n8964_), .A2(\A[882] ), .ZN(new_n8984_));
  NAND2_X1   g07968(.A1(new_n8962_), .A2(\A[881] ), .ZN(new_n8985_));
  AOI21_X1   g07969(.A1(new_n8984_), .A2(new_n8985_), .B(new_n8967_), .ZN(new_n8986_));
  OR2_X2     g07970(.A1(\A[881] ), .A2(\A[882] ), .Z(new_n8987_));
  AOI21_X1   g07971(.A1(new_n8987_), .A2(new_n8972_), .B(\A[880] ), .ZN(new_n8988_));
  NOR2_X1    g07972(.A1(new_n8986_), .A2(new_n8988_), .ZN(new_n8989_));
  NOR2_X1    g07973(.A1(new_n8983_), .A2(new_n8989_), .ZN(new_n8990_));
  NOR2_X1    g07974(.A1(new_n8990_), .A2(new_n8977_), .ZN(new_n8991_));
  INV_X1     g07975(.I(\A[871] ), .ZN(new_n8992_));
  INV_X1     g07976(.I(\A[872] ), .ZN(new_n8993_));
  NAND2_X1   g07977(.A1(new_n8993_), .A2(\A[873] ), .ZN(new_n8994_));
  INV_X1     g07978(.I(\A[873] ), .ZN(new_n8995_));
  NAND2_X1   g07979(.A1(new_n8995_), .A2(\A[872] ), .ZN(new_n8996_));
  AOI21_X1   g07980(.A1(new_n8994_), .A2(new_n8996_), .B(new_n8992_), .ZN(new_n8997_));
  NOR2_X1    g07981(.A1(\A[872] ), .A2(\A[873] ), .ZN(new_n8998_));
  INV_X1     g07982(.I(new_n8998_), .ZN(new_n8999_));
  NAND2_X1   g07983(.A1(\A[872] ), .A2(\A[873] ), .ZN(new_n9000_));
  AOI21_X1   g07984(.A1(new_n8999_), .A2(new_n9000_), .B(\A[871] ), .ZN(new_n9001_));
  NOR2_X1    g07985(.A1(new_n9001_), .A2(new_n8997_), .ZN(new_n9002_));
  INV_X1     g07986(.I(\A[874] ), .ZN(new_n9003_));
  INV_X1     g07987(.I(\A[875] ), .ZN(new_n9004_));
  NAND2_X1   g07988(.A1(new_n9004_), .A2(\A[876] ), .ZN(new_n9005_));
  INV_X1     g07989(.I(\A[876] ), .ZN(new_n9006_));
  NAND2_X1   g07990(.A1(new_n9006_), .A2(\A[875] ), .ZN(new_n9007_));
  AOI21_X1   g07991(.A1(new_n9005_), .A2(new_n9007_), .B(new_n9003_), .ZN(new_n9008_));
  OR2_X2     g07992(.A1(\A[875] ), .A2(\A[876] ), .Z(new_n9009_));
  NAND2_X1   g07993(.A1(\A[875] ), .A2(\A[876] ), .ZN(new_n9010_));
  AOI21_X1   g07994(.A1(new_n9009_), .A2(new_n9010_), .B(\A[874] ), .ZN(new_n9011_));
  NOR2_X1    g07995(.A1(new_n9008_), .A2(new_n9011_), .ZN(new_n9012_));
  NOR2_X1    g07996(.A1(\A[875] ), .A2(\A[876] ), .ZN(new_n9013_));
  AOI21_X1   g07997(.A1(new_n9003_), .A2(new_n9010_), .B(new_n9013_), .ZN(new_n9014_));
  AOI21_X1   g07998(.A1(new_n8992_), .A2(new_n9000_), .B(new_n8998_), .ZN(new_n9015_));
  NAND2_X1   g07999(.A1(new_n9014_), .A2(new_n9015_), .ZN(new_n9016_));
  AND2_X2    g08000(.A1(new_n8991_), .A2(new_n8976_), .Z(new_n9018_));
  NOR3_X1    g08001(.A1(new_n8947_), .A2(new_n9018_), .A3(new_n8950_), .ZN(new_n9019_));
  INV_X1     g08002(.I(new_n9019_), .ZN(new_n9020_));
  OAI21_X1   g08003(.A1(new_n8935_), .A2(new_n8944_), .B(new_n9020_), .ZN(new_n9021_));
  NAND3_X1   g08004(.A1(new_n8930_), .A2(new_n8922_), .A3(new_n9019_), .ZN(new_n9022_));
  NAND2_X1   g08005(.A1(new_n8983_), .A2(new_n8989_), .ZN(new_n9023_));
  NAND2_X1   g08006(.A1(new_n8961_), .A2(new_n8971_), .ZN(new_n9024_));
  NAND3_X1   g08007(.A1(new_n8976_), .A2(new_n9023_), .A3(new_n9024_), .ZN(new_n9025_));
  NAND2_X1   g08008(.A1(new_n9002_), .A2(new_n9012_), .ZN(new_n9026_));
  NOR2_X1    g08009(.A1(new_n8995_), .A2(\A[872] ), .ZN(new_n9027_));
  NOR2_X1    g08010(.A1(new_n8993_), .A2(\A[873] ), .ZN(new_n9028_));
  OAI21_X1   g08011(.A1(new_n9027_), .A2(new_n9028_), .B(\A[871] ), .ZN(new_n9029_));
  INV_X1     g08012(.I(new_n9000_), .ZN(new_n9030_));
  OAI21_X1   g08013(.A1(new_n9030_), .A2(new_n8998_), .B(new_n8992_), .ZN(new_n9031_));
  NAND2_X1   g08014(.A1(new_n9029_), .A2(new_n9031_), .ZN(new_n9032_));
  NOR2_X1    g08015(.A1(new_n9006_), .A2(\A[875] ), .ZN(new_n9033_));
  NOR2_X1    g08016(.A1(new_n9004_), .A2(\A[876] ), .ZN(new_n9034_));
  OAI21_X1   g08017(.A1(new_n9033_), .A2(new_n9034_), .B(\A[874] ), .ZN(new_n9035_));
  AND2_X2    g08018(.A1(\A[875] ), .A2(\A[876] ), .Z(new_n9036_));
  OAI21_X1   g08019(.A1(new_n9036_), .A2(new_n9013_), .B(new_n9003_), .ZN(new_n9037_));
  NAND2_X1   g08020(.A1(new_n9035_), .A2(new_n9037_), .ZN(new_n9038_));
  NAND2_X1   g08021(.A1(new_n9032_), .A2(new_n9038_), .ZN(new_n9039_));
  NAND2_X1   g08022(.A1(new_n9026_), .A2(new_n9039_), .ZN(new_n9040_));
  INV_X1     g08023(.I(new_n8973_), .ZN(new_n9041_));
  OAI21_X1   g08024(.A1(new_n8961_), .A2(new_n8971_), .B(new_n8974_), .ZN(new_n9042_));
  INV_X1     g08025(.I(new_n8974_), .ZN(new_n9043_));
  NAND3_X1   g08026(.A1(new_n8983_), .A2(new_n8989_), .A3(new_n9043_), .ZN(new_n9044_));
  AOI21_X1   g08027(.A1(new_n9042_), .A2(new_n9044_), .B(new_n9041_), .ZN(new_n9045_));
  AOI21_X1   g08028(.A1(new_n8983_), .A2(new_n8989_), .B(new_n9043_), .ZN(new_n9046_));
  NOR3_X1    g08029(.A1(new_n8961_), .A2(new_n8971_), .A3(new_n8974_), .ZN(new_n9047_));
  NOR3_X1    g08030(.A1(new_n9046_), .A2(new_n9047_), .A3(new_n8973_), .ZN(new_n9048_));
  NOR4_X1    g08031(.A1(new_n9045_), .A2(new_n9048_), .A3(new_n9025_), .A4(new_n9040_), .ZN(new_n9049_));
  NOR3_X1    g08032(.A1(new_n9032_), .A2(new_n9038_), .A3(new_n9016_), .ZN(new_n9050_));
  INV_X1     g08033(.I(new_n8975_), .ZN(new_n9051_));
  NOR2_X1    g08034(.A1(new_n8961_), .A2(new_n8989_), .ZN(new_n9052_));
  NOR2_X1    g08035(.A1(new_n8983_), .A2(new_n8971_), .ZN(new_n9053_));
  OAI21_X1   g08036(.A1(new_n9052_), .A2(new_n9053_), .B(new_n9051_), .ZN(new_n9054_));
  NAND2_X1   g08037(.A1(new_n9054_), .A2(new_n9050_), .ZN(new_n9055_));
  INV_X1     g08038(.I(new_n9014_), .ZN(new_n9056_));
  OAI21_X1   g08039(.A1(new_n9032_), .A2(new_n9038_), .B(new_n9015_), .ZN(new_n9057_));
  INV_X1     g08040(.I(new_n9015_), .ZN(new_n9058_));
  NAND3_X1   g08041(.A1(new_n9002_), .A2(new_n9012_), .A3(new_n9058_), .ZN(new_n9059_));
  AOI21_X1   g08042(.A1(new_n9057_), .A2(new_n9059_), .B(new_n9056_), .ZN(new_n9060_));
  NOR4_X1    g08043(.A1(new_n8997_), .A2(new_n9001_), .A3(new_n9008_), .A4(new_n9011_), .ZN(new_n9061_));
  NOR2_X1    g08044(.A1(new_n9061_), .A2(new_n9058_), .ZN(new_n9062_));
  NOR3_X1    g08045(.A1(new_n9032_), .A2(new_n9038_), .A3(new_n9015_), .ZN(new_n9063_));
  NOR3_X1    g08046(.A1(new_n9062_), .A2(new_n9014_), .A3(new_n9063_), .ZN(new_n9064_));
  NOR2_X1    g08047(.A1(new_n9064_), .A2(new_n9060_), .ZN(new_n9065_));
  NOR3_X1    g08048(.A1(new_n9049_), .A2(new_n9055_), .A3(new_n9065_), .ZN(new_n9066_));
  INV_X1     g08049(.I(new_n9066_), .ZN(new_n9067_));
  OAI21_X1   g08050(.A1(new_n9062_), .A2(new_n9063_), .B(new_n9014_), .ZN(new_n9068_));
  NAND3_X1   g08051(.A1(new_n9057_), .A2(new_n9059_), .A3(new_n9056_), .ZN(new_n9069_));
  NAND2_X1   g08052(.A1(new_n9068_), .A2(new_n9069_), .ZN(new_n9070_));
  NOR2_X1    g08053(.A1(new_n9002_), .A2(new_n9012_), .ZN(new_n9071_));
  NOR2_X1    g08054(.A1(new_n9071_), .A2(new_n9061_), .ZN(new_n9072_));
  NAND4_X1   g08055(.A1(new_n8991_), .A2(new_n9072_), .A3(new_n8976_), .A4(new_n9050_), .ZN(new_n9073_));
  NAND2_X1   g08056(.A1(new_n9070_), .A2(new_n9073_), .ZN(new_n9074_));
  NAND2_X1   g08057(.A1(new_n8983_), .A2(new_n8971_), .ZN(new_n9075_));
  NAND2_X1   g08058(.A1(new_n8961_), .A2(new_n8989_), .ZN(new_n9076_));
  AOI21_X1   g08059(.A1(new_n9076_), .A2(new_n9075_), .B(new_n8975_), .ZN(new_n9077_));
  NOR3_X1    g08060(.A1(new_n9045_), .A2(new_n9048_), .A3(new_n9077_), .ZN(new_n9078_));
  NAND3_X1   g08061(.A1(new_n9050_), .A2(new_n9026_), .A3(new_n9039_), .ZN(new_n9079_));
  NOR4_X1    g08062(.A1(new_n9025_), .A2(new_n9064_), .A3(new_n9060_), .A4(new_n9079_), .ZN(new_n9080_));
  NOR2_X1    g08063(.A1(new_n9080_), .A2(new_n9078_), .ZN(new_n9081_));
  OAI21_X1   g08064(.A1(new_n9046_), .A2(new_n9047_), .B(new_n8973_), .ZN(new_n9082_));
  NAND3_X1   g08065(.A1(new_n9042_), .A2(new_n9044_), .A3(new_n9041_), .ZN(new_n9083_));
  NAND3_X1   g08066(.A1(new_n9082_), .A2(new_n9083_), .A3(new_n9054_), .ZN(new_n9084_));
  NOR3_X1    g08067(.A1(new_n9084_), .A2(new_n9070_), .A3(new_n9073_), .ZN(new_n9085_));
  OAI21_X1   g08068(.A1(new_n9081_), .A2(new_n9085_), .B(new_n9074_), .ZN(new_n9086_));
  NAND2_X1   g08069(.A1(new_n9086_), .A2(new_n9067_), .ZN(new_n9087_));
  AOI22_X1   g08070(.A1(new_n9021_), .A2(new_n9022_), .B1(new_n9087_), .B2(new_n8931_), .ZN(new_n9088_));
  NOR2_X1    g08071(.A1(new_n8936_), .A2(new_n8852_), .ZN(new_n9089_));
  NOR2_X1    g08072(.A1(new_n8856_), .A2(new_n8860_), .ZN(new_n9090_));
  OAI21_X1   g08073(.A1(new_n8894_), .A2(new_n9090_), .B(new_n8861_), .ZN(new_n9091_));
  NOR2_X1    g08074(.A1(new_n8813_), .A2(new_n8818_), .ZN(new_n9092_));
  OAI21_X1   g08075(.A1(new_n8833_), .A2(new_n9092_), .B(new_n8908_), .ZN(new_n9093_));
  XNOR2_X1   g08076(.A1(new_n9093_), .A2(new_n9091_), .ZN(new_n9094_));
  INV_X1     g08077(.I(new_n9094_), .ZN(new_n9095_));
  NOR3_X1    g08078(.A1(new_n9089_), .A2(new_n9095_), .A3(new_n8943_), .ZN(new_n9096_));
  NOR2_X1    g08079(.A1(new_n9049_), .A2(new_n9055_), .ZN(new_n9097_));
  NOR2_X1    g08080(.A1(new_n9025_), .A2(new_n9079_), .ZN(new_n9098_));
  AOI21_X1   g08081(.A1(new_n9084_), .A2(new_n9098_), .B(new_n9065_), .ZN(new_n9099_));
  NOR2_X1    g08082(.A1(new_n8973_), .A2(new_n8974_), .ZN(new_n9100_));
  OAI21_X1   g08083(.A1(new_n9023_), .A2(new_n9100_), .B(new_n8975_), .ZN(new_n9101_));
  NOR2_X1    g08084(.A1(new_n9014_), .A2(new_n9015_), .ZN(new_n9102_));
  OAI21_X1   g08085(.A1(new_n9026_), .A2(new_n9102_), .B(new_n9016_), .ZN(new_n9103_));
  XOR2_X1    g08086(.A1(new_n9101_), .A2(new_n9103_), .Z(new_n9104_));
  NOR3_X1    g08087(.A1(new_n9099_), .A2(new_n9097_), .A3(new_n9104_), .ZN(new_n9105_));
  XOR2_X1    g08088(.A1(new_n9096_), .A2(new_n9105_), .Z(new_n9106_));
  NAND2_X1   g08089(.A1(new_n9106_), .A2(new_n9088_), .ZN(new_n9107_));
  NOR2_X1    g08090(.A1(new_n8935_), .A2(new_n8944_), .ZN(new_n9108_));
  AOI21_X1   g08091(.A1(new_n8930_), .A2(new_n8922_), .B(new_n9019_), .ZN(new_n9109_));
  NOR3_X1    g08092(.A1(new_n8935_), .A2(new_n8944_), .A3(new_n9020_), .ZN(new_n9110_));
  OAI21_X1   g08093(.A1(new_n9070_), .A2(new_n9073_), .B(new_n9084_), .ZN(new_n9111_));
  NAND3_X1   g08094(.A1(new_n9078_), .A2(new_n9065_), .A3(new_n9098_), .ZN(new_n9112_));
  NAND2_X1   g08095(.A1(new_n9111_), .A2(new_n9112_), .ZN(new_n9113_));
  AOI21_X1   g08096(.A1(new_n9113_), .A2(new_n9074_), .B(new_n9066_), .ZN(new_n9114_));
  OAI22_X1   g08097(.A1(new_n9110_), .A2(new_n9109_), .B1(new_n9114_), .B2(new_n9108_), .ZN(new_n9115_));
  NAND2_X1   g08098(.A1(new_n8926_), .A2(new_n8932_), .ZN(new_n9116_));
  NAND3_X1   g08099(.A1(new_n9116_), .A2(new_n9094_), .A3(new_n8929_), .ZN(new_n9117_));
  INV_X1     g08100(.I(new_n9105_), .ZN(new_n9118_));
  NAND2_X1   g08101(.A1(new_n9118_), .A2(new_n9117_), .ZN(new_n9119_));
  INV_X1     g08102(.I(new_n9119_), .ZN(new_n9120_));
  NOR2_X1    g08103(.A1(new_n9118_), .A2(new_n9117_), .ZN(new_n9121_));
  OAI21_X1   g08104(.A1(new_n9120_), .A2(new_n9121_), .B(new_n9115_), .ZN(new_n9122_));
  NAND2_X1   g08105(.A1(new_n9122_), .A2(new_n9107_), .ZN(new_n9123_));
  NOR2_X1    g08106(.A1(new_n9123_), .A2(new_n8809_), .ZN(new_n9124_));
  NOR3_X1    g08107(.A1(new_n9110_), .A2(new_n9109_), .A3(new_n9087_), .ZN(new_n9125_));
  NOR2_X1    g08108(.A1(new_n8947_), .A2(new_n8950_), .ZN(new_n9126_));
  NOR2_X1    g08109(.A1(new_n9126_), .A2(new_n9025_), .ZN(new_n9127_));
  NOR2_X1    g08110(.A1(new_n9127_), .A2(new_n9019_), .ZN(new_n9128_));
  NOR2_X1    g08111(.A1(new_n8634_), .A2(new_n8702_), .ZN(new_n9129_));
  NOR2_X1    g08112(.A1(new_n9129_), .A2(new_n8706_), .ZN(new_n9130_));
  NAND2_X1   g08113(.A1(new_n9130_), .A2(new_n9128_), .ZN(new_n9131_));
  INV_X1     g08114(.I(new_n9131_), .ZN(new_n9132_));
  NOR2_X1    g08115(.A1(new_n9132_), .A2(new_n9125_), .ZN(new_n9133_));
  INV_X1     g08116(.I(new_n9125_), .ZN(new_n9134_));
  NOR2_X1    g08117(.A1(new_n9134_), .A2(new_n9131_), .ZN(new_n9135_));
  OAI21_X1   g08118(.A1(new_n8792_), .A2(new_n8791_), .B(new_n8799_), .ZN(new_n9136_));
  NAND3_X1   g08119(.A1(new_n8704_), .A2(new_n8771_), .A3(new_n8707_), .ZN(new_n9137_));
  NAND2_X1   g08120(.A1(new_n9136_), .A2(new_n9137_), .ZN(new_n9138_));
  INV_X1     g08121(.I(new_n9138_), .ZN(new_n9139_));
  OAI22_X1   g08122(.A1(new_n9139_), .A2(new_n9125_), .B1(new_n9135_), .B2(new_n9133_), .ZN(new_n9140_));
  INV_X1     g08123(.I(new_n9140_), .ZN(new_n9141_));
  NAND2_X1   g08124(.A1(new_n9123_), .A2(new_n8809_), .ZN(new_n9142_));
  AOI21_X1   g08125(.A1(new_n9141_), .A2(new_n9142_), .B(new_n9124_), .ZN(new_n9143_));
  NAND2_X1   g08126(.A1(new_n8775_), .A2(new_n8777_), .ZN(new_n9144_));
  NOR2_X1    g08127(.A1(new_n8802_), .A2(new_n8626_), .ZN(new_n9145_));
  OAI21_X1   g08128(.A1(new_n8775_), .A2(new_n8777_), .B(new_n9145_), .ZN(new_n9146_));
  NAND2_X1   g08129(.A1(new_n9146_), .A2(new_n9144_), .ZN(new_n9147_));
  AND2_X2    g08130(.A1(new_n8781_), .A2(new_n8780_), .Z(new_n9148_));
  INV_X1     g08131(.I(new_n8783_), .ZN(new_n9149_));
  NAND2_X1   g08132(.A1(new_n9149_), .A2(new_n8785_), .ZN(new_n9150_));
  INV_X1     g08133(.I(new_n9150_), .ZN(new_n9151_));
  OR2_X2     g08134(.A1(new_n9149_), .A2(new_n8785_), .Z(new_n9152_));
  AOI21_X1   g08135(.A1(new_n9148_), .A2(new_n9152_), .B(new_n9151_), .ZN(new_n9153_));
  AOI21_X1   g08136(.A1(new_n8800_), .A2(new_n8801_), .B(new_n8806_), .ZN(new_n9154_));
  NOR2_X1    g08137(.A1(new_n9154_), .A2(new_n9153_), .ZN(new_n9155_));
  NAND4_X1   g08138(.A1(new_n8772_), .A2(new_n8804_), .A3(new_n8805_), .A4(new_n9153_), .ZN(new_n9156_));
  INV_X1     g08139(.I(new_n9156_), .ZN(new_n9157_));
  OAI21_X1   g08140(.A1(new_n9155_), .A2(new_n9157_), .B(new_n9147_), .ZN(new_n9158_));
  INV_X1     g08141(.I(new_n9147_), .ZN(new_n9159_));
  INV_X1     g08142(.I(new_n9153_), .ZN(new_n9160_));
  NAND3_X1   g08143(.A1(new_n8772_), .A2(new_n8804_), .A3(new_n8805_), .ZN(new_n9161_));
  NAND2_X1   g08144(.A1(new_n9161_), .A2(new_n9160_), .ZN(new_n9162_));
  NAND3_X1   g08145(.A1(new_n9162_), .A2(new_n9159_), .A3(new_n9156_), .ZN(new_n9163_));
  NAND2_X1   g08146(.A1(new_n9158_), .A2(new_n9163_), .ZN(new_n9164_));
  NAND2_X1   g08147(.A1(new_n9093_), .A2(new_n9091_), .ZN(new_n9165_));
  NOR2_X1    g08148(.A1(new_n9089_), .A2(new_n8943_), .ZN(new_n9166_));
  OAI21_X1   g08149(.A1(new_n9091_), .A2(new_n9093_), .B(new_n9166_), .ZN(new_n9167_));
  NAND2_X1   g08150(.A1(new_n9167_), .A2(new_n9165_), .ZN(new_n9168_));
  INV_X1     g08151(.I(new_n9168_), .ZN(new_n9169_));
  NAND2_X1   g08152(.A1(new_n9101_), .A2(new_n9103_), .ZN(new_n9170_));
  NOR2_X1    g08153(.A1(new_n9101_), .A2(new_n9103_), .ZN(new_n9171_));
  OR3_X2     g08154(.A1(new_n9099_), .A2(new_n9097_), .A3(new_n9171_), .Z(new_n9172_));
  NAND2_X1   g08155(.A1(new_n9172_), .A2(new_n9170_), .ZN(new_n9173_));
  NAND3_X1   g08156(.A1(new_n9088_), .A2(new_n9096_), .A3(new_n9105_), .ZN(new_n9174_));
  NAND2_X1   g08157(.A1(new_n9174_), .A2(new_n9173_), .ZN(new_n9175_));
  INV_X1     g08158(.I(new_n9173_), .ZN(new_n9176_));
  NAND4_X1   g08159(.A1(new_n9088_), .A2(new_n9176_), .A3(new_n9096_), .A4(new_n9105_), .ZN(new_n9177_));
  AOI21_X1   g08160(.A1(new_n9175_), .A2(new_n9177_), .B(new_n9169_), .ZN(new_n9178_));
  NAND2_X1   g08161(.A1(new_n9108_), .A2(new_n9019_), .ZN(new_n9179_));
  OAI21_X1   g08162(.A1(new_n9110_), .A2(new_n9109_), .B(new_n9114_), .ZN(new_n9180_));
  NAND3_X1   g08163(.A1(new_n9180_), .A2(new_n9179_), .A3(new_n9119_), .ZN(new_n9181_));
  AOI21_X1   g08164(.A1(new_n9181_), .A2(new_n9121_), .B(new_n9176_), .ZN(new_n9182_));
  NOR4_X1    g08165(.A1(new_n9115_), .A2(new_n9173_), .A3(new_n9117_), .A4(new_n9118_), .ZN(new_n9183_));
  NOR3_X1    g08166(.A1(new_n9182_), .A2(new_n9168_), .A3(new_n9183_), .ZN(new_n9184_));
  NOR2_X1    g08167(.A1(new_n9184_), .A2(new_n9178_), .ZN(new_n9185_));
  NAND2_X1   g08168(.A1(new_n9164_), .A2(new_n9185_), .ZN(new_n9186_));
  OAI21_X1   g08169(.A1(new_n9182_), .A2(new_n9183_), .B(new_n9168_), .ZN(new_n9187_));
  NAND3_X1   g08170(.A1(new_n9175_), .A2(new_n9169_), .A3(new_n9177_), .ZN(new_n9188_));
  NAND2_X1   g08171(.A1(new_n9187_), .A2(new_n9188_), .ZN(new_n9189_));
  NAND3_X1   g08172(.A1(new_n9189_), .A2(new_n9158_), .A3(new_n9163_), .ZN(new_n9190_));
  AOI21_X1   g08173(.A1(new_n9186_), .A2(new_n9190_), .B(new_n9143_), .ZN(new_n9191_));
  NAND4_X1   g08174(.A1(new_n8789_), .A2(new_n9122_), .A3(new_n9107_), .A4(new_n8808_), .ZN(new_n9192_));
  AOI22_X1   g08175(.A1(new_n9107_), .A2(new_n9122_), .B1(new_n8789_), .B2(new_n8808_), .ZN(new_n9193_));
  OAI21_X1   g08176(.A1(new_n9140_), .A2(new_n9193_), .B(new_n9192_), .ZN(new_n9194_));
  NAND4_X1   g08177(.A1(new_n9158_), .A2(new_n9163_), .A3(new_n9187_), .A4(new_n9188_), .ZN(new_n9195_));
  AOI21_X1   g08178(.A1(new_n9162_), .A2(new_n9156_), .B(new_n9159_), .ZN(new_n9196_));
  NOR3_X1    g08179(.A1(new_n9155_), .A2(new_n9157_), .A3(new_n9147_), .ZN(new_n9197_));
  OAI22_X1   g08180(.A1(new_n9197_), .A2(new_n9196_), .B1(new_n9184_), .B2(new_n9178_), .ZN(new_n9198_));
  AOI21_X1   g08181(.A1(new_n9198_), .A2(new_n9195_), .B(new_n9194_), .ZN(new_n9199_));
  NOR4_X1    g08182(.A1(new_n8484_), .A2(new_n9191_), .A3(new_n8492_), .A4(new_n9199_), .ZN(new_n9200_));
  INV_X1     g08183(.I(new_n9123_), .ZN(new_n9201_));
  NOR2_X1    g08184(.A1(new_n9201_), .A2(new_n8809_), .ZN(new_n9202_));
  AND2_X2    g08185(.A1(new_n8789_), .A2(new_n8808_), .Z(new_n9203_));
  NOR2_X1    g08186(.A1(new_n9203_), .A2(new_n9123_), .ZN(new_n9204_));
  OAI21_X1   g08187(.A1(new_n9202_), .A2(new_n9204_), .B(new_n9141_), .ZN(new_n9205_));
  OAI21_X1   g08188(.A1(new_n9124_), .A2(new_n9193_), .B(new_n9140_), .ZN(new_n9206_));
  NOR2_X1    g08189(.A1(new_n8414_), .A2(new_n8410_), .ZN(new_n9207_));
  NOR2_X1    g08190(.A1(new_n9207_), .A2(new_n8383_), .ZN(new_n9208_));
  AOI21_X1   g08191(.A1(new_n8383_), .A2(new_n8400_), .B(new_n9208_), .ZN(new_n9209_));
  NOR2_X1    g08192(.A1(new_n9209_), .A2(new_n8105_), .ZN(new_n9210_));
  XOR2_X1    g08193(.A1(new_n8099_), .A2(new_n8087_), .Z(new_n9211_));
  NOR2_X1    g08194(.A1(new_n9211_), .A2(new_n8097_), .ZN(new_n9212_));
  AOI21_X1   g08195(.A1(new_n8097_), .A2(new_n8103_), .B(new_n9212_), .ZN(new_n9213_));
  NOR2_X1    g08196(.A1(new_n9213_), .A2(new_n8416_), .ZN(new_n9214_));
  OAI21_X1   g08197(.A1(new_n9214_), .A2(new_n9210_), .B(new_n8431_), .ZN(new_n9215_));
  OAI21_X1   g08198(.A1(new_n8417_), .A2(new_n8432_), .B(new_n8488_), .ZN(new_n9216_));
  NAND4_X1   g08199(.A1(new_n9205_), .A2(new_n9215_), .A3(new_n9216_), .A4(new_n9206_), .ZN(new_n9217_));
  NOR3_X1    g08200(.A1(new_n8486_), .A2(new_n8425_), .A3(new_n8430_), .ZN(new_n9218_));
  INV_X1     g08201(.I(new_n9218_), .ZN(new_n9219_));
  NAND2_X1   g08202(.A1(new_n8315_), .A2(new_n8420_), .ZN(new_n9220_));
  OAI21_X1   g08203(.A1(new_n8005_), .A2(new_n8421_), .B(new_n9220_), .ZN(new_n9221_));
  NOR2_X1    g08204(.A1(new_n9130_), .A2(new_n9128_), .ZN(new_n9222_));
  NOR2_X1    g08205(.A1(new_n9132_), .A2(new_n9222_), .ZN(new_n9223_));
  NAND3_X1   g08206(.A1(new_n9223_), .A2(new_n8423_), .A3(new_n9221_), .ZN(new_n9224_));
  NAND2_X1   g08207(.A1(new_n9219_), .A2(new_n9224_), .ZN(new_n9225_));
  INV_X1     g08208(.I(new_n9224_), .ZN(new_n9226_));
  NAND2_X1   g08209(.A1(new_n9218_), .A2(new_n9226_), .ZN(new_n9227_));
  NAND2_X1   g08210(.A1(new_n9225_), .A2(new_n9227_), .ZN(new_n9228_));
  NOR2_X1    g08211(.A1(new_n9219_), .A2(new_n9224_), .ZN(new_n9229_));
  INV_X1     g08212(.I(new_n9133_), .ZN(new_n9230_));
  INV_X1     g08213(.I(new_n9135_), .ZN(new_n9231_));
  AOI21_X1   g08214(.A1(new_n9231_), .A2(new_n9230_), .B(new_n9138_), .ZN(new_n9232_));
  NOR3_X1    g08215(.A1(new_n9139_), .A2(new_n9135_), .A3(new_n9133_), .ZN(new_n9233_));
  NOR2_X1    g08216(.A1(new_n9232_), .A2(new_n9233_), .ZN(new_n9234_));
  AOI21_X1   g08217(.A1(new_n9228_), .A2(new_n9234_), .B(new_n9229_), .ZN(new_n9235_));
  AOI22_X1   g08218(.A1(new_n9205_), .A2(new_n9206_), .B1(new_n9215_), .B2(new_n9216_), .ZN(new_n9236_));
  OAI21_X1   g08219(.A1(new_n9236_), .A2(new_n9235_), .B(new_n9217_), .ZN(new_n9237_));
  OAI22_X1   g08220(.A1(new_n8484_), .A2(new_n8492_), .B1(new_n9191_), .B2(new_n9199_), .ZN(new_n9238_));
  AOI21_X1   g08221(.A1(new_n9238_), .A2(new_n9237_), .B(new_n9200_), .ZN(new_n9239_));
  NAND2_X1   g08222(.A1(new_n8459_), .A2(new_n8467_), .ZN(new_n9240_));
  NAND2_X1   g08223(.A1(new_n8458_), .A2(new_n8464_), .ZN(new_n9241_));
  NAND3_X1   g08224(.A1(new_n9241_), .A2(new_n8471_), .A3(new_n8414_), .ZN(new_n9242_));
  NAND2_X1   g08225(.A1(new_n9242_), .A2(new_n9240_), .ZN(new_n9243_));
  INV_X1     g08226(.I(new_n9243_), .ZN(new_n9244_));
  NAND2_X1   g08227(.A1(new_n8434_), .A2(new_n8490_), .ZN(new_n9245_));
  XOR2_X1    g08228(.A1(new_n8438_), .A2(new_n8443_), .Z(new_n9246_));
  XOR2_X1    g08229(.A1(new_n8458_), .A2(new_n8464_), .Z(new_n9247_));
  NOR4_X1    g08230(.A1(new_n9246_), .A2(new_n9247_), .A3(new_n8447_), .A4(new_n8465_), .ZN(new_n9248_));
  NAND2_X1   g08231(.A1(new_n8450_), .A2(new_n8444_), .ZN(new_n9249_));
  NAND2_X1   g08232(.A1(new_n8438_), .A2(new_n8443_), .ZN(new_n9250_));
  NAND2_X1   g08233(.A1(new_n8445_), .A2(new_n9250_), .ZN(new_n9251_));
  NAND2_X1   g08234(.A1(new_n9251_), .A2(new_n9249_), .ZN(new_n9252_));
  AOI21_X1   g08235(.A1(new_n9245_), .A2(new_n9248_), .B(new_n9252_), .ZN(new_n9253_));
  NAND3_X1   g08236(.A1(new_n9245_), .A2(new_n9248_), .A3(new_n9252_), .ZN(new_n9254_));
  INV_X1     g08237(.I(new_n9254_), .ZN(new_n9255_));
  OAI21_X1   g08238(.A1(new_n9255_), .A2(new_n9253_), .B(new_n9244_), .ZN(new_n9256_));
  NOR2_X1    g08239(.A1(new_n8454_), .A2(new_n8482_), .ZN(new_n9257_));
  NOR2_X1    g08240(.A1(new_n9257_), .A2(new_n8489_), .ZN(new_n9258_));
  INV_X1     g08241(.I(new_n9248_), .ZN(new_n9259_));
  INV_X1     g08242(.I(new_n9252_), .ZN(new_n9260_));
  OAI21_X1   g08243(.A1(new_n9258_), .A2(new_n9259_), .B(new_n9260_), .ZN(new_n9261_));
  NAND3_X1   g08244(.A1(new_n9261_), .A2(new_n9243_), .A3(new_n9254_), .ZN(new_n9262_));
  NAND2_X1   g08245(.A1(new_n9169_), .A2(new_n9176_), .ZN(new_n9263_));
  NAND2_X1   g08246(.A1(new_n9168_), .A2(new_n9173_), .ZN(new_n9264_));
  NAND3_X1   g08247(.A1(new_n9264_), .A2(new_n9181_), .A3(new_n9121_), .ZN(new_n9265_));
  NAND2_X1   g08248(.A1(new_n9265_), .A2(new_n9263_), .ZN(new_n9266_));
  INV_X1     g08249(.I(new_n9266_), .ZN(new_n9267_));
  NAND2_X1   g08250(.A1(new_n9143_), .A2(new_n9195_), .ZN(new_n9268_));
  XOR2_X1    g08251(.A1(new_n9147_), .A2(new_n9160_), .Z(new_n9269_));
  XOR2_X1    g08252(.A1(new_n9168_), .A2(new_n9173_), .Z(new_n9270_));
  NOR4_X1    g08253(.A1(new_n9269_), .A2(new_n9270_), .A3(new_n9161_), .A4(new_n9174_), .ZN(new_n9271_));
  NAND2_X1   g08254(.A1(new_n9159_), .A2(new_n9153_), .ZN(new_n9272_));
  NAND2_X1   g08255(.A1(new_n9147_), .A2(new_n9160_), .ZN(new_n9273_));
  NAND2_X1   g08256(.A1(new_n9154_), .A2(new_n9273_), .ZN(new_n9274_));
  NAND2_X1   g08257(.A1(new_n9274_), .A2(new_n9272_), .ZN(new_n9275_));
  AOI21_X1   g08258(.A1(new_n9268_), .A2(new_n9271_), .B(new_n9275_), .ZN(new_n9276_));
  NOR2_X1    g08259(.A1(new_n9164_), .A2(new_n9189_), .ZN(new_n9277_));
  NOR2_X1    g08260(.A1(new_n9277_), .A2(new_n9194_), .ZN(new_n9278_));
  INV_X1     g08261(.I(new_n9271_), .ZN(new_n9279_));
  INV_X1     g08262(.I(new_n9275_), .ZN(new_n9280_));
  NOR3_X1    g08263(.A1(new_n9278_), .A2(new_n9279_), .A3(new_n9280_), .ZN(new_n9281_));
  OAI21_X1   g08264(.A1(new_n9281_), .A2(new_n9276_), .B(new_n9267_), .ZN(new_n9282_));
  OAI21_X1   g08265(.A1(new_n9278_), .A2(new_n9279_), .B(new_n9280_), .ZN(new_n9283_));
  NAND3_X1   g08266(.A1(new_n9268_), .A2(new_n9271_), .A3(new_n9275_), .ZN(new_n9284_));
  NAND3_X1   g08267(.A1(new_n9283_), .A2(new_n9266_), .A3(new_n9284_), .ZN(new_n9285_));
  NAND4_X1   g08268(.A1(new_n9256_), .A2(new_n9262_), .A3(new_n9282_), .A4(new_n9285_), .ZN(new_n9286_));
  NAND2_X1   g08269(.A1(new_n9286_), .A2(new_n9239_), .ZN(new_n9287_));
  NAND2_X1   g08270(.A1(new_n9245_), .A2(new_n9248_), .ZN(new_n9288_));
  INV_X1     g08271(.I(new_n9288_), .ZN(new_n9289_));
  NOR2_X1    g08272(.A1(new_n9278_), .A2(new_n9279_), .ZN(new_n9290_));
  XNOR2_X1   g08273(.A1(new_n9275_), .A2(new_n9266_), .ZN(new_n9291_));
  XNOR2_X1   g08274(.A1(new_n9252_), .A2(new_n9243_), .ZN(new_n9292_));
  AND4_X2    g08275(.A1(new_n9289_), .A2(new_n9290_), .A3(new_n9291_), .A4(new_n9292_), .Z(new_n9293_));
  NAND2_X1   g08276(.A1(new_n9287_), .A2(new_n9293_), .ZN(new_n9294_));
  AOI22_X1   g08277(.A1(new_n9272_), .A2(new_n9161_), .B1(new_n9263_), .B2(new_n9174_), .ZN(new_n9295_));
  AOI21_X1   g08278(.A1(new_n9264_), .A2(new_n9273_), .B(new_n9295_), .ZN(new_n9296_));
  OR2_X2     g08279(.A1(new_n9290_), .A2(new_n9296_), .Z(new_n9297_));
  AOI22_X1   g08280(.A1(new_n9249_), .A2(new_n8447_), .B1(new_n9240_), .B2(new_n8465_), .ZN(new_n9298_));
  AOI21_X1   g08281(.A1(new_n9241_), .A2(new_n9250_), .B(new_n9298_), .ZN(new_n9299_));
  NOR2_X1    g08282(.A1(new_n9289_), .A2(new_n9299_), .ZN(new_n9300_));
  INV_X1     g08283(.I(new_n9300_), .ZN(new_n9301_));
  NOR2_X1    g08284(.A1(new_n9252_), .A2(new_n9243_), .ZN(new_n9302_));
  NOR2_X1    g08285(.A1(new_n9275_), .A2(new_n9266_), .ZN(new_n9303_));
  NOR4_X1    g08286(.A1(new_n9301_), .A2(new_n9297_), .A3(new_n9302_), .A4(new_n9303_), .ZN(new_n9304_));
  NOR2_X1    g08287(.A1(new_n9297_), .A2(new_n9303_), .ZN(new_n9305_));
  INV_X1     g08288(.I(new_n9305_), .ZN(new_n9306_));
  NOR2_X1    g08289(.A1(new_n9301_), .A2(new_n9302_), .ZN(new_n9307_));
  INV_X1     g08290(.I(new_n9307_), .ZN(new_n9308_));
  AOI22_X1   g08291(.A1(new_n9294_), .A2(new_n9304_), .B1(new_n9306_), .B2(new_n9308_), .ZN(new_n9309_));
  NOR2_X1    g08292(.A1(\A[41] ), .A2(\A[42] ), .ZN(new_n9310_));
  AOI21_X1   g08293(.A1(\A[41] ), .A2(\A[42] ), .B(\A[40] ), .ZN(new_n9311_));
  NOR2_X1    g08294(.A1(new_n9311_), .A2(new_n9310_), .ZN(new_n9312_));
  NOR2_X1    g08295(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n9313_));
  AOI21_X1   g08296(.A1(\A[38] ), .A2(\A[39] ), .B(\A[37] ), .ZN(new_n9314_));
  NOR2_X1    g08297(.A1(new_n9314_), .A2(new_n9313_), .ZN(new_n9315_));
  NAND2_X1   g08298(.A1(new_n9312_), .A2(new_n9315_), .ZN(new_n9316_));
  INV_X1     g08299(.I(\A[39] ), .ZN(new_n9317_));
  NOR2_X1    g08300(.A1(new_n9317_), .A2(\A[38] ), .ZN(new_n9318_));
  INV_X1     g08301(.I(\A[38] ), .ZN(new_n9319_));
  NOR2_X1    g08302(.A1(new_n9319_), .A2(\A[39] ), .ZN(new_n9320_));
  OAI21_X1   g08303(.A1(new_n9318_), .A2(new_n9320_), .B(\A[37] ), .ZN(new_n9321_));
  INV_X1     g08304(.I(\A[37] ), .ZN(new_n9322_));
  NAND2_X1   g08305(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n9323_));
  INV_X1     g08306(.I(new_n9323_), .ZN(new_n9324_));
  OAI21_X1   g08307(.A1(new_n9324_), .A2(new_n9313_), .B(new_n9322_), .ZN(new_n9325_));
  INV_X1     g08308(.I(\A[42] ), .ZN(new_n9326_));
  NOR2_X1    g08309(.A1(new_n9326_), .A2(\A[41] ), .ZN(new_n9327_));
  INV_X1     g08310(.I(\A[41] ), .ZN(new_n9328_));
  NOR2_X1    g08311(.A1(new_n9328_), .A2(\A[42] ), .ZN(new_n9329_));
  OAI21_X1   g08312(.A1(new_n9327_), .A2(new_n9329_), .B(\A[40] ), .ZN(new_n9330_));
  INV_X1     g08313(.I(\A[40] ), .ZN(new_n9331_));
  NAND2_X1   g08314(.A1(\A[41] ), .A2(\A[42] ), .ZN(new_n9332_));
  INV_X1     g08315(.I(new_n9332_), .ZN(new_n9333_));
  OAI21_X1   g08316(.A1(new_n9333_), .A2(new_n9310_), .B(new_n9331_), .ZN(new_n9334_));
  NAND4_X1   g08317(.A1(new_n9321_), .A2(new_n9325_), .A3(new_n9330_), .A4(new_n9334_), .ZN(new_n9335_));
  OAI22_X1   g08318(.A1(new_n9310_), .A2(new_n9311_), .B1(new_n9314_), .B2(new_n9313_), .ZN(new_n9336_));
  INV_X1     g08319(.I(new_n9336_), .ZN(new_n9337_));
  OAI21_X1   g08320(.A1(new_n9335_), .A2(new_n9337_), .B(new_n9316_), .ZN(new_n9338_));
  INV_X1     g08321(.I(new_n9315_), .ZN(new_n9339_));
  NAND2_X1   g08322(.A1(new_n9319_), .A2(\A[39] ), .ZN(new_n9340_));
  NAND2_X1   g08323(.A1(new_n9317_), .A2(\A[38] ), .ZN(new_n9341_));
  AOI21_X1   g08324(.A1(new_n9340_), .A2(new_n9341_), .B(new_n9322_), .ZN(new_n9342_));
  INV_X1     g08325(.I(new_n9313_), .ZN(new_n9343_));
  AOI21_X1   g08326(.A1(new_n9343_), .A2(new_n9323_), .B(\A[37] ), .ZN(new_n9344_));
  NAND2_X1   g08327(.A1(new_n9328_), .A2(\A[42] ), .ZN(new_n9345_));
  NAND2_X1   g08328(.A1(new_n9326_), .A2(\A[41] ), .ZN(new_n9346_));
  AOI21_X1   g08329(.A1(new_n9345_), .A2(new_n9346_), .B(new_n9331_), .ZN(new_n9347_));
  INV_X1     g08330(.I(new_n9310_), .ZN(new_n9348_));
  AOI21_X1   g08331(.A1(new_n9348_), .A2(new_n9332_), .B(\A[40] ), .ZN(new_n9349_));
  NOR4_X1    g08332(.A1(new_n9342_), .A2(new_n9344_), .A3(new_n9349_), .A4(new_n9347_), .ZN(new_n9350_));
  NOR2_X1    g08333(.A1(new_n9350_), .A2(new_n9339_), .ZN(new_n9351_));
  NAND2_X1   g08334(.A1(new_n9321_), .A2(new_n9325_), .ZN(new_n9352_));
  NAND2_X1   g08335(.A1(new_n9330_), .A2(new_n9334_), .ZN(new_n9353_));
  NOR3_X1    g08336(.A1(new_n9352_), .A2(new_n9353_), .A3(new_n9315_), .ZN(new_n9354_));
  OAI21_X1   g08337(.A1(new_n9351_), .A2(new_n9354_), .B(new_n9312_), .ZN(new_n9355_));
  INV_X1     g08338(.I(new_n9312_), .ZN(new_n9356_));
  NAND2_X1   g08339(.A1(new_n9335_), .A2(new_n9315_), .ZN(new_n9357_));
  NAND2_X1   g08340(.A1(new_n9350_), .A2(new_n9339_), .ZN(new_n9358_));
  NAND3_X1   g08341(.A1(new_n9358_), .A2(new_n9357_), .A3(new_n9356_), .ZN(new_n9359_));
  NAND2_X1   g08342(.A1(new_n9359_), .A2(new_n9355_), .ZN(new_n9360_));
  NOR2_X1    g08343(.A1(new_n9344_), .A2(new_n9342_), .ZN(new_n9361_));
  NOR2_X1    g08344(.A1(new_n9349_), .A2(new_n9347_), .ZN(new_n9362_));
  NOR2_X1    g08345(.A1(new_n9361_), .A2(new_n9362_), .ZN(new_n9363_));
  NOR2_X1    g08346(.A1(new_n9363_), .A2(new_n9350_), .ZN(new_n9364_));
  INV_X1     g08347(.I(new_n9364_), .ZN(new_n9365_));
  OAI21_X1   g08348(.A1(new_n9360_), .A2(new_n9365_), .B(new_n9338_), .ZN(new_n9366_));
  INV_X1     g08349(.I(new_n9366_), .ZN(new_n9367_));
  INV_X1     g08350(.I(\A[34] ), .ZN(new_n9368_));
  NOR2_X1    g08351(.A1(\A[35] ), .A2(\A[36] ), .ZN(new_n9369_));
  NAND2_X1   g08352(.A1(\A[35] ), .A2(\A[36] ), .ZN(new_n9370_));
  AOI21_X1   g08353(.A1(new_n9368_), .A2(new_n9370_), .B(new_n9369_), .ZN(new_n9371_));
  INV_X1     g08354(.I(\A[31] ), .ZN(new_n9372_));
  NOR2_X1    g08355(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n9373_));
  NAND2_X1   g08356(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n9374_));
  AOI21_X1   g08357(.A1(new_n9372_), .A2(new_n9374_), .B(new_n9373_), .ZN(new_n9375_));
  NAND2_X1   g08358(.A1(new_n9371_), .A2(new_n9375_), .ZN(new_n9376_));
  NOR2_X1    g08359(.A1(new_n9371_), .A2(new_n9375_), .ZN(new_n9377_));
  INV_X1     g08360(.I(\A[33] ), .ZN(new_n9378_));
  NOR2_X1    g08361(.A1(new_n9378_), .A2(\A[32] ), .ZN(new_n9379_));
  INV_X1     g08362(.I(\A[32] ), .ZN(new_n9380_));
  NOR2_X1    g08363(.A1(new_n9380_), .A2(\A[33] ), .ZN(new_n9381_));
  OAI21_X1   g08364(.A1(new_n9379_), .A2(new_n9381_), .B(\A[31] ), .ZN(new_n9382_));
  INV_X1     g08365(.I(new_n9374_), .ZN(new_n9383_));
  OAI21_X1   g08366(.A1(new_n9383_), .A2(new_n9373_), .B(new_n9372_), .ZN(new_n9384_));
  INV_X1     g08367(.I(\A[36] ), .ZN(new_n9385_));
  NOR2_X1    g08368(.A1(new_n9385_), .A2(\A[35] ), .ZN(new_n9386_));
  INV_X1     g08369(.I(\A[35] ), .ZN(new_n9387_));
  NOR2_X1    g08370(.A1(new_n9387_), .A2(\A[36] ), .ZN(new_n9388_));
  OAI21_X1   g08371(.A1(new_n9386_), .A2(new_n9388_), .B(\A[34] ), .ZN(new_n9389_));
  INV_X1     g08372(.I(new_n9370_), .ZN(new_n9390_));
  OAI21_X1   g08373(.A1(new_n9390_), .A2(new_n9369_), .B(new_n9368_), .ZN(new_n9391_));
  NAND4_X1   g08374(.A1(new_n9382_), .A2(new_n9384_), .A3(new_n9389_), .A4(new_n9391_), .ZN(new_n9392_));
  OAI21_X1   g08375(.A1(new_n9392_), .A2(new_n9377_), .B(new_n9376_), .ZN(new_n9393_));
  NAND2_X1   g08376(.A1(new_n9352_), .A2(new_n9353_), .ZN(new_n9394_));
  NAND4_X1   g08377(.A1(new_n9394_), .A2(new_n9312_), .A3(new_n9315_), .A4(new_n9335_), .ZN(new_n9395_));
  NAND2_X1   g08378(.A1(new_n9361_), .A2(new_n9353_), .ZN(new_n9396_));
  NAND2_X1   g08379(.A1(new_n9362_), .A2(new_n9352_), .ZN(new_n9397_));
  NAND2_X1   g08380(.A1(new_n9380_), .A2(\A[33] ), .ZN(new_n9398_));
  NAND2_X1   g08381(.A1(new_n9378_), .A2(\A[32] ), .ZN(new_n9399_));
  AOI21_X1   g08382(.A1(new_n9398_), .A2(new_n9399_), .B(new_n9372_), .ZN(new_n9400_));
  INV_X1     g08383(.I(new_n9373_), .ZN(new_n9401_));
  AOI21_X1   g08384(.A1(new_n9401_), .A2(new_n9374_), .B(\A[31] ), .ZN(new_n9402_));
  NOR2_X1    g08385(.A1(new_n9402_), .A2(new_n9400_), .ZN(new_n9403_));
  NAND2_X1   g08386(.A1(new_n9389_), .A2(new_n9391_), .ZN(new_n9404_));
  NAND2_X1   g08387(.A1(new_n9403_), .A2(new_n9404_), .ZN(new_n9405_));
  NAND2_X1   g08388(.A1(new_n9382_), .A2(new_n9384_), .ZN(new_n9406_));
  NAND2_X1   g08389(.A1(new_n9387_), .A2(\A[36] ), .ZN(new_n9407_));
  NAND2_X1   g08390(.A1(new_n9385_), .A2(\A[35] ), .ZN(new_n9408_));
  AOI21_X1   g08391(.A1(new_n9407_), .A2(new_n9408_), .B(new_n9368_), .ZN(new_n9409_));
  INV_X1     g08392(.I(new_n9369_), .ZN(new_n9410_));
  AOI21_X1   g08393(.A1(new_n9410_), .A2(new_n9370_), .B(\A[34] ), .ZN(new_n9411_));
  NOR2_X1    g08394(.A1(new_n9411_), .A2(new_n9409_), .ZN(new_n9412_));
  NAND2_X1   g08395(.A1(new_n9412_), .A2(new_n9406_), .ZN(new_n9413_));
  AOI22_X1   g08396(.A1(new_n9396_), .A2(new_n9397_), .B1(new_n9405_), .B2(new_n9413_), .ZN(new_n9414_));
  NOR3_X1    g08397(.A1(new_n9338_), .A2(new_n9376_), .A3(new_n9392_), .ZN(new_n9415_));
  NAND3_X1   g08398(.A1(new_n9415_), .A2(new_n9414_), .A3(new_n9395_), .ZN(new_n9416_));
  NOR2_X1    g08399(.A1(new_n9416_), .A2(new_n9360_), .ZN(new_n9417_));
  NOR4_X1    g08400(.A1(new_n9335_), .A2(new_n9392_), .A3(new_n9316_), .A4(new_n9376_), .ZN(new_n9418_));
  NOR2_X1    g08401(.A1(new_n9414_), .A2(new_n9418_), .ZN(new_n9419_));
  INV_X1     g08402(.I(new_n9371_), .ZN(new_n9420_));
  NAND2_X1   g08403(.A1(new_n9392_), .A2(new_n9375_), .ZN(new_n9421_));
  INV_X1     g08404(.I(new_n9375_), .ZN(new_n9422_));
  NOR4_X1    g08405(.A1(new_n9400_), .A2(new_n9402_), .A3(new_n9411_), .A4(new_n9409_), .ZN(new_n9423_));
  NAND2_X1   g08406(.A1(new_n9423_), .A2(new_n9422_), .ZN(new_n9424_));
  AOI21_X1   g08407(.A1(new_n9424_), .A2(new_n9421_), .B(new_n9420_), .ZN(new_n9425_));
  NOR2_X1    g08408(.A1(new_n9423_), .A2(new_n9422_), .ZN(new_n9426_));
  NOR2_X1    g08409(.A1(new_n9392_), .A2(new_n9375_), .ZN(new_n9427_));
  NOR3_X1    g08410(.A1(new_n9426_), .A2(new_n9427_), .A3(new_n9371_), .ZN(new_n9428_));
  NOR2_X1    g08411(.A1(new_n9425_), .A2(new_n9428_), .ZN(new_n9429_));
  NOR3_X1    g08412(.A1(new_n9429_), .A2(new_n9360_), .A3(new_n9419_), .ZN(new_n9430_));
  OAI21_X1   g08413(.A1(new_n9430_), .A2(new_n9417_), .B(new_n9393_), .ZN(new_n9431_));
  INV_X1     g08414(.I(new_n9393_), .ZN(new_n9432_));
  AOI21_X1   g08415(.A1(new_n9358_), .A2(new_n9357_), .B(new_n9356_), .ZN(new_n9433_));
  NOR3_X1    g08416(.A1(new_n9351_), .A2(new_n9354_), .A3(new_n9312_), .ZN(new_n9434_));
  NOR2_X1    g08417(.A1(new_n9433_), .A2(new_n9434_), .ZN(new_n9435_));
  NOR4_X1    g08418(.A1(new_n9363_), .A2(new_n9350_), .A3(new_n9356_), .A4(new_n9339_), .ZN(new_n9436_));
  NOR2_X1    g08419(.A1(new_n9362_), .A2(new_n9352_), .ZN(new_n9437_));
  NOR2_X1    g08420(.A1(new_n9361_), .A2(new_n9353_), .ZN(new_n9438_));
  NOR2_X1    g08421(.A1(new_n9412_), .A2(new_n9406_), .ZN(new_n9439_));
  NOR2_X1    g08422(.A1(new_n9403_), .A2(new_n9404_), .ZN(new_n9440_));
  OAI22_X1   g08423(.A1(new_n9437_), .A2(new_n9438_), .B1(new_n9439_), .B2(new_n9440_), .ZN(new_n9441_));
  NAND3_X1   g08424(.A1(new_n9361_), .A2(new_n9362_), .A3(new_n9336_), .ZN(new_n9442_));
  INV_X1     g08425(.I(new_n9376_), .ZN(new_n9443_));
  NAND4_X1   g08426(.A1(new_n9442_), .A2(new_n9316_), .A3(new_n9443_), .A4(new_n9423_), .ZN(new_n9444_));
  NOR3_X1    g08427(.A1(new_n9441_), .A2(new_n9436_), .A3(new_n9444_), .ZN(new_n9445_));
  NAND2_X1   g08428(.A1(new_n9445_), .A2(new_n9435_), .ZN(new_n9446_));
  INV_X1     g08429(.I(new_n9316_), .ZN(new_n9447_));
  NAND4_X1   g08430(.A1(new_n9350_), .A2(new_n9423_), .A3(new_n9447_), .A4(new_n9443_), .ZN(new_n9448_));
  NAND2_X1   g08431(.A1(new_n9441_), .A2(new_n9448_), .ZN(new_n9449_));
  OAI21_X1   g08432(.A1(new_n9426_), .A2(new_n9427_), .B(new_n9371_), .ZN(new_n9450_));
  NAND3_X1   g08433(.A1(new_n9424_), .A2(new_n9421_), .A3(new_n9420_), .ZN(new_n9451_));
  NAND2_X1   g08434(.A1(new_n9450_), .A2(new_n9451_), .ZN(new_n9452_));
  NAND3_X1   g08435(.A1(new_n9452_), .A2(new_n9435_), .A3(new_n9449_), .ZN(new_n9453_));
  NAND3_X1   g08436(.A1(new_n9453_), .A2(new_n9446_), .A3(new_n9432_), .ZN(new_n9454_));
  AOI21_X1   g08437(.A1(new_n9431_), .A2(new_n9454_), .B(new_n9367_), .ZN(new_n9455_));
  AOI21_X1   g08438(.A1(new_n9453_), .A2(new_n9446_), .B(new_n9432_), .ZN(new_n9456_));
  NOR3_X1    g08439(.A1(new_n9430_), .A2(new_n9417_), .A3(new_n9393_), .ZN(new_n9457_));
  NOR3_X1    g08440(.A1(new_n9457_), .A2(new_n9456_), .A3(new_n9366_), .ZN(new_n9458_));
  NOR2_X1    g08441(.A1(new_n9458_), .A2(new_n9455_), .ZN(new_n9459_));
  INV_X1     g08442(.I(\A[43] ), .ZN(new_n9460_));
  INV_X1     g08443(.I(\A[44] ), .ZN(new_n9461_));
  NAND2_X1   g08444(.A1(new_n9461_), .A2(\A[45] ), .ZN(new_n9462_));
  INV_X1     g08445(.I(\A[45] ), .ZN(new_n9463_));
  NAND2_X1   g08446(.A1(new_n9463_), .A2(\A[44] ), .ZN(new_n9464_));
  AOI21_X1   g08447(.A1(new_n9462_), .A2(new_n9464_), .B(new_n9460_), .ZN(new_n9465_));
  NOR2_X1    g08448(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n9466_));
  INV_X1     g08449(.I(new_n9466_), .ZN(new_n9467_));
  NAND2_X1   g08450(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n9468_));
  AOI21_X1   g08451(.A1(new_n9467_), .A2(new_n9468_), .B(\A[43] ), .ZN(new_n9469_));
  NOR2_X1    g08452(.A1(new_n9469_), .A2(new_n9465_), .ZN(new_n9470_));
  INV_X1     g08453(.I(\A[48] ), .ZN(new_n9471_));
  NOR2_X1    g08454(.A1(new_n9471_), .A2(\A[47] ), .ZN(new_n9472_));
  INV_X1     g08455(.I(\A[47] ), .ZN(new_n9473_));
  NOR2_X1    g08456(.A1(new_n9473_), .A2(\A[48] ), .ZN(new_n9474_));
  OAI21_X1   g08457(.A1(new_n9472_), .A2(new_n9474_), .B(\A[46] ), .ZN(new_n9475_));
  INV_X1     g08458(.I(\A[46] ), .ZN(new_n9476_));
  NOR2_X1    g08459(.A1(\A[47] ), .A2(\A[48] ), .ZN(new_n9477_));
  NAND2_X1   g08460(.A1(\A[47] ), .A2(\A[48] ), .ZN(new_n9478_));
  INV_X1     g08461(.I(new_n9478_), .ZN(new_n9479_));
  OAI21_X1   g08462(.A1(new_n9479_), .A2(new_n9477_), .B(new_n9476_), .ZN(new_n9480_));
  NAND2_X1   g08463(.A1(new_n9475_), .A2(new_n9480_), .ZN(new_n9481_));
  NAND2_X1   g08464(.A1(new_n9470_), .A2(new_n9481_), .ZN(new_n9482_));
  NOR2_X1    g08465(.A1(new_n9463_), .A2(\A[44] ), .ZN(new_n9483_));
  NOR2_X1    g08466(.A1(new_n9461_), .A2(\A[45] ), .ZN(new_n9484_));
  OAI21_X1   g08467(.A1(new_n9483_), .A2(new_n9484_), .B(\A[43] ), .ZN(new_n9485_));
  INV_X1     g08468(.I(new_n9468_), .ZN(new_n9486_));
  OAI21_X1   g08469(.A1(new_n9486_), .A2(new_n9466_), .B(new_n9460_), .ZN(new_n9487_));
  NAND2_X1   g08470(.A1(new_n9485_), .A2(new_n9487_), .ZN(new_n9488_));
  NAND2_X1   g08471(.A1(new_n9473_), .A2(\A[48] ), .ZN(new_n9489_));
  NAND2_X1   g08472(.A1(new_n9471_), .A2(\A[47] ), .ZN(new_n9490_));
  AOI21_X1   g08473(.A1(new_n9489_), .A2(new_n9490_), .B(new_n9476_), .ZN(new_n9491_));
  INV_X1     g08474(.I(new_n9477_), .ZN(new_n9492_));
  AOI21_X1   g08475(.A1(new_n9492_), .A2(new_n9478_), .B(\A[46] ), .ZN(new_n9493_));
  NOR2_X1    g08476(.A1(new_n9493_), .A2(new_n9491_), .ZN(new_n9494_));
  NAND2_X1   g08477(.A1(new_n9494_), .A2(new_n9488_), .ZN(new_n9495_));
  NAND2_X1   g08478(.A1(new_n9482_), .A2(new_n9495_), .ZN(new_n9496_));
  INV_X1     g08479(.I(\A[51] ), .ZN(new_n9497_));
  NOR2_X1    g08480(.A1(new_n9497_), .A2(\A[50] ), .ZN(new_n9498_));
  INV_X1     g08481(.I(\A[50] ), .ZN(new_n9499_));
  NOR2_X1    g08482(.A1(new_n9499_), .A2(\A[51] ), .ZN(new_n9500_));
  OAI21_X1   g08483(.A1(new_n9498_), .A2(new_n9500_), .B(\A[49] ), .ZN(new_n9501_));
  INV_X1     g08484(.I(\A[49] ), .ZN(new_n9502_));
  NOR2_X1    g08485(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n9503_));
  AND2_X2    g08486(.A1(\A[50] ), .A2(\A[51] ), .Z(new_n9504_));
  OAI21_X1   g08487(.A1(new_n9504_), .A2(new_n9503_), .B(new_n9502_), .ZN(new_n9505_));
  NAND2_X1   g08488(.A1(new_n9501_), .A2(new_n9505_), .ZN(new_n9506_));
  INV_X1     g08489(.I(\A[52] ), .ZN(new_n9507_));
  INV_X1     g08490(.I(\A[53] ), .ZN(new_n9508_));
  NAND2_X1   g08491(.A1(new_n9508_), .A2(\A[54] ), .ZN(new_n9509_));
  INV_X1     g08492(.I(\A[54] ), .ZN(new_n9510_));
  NAND2_X1   g08493(.A1(new_n9510_), .A2(\A[53] ), .ZN(new_n9511_));
  AOI21_X1   g08494(.A1(new_n9509_), .A2(new_n9511_), .B(new_n9507_), .ZN(new_n9512_));
  OR2_X2     g08495(.A1(\A[53] ), .A2(\A[54] ), .Z(new_n9513_));
  NAND2_X1   g08496(.A1(\A[53] ), .A2(\A[54] ), .ZN(new_n9514_));
  AOI21_X1   g08497(.A1(new_n9513_), .A2(new_n9514_), .B(\A[52] ), .ZN(new_n9515_));
  NOR2_X1    g08498(.A1(new_n9512_), .A2(new_n9515_), .ZN(new_n9516_));
  NOR2_X1    g08499(.A1(new_n9516_), .A2(new_n9506_), .ZN(new_n9517_));
  NAND2_X1   g08500(.A1(new_n9499_), .A2(\A[51] ), .ZN(new_n9518_));
  NAND2_X1   g08501(.A1(new_n9497_), .A2(\A[50] ), .ZN(new_n9519_));
  AOI21_X1   g08502(.A1(new_n9518_), .A2(new_n9519_), .B(new_n9502_), .ZN(new_n9520_));
  INV_X1     g08503(.I(new_n9503_), .ZN(new_n9521_));
  NAND2_X1   g08504(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n9522_));
  AOI21_X1   g08505(.A1(new_n9521_), .A2(new_n9522_), .B(\A[49] ), .ZN(new_n9523_));
  NOR2_X1    g08506(.A1(new_n9523_), .A2(new_n9520_), .ZN(new_n9524_));
  NOR2_X1    g08507(.A1(new_n9510_), .A2(\A[53] ), .ZN(new_n9525_));
  NOR2_X1    g08508(.A1(new_n9508_), .A2(\A[54] ), .ZN(new_n9526_));
  OAI21_X1   g08509(.A1(new_n9525_), .A2(new_n9526_), .B(\A[52] ), .ZN(new_n9527_));
  NOR2_X1    g08510(.A1(\A[53] ), .A2(\A[54] ), .ZN(new_n9528_));
  AND2_X2    g08511(.A1(\A[53] ), .A2(\A[54] ), .Z(new_n9529_));
  OAI21_X1   g08512(.A1(new_n9529_), .A2(new_n9528_), .B(new_n9507_), .ZN(new_n9530_));
  NAND2_X1   g08513(.A1(new_n9527_), .A2(new_n9530_), .ZN(new_n9531_));
  NOR2_X1    g08514(.A1(new_n9524_), .A2(new_n9531_), .ZN(new_n9532_));
  NOR2_X1    g08515(.A1(new_n9517_), .A2(new_n9532_), .ZN(new_n9533_));
  NAND2_X1   g08516(.A1(new_n9496_), .A2(new_n9533_), .ZN(new_n9534_));
  NOR2_X1    g08517(.A1(new_n9494_), .A2(new_n9488_), .ZN(new_n9535_));
  NOR2_X1    g08518(.A1(new_n9470_), .A2(new_n9481_), .ZN(new_n9536_));
  NOR2_X1    g08519(.A1(new_n9535_), .A2(new_n9536_), .ZN(new_n9537_));
  NAND2_X1   g08520(.A1(new_n9524_), .A2(new_n9531_), .ZN(new_n9538_));
  NAND3_X1   g08521(.A1(new_n9506_), .A2(new_n9527_), .A3(new_n9530_), .ZN(new_n9539_));
  NAND2_X1   g08522(.A1(new_n9538_), .A2(new_n9539_), .ZN(new_n9540_));
  NAND2_X1   g08523(.A1(new_n9537_), .A2(new_n9540_), .ZN(new_n9541_));
  NAND2_X1   g08524(.A1(new_n9534_), .A2(new_n9541_), .ZN(new_n9542_));
  NOR2_X1    g08525(.A1(new_n9437_), .A2(new_n9438_), .ZN(new_n9543_));
  NAND2_X1   g08526(.A1(new_n9405_), .A2(new_n9413_), .ZN(new_n9544_));
  NAND2_X1   g08527(.A1(new_n9543_), .A2(new_n9544_), .ZN(new_n9545_));
  NAND2_X1   g08528(.A1(new_n9396_), .A2(new_n9397_), .ZN(new_n9546_));
  NOR2_X1    g08529(.A1(new_n9439_), .A2(new_n9440_), .ZN(new_n9547_));
  NAND2_X1   g08530(.A1(new_n9547_), .A2(new_n9546_), .ZN(new_n9548_));
  NAND2_X1   g08531(.A1(new_n9545_), .A2(new_n9548_), .ZN(new_n9549_));
  NAND2_X1   g08532(.A1(new_n9549_), .A2(new_n9542_), .ZN(new_n9550_));
  AOI21_X1   g08533(.A1(new_n9476_), .A2(new_n9478_), .B(new_n9477_), .ZN(new_n9551_));
  AOI21_X1   g08534(.A1(new_n9460_), .A2(new_n9468_), .B(new_n9466_), .ZN(new_n9552_));
  INV_X1     g08535(.I(new_n9552_), .ZN(new_n9553_));
  NOR4_X1    g08536(.A1(new_n9465_), .A2(new_n9469_), .A3(new_n9493_), .A4(new_n9491_), .ZN(new_n9554_));
  NOR2_X1    g08537(.A1(new_n9554_), .A2(new_n9553_), .ZN(new_n9555_));
  NAND4_X1   g08538(.A1(new_n9485_), .A2(new_n9487_), .A3(new_n9475_), .A4(new_n9480_), .ZN(new_n9556_));
  NOR2_X1    g08539(.A1(new_n9556_), .A2(new_n9552_), .ZN(new_n9557_));
  OAI21_X1   g08540(.A1(new_n9555_), .A2(new_n9557_), .B(new_n9551_), .ZN(new_n9558_));
  INV_X1     g08541(.I(new_n9551_), .ZN(new_n9559_));
  NAND2_X1   g08542(.A1(new_n9556_), .A2(new_n9552_), .ZN(new_n9560_));
  NAND3_X1   g08543(.A1(new_n9470_), .A2(new_n9494_), .A3(new_n9553_), .ZN(new_n9561_));
  NAND3_X1   g08544(.A1(new_n9560_), .A2(new_n9561_), .A3(new_n9559_), .ZN(new_n9562_));
  NAND2_X1   g08545(.A1(new_n9558_), .A2(new_n9562_), .ZN(new_n9563_));
  AOI21_X1   g08546(.A1(new_n9507_), .A2(new_n9514_), .B(new_n9528_), .ZN(new_n9564_));
  INV_X1     g08547(.I(new_n9564_), .ZN(new_n9565_));
  AOI21_X1   g08548(.A1(new_n9502_), .A2(new_n9522_), .B(new_n9503_), .ZN(new_n9566_));
  NAND4_X1   g08549(.A1(new_n9501_), .A2(new_n9527_), .A3(new_n9505_), .A4(new_n9530_), .ZN(new_n9567_));
  NAND2_X1   g08550(.A1(new_n9567_), .A2(new_n9566_), .ZN(new_n9568_));
  INV_X1     g08551(.I(new_n9566_), .ZN(new_n9569_));
  NAND3_X1   g08552(.A1(new_n9524_), .A2(new_n9516_), .A3(new_n9569_), .ZN(new_n9570_));
  AOI21_X1   g08553(.A1(new_n9568_), .A2(new_n9570_), .B(new_n9565_), .ZN(new_n9571_));
  AOI21_X1   g08554(.A1(new_n9524_), .A2(new_n9516_), .B(new_n9569_), .ZN(new_n9572_));
  NOR3_X1    g08555(.A1(new_n9506_), .A2(new_n9531_), .A3(new_n9566_), .ZN(new_n9573_));
  NOR3_X1    g08556(.A1(new_n9572_), .A2(new_n9573_), .A3(new_n9564_), .ZN(new_n9574_));
  NOR2_X1    g08557(.A1(new_n9571_), .A2(new_n9574_), .ZN(new_n9575_));
  NOR4_X1    g08558(.A1(new_n9520_), .A2(new_n9523_), .A3(new_n9512_), .A4(new_n9515_), .ZN(new_n9576_));
  NAND2_X1   g08559(.A1(new_n9551_), .A2(new_n9552_), .ZN(new_n9577_));
  INV_X1     g08560(.I(new_n9577_), .ZN(new_n9578_));
  NAND2_X1   g08561(.A1(new_n9564_), .A2(new_n9566_), .ZN(new_n9579_));
  INV_X1     g08562(.I(new_n9579_), .ZN(new_n9580_));
  NAND4_X1   g08563(.A1(new_n9554_), .A2(new_n9576_), .A3(new_n9578_), .A4(new_n9580_), .ZN(new_n9581_));
  OAI21_X1   g08564(.A1(new_n9537_), .A2(new_n9533_), .B(new_n9581_), .ZN(new_n9582_));
  NAND2_X1   g08565(.A1(new_n9575_), .A2(new_n9582_), .ZN(new_n9583_));
  OAI22_X1   g08566(.A1(new_n9535_), .A2(new_n9536_), .B1(new_n9517_), .B2(new_n9532_), .ZN(new_n9584_));
  OAI21_X1   g08567(.A1(new_n9524_), .A2(new_n9516_), .B(new_n9580_), .ZN(new_n9585_));
  NAND3_X1   g08568(.A1(new_n9585_), .A2(new_n9554_), .A3(new_n9578_), .ZN(new_n9586_));
  NOR4_X1    g08569(.A1(new_n9586_), .A2(new_n9584_), .A3(new_n9571_), .A4(new_n9574_), .ZN(new_n9587_));
  OAI21_X1   g08570(.A1(new_n9583_), .A2(new_n9587_), .B(new_n9563_), .ZN(new_n9588_));
  AOI21_X1   g08571(.A1(new_n9560_), .A2(new_n9561_), .B(new_n9559_), .ZN(new_n9589_));
  NOR3_X1    g08572(.A1(new_n9555_), .A2(new_n9557_), .A3(new_n9551_), .ZN(new_n9590_));
  NOR2_X1    g08573(.A1(new_n9590_), .A2(new_n9589_), .ZN(new_n9591_));
  OAI21_X1   g08574(.A1(new_n9572_), .A2(new_n9573_), .B(new_n9564_), .ZN(new_n9592_));
  NAND3_X1   g08575(.A1(new_n9568_), .A2(new_n9570_), .A3(new_n9565_), .ZN(new_n9593_));
  AOI22_X1   g08576(.A1(new_n9482_), .A2(new_n9495_), .B1(new_n9538_), .B2(new_n9539_), .ZN(new_n9594_));
  NOR4_X1    g08577(.A1(new_n9556_), .A2(new_n9567_), .A3(new_n9577_), .A4(new_n9579_), .ZN(new_n9595_));
  AOI22_X1   g08578(.A1(new_n9594_), .A2(new_n9595_), .B1(new_n9592_), .B2(new_n9593_), .ZN(new_n9596_));
  NOR4_X1    g08579(.A1(new_n9584_), .A2(new_n9571_), .A3(new_n9574_), .A4(new_n9581_), .ZN(new_n9597_));
  OAI21_X1   g08580(.A1(new_n9596_), .A2(new_n9597_), .B(new_n9591_), .ZN(new_n9598_));
  AOI21_X1   g08581(.A1(new_n9588_), .A2(new_n9598_), .B(new_n9550_), .ZN(new_n9599_));
  NAND3_X1   g08582(.A1(new_n9416_), .A2(new_n9435_), .A3(new_n9449_), .ZN(new_n9600_));
  OAI22_X1   g08583(.A1(new_n9441_), .A2(new_n9448_), .B1(new_n9433_), .B2(new_n9434_), .ZN(new_n9601_));
  NAND4_X1   g08584(.A1(new_n9414_), .A2(new_n9359_), .A3(new_n9355_), .A4(new_n9418_), .ZN(new_n9602_));
  AOI21_X1   g08585(.A1(new_n9601_), .A2(new_n9602_), .B(new_n9452_), .ZN(new_n9603_));
  AOI21_X1   g08586(.A1(new_n9452_), .A2(new_n9600_), .B(new_n9603_), .ZN(new_n9604_));
  OAI22_X1   g08587(.A1(new_n9584_), .A2(new_n9581_), .B1(new_n9571_), .B2(new_n9574_), .ZN(new_n9605_));
  NAND4_X1   g08588(.A1(new_n9594_), .A2(new_n9592_), .A3(new_n9593_), .A4(new_n9595_), .ZN(new_n9606_));
  AOI21_X1   g08589(.A1(new_n9605_), .A2(new_n9606_), .B(new_n9563_), .ZN(new_n9607_));
  AOI21_X1   g08590(.A1(new_n9588_), .A2(new_n9550_), .B(new_n9607_), .ZN(new_n9608_));
  AOI21_X1   g08591(.A1(new_n9604_), .A2(new_n9608_), .B(new_n9599_), .ZN(new_n9609_));
  OAI21_X1   g08592(.A1(new_n9564_), .A2(new_n9566_), .B(new_n9576_), .ZN(new_n9610_));
  NAND2_X1   g08593(.A1(new_n9610_), .A2(new_n9579_), .ZN(new_n9611_));
  AOI21_X1   g08594(.A1(new_n9506_), .A2(new_n9531_), .B(new_n9579_), .ZN(new_n9612_));
  NOR3_X1    g08595(.A1(new_n9612_), .A2(new_n9556_), .A3(new_n9577_), .ZN(new_n9613_));
  NAND4_X1   g08596(.A1(new_n9594_), .A2(new_n9592_), .A3(new_n9593_), .A4(new_n9613_), .ZN(new_n9614_));
  OAI21_X1   g08597(.A1(new_n9551_), .A2(new_n9552_), .B(new_n9554_), .ZN(new_n9615_));
  NAND2_X1   g08598(.A1(new_n9615_), .A2(new_n9577_), .ZN(new_n9616_));
  INV_X1     g08599(.I(new_n9616_), .ZN(new_n9617_));
  NAND3_X1   g08600(.A1(new_n9563_), .A2(new_n9575_), .A3(new_n9582_), .ZN(new_n9618_));
  AOI21_X1   g08601(.A1(new_n9618_), .A2(new_n9614_), .B(new_n9617_), .ZN(new_n9619_));
  NAND2_X1   g08602(.A1(new_n9592_), .A2(new_n9593_), .ZN(new_n9620_));
  AOI21_X1   g08603(.A1(new_n9496_), .A2(new_n9540_), .B(new_n9595_), .ZN(new_n9621_));
  NOR3_X1    g08604(.A1(new_n9591_), .A2(new_n9620_), .A3(new_n9621_), .ZN(new_n9622_));
  NOR3_X1    g08605(.A1(new_n9622_), .A2(new_n9587_), .A3(new_n9616_), .ZN(new_n9623_));
  OAI21_X1   g08606(.A1(new_n9623_), .A2(new_n9619_), .B(new_n9611_), .ZN(new_n9624_));
  INV_X1     g08607(.I(new_n9611_), .ZN(new_n9625_));
  OAI21_X1   g08608(.A1(new_n9622_), .A2(new_n9587_), .B(new_n9616_), .ZN(new_n9626_));
  NAND3_X1   g08609(.A1(new_n9618_), .A2(new_n9614_), .A3(new_n9617_), .ZN(new_n9627_));
  NAND3_X1   g08610(.A1(new_n9626_), .A2(new_n9627_), .A3(new_n9625_), .ZN(new_n9628_));
  NAND2_X1   g08611(.A1(new_n9624_), .A2(new_n9628_), .ZN(new_n9629_));
  NOR2_X1    g08612(.A1(new_n9629_), .A2(new_n9609_), .ZN(new_n9630_));
  AOI22_X1   g08613(.A1(new_n9545_), .A2(new_n9548_), .B1(new_n9534_), .B2(new_n9541_), .ZN(new_n9631_));
  NOR2_X1    g08614(.A1(new_n9620_), .A2(new_n9621_), .ZN(new_n9632_));
  AOI21_X1   g08615(.A1(new_n9632_), .A2(new_n9614_), .B(new_n9591_), .ZN(new_n9633_));
  OAI21_X1   g08616(.A1(new_n9633_), .A2(new_n9607_), .B(new_n9631_), .ZN(new_n9634_));
  NAND2_X1   g08617(.A1(new_n9600_), .A2(new_n9452_), .ZN(new_n9635_));
  AOI22_X1   g08618(.A1(new_n9414_), .A2(new_n9418_), .B1(new_n9359_), .B2(new_n9355_), .ZN(new_n9636_));
  NOR4_X1    g08619(.A1(new_n9441_), .A2(new_n9433_), .A3(new_n9434_), .A4(new_n9448_), .ZN(new_n9637_));
  OAI21_X1   g08620(.A1(new_n9636_), .A2(new_n9637_), .B(new_n9429_), .ZN(new_n9638_));
  NAND2_X1   g08621(.A1(new_n9635_), .A2(new_n9638_), .ZN(new_n9639_));
  OAI21_X1   g08622(.A1(new_n9633_), .A2(new_n9631_), .B(new_n9598_), .ZN(new_n9640_));
  OAI21_X1   g08623(.A1(new_n9639_), .A2(new_n9640_), .B(new_n9634_), .ZN(new_n9641_));
  AOI21_X1   g08624(.A1(new_n9626_), .A2(new_n9627_), .B(new_n9625_), .ZN(new_n9642_));
  NOR3_X1    g08625(.A1(new_n9623_), .A2(new_n9619_), .A3(new_n9611_), .ZN(new_n9643_));
  NOR2_X1    g08626(.A1(new_n9643_), .A2(new_n9642_), .ZN(new_n9644_));
  NOR2_X1    g08627(.A1(new_n9644_), .A2(new_n9641_), .ZN(new_n9645_));
  OAI21_X1   g08628(.A1(new_n9630_), .A2(new_n9645_), .B(new_n9459_), .ZN(new_n9646_));
  OAI21_X1   g08629(.A1(new_n9457_), .A2(new_n9456_), .B(new_n9366_), .ZN(new_n9647_));
  NAND3_X1   g08630(.A1(new_n9431_), .A2(new_n9454_), .A3(new_n9367_), .ZN(new_n9648_));
  NAND2_X1   g08631(.A1(new_n9647_), .A2(new_n9648_), .ZN(new_n9649_));
  NAND3_X1   g08632(.A1(new_n9641_), .A2(new_n9624_), .A3(new_n9628_), .ZN(new_n9650_));
  NAND2_X1   g08633(.A1(new_n9629_), .A2(new_n9609_), .ZN(new_n9651_));
  NAND3_X1   g08634(.A1(new_n9651_), .A2(new_n9650_), .A3(new_n9649_), .ZN(new_n9652_));
  INV_X1     g08635(.I(\A[76] ), .ZN(new_n9653_));
  NOR2_X1    g08636(.A1(\A[77] ), .A2(\A[78] ), .ZN(new_n9654_));
  NAND2_X1   g08637(.A1(\A[77] ), .A2(\A[78] ), .ZN(new_n9655_));
  AOI21_X1   g08638(.A1(new_n9653_), .A2(new_n9655_), .B(new_n9654_), .ZN(new_n9656_));
  INV_X1     g08639(.I(\A[73] ), .ZN(new_n9657_));
  NOR2_X1    g08640(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n9658_));
  NAND2_X1   g08641(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n9659_));
  AOI21_X1   g08642(.A1(new_n9657_), .A2(new_n9659_), .B(new_n9658_), .ZN(new_n9660_));
  INV_X1     g08643(.I(new_n9660_), .ZN(new_n9661_));
  INV_X1     g08644(.I(\A[74] ), .ZN(new_n9662_));
  NAND2_X1   g08645(.A1(new_n9662_), .A2(\A[75] ), .ZN(new_n9663_));
  INV_X1     g08646(.I(\A[75] ), .ZN(new_n9664_));
  NAND2_X1   g08647(.A1(new_n9664_), .A2(\A[74] ), .ZN(new_n9665_));
  AOI21_X1   g08648(.A1(new_n9663_), .A2(new_n9665_), .B(new_n9657_), .ZN(new_n9666_));
  INV_X1     g08649(.I(new_n9658_), .ZN(new_n9667_));
  AOI21_X1   g08650(.A1(new_n9667_), .A2(new_n9659_), .B(\A[73] ), .ZN(new_n9668_));
  NOR2_X1    g08651(.A1(new_n9668_), .A2(new_n9666_), .ZN(new_n9669_));
  INV_X1     g08652(.I(\A[77] ), .ZN(new_n9670_));
  NAND2_X1   g08653(.A1(new_n9670_), .A2(\A[78] ), .ZN(new_n9671_));
  INV_X1     g08654(.I(\A[78] ), .ZN(new_n9672_));
  NAND2_X1   g08655(.A1(new_n9672_), .A2(\A[77] ), .ZN(new_n9673_));
  AOI21_X1   g08656(.A1(new_n9671_), .A2(new_n9673_), .B(new_n9653_), .ZN(new_n9674_));
  INV_X1     g08657(.I(new_n9654_), .ZN(new_n9675_));
  AOI21_X1   g08658(.A1(new_n9675_), .A2(new_n9655_), .B(\A[76] ), .ZN(new_n9676_));
  NOR2_X1    g08659(.A1(new_n9676_), .A2(new_n9674_), .ZN(new_n9677_));
  AOI21_X1   g08660(.A1(new_n9669_), .A2(new_n9677_), .B(new_n9661_), .ZN(new_n9678_));
  NOR2_X1    g08661(.A1(new_n9664_), .A2(\A[74] ), .ZN(new_n9679_));
  NOR2_X1    g08662(.A1(new_n9662_), .A2(\A[75] ), .ZN(new_n9680_));
  OAI21_X1   g08663(.A1(new_n9679_), .A2(new_n9680_), .B(\A[73] ), .ZN(new_n9681_));
  INV_X1     g08664(.I(new_n9659_), .ZN(new_n9682_));
  OAI21_X1   g08665(.A1(new_n9682_), .A2(new_n9658_), .B(new_n9657_), .ZN(new_n9683_));
  NAND2_X1   g08666(.A1(new_n9681_), .A2(new_n9683_), .ZN(new_n9684_));
  NOR2_X1    g08667(.A1(new_n9672_), .A2(\A[77] ), .ZN(new_n9685_));
  NOR2_X1    g08668(.A1(new_n9670_), .A2(\A[78] ), .ZN(new_n9686_));
  OAI21_X1   g08669(.A1(new_n9685_), .A2(new_n9686_), .B(\A[76] ), .ZN(new_n9687_));
  AND2_X2    g08670(.A1(\A[77] ), .A2(\A[78] ), .Z(new_n9688_));
  OAI21_X1   g08671(.A1(new_n9688_), .A2(new_n9654_), .B(new_n9653_), .ZN(new_n9689_));
  NAND2_X1   g08672(.A1(new_n9687_), .A2(new_n9689_), .ZN(new_n9690_));
  NOR3_X1    g08673(.A1(new_n9684_), .A2(new_n9690_), .A3(new_n9660_), .ZN(new_n9691_));
  OAI21_X1   g08674(.A1(new_n9678_), .A2(new_n9691_), .B(new_n9656_), .ZN(new_n9692_));
  INV_X1     g08675(.I(new_n9656_), .ZN(new_n9693_));
  OAI21_X1   g08676(.A1(new_n9684_), .A2(new_n9690_), .B(new_n9660_), .ZN(new_n9694_));
  NAND3_X1   g08677(.A1(new_n9669_), .A2(new_n9677_), .A3(new_n9661_), .ZN(new_n9695_));
  NAND3_X1   g08678(.A1(new_n9695_), .A2(new_n9694_), .A3(new_n9693_), .ZN(new_n9696_));
  INV_X1     g08679(.I(\A[69] ), .ZN(new_n9697_));
  NOR2_X1    g08680(.A1(new_n9697_), .A2(\A[68] ), .ZN(new_n9698_));
  INV_X1     g08681(.I(\A[68] ), .ZN(new_n9699_));
  NOR2_X1    g08682(.A1(new_n9699_), .A2(\A[69] ), .ZN(new_n9700_));
  OAI21_X1   g08683(.A1(new_n9698_), .A2(new_n9700_), .B(\A[67] ), .ZN(new_n9701_));
  INV_X1     g08684(.I(\A[67] ), .ZN(new_n9702_));
  NOR2_X1    g08685(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n9703_));
  NAND2_X1   g08686(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n9704_));
  INV_X1     g08687(.I(new_n9704_), .ZN(new_n9705_));
  OAI21_X1   g08688(.A1(new_n9705_), .A2(new_n9703_), .B(new_n9702_), .ZN(new_n9706_));
  NAND2_X1   g08689(.A1(new_n9701_), .A2(new_n9706_), .ZN(new_n9707_));
  INV_X1     g08690(.I(\A[70] ), .ZN(new_n9708_));
  INV_X1     g08691(.I(\A[71] ), .ZN(new_n9709_));
  NAND2_X1   g08692(.A1(new_n9709_), .A2(\A[72] ), .ZN(new_n9710_));
  INV_X1     g08693(.I(\A[72] ), .ZN(new_n9711_));
  NAND2_X1   g08694(.A1(new_n9711_), .A2(\A[71] ), .ZN(new_n9712_));
  AOI21_X1   g08695(.A1(new_n9710_), .A2(new_n9712_), .B(new_n9708_), .ZN(new_n9713_));
  OR2_X2     g08696(.A1(\A[71] ), .A2(\A[72] ), .Z(new_n9714_));
  NAND2_X1   g08697(.A1(\A[71] ), .A2(\A[72] ), .ZN(new_n9715_));
  AOI21_X1   g08698(.A1(new_n9714_), .A2(new_n9715_), .B(\A[70] ), .ZN(new_n9716_));
  NOR2_X1    g08699(.A1(new_n9713_), .A2(new_n9716_), .ZN(new_n9717_));
  NOR2_X1    g08700(.A1(new_n9707_), .A2(new_n9717_), .ZN(new_n9718_));
  NAND2_X1   g08701(.A1(new_n9699_), .A2(\A[69] ), .ZN(new_n9719_));
  NAND2_X1   g08702(.A1(new_n9697_), .A2(\A[68] ), .ZN(new_n9720_));
  AOI21_X1   g08703(.A1(new_n9719_), .A2(new_n9720_), .B(new_n9702_), .ZN(new_n9721_));
  INV_X1     g08704(.I(new_n9703_), .ZN(new_n9722_));
  AOI21_X1   g08705(.A1(new_n9722_), .A2(new_n9704_), .B(\A[67] ), .ZN(new_n9723_));
  NOR2_X1    g08706(.A1(new_n9723_), .A2(new_n9721_), .ZN(new_n9724_));
  NOR2_X1    g08707(.A1(new_n9711_), .A2(\A[71] ), .ZN(new_n9725_));
  NOR2_X1    g08708(.A1(new_n9709_), .A2(\A[72] ), .ZN(new_n9726_));
  OAI21_X1   g08709(.A1(new_n9725_), .A2(new_n9726_), .B(\A[70] ), .ZN(new_n9727_));
  NOR2_X1    g08710(.A1(\A[71] ), .A2(\A[72] ), .ZN(new_n9728_));
  INV_X1     g08711(.I(new_n9715_), .ZN(new_n9729_));
  OAI21_X1   g08712(.A1(new_n9729_), .A2(new_n9728_), .B(new_n9708_), .ZN(new_n9730_));
  NAND2_X1   g08713(.A1(new_n9727_), .A2(new_n9730_), .ZN(new_n9731_));
  NOR2_X1    g08714(.A1(new_n9724_), .A2(new_n9731_), .ZN(new_n9732_));
  NOR2_X1    g08715(.A1(new_n9732_), .A2(new_n9718_), .ZN(new_n9733_));
  NOR2_X1    g08716(.A1(new_n9677_), .A2(new_n9684_), .ZN(new_n9734_));
  NOR2_X1    g08717(.A1(new_n9669_), .A2(new_n9690_), .ZN(new_n9735_));
  NOR2_X1    g08718(.A1(new_n9734_), .A2(new_n9735_), .ZN(new_n9736_));
  NOR2_X1    g08719(.A1(new_n9733_), .A2(new_n9736_), .ZN(new_n9737_));
  NOR4_X1    g08720(.A1(new_n9721_), .A2(new_n9723_), .A3(new_n9713_), .A4(new_n9716_), .ZN(new_n9738_));
  AOI21_X1   g08721(.A1(new_n9708_), .A2(new_n9715_), .B(new_n9728_), .ZN(new_n9739_));
  AOI21_X1   g08722(.A1(new_n9702_), .A2(new_n9704_), .B(new_n9703_), .ZN(new_n9740_));
  NAND2_X1   g08723(.A1(new_n9739_), .A2(new_n9740_), .ZN(new_n9741_));
  INV_X1     g08724(.I(new_n9741_), .ZN(new_n9742_));
  NAND2_X1   g08725(.A1(new_n9738_), .A2(new_n9742_), .ZN(new_n9743_));
  NAND2_X1   g08726(.A1(new_n9656_), .A2(new_n9660_), .ZN(new_n9744_));
  AOI21_X1   g08727(.A1(new_n9684_), .A2(new_n9690_), .B(new_n9744_), .ZN(new_n9745_));
  NOR2_X1    g08728(.A1(new_n9743_), .A2(new_n9745_), .ZN(new_n9746_));
  NAND4_X1   g08729(.A1(new_n9737_), .A2(new_n9692_), .A3(new_n9746_), .A4(new_n9696_), .ZN(new_n9747_));
  INV_X1     g08730(.I(new_n9740_), .ZN(new_n9748_));
  NOR2_X1    g08731(.A1(new_n9738_), .A2(new_n9748_), .ZN(new_n9749_));
  NOR3_X1    g08732(.A1(new_n9707_), .A2(new_n9731_), .A3(new_n9740_), .ZN(new_n9750_));
  OAI21_X1   g08733(.A1(new_n9749_), .A2(new_n9750_), .B(new_n9739_), .ZN(new_n9751_));
  INV_X1     g08734(.I(new_n9739_), .ZN(new_n9752_));
  OAI21_X1   g08735(.A1(new_n9707_), .A2(new_n9731_), .B(new_n9740_), .ZN(new_n9753_));
  NAND3_X1   g08736(.A1(new_n9724_), .A2(new_n9717_), .A3(new_n9748_), .ZN(new_n9754_));
  NAND3_X1   g08737(.A1(new_n9753_), .A2(new_n9754_), .A3(new_n9752_), .ZN(new_n9755_));
  NAND2_X1   g08738(.A1(new_n9751_), .A2(new_n9755_), .ZN(new_n9756_));
  INV_X1     g08739(.I(new_n9756_), .ZN(new_n9757_));
  AOI21_X1   g08740(.A1(new_n9695_), .A2(new_n9694_), .B(new_n9693_), .ZN(new_n9758_));
  NOR3_X1    g08741(.A1(new_n9678_), .A2(new_n9691_), .A3(new_n9656_), .ZN(new_n9759_));
  NOR2_X1    g08742(.A1(new_n9759_), .A2(new_n9758_), .ZN(new_n9760_));
  NAND2_X1   g08743(.A1(new_n9724_), .A2(new_n9731_), .ZN(new_n9761_));
  NAND2_X1   g08744(.A1(new_n9707_), .A2(new_n9717_), .ZN(new_n9762_));
  NAND2_X1   g08745(.A1(new_n9761_), .A2(new_n9762_), .ZN(new_n9763_));
  NAND2_X1   g08746(.A1(new_n9669_), .A2(new_n9690_), .ZN(new_n9764_));
  NAND2_X1   g08747(.A1(new_n9677_), .A2(new_n9684_), .ZN(new_n9765_));
  NAND2_X1   g08748(.A1(new_n9765_), .A2(new_n9764_), .ZN(new_n9766_));
  NAND4_X1   g08749(.A1(new_n9681_), .A2(new_n9687_), .A3(new_n9683_), .A4(new_n9689_), .ZN(new_n9767_));
  NAND4_X1   g08750(.A1(new_n9701_), .A2(new_n9706_), .A3(new_n9727_), .A4(new_n9730_), .ZN(new_n9768_));
  NOR4_X1    g08751(.A1(new_n9768_), .A2(new_n9767_), .A3(new_n9741_), .A4(new_n9744_), .ZN(new_n9769_));
  NAND3_X1   g08752(.A1(new_n9763_), .A2(new_n9766_), .A3(new_n9769_), .ZN(new_n9770_));
  NAND2_X1   g08753(.A1(new_n9760_), .A2(new_n9770_), .ZN(new_n9771_));
  NAND3_X1   g08754(.A1(new_n9771_), .A2(new_n9747_), .A3(new_n9757_), .ZN(new_n9772_));
  INV_X1     g08755(.I(new_n9767_), .ZN(new_n9773_));
  INV_X1     g08756(.I(new_n9744_), .ZN(new_n9774_));
  NAND4_X1   g08757(.A1(new_n9773_), .A2(new_n9738_), .A3(new_n9742_), .A4(new_n9774_), .ZN(new_n9775_));
  NOR3_X1    g08758(.A1(new_n9775_), .A2(new_n9733_), .A3(new_n9736_), .ZN(new_n9776_));
  NOR2_X1    g08759(.A1(new_n9760_), .A2(new_n9776_), .ZN(new_n9777_));
  NAND2_X1   g08760(.A1(new_n9692_), .A2(new_n9696_), .ZN(new_n9778_));
  NOR2_X1    g08761(.A1(new_n9778_), .A2(new_n9770_), .ZN(new_n9779_));
  OAI21_X1   g08762(.A1(new_n9777_), .A2(new_n9779_), .B(new_n9757_), .ZN(new_n9780_));
  NAND2_X1   g08763(.A1(new_n9780_), .A2(new_n9772_), .ZN(new_n9781_));
  NAND2_X1   g08764(.A1(new_n9763_), .A2(new_n9766_), .ZN(new_n9782_));
  INV_X1     g08765(.I(new_n9746_), .ZN(new_n9783_));
  NOR3_X1    g08766(.A1(new_n9778_), .A2(new_n9782_), .A3(new_n9783_), .ZN(new_n9784_));
  NOR2_X1    g08767(.A1(new_n9776_), .A2(new_n9778_), .ZN(new_n9785_));
  NOR3_X1    g08768(.A1(new_n9784_), .A2(new_n9785_), .A3(new_n9756_), .ZN(new_n9786_));
  NAND2_X1   g08769(.A1(new_n9778_), .A2(new_n9770_), .ZN(new_n9787_));
  NAND3_X1   g08770(.A1(new_n9776_), .A2(new_n9692_), .A3(new_n9696_), .ZN(new_n9788_));
  AOI21_X1   g08771(.A1(new_n9788_), .A2(new_n9787_), .B(new_n9756_), .ZN(new_n9789_));
  NOR3_X1    g08772(.A1(new_n9736_), .A2(new_n9767_), .A3(new_n9744_), .ZN(new_n9790_));
  NAND3_X1   g08773(.A1(new_n9763_), .A2(new_n9738_), .A3(new_n9742_), .ZN(new_n9791_));
  NOR2_X1    g08774(.A1(new_n9790_), .A2(new_n9791_), .ZN(new_n9792_));
  NAND3_X1   g08775(.A1(new_n9766_), .A2(new_n9773_), .A3(new_n9774_), .ZN(new_n9793_));
  NOR2_X1    g08776(.A1(new_n9733_), .A2(new_n9743_), .ZN(new_n9794_));
  NOR2_X1    g08777(.A1(new_n9793_), .A2(new_n9794_), .ZN(new_n9795_));
  INV_X1     g08778(.I(\A[66] ), .ZN(new_n9796_));
  NOR2_X1    g08779(.A1(new_n9796_), .A2(\A[65] ), .ZN(new_n9797_));
  INV_X1     g08780(.I(\A[65] ), .ZN(new_n9798_));
  NOR2_X1    g08781(.A1(new_n9798_), .A2(\A[66] ), .ZN(new_n9799_));
  OAI21_X1   g08782(.A1(new_n9797_), .A2(new_n9799_), .B(\A[64] ), .ZN(new_n9800_));
  INV_X1     g08783(.I(\A[64] ), .ZN(new_n9801_));
  NOR2_X1    g08784(.A1(\A[65] ), .A2(\A[66] ), .ZN(new_n9802_));
  NAND2_X1   g08785(.A1(\A[65] ), .A2(\A[66] ), .ZN(new_n9803_));
  INV_X1     g08786(.I(new_n9803_), .ZN(new_n9804_));
  OAI21_X1   g08787(.A1(new_n9804_), .A2(new_n9802_), .B(new_n9801_), .ZN(new_n9805_));
  NAND2_X1   g08788(.A1(new_n9800_), .A2(new_n9805_), .ZN(new_n9806_));
  AOI21_X1   g08789(.A1(new_n9801_), .A2(new_n9803_), .B(new_n9802_), .ZN(new_n9807_));
  NAND4_X1   g08790(.A1(new_n9807_), .A2(\A[61] ), .A3(\A[62] ), .A4(\A[63] ), .ZN(new_n9808_));
  NOR2_X1    g08791(.A1(new_n9806_), .A2(new_n9808_), .ZN(new_n9809_));
  INV_X1     g08792(.I(\A[63] ), .ZN(new_n9810_));
  NOR2_X1    g08793(.A1(new_n9810_), .A2(\A[62] ), .ZN(new_n9811_));
  INV_X1     g08794(.I(\A[62] ), .ZN(new_n9812_));
  NOR2_X1    g08795(.A1(new_n9812_), .A2(\A[63] ), .ZN(new_n9813_));
  OAI21_X1   g08796(.A1(new_n9811_), .A2(new_n9813_), .B(\A[61] ), .ZN(new_n9814_));
  INV_X1     g08797(.I(\A[61] ), .ZN(new_n9815_));
  NOR2_X1    g08798(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n9816_));
  NAND2_X1   g08799(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n9817_));
  INV_X1     g08800(.I(new_n9817_), .ZN(new_n9818_));
  OAI21_X1   g08801(.A1(new_n9818_), .A2(new_n9816_), .B(new_n9815_), .ZN(new_n9819_));
  NAND2_X1   g08802(.A1(new_n9814_), .A2(new_n9819_), .ZN(new_n9820_));
  XOR2_X1    g08803(.A1(new_n9806_), .A2(new_n9820_), .Z(new_n9821_));
  INV_X1     g08804(.I(\A[55] ), .ZN(new_n9822_));
  INV_X1     g08805(.I(\A[56] ), .ZN(new_n9823_));
  NAND2_X1   g08806(.A1(new_n9823_), .A2(\A[57] ), .ZN(new_n9824_));
  INV_X1     g08807(.I(\A[57] ), .ZN(new_n9825_));
  NAND2_X1   g08808(.A1(new_n9825_), .A2(\A[56] ), .ZN(new_n9826_));
  AOI21_X1   g08809(.A1(new_n9824_), .A2(new_n9826_), .B(new_n9822_), .ZN(new_n9827_));
  NOR2_X1    g08810(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n9828_));
  INV_X1     g08811(.I(new_n9828_), .ZN(new_n9829_));
  NAND2_X1   g08812(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n9830_));
  AOI21_X1   g08813(.A1(new_n9829_), .A2(new_n9830_), .B(\A[55] ), .ZN(new_n9831_));
  NOR2_X1    g08814(.A1(new_n9831_), .A2(new_n9827_), .ZN(new_n9832_));
  INV_X1     g08815(.I(\A[58] ), .ZN(new_n9833_));
  INV_X1     g08816(.I(\A[59] ), .ZN(new_n9834_));
  NAND2_X1   g08817(.A1(new_n9834_), .A2(\A[60] ), .ZN(new_n9835_));
  INV_X1     g08818(.I(\A[60] ), .ZN(new_n9836_));
  NAND2_X1   g08819(.A1(new_n9836_), .A2(\A[59] ), .ZN(new_n9837_));
  AOI21_X1   g08820(.A1(new_n9835_), .A2(new_n9837_), .B(new_n9833_), .ZN(new_n9838_));
  NOR2_X1    g08821(.A1(\A[59] ), .A2(\A[60] ), .ZN(new_n9839_));
  INV_X1     g08822(.I(new_n9839_), .ZN(new_n9840_));
  NAND2_X1   g08823(.A1(\A[59] ), .A2(\A[60] ), .ZN(new_n9841_));
  AOI21_X1   g08824(.A1(new_n9840_), .A2(new_n9841_), .B(\A[58] ), .ZN(new_n9842_));
  NOR2_X1    g08825(.A1(new_n9842_), .A2(new_n9838_), .ZN(new_n9843_));
  AOI21_X1   g08826(.A1(new_n9833_), .A2(new_n9841_), .B(new_n9839_), .ZN(new_n9844_));
  AOI21_X1   g08827(.A1(new_n9822_), .A2(new_n9830_), .B(new_n9828_), .ZN(new_n9845_));
  NAND2_X1   g08828(.A1(new_n9844_), .A2(new_n9845_), .ZN(new_n9846_));
  NAND2_X1   g08829(.A1(new_n9821_), .A2(new_n9809_), .ZN(new_n9848_));
  INV_X1     g08830(.I(new_n9848_), .ZN(new_n9849_));
  OAI21_X1   g08831(.A1(new_n9792_), .A2(new_n9795_), .B(new_n9849_), .ZN(new_n9850_));
  OAI21_X1   g08832(.A1(new_n9786_), .A2(new_n9789_), .B(new_n9850_), .ZN(new_n9851_));
  NAND2_X1   g08833(.A1(new_n9793_), .A2(new_n9794_), .ZN(new_n9852_));
  NAND2_X1   g08834(.A1(new_n9790_), .A2(new_n9791_), .ZN(new_n9853_));
  AOI21_X1   g08835(.A1(new_n9853_), .A2(new_n9852_), .B(new_n9848_), .ZN(new_n9854_));
  NAND3_X1   g08836(.A1(new_n9780_), .A2(new_n9772_), .A3(new_n9854_), .ZN(new_n9855_));
  INV_X1     g08837(.I(new_n9845_), .ZN(new_n9856_));
  AOI21_X1   g08838(.A1(new_n9832_), .A2(new_n9843_), .B(new_n9856_), .ZN(new_n9857_));
  NOR2_X1    g08839(.A1(new_n9825_), .A2(\A[56] ), .ZN(new_n9858_));
  NOR2_X1    g08840(.A1(new_n9823_), .A2(\A[57] ), .ZN(new_n9859_));
  OAI21_X1   g08841(.A1(new_n9858_), .A2(new_n9859_), .B(\A[55] ), .ZN(new_n9860_));
  INV_X1     g08842(.I(new_n9830_), .ZN(new_n9861_));
  OAI21_X1   g08843(.A1(new_n9861_), .A2(new_n9828_), .B(new_n9822_), .ZN(new_n9862_));
  NAND2_X1   g08844(.A1(new_n9860_), .A2(new_n9862_), .ZN(new_n9863_));
  NOR2_X1    g08845(.A1(new_n9836_), .A2(\A[59] ), .ZN(new_n9864_));
  NOR2_X1    g08846(.A1(new_n9834_), .A2(\A[60] ), .ZN(new_n9865_));
  OAI21_X1   g08847(.A1(new_n9864_), .A2(new_n9865_), .B(\A[58] ), .ZN(new_n9866_));
  INV_X1     g08848(.I(new_n9841_), .ZN(new_n9867_));
  OAI21_X1   g08849(.A1(new_n9867_), .A2(new_n9839_), .B(new_n9833_), .ZN(new_n9868_));
  NAND2_X1   g08850(.A1(new_n9866_), .A2(new_n9868_), .ZN(new_n9869_));
  NOR3_X1    g08851(.A1(new_n9863_), .A2(new_n9869_), .A3(new_n9845_), .ZN(new_n9870_));
  OAI21_X1   g08852(.A1(new_n9857_), .A2(new_n9870_), .B(new_n9844_), .ZN(new_n9871_));
  INV_X1     g08853(.I(new_n9844_), .ZN(new_n9872_));
  OAI21_X1   g08854(.A1(new_n9863_), .A2(new_n9869_), .B(new_n9845_), .ZN(new_n9873_));
  NAND3_X1   g08855(.A1(new_n9832_), .A2(new_n9843_), .A3(new_n9856_), .ZN(new_n9874_));
  NAND3_X1   g08856(.A1(new_n9873_), .A2(new_n9874_), .A3(new_n9872_), .ZN(new_n9875_));
  NAND2_X1   g08857(.A1(new_n9871_), .A2(new_n9875_), .ZN(new_n9876_));
  NOR3_X1    g08858(.A1(new_n9863_), .A2(new_n9869_), .A3(new_n9846_), .ZN(new_n9877_));
  INV_X1     g08859(.I(new_n9877_), .ZN(new_n9878_));
  NAND2_X1   g08860(.A1(new_n9798_), .A2(\A[66] ), .ZN(new_n9879_));
  NAND2_X1   g08861(.A1(new_n9796_), .A2(\A[65] ), .ZN(new_n9880_));
  AOI21_X1   g08862(.A1(new_n9879_), .A2(new_n9880_), .B(new_n9801_), .ZN(new_n9881_));
  INV_X1     g08863(.I(new_n9802_), .ZN(new_n9882_));
  AOI21_X1   g08864(.A1(new_n9882_), .A2(new_n9803_), .B(\A[64] ), .ZN(new_n9883_));
  NOR2_X1    g08865(.A1(new_n9883_), .A2(new_n9881_), .ZN(new_n9884_));
  NAND2_X1   g08866(.A1(new_n9812_), .A2(\A[63] ), .ZN(new_n9885_));
  NAND2_X1   g08867(.A1(new_n9810_), .A2(\A[62] ), .ZN(new_n9886_));
  AOI21_X1   g08868(.A1(new_n9885_), .A2(new_n9886_), .B(new_n9815_), .ZN(new_n9887_));
  INV_X1     g08869(.I(new_n9816_), .ZN(new_n9888_));
  AOI21_X1   g08870(.A1(new_n9888_), .A2(new_n9817_), .B(\A[61] ), .ZN(new_n9889_));
  NOR2_X1    g08871(.A1(new_n9889_), .A2(new_n9887_), .ZN(new_n9890_));
  AOI21_X1   g08872(.A1(new_n9815_), .A2(new_n9817_), .B(new_n9816_), .ZN(new_n9891_));
  INV_X1     g08873(.I(new_n9891_), .ZN(new_n9892_));
  AOI21_X1   g08874(.A1(new_n9884_), .A2(new_n9890_), .B(new_n9892_), .ZN(new_n9893_));
  NOR3_X1    g08875(.A1(new_n9806_), .A2(new_n9820_), .A3(new_n9891_), .ZN(new_n9894_));
  OAI21_X1   g08876(.A1(new_n9893_), .A2(new_n9894_), .B(new_n9807_), .ZN(new_n9895_));
  INV_X1     g08877(.I(new_n9807_), .ZN(new_n9896_));
  OAI21_X1   g08878(.A1(new_n9806_), .A2(new_n9820_), .B(new_n9891_), .ZN(new_n9897_));
  NAND3_X1   g08879(.A1(new_n9884_), .A2(new_n9890_), .A3(new_n9892_), .ZN(new_n9898_));
  NAND3_X1   g08880(.A1(new_n9897_), .A2(new_n9898_), .A3(new_n9896_), .ZN(new_n9899_));
  NAND2_X1   g08881(.A1(new_n9895_), .A2(new_n9899_), .ZN(new_n9900_));
  NAND2_X1   g08882(.A1(new_n9832_), .A2(new_n9869_), .ZN(new_n9901_));
  NAND2_X1   g08883(.A1(new_n9843_), .A2(new_n9863_), .ZN(new_n9902_));
  NAND2_X1   g08884(.A1(new_n9901_), .A2(new_n9902_), .ZN(new_n9903_));
  NAND2_X1   g08885(.A1(new_n9821_), .A2(new_n9903_), .ZN(new_n9904_));
  NAND2_X1   g08886(.A1(new_n9807_), .A2(new_n9891_), .ZN(new_n9905_));
  AOI21_X1   g08887(.A1(new_n9806_), .A2(new_n9820_), .B(new_n9905_), .ZN(new_n9906_));
  NOR4_X1    g08888(.A1(new_n9900_), .A2(new_n9904_), .A3(new_n9878_), .A4(new_n9906_), .ZN(new_n9907_));
  NAND2_X1   g08889(.A1(new_n9907_), .A2(new_n9876_), .ZN(new_n9908_));
  XOR2_X1    g08890(.A1(new_n9884_), .A2(new_n9820_), .Z(new_n9909_));
  XOR2_X1    g08891(.A1(new_n9832_), .A2(new_n9869_), .Z(new_n9910_));
  NAND2_X1   g08892(.A1(new_n9877_), .A2(new_n9809_), .ZN(new_n9911_));
  NOR3_X1    g08893(.A1(new_n9909_), .A2(new_n9910_), .A3(new_n9911_), .ZN(new_n9912_));
  NAND2_X1   g08894(.A1(new_n9912_), .A2(new_n9876_), .ZN(new_n9913_));
  AOI21_X1   g08895(.A1(new_n9873_), .A2(new_n9874_), .B(new_n9872_), .ZN(new_n9914_));
  NOR3_X1    g08896(.A1(new_n9857_), .A2(new_n9870_), .A3(new_n9844_), .ZN(new_n9915_));
  NOR2_X1    g08897(.A1(new_n9915_), .A2(new_n9914_), .ZN(new_n9916_));
  NAND4_X1   g08898(.A1(new_n9821_), .A2(new_n9903_), .A3(new_n9809_), .A4(new_n9877_), .ZN(new_n9917_));
  AOI21_X1   g08899(.A1(new_n9917_), .A2(new_n9916_), .B(new_n9900_), .ZN(new_n9918_));
  AOI21_X1   g08900(.A1(new_n9897_), .A2(new_n9898_), .B(new_n9896_), .ZN(new_n9919_));
  NOR3_X1    g08901(.A1(new_n9893_), .A2(new_n9894_), .A3(new_n9807_), .ZN(new_n9920_));
  NOR2_X1    g08902(.A1(new_n9920_), .A2(new_n9919_), .ZN(new_n9921_));
  NOR3_X1    g08903(.A1(new_n9912_), .A2(new_n9921_), .A3(new_n9876_), .ZN(new_n9922_));
  OAI21_X1   g08904(.A1(new_n9922_), .A2(new_n9918_), .B(new_n9913_), .ZN(new_n9923_));
  NAND2_X1   g08905(.A1(new_n9923_), .A2(new_n9908_), .ZN(new_n9924_));
  AOI22_X1   g08906(.A1(new_n9924_), .A2(new_n9781_), .B1(new_n9851_), .B2(new_n9855_), .ZN(new_n9925_));
  OAI21_X1   g08907(.A1(new_n9656_), .A2(new_n9660_), .B(new_n9773_), .ZN(new_n9926_));
  NAND2_X1   g08908(.A1(new_n9926_), .A2(new_n9744_), .ZN(new_n9927_));
  INV_X1     g08909(.I(new_n9927_), .ZN(new_n9928_));
  OAI21_X1   g08910(.A1(new_n9739_), .A2(new_n9740_), .B(new_n9738_), .ZN(new_n9929_));
  NAND2_X1   g08911(.A1(new_n9929_), .A2(new_n9741_), .ZN(new_n9930_));
  AOI22_X1   g08912(.A1(new_n9760_), .A2(new_n9770_), .B1(new_n9751_), .B2(new_n9755_), .ZN(new_n9931_));
  OAI21_X1   g08913(.A1(new_n9931_), .A2(new_n9784_), .B(new_n9930_), .ZN(new_n9932_));
  INV_X1     g08914(.I(new_n9930_), .ZN(new_n9933_));
  OAI21_X1   g08915(.A1(new_n9778_), .A2(new_n9776_), .B(new_n9756_), .ZN(new_n9934_));
  NAND3_X1   g08916(.A1(new_n9934_), .A2(new_n9747_), .A3(new_n9933_), .ZN(new_n9935_));
  AOI21_X1   g08917(.A1(new_n9932_), .A2(new_n9935_), .B(new_n9928_), .ZN(new_n9936_));
  AOI21_X1   g08918(.A1(new_n9934_), .A2(new_n9747_), .B(new_n9933_), .ZN(new_n9937_));
  NOR3_X1    g08919(.A1(new_n9931_), .A2(new_n9784_), .A3(new_n9930_), .ZN(new_n9938_));
  NOR3_X1    g08920(.A1(new_n9938_), .A2(new_n9937_), .A3(new_n9927_), .ZN(new_n9939_));
  NOR2_X1    g08921(.A1(new_n9939_), .A2(new_n9936_), .ZN(new_n9940_));
  NAND2_X1   g08922(.A1(new_n9896_), .A2(new_n9892_), .ZN(new_n9941_));
  NAND3_X1   g08923(.A1(new_n9941_), .A2(new_n9884_), .A3(new_n9890_), .ZN(new_n9942_));
  NAND2_X1   g08924(.A1(new_n9942_), .A2(new_n9905_), .ZN(new_n9943_));
  NOR2_X1    g08925(.A1(new_n9909_), .A2(new_n9910_), .ZN(new_n9944_));
  NOR2_X1    g08926(.A1(new_n9878_), .A2(new_n9906_), .ZN(new_n9945_));
  NAND3_X1   g08927(.A1(new_n9921_), .A2(new_n9944_), .A3(new_n9945_), .ZN(new_n9946_));
  NAND2_X1   g08928(.A1(new_n9872_), .A2(new_n9856_), .ZN(new_n9947_));
  NAND3_X1   g08929(.A1(new_n9947_), .A2(new_n9832_), .A3(new_n9843_), .ZN(new_n9948_));
  NAND2_X1   g08930(.A1(new_n9948_), .A2(new_n9846_), .ZN(new_n9949_));
  INV_X1     g08931(.I(new_n9949_), .ZN(new_n9950_));
  OAI21_X1   g08932(.A1(new_n9912_), .A2(new_n9900_), .B(new_n9876_), .ZN(new_n9951_));
  AOI21_X1   g08933(.A1(new_n9951_), .A2(new_n9946_), .B(new_n9950_), .ZN(new_n9952_));
  AOI21_X1   g08934(.A1(new_n9917_), .A2(new_n9921_), .B(new_n9916_), .ZN(new_n9953_));
  NOR3_X1    g08935(.A1(new_n9953_), .A2(new_n9907_), .A3(new_n9949_), .ZN(new_n9954_));
  OAI21_X1   g08936(.A1(new_n9954_), .A2(new_n9952_), .B(new_n9943_), .ZN(new_n9955_));
  INV_X1     g08937(.I(new_n9943_), .ZN(new_n9956_));
  OAI21_X1   g08938(.A1(new_n9953_), .A2(new_n9907_), .B(new_n9949_), .ZN(new_n9957_));
  NAND3_X1   g08939(.A1(new_n9951_), .A2(new_n9946_), .A3(new_n9950_), .ZN(new_n9958_));
  NAND3_X1   g08940(.A1(new_n9957_), .A2(new_n9958_), .A3(new_n9956_), .ZN(new_n9959_));
  NAND2_X1   g08941(.A1(new_n9955_), .A2(new_n9959_), .ZN(new_n9960_));
  NOR2_X1    g08942(.A1(new_n9960_), .A2(new_n9940_), .ZN(new_n9961_));
  OAI21_X1   g08943(.A1(new_n9938_), .A2(new_n9937_), .B(new_n9927_), .ZN(new_n9962_));
  NAND3_X1   g08944(.A1(new_n9932_), .A2(new_n9935_), .A3(new_n9928_), .ZN(new_n9963_));
  NAND2_X1   g08945(.A1(new_n9962_), .A2(new_n9963_), .ZN(new_n9964_));
  AOI21_X1   g08946(.A1(new_n9957_), .A2(new_n9958_), .B(new_n9956_), .ZN(new_n9965_));
  NOR3_X1    g08947(.A1(new_n9954_), .A2(new_n9952_), .A3(new_n9943_), .ZN(new_n9966_));
  NOR2_X1    g08948(.A1(new_n9966_), .A2(new_n9965_), .ZN(new_n9967_));
  NOR2_X1    g08949(.A1(new_n9967_), .A2(new_n9964_), .ZN(new_n9968_));
  OAI21_X1   g08950(.A1(new_n9961_), .A2(new_n9968_), .B(new_n9925_), .ZN(new_n9969_));
  NOR2_X1    g08951(.A1(new_n9786_), .A2(new_n9789_), .ZN(new_n9970_));
  AOI21_X1   g08952(.A1(new_n9780_), .A2(new_n9772_), .B(new_n9854_), .ZN(new_n9971_));
  NOR3_X1    g08953(.A1(new_n9786_), .A2(new_n9789_), .A3(new_n9850_), .ZN(new_n9972_));
  OAI21_X1   g08954(.A1(new_n9912_), .A2(new_n9876_), .B(new_n9921_), .ZN(new_n9973_));
  NAND3_X1   g08955(.A1(new_n9917_), .A2(new_n9916_), .A3(new_n9900_), .ZN(new_n9974_));
  NAND2_X1   g08956(.A1(new_n9973_), .A2(new_n9974_), .ZN(new_n9975_));
  AOI22_X1   g08957(.A1(new_n9975_), .A2(new_n9913_), .B1(new_n9876_), .B2(new_n9907_), .ZN(new_n9976_));
  OAI22_X1   g08958(.A1(new_n9976_), .A2(new_n9970_), .B1(new_n9972_), .B2(new_n9971_), .ZN(new_n9977_));
  NOR2_X1    g08959(.A1(new_n9960_), .A2(new_n9964_), .ZN(new_n9978_));
  AOI22_X1   g08960(.A1(new_n9955_), .A2(new_n9959_), .B1(new_n9962_), .B2(new_n9963_), .ZN(new_n9979_));
  OAI21_X1   g08961(.A1(new_n9978_), .A2(new_n9979_), .B(new_n9977_), .ZN(new_n9980_));
  NAND4_X1   g08962(.A1(new_n9969_), .A2(new_n9646_), .A3(new_n9980_), .A4(new_n9652_), .ZN(new_n9981_));
  NOR3_X1    g08963(.A1(new_n9924_), .A2(new_n9971_), .A3(new_n9972_), .ZN(new_n9982_));
  NAND3_X1   g08964(.A1(new_n9976_), .A2(new_n9851_), .A3(new_n9855_), .ZN(new_n9983_));
  NOR2_X1    g08965(.A1(new_n9792_), .A2(new_n9795_), .ZN(new_n9984_));
  INV_X1     g08966(.I(new_n9809_), .ZN(new_n9985_));
  NOR2_X1    g08967(.A1(new_n9909_), .A2(new_n9985_), .ZN(new_n9986_));
  NOR2_X1    g08968(.A1(new_n9984_), .A2(new_n9986_), .ZN(new_n9987_));
  AND2_X2    g08969(.A1(new_n9984_), .A2(new_n9986_), .Z(new_n9988_));
  AOI21_X1   g08970(.A1(new_n9534_), .A2(new_n9541_), .B(new_n9544_), .ZN(new_n9989_));
  NOR2_X1    g08971(.A1(new_n9542_), .A2(new_n9547_), .ZN(new_n9990_));
  NOR2_X1    g08972(.A1(new_n9990_), .A2(new_n9989_), .ZN(new_n9991_));
  NOR2_X1    g08973(.A1(new_n9991_), .A2(new_n9546_), .ZN(new_n9992_));
  NOR3_X1    g08974(.A1(new_n9990_), .A2(new_n9543_), .A3(new_n9989_), .ZN(new_n9993_));
  NOR4_X1    g08975(.A1(new_n9992_), .A2(new_n9988_), .A3(new_n9987_), .A4(new_n9993_), .ZN(new_n9994_));
  INV_X1     g08976(.I(new_n9994_), .ZN(new_n9995_));
  NAND2_X1   g08977(.A1(new_n9995_), .A2(new_n9983_), .ZN(new_n9996_));
  NAND2_X1   g08978(.A1(new_n9982_), .A2(new_n9994_), .ZN(new_n9997_));
  NAND2_X1   g08979(.A1(new_n9996_), .A2(new_n9997_), .ZN(new_n9998_));
  OAI21_X1   g08980(.A1(new_n9633_), .A2(new_n9607_), .B(new_n9550_), .ZN(new_n9999_));
  NAND3_X1   g08981(.A1(new_n9588_), .A2(new_n9631_), .A3(new_n9598_), .ZN(new_n10000_));
  NAND2_X1   g08982(.A1(new_n9999_), .A2(new_n10000_), .ZN(new_n10001_));
  XOR2_X1    g08983(.A1(new_n10001_), .A2(new_n9639_), .Z(new_n10002_));
  OAI21_X1   g08984(.A1(new_n9982_), .A2(new_n10002_), .B(new_n9998_), .ZN(new_n10003_));
  AOI21_X1   g08985(.A1(new_n9651_), .A2(new_n9650_), .B(new_n9649_), .ZN(new_n10004_));
  NOR3_X1    g08986(.A1(new_n9630_), .A2(new_n9645_), .A3(new_n9459_), .ZN(new_n10005_));
  NOR2_X1    g08987(.A1(new_n10005_), .A2(new_n10004_), .ZN(new_n10006_));
  NAND2_X1   g08988(.A1(new_n9967_), .A2(new_n9964_), .ZN(new_n10007_));
  NAND2_X1   g08989(.A1(new_n9960_), .A2(new_n9940_), .ZN(new_n10008_));
  AOI21_X1   g08990(.A1(new_n10008_), .A2(new_n10007_), .B(new_n9977_), .ZN(new_n10009_));
  NAND4_X1   g08991(.A1(new_n9955_), .A2(new_n9959_), .A3(new_n9962_), .A4(new_n9963_), .ZN(new_n10010_));
  NAND2_X1   g08992(.A1(new_n9960_), .A2(new_n9964_), .ZN(new_n10011_));
  AOI21_X1   g08993(.A1(new_n10011_), .A2(new_n10010_), .B(new_n9925_), .ZN(new_n10012_));
  NOR2_X1    g08994(.A1(new_n10009_), .A2(new_n10012_), .ZN(new_n10013_));
  NOR2_X1    g08995(.A1(new_n10013_), .A2(new_n10006_), .ZN(new_n10014_));
  OAI21_X1   g08996(.A1(new_n10014_), .A2(new_n10003_), .B(new_n9981_), .ZN(new_n10015_));
  NOR2_X1    g08997(.A1(new_n9928_), .A2(new_n9933_), .ZN(new_n10016_));
  NAND2_X1   g08998(.A1(new_n9934_), .A2(new_n9747_), .ZN(new_n10017_));
  AOI21_X1   g08999(.A1(new_n9928_), .A2(new_n9933_), .B(new_n10017_), .ZN(new_n10018_));
  NOR2_X1    g09000(.A1(new_n10018_), .A2(new_n10016_), .ZN(new_n10019_));
  INV_X1     g09001(.I(new_n10019_), .ZN(new_n10020_));
  NOR2_X1    g09002(.A1(new_n9956_), .A2(new_n9950_), .ZN(new_n10021_));
  NAND2_X1   g09003(.A1(new_n9951_), .A2(new_n9946_), .ZN(new_n10022_));
  AOI21_X1   g09004(.A1(new_n9956_), .A2(new_n9950_), .B(new_n10022_), .ZN(new_n10023_));
  NOR2_X1    g09005(.A1(new_n10023_), .A2(new_n10021_), .ZN(new_n10024_));
  NAND2_X1   g09006(.A1(new_n10010_), .A2(new_n9977_), .ZN(new_n10025_));
  XOR2_X1    g09007(.A1(new_n9927_), .A2(new_n9930_), .Z(new_n10026_));
  XNOR2_X1   g09008(.A1(new_n9943_), .A2(new_n9949_), .ZN(new_n10027_));
  INV_X1     g09009(.I(new_n10027_), .ZN(new_n10028_));
  NOR4_X1    g09010(.A1(new_n10022_), .A2(new_n10026_), .A3(new_n10017_), .A4(new_n10028_), .ZN(new_n10029_));
  AOI21_X1   g09011(.A1(new_n10025_), .A2(new_n10029_), .B(new_n10024_), .ZN(new_n10030_));
  INV_X1     g09012(.I(new_n10024_), .ZN(new_n10031_));
  AOI21_X1   g09013(.A1(new_n9940_), .A2(new_n9967_), .B(new_n9925_), .ZN(new_n10032_));
  INV_X1     g09014(.I(new_n10029_), .ZN(new_n10033_));
  NOR3_X1    g09015(.A1(new_n10032_), .A2(new_n10031_), .A3(new_n10033_), .ZN(new_n10034_));
  OAI21_X1   g09016(.A1(new_n10034_), .A2(new_n10030_), .B(new_n10020_), .ZN(new_n10035_));
  OAI21_X1   g09017(.A1(new_n10032_), .A2(new_n10033_), .B(new_n10031_), .ZN(new_n10036_));
  NAND3_X1   g09018(.A1(new_n10025_), .A2(new_n10024_), .A3(new_n10029_), .ZN(new_n10037_));
  NAND3_X1   g09019(.A1(new_n10036_), .A2(new_n10037_), .A3(new_n10019_), .ZN(new_n10038_));
  NAND2_X1   g09020(.A1(new_n10035_), .A2(new_n10038_), .ZN(new_n10039_));
  NOR2_X1    g09021(.A1(new_n9617_), .A2(new_n9625_), .ZN(new_n10040_));
  NAND2_X1   g09022(.A1(new_n9618_), .A2(new_n9614_), .ZN(new_n10041_));
  AOI21_X1   g09023(.A1(new_n9625_), .A2(new_n9617_), .B(new_n10041_), .ZN(new_n10042_));
  NOR2_X1    g09024(.A1(new_n10042_), .A2(new_n10040_), .ZN(new_n10043_));
  NAND2_X1   g09025(.A1(new_n9366_), .A2(new_n9393_), .ZN(new_n10044_));
  NOR2_X1    g09026(.A1(new_n9430_), .A2(new_n9417_), .ZN(new_n10045_));
  OAI21_X1   g09027(.A1(new_n9366_), .A2(new_n9393_), .B(new_n10045_), .ZN(new_n10046_));
  NAND2_X1   g09028(.A1(new_n10046_), .A2(new_n10044_), .ZN(new_n10047_));
  AOI21_X1   g09029(.A1(new_n9459_), .A2(new_n9644_), .B(new_n9609_), .ZN(new_n10048_));
  INV_X1     g09030(.I(new_n10045_), .ZN(new_n10049_));
  XOR2_X1    g09031(.A1(new_n9366_), .A2(new_n9393_), .Z(new_n10050_));
  XOR2_X1    g09032(.A1(new_n9616_), .A2(new_n9611_), .Z(new_n10051_));
  NOR4_X1    g09033(.A1(new_n10050_), .A2(new_n10049_), .A3(new_n10041_), .A4(new_n10051_), .ZN(new_n10052_));
  INV_X1     g09034(.I(new_n10052_), .ZN(new_n10053_));
  OAI21_X1   g09035(.A1(new_n10048_), .A2(new_n10053_), .B(new_n10047_), .ZN(new_n10054_));
  INV_X1     g09036(.I(new_n10047_), .ZN(new_n10055_));
  OAI21_X1   g09037(.A1(new_n9649_), .A2(new_n9629_), .B(new_n9641_), .ZN(new_n10056_));
  NAND3_X1   g09038(.A1(new_n10056_), .A2(new_n10052_), .A3(new_n10055_), .ZN(new_n10057_));
  AOI21_X1   g09039(.A1(new_n10054_), .A2(new_n10057_), .B(new_n10043_), .ZN(new_n10058_));
  INV_X1     g09040(.I(new_n10043_), .ZN(new_n10059_));
  AOI21_X1   g09041(.A1(new_n10056_), .A2(new_n10052_), .B(new_n10055_), .ZN(new_n10060_));
  NOR3_X1    g09042(.A1(new_n10048_), .A2(new_n10047_), .A3(new_n10053_), .ZN(new_n10061_));
  NOR3_X1    g09043(.A1(new_n10061_), .A2(new_n10060_), .A3(new_n10059_), .ZN(new_n10062_));
  NOR2_X1    g09044(.A1(new_n10062_), .A2(new_n10058_), .ZN(new_n10063_));
  NOR2_X1    g09045(.A1(new_n10039_), .A2(new_n10063_), .ZN(new_n10064_));
  OAI21_X1   g09046(.A1(new_n10061_), .A2(new_n10060_), .B(new_n10059_), .ZN(new_n10065_));
  NAND3_X1   g09047(.A1(new_n10054_), .A2(new_n10057_), .A3(new_n10043_), .ZN(new_n10066_));
  NAND2_X1   g09048(.A1(new_n10065_), .A2(new_n10066_), .ZN(new_n10067_));
  AOI21_X1   g09049(.A1(new_n10035_), .A2(new_n10038_), .B(new_n10067_), .ZN(new_n10068_));
  OAI21_X1   g09050(.A1(new_n10068_), .A2(new_n10064_), .B(new_n10015_), .ZN(new_n10069_));
  NOR4_X1    g09051(.A1(new_n10009_), .A2(new_n10005_), .A3(new_n10012_), .A4(new_n10004_), .ZN(new_n10070_));
  XOR2_X1    g09052(.A1(new_n9982_), .A2(new_n9994_), .Z(new_n10071_));
  INV_X1     g09053(.I(new_n10002_), .ZN(new_n10072_));
  AOI21_X1   g09054(.A1(new_n9983_), .A2(new_n10072_), .B(new_n10071_), .ZN(new_n10073_));
  NAND2_X1   g09055(.A1(new_n9646_), .A2(new_n9652_), .ZN(new_n10074_));
  NAND2_X1   g09056(.A1(new_n9969_), .A2(new_n9980_), .ZN(new_n10075_));
  NAND2_X1   g09057(.A1(new_n10075_), .A2(new_n10074_), .ZN(new_n10076_));
  AOI21_X1   g09058(.A1(new_n10076_), .A2(new_n10073_), .B(new_n10070_), .ZN(new_n10077_));
  AOI21_X1   g09059(.A1(new_n10036_), .A2(new_n10037_), .B(new_n10019_), .ZN(new_n10078_));
  NOR3_X1    g09060(.A1(new_n10034_), .A2(new_n10030_), .A3(new_n10020_), .ZN(new_n10079_));
  NOR4_X1    g09061(.A1(new_n10079_), .A2(new_n10078_), .A3(new_n10058_), .A4(new_n10062_), .ZN(new_n10080_));
  AOI22_X1   g09062(.A1(new_n10035_), .A2(new_n10038_), .B1(new_n10065_), .B2(new_n10066_), .ZN(new_n10081_));
  OAI21_X1   g09063(.A1(new_n10080_), .A2(new_n10081_), .B(new_n10077_), .ZN(new_n10082_));
  INV_X1     g09064(.I(\A[16] ), .ZN(new_n10083_));
  NOR2_X1    g09065(.A1(\A[17] ), .A2(\A[18] ), .ZN(new_n10084_));
  NAND2_X1   g09066(.A1(\A[17] ), .A2(\A[18] ), .ZN(new_n10085_));
  AOI21_X1   g09067(.A1(new_n10083_), .A2(new_n10085_), .B(new_n10084_), .ZN(new_n10086_));
  NOR2_X1    g09068(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n10087_));
  INV_X1     g09069(.I(new_n10087_), .ZN(new_n10088_));
  INV_X1     g09070(.I(\A[14] ), .ZN(new_n10089_));
  INV_X1     g09071(.I(\A[15] ), .ZN(new_n10090_));
  NOR2_X1    g09072(.A1(new_n10089_), .A2(new_n10090_), .ZN(new_n10091_));
  OAI21_X1   g09073(.A1(\A[13] ), .A2(new_n10091_), .B(new_n10088_), .ZN(new_n10092_));
  INV_X1     g09074(.I(new_n10092_), .ZN(new_n10093_));
  NAND2_X1   g09075(.A1(new_n10093_), .A2(new_n10086_), .ZN(new_n10094_));
  INV_X1     g09076(.I(new_n10086_), .ZN(new_n10095_));
  NAND2_X1   g09077(.A1(new_n10095_), .A2(new_n10092_), .ZN(new_n10096_));
  NOR2_X1    g09078(.A1(new_n10090_), .A2(\A[14] ), .ZN(new_n10097_));
  NOR2_X1    g09079(.A1(new_n10089_), .A2(\A[15] ), .ZN(new_n10098_));
  OAI21_X1   g09080(.A1(new_n10097_), .A2(new_n10098_), .B(\A[13] ), .ZN(new_n10099_));
  INV_X1     g09081(.I(\A[13] ), .ZN(new_n10100_));
  OAI21_X1   g09082(.A1(new_n10091_), .A2(new_n10087_), .B(new_n10100_), .ZN(new_n10101_));
  AND2_X2    g09083(.A1(new_n10101_), .A2(new_n10099_), .Z(new_n10102_));
  INV_X1     g09084(.I(\A[17] ), .ZN(new_n10103_));
  NAND2_X1   g09085(.A1(new_n10103_), .A2(\A[18] ), .ZN(new_n10104_));
  INV_X1     g09086(.I(\A[18] ), .ZN(new_n10105_));
  NAND2_X1   g09087(.A1(new_n10105_), .A2(\A[17] ), .ZN(new_n10106_));
  AOI21_X1   g09088(.A1(new_n10104_), .A2(new_n10106_), .B(new_n10083_), .ZN(new_n10107_));
  INV_X1     g09089(.I(new_n10084_), .ZN(new_n10108_));
  AOI21_X1   g09090(.A1(new_n10108_), .A2(new_n10085_), .B(\A[16] ), .ZN(new_n10109_));
  NOR2_X1    g09091(.A1(new_n10109_), .A2(new_n10107_), .ZN(new_n10110_));
  NAND3_X1   g09092(.A1(new_n10102_), .A2(new_n10096_), .A3(new_n10110_), .ZN(new_n10111_));
  NAND2_X1   g09093(.A1(new_n10111_), .A2(new_n10094_), .ZN(new_n10112_));
  NOR2_X1    g09094(.A1(\A[11] ), .A2(\A[12] ), .ZN(new_n10113_));
  INV_X1     g09095(.I(\A[11] ), .ZN(new_n10114_));
  INV_X1     g09096(.I(\A[12] ), .ZN(new_n10115_));
  NOR2_X1    g09097(.A1(new_n10114_), .A2(new_n10115_), .ZN(new_n10116_));
  NOR2_X1    g09098(.A1(new_n10116_), .A2(\A[10] ), .ZN(new_n10117_));
  NOR2_X1    g09099(.A1(new_n10117_), .A2(new_n10113_), .ZN(new_n10118_));
  NOR2_X1    g09100(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n10119_));
  INV_X1     g09101(.I(\A[8] ), .ZN(new_n10120_));
  INV_X1     g09102(.I(\A[9] ), .ZN(new_n10121_));
  NOR2_X1    g09103(.A1(new_n10120_), .A2(new_n10121_), .ZN(new_n10122_));
  NOR2_X1    g09104(.A1(new_n10122_), .A2(\A[7] ), .ZN(new_n10123_));
  NOR2_X1    g09105(.A1(new_n10123_), .A2(new_n10119_), .ZN(new_n10124_));
  NAND2_X1   g09106(.A1(new_n10118_), .A2(new_n10124_), .ZN(new_n10125_));
  NOR2_X1    g09107(.A1(new_n10121_), .A2(\A[8] ), .ZN(new_n10126_));
  NOR2_X1    g09108(.A1(new_n10120_), .A2(\A[9] ), .ZN(new_n10127_));
  OAI21_X1   g09109(.A1(new_n10126_), .A2(new_n10127_), .B(\A[7] ), .ZN(new_n10128_));
  INV_X1     g09110(.I(\A[7] ), .ZN(new_n10129_));
  OAI21_X1   g09111(.A1(new_n10122_), .A2(new_n10119_), .B(new_n10129_), .ZN(new_n10130_));
  NOR2_X1    g09112(.A1(new_n10115_), .A2(\A[11] ), .ZN(new_n10131_));
  NOR2_X1    g09113(.A1(new_n10114_), .A2(\A[12] ), .ZN(new_n10132_));
  OAI21_X1   g09114(.A1(new_n10131_), .A2(new_n10132_), .B(\A[10] ), .ZN(new_n10133_));
  INV_X1     g09115(.I(\A[10] ), .ZN(new_n10134_));
  OAI21_X1   g09116(.A1(new_n10116_), .A2(new_n10113_), .B(new_n10134_), .ZN(new_n10135_));
  NAND4_X1   g09117(.A1(new_n10128_), .A2(new_n10130_), .A3(new_n10135_), .A4(new_n10133_), .ZN(new_n10136_));
  INV_X1     g09118(.I(new_n10136_), .ZN(new_n10137_));
  OAI21_X1   g09119(.A1(new_n10118_), .A2(new_n10124_), .B(new_n10137_), .ZN(new_n10138_));
  NAND2_X1   g09120(.A1(new_n10138_), .A2(new_n10125_), .ZN(new_n10139_));
  INV_X1     g09121(.I(new_n10139_), .ZN(new_n10140_));
  INV_X1     g09122(.I(new_n10124_), .ZN(new_n10141_));
  NAND2_X1   g09123(.A1(new_n10130_), .A2(new_n10128_), .ZN(new_n10142_));
  INV_X1     g09124(.I(new_n10142_), .ZN(new_n10143_));
  AND2_X2    g09125(.A1(new_n10135_), .A2(new_n10133_), .Z(new_n10144_));
  AOI21_X1   g09126(.A1(new_n10143_), .A2(new_n10144_), .B(new_n10141_), .ZN(new_n10145_));
  NOR2_X1    g09127(.A1(new_n10136_), .A2(new_n10124_), .ZN(new_n10146_));
  OAI21_X1   g09128(.A1(new_n10145_), .A2(new_n10146_), .B(new_n10118_), .ZN(new_n10147_));
  INV_X1     g09129(.I(new_n10118_), .ZN(new_n10148_));
  NAND2_X1   g09130(.A1(new_n10136_), .A2(new_n10124_), .ZN(new_n10149_));
  NAND3_X1   g09131(.A1(new_n10143_), .A2(new_n10144_), .A3(new_n10141_), .ZN(new_n10150_));
  NAND3_X1   g09132(.A1(new_n10150_), .A2(new_n10148_), .A3(new_n10149_), .ZN(new_n10151_));
  NAND2_X1   g09133(.A1(new_n10147_), .A2(new_n10151_), .ZN(new_n10152_));
  AOI21_X1   g09134(.A1(new_n10102_), .A2(new_n10110_), .B(new_n10092_), .ZN(new_n10153_));
  NAND2_X1   g09135(.A1(new_n10101_), .A2(new_n10099_), .ZN(new_n10154_));
  NOR2_X1    g09136(.A1(new_n10105_), .A2(\A[17] ), .ZN(new_n10155_));
  NOR2_X1    g09137(.A1(new_n10103_), .A2(\A[18] ), .ZN(new_n10156_));
  OAI21_X1   g09138(.A1(new_n10155_), .A2(new_n10156_), .B(\A[16] ), .ZN(new_n10157_));
  INV_X1     g09139(.I(new_n10085_), .ZN(new_n10158_));
  OAI21_X1   g09140(.A1(new_n10158_), .A2(new_n10084_), .B(new_n10083_), .ZN(new_n10159_));
  NAND2_X1   g09141(.A1(new_n10157_), .A2(new_n10159_), .ZN(new_n10160_));
  NOR3_X1    g09142(.A1(new_n10154_), .A2(new_n10160_), .A3(new_n10093_), .ZN(new_n10161_));
  OAI21_X1   g09143(.A1(new_n10153_), .A2(new_n10161_), .B(new_n10086_), .ZN(new_n10162_));
  OAI21_X1   g09144(.A1(new_n10154_), .A2(new_n10160_), .B(new_n10093_), .ZN(new_n10163_));
  NAND3_X1   g09145(.A1(new_n10102_), .A2(new_n10092_), .A3(new_n10110_), .ZN(new_n10164_));
  NAND3_X1   g09146(.A1(new_n10164_), .A2(new_n10095_), .A3(new_n10163_), .ZN(new_n10165_));
  NAND2_X1   g09147(.A1(new_n10162_), .A2(new_n10165_), .ZN(new_n10166_));
  NAND2_X1   g09148(.A1(new_n10135_), .A2(new_n10133_), .ZN(new_n10167_));
  XNOR2_X1   g09149(.A1(new_n10142_), .A2(new_n10167_), .ZN(new_n10168_));
  XOR2_X1    g09150(.A1(new_n10110_), .A2(new_n10154_), .Z(new_n10169_));
  NAND4_X1   g09151(.A1(new_n10086_), .A2(\A[13] ), .A3(\A[14] ), .A4(\A[15] ), .ZN(new_n10170_));
  NOR2_X1    g09152(.A1(new_n10160_), .A2(new_n10170_), .ZN(new_n10171_));
  NOR2_X1    g09153(.A1(new_n10125_), .A2(new_n10136_), .ZN(new_n10172_));
  NAND2_X1   g09154(.A1(new_n10172_), .A2(new_n10171_), .ZN(new_n10173_));
  NOR3_X1    g09155(.A1(new_n10168_), .A2(new_n10173_), .A3(new_n10169_), .ZN(new_n10174_));
  OAI21_X1   g09156(.A1(new_n10166_), .A2(new_n10174_), .B(new_n10152_), .ZN(new_n10175_));
  AOI21_X1   g09157(.A1(new_n10164_), .A2(new_n10163_), .B(new_n10095_), .ZN(new_n10176_));
  NOR3_X1    g09158(.A1(new_n10153_), .A2(new_n10086_), .A3(new_n10161_), .ZN(new_n10177_));
  NOR2_X1    g09159(.A1(new_n10177_), .A2(new_n10176_), .ZN(new_n10178_));
  NOR2_X1    g09160(.A1(new_n10168_), .A2(new_n10169_), .ZN(new_n10179_));
  INV_X1     g09161(.I(new_n10172_), .ZN(new_n10180_));
  AOI21_X1   g09162(.A1(new_n10154_), .A2(new_n10160_), .B(new_n10094_), .ZN(new_n10181_));
  NOR2_X1    g09163(.A1(new_n10180_), .A2(new_n10181_), .ZN(new_n10182_));
  NAND3_X1   g09164(.A1(new_n10178_), .A2(new_n10179_), .A3(new_n10182_), .ZN(new_n10183_));
  AOI21_X1   g09165(.A1(new_n10175_), .A2(new_n10183_), .B(new_n10140_), .ZN(new_n10184_));
  AOI21_X1   g09166(.A1(new_n10150_), .A2(new_n10149_), .B(new_n10148_), .ZN(new_n10185_));
  NOR3_X1    g09167(.A1(new_n10145_), .A2(new_n10118_), .A3(new_n10146_), .ZN(new_n10186_));
  NOR2_X1    g09168(.A1(new_n10186_), .A2(new_n10185_), .ZN(new_n10187_));
  XOR2_X1    g09169(.A1(new_n10142_), .A2(new_n10167_), .Z(new_n10188_));
  XOR2_X1    g09170(.A1(new_n10154_), .A2(new_n10160_), .Z(new_n10189_));
  NAND4_X1   g09171(.A1(new_n10188_), .A2(new_n10189_), .A3(new_n10171_), .A4(new_n10172_), .ZN(new_n10190_));
  AOI21_X1   g09172(.A1(new_n10178_), .A2(new_n10190_), .B(new_n10187_), .ZN(new_n10191_));
  NAND2_X1   g09173(.A1(new_n10188_), .A2(new_n10189_), .ZN(new_n10192_));
  NOR4_X1    g09174(.A1(new_n10166_), .A2(new_n10192_), .A3(new_n10180_), .A4(new_n10181_), .ZN(new_n10193_));
  NOR3_X1    g09175(.A1(new_n10191_), .A2(new_n10193_), .A3(new_n10139_), .ZN(new_n10194_));
  OAI21_X1   g09176(.A1(new_n10194_), .A2(new_n10184_), .B(new_n10112_), .ZN(new_n10195_));
  INV_X1     g09177(.I(new_n10112_), .ZN(new_n10196_));
  OAI21_X1   g09178(.A1(new_n10191_), .A2(new_n10193_), .B(new_n10139_), .ZN(new_n10197_));
  NAND3_X1   g09179(.A1(new_n10175_), .A2(new_n10140_), .A3(new_n10183_), .ZN(new_n10198_));
  NAND3_X1   g09180(.A1(new_n10197_), .A2(new_n10198_), .A3(new_n10196_), .ZN(new_n10199_));
  NOR2_X1    g09181(.A1(\A[29] ), .A2(\A[30] ), .ZN(new_n10200_));
  INV_X1     g09182(.I(new_n10200_), .ZN(new_n10201_));
  INV_X1     g09183(.I(\A[29] ), .ZN(new_n10202_));
  INV_X1     g09184(.I(\A[30] ), .ZN(new_n10203_));
  NOR2_X1    g09185(.A1(new_n10202_), .A2(new_n10203_), .ZN(new_n10204_));
  OAI21_X1   g09186(.A1(\A[28] ), .A2(new_n10204_), .B(new_n10201_), .ZN(new_n10205_));
  INV_X1     g09187(.I(new_n10205_), .ZN(new_n10206_));
  NOR2_X1    g09188(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n10207_));
  INV_X1     g09189(.I(new_n10207_), .ZN(new_n10208_));
  INV_X1     g09190(.I(\A[26] ), .ZN(new_n10209_));
  INV_X1     g09191(.I(\A[27] ), .ZN(new_n10210_));
  NOR2_X1    g09192(.A1(new_n10209_), .A2(new_n10210_), .ZN(new_n10211_));
  OAI21_X1   g09193(.A1(\A[25] ), .A2(new_n10211_), .B(new_n10208_), .ZN(new_n10212_));
  INV_X1     g09194(.I(new_n10212_), .ZN(new_n10213_));
  NAND2_X1   g09195(.A1(new_n10206_), .A2(new_n10213_), .ZN(new_n10214_));
  NAND2_X1   g09196(.A1(new_n10205_), .A2(new_n10212_), .ZN(new_n10215_));
  NOR2_X1    g09197(.A1(new_n10210_), .A2(\A[26] ), .ZN(new_n10216_));
  NOR2_X1    g09198(.A1(new_n10209_), .A2(\A[27] ), .ZN(new_n10217_));
  OAI21_X1   g09199(.A1(new_n10216_), .A2(new_n10217_), .B(\A[25] ), .ZN(new_n10218_));
  INV_X1     g09200(.I(\A[25] ), .ZN(new_n10219_));
  OAI21_X1   g09201(.A1(new_n10211_), .A2(new_n10207_), .B(new_n10219_), .ZN(new_n10220_));
  NAND2_X1   g09202(.A1(new_n10220_), .A2(new_n10218_), .ZN(new_n10221_));
  INV_X1     g09203(.I(new_n10221_), .ZN(new_n10222_));
  NOR2_X1    g09204(.A1(new_n10203_), .A2(\A[29] ), .ZN(new_n10223_));
  NOR2_X1    g09205(.A1(new_n10202_), .A2(\A[30] ), .ZN(new_n10224_));
  OAI21_X1   g09206(.A1(new_n10223_), .A2(new_n10224_), .B(\A[28] ), .ZN(new_n10225_));
  INV_X1     g09207(.I(\A[28] ), .ZN(new_n10226_));
  OAI21_X1   g09208(.A1(new_n10204_), .A2(new_n10200_), .B(new_n10226_), .ZN(new_n10227_));
  NAND2_X1   g09209(.A1(new_n10227_), .A2(new_n10225_), .ZN(new_n10228_));
  INV_X1     g09210(.I(new_n10228_), .ZN(new_n10229_));
  NAND3_X1   g09211(.A1(new_n10222_), .A2(new_n10229_), .A3(new_n10215_), .ZN(new_n10230_));
  NAND2_X1   g09212(.A1(new_n10230_), .A2(new_n10214_), .ZN(new_n10231_));
  NOR2_X1    g09213(.A1(\A[23] ), .A2(\A[24] ), .ZN(new_n10232_));
  INV_X1     g09214(.I(\A[23] ), .ZN(new_n10233_));
  INV_X1     g09215(.I(\A[24] ), .ZN(new_n10234_));
  NOR2_X1    g09216(.A1(new_n10233_), .A2(new_n10234_), .ZN(new_n10235_));
  NOR2_X1    g09217(.A1(new_n10235_), .A2(\A[22] ), .ZN(new_n10236_));
  NOR2_X1    g09218(.A1(new_n10236_), .A2(new_n10232_), .ZN(new_n10237_));
  NOR2_X1    g09219(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n10238_));
  INV_X1     g09220(.I(\A[20] ), .ZN(new_n10239_));
  INV_X1     g09221(.I(\A[21] ), .ZN(new_n10240_));
  NOR2_X1    g09222(.A1(new_n10239_), .A2(new_n10240_), .ZN(new_n10241_));
  NOR2_X1    g09223(.A1(new_n10241_), .A2(\A[19] ), .ZN(new_n10242_));
  NOR2_X1    g09224(.A1(new_n10242_), .A2(new_n10238_), .ZN(new_n10243_));
  NAND2_X1   g09225(.A1(new_n10243_), .A2(new_n10237_), .ZN(new_n10244_));
  NOR2_X1    g09226(.A1(new_n10240_), .A2(\A[20] ), .ZN(new_n10245_));
  NOR2_X1    g09227(.A1(new_n10239_), .A2(\A[21] ), .ZN(new_n10246_));
  OAI21_X1   g09228(.A1(new_n10245_), .A2(new_n10246_), .B(\A[19] ), .ZN(new_n10247_));
  INV_X1     g09229(.I(\A[19] ), .ZN(new_n10248_));
  OAI21_X1   g09230(.A1(new_n10241_), .A2(new_n10238_), .B(new_n10248_), .ZN(new_n10249_));
  NAND2_X1   g09231(.A1(new_n10249_), .A2(new_n10247_), .ZN(new_n10250_));
  NOR2_X1    g09232(.A1(new_n10234_), .A2(\A[23] ), .ZN(new_n10251_));
  NOR2_X1    g09233(.A1(new_n10233_), .A2(\A[24] ), .ZN(new_n10252_));
  OAI21_X1   g09234(.A1(new_n10251_), .A2(new_n10252_), .B(\A[22] ), .ZN(new_n10253_));
  INV_X1     g09235(.I(\A[22] ), .ZN(new_n10254_));
  OAI21_X1   g09236(.A1(new_n10235_), .A2(new_n10232_), .B(new_n10254_), .ZN(new_n10255_));
  NAND2_X1   g09237(.A1(new_n10255_), .A2(new_n10253_), .ZN(new_n10256_));
  NOR2_X1    g09238(.A1(new_n10250_), .A2(new_n10256_), .ZN(new_n10257_));
  OAI21_X1   g09239(.A1(new_n10237_), .A2(new_n10243_), .B(new_n10257_), .ZN(new_n10258_));
  NAND2_X1   g09240(.A1(new_n10258_), .A2(new_n10244_), .ZN(new_n10259_));
  INV_X1     g09241(.I(new_n10259_), .ZN(new_n10260_));
  OAI21_X1   g09242(.A1(new_n10250_), .A2(new_n10256_), .B(new_n10243_), .ZN(new_n10261_));
  INV_X1     g09243(.I(new_n10261_), .ZN(new_n10262_));
  NOR3_X1    g09244(.A1(new_n10250_), .A2(new_n10256_), .A3(new_n10243_), .ZN(new_n10263_));
  OAI21_X1   g09245(.A1(new_n10262_), .A2(new_n10263_), .B(new_n10237_), .ZN(new_n10264_));
  INV_X1     g09246(.I(new_n10237_), .ZN(new_n10265_));
  INV_X1     g09247(.I(new_n10263_), .ZN(new_n10266_));
  NAND3_X1   g09248(.A1(new_n10266_), .A2(new_n10265_), .A3(new_n10261_), .ZN(new_n10267_));
  NAND2_X1   g09249(.A1(new_n10264_), .A2(new_n10267_), .ZN(new_n10268_));
  OAI21_X1   g09250(.A1(new_n10221_), .A2(new_n10228_), .B(new_n10213_), .ZN(new_n10269_));
  INV_X1     g09251(.I(new_n10269_), .ZN(new_n10270_));
  NOR3_X1    g09252(.A1(new_n10221_), .A2(new_n10228_), .A3(new_n10213_), .ZN(new_n10271_));
  OAI21_X1   g09253(.A1(new_n10270_), .A2(new_n10271_), .B(new_n10206_), .ZN(new_n10272_));
  NAND3_X1   g09254(.A1(new_n10222_), .A2(new_n10229_), .A3(new_n10212_), .ZN(new_n10273_));
  NAND3_X1   g09255(.A1(new_n10273_), .A2(new_n10205_), .A3(new_n10269_), .ZN(new_n10274_));
  NAND2_X1   g09256(.A1(new_n10272_), .A2(new_n10274_), .ZN(new_n10275_));
  XNOR2_X1   g09257(.A1(new_n10250_), .A2(new_n10256_), .ZN(new_n10276_));
  XNOR2_X1   g09258(.A1(new_n10221_), .A2(new_n10228_), .ZN(new_n10277_));
  NOR3_X1    g09259(.A1(new_n10221_), .A2(new_n10205_), .A3(new_n10212_), .ZN(new_n10278_));
  NAND2_X1   g09260(.A1(new_n10278_), .A2(new_n10229_), .ZN(new_n10279_));
  NAND3_X1   g09261(.A1(new_n10257_), .A2(new_n10237_), .A3(new_n10243_), .ZN(new_n10280_));
  NOR4_X1    g09262(.A1(new_n10276_), .A2(new_n10277_), .A3(new_n10279_), .A4(new_n10280_), .ZN(new_n10281_));
  OAI21_X1   g09263(.A1(new_n10275_), .A2(new_n10281_), .B(new_n10268_), .ZN(new_n10282_));
  AOI21_X1   g09264(.A1(new_n10273_), .A2(new_n10269_), .B(new_n10205_), .ZN(new_n10283_));
  NOR3_X1    g09265(.A1(new_n10270_), .A2(new_n10206_), .A3(new_n10271_), .ZN(new_n10284_));
  NOR2_X1    g09266(.A1(new_n10284_), .A2(new_n10283_), .ZN(new_n10285_));
  XOR2_X1    g09267(.A1(new_n10250_), .A2(new_n10256_), .Z(new_n10286_));
  XOR2_X1    g09268(.A1(new_n10221_), .A2(new_n10228_), .Z(new_n10287_));
  AOI21_X1   g09269(.A1(new_n10221_), .A2(new_n10228_), .B(new_n10214_), .ZN(new_n10288_));
  NOR2_X1    g09270(.A1(new_n10288_), .A2(new_n10280_), .ZN(new_n10289_));
  NAND4_X1   g09271(.A1(new_n10285_), .A2(new_n10286_), .A3(new_n10287_), .A4(new_n10289_), .ZN(new_n10290_));
  AOI21_X1   g09272(.A1(new_n10282_), .A2(new_n10290_), .B(new_n10260_), .ZN(new_n10291_));
  AOI21_X1   g09273(.A1(new_n10266_), .A2(new_n10261_), .B(new_n10265_), .ZN(new_n10292_));
  NOR3_X1    g09274(.A1(new_n10262_), .A2(new_n10237_), .A3(new_n10263_), .ZN(new_n10293_));
  NOR2_X1    g09275(.A1(new_n10293_), .A2(new_n10292_), .ZN(new_n10294_));
  NOR2_X1    g09276(.A1(new_n10280_), .A2(new_n10279_), .ZN(new_n10295_));
  NAND3_X1   g09277(.A1(new_n10295_), .A2(new_n10286_), .A3(new_n10287_), .ZN(new_n10296_));
  AOI21_X1   g09278(.A1(new_n10285_), .A2(new_n10296_), .B(new_n10294_), .ZN(new_n10297_));
  NAND2_X1   g09279(.A1(new_n10286_), .A2(new_n10287_), .ZN(new_n10298_));
  NOR4_X1    g09280(.A1(new_n10275_), .A2(new_n10298_), .A3(new_n10280_), .A4(new_n10288_), .ZN(new_n10299_));
  NOR3_X1    g09281(.A1(new_n10297_), .A2(new_n10299_), .A3(new_n10259_), .ZN(new_n10300_));
  OAI21_X1   g09282(.A1(new_n10300_), .A2(new_n10291_), .B(new_n10231_), .ZN(new_n10301_));
  INV_X1     g09283(.I(new_n10231_), .ZN(new_n10302_));
  OAI21_X1   g09284(.A1(new_n10297_), .A2(new_n10299_), .B(new_n10259_), .ZN(new_n10303_));
  NAND3_X1   g09285(.A1(new_n10282_), .A2(new_n10290_), .A3(new_n10260_), .ZN(new_n10304_));
  NAND3_X1   g09286(.A1(new_n10303_), .A2(new_n10304_), .A3(new_n10302_), .ZN(new_n10305_));
  AOI22_X1   g09287(.A1(new_n10301_), .A2(new_n10305_), .B1(new_n10195_), .B2(new_n10199_), .ZN(new_n10306_));
  NAND2_X1   g09288(.A1(new_n10195_), .A2(new_n10199_), .ZN(new_n10307_));
  NAND2_X1   g09289(.A1(new_n10301_), .A2(new_n10305_), .ZN(new_n10308_));
  NOR2_X1    g09290(.A1(new_n10308_), .A2(new_n10307_), .ZN(new_n10309_));
  AOI21_X1   g09291(.A1(new_n10285_), .A2(new_n10296_), .B(new_n10268_), .ZN(new_n10311_));
  NAND4_X1   g09292(.A1(new_n10206_), .A2(\A[25] ), .A3(\A[26] ), .A4(\A[27] ), .ZN(new_n10312_));
  NOR3_X1    g09293(.A1(new_n10312_), .A2(new_n10222_), .A3(new_n10228_), .ZN(new_n10313_));
  NOR3_X1    g09294(.A1(new_n10276_), .A2(new_n10280_), .A3(new_n10313_), .ZN(new_n10314_));
  NOR3_X1    g09295(.A1(new_n10244_), .A2(new_n10250_), .A3(new_n10256_), .ZN(new_n10315_));
  NAND3_X1   g09296(.A1(new_n10278_), .A2(new_n10221_), .A3(new_n10229_), .ZN(new_n10316_));
  AOI21_X1   g09297(.A1(new_n10286_), .A2(new_n10315_), .B(new_n10316_), .ZN(new_n10317_));
  NOR3_X1    g09298(.A1(new_n10102_), .A2(new_n10160_), .A3(new_n10170_), .ZN(new_n10318_));
  NOR3_X1    g09299(.A1(new_n10168_), .A2(new_n10180_), .A3(new_n10318_), .ZN(new_n10319_));
  OR3_X2     g09300(.A1(new_n10102_), .A2(new_n10160_), .A3(new_n10170_), .Z(new_n10320_));
  AOI21_X1   g09301(.A1(new_n10188_), .A2(new_n10172_), .B(new_n10320_), .ZN(new_n10321_));
  OAI22_X1   g09302(.A1(new_n10319_), .A2(new_n10321_), .B1(new_n10314_), .B2(new_n10317_), .ZN(new_n10322_));
  NAND2_X1   g09303(.A1(new_n10311_), .A2(new_n10322_), .ZN(new_n10323_));
  OAI21_X1   g09304(.A1(new_n10275_), .A2(new_n10281_), .B(new_n10294_), .ZN(new_n10324_));
  NAND3_X1   g09305(.A1(new_n10286_), .A2(new_n10315_), .A3(new_n10316_), .ZN(new_n10325_));
  OAI21_X1   g09306(.A1(new_n10276_), .A2(new_n10280_), .B(new_n10313_), .ZN(new_n10326_));
  NAND3_X1   g09307(.A1(new_n10188_), .A2(new_n10320_), .A3(new_n10172_), .ZN(new_n10327_));
  OAI21_X1   g09308(.A1(new_n10168_), .A2(new_n10180_), .B(new_n10318_), .ZN(new_n10328_));
  AOI22_X1   g09309(.A1(new_n10327_), .A2(new_n10328_), .B1(new_n10326_), .B2(new_n10325_), .ZN(new_n10329_));
  NAND2_X1   g09310(.A1(new_n10324_), .A2(new_n10329_), .ZN(new_n10330_));
  NAND2_X1   g09311(.A1(new_n10330_), .A2(new_n10323_), .ZN(new_n10331_));
  NOR2_X1    g09312(.A1(new_n10311_), .A2(new_n10322_), .ZN(new_n10332_));
  NOR2_X1    g09313(.A1(new_n10183_), .A2(new_n10187_), .ZN(new_n10333_));
  NAND2_X1   g09314(.A1(new_n10152_), .A2(new_n10174_), .ZN(new_n10334_));
  OAI21_X1   g09315(.A1(new_n10152_), .A2(new_n10174_), .B(new_n10178_), .ZN(new_n10335_));
  NAND3_X1   g09316(.A1(new_n10187_), .A2(new_n10190_), .A3(new_n10166_), .ZN(new_n10336_));
  NAND2_X1   g09317(.A1(new_n10335_), .A2(new_n10336_), .ZN(new_n10337_));
  AOI21_X1   g09318(.A1(new_n10337_), .A2(new_n10334_), .B(new_n10333_), .ZN(new_n10338_));
  AOI21_X1   g09319(.A1(new_n10331_), .A2(new_n10338_), .B(new_n10332_), .ZN(new_n10339_));
  NOR3_X1    g09320(.A1(new_n10309_), .A2(new_n10306_), .A3(new_n10339_), .ZN(new_n10340_));
  NAND2_X1   g09321(.A1(new_n10308_), .A2(new_n10307_), .ZN(new_n10341_));
  NAND4_X1   g09322(.A1(new_n10301_), .A2(new_n10305_), .A3(new_n10195_), .A4(new_n10199_), .ZN(new_n10342_));
  NAND2_X1   g09323(.A1(new_n10193_), .A2(new_n10152_), .ZN(new_n10343_));
  AOI21_X1   g09324(.A1(new_n10187_), .A2(new_n10190_), .B(new_n10166_), .ZN(new_n10344_));
  NOR3_X1    g09325(.A1(new_n10152_), .A2(new_n10174_), .A3(new_n10178_), .ZN(new_n10345_));
  OAI21_X1   g09326(.A1(new_n10345_), .A2(new_n10344_), .B(new_n10334_), .ZN(new_n10346_));
  NAND2_X1   g09327(.A1(new_n10346_), .A2(new_n10343_), .ZN(new_n10347_));
  AOI22_X1   g09328(.A1(new_n10347_), .A2(new_n10311_), .B1(new_n10323_), .B2(new_n10330_), .ZN(new_n10348_));
  AOI21_X1   g09329(.A1(new_n10341_), .A2(new_n10342_), .B(new_n10348_), .ZN(new_n10349_));
  NOR2_X1    g09330(.A1(\A[995] ), .A2(\A[996] ), .ZN(new_n10350_));
  INV_X1     g09331(.I(\A[995] ), .ZN(new_n10351_));
  INV_X1     g09332(.I(\A[996] ), .ZN(new_n10352_));
  NOR2_X1    g09333(.A1(new_n10351_), .A2(new_n10352_), .ZN(new_n10353_));
  NOR2_X1    g09334(.A1(new_n10353_), .A2(\A[994] ), .ZN(new_n10354_));
  NOR2_X1    g09335(.A1(new_n10354_), .A2(new_n10350_), .ZN(new_n10355_));
  INV_X1     g09336(.I(new_n10355_), .ZN(new_n10356_));
  NOR2_X1    g09337(.A1(\A[992] ), .A2(\A[993] ), .ZN(new_n10357_));
  INV_X1     g09338(.I(new_n10357_), .ZN(new_n10358_));
  INV_X1     g09339(.I(\A[992] ), .ZN(new_n10359_));
  INV_X1     g09340(.I(\A[993] ), .ZN(new_n10360_));
  NOR2_X1    g09341(.A1(new_n10359_), .A2(new_n10360_), .ZN(new_n10361_));
  OAI21_X1   g09342(.A1(\A[991] ), .A2(new_n10361_), .B(new_n10358_), .ZN(new_n10362_));
  NOR2_X1    g09343(.A1(new_n10356_), .A2(new_n10362_), .ZN(new_n10363_));
  INV_X1     g09344(.I(new_n10363_), .ZN(new_n10364_));
  INV_X1     g09345(.I(new_n10362_), .ZN(new_n10365_));
  NOR2_X1    g09346(.A1(new_n10365_), .A2(new_n10355_), .ZN(new_n10366_));
  NOR2_X1    g09347(.A1(new_n10360_), .A2(\A[992] ), .ZN(new_n10367_));
  NOR2_X1    g09348(.A1(new_n10359_), .A2(\A[993] ), .ZN(new_n10368_));
  OAI21_X1   g09349(.A1(new_n10367_), .A2(new_n10368_), .B(\A[991] ), .ZN(new_n10369_));
  NOR2_X1    g09350(.A1(new_n10361_), .A2(new_n10357_), .ZN(new_n10370_));
  OAI21_X1   g09351(.A1(\A[991] ), .A2(new_n10370_), .B(new_n10369_), .ZN(new_n10371_));
  NOR2_X1    g09352(.A1(new_n10352_), .A2(\A[995] ), .ZN(new_n10372_));
  NOR2_X1    g09353(.A1(new_n10351_), .A2(\A[996] ), .ZN(new_n10373_));
  OAI21_X1   g09354(.A1(new_n10372_), .A2(new_n10373_), .B(\A[994] ), .ZN(new_n10374_));
  NOR2_X1    g09355(.A1(new_n10353_), .A2(new_n10350_), .ZN(new_n10375_));
  OAI21_X1   g09356(.A1(\A[994] ), .A2(new_n10375_), .B(new_n10374_), .ZN(new_n10376_));
  NOR2_X1    g09357(.A1(new_n10371_), .A2(new_n10376_), .ZN(new_n10377_));
  INV_X1     g09358(.I(new_n10377_), .ZN(new_n10378_));
  OAI21_X1   g09359(.A1(new_n10378_), .A2(new_n10366_), .B(new_n10364_), .ZN(new_n10379_));
  INV_X1     g09360(.I(new_n10379_), .ZN(new_n10380_));
  NOR2_X1    g09361(.A1(\A[1] ), .A2(\A[2] ), .ZN(new_n10381_));
  AOI21_X1   g09362(.A1(\A[1] ), .A2(\A[2] ), .B(\A[0] ), .ZN(new_n10382_));
  NOR2_X1    g09363(.A1(new_n10382_), .A2(new_n10381_), .ZN(new_n10383_));
  INV_X1     g09364(.I(\A[3] ), .ZN(new_n10384_));
  NOR2_X1    g09365(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n10385_));
  NAND2_X1   g09366(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n10386_));
  AOI21_X1   g09367(.A1(new_n10384_), .A2(new_n10386_), .B(new_n10385_), .ZN(new_n10387_));
  INV_X1     g09368(.I(new_n10387_), .ZN(new_n10388_));
  XOR2_X1    g09369(.A1(\A[4] ), .A2(\A[5] ), .Z(new_n10389_));
  INV_X1     g09370(.I(new_n10385_), .ZN(new_n10390_));
  AOI21_X1   g09371(.A1(new_n10390_), .A2(new_n10386_), .B(\A[3] ), .ZN(new_n10391_));
  AOI21_X1   g09372(.A1(\A[3] ), .A2(new_n10389_), .B(new_n10391_), .ZN(new_n10392_));
  INV_X1     g09373(.I(\A[2] ), .ZN(new_n10393_));
  XOR2_X1    g09374(.A1(\A[0] ), .A2(\A[1] ), .Z(new_n10394_));
  NAND2_X1   g09375(.A1(new_n10394_), .A2(new_n10393_), .ZN(new_n10395_));
  XNOR2_X1   g09376(.A1(\A[0] ), .A2(\A[1] ), .ZN(new_n10396_));
  NAND2_X1   g09377(.A1(new_n10396_), .A2(\A[2] ), .ZN(new_n10397_));
  AOI21_X1   g09378(.A1(new_n10397_), .A2(new_n10395_), .B(\A[6] ), .ZN(new_n10398_));
  INV_X1     g09379(.I(\A[0] ), .ZN(new_n10399_));
  XOR2_X1    g09380(.A1(\A[1] ), .A2(\A[2] ), .Z(new_n10400_));
  NAND2_X1   g09381(.A1(new_n10400_), .A2(new_n10399_), .ZN(new_n10401_));
  XNOR2_X1   g09382(.A1(\A[1] ), .A2(\A[2] ), .ZN(new_n10402_));
  NAND2_X1   g09383(.A1(new_n10402_), .A2(\A[0] ), .ZN(new_n10403_));
  AOI21_X1   g09384(.A1(new_n10403_), .A2(new_n10401_), .B(\A[6] ), .ZN(new_n10404_));
  OAI21_X1   g09385(.A1(new_n10398_), .A2(new_n10404_), .B(new_n10392_), .ZN(new_n10405_));
  XNOR2_X1   g09386(.A1(new_n10387_), .A2(new_n10383_), .ZN(new_n10406_));
  INV_X1     g09387(.I(\A[6] ), .ZN(new_n10407_));
  AOI21_X1   g09388(.A1(new_n10397_), .A2(new_n10395_), .B(new_n10407_), .ZN(new_n10408_));
  NOR2_X1    g09389(.A1(new_n10406_), .A2(new_n10408_), .ZN(new_n10409_));
  AOI22_X1   g09390(.A1(new_n10405_), .A2(new_n10409_), .B1(new_n10383_), .B2(new_n10388_), .ZN(new_n10410_));
  XOR2_X1    g09391(.A1(new_n10387_), .A2(new_n10383_), .Z(new_n10411_));
  INV_X1     g09392(.I(new_n10408_), .ZN(new_n10412_));
  NAND2_X1   g09393(.A1(new_n10405_), .A2(new_n10412_), .ZN(new_n10413_));
  NAND2_X1   g09394(.A1(new_n10413_), .A2(new_n10411_), .ZN(new_n10414_));
  INV_X1     g09395(.I(new_n10411_), .ZN(new_n10415_));
  NAND3_X1   g09396(.A1(new_n10405_), .A2(new_n10412_), .A3(new_n10415_), .ZN(new_n10416_));
  INV_X1     g09397(.I(new_n10392_), .ZN(new_n10417_));
  INV_X1     g09398(.I(new_n10398_), .ZN(new_n10418_));
  NOR2_X1    g09399(.A1(new_n10402_), .A2(\A[0] ), .ZN(new_n10419_));
  NOR2_X1    g09400(.A1(new_n10400_), .A2(new_n10399_), .ZN(new_n10420_));
  OAI21_X1   g09401(.A1(new_n10419_), .A2(new_n10420_), .B(new_n10407_), .ZN(new_n10421_));
  NAND3_X1   g09402(.A1(new_n10418_), .A2(new_n10417_), .A3(new_n10421_), .ZN(new_n10422_));
  XOR2_X1    g09403(.A1(\A[998] ), .A2(\A[999] ), .Z(new_n10423_));
  NAND2_X1   g09404(.A1(new_n10423_), .A2(\A[997] ), .ZN(new_n10424_));
  INV_X1     g09405(.I(\A[997] ), .ZN(new_n10425_));
  AND2_X2    g09406(.A1(\A[998] ), .A2(\A[999] ), .Z(new_n10426_));
  NOR2_X1    g09407(.A1(\A[998] ), .A2(\A[999] ), .ZN(new_n10427_));
  OAI21_X1   g09408(.A1(new_n10426_), .A2(new_n10427_), .B(new_n10425_), .ZN(new_n10428_));
  NAND2_X1   g09409(.A1(new_n10424_), .A2(new_n10428_), .ZN(new_n10429_));
  INV_X1     g09410(.I(new_n10429_), .ZN(new_n10430_));
  NAND3_X1   g09411(.A1(new_n10422_), .A2(new_n10405_), .A3(new_n10430_), .ZN(new_n10431_));
  AOI21_X1   g09412(.A1(new_n10414_), .A2(new_n10416_), .B(new_n10431_), .ZN(new_n10432_));
  NOR2_X1    g09413(.A1(new_n10426_), .A2(\A[997] ), .ZN(new_n10433_));
  NOR2_X1    g09414(.A1(new_n10433_), .A2(new_n10427_), .ZN(new_n10434_));
  OAI21_X1   g09415(.A1(new_n10432_), .A2(new_n10434_), .B(new_n10410_), .ZN(new_n10435_));
  INV_X1     g09416(.I(new_n10410_), .ZN(new_n10436_));
  AOI21_X1   g09417(.A1(new_n10405_), .A2(new_n10412_), .B(new_n10415_), .ZN(new_n10437_));
  INV_X1     g09418(.I(new_n10416_), .ZN(new_n10438_));
  AOI21_X1   g09419(.A1(new_n10418_), .A2(new_n10421_), .B(new_n10417_), .ZN(new_n10439_));
  NOR3_X1    g09420(.A1(new_n10398_), .A2(new_n10404_), .A3(new_n10392_), .ZN(new_n10440_));
  NOR3_X1    g09421(.A1(new_n10439_), .A2(new_n10440_), .A3(new_n10429_), .ZN(new_n10441_));
  OAI21_X1   g09422(.A1(new_n10438_), .A2(new_n10437_), .B(new_n10441_), .ZN(new_n10442_));
  INV_X1     g09423(.I(new_n10434_), .ZN(new_n10443_));
  NAND3_X1   g09424(.A1(new_n10442_), .A2(new_n10436_), .A3(new_n10443_), .ZN(new_n10444_));
  NAND2_X1   g09425(.A1(new_n10444_), .A2(new_n10435_), .ZN(new_n10445_));
  NAND2_X1   g09426(.A1(new_n10445_), .A2(new_n10380_), .ZN(new_n10446_));
  NOR3_X1    g09427(.A1(new_n10432_), .A2(new_n10436_), .A3(new_n10434_), .ZN(new_n10447_));
  INV_X1     g09428(.I(new_n10447_), .ZN(new_n10448_));
  OAI21_X1   g09429(.A1(new_n10432_), .A2(new_n10434_), .B(new_n10436_), .ZN(new_n10449_));
  NAND3_X1   g09430(.A1(new_n10448_), .A2(new_n10449_), .A3(new_n10379_), .ZN(new_n10450_));
  NAND2_X1   g09431(.A1(new_n10446_), .A2(new_n10450_), .ZN(new_n10451_));
  AOI21_X1   g09432(.A1(new_n10418_), .A2(new_n10421_), .B(new_n10429_), .ZN(new_n10452_));
  NOR3_X1    g09433(.A1(new_n10430_), .A2(new_n10398_), .A3(new_n10404_), .ZN(new_n10453_));
  OAI21_X1   g09434(.A1(new_n10452_), .A2(new_n10453_), .B(new_n10392_), .ZN(new_n10454_));
  NOR3_X1    g09435(.A1(new_n10452_), .A2(new_n10392_), .A3(new_n10453_), .ZN(new_n10455_));
  INV_X1     g09436(.I(new_n10455_), .ZN(new_n10456_));
  XNOR2_X1   g09437(.A1(new_n10371_), .A2(new_n10376_), .ZN(new_n10457_));
  INV_X1     g09438(.I(new_n10457_), .ZN(new_n10458_));
  NAND3_X1   g09439(.A1(new_n10456_), .A2(new_n10454_), .A3(new_n10458_), .ZN(new_n10459_));
  NAND2_X1   g09440(.A1(new_n10442_), .A2(new_n10443_), .ZN(new_n10460_));
  NAND2_X1   g09441(.A1(new_n10432_), .A2(new_n10434_), .ZN(new_n10461_));
  AOI21_X1   g09442(.A1(new_n10460_), .A2(new_n10461_), .B(new_n10459_), .ZN(new_n10462_));
  INV_X1     g09443(.I(new_n10454_), .ZN(new_n10463_));
  NOR3_X1    g09444(.A1(new_n10463_), .A2(new_n10455_), .A3(new_n10457_), .ZN(new_n10464_));
  NAND2_X1   g09445(.A1(new_n10414_), .A2(new_n10416_), .ZN(new_n10465_));
  AOI21_X1   g09446(.A1(new_n10465_), .A2(new_n10441_), .B(new_n10434_), .ZN(new_n10466_));
  NOR2_X1    g09447(.A1(new_n10442_), .A2(new_n10443_), .ZN(new_n10467_));
  NOR2_X1    g09448(.A1(new_n10377_), .A2(new_n10362_), .ZN(new_n10468_));
  NAND2_X1   g09449(.A1(new_n10377_), .A2(new_n10362_), .ZN(new_n10469_));
  INV_X1     g09450(.I(new_n10469_), .ZN(new_n10470_));
  OAI21_X1   g09451(.A1(new_n10470_), .A2(new_n10468_), .B(new_n10355_), .ZN(new_n10471_));
  INV_X1     g09452(.I(new_n10468_), .ZN(new_n10472_));
  NAND3_X1   g09453(.A1(new_n10472_), .A2(new_n10356_), .A3(new_n10469_), .ZN(new_n10473_));
  AND2_X2    g09454(.A1(new_n10471_), .A2(new_n10473_), .Z(new_n10474_));
  NOR4_X1    g09455(.A1(new_n10467_), .A2(new_n10474_), .A3(new_n10466_), .A4(new_n10464_), .ZN(new_n10475_));
  NOR2_X1    g09456(.A1(new_n10475_), .A2(new_n10462_), .ZN(new_n10476_));
  NOR2_X1    g09457(.A1(new_n10451_), .A2(new_n10476_), .ZN(new_n10477_));
  AOI21_X1   g09458(.A1(new_n10444_), .A2(new_n10435_), .B(new_n10379_), .ZN(new_n10478_));
  AOI21_X1   g09459(.A1(new_n10442_), .A2(new_n10443_), .B(new_n10410_), .ZN(new_n10479_));
  NOR2_X1    g09460(.A1(new_n10479_), .A2(new_n10447_), .ZN(new_n10480_));
  AOI21_X1   g09461(.A1(new_n10379_), .A2(new_n10480_), .B(new_n10478_), .ZN(new_n10481_));
  OAI21_X1   g09462(.A1(new_n10467_), .A2(new_n10466_), .B(new_n10464_), .ZN(new_n10482_));
  NAND2_X1   g09463(.A1(new_n10471_), .A2(new_n10473_), .ZN(new_n10483_));
  NAND4_X1   g09464(.A1(new_n10460_), .A2(new_n10461_), .A3(new_n10459_), .A4(new_n10483_), .ZN(new_n10484_));
  NAND2_X1   g09465(.A1(new_n10484_), .A2(new_n10482_), .ZN(new_n10485_));
  NOR2_X1    g09466(.A1(new_n10481_), .A2(new_n10485_), .ZN(new_n10486_));
  NOR2_X1    g09467(.A1(new_n10477_), .A2(new_n10486_), .ZN(new_n10487_));
  OAI21_X1   g09468(.A1(new_n10340_), .A2(new_n10349_), .B(new_n10487_), .ZN(new_n10488_));
  NAND3_X1   g09469(.A1(new_n10341_), .A2(new_n10342_), .A3(new_n10348_), .ZN(new_n10489_));
  OAI21_X1   g09470(.A1(new_n10309_), .A2(new_n10306_), .B(new_n10339_), .ZN(new_n10490_));
  NAND2_X1   g09471(.A1(new_n10481_), .A2(new_n10485_), .ZN(new_n10491_));
  NAND2_X1   g09472(.A1(new_n10451_), .A2(new_n10476_), .ZN(new_n10492_));
  NAND2_X1   g09473(.A1(new_n10492_), .A2(new_n10491_), .ZN(new_n10493_));
  NAND3_X1   g09474(.A1(new_n10490_), .A2(new_n10489_), .A3(new_n10493_), .ZN(new_n10494_));
  NAND3_X1   g09475(.A1(new_n10490_), .A2(new_n10489_), .A3(new_n10493_), .ZN(new_n10495_));
  NAND3_X1   g09476(.A1(new_n10488_), .A2(new_n10494_), .A3(new_n10495_), .ZN(new_n10496_));
  NAND2_X1   g09477(.A1(new_n10485_), .A2(new_n10480_), .ZN(new_n10497_));
  INV_X1     g09478(.I(new_n10480_), .ZN(new_n10498_));
  NOR2_X1    g09479(.A1(new_n10476_), .A2(new_n10498_), .ZN(new_n10499_));
  NAND2_X1   g09480(.A1(new_n10499_), .A2(new_n10379_), .ZN(new_n10500_));
  NAND3_X1   g09481(.A1(new_n10500_), .A2(new_n10435_), .A3(new_n10497_), .ZN(new_n10501_));
  INV_X1     g09482(.I(new_n10435_), .ZN(new_n10502_));
  NOR2_X1    g09483(.A1(new_n10497_), .A2(new_n10380_), .ZN(new_n10503_));
  OAI21_X1   g09484(.A1(new_n10503_), .A2(new_n10499_), .B(new_n10502_), .ZN(new_n10504_));
  NAND2_X1   g09485(.A1(new_n10501_), .A2(new_n10504_), .ZN(new_n10505_));
  NOR2_X1    g09486(.A1(new_n10260_), .A2(new_n10302_), .ZN(new_n10506_));
  NAND2_X1   g09487(.A1(new_n10282_), .A2(new_n10290_), .ZN(new_n10507_));
  AOI21_X1   g09488(.A1(new_n10302_), .A2(new_n10260_), .B(new_n10507_), .ZN(new_n10508_));
  NOR2_X1    g09489(.A1(new_n10508_), .A2(new_n10506_), .ZN(new_n10509_));
  INV_X1     g09490(.I(new_n10509_), .ZN(new_n10510_));
  NOR2_X1    g09491(.A1(new_n10140_), .A2(new_n10196_), .ZN(new_n10511_));
  NAND2_X1   g09492(.A1(new_n10175_), .A2(new_n10183_), .ZN(new_n10512_));
  AOI21_X1   g09493(.A1(new_n10196_), .A2(new_n10140_), .B(new_n10512_), .ZN(new_n10513_));
  NOR2_X1    g09494(.A1(new_n10513_), .A2(new_n10511_), .ZN(new_n10514_));
  OAI21_X1   g09495(.A1(new_n10308_), .A2(new_n10307_), .B(new_n10339_), .ZN(new_n10515_));
  XOR2_X1    g09496(.A1(new_n10259_), .A2(new_n10231_), .Z(new_n10516_));
  XOR2_X1    g09497(.A1(new_n10139_), .A2(new_n10112_), .Z(new_n10517_));
  NOR4_X1    g09498(.A1(new_n10507_), .A2(new_n10512_), .A3(new_n10516_), .A4(new_n10517_), .ZN(new_n10518_));
  AOI21_X1   g09499(.A1(new_n10515_), .A2(new_n10518_), .B(new_n10514_), .ZN(new_n10519_));
  INV_X1     g09500(.I(new_n10514_), .ZN(new_n10520_));
  AOI21_X1   g09501(.A1(new_n10197_), .A2(new_n10198_), .B(new_n10196_), .ZN(new_n10521_));
  NOR3_X1    g09502(.A1(new_n10194_), .A2(new_n10184_), .A3(new_n10112_), .ZN(new_n10522_));
  NOR2_X1    g09503(.A1(new_n10522_), .A2(new_n10521_), .ZN(new_n10523_));
  AOI21_X1   g09504(.A1(new_n10303_), .A2(new_n10304_), .B(new_n10302_), .ZN(new_n10524_));
  NOR3_X1    g09505(.A1(new_n10300_), .A2(new_n10291_), .A3(new_n10231_), .ZN(new_n10525_));
  NOR2_X1    g09506(.A1(new_n10525_), .A2(new_n10524_), .ZN(new_n10526_));
  AOI21_X1   g09507(.A1(new_n10526_), .A2(new_n10523_), .B(new_n10348_), .ZN(new_n10527_));
  INV_X1     g09508(.I(new_n10518_), .ZN(new_n10528_));
  NOR3_X1    g09509(.A1(new_n10527_), .A2(new_n10520_), .A3(new_n10528_), .ZN(new_n10529_));
  OAI21_X1   g09510(.A1(new_n10529_), .A2(new_n10519_), .B(new_n10510_), .ZN(new_n10530_));
  OAI21_X1   g09511(.A1(new_n10527_), .A2(new_n10528_), .B(new_n10520_), .ZN(new_n10531_));
  NAND3_X1   g09512(.A1(new_n10515_), .A2(new_n10514_), .A3(new_n10518_), .ZN(new_n10532_));
  NAND3_X1   g09513(.A1(new_n10531_), .A2(new_n10532_), .A3(new_n10509_), .ZN(new_n10533_));
  AOI21_X1   g09514(.A1(new_n10530_), .A2(new_n10533_), .B(new_n10505_), .ZN(new_n10534_));
  NOR3_X1    g09515(.A1(new_n10503_), .A2(new_n10502_), .A3(new_n10499_), .ZN(new_n10535_));
  AOI21_X1   g09516(.A1(new_n10500_), .A2(new_n10497_), .B(new_n10435_), .ZN(new_n10536_));
  NOR2_X1    g09517(.A1(new_n10536_), .A2(new_n10535_), .ZN(new_n10537_));
  AOI21_X1   g09518(.A1(new_n10531_), .A2(new_n10532_), .B(new_n10509_), .ZN(new_n10538_));
  NOR3_X1    g09519(.A1(new_n10529_), .A2(new_n10519_), .A3(new_n10510_), .ZN(new_n10539_));
  NOR3_X1    g09520(.A1(new_n10539_), .A2(new_n10538_), .A3(new_n10537_), .ZN(new_n10540_));
  OAI21_X1   g09521(.A1(new_n10540_), .A2(new_n10534_), .B(new_n10496_), .ZN(new_n10541_));
  AOI21_X1   g09522(.A1(new_n10490_), .A2(new_n10489_), .B(new_n10493_), .ZN(new_n10542_));
  NOR3_X1    g09523(.A1(new_n10340_), .A2(new_n10349_), .A3(new_n10487_), .ZN(new_n10543_));
  NOR3_X1    g09524(.A1(new_n10340_), .A2(new_n10349_), .A3(new_n10487_), .ZN(new_n10544_));
  NOR3_X1    g09525(.A1(new_n10543_), .A2(new_n10544_), .A3(new_n10542_), .ZN(new_n10545_));
  NOR3_X1    g09526(.A1(new_n10539_), .A2(new_n10538_), .A3(new_n10505_), .ZN(new_n10546_));
  AOI21_X1   g09527(.A1(new_n10530_), .A2(new_n10533_), .B(new_n10537_), .ZN(new_n10547_));
  OAI21_X1   g09528(.A1(new_n10546_), .A2(new_n10547_), .B(new_n10545_), .ZN(new_n10548_));
  NAND4_X1   g09529(.A1(new_n10069_), .A2(new_n10082_), .A3(new_n10541_), .A4(new_n10548_), .ZN(new_n10549_));
  NAND2_X1   g09530(.A1(new_n10075_), .A2(new_n10006_), .ZN(new_n10550_));
  NAND3_X1   g09531(.A1(new_n10074_), .A2(new_n9969_), .A3(new_n9980_), .ZN(new_n10551_));
  AOI21_X1   g09532(.A1(new_n10550_), .A2(new_n10551_), .B(new_n10003_), .ZN(new_n10552_));
  AOI21_X1   g09533(.A1(new_n10076_), .A2(new_n9981_), .B(new_n10073_), .ZN(new_n10553_));
  NOR2_X1    g09534(.A1(new_n10309_), .A2(new_n10306_), .ZN(new_n10554_));
  AOI21_X1   g09535(.A1(new_n10492_), .A2(new_n10491_), .B(new_n10348_), .ZN(new_n10555_));
  NOR3_X1    g09536(.A1(new_n10477_), .A2(new_n10486_), .A3(new_n10339_), .ZN(new_n10556_));
  OAI21_X1   g09537(.A1(new_n10556_), .A2(new_n10555_), .B(new_n10554_), .ZN(new_n10557_));
  NAND2_X1   g09538(.A1(new_n10341_), .A2(new_n10342_), .ZN(new_n10558_));
  OAI21_X1   g09539(.A1(new_n10477_), .A2(new_n10486_), .B(new_n10339_), .ZN(new_n10559_));
  NAND3_X1   g09540(.A1(new_n10492_), .A2(new_n10491_), .A3(new_n10348_), .ZN(new_n10560_));
  NAND3_X1   g09541(.A1(new_n10559_), .A2(new_n10560_), .A3(new_n10558_), .ZN(new_n10561_));
  NAND2_X1   g09542(.A1(new_n10557_), .A2(new_n10561_), .ZN(new_n10562_));
  NOR3_X1    g09543(.A1(new_n10552_), .A2(new_n10553_), .A3(new_n10562_), .ZN(new_n10563_));
  NAND2_X1   g09544(.A1(new_n10071_), .A2(new_n10002_), .ZN(new_n10564_));
  NOR2_X1    g09545(.A1(new_n9988_), .A2(new_n9987_), .ZN(new_n10565_));
  NOR2_X1    g09546(.A1(new_n9992_), .A2(new_n9993_), .ZN(new_n10566_));
  NOR2_X1    g09547(.A1(new_n10566_), .A2(new_n10565_), .ZN(new_n10567_));
  NOR2_X1    g09548(.A1(new_n10567_), .A2(new_n9994_), .ZN(new_n10568_));
  NOR2_X1    g09549(.A1(new_n10276_), .A2(new_n10280_), .ZN(new_n10569_));
  XOR2_X1    g09550(.A1(new_n10569_), .A2(new_n10313_), .Z(new_n10570_));
  OAI21_X1   g09551(.A1(new_n10463_), .A2(new_n10455_), .B(new_n10457_), .ZN(new_n10571_));
  NAND2_X1   g09552(.A1(new_n10571_), .A2(new_n10459_), .ZN(new_n10572_));
  NOR2_X1    g09553(.A1(new_n10168_), .A2(new_n10180_), .ZN(new_n10573_));
  XOR2_X1    g09554(.A1(new_n10573_), .A2(new_n10320_), .Z(new_n10574_));
  NAND2_X1   g09555(.A1(new_n10572_), .A2(new_n10574_), .ZN(new_n10575_));
  XOR2_X1    g09556(.A1(new_n10573_), .A2(new_n10318_), .Z(new_n10576_));
  NAND3_X1   g09557(.A1(new_n10576_), .A2(new_n10571_), .A3(new_n10459_), .ZN(new_n10577_));
  AOI21_X1   g09558(.A1(new_n10575_), .A2(new_n10577_), .B(new_n10570_), .ZN(new_n10578_));
  INV_X1     g09559(.I(new_n10570_), .ZN(new_n10579_));
  NAND2_X1   g09560(.A1(new_n10572_), .A2(new_n10576_), .ZN(new_n10580_));
  NAND3_X1   g09561(.A1(new_n10574_), .A2(new_n10571_), .A3(new_n10459_), .ZN(new_n10581_));
  AOI21_X1   g09562(.A1(new_n10580_), .A2(new_n10581_), .B(new_n10579_), .ZN(new_n10582_));
  NOR2_X1    g09563(.A1(new_n10578_), .A2(new_n10582_), .ZN(new_n10583_));
  NAND2_X1   g09564(.A1(new_n10568_), .A2(new_n10583_), .ZN(new_n10584_));
  OAI21_X1   g09565(.A1(new_n9998_), .A2(new_n10072_), .B(new_n10584_), .ZN(new_n10585_));
  NAND4_X1   g09566(.A1(new_n10071_), .A2(new_n10002_), .A3(new_n10568_), .A4(new_n10583_), .ZN(new_n10586_));
  XOR2_X1    g09567(.A1(new_n10574_), .A2(new_n10570_), .Z(new_n10587_));
  NOR2_X1    g09568(.A1(new_n10587_), .A2(new_n10572_), .ZN(new_n10588_));
  INV_X1     g09569(.I(new_n10588_), .ZN(new_n10589_));
  NAND3_X1   g09570(.A1(new_n10338_), .A2(new_n10323_), .A3(new_n10330_), .ZN(new_n10590_));
  AOI21_X1   g09571(.A1(new_n10460_), .A2(new_n10461_), .B(new_n10483_), .ZN(new_n10591_));
  NOR3_X1    g09572(.A1(new_n10467_), .A2(new_n10474_), .A3(new_n10466_), .ZN(new_n10592_));
  OAI21_X1   g09573(.A1(new_n10592_), .A2(new_n10591_), .B(new_n10459_), .ZN(new_n10593_));
  OAI21_X1   g09574(.A1(new_n10467_), .A2(new_n10466_), .B(new_n10474_), .ZN(new_n10594_));
  NAND3_X1   g09575(.A1(new_n10460_), .A2(new_n10461_), .A3(new_n10483_), .ZN(new_n10595_));
  NAND3_X1   g09576(.A1(new_n10594_), .A2(new_n10595_), .A3(new_n10464_), .ZN(new_n10596_));
  NAND3_X1   g09577(.A1(new_n10590_), .A2(new_n10593_), .A3(new_n10596_), .ZN(new_n10597_));
  NOR2_X1    g09578(.A1(new_n10331_), .A2(new_n10347_), .ZN(new_n10598_));
  AOI21_X1   g09579(.A1(new_n10594_), .A2(new_n10595_), .B(new_n10464_), .ZN(new_n10599_));
  NOR3_X1    g09580(.A1(new_n10592_), .A2(new_n10591_), .A3(new_n10459_), .ZN(new_n10600_));
  OAI21_X1   g09581(.A1(new_n10599_), .A2(new_n10600_), .B(new_n10598_), .ZN(new_n10601_));
  NAND2_X1   g09582(.A1(new_n10601_), .A2(new_n10597_), .ZN(new_n10602_));
  NAND2_X1   g09583(.A1(new_n10602_), .A2(new_n10589_), .ZN(new_n10603_));
  NAND3_X1   g09584(.A1(new_n10601_), .A2(new_n10597_), .A3(new_n10588_), .ZN(new_n10604_));
  NAND2_X1   g09585(.A1(new_n10603_), .A2(new_n10604_), .ZN(new_n10605_));
  AOI22_X1   g09586(.A1(new_n10605_), .A2(new_n10564_), .B1(new_n10585_), .B2(new_n10586_), .ZN(new_n10606_));
  OAI21_X1   g09587(.A1(new_n10552_), .A2(new_n10553_), .B(new_n10562_), .ZN(new_n10607_));
  AOI21_X1   g09588(.A1(new_n10606_), .A2(new_n10607_), .B(new_n10563_), .ZN(new_n10608_));
  AOI22_X1   g09589(.A1(new_n10069_), .A2(new_n10082_), .B1(new_n10541_), .B2(new_n10548_), .ZN(new_n10609_));
  OAI21_X1   g09590(.A1(new_n10608_), .A2(new_n10609_), .B(new_n10549_), .ZN(new_n10610_));
  NAND2_X1   g09591(.A1(new_n10025_), .A2(new_n10029_), .ZN(new_n10611_));
  NAND2_X1   g09592(.A1(new_n10024_), .A2(new_n10019_), .ZN(new_n10612_));
  NAND2_X1   g09593(.A1(new_n10611_), .A2(new_n10612_), .ZN(new_n10613_));
  NOR2_X1    g09594(.A1(new_n10024_), .A2(new_n10019_), .ZN(new_n10614_));
  INV_X1     g09595(.I(new_n10614_), .ZN(new_n10615_));
  NAND2_X1   g09596(.A1(new_n10613_), .A2(new_n10615_), .ZN(new_n10616_));
  INV_X1     g09597(.I(new_n10616_), .ZN(new_n10617_));
  NAND2_X1   g09598(.A1(new_n10056_), .A2(new_n10052_), .ZN(new_n10618_));
  OAI21_X1   g09599(.A1(new_n10059_), .A2(new_n10047_), .B(new_n10618_), .ZN(new_n10619_));
  NAND2_X1   g09600(.A1(new_n10059_), .A2(new_n10047_), .ZN(new_n10620_));
  NAND2_X1   g09601(.A1(new_n10619_), .A2(new_n10620_), .ZN(new_n10621_));
  XNOR2_X1   g09602(.A1(new_n10047_), .A2(new_n10043_), .ZN(new_n10622_));
  XOR2_X1    g09603(.A1(new_n10024_), .A2(new_n10019_), .Z(new_n10623_));
  NOR4_X1    g09604(.A1(new_n10622_), .A2(new_n10611_), .A3(new_n10623_), .A4(new_n10618_), .ZN(new_n10624_));
  OAI21_X1   g09605(.A1(new_n10015_), .A2(new_n10080_), .B(new_n10624_), .ZN(new_n10625_));
  NAND2_X1   g09606(.A1(new_n10625_), .A2(new_n10621_), .ZN(new_n10626_));
  AND2_X2    g09607(.A1(new_n10619_), .A2(new_n10620_), .Z(new_n10627_));
  NAND4_X1   g09608(.A1(new_n10035_), .A2(new_n10038_), .A3(new_n10065_), .A4(new_n10066_), .ZN(new_n10628_));
  INV_X1     g09609(.I(new_n10624_), .ZN(new_n10629_));
  AOI21_X1   g09610(.A1(new_n10077_), .A2(new_n10628_), .B(new_n10629_), .ZN(new_n10630_));
  NAND2_X1   g09611(.A1(new_n10630_), .A2(new_n10627_), .ZN(new_n10631_));
  AOI21_X1   g09612(.A1(new_n10626_), .A2(new_n10631_), .B(new_n10617_), .ZN(new_n10632_));
  NOR2_X1    g09613(.A1(new_n10630_), .A2(new_n10627_), .ZN(new_n10633_));
  NOR2_X1    g09614(.A1(new_n10625_), .A2(new_n10621_), .ZN(new_n10634_));
  NOR3_X1    g09615(.A1(new_n10634_), .A2(new_n10633_), .A3(new_n10616_), .ZN(new_n10635_));
  NOR2_X1    g09616(.A1(new_n10547_), .A2(new_n10545_), .ZN(new_n10636_));
  AOI21_X1   g09617(.A1(new_n10484_), .A2(new_n10482_), .B(new_n10380_), .ZN(new_n10637_));
  NOR3_X1    g09618(.A1(new_n10475_), .A2(new_n10462_), .A3(new_n10379_), .ZN(new_n10638_));
  OAI21_X1   g09619(.A1(new_n10638_), .A2(new_n10637_), .B(new_n10480_), .ZN(new_n10639_));
  AOI21_X1   g09620(.A1(new_n10476_), .A2(new_n10380_), .B(new_n10435_), .ZN(new_n10640_));
  NAND2_X1   g09621(.A1(new_n10639_), .A2(new_n10640_), .ZN(new_n10641_));
  NAND4_X1   g09622(.A1(new_n10641_), .A2(new_n10509_), .A3(new_n10515_), .A4(new_n10518_), .ZN(new_n10642_));
  OAI21_X1   g09623(.A1(new_n10475_), .A2(new_n10462_), .B(new_n10379_), .ZN(new_n10643_));
  NAND3_X1   g09624(.A1(new_n10484_), .A2(new_n10482_), .A3(new_n10380_), .ZN(new_n10644_));
  AOI21_X1   g09625(.A1(new_n10643_), .A2(new_n10644_), .B(new_n10498_), .ZN(new_n10645_));
  OAI21_X1   g09626(.A1(new_n10485_), .A2(new_n10379_), .B(new_n10502_), .ZN(new_n10646_));
  NOR2_X1    g09627(.A1(new_n10645_), .A2(new_n10646_), .ZN(new_n10647_));
  NAND3_X1   g09628(.A1(new_n10515_), .A2(new_n10509_), .A3(new_n10518_), .ZN(new_n10648_));
  NAND2_X1   g09629(.A1(new_n10648_), .A2(new_n10647_), .ZN(new_n10649_));
  OAI21_X1   g09630(.A1(new_n10527_), .A2(new_n10528_), .B(new_n10509_), .ZN(new_n10650_));
  NAND3_X1   g09631(.A1(new_n10515_), .A2(new_n10510_), .A3(new_n10518_), .ZN(new_n10651_));
  AOI21_X1   g09632(.A1(new_n10650_), .A2(new_n10651_), .B(new_n10520_), .ZN(new_n10652_));
  NAND3_X1   g09633(.A1(new_n10652_), .A2(new_n10642_), .A3(new_n10649_), .ZN(new_n10653_));
  INV_X1     g09634(.I(new_n10653_), .ZN(new_n10654_));
  AOI21_X1   g09635(.A1(new_n10642_), .A2(new_n10649_), .B(new_n10652_), .ZN(new_n10655_));
  NOR2_X1    g09636(.A1(new_n10654_), .A2(new_n10655_), .ZN(new_n10656_));
  NOR3_X1    g09637(.A1(new_n10656_), .A2(new_n10636_), .A3(new_n10546_), .ZN(new_n10657_));
  OAI22_X1   g09638(.A1(new_n10496_), .A2(new_n10537_), .B1(new_n10538_), .B2(new_n10539_), .ZN(new_n10658_));
  NAND2_X1   g09639(.A1(new_n10656_), .A2(new_n10658_), .ZN(new_n10659_));
  NOR2_X1    g09640(.A1(new_n10657_), .A2(new_n10659_), .ZN(new_n10660_));
  NOR3_X1    g09641(.A1(new_n10660_), .A2(new_n10632_), .A3(new_n10635_), .ZN(new_n10661_));
  XOR2_X1    g09642(.A1(new_n10621_), .A2(new_n10616_), .Z(new_n10662_));
  NAND2_X1   g09643(.A1(new_n10662_), .A2(new_n10625_), .ZN(new_n10663_));
  NAND2_X1   g09644(.A1(new_n10077_), .A2(new_n10628_), .ZN(new_n10664_));
  NAND3_X1   g09645(.A1(new_n10530_), .A2(new_n10533_), .A3(new_n10537_), .ZN(new_n10665_));
  OAI21_X1   g09646(.A1(new_n10539_), .A2(new_n10538_), .B(new_n10505_), .ZN(new_n10666_));
  NAND2_X1   g09647(.A1(new_n10666_), .A2(new_n10496_), .ZN(new_n10667_));
  NAND2_X1   g09648(.A1(new_n10667_), .A2(new_n10665_), .ZN(new_n10668_));
  NOR2_X1    g09649(.A1(new_n10621_), .A2(new_n10616_), .ZN(new_n10669_));
  INV_X1     g09650(.I(new_n10669_), .ZN(new_n10670_));
  NAND2_X1   g09651(.A1(new_n10621_), .A2(new_n10616_), .ZN(new_n10671_));
  AOI21_X1   g09652(.A1(new_n10670_), .A2(new_n10671_), .B(new_n10629_), .ZN(new_n10672_));
  OAI22_X1   g09653(.A1(new_n10664_), .A2(new_n10672_), .B1(new_n10668_), .B2(new_n10656_), .ZN(new_n10673_));
  OAI21_X1   g09654(.A1(new_n10673_), .A2(new_n10659_), .B(new_n10663_), .ZN(new_n10674_));
  OAI21_X1   g09655(.A1(new_n10661_), .A2(new_n10610_), .B(new_n10674_), .ZN(new_n10675_));
  AND4_X2    g09656(.A1(new_n10613_), .A2(new_n10619_), .A3(new_n10615_), .A4(new_n10620_), .Z(new_n10676_));
  NAND2_X1   g09657(.A1(new_n10625_), .A2(new_n10676_), .ZN(new_n10677_));
  INV_X1     g09658(.I(new_n10677_), .ZN(new_n10678_));
  NOR2_X1    g09659(.A1(new_n10636_), .A2(new_n10546_), .ZN(new_n10679_));
  AOI22_X1   g09660(.A1(new_n10515_), .A2(new_n10518_), .B1(new_n10509_), .B2(new_n10514_), .ZN(new_n10680_));
  NOR2_X1    g09661(.A1(new_n10509_), .A2(new_n10514_), .ZN(new_n10681_));
  NOR3_X1    g09662(.A1(new_n10680_), .A2(new_n10647_), .A3(new_n10681_), .ZN(new_n10682_));
  INV_X1     g09663(.I(new_n10682_), .ZN(new_n10683_));
  NAND2_X1   g09664(.A1(new_n10679_), .A2(new_n10683_), .ZN(new_n10684_));
  OAI21_X1   g09665(.A1(new_n10680_), .A2(new_n10681_), .B(new_n10647_), .ZN(new_n10685_));
  NAND4_X1   g09666(.A1(new_n10684_), .A2(new_n10678_), .A3(new_n10671_), .A4(new_n10685_), .ZN(new_n10686_));
  NAND3_X1   g09667(.A1(new_n10625_), .A2(new_n10671_), .A3(new_n10676_), .ZN(new_n10687_));
  OAI21_X1   g09668(.A1(new_n10668_), .A2(new_n10682_), .B(new_n10685_), .ZN(new_n10688_));
  AOI22_X1   g09669(.A1(new_n10675_), .A2(new_n10686_), .B1(new_n10687_), .B2(new_n10688_), .ZN(new_n10689_));
  INV_X1     g09670(.I(\A[958] ), .ZN(new_n10690_));
  NOR2_X1    g09671(.A1(\A[959] ), .A2(\A[960] ), .ZN(new_n10691_));
  NAND2_X1   g09672(.A1(\A[959] ), .A2(\A[960] ), .ZN(new_n10692_));
  AOI21_X1   g09673(.A1(new_n10690_), .A2(new_n10692_), .B(new_n10691_), .ZN(new_n10693_));
  INV_X1     g09674(.I(new_n10693_), .ZN(new_n10694_));
  INV_X1     g09675(.I(\A[955] ), .ZN(new_n10695_));
  NOR2_X1    g09676(.A1(\A[956] ), .A2(\A[957] ), .ZN(new_n10696_));
  NAND2_X1   g09677(.A1(\A[956] ), .A2(\A[957] ), .ZN(new_n10697_));
  AOI21_X1   g09678(.A1(new_n10695_), .A2(new_n10697_), .B(new_n10696_), .ZN(new_n10698_));
  INV_X1     g09679(.I(\A[956] ), .ZN(new_n10699_));
  NAND2_X1   g09680(.A1(new_n10699_), .A2(\A[957] ), .ZN(new_n10700_));
  INV_X1     g09681(.I(\A[957] ), .ZN(new_n10701_));
  NAND2_X1   g09682(.A1(new_n10701_), .A2(\A[956] ), .ZN(new_n10702_));
  AOI21_X1   g09683(.A1(new_n10700_), .A2(new_n10702_), .B(new_n10695_), .ZN(new_n10703_));
  INV_X1     g09684(.I(new_n10696_), .ZN(new_n10704_));
  AOI21_X1   g09685(.A1(new_n10704_), .A2(new_n10697_), .B(\A[955] ), .ZN(new_n10705_));
  NOR2_X1    g09686(.A1(new_n10705_), .A2(new_n10703_), .ZN(new_n10706_));
  INV_X1     g09687(.I(\A[959] ), .ZN(new_n10707_));
  NAND2_X1   g09688(.A1(new_n10707_), .A2(\A[960] ), .ZN(new_n10708_));
  INV_X1     g09689(.I(\A[960] ), .ZN(new_n10709_));
  NAND2_X1   g09690(.A1(new_n10709_), .A2(\A[959] ), .ZN(new_n10710_));
  AOI21_X1   g09691(.A1(new_n10708_), .A2(new_n10710_), .B(new_n10690_), .ZN(new_n10711_));
  INV_X1     g09692(.I(new_n10691_), .ZN(new_n10712_));
  AOI21_X1   g09693(.A1(new_n10712_), .A2(new_n10692_), .B(\A[958] ), .ZN(new_n10713_));
  NOR2_X1    g09694(.A1(new_n10713_), .A2(new_n10711_), .ZN(new_n10714_));
  NAND2_X1   g09695(.A1(new_n10706_), .A2(new_n10714_), .ZN(new_n10715_));
  NAND2_X1   g09696(.A1(new_n10715_), .A2(new_n10698_), .ZN(new_n10716_));
  INV_X1     g09697(.I(new_n10698_), .ZN(new_n10717_));
  NOR2_X1    g09698(.A1(new_n10701_), .A2(\A[956] ), .ZN(new_n10718_));
  NOR2_X1    g09699(.A1(new_n10699_), .A2(\A[957] ), .ZN(new_n10719_));
  OAI21_X1   g09700(.A1(new_n10718_), .A2(new_n10719_), .B(\A[955] ), .ZN(new_n10720_));
  INV_X1     g09701(.I(new_n10697_), .ZN(new_n10721_));
  OAI21_X1   g09702(.A1(new_n10721_), .A2(new_n10696_), .B(new_n10695_), .ZN(new_n10722_));
  NAND2_X1   g09703(.A1(new_n10720_), .A2(new_n10722_), .ZN(new_n10723_));
  NOR2_X1    g09704(.A1(new_n10709_), .A2(\A[959] ), .ZN(new_n10724_));
  NOR2_X1    g09705(.A1(new_n10707_), .A2(\A[960] ), .ZN(new_n10725_));
  OAI21_X1   g09706(.A1(new_n10724_), .A2(new_n10725_), .B(\A[958] ), .ZN(new_n10726_));
  INV_X1     g09707(.I(new_n10692_), .ZN(new_n10727_));
  OAI21_X1   g09708(.A1(new_n10727_), .A2(new_n10691_), .B(new_n10690_), .ZN(new_n10728_));
  NAND2_X1   g09709(.A1(new_n10726_), .A2(new_n10728_), .ZN(new_n10729_));
  NOR2_X1    g09710(.A1(new_n10723_), .A2(new_n10729_), .ZN(new_n10730_));
  NAND2_X1   g09711(.A1(new_n10730_), .A2(new_n10717_), .ZN(new_n10731_));
  AOI21_X1   g09712(.A1(new_n10731_), .A2(new_n10716_), .B(new_n10694_), .ZN(new_n10732_));
  NOR2_X1    g09713(.A1(new_n10730_), .A2(new_n10717_), .ZN(new_n10733_));
  NOR2_X1    g09714(.A1(new_n10715_), .A2(new_n10698_), .ZN(new_n10734_));
  NOR3_X1    g09715(.A1(new_n10733_), .A2(new_n10734_), .A3(new_n10693_), .ZN(new_n10735_));
  NOR2_X1    g09716(.A1(new_n10732_), .A2(new_n10735_), .ZN(new_n10736_));
  INV_X1     g09717(.I(new_n10736_), .ZN(new_n10737_));
  INV_X1     g09718(.I(\A[964] ), .ZN(new_n10738_));
  NOR2_X1    g09719(.A1(\A[965] ), .A2(\A[966] ), .ZN(new_n10739_));
  NAND2_X1   g09720(.A1(\A[965] ), .A2(\A[966] ), .ZN(new_n10740_));
  AOI21_X1   g09721(.A1(new_n10738_), .A2(new_n10740_), .B(new_n10739_), .ZN(new_n10741_));
  INV_X1     g09722(.I(new_n10741_), .ZN(new_n10742_));
  INV_X1     g09723(.I(\A[961] ), .ZN(new_n10743_));
  NOR2_X1    g09724(.A1(\A[962] ), .A2(\A[963] ), .ZN(new_n10744_));
  NAND2_X1   g09725(.A1(\A[962] ), .A2(\A[963] ), .ZN(new_n10745_));
  AOI21_X1   g09726(.A1(new_n10743_), .A2(new_n10745_), .B(new_n10744_), .ZN(new_n10746_));
  INV_X1     g09727(.I(new_n10746_), .ZN(new_n10747_));
  NOR2_X1    g09728(.A1(new_n10742_), .A2(new_n10747_), .ZN(new_n10748_));
  INV_X1     g09729(.I(new_n10748_), .ZN(new_n10749_));
  INV_X1     g09730(.I(\A[962] ), .ZN(new_n10750_));
  NAND2_X1   g09731(.A1(new_n10750_), .A2(\A[963] ), .ZN(new_n10751_));
  INV_X1     g09732(.I(\A[963] ), .ZN(new_n10752_));
  NAND2_X1   g09733(.A1(new_n10752_), .A2(\A[962] ), .ZN(new_n10753_));
  AOI21_X1   g09734(.A1(new_n10751_), .A2(new_n10753_), .B(new_n10743_), .ZN(new_n10754_));
  INV_X1     g09735(.I(new_n10744_), .ZN(new_n10755_));
  AOI21_X1   g09736(.A1(new_n10755_), .A2(new_n10745_), .B(\A[961] ), .ZN(new_n10756_));
  NOR2_X1    g09737(.A1(new_n10756_), .A2(new_n10754_), .ZN(new_n10757_));
  INV_X1     g09738(.I(\A[966] ), .ZN(new_n10758_));
  NOR2_X1    g09739(.A1(new_n10758_), .A2(\A[965] ), .ZN(new_n10759_));
  INV_X1     g09740(.I(\A[965] ), .ZN(new_n10760_));
  NOR2_X1    g09741(.A1(new_n10760_), .A2(\A[966] ), .ZN(new_n10761_));
  OAI21_X1   g09742(.A1(new_n10759_), .A2(new_n10761_), .B(\A[964] ), .ZN(new_n10762_));
  INV_X1     g09743(.I(new_n10740_), .ZN(new_n10763_));
  OAI21_X1   g09744(.A1(new_n10763_), .A2(new_n10739_), .B(new_n10738_), .ZN(new_n10764_));
  NAND2_X1   g09745(.A1(new_n10762_), .A2(new_n10764_), .ZN(new_n10765_));
  NAND2_X1   g09746(.A1(new_n10757_), .A2(new_n10765_), .ZN(new_n10766_));
  NOR2_X1    g09747(.A1(new_n10752_), .A2(\A[962] ), .ZN(new_n10767_));
  NOR2_X1    g09748(.A1(new_n10750_), .A2(\A[963] ), .ZN(new_n10768_));
  OAI21_X1   g09749(.A1(new_n10767_), .A2(new_n10768_), .B(\A[961] ), .ZN(new_n10769_));
  INV_X1     g09750(.I(new_n10745_), .ZN(new_n10770_));
  OAI21_X1   g09751(.A1(new_n10770_), .A2(new_n10744_), .B(new_n10743_), .ZN(new_n10771_));
  NAND2_X1   g09752(.A1(new_n10769_), .A2(new_n10771_), .ZN(new_n10772_));
  NAND2_X1   g09753(.A1(new_n10760_), .A2(\A[966] ), .ZN(new_n10773_));
  NAND2_X1   g09754(.A1(new_n10758_), .A2(\A[965] ), .ZN(new_n10774_));
  AOI21_X1   g09755(.A1(new_n10773_), .A2(new_n10774_), .B(new_n10738_), .ZN(new_n10775_));
  INV_X1     g09756(.I(new_n10739_), .ZN(new_n10776_));
  AOI21_X1   g09757(.A1(new_n10776_), .A2(new_n10740_), .B(\A[964] ), .ZN(new_n10777_));
  NOR2_X1    g09758(.A1(new_n10777_), .A2(new_n10775_), .ZN(new_n10778_));
  NAND2_X1   g09759(.A1(new_n10778_), .A2(new_n10772_), .ZN(new_n10779_));
  AOI21_X1   g09760(.A1(new_n10766_), .A2(new_n10779_), .B(new_n10749_), .ZN(new_n10780_));
  AOI21_X1   g09761(.A1(new_n10757_), .A2(new_n10778_), .B(new_n10747_), .ZN(new_n10781_));
  NOR3_X1    g09762(.A1(new_n10772_), .A2(new_n10765_), .A3(new_n10746_), .ZN(new_n10782_));
  OAI21_X1   g09763(.A1(new_n10781_), .A2(new_n10782_), .B(new_n10741_), .ZN(new_n10783_));
  INV_X1     g09764(.I(new_n10783_), .ZN(new_n10784_));
  NOR3_X1    g09765(.A1(new_n10781_), .A2(new_n10782_), .A3(new_n10741_), .ZN(new_n10785_));
  NOR3_X1    g09766(.A1(new_n10784_), .A2(new_n10780_), .A3(new_n10785_), .ZN(new_n10786_));
  NAND3_X1   g09767(.A1(new_n10748_), .A2(new_n10757_), .A3(new_n10778_), .ZN(new_n10787_));
  NAND2_X1   g09768(.A1(new_n10757_), .A2(new_n10778_), .ZN(new_n10788_));
  NAND2_X1   g09769(.A1(new_n10772_), .A2(new_n10765_), .ZN(new_n10789_));
  NAND2_X1   g09770(.A1(new_n10788_), .A2(new_n10789_), .ZN(new_n10790_));
  NAND2_X1   g09771(.A1(new_n10723_), .A2(new_n10729_), .ZN(new_n10791_));
  NAND2_X1   g09772(.A1(new_n10715_), .A2(new_n10791_), .ZN(new_n10792_));
  NAND3_X1   g09773(.A1(new_n10730_), .A2(new_n10693_), .A3(new_n10698_), .ZN(new_n10793_));
  NOR4_X1    g09774(.A1(new_n10790_), .A2(new_n10793_), .A3(new_n10792_), .A4(new_n10787_), .ZN(new_n10794_));
  NAND2_X1   g09775(.A1(new_n10786_), .A2(new_n10794_), .ZN(new_n10795_));
  OR3_X2     g09776(.A1(new_n10781_), .A2(new_n10782_), .A3(new_n10741_), .Z(new_n10796_));
  NAND2_X1   g09777(.A1(new_n10796_), .A2(new_n10783_), .ZN(new_n10797_));
  NOR2_X1    g09778(.A1(new_n10790_), .A2(new_n10787_), .ZN(new_n10798_));
  NOR2_X1    g09779(.A1(new_n10706_), .A2(new_n10714_), .ZN(new_n10799_));
  NOR2_X1    g09780(.A1(new_n10799_), .A2(new_n10730_), .ZN(new_n10800_));
  NAND2_X1   g09781(.A1(new_n10693_), .A2(new_n10698_), .ZN(new_n10801_));
  NOR2_X1    g09782(.A1(new_n10715_), .A2(new_n10801_), .ZN(new_n10802_));
  NAND3_X1   g09783(.A1(new_n10798_), .A2(new_n10800_), .A3(new_n10802_), .ZN(new_n10803_));
  OAI21_X1   g09784(.A1(new_n10797_), .A2(new_n10780_), .B(new_n10803_), .ZN(new_n10804_));
  AOI21_X1   g09785(.A1(new_n10804_), .A2(new_n10795_), .B(new_n10737_), .ZN(new_n10805_));
  NOR2_X1    g09786(.A1(new_n10786_), .A2(new_n10803_), .ZN(new_n10806_));
  NOR2_X1    g09787(.A1(new_n10784_), .A2(new_n10785_), .ZN(new_n10807_));
  NOR3_X1    g09788(.A1(new_n10790_), .A2(new_n10792_), .A3(new_n10787_), .ZN(new_n10808_));
  NOR2_X1    g09789(.A1(new_n10780_), .A2(new_n10793_), .ZN(new_n10809_));
  INV_X1     g09790(.I(new_n10809_), .ZN(new_n10810_));
  AOI21_X1   g09791(.A1(new_n10807_), .A2(new_n10808_), .B(new_n10810_), .ZN(new_n10811_));
  NOR3_X1    g09792(.A1(new_n10811_), .A2(new_n10806_), .A3(new_n10737_), .ZN(new_n10812_));
  NOR2_X1    g09793(.A1(new_n10805_), .A2(new_n10812_), .ZN(new_n10813_));
  NOR3_X1    g09794(.A1(new_n10803_), .A2(new_n10797_), .A3(new_n10780_), .ZN(new_n10814_));
  NOR2_X1    g09795(.A1(new_n10786_), .A2(new_n10794_), .ZN(new_n10815_));
  OAI21_X1   g09796(.A1(new_n10815_), .A2(new_n10814_), .B(new_n10736_), .ZN(new_n10816_));
  OAI21_X1   g09797(.A1(new_n10797_), .A2(new_n10780_), .B(new_n10794_), .ZN(new_n10817_));
  INV_X1     g09798(.I(new_n10787_), .ZN(new_n10818_));
  AND2_X2    g09799(.A1(new_n10788_), .A2(new_n10789_), .Z(new_n10819_));
  NAND3_X1   g09800(.A1(new_n10819_), .A2(new_n10818_), .A3(new_n10800_), .ZN(new_n10820_));
  OAI21_X1   g09801(.A1(new_n10797_), .A2(new_n10820_), .B(new_n10809_), .ZN(new_n10821_));
  NAND3_X1   g09802(.A1(new_n10821_), .A2(new_n10817_), .A3(new_n10736_), .ZN(new_n10822_));
  NOR2_X1    g09803(.A1(new_n10793_), .A2(new_n10792_), .ZN(new_n10823_));
  XOR2_X1    g09804(.A1(new_n10823_), .A2(new_n10798_), .Z(new_n10824_));
  INV_X1     g09805(.I(\A[949] ), .ZN(new_n10825_));
  INV_X1     g09806(.I(\A[950] ), .ZN(new_n10826_));
  NAND2_X1   g09807(.A1(new_n10826_), .A2(\A[951] ), .ZN(new_n10827_));
  INV_X1     g09808(.I(\A[951] ), .ZN(new_n10828_));
  NAND2_X1   g09809(.A1(new_n10828_), .A2(\A[950] ), .ZN(new_n10829_));
  AOI21_X1   g09810(.A1(new_n10827_), .A2(new_n10829_), .B(new_n10825_), .ZN(new_n10830_));
  NOR2_X1    g09811(.A1(\A[950] ), .A2(\A[951] ), .ZN(new_n10831_));
  INV_X1     g09812(.I(new_n10831_), .ZN(new_n10832_));
  NAND2_X1   g09813(.A1(\A[950] ), .A2(\A[951] ), .ZN(new_n10833_));
  AOI21_X1   g09814(.A1(new_n10832_), .A2(new_n10833_), .B(\A[949] ), .ZN(new_n10834_));
  NOR2_X1    g09815(.A1(new_n10834_), .A2(new_n10830_), .ZN(new_n10835_));
  INV_X1     g09816(.I(\A[952] ), .ZN(new_n10836_));
  INV_X1     g09817(.I(\A[953] ), .ZN(new_n10837_));
  NAND2_X1   g09818(.A1(new_n10837_), .A2(\A[954] ), .ZN(new_n10838_));
  INV_X1     g09819(.I(\A[954] ), .ZN(new_n10839_));
  NAND2_X1   g09820(.A1(new_n10839_), .A2(\A[953] ), .ZN(new_n10840_));
  AOI21_X1   g09821(.A1(new_n10838_), .A2(new_n10840_), .B(new_n10836_), .ZN(new_n10841_));
  NOR2_X1    g09822(.A1(\A[953] ), .A2(\A[954] ), .ZN(new_n10842_));
  INV_X1     g09823(.I(new_n10842_), .ZN(new_n10843_));
  NAND2_X1   g09824(.A1(\A[953] ), .A2(\A[954] ), .ZN(new_n10844_));
  AOI21_X1   g09825(.A1(new_n10843_), .A2(new_n10844_), .B(\A[952] ), .ZN(new_n10845_));
  NOR2_X1    g09826(.A1(new_n10845_), .A2(new_n10841_), .ZN(new_n10846_));
  NAND2_X1   g09827(.A1(new_n10835_), .A2(new_n10846_), .ZN(new_n10847_));
  AOI21_X1   g09828(.A1(new_n10836_), .A2(new_n10844_), .B(new_n10842_), .ZN(new_n10848_));
  AOI21_X1   g09829(.A1(new_n10825_), .A2(new_n10833_), .B(new_n10831_), .ZN(new_n10849_));
  NAND2_X1   g09830(.A1(new_n10848_), .A2(new_n10849_), .ZN(new_n10850_));
  NOR2_X1    g09831(.A1(new_n10828_), .A2(\A[950] ), .ZN(new_n10851_));
  NOR2_X1    g09832(.A1(new_n10826_), .A2(\A[951] ), .ZN(new_n10852_));
  OAI21_X1   g09833(.A1(new_n10851_), .A2(new_n10852_), .B(\A[949] ), .ZN(new_n10853_));
  INV_X1     g09834(.I(new_n10833_), .ZN(new_n10854_));
  OAI21_X1   g09835(.A1(new_n10854_), .A2(new_n10831_), .B(new_n10825_), .ZN(new_n10855_));
  NAND2_X1   g09836(.A1(new_n10853_), .A2(new_n10855_), .ZN(new_n10856_));
  NOR2_X1    g09837(.A1(new_n10839_), .A2(\A[953] ), .ZN(new_n10857_));
  NOR2_X1    g09838(.A1(new_n10837_), .A2(\A[954] ), .ZN(new_n10858_));
  OAI21_X1   g09839(.A1(new_n10857_), .A2(new_n10858_), .B(\A[952] ), .ZN(new_n10859_));
  INV_X1     g09840(.I(new_n10844_), .ZN(new_n10860_));
  OAI21_X1   g09841(.A1(new_n10860_), .A2(new_n10842_), .B(new_n10836_), .ZN(new_n10861_));
  NAND2_X1   g09842(.A1(new_n10859_), .A2(new_n10861_), .ZN(new_n10862_));
  NAND2_X1   g09843(.A1(new_n10856_), .A2(new_n10862_), .ZN(new_n10863_));
  NAND2_X1   g09844(.A1(new_n10847_), .A2(new_n10863_), .ZN(new_n10864_));
  NOR3_X1    g09845(.A1(new_n10864_), .A2(new_n10847_), .A3(new_n10850_), .ZN(new_n10865_));
  INV_X1     g09846(.I(\A[943] ), .ZN(new_n10866_));
  INV_X1     g09847(.I(\A[944] ), .ZN(new_n10867_));
  NAND2_X1   g09848(.A1(new_n10867_), .A2(\A[945] ), .ZN(new_n10868_));
  INV_X1     g09849(.I(\A[945] ), .ZN(new_n10869_));
  NAND2_X1   g09850(.A1(new_n10869_), .A2(\A[944] ), .ZN(new_n10870_));
  AOI21_X1   g09851(.A1(new_n10868_), .A2(new_n10870_), .B(new_n10866_), .ZN(new_n10871_));
  NOR2_X1    g09852(.A1(\A[944] ), .A2(\A[945] ), .ZN(new_n10872_));
  INV_X1     g09853(.I(new_n10872_), .ZN(new_n10873_));
  NAND2_X1   g09854(.A1(\A[944] ), .A2(\A[945] ), .ZN(new_n10874_));
  AOI21_X1   g09855(.A1(new_n10873_), .A2(new_n10874_), .B(\A[943] ), .ZN(new_n10875_));
  NOR2_X1    g09856(.A1(new_n10875_), .A2(new_n10871_), .ZN(new_n10876_));
  INV_X1     g09857(.I(\A[946] ), .ZN(new_n10877_));
  INV_X1     g09858(.I(\A[947] ), .ZN(new_n10878_));
  NAND2_X1   g09859(.A1(new_n10878_), .A2(\A[948] ), .ZN(new_n10879_));
  INV_X1     g09860(.I(\A[948] ), .ZN(new_n10880_));
  NAND2_X1   g09861(.A1(new_n10880_), .A2(\A[947] ), .ZN(new_n10881_));
  AOI21_X1   g09862(.A1(new_n10879_), .A2(new_n10881_), .B(new_n10877_), .ZN(new_n10882_));
  NOR2_X1    g09863(.A1(\A[947] ), .A2(\A[948] ), .ZN(new_n10883_));
  INV_X1     g09864(.I(new_n10883_), .ZN(new_n10884_));
  NAND2_X1   g09865(.A1(\A[947] ), .A2(\A[948] ), .ZN(new_n10885_));
  AOI21_X1   g09866(.A1(new_n10884_), .A2(new_n10885_), .B(\A[946] ), .ZN(new_n10886_));
  NOR2_X1    g09867(.A1(new_n10886_), .A2(new_n10882_), .ZN(new_n10887_));
  AOI21_X1   g09868(.A1(new_n10877_), .A2(new_n10885_), .B(new_n10883_), .ZN(new_n10888_));
  AOI21_X1   g09869(.A1(new_n10866_), .A2(new_n10874_), .B(new_n10872_), .ZN(new_n10889_));
  NAND2_X1   g09870(.A1(new_n10888_), .A2(new_n10889_), .ZN(new_n10890_));
  NOR2_X1    g09871(.A1(new_n10824_), .A2(new_n10865_), .ZN(new_n10892_));
  AOI21_X1   g09872(.A1(new_n10816_), .A2(new_n10822_), .B(new_n10892_), .ZN(new_n10893_));
  NAND2_X1   g09873(.A1(new_n10800_), .A2(new_n10802_), .ZN(new_n10894_));
  XOR2_X1    g09874(.A1(new_n10798_), .A2(new_n10894_), .Z(new_n10895_));
  NOR2_X1    g09875(.A1(new_n10847_), .A2(new_n10850_), .ZN(new_n10896_));
  NAND3_X1   g09876(.A1(new_n10896_), .A2(new_n10847_), .A3(new_n10863_), .ZN(new_n10897_));
  NAND2_X1   g09877(.A1(new_n10895_), .A2(new_n10897_), .ZN(new_n10898_));
  NOR3_X1    g09878(.A1(new_n10812_), .A2(new_n10805_), .A3(new_n10898_), .ZN(new_n10899_));
  NAND2_X1   g09879(.A1(new_n10876_), .A2(new_n10887_), .ZN(new_n10900_));
  NOR2_X1    g09880(.A1(new_n10869_), .A2(\A[944] ), .ZN(new_n10901_));
  NOR2_X1    g09881(.A1(new_n10867_), .A2(\A[945] ), .ZN(new_n10902_));
  OAI21_X1   g09882(.A1(new_n10901_), .A2(new_n10902_), .B(\A[943] ), .ZN(new_n10903_));
  INV_X1     g09883(.I(new_n10874_), .ZN(new_n10904_));
  OAI21_X1   g09884(.A1(new_n10904_), .A2(new_n10872_), .B(new_n10866_), .ZN(new_n10905_));
  NAND2_X1   g09885(.A1(new_n10903_), .A2(new_n10905_), .ZN(new_n10906_));
  NOR2_X1    g09886(.A1(new_n10880_), .A2(\A[947] ), .ZN(new_n10907_));
  NOR2_X1    g09887(.A1(new_n10878_), .A2(\A[948] ), .ZN(new_n10908_));
  OAI21_X1   g09888(.A1(new_n10907_), .A2(new_n10908_), .B(\A[946] ), .ZN(new_n10909_));
  INV_X1     g09889(.I(new_n10885_), .ZN(new_n10910_));
  OAI21_X1   g09890(.A1(new_n10910_), .A2(new_n10883_), .B(new_n10877_), .ZN(new_n10911_));
  NAND2_X1   g09891(.A1(new_n10909_), .A2(new_n10911_), .ZN(new_n10912_));
  NAND2_X1   g09892(.A1(new_n10906_), .A2(new_n10912_), .ZN(new_n10913_));
  AND2_X2    g09893(.A1(new_n10900_), .A2(new_n10913_), .Z(new_n10914_));
  INV_X1     g09894(.I(new_n10849_), .ZN(new_n10915_));
  AOI21_X1   g09895(.A1(new_n10835_), .A2(new_n10846_), .B(new_n10915_), .ZN(new_n10916_));
  NAND3_X1   g09896(.A1(new_n10835_), .A2(new_n10846_), .A3(new_n10915_), .ZN(new_n10917_));
  INV_X1     g09897(.I(new_n10917_), .ZN(new_n10918_));
  OAI21_X1   g09898(.A1(new_n10918_), .A2(new_n10916_), .B(new_n10848_), .ZN(new_n10919_));
  INV_X1     g09899(.I(new_n10848_), .ZN(new_n10920_));
  INV_X1     g09900(.I(new_n10916_), .ZN(new_n10921_));
  NAND3_X1   g09901(.A1(new_n10921_), .A2(new_n10920_), .A3(new_n10917_), .ZN(new_n10922_));
  NAND4_X1   g09902(.A1(new_n10865_), .A2(new_n10922_), .A3(new_n10919_), .A4(new_n10914_), .ZN(new_n10923_));
  NOR2_X1    g09903(.A1(new_n10900_), .A2(new_n10890_), .ZN(new_n10924_));
  INV_X1     g09904(.I(new_n10850_), .ZN(new_n10925_));
  NOR2_X1    g09905(.A1(new_n10846_), .A2(new_n10856_), .ZN(new_n10926_));
  NOR2_X1    g09906(.A1(new_n10835_), .A2(new_n10862_), .ZN(new_n10927_));
  OAI21_X1   g09907(.A1(new_n10926_), .A2(new_n10927_), .B(new_n10925_), .ZN(new_n10928_));
  AND2_X2    g09908(.A1(new_n10928_), .A2(new_n10924_), .Z(new_n10929_));
  INV_X1     g09909(.I(new_n10888_), .ZN(new_n10930_));
  OAI21_X1   g09910(.A1(new_n10906_), .A2(new_n10912_), .B(new_n10889_), .ZN(new_n10931_));
  INV_X1     g09911(.I(new_n10889_), .ZN(new_n10932_));
  NAND3_X1   g09912(.A1(new_n10876_), .A2(new_n10887_), .A3(new_n10932_), .ZN(new_n10933_));
  AOI21_X1   g09913(.A1(new_n10931_), .A2(new_n10933_), .B(new_n10930_), .ZN(new_n10934_));
  INV_X1     g09914(.I(new_n10934_), .ZN(new_n10935_));
  NAND3_X1   g09915(.A1(new_n10931_), .A2(new_n10933_), .A3(new_n10930_), .ZN(new_n10936_));
  NAND2_X1   g09916(.A1(new_n10935_), .A2(new_n10936_), .ZN(new_n10937_));
  NAND3_X1   g09917(.A1(new_n10923_), .A2(new_n10929_), .A3(new_n10937_), .ZN(new_n10938_));
  INV_X1     g09918(.I(new_n10938_), .ZN(new_n10939_));
  AND2_X2    g09919(.A1(new_n10847_), .A2(new_n10863_), .Z(new_n10940_));
  NAND4_X1   g09920(.A1(new_n10914_), .A2(new_n10940_), .A3(new_n10896_), .A4(new_n10924_), .ZN(new_n10941_));
  NAND2_X1   g09921(.A1(new_n10937_), .A2(new_n10941_), .ZN(new_n10942_));
  NAND3_X1   g09922(.A1(new_n10922_), .A2(new_n10919_), .A3(new_n10928_), .ZN(new_n10943_));
  OAI21_X1   g09923(.A1(new_n10937_), .A2(new_n10941_), .B(new_n10943_), .ZN(new_n10944_));
  AOI21_X1   g09924(.A1(new_n10921_), .A2(new_n10917_), .B(new_n10920_), .ZN(new_n10945_));
  NOR3_X1    g09925(.A1(new_n10918_), .A2(new_n10848_), .A3(new_n10916_), .ZN(new_n10946_));
  INV_X1     g09926(.I(new_n10928_), .ZN(new_n10947_));
  NOR3_X1    g09927(.A1(new_n10945_), .A2(new_n10947_), .A3(new_n10946_), .ZN(new_n10948_));
  NAND3_X1   g09928(.A1(new_n10924_), .A2(new_n10900_), .A3(new_n10913_), .ZN(new_n10949_));
  INV_X1     g09929(.I(new_n10936_), .ZN(new_n10950_));
  NOR4_X1    g09930(.A1(new_n10950_), .A2(new_n10897_), .A3(new_n10949_), .A4(new_n10934_), .ZN(new_n10951_));
  NAND2_X1   g09931(.A1(new_n10951_), .A2(new_n10948_), .ZN(new_n10952_));
  NAND2_X1   g09932(.A1(new_n10944_), .A2(new_n10952_), .ZN(new_n10953_));
  AOI21_X1   g09933(.A1(new_n10953_), .A2(new_n10942_), .B(new_n10939_), .ZN(new_n10954_));
  OAI22_X1   g09934(.A1(new_n10893_), .A2(new_n10899_), .B1(new_n10954_), .B2(new_n10813_), .ZN(new_n10955_));
  AOI21_X1   g09935(.A1(new_n10737_), .A2(new_n10817_), .B(new_n10811_), .ZN(new_n10956_));
  NOR2_X1    g09936(.A1(new_n10741_), .A2(new_n10746_), .ZN(new_n10957_));
  OAI21_X1   g09937(.A1(new_n10788_), .A2(new_n10957_), .B(new_n10749_), .ZN(new_n10958_));
  NOR2_X1    g09938(.A1(new_n10693_), .A2(new_n10698_), .ZN(new_n10959_));
  OAI21_X1   g09939(.A1(new_n10715_), .A2(new_n10959_), .B(new_n10801_), .ZN(new_n10960_));
  XNOR2_X1   g09940(.A1(new_n10958_), .A2(new_n10960_), .ZN(new_n10961_));
  NAND2_X1   g09941(.A1(new_n10956_), .A2(new_n10961_), .ZN(new_n10962_));
  NAND2_X1   g09942(.A1(new_n10923_), .A2(new_n10929_), .ZN(new_n10963_));
  OAI21_X1   g09943(.A1(new_n10948_), .A2(new_n10941_), .B(new_n10937_), .ZN(new_n10964_));
  NOR2_X1    g09944(.A1(new_n10848_), .A2(new_n10849_), .ZN(new_n10965_));
  OAI21_X1   g09945(.A1(new_n10847_), .A2(new_n10965_), .B(new_n10850_), .ZN(new_n10966_));
  NOR2_X1    g09946(.A1(new_n10888_), .A2(new_n10889_), .ZN(new_n10967_));
  OAI21_X1   g09947(.A1(new_n10900_), .A2(new_n10967_), .B(new_n10890_), .ZN(new_n10968_));
  XNOR2_X1   g09948(.A1(new_n10966_), .A2(new_n10968_), .ZN(new_n10969_));
  NAND3_X1   g09949(.A1(new_n10964_), .A2(new_n10963_), .A3(new_n10969_), .ZN(new_n10970_));
  INV_X1     g09950(.I(new_n10970_), .ZN(new_n10971_));
  XOR2_X1    g09951(.A1(new_n10962_), .A2(new_n10971_), .Z(new_n10972_));
  NOR2_X1    g09952(.A1(new_n10972_), .A2(new_n10955_), .ZN(new_n10973_));
  NAND2_X1   g09953(.A1(new_n10816_), .A2(new_n10822_), .ZN(new_n10974_));
  OAI21_X1   g09954(.A1(new_n10805_), .A2(new_n10812_), .B(new_n10898_), .ZN(new_n10975_));
  NAND3_X1   g09955(.A1(new_n10816_), .A2(new_n10892_), .A3(new_n10822_), .ZN(new_n10976_));
  NOR2_X1    g09956(.A1(new_n10951_), .A2(new_n10948_), .ZN(new_n10977_));
  NOR3_X1    g09957(.A1(new_n10943_), .A2(new_n10937_), .A3(new_n10941_), .ZN(new_n10978_));
  OAI21_X1   g09958(.A1(new_n10977_), .A2(new_n10978_), .B(new_n10942_), .ZN(new_n10979_));
  NAND2_X1   g09959(.A1(new_n10979_), .A2(new_n10938_), .ZN(new_n10980_));
  AOI22_X1   g09960(.A1(new_n10975_), .A2(new_n10976_), .B1(new_n10980_), .B2(new_n10974_), .ZN(new_n10981_));
  NAND2_X1   g09961(.A1(new_n10962_), .A2(new_n10970_), .ZN(new_n10982_));
  NOR2_X1    g09962(.A1(new_n10962_), .A2(new_n10970_), .ZN(new_n10983_));
  INV_X1     g09963(.I(new_n10983_), .ZN(new_n10984_));
  AOI21_X1   g09964(.A1(new_n10984_), .A2(new_n10982_), .B(new_n10981_), .ZN(new_n10985_));
  INV_X1     g09965(.I(\A[988] ), .ZN(new_n10986_));
  NOR2_X1    g09966(.A1(\A[989] ), .A2(\A[990] ), .ZN(new_n10987_));
  NAND2_X1   g09967(.A1(\A[989] ), .A2(\A[990] ), .ZN(new_n10988_));
  AOI21_X1   g09968(.A1(new_n10986_), .A2(new_n10988_), .B(new_n10987_), .ZN(new_n10989_));
  INV_X1     g09969(.I(new_n10989_), .ZN(new_n10990_));
  INV_X1     g09970(.I(\A[985] ), .ZN(new_n10991_));
  NOR2_X1    g09971(.A1(\A[986] ), .A2(\A[987] ), .ZN(new_n10992_));
  NAND2_X1   g09972(.A1(\A[986] ), .A2(\A[987] ), .ZN(new_n10993_));
  AOI21_X1   g09973(.A1(new_n10991_), .A2(new_n10993_), .B(new_n10992_), .ZN(new_n10994_));
  INV_X1     g09974(.I(\A[986] ), .ZN(new_n10995_));
  NAND2_X1   g09975(.A1(new_n10995_), .A2(\A[987] ), .ZN(new_n10996_));
  INV_X1     g09976(.I(\A[987] ), .ZN(new_n10997_));
  NAND2_X1   g09977(.A1(new_n10997_), .A2(\A[986] ), .ZN(new_n10998_));
  AOI21_X1   g09978(.A1(new_n10996_), .A2(new_n10998_), .B(new_n10991_), .ZN(new_n10999_));
  INV_X1     g09979(.I(new_n10992_), .ZN(new_n11000_));
  AOI21_X1   g09980(.A1(new_n11000_), .A2(new_n10993_), .B(\A[985] ), .ZN(new_n11001_));
  NOR2_X1    g09981(.A1(new_n11001_), .A2(new_n10999_), .ZN(new_n11002_));
  INV_X1     g09982(.I(\A[989] ), .ZN(new_n11003_));
  NAND2_X1   g09983(.A1(new_n11003_), .A2(\A[990] ), .ZN(new_n11004_));
  INV_X1     g09984(.I(\A[990] ), .ZN(new_n11005_));
  NAND2_X1   g09985(.A1(new_n11005_), .A2(\A[989] ), .ZN(new_n11006_));
  AOI21_X1   g09986(.A1(new_n11004_), .A2(new_n11006_), .B(new_n10986_), .ZN(new_n11007_));
  INV_X1     g09987(.I(new_n10987_), .ZN(new_n11008_));
  AOI21_X1   g09988(.A1(new_n11008_), .A2(new_n10988_), .B(\A[988] ), .ZN(new_n11009_));
  NOR2_X1    g09989(.A1(new_n11009_), .A2(new_n11007_), .ZN(new_n11010_));
  NAND2_X1   g09990(.A1(new_n11002_), .A2(new_n11010_), .ZN(new_n11011_));
  NAND2_X1   g09991(.A1(new_n11011_), .A2(new_n10994_), .ZN(new_n11012_));
  INV_X1     g09992(.I(new_n10994_), .ZN(new_n11013_));
  NOR2_X1    g09993(.A1(new_n10997_), .A2(\A[986] ), .ZN(new_n11014_));
  NOR2_X1    g09994(.A1(new_n10995_), .A2(\A[987] ), .ZN(new_n11015_));
  OAI21_X1   g09995(.A1(new_n11014_), .A2(new_n11015_), .B(\A[985] ), .ZN(new_n11016_));
  INV_X1     g09996(.I(new_n10993_), .ZN(new_n11017_));
  OAI21_X1   g09997(.A1(new_n11017_), .A2(new_n10992_), .B(new_n10991_), .ZN(new_n11018_));
  NAND2_X1   g09998(.A1(new_n11016_), .A2(new_n11018_), .ZN(new_n11019_));
  NOR2_X1    g09999(.A1(new_n11005_), .A2(\A[989] ), .ZN(new_n11020_));
  NOR2_X1    g10000(.A1(new_n11003_), .A2(\A[990] ), .ZN(new_n11021_));
  OAI21_X1   g10001(.A1(new_n11020_), .A2(new_n11021_), .B(\A[988] ), .ZN(new_n11022_));
  INV_X1     g10002(.I(new_n10988_), .ZN(new_n11023_));
  OAI21_X1   g10003(.A1(new_n11023_), .A2(new_n10987_), .B(new_n10986_), .ZN(new_n11024_));
  NAND2_X1   g10004(.A1(new_n11022_), .A2(new_n11024_), .ZN(new_n11025_));
  NOR2_X1    g10005(.A1(new_n11019_), .A2(new_n11025_), .ZN(new_n11026_));
  NAND2_X1   g10006(.A1(new_n11026_), .A2(new_n11013_), .ZN(new_n11027_));
  AOI21_X1   g10007(.A1(new_n11027_), .A2(new_n11012_), .B(new_n10990_), .ZN(new_n11028_));
  NOR2_X1    g10008(.A1(new_n11026_), .A2(new_n11013_), .ZN(new_n11029_));
  NOR2_X1    g10009(.A1(new_n11011_), .A2(new_n10994_), .ZN(new_n11030_));
  NOR3_X1    g10010(.A1(new_n11029_), .A2(new_n11030_), .A3(new_n10989_), .ZN(new_n11031_));
  INV_X1     g10011(.I(\A[979] ), .ZN(new_n11032_));
  INV_X1     g10012(.I(\A[980] ), .ZN(new_n11033_));
  NAND2_X1   g10013(.A1(new_n11033_), .A2(\A[981] ), .ZN(new_n11034_));
  INV_X1     g10014(.I(\A[981] ), .ZN(new_n11035_));
  NAND2_X1   g10015(.A1(new_n11035_), .A2(\A[980] ), .ZN(new_n11036_));
  AOI21_X1   g10016(.A1(new_n11034_), .A2(new_n11036_), .B(new_n11032_), .ZN(new_n11037_));
  NOR2_X1    g10017(.A1(\A[980] ), .A2(\A[981] ), .ZN(new_n11038_));
  INV_X1     g10018(.I(new_n11038_), .ZN(new_n11039_));
  NAND2_X1   g10019(.A1(\A[980] ), .A2(\A[981] ), .ZN(new_n11040_));
  AOI21_X1   g10020(.A1(new_n11039_), .A2(new_n11040_), .B(\A[979] ), .ZN(new_n11041_));
  NOR2_X1    g10021(.A1(new_n11041_), .A2(new_n11037_), .ZN(new_n11042_));
  INV_X1     g10022(.I(\A[982] ), .ZN(new_n11043_));
  INV_X1     g10023(.I(\A[983] ), .ZN(new_n11044_));
  NAND2_X1   g10024(.A1(new_n11044_), .A2(\A[984] ), .ZN(new_n11045_));
  INV_X1     g10025(.I(\A[984] ), .ZN(new_n11046_));
  NAND2_X1   g10026(.A1(new_n11046_), .A2(\A[983] ), .ZN(new_n11047_));
  AOI21_X1   g10027(.A1(new_n11045_), .A2(new_n11047_), .B(new_n11043_), .ZN(new_n11048_));
  NOR2_X1    g10028(.A1(\A[983] ), .A2(\A[984] ), .ZN(new_n11049_));
  INV_X1     g10029(.I(new_n11049_), .ZN(new_n11050_));
  NAND2_X1   g10030(.A1(\A[983] ), .A2(\A[984] ), .ZN(new_n11051_));
  AOI21_X1   g10031(.A1(new_n11050_), .A2(new_n11051_), .B(\A[982] ), .ZN(new_n11052_));
  NOR2_X1    g10032(.A1(new_n11052_), .A2(new_n11048_), .ZN(new_n11053_));
  NAND2_X1   g10033(.A1(new_n11042_), .A2(new_n11053_), .ZN(new_n11054_));
  NOR2_X1    g10034(.A1(new_n11035_), .A2(\A[980] ), .ZN(new_n11055_));
  NOR2_X1    g10035(.A1(new_n11033_), .A2(\A[981] ), .ZN(new_n11056_));
  OAI21_X1   g10036(.A1(new_n11055_), .A2(new_n11056_), .B(\A[979] ), .ZN(new_n11057_));
  INV_X1     g10037(.I(new_n11040_), .ZN(new_n11058_));
  OAI21_X1   g10038(.A1(new_n11058_), .A2(new_n11038_), .B(new_n11032_), .ZN(new_n11059_));
  NAND2_X1   g10039(.A1(new_n11057_), .A2(new_n11059_), .ZN(new_n11060_));
  NOR2_X1    g10040(.A1(new_n11046_), .A2(\A[983] ), .ZN(new_n11061_));
  NOR2_X1    g10041(.A1(new_n11044_), .A2(\A[984] ), .ZN(new_n11062_));
  OAI21_X1   g10042(.A1(new_n11061_), .A2(new_n11062_), .B(\A[982] ), .ZN(new_n11063_));
  INV_X1     g10043(.I(new_n11051_), .ZN(new_n11064_));
  OAI21_X1   g10044(.A1(new_n11064_), .A2(new_n11049_), .B(new_n11043_), .ZN(new_n11065_));
  NAND2_X1   g10045(.A1(new_n11063_), .A2(new_n11065_), .ZN(new_n11066_));
  NAND2_X1   g10046(.A1(new_n11060_), .A2(new_n11066_), .ZN(new_n11067_));
  NAND2_X1   g10047(.A1(new_n11019_), .A2(new_n11025_), .ZN(new_n11068_));
  NAND4_X1   g10048(.A1(new_n11011_), .A2(new_n11054_), .A3(new_n11067_), .A4(new_n11068_), .ZN(new_n11069_));
  NAND2_X1   g10049(.A1(new_n10989_), .A2(new_n10994_), .ZN(new_n11070_));
  NOR2_X1    g10050(.A1(new_n11011_), .A2(new_n11070_), .ZN(new_n11071_));
  AOI21_X1   g10051(.A1(new_n11043_), .A2(new_n11051_), .B(new_n11049_), .ZN(new_n11072_));
  AOI21_X1   g10052(.A1(new_n11032_), .A2(new_n11040_), .B(new_n11038_), .ZN(new_n11073_));
  NAND4_X1   g10053(.A1(new_n11042_), .A2(new_n11053_), .A3(new_n11072_), .A4(new_n11073_), .ZN(new_n11074_));
  NOR3_X1    g10054(.A1(new_n11069_), .A2(new_n11071_), .A3(new_n11074_), .ZN(new_n11075_));
  NOR3_X1    g10055(.A1(new_n11075_), .A2(new_n11028_), .A3(new_n11031_), .ZN(new_n11076_));
  NOR2_X1    g10056(.A1(new_n11060_), .A2(new_n11066_), .ZN(new_n11077_));
  INV_X1     g10057(.I(new_n11073_), .ZN(new_n11078_));
  NOR2_X1    g10058(.A1(new_n11077_), .A2(new_n11078_), .ZN(new_n11079_));
  NOR2_X1    g10059(.A1(new_n11054_), .A2(new_n11073_), .ZN(new_n11080_));
  OAI21_X1   g10060(.A1(new_n11079_), .A2(new_n11080_), .B(new_n11072_), .ZN(new_n11081_));
  INV_X1     g10061(.I(new_n11072_), .ZN(new_n11082_));
  NAND2_X1   g10062(.A1(new_n11054_), .A2(new_n11073_), .ZN(new_n11083_));
  NAND2_X1   g10063(.A1(new_n11077_), .A2(new_n11078_), .ZN(new_n11084_));
  NAND3_X1   g10064(.A1(new_n11084_), .A2(new_n11083_), .A3(new_n11082_), .ZN(new_n11085_));
  NAND2_X1   g10065(.A1(new_n11081_), .A2(new_n11085_), .ZN(new_n11086_));
  NAND2_X1   g10066(.A1(new_n11072_), .A2(new_n11073_), .ZN(new_n11087_));
  NOR2_X1    g10067(.A1(new_n11054_), .A2(new_n11087_), .ZN(new_n11088_));
  INV_X1     g10068(.I(new_n11070_), .ZN(new_n11089_));
  NAND2_X1   g10069(.A1(new_n11068_), .A2(new_n11089_), .ZN(new_n11090_));
  NAND2_X1   g10070(.A1(new_n11088_), .A2(new_n11090_), .ZN(new_n11091_));
  XNOR2_X1   g10071(.A1(new_n10989_), .A2(new_n10994_), .ZN(new_n11092_));
  NOR2_X1    g10072(.A1(new_n11011_), .A2(new_n11092_), .ZN(new_n11093_));
  NAND2_X1   g10073(.A1(new_n10990_), .A2(new_n11013_), .ZN(new_n11094_));
  AOI21_X1   g10074(.A1(new_n11070_), .A2(new_n11094_), .B(new_n11026_), .ZN(new_n11095_));
  NOR4_X1    g10075(.A1(new_n11091_), .A2(new_n11069_), .A3(new_n11093_), .A4(new_n11095_), .ZN(new_n11096_));
  NOR3_X1    g10076(.A1(new_n11076_), .A2(new_n11096_), .A3(new_n11086_), .ZN(new_n11097_));
  NAND2_X1   g10077(.A1(new_n11026_), .A2(new_n11089_), .ZN(new_n11098_));
  NAND2_X1   g10078(.A1(new_n11088_), .A2(new_n11098_), .ZN(new_n11099_));
  OAI22_X1   g10079(.A1(new_n11028_), .A2(new_n11031_), .B1(new_n11099_), .B2(new_n11069_), .ZN(new_n11100_));
  OAI21_X1   g10080(.A1(new_n11029_), .A2(new_n11030_), .B(new_n10989_), .ZN(new_n11101_));
  NAND3_X1   g10081(.A1(new_n11027_), .A2(new_n11012_), .A3(new_n10990_), .ZN(new_n11102_));
  NOR2_X1    g10082(.A1(new_n11042_), .A2(new_n11053_), .ZN(new_n11103_));
  NOR2_X1    g10083(.A1(new_n11002_), .A2(new_n11010_), .ZN(new_n11104_));
  NOR4_X1    g10084(.A1(new_n11026_), .A2(new_n11103_), .A3(new_n11104_), .A4(new_n11077_), .ZN(new_n11105_));
  NOR2_X1    g10085(.A1(new_n11071_), .A2(new_n11074_), .ZN(new_n11106_));
  NAND4_X1   g10086(.A1(new_n11101_), .A2(new_n11102_), .A3(new_n11106_), .A4(new_n11105_), .ZN(new_n11107_));
  AOI21_X1   g10087(.A1(new_n11100_), .A2(new_n11107_), .B(new_n11086_), .ZN(new_n11108_));
  NOR2_X1    g10088(.A1(new_n11097_), .A2(new_n11108_), .ZN(new_n11109_));
  NAND2_X1   g10089(.A1(new_n11106_), .A2(new_n11105_), .ZN(new_n11110_));
  NAND3_X1   g10090(.A1(new_n11110_), .A2(new_n11101_), .A3(new_n11102_), .ZN(new_n11111_));
  AOI21_X1   g10091(.A1(new_n11084_), .A2(new_n11083_), .B(new_n11082_), .ZN(new_n11112_));
  NOR3_X1    g10092(.A1(new_n11079_), .A2(new_n11080_), .A3(new_n11072_), .ZN(new_n11113_));
  NOR2_X1    g10093(.A1(new_n11112_), .A2(new_n11113_), .ZN(new_n11114_));
  NOR2_X1    g10094(.A1(new_n11095_), .A2(new_n11093_), .ZN(new_n11115_));
  NAND4_X1   g10095(.A1(new_n11115_), .A2(new_n11105_), .A3(new_n11088_), .A4(new_n11090_), .ZN(new_n11116_));
  NAND3_X1   g10096(.A1(new_n11111_), .A2(new_n11116_), .A3(new_n11114_), .ZN(new_n11117_));
  AOI22_X1   g10097(.A1(new_n11101_), .A2(new_n11102_), .B1(new_n11106_), .B2(new_n11105_), .ZN(new_n11118_));
  NOR3_X1    g10098(.A1(new_n11110_), .A2(new_n11028_), .A3(new_n11031_), .ZN(new_n11119_));
  OAI21_X1   g10099(.A1(new_n11119_), .A2(new_n11118_), .B(new_n11114_), .ZN(new_n11120_));
  NAND2_X1   g10100(.A1(new_n11011_), .A2(new_n11068_), .ZN(new_n11121_));
  NOR3_X1    g10101(.A1(new_n11074_), .A2(new_n11103_), .A3(new_n11077_), .ZN(new_n11122_));
  NAND2_X1   g10102(.A1(new_n11122_), .A2(new_n11121_), .ZN(new_n11123_));
  INV_X1     g10103(.I(new_n11121_), .ZN(new_n11124_));
  NAND3_X1   g10104(.A1(new_n11088_), .A2(new_n11054_), .A3(new_n11067_), .ZN(new_n11125_));
  NAND2_X1   g10105(.A1(new_n11125_), .A2(new_n11124_), .ZN(new_n11126_));
  INV_X1     g10106(.I(\A[976] ), .ZN(new_n11127_));
  NOR2_X1    g10107(.A1(\A[977] ), .A2(\A[978] ), .ZN(new_n11128_));
  NAND2_X1   g10108(.A1(\A[977] ), .A2(\A[978] ), .ZN(new_n11129_));
  AOI21_X1   g10109(.A1(new_n11127_), .A2(new_n11129_), .B(new_n11128_), .ZN(new_n11130_));
  INV_X1     g10110(.I(new_n11130_), .ZN(new_n11131_));
  INV_X1     g10111(.I(\A[973] ), .ZN(new_n11132_));
  NOR2_X1    g10112(.A1(\A[974] ), .A2(\A[975] ), .ZN(new_n11133_));
  NAND2_X1   g10113(.A1(\A[974] ), .A2(\A[975] ), .ZN(new_n11134_));
  AOI21_X1   g10114(.A1(new_n11132_), .A2(new_n11134_), .B(new_n11133_), .ZN(new_n11135_));
  INV_X1     g10115(.I(new_n11135_), .ZN(new_n11136_));
  NOR2_X1    g10116(.A1(new_n11131_), .A2(new_n11136_), .ZN(new_n11137_));
  INV_X1     g10117(.I(\A[975] ), .ZN(new_n11138_));
  NOR2_X1    g10118(.A1(new_n11138_), .A2(\A[974] ), .ZN(new_n11139_));
  INV_X1     g10119(.I(\A[974] ), .ZN(new_n11140_));
  NOR2_X1    g10120(.A1(new_n11140_), .A2(\A[975] ), .ZN(new_n11141_));
  OAI21_X1   g10121(.A1(new_n11139_), .A2(new_n11141_), .B(\A[973] ), .ZN(new_n11142_));
  INV_X1     g10122(.I(new_n11134_), .ZN(new_n11143_));
  OAI21_X1   g10123(.A1(new_n11143_), .A2(new_n11133_), .B(new_n11132_), .ZN(new_n11144_));
  NAND2_X1   g10124(.A1(new_n11142_), .A2(new_n11144_), .ZN(new_n11145_));
  INV_X1     g10125(.I(\A[978] ), .ZN(new_n11146_));
  NOR2_X1    g10126(.A1(new_n11146_), .A2(\A[977] ), .ZN(new_n11147_));
  INV_X1     g10127(.I(\A[977] ), .ZN(new_n11148_));
  NOR2_X1    g10128(.A1(new_n11148_), .A2(\A[978] ), .ZN(new_n11149_));
  OAI21_X1   g10129(.A1(new_n11147_), .A2(new_n11149_), .B(\A[976] ), .ZN(new_n11150_));
  INV_X1     g10130(.I(new_n11129_), .ZN(new_n11151_));
  OAI21_X1   g10131(.A1(new_n11151_), .A2(new_n11128_), .B(new_n11127_), .ZN(new_n11152_));
  NAND2_X1   g10132(.A1(new_n11150_), .A2(new_n11152_), .ZN(new_n11153_));
  NOR2_X1    g10133(.A1(new_n11145_), .A2(new_n11153_), .ZN(new_n11154_));
  NAND2_X1   g10134(.A1(new_n11154_), .A2(new_n11137_), .ZN(new_n11155_));
  NAND2_X1   g10135(.A1(new_n11140_), .A2(\A[975] ), .ZN(new_n11156_));
  NAND2_X1   g10136(.A1(new_n11138_), .A2(\A[974] ), .ZN(new_n11157_));
  AOI21_X1   g10137(.A1(new_n11156_), .A2(new_n11157_), .B(new_n11132_), .ZN(new_n11158_));
  INV_X1     g10138(.I(new_n11133_), .ZN(new_n11159_));
  AOI21_X1   g10139(.A1(new_n11159_), .A2(new_n11134_), .B(\A[973] ), .ZN(new_n11160_));
  NOR2_X1    g10140(.A1(new_n11160_), .A2(new_n11158_), .ZN(new_n11161_));
  NAND2_X1   g10141(.A1(new_n11148_), .A2(\A[978] ), .ZN(new_n11162_));
  NAND2_X1   g10142(.A1(new_n11146_), .A2(\A[977] ), .ZN(new_n11163_));
  AOI21_X1   g10143(.A1(new_n11162_), .A2(new_n11163_), .B(new_n11127_), .ZN(new_n11164_));
  INV_X1     g10144(.I(new_n11128_), .ZN(new_n11165_));
  AOI21_X1   g10145(.A1(new_n11165_), .A2(new_n11129_), .B(\A[976] ), .ZN(new_n11166_));
  NOR2_X1    g10146(.A1(new_n11166_), .A2(new_n11164_), .ZN(new_n11167_));
  NOR2_X1    g10147(.A1(new_n11161_), .A2(new_n11167_), .ZN(new_n11168_));
  NOR2_X1    g10148(.A1(new_n11168_), .A2(new_n11154_), .ZN(new_n11169_));
  INV_X1     g10149(.I(\A[967] ), .ZN(new_n11170_));
  INV_X1     g10150(.I(\A[968] ), .ZN(new_n11171_));
  NAND2_X1   g10151(.A1(new_n11171_), .A2(\A[969] ), .ZN(new_n11172_));
  INV_X1     g10152(.I(\A[969] ), .ZN(new_n11173_));
  NAND2_X1   g10153(.A1(new_n11173_), .A2(\A[968] ), .ZN(new_n11174_));
  AOI21_X1   g10154(.A1(new_n11172_), .A2(new_n11174_), .B(new_n11170_), .ZN(new_n11175_));
  NOR2_X1    g10155(.A1(\A[968] ), .A2(\A[969] ), .ZN(new_n11176_));
  INV_X1     g10156(.I(new_n11176_), .ZN(new_n11177_));
  NAND2_X1   g10157(.A1(\A[968] ), .A2(\A[969] ), .ZN(new_n11178_));
  AOI21_X1   g10158(.A1(new_n11177_), .A2(new_n11178_), .B(\A[967] ), .ZN(new_n11179_));
  NOR2_X1    g10159(.A1(new_n11179_), .A2(new_n11175_), .ZN(new_n11180_));
  INV_X1     g10160(.I(\A[970] ), .ZN(new_n11181_));
  INV_X1     g10161(.I(\A[971] ), .ZN(new_n11182_));
  NAND2_X1   g10162(.A1(new_n11182_), .A2(\A[972] ), .ZN(new_n11183_));
  INV_X1     g10163(.I(\A[972] ), .ZN(new_n11184_));
  NAND2_X1   g10164(.A1(new_n11184_), .A2(\A[971] ), .ZN(new_n11185_));
  AOI21_X1   g10165(.A1(new_n11183_), .A2(new_n11185_), .B(new_n11181_), .ZN(new_n11186_));
  NOR2_X1    g10166(.A1(\A[971] ), .A2(\A[972] ), .ZN(new_n11187_));
  INV_X1     g10167(.I(new_n11187_), .ZN(new_n11188_));
  NAND2_X1   g10168(.A1(\A[971] ), .A2(\A[972] ), .ZN(new_n11189_));
  AOI21_X1   g10169(.A1(new_n11188_), .A2(new_n11189_), .B(\A[970] ), .ZN(new_n11190_));
  NOR2_X1    g10170(.A1(new_n11190_), .A2(new_n11186_), .ZN(new_n11191_));
  AOI21_X1   g10171(.A1(new_n11181_), .A2(new_n11189_), .B(new_n11187_), .ZN(new_n11192_));
  INV_X1     g10172(.I(new_n11192_), .ZN(new_n11193_));
  AOI21_X1   g10173(.A1(new_n11170_), .A2(new_n11178_), .B(new_n11176_), .ZN(new_n11194_));
  INV_X1     g10174(.I(new_n11194_), .ZN(new_n11195_));
  NOR2_X1    g10175(.A1(new_n11193_), .A2(new_n11195_), .ZN(new_n11196_));
  NAND2_X1   g10176(.A1(new_n11169_), .A2(new_n11155_), .ZN(new_n11197_));
  AOI21_X1   g10177(.A1(new_n11126_), .A2(new_n11123_), .B(new_n11197_), .ZN(new_n11198_));
  AOI21_X1   g10178(.A1(new_n11120_), .A2(new_n11117_), .B(new_n11198_), .ZN(new_n11199_));
  INV_X1     g10179(.I(new_n11198_), .ZN(new_n11200_));
  NOR3_X1    g10180(.A1(new_n11097_), .A2(new_n11200_), .A3(new_n11108_), .ZN(new_n11201_));
  NAND2_X1   g10181(.A1(new_n11180_), .A2(new_n11191_), .ZN(new_n11202_));
  NAND2_X1   g10182(.A1(new_n11202_), .A2(new_n11194_), .ZN(new_n11203_));
  NAND3_X1   g10183(.A1(new_n11180_), .A2(new_n11191_), .A3(new_n11195_), .ZN(new_n11204_));
  AOI21_X1   g10184(.A1(new_n11203_), .A2(new_n11204_), .B(new_n11193_), .ZN(new_n11205_));
  NOR2_X1    g10185(.A1(new_n11173_), .A2(\A[968] ), .ZN(new_n11206_));
  NOR2_X1    g10186(.A1(new_n11171_), .A2(\A[969] ), .ZN(new_n11207_));
  OAI21_X1   g10187(.A1(new_n11206_), .A2(new_n11207_), .B(\A[967] ), .ZN(new_n11208_));
  INV_X1     g10188(.I(new_n11178_), .ZN(new_n11209_));
  OAI21_X1   g10189(.A1(new_n11209_), .A2(new_n11176_), .B(new_n11170_), .ZN(new_n11210_));
  NAND2_X1   g10190(.A1(new_n11208_), .A2(new_n11210_), .ZN(new_n11211_));
  NOR2_X1    g10191(.A1(new_n11184_), .A2(\A[971] ), .ZN(new_n11212_));
  NOR2_X1    g10192(.A1(new_n11182_), .A2(\A[972] ), .ZN(new_n11213_));
  OAI21_X1   g10193(.A1(new_n11212_), .A2(new_n11213_), .B(\A[970] ), .ZN(new_n11214_));
  INV_X1     g10194(.I(new_n11189_), .ZN(new_n11215_));
  OAI21_X1   g10195(.A1(new_n11215_), .A2(new_n11187_), .B(new_n11181_), .ZN(new_n11216_));
  NAND2_X1   g10196(.A1(new_n11214_), .A2(new_n11216_), .ZN(new_n11217_));
  NOR2_X1    g10197(.A1(new_n11211_), .A2(new_n11217_), .ZN(new_n11218_));
  NOR2_X1    g10198(.A1(new_n11218_), .A2(new_n11195_), .ZN(new_n11219_));
  INV_X1     g10199(.I(new_n11204_), .ZN(new_n11220_));
  NOR3_X1    g10200(.A1(new_n11219_), .A2(new_n11220_), .A3(new_n11192_), .ZN(new_n11221_));
  NOR2_X1    g10201(.A1(new_n11221_), .A2(new_n11205_), .ZN(new_n11222_));
  OR2_X2     g10202(.A1(new_n11168_), .A2(new_n11154_), .Z(new_n11223_));
  NAND2_X1   g10203(.A1(new_n11211_), .A2(new_n11217_), .ZN(new_n11224_));
  NAND2_X1   g10204(.A1(new_n11202_), .A2(new_n11224_), .ZN(new_n11225_));
  NOR2_X1    g10205(.A1(new_n11223_), .A2(new_n11225_), .ZN(new_n11226_));
  NAND2_X1   g10206(.A1(new_n11218_), .A2(new_n11196_), .ZN(new_n11227_));
  INV_X1     g10207(.I(new_n11137_), .ZN(new_n11228_));
  NOR2_X1    g10208(.A1(new_n11168_), .A2(new_n11228_), .ZN(new_n11229_));
  NAND2_X1   g10209(.A1(new_n11161_), .A2(new_n11167_), .ZN(new_n11230_));
  XNOR2_X1   g10210(.A1(new_n11130_), .A2(new_n11135_), .ZN(new_n11231_));
  NOR2_X1    g10211(.A1(new_n11230_), .A2(new_n11231_), .ZN(new_n11232_));
  NAND2_X1   g10212(.A1(new_n11131_), .A2(new_n11136_), .ZN(new_n11233_));
  AOI21_X1   g10213(.A1(new_n11228_), .A2(new_n11233_), .B(new_n11154_), .ZN(new_n11234_));
  NOR4_X1    g10214(.A1(new_n11234_), .A2(new_n11229_), .A3(new_n11232_), .A4(new_n11227_), .ZN(new_n11235_));
  NAND2_X1   g10215(.A1(new_n11235_), .A2(new_n11226_), .ZN(new_n11236_));
  NOR2_X1    g10216(.A1(new_n11236_), .A2(new_n11222_), .ZN(new_n11237_));
  OAI21_X1   g10217(.A1(new_n11219_), .A2(new_n11220_), .B(new_n11192_), .ZN(new_n11238_));
  NAND3_X1   g10218(.A1(new_n11203_), .A2(new_n11193_), .A3(new_n11204_), .ZN(new_n11239_));
  NAND2_X1   g10219(.A1(new_n11238_), .A2(new_n11239_), .ZN(new_n11240_));
  NOR2_X1    g10220(.A1(new_n11230_), .A2(new_n11228_), .ZN(new_n11241_));
  NOR4_X1    g10221(.A1(new_n11223_), .A2(new_n11225_), .A3(new_n11241_), .A4(new_n11227_), .ZN(new_n11242_));
  NAND2_X1   g10222(.A1(new_n11240_), .A2(new_n11242_), .ZN(new_n11243_));
  AOI21_X1   g10223(.A1(new_n11161_), .A2(new_n11167_), .B(new_n11136_), .ZN(new_n11244_));
  NOR3_X1    g10224(.A1(new_n11145_), .A2(new_n11153_), .A3(new_n11135_), .ZN(new_n11245_));
  OAI21_X1   g10225(.A1(new_n11244_), .A2(new_n11245_), .B(new_n11130_), .ZN(new_n11246_));
  INV_X1     g10226(.I(new_n11246_), .ZN(new_n11247_));
  NOR3_X1    g10227(.A1(new_n11244_), .A2(new_n11245_), .A3(new_n11130_), .ZN(new_n11248_));
  NOR2_X1    g10228(.A1(new_n11247_), .A2(new_n11248_), .ZN(new_n11249_));
  OAI21_X1   g10229(.A1(new_n11240_), .A2(new_n11242_), .B(new_n11249_), .ZN(new_n11250_));
  INV_X1     g10230(.I(new_n11196_), .ZN(new_n11251_));
  NOR2_X1    g10231(.A1(new_n11202_), .A2(new_n11251_), .ZN(new_n11252_));
  NOR2_X1    g10232(.A1(new_n11180_), .A2(new_n11191_), .ZN(new_n11253_));
  NOR2_X1    g10233(.A1(new_n11253_), .A2(new_n11218_), .ZN(new_n11254_));
  NAND4_X1   g10234(.A1(new_n11169_), .A2(new_n11254_), .A3(new_n11252_), .A4(new_n11155_), .ZN(new_n11255_));
  INV_X1     g10235(.I(new_n11248_), .ZN(new_n11256_));
  NAND2_X1   g10236(.A1(new_n11256_), .A2(new_n11246_), .ZN(new_n11257_));
  NAND3_X1   g10237(.A1(new_n11222_), .A2(new_n11257_), .A3(new_n11255_), .ZN(new_n11258_));
  NAND2_X1   g10238(.A1(new_n11250_), .A2(new_n11258_), .ZN(new_n11259_));
  AOI21_X1   g10239(.A1(new_n11259_), .A2(new_n11243_), .B(new_n11237_), .ZN(new_n11260_));
  OAI22_X1   g10240(.A1(new_n11260_), .A2(new_n11109_), .B1(new_n11199_), .B2(new_n11201_), .ZN(new_n11261_));
  AOI21_X1   g10241(.A1(new_n11026_), .A2(new_n11094_), .B(new_n11089_), .ZN(new_n11262_));
  INV_X1     g10242(.I(new_n11262_), .ZN(new_n11263_));
  OAI21_X1   g10243(.A1(new_n11072_), .A2(new_n11073_), .B(new_n11077_), .ZN(new_n11264_));
  NAND2_X1   g10244(.A1(new_n11264_), .A2(new_n11087_), .ZN(new_n11265_));
  INV_X1     g10245(.I(new_n11265_), .ZN(new_n11266_));
  NAND2_X1   g10246(.A1(new_n11101_), .A2(new_n11102_), .ZN(new_n11267_));
  OAI21_X1   g10247(.A1(new_n11267_), .A2(new_n11075_), .B(new_n11086_), .ZN(new_n11268_));
  AOI21_X1   g10248(.A1(new_n11268_), .A2(new_n11116_), .B(new_n11266_), .ZN(new_n11269_));
  NOR2_X1    g10249(.A1(new_n11076_), .A2(new_n11114_), .ZN(new_n11270_));
  NOR3_X1    g10250(.A1(new_n11270_), .A2(new_n11096_), .A3(new_n11265_), .ZN(new_n11271_));
  OAI21_X1   g10251(.A1(new_n11271_), .A2(new_n11269_), .B(new_n11263_), .ZN(new_n11272_));
  OAI21_X1   g10252(.A1(new_n11270_), .A2(new_n11096_), .B(new_n11265_), .ZN(new_n11273_));
  NAND3_X1   g10253(.A1(new_n11268_), .A2(new_n11116_), .A3(new_n11266_), .ZN(new_n11274_));
  NAND3_X1   g10254(.A1(new_n11273_), .A2(new_n11274_), .A3(new_n11262_), .ZN(new_n11275_));
  NAND2_X1   g10255(.A1(new_n11272_), .A2(new_n11275_), .ZN(new_n11276_));
  AOI21_X1   g10256(.A1(new_n11154_), .A2(new_n11233_), .B(new_n11137_), .ZN(new_n11277_));
  INV_X1     g10257(.I(new_n11236_), .ZN(new_n11278_));
  OAI21_X1   g10258(.A1(new_n11192_), .A2(new_n11194_), .B(new_n11218_), .ZN(new_n11279_));
  NAND2_X1   g10259(.A1(new_n11279_), .A2(new_n11251_), .ZN(new_n11280_));
  AOI21_X1   g10260(.A1(new_n11255_), .A2(new_n11249_), .B(new_n11222_), .ZN(new_n11281_));
  OAI21_X1   g10261(.A1(new_n11281_), .A2(new_n11278_), .B(new_n11280_), .ZN(new_n11282_));
  INV_X1     g10262(.I(new_n11280_), .ZN(new_n11283_));
  OAI21_X1   g10263(.A1(new_n11242_), .A2(new_n11257_), .B(new_n11240_), .ZN(new_n11284_));
  NAND3_X1   g10264(.A1(new_n11284_), .A2(new_n11236_), .A3(new_n11283_), .ZN(new_n11285_));
  AOI21_X1   g10265(.A1(new_n11282_), .A2(new_n11285_), .B(new_n11277_), .ZN(new_n11286_));
  INV_X1     g10266(.I(new_n11277_), .ZN(new_n11287_));
  AOI21_X1   g10267(.A1(new_n11284_), .A2(new_n11236_), .B(new_n11283_), .ZN(new_n11288_));
  NOR3_X1    g10268(.A1(new_n11281_), .A2(new_n11278_), .A3(new_n11280_), .ZN(new_n11289_));
  NOR3_X1    g10269(.A1(new_n11289_), .A2(new_n11288_), .A3(new_n11287_), .ZN(new_n11290_));
  NOR2_X1    g10270(.A1(new_n11286_), .A2(new_n11290_), .ZN(new_n11291_));
  XOR2_X1    g10271(.A1(new_n11276_), .A2(new_n11291_), .Z(new_n11292_));
  NOR2_X1    g10272(.A1(new_n11292_), .A2(new_n11261_), .ZN(new_n11293_));
  OAI21_X1   g10273(.A1(new_n11289_), .A2(new_n11288_), .B(new_n11287_), .ZN(new_n11294_));
  NAND3_X1   g10274(.A1(new_n11282_), .A2(new_n11285_), .A3(new_n11277_), .ZN(new_n11295_));
  NAND2_X1   g10275(.A1(new_n11294_), .A2(new_n11295_), .ZN(new_n11296_));
  NOR2_X1    g10276(.A1(new_n11276_), .A2(new_n11296_), .ZN(new_n11297_));
  AOI21_X1   g10277(.A1(new_n11273_), .A2(new_n11274_), .B(new_n11262_), .ZN(new_n11298_));
  NOR3_X1    g10278(.A1(new_n11271_), .A2(new_n11269_), .A3(new_n11263_), .ZN(new_n11299_));
  NOR2_X1    g10279(.A1(new_n11299_), .A2(new_n11298_), .ZN(new_n11300_));
  NOR2_X1    g10280(.A1(new_n11300_), .A2(new_n11291_), .ZN(new_n11301_));
  OAI21_X1   g10281(.A1(new_n11301_), .A2(new_n11297_), .B(new_n11261_), .ZN(new_n11302_));
  INV_X1     g10282(.I(new_n11302_), .ZN(new_n11303_));
  NOR4_X1    g10283(.A1(new_n11293_), .A2(new_n10973_), .A3(new_n11303_), .A4(new_n10985_), .ZN(new_n11304_));
  NAND2_X1   g10284(.A1(new_n10958_), .A2(new_n10960_), .ZN(new_n11305_));
  OAI21_X1   g10285(.A1(new_n10958_), .A2(new_n10960_), .B(new_n10956_), .ZN(new_n11306_));
  NAND2_X1   g10286(.A1(new_n11306_), .A2(new_n11305_), .ZN(new_n11307_));
  NAND2_X1   g10287(.A1(new_n10966_), .A2(new_n10968_), .ZN(new_n11308_));
  OR2_X2     g10288(.A1(new_n10966_), .A2(new_n10968_), .Z(new_n11309_));
  NAND3_X1   g10289(.A1(new_n10964_), .A2(new_n10963_), .A3(new_n11309_), .ZN(new_n11310_));
  NAND2_X1   g10290(.A1(new_n11310_), .A2(new_n11308_), .ZN(new_n11311_));
  INV_X1     g10291(.I(new_n11311_), .ZN(new_n11312_));
  NAND2_X1   g10292(.A1(new_n10955_), .A2(new_n10982_), .ZN(new_n11313_));
  AOI21_X1   g10293(.A1(new_n11313_), .A2(new_n10983_), .B(new_n11312_), .ZN(new_n11314_));
  NOR4_X1    g10294(.A1(new_n10955_), .A2(new_n10962_), .A3(new_n10970_), .A4(new_n11311_), .ZN(new_n11315_));
  OAI21_X1   g10295(.A1(new_n11314_), .A2(new_n11315_), .B(new_n11307_), .ZN(new_n11316_));
  INV_X1     g10296(.I(new_n11307_), .ZN(new_n11317_));
  INV_X1     g10297(.I(new_n10962_), .ZN(new_n11318_));
  NAND3_X1   g10298(.A1(new_n10981_), .A2(new_n11318_), .A3(new_n10971_), .ZN(new_n11319_));
  NAND2_X1   g10299(.A1(new_n11319_), .A2(new_n11311_), .ZN(new_n11320_));
  NAND4_X1   g10300(.A1(new_n10981_), .A2(new_n11312_), .A3(new_n11318_), .A4(new_n10971_), .ZN(new_n11321_));
  NAND3_X1   g10301(.A1(new_n11320_), .A2(new_n11317_), .A3(new_n11321_), .ZN(new_n11322_));
  NAND2_X1   g10302(.A1(new_n11316_), .A2(new_n11322_), .ZN(new_n11323_));
  NAND2_X1   g10303(.A1(new_n11268_), .A2(new_n11116_), .ZN(new_n11324_));
  NAND2_X1   g10304(.A1(new_n11265_), .A2(new_n11263_), .ZN(new_n11325_));
  NOR2_X1    g10305(.A1(new_n11265_), .A2(new_n11263_), .ZN(new_n11326_));
  OAI21_X1   g10306(.A1(new_n11324_), .A2(new_n11326_), .B(new_n11325_), .ZN(new_n11327_));
  NAND2_X1   g10307(.A1(new_n11284_), .A2(new_n11236_), .ZN(new_n11328_));
  NOR2_X1    g10308(.A1(new_n11280_), .A2(new_n11287_), .ZN(new_n11329_));
  NOR2_X1    g10309(.A1(new_n11328_), .A2(new_n11329_), .ZN(new_n11330_));
  AOI21_X1   g10310(.A1(new_n11287_), .A2(new_n11280_), .B(new_n11330_), .ZN(new_n11331_));
  OAI21_X1   g10311(.A1(new_n11276_), .A2(new_n11296_), .B(new_n11261_), .ZN(new_n11332_));
  XOR2_X1    g10312(.A1(new_n11265_), .A2(new_n11263_), .Z(new_n11333_));
  XOR2_X1    g10313(.A1(new_n11280_), .A2(new_n11287_), .Z(new_n11334_));
  NOR4_X1    g10314(.A1(new_n11324_), .A2(new_n11328_), .A3(new_n11333_), .A4(new_n11334_), .ZN(new_n11335_));
  AOI21_X1   g10315(.A1(new_n11332_), .A2(new_n11335_), .B(new_n11331_), .ZN(new_n11336_));
  INV_X1     g10316(.I(new_n11331_), .ZN(new_n11337_));
  NAND2_X1   g10317(.A1(new_n11120_), .A2(new_n11117_), .ZN(new_n11338_));
  OAI21_X1   g10318(.A1(new_n11097_), .A2(new_n11108_), .B(new_n11200_), .ZN(new_n11339_));
  NAND3_X1   g10319(.A1(new_n11120_), .A2(new_n11117_), .A3(new_n11198_), .ZN(new_n11340_));
  INV_X1     g10320(.I(new_n11237_), .ZN(new_n11341_));
  AOI21_X1   g10321(.A1(new_n11222_), .A2(new_n11255_), .B(new_n11257_), .ZN(new_n11342_));
  NOR3_X1    g10322(.A1(new_n11240_), .A2(new_n11249_), .A3(new_n11242_), .ZN(new_n11343_));
  OAI21_X1   g10323(.A1(new_n11342_), .A2(new_n11343_), .B(new_n11243_), .ZN(new_n11344_));
  NAND2_X1   g10324(.A1(new_n11344_), .A2(new_n11341_), .ZN(new_n11345_));
  AOI22_X1   g10325(.A1(new_n11345_), .A2(new_n11338_), .B1(new_n11340_), .B2(new_n11339_), .ZN(new_n11346_));
  AOI21_X1   g10326(.A1(new_n11300_), .A2(new_n11291_), .B(new_n11346_), .ZN(new_n11347_));
  INV_X1     g10327(.I(new_n11335_), .ZN(new_n11348_));
  NOR3_X1    g10328(.A1(new_n11347_), .A2(new_n11337_), .A3(new_n11348_), .ZN(new_n11349_));
  OAI21_X1   g10329(.A1(new_n11349_), .A2(new_n11336_), .B(new_n11327_), .ZN(new_n11350_));
  INV_X1     g10330(.I(new_n11327_), .ZN(new_n11351_));
  OAI21_X1   g10331(.A1(new_n11347_), .A2(new_n11348_), .B(new_n11337_), .ZN(new_n11352_));
  NAND3_X1   g10332(.A1(new_n11332_), .A2(new_n11331_), .A3(new_n11335_), .ZN(new_n11353_));
  NAND3_X1   g10333(.A1(new_n11352_), .A2(new_n11353_), .A3(new_n11351_), .ZN(new_n11354_));
  NAND2_X1   g10334(.A1(new_n11350_), .A2(new_n11354_), .ZN(new_n11355_));
  NOR2_X1    g10335(.A1(new_n11355_), .A2(new_n11323_), .ZN(new_n11356_));
  NOR2_X1    g10336(.A1(new_n11356_), .A2(new_n11304_), .ZN(new_n11357_));
  INV_X1     g10337(.I(new_n11319_), .ZN(new_n11358_));
  NOR2_X1    g10338(.A1(new_n11347_), .A2(new_n11348_), .ZN(new_n11359_));
  XOR2_X1    g10339(.A1(new_n11307_), .A2(new_n11312_), .Z(new_n11360_));
  XOR2_X1    g10340(.A1(new_n11331_), .A2(new_n11327_), .Z(new_n11361_));
  NAND4_X1   g10341(.A1(new_n11360_), .A2(new_n11359_), .A3(new_n11361_), .A4(new_n11358_), .ZN(new_n11362_));
  NOR2_X1    g10342(.A1(new_n11357_), .A2(new_n11362_), .ZN(new_n11363_));
  AOI21_X1   g10343(.A1(new_n11351_), .A2(new_n11331_), .B(new_n11359_), .ZN(new_n11364_));
  NOR2_X1    g10344(.A1(new_n11331_), .A2(new_n11351_), .ZN(new_n11365_));
  NOR2_X1    g10345(.A1(new_n11364_), .A2(new_n11365_), .ZN(new_n11366_));
  NOR4_X1    g10346(.A1(new_n11366_), .A2(new_n11317_), .A3(new_n11312_), .A4(new_n11319_), .ZN(new_n11367_));
  NOR2_X1    g10347(.A1(new_n11307_), .A2(new_n11311_), .ZN(new_n11368_));
  AOI21_X1   g10348(.A1(new_n11307_), .A2(new_n11311_), .B(new_n11319_), .ZN(new_n11369_));
  NOR2_X1    g10349(.A1(new_n11369_), .A2(new_n11368_), .ZN(new_n11370_));
  INV_X1     g10350(.I(new_n11370_), .ZN(new_n11371_));
  OAI22_X1   g10351(.A1(new_n11363_), .A2(new_n11367_), .B1(new_n11366_), .B2(new_n11371_), .ZN(new_n11372_));
  INV_X1     g10352(.I(new_n11372_), .ZN(new_n11373_));
  NOR2_X1    g10353(.A1(new_n10661_), .A2(new_n10610_), .ZN(new_n11374_));
  INV_X1     g10354(.I(new_n10687_), .ZN(new_n11375_));
  NOR2_X1    g10355(.A1(new_n11375_), .A2(new_n10688_), .ZN(new_n11376_));
  INV_X1     g10356(.I(new_n10685_), .ZN(new_n11377_));
  AOI21_X1   g10357(.A1(new_n10679_), .A2(new_n10683_), .B(new_n11377_), .ZN(new_n11378_));
  NOR2_X1    g10358(.A1(new_n11378_), .A2(new_n10687_), .ZN(new_n11379_));
  NOR2_X1    g10359(.A1(new_n11376_), .A2(new_n11379_), .ZN(new_n11380_));
  OAI21_X1   g10360(.A1(new_n11374_), .A2(new_n10674_), .B(new_n11380_), .ZN(new_n11381_));
  OR2_X2     g10361(.A1(new_n11381_), .A2(new_n11373_), .Z(new_n11382_));
  NAND2_X1   g10362(.A1(new_n10675_), .A2(new_n10688_), .ZN(new_n11383_));
  NAND3_X1   g10363(.A1(new_n10067_), .A2(new_n10035_), .A3(new_n10038_), .ZN(new_n11384_));
  NAND2_X1   g10364(.A1(new_n10039_), .A2(new_n10063_), .ZN(new_n11385_));
  AOI21_X1   g10365(.A1(new_n11385_), .A2(new_n11384_), .B(new_n10077_), .ZN(new_n11386_));
  OAI22_X1   g10366(.A1(new_n10079_), .A2(new_n10078_), .B1(new_n10058_), .B2(new_n10062_), .ZN(new_n11387_));
  AOI21_X1   g10367(.A1(new_n10628_), .A2(new_n11387_), .B(new_n10015_), .ZN(new_n11388_));
  OAI21_X1   g10368(.A1(new_n10539_), .A2(new_n10538_), .B(new_n10537_), .ZN(new_n11389_));
  NAND3_X1   g10369(.A1(new_n10530_), .A2(new_n10533_), .A3(new_n10505_), .ZN(new_n11390_));
  AOI21_X1   g10370(.A1(new_n11389_), .A2(new_n11390_), .B(new_n10545_), .ZN(new_n11391_));
  AOI21_X1   g10371(.A1(new_n10666_), .A2(new_n10665_), .B(new_n10496_), .ZN(new_n11392_));
  NOR4_X1    g10372(.A1(new_n11386_), .A2(new_n11388_), .A3(new_n11391_), .A4(new_n11392_), .ZN(new_n11393_));
  NOR2_X1    g10373(.A1(new_n10013_), .A2(new_n10074_), .ZN(new_n11394_));
  NOR2_X1    g10374(.A1(new_n10075_), .A2(new_n10006_), .ZN(new_n11395_));
  OAI21_X1   g10375(.A1(new_n11395_), .A2(new_n11394_), .B(new_n10073_), .ZN(new_n11396_));
  OAI21_X1   g10376(.A1(new_n10014_), .A2(new_n10070_), .B(new_n10003_), .ZN(new_n11397_));
  AOI21_X1   g10377(.A1(new_n10559_), .A2(new_n10560_), .B(new_n10558_), .ZN(new_n11398_));
  NOR3_X1    g10378(.A1(new_n10556_), .A2(new_n10555_), .A3(new_n10554_), .ZN(new_n11399_));
  NOR2_X1    g10379(.A1(new_n11399_), .A2(new_n11398_), .ZN(new_n11400_));
  NAND3_X1   g10380(.A1(new_n11396_), .A2(new_n11397_), .A3(new_n11400_), .ZN(new_n11401_));
  INV_X1     g10381(.I(new_n10606_), .ZN(new_n11402_));
  AOI21_X1   g10382(.A1(new_n11396_), .A2(new_n11397_), .B(new_n11400_), .ZN(new_n11403_));
  OAI21_X1   g10383(.A1(new_n11402_), .A2(new_n11403_), .B(new_n11401_), .ZN(new_n11404_));
  OAI22_X1   g10384(.A1(new_n11386_), .A2(new_n11388_), .B1(new_n11391_), .B2(new_n11392_), .ZN(new_n11405_));
  AOI21_X1   g10385(.A1(new_n11404_), .A2(new_n11405_), .B(new_n11393_), .ZN(new_n11406_));
  OAI21_X1   g10386(.A1(new_n10634_), .A2(new_n10633_), .B(new_n10616_), .ZN(new_n11407_));
  NAND3_X1   g10387(.A1(new_n10626_), .A2(new_n10631_), .A3(new_n10617_), .ZN(new_n11408_));
  NAND2_X1   g10388(.A1(new_n10649_), .A2(new_n10642_), .ZN(new_n11409_));
  AOI21_X1   g10389(.A1(new_n10515_), .A2(new_n10518_), .B(new_n10510_), .ZN(new_n11410_));
  INV_X1     g10390(.I(new_n10651_), .ZN(new_n11411_));
  OAI21_X1   g10391(.A1(new_n11411_), .A2(new_n11410_), .B(new_n10514_), .ZN(new_n11412_));
  NAND2_X1   g10392(.A1(new_n11412_), .A2(new_n11409_), .ZN(new_n11413_));
  NAND2_X1   g10393(.A1(new_n11413_), .A2(new_n10653_), .ZN(new_n11414_));
  NAND3_X1   g10394(.A1(new_n11414_), .A2(new_n10667_), .A3(new_n10665_), .ZN(new_n11415_));
  AOI22_X1   g10395(.A1(new_n10545_), .A2(new_n10505_), .B1(new_n10530_), .B2(new_n10533_), .ZN(new_n11416_));
  NOR2_X1    g10396(.A1(new_n11414_), .A2(new_n11416_), .ZN(new_n11417_));
  NAND2_X1   g10397(.A1(new_n11417_), .A2(new_n11415_), .ZN(new_n11418_));
  NAND3_X1   g10398(.A1(new_n11418_), .A2(new_n11407_), .A3(new_n11408_), .ZN(new_n11419_));
  NAND2_X1   g10399(.A1(new_n11419_), .A2(new_n11406_), .ZN(new_n11420_));
  NAND3_X1   g10400(.A1(new_n11420_), .A2(new_n10674_), .A3(new_n11378_), .ZN(new_n11421_));
  AOI21_X1   g10401(.A1(new_n11383_), .A2(new_n11421_), .B(new_n11375_), .ZN(new_n11422_));
  AOI21_X1   g10402(.A1(new_n11420_), .A2(new_n10674_), .B(new_n11378_), .ZN(new_n11423_));
  NOR2_X1    g10403(.A1(new_n10675_), .A2(new_n10688_), .ZN(new_n11424_));
  NOR3_X1    g10404(.A1(new_n11424_), .A2(new_n11423_), .A3(new_n10687_), .ZN(new_n11425_));
  NOR2_X1    g10405(.A1(new_n11425_), .A2(new_n11422_), .ZN(new_n11426_));
  NAND3_X1   g10406(.A1(new_n11426_), .A2(new_n11373_), .A3(new_n11382_), .ZN(new_n11427_));
  INV_X1     g10407(.I(new_n11427_), .ZN(new_n11428_));
  NAND2_X1   g10408(.A1(new_n7787_), .A2(new_n7791_), .ZN(new_n11429_));
  NAND3_X1   g10409(.A1(new_n11429_), .A2(new_n7787_), .A3(new_n7791_), .ZN(new_n11430_));
  XOR2_X1    g10410(.A1(new_n11427_), .A2(new_n10689_), .Z(new_n11431_));
  XNOR2_X1   g10411(.A1(new_n11431_), .A2(new_n9309_), .ZN(new_n11432_));
  OAI21_X1   g10412(.A1(new_n10609_), .A2(new_n11393_), .B(new_n10608_), .ZN(new_n11433_));
  NAND3_X1   g10413(.A1(new_n10549_), .A2(new_n11405_), .A3(new_n11404_), .ZN(new_n11434_));
  AOI21_X1   g10414(.A1(new_n11320_), .A2(new_n11321_), .B(new_n11317_), .ZN(new_n11435_));
  NOR3_X1    g10415(.A1(new_n11314_), .A2(new_n11307_), .A3(new_n11315_), .ZN(new_n11436_));
  NOR2_X1    g10416(.A1(new_n11436_), .A2(new_n11435_), .ZN(new_n11437_));
  NOR2_X1    g10417(.A1(new_n11355_), .A2(new_n11437_), .ZN(new_n11438_));
  AOI21_X1   g10418(.A1(new_n11352_), .A2(new_n11353_), .B(new_n11351_), .ZN(new_n11439_));
  NOR3_X1    g10419(.A1(new_n11349_), .A2(new_n11336_), .A3(new_n11327_), .ZN(new_n11440_));
  NOR2_X1    g10420(.A1(new_n11440_), .A2(new_n11439_), .ZN(new_n11441_));
  NOR2_X1    g10421(.A1(new_n11441_), .A2(new_n11323_), .ZN(new_n11442_));
  OAI21_X1   g10422(.A1(new_n11442_), .A2(new_n11438_), .B(new_n11304_), .ZN(new_n11443_));
  XOR2_X1    g10423(.A1(new_n10962_), .A2(new_n10970_), .Z(new_n11444_));
  AOI21_X1   g10424(.A1(new_n10981_), .A2(new_n11444_), .B(new_n10985_), .ZN(new_n11445_));
  NOR2_X1    g10425(.A1(new_n11293_), .A2(new_n11303_), .ZN(new_n11446_));
  NAND2_X1   g10426(.A1(new_n11446_), .A2(new_n11445_), .ZN(new_n11447_));
  AOI22_X1   g10427(.A1(new_n11350_), .A2(new_n11354_), .B1(new_n11316_), .B2(new_n11322_), .ZN(new_n11448_));
  OAI21_X1   g10428(.A1(new_n11356_), .A2(new_n11448_), .B(new_n11447_), .ZN(new_n11449_));
  NAND2_X1   g10429(.A1(new_n11443_), .A2(new_n11449_), .ZN(new_n11450_));
  AOI21_X1   g10430(.A1(new_n11433_), .A2(new_n11434_), .B(new_n11450_), .ZN(new_n11451_));
  NAND3_X1   g10431(.A1(new_n11433_), .A2(new_n11434_), .A3(new_n11450_), .ZN(new_n11452_));
  INV_X1     g10432(.I(new_n11452_), .ZN(new_n11453_));
  NAND3_X1   g10433(.A1(new_n11433_), .A2(new_n11434_), .A3(new_n11450_), .ZN(new_n11454_));
  INV_X1     g10434(.I(new_n11454_), .ZN(new_n11455_));
  NOR3_X1    g10435(.A1(new_n11453_), .A2(new_n11455_), .A3(new_n11451_), .ZN(new_n11456_));
  AOI21_X1   g10436(.A1(new_n11407_), .A2(new_n11408_), .B(new_n10660_), .ZN(new_n11457_));
  NOR3_X1    g10437(.A1(new_n11418_), .A2(new_n10632_), .A3(new_n10635_), .ZN(new_n11458_));
  OAI21_X1   g10438(.A1(new_n11457_), .A2(new_n11458_), .B(new_n11406_), .ZN(new_n11459_));
  AOI21_X1   g10439(.A1(new_n11407_), .A2(new_n11408_), .B(new_n11418_), .ZN(new_n11460_));
  OAI21_X1   g10440(.A1(new_n11460_), .A2(new_n10661_), .B(new_n10610_), .ZN(new_n11461_));
  INV_X1     g10441(.I(new_n11366_), .ZN(new_n11462_));
  OAI21_X1   g10442(.A1(new_n11357_), .A2(new_n11362_), .B(new_n11370_), .ZN(new_n11463_));
  INV_X1     g10443(.I(new_n11463_), .ZN(new_n11464_));
  NOR3_X1    g10444(.A1(new_n11357_), .A2(new_n11362_), .A3(new_n11370_), .ZN(new_n11465_));
  OAI21_X1   g10445(.A1(new_n11464_), .A2(new_n11465_), .B(new_n11462_), .ZN(new_n11466_));
  NAND2_X1   g10446(.A1(new_n11363_), .A2(new_n11371_), .ZN(new_n11467_));
  NAND3_X1   g10447(.A1(new_n11467_), .A2(new_n11366_), .A3(new_n11463_), .ZN(new_n11468_));
  NAND2_X1   g10448(.A1(new_n11466_), .A2(new_n11468_), .ZN(new_n11469_));
  AOI21_X1   g10449(.A1(new_n11459_), .A2(new_n11461_), .B(new_n11469_), .ZN(new_n11470_));
  OAI21_X1   g10450(.A1(new_n10632_), .A2(new_n10635_), .B(new_n11418_), .ZN(new_n11471_));
  NAND3_X1   g10451(.A1(new_n10660_), .A2(new_n11407_), .A3(new_n11408_), .ZN(new_n11472_));
  AOI21_X1   g10452(.A1(new_n11471_), .A2(new_n11472_), .B(new_n10610_), .ZN(new_n11473_));
  OAI21_X1   g10453(.A1(new_n10632_), .A2(new_n10635_), .B(new_n10660_), .ZN(new_n11474_));
  AOI21_X1   g10454(.A1(new_n11474_), .A2(new_n11419_), .B(new_n11406_), .ZN(new_n11475_));
  AOI21_X1   g10455(.A1(new_n11467_), .A2(new_n11463_), .B(new_n11366_), .ZN(new_n11476_));
  NOR3_X1    g10456(.A1(new_n11464_), .A2(new_n11462_), .A3(new_n11465_), .ZN(new_n11477_));
  NOR2_X1    g10457(.A1(new_n11477_), .A2(new_n11476_), .ZN(new_n11478_));
  NOR3_X1    g10458(.A1(new_n11475_), .A2(new_n11478_), .A3(new_n11473_), .ZN(new_n11479_));
  OAI21_X1   g10459(.A1(new_n11470_), .A2(new_n11479_), .B(new_n11456_), .ZN(new_n11480_));
  INV_X1     g10460(.I(new_n11433_), .ZN(new_n11481_));
  NOR3_X1    g10461(.A1(new_n10609_), .A2(new_n11393_), .A3(new_n10608_), .ZN(new_n11482_));
  NAND2_X1   g10462(.A1(new_n11441_), .A2(new_n11323_), .ZN(new_n11483_));
  NAND2_X1   g10463(.A1(new_n11355_), .A2(new_n11437_), .ZN(new_n11484_));
  AOI21_X1   g10464(.A1(new_n11483_), .A2(new_n11484_), .B(new_n11447_), .ZN(new_n11485_));
  NAND3_X1   g10465(.A1(new_n11437_), .A2(new_n11350_), .A3(new_n11354_), .ZN(new_n11486_));
  NAND2_X1   g10466(.A1(new_n11355_), .A2(new_n11323_), .ZN(new_n11487_));
  AOI21_X1   g10467(.A1(new_n11487_), .A2(new_n11486_), .B(new_n11304_), .ZN(new_n11488_));
  NOR2_X1    g10468(.A1(new_n11485_), .A2(new_n11488_), .ZN(new_n11489_));
  OAI21_X1   g10469(.A1(new_n11481_), .A2(new_n11482_), .B(new_n11489_), .ZN(new_n11490_));
  NAND3_X1   g10470(.A1(new_n11490_), .A2(new_n11452_), .A3(new_n11454_), .ZN(new_n11491_));
  OAI21_X1   g10471(.A1(new_n11475_), .A2(new_n11473_), .B(new_n11478_), .ZN(new_n11492_));
  NAND3_X1   g10472(.A1(new_n11459_), .A2(new_n11461_), .A3(new_n11469_), .ZN(new_n11493_));
  NAND3_X1   g10473(.A1(new_n11492_), .A2(new_n11493_), .A3(new_n11491_), .ZN(new_n11494_));
  NAND2_X1   g10474(.A1(new_n11480_), .A2(new_n11494_), .ZN(new_n11495_));
  AOI21_X1   g10475(.A1(new_n11492_), .A2(new_n11493_), .B(new_n11491_), .ZN(new_n11496_));
  NOR3_X1    g10476(.A1(new_n11456_), .A2(new_n11479_), .A3(new_n11470_), .ZN(new_n11497_));
  INV_X1     g10477(.I(new_n9239_), .ZN(new_n11498_));
  NAND2_X1   g10478(.A1(new_n9256_), .A2(new_n9262_), .ZN(new_n11499_));
  NAND2_X1   g10479(.A1(new_n9282_), .A2(new_n9285_), .ZN(new_n11500_));
  XOR2_X1    g10480(.A1(new_n11499_), .A2(new_n11500_), .Z(new_n11501_));
  AOI22_X1   g10481(.A1(new_n9256_), .A2(new_n9262_), .B1(new_n9282_), .B2(new_n9285_), .ZN(new_n11502_));
  INV_X1     g10482(.I(new_n11502_), .ZN(new_n11503_));
  AOI21_X1   g10483(.A1(new_n11503_), .A2(new_n9286_), .B(new_n11498_), .ZN(new_n11504_));
  AOI21_X1   g10484(.A1(new_n11501_), .A2(new_n11498_), .B(new_n11504_), .ZN(new_n11505_));
  OAI21_X1   g10485(.A1(new_n11497_), .A2(new_n11496_), .B(new_n11505_), .ZN(new_n11506_));
  XNOR2_X1   g10486(.A1(new_n11499_), .A2(new_n11500_), .ZN(new_n11507_));
  INV_X1     g10487(.I(new_n9286_), .ZN(new_n11508_));
  OAI21_X1   g10488(.A1(new_n11508_), .A2(new_n11502_), .B(new_n9239_), .ZN(new_n11509_));
  OAI21_X1   g10489(.A1(new_n11507_), .A2(new_n9239_), .B(new_n11509_), .ZN(new_n11510_));
  NAND3_X1   g10490(.A1(new_n11480_), .A2(new_n11494_), .A3(new_n11510_), .ZN(new_n11511_));
  NOR2_X1    g10491(.A1(new_n10609_), .A2(new_n11393_), .ZN(new_n11512_));
  NAND2_X1   g10492(.A1(new_n11450_), .A2(new_n10608_), .ZN(new_n11513_));
  NAND2_X1   g10493(.A1(new_n11489_), .A2(new_n11404_), .ZN(new_n11514_));
  AOI21_X1   g10494(.A1(new_n11514_), .A2(new_n11513_), .B(new_n11512_), .ZN(new_n11515_));
  NAND2_X1   g10495(.A1(new_n10549_), .A2(new_n11405_), .ZN(new_n11516_));
  NAND2_X1   g10496(.A1(new_n11450_), .A2(new_n11404_), .ZN(new_n11517_));
  NAND2_X1   g10497(.A1(new_n11489_), .A2(new_n10608_), .ZN(new_n11518_));
  AOI21_X1   g10498(.A1(new_n11518_), .A2(new_n11517_), .B(new_n11516_), .ZN(new_n11519_));
  NOR2_X1    g10499(.A1(new_n11515_), .A2(new_n11519_), .ZN(new_n11520_));
  INV_X1     g10500(.I(new_n11520_), .ZN(new_n11521_));
  NOR2_X1    g10501(.A1(new_n8484_), .A2(new_n8492_), .ZN(new_n11522_));
  AOI21_X1   g10502(.A1(new_n9158_), .A2(new_n9163_), .B(new_n9189_), .ZN(new_n11523_));
  NOR2_X1    g10503(.A1(new_n9164_), .A2(new_n9185_), .ZN(new_n11524_));
  OAI21_X1   g10504(.A1(new_n11523_), .A2(new_n11524_), .B(new_n9194_), .ZN(new_n11525_));
  AOI22_X1   g10505(.A1(new_n9158_), .A2(new_n9163_), .B1(new_n9187_), .B2(new_n9188_), .ZN(new_n11526_));
  OAI21_X1   g10506(.A1(new_n9277_), .A2(new_n11526_), .B(new_n9143_), .ZN(new_n11527_));
  NAND2_X1   g10507(.A1(new_n11525_), .A2(new_n11527_), .ZN(new_n11528_));
  NAND2_X1   g10508(.A1(new_n11522_), .A2(new_n11528_), .ZN(new_n11529_));
  NOR2_X1    g10509(.A1(new_n8479_), .A2(new_n8482_), .ZN(new_n11530_));
  NOR2_X1    g10510(.A1(new_n8454_), .A2(new_n8475_), .ZN(new_n11531_));
  OAI21_X1   g10511(.A1(new_n11531_), .A2(new_n11530_), .B(new_n8489_), .ZN(new_n11532_));
  AOI22_X1   g10512(.A1(new_n8449_), .A2(new_n8453_), .B1(new_n8480_), .B2(new_n8481_), .ZN(new_n11533_));
  OAI21_X1   g10513(.A1(new_n9257_), .A2(new_n11533_), .B(new_n8434_), .ZN(new_n11534_));
  NAND2_X1   g10514(.A1(new_n11532_), .A2(new_n11534_), .ZN(new_n11535_));
  NAND2_X1   g10515(.A1(new_n9186_), .A2(new_n9190_), .ZN(new_n11536_));
  AOI21_X1   g10516(.A1(new_n11536_), .A2(new_n9194_), .B(new_n9199_), .ZN(new_n11537_));
  NAND2_X1   g10517(.A1(new_n11535_), .A2(new_n11537_), .ZN(new_n11538_));
  NAND2_X1   g10518(.A1(new_n11529_), .A2(new_n11538_), .ZN(new_n11539_));
  NAND4_X1   g10519(.A1(new_n11532_), .A2(new_n11525_), .A3(new_n11534_), .A4(new_n11527_), .ZN(new_n11540_));
  AOI21_X1   g10520(.A1(new_n9238_), .A2(new_n11540_), .B(new_n9237_), .ZN(new_n11541_));
  AOI21_X1   g10521(.A1(new_n11539_), .A2(new_n9237_), .B(new_n11541_), .ZN(new_n11542_));
  OAI21_X1   g10522(.A1(new_n11515_), .A2(new_n11519_), .B(new_n11542_), .ZN(new_n11543_));
  NOR2_X1    g10523(.A1(new_n11489_), .A2(new_n11404_), .ZN(new_n11544_));
  NOR2_X1    g10524(.A1(new_n11450_), .A2(new_n10608_), .ZN(new_n11545_));
  OAI21_X1   g10525(.A1(new_n11544_), .A2(new_n11545_), .B(new_n11516_), .ZN(new_n11546_));
  NOR2_X1    g10526(.A1(new_n11489_), .A2(new_n10608_), .ZN(new_n11547_));
  NOR2_X1    g10527(.A1(new_n11450_), .A2(new_n11404_), .ZN(new_n11548_));
  OAI21_X1   g10528(.A1(new_n11547_), .A2(new_n11548_), .B(new_n11512_), .ZN(new_n11549_));
  NOR2_X1    g10529(.A1(new_n11535_), .A2(new_n11537_), .ZN(new_n11550_));
  NOR2_X1    g10530(.A1(new_n11522_), .A2(new_n11528_), .ZN(new_n11551_));
  OAI21_X1   g10531(.A1(new_n11551_), .A2(new_n11550_), .B(new_n9237_), .ZN(new_n11552_));
  NAND2_X1   g10532(.A1(new_n9203_), .A2(new_n9123_), .ZN(new_n11553_));
  NAND2_X1   g10533(.A1(new_n9201_), .A2(new_n8809_), .ZN(new_n11554_));
  AOI21_X1   g10534(.A1(new_n11554_), .A2(new_n11553_), .B(new_n9140_), .ZN(new_n11555_));
  AOI21_X1   g10535(.A1(new_n9142_), .A2(new_n9192_), .B(new_n9141_), .ZN(new_n11556_));
  NAND2_X1   g10536(.A1(new_n9215_), .A2(new_n9216_), .ZN(new_n11557_));
  NOR3_X1    g10537(.A1(new_n11557_), .A2(new_n11555_), .A3(new_n11556_), .ZN(new_n11558_));
  INV_X1     g10538(.I(new_n9234_), .ZN(new_n11559_));
  AOI22_X1   g10539(.A1(new_n11559_), .A2(new_n9219_), .B1(new_n9225_), .B2(new_n9227_), .ZN(new_n11560_));
  NAND2_X1   g10540(.A1(new_n9213_), .A2(new_n8416_), .ZN(new_n11561_));
  NAND2_X1   g10541(.A1(new_n9209_), .A2(new_n8105_), .ZN(new_n11562_));
  AOI21_X1   g10542(.A1(new_n11561_), .A2(new_n11562_), .B(new_n8488_), .ZN(new_n11563_));
  AOI21_X1   g10543(.A1(new_n8433_), .A2(new_n8485_), .B(new_n8431_), .ZN(new_n11564_));
  OAI22_X1   g10544(.A1(new_n11555_), .A2(new_n11556_), .B1(new_n11563_), .B2(new_n11564_), .ZN(new_n11565_));
  AOI21_X1   g10545(.A1(new_n11560_), .A2(new_n11565_), .B(new_n11558_), .ZN(new_n11566_));
  NOR2_X1    g10546(.A1(new_n11522_), .A2(new_n11537_), .ZN(new_n11567_));
  OAI21_X1   g10547(.A1(new_n11567_), .A2(new_n9200_), .B(new_n11566_), .ZN(new_n11568_));
  NAND2_X1   g10548(.A1(new_n11552_), .A2(new_n11568_), .ZN(new_n11569_));
  NAND3_X1   g10549(.A1(new_n11569_), .A2(new_n11549_), .A3(new_n11546_), .ZN(new_n11570_));
  NAND2_X1   g10550(.A1(new_n10585_), .A2(new_n10586_), .ZN(new_n11571_));
  NOR2_X1    g10551(.A1(new_n11571_), .A2(new_n10605_), .ZN(new_n11572_));
  NAND2_X1   g10552(.A1(new_n11169_), .A2(new_n11155_), .ZN(new_n11573_));
  XOR2_X1    g10553(.A1(new_n11573_), .A2(new_n11121_), .Z(new_n11574_));
  XOR2_X1    g10554(.A1(new_n11574_), .A2(new_n11122_), .Z(new_n11575_));
  NAND2_X1   g10555(.A1(new_n10824_), .A2(new_n10865_), .ZN(new_n11576_));
  NAND2_X1   g10556(.A1(new_n10898_), .A2(new_n11576_), .ZN(new_n11577_));
  NOR2_X1    g10557(.A1(new_n11575_), .A2(new_n11577_), .ZN(new_n11578_));
  INV_X1     g10558(.I(new_n11578_), .ZN(new_n11579_));
  NAND2_X1   g10559(.A1(new_n11575_), .A2(new_n11577_), .ZN(new_n11580_));
  NAND2_X1   g10560(.A1(new_n11579_), .A2(new_n11580_), .ZN(new_n11581_));
  INV_X1     g10561(.I(new_n11581_), .ZN(new_n11582_));
  NOR3_X1    g10562(.A1(new_n10583_), .A2(new_n10567_), .A3(new_n9994_), .ZN(new_n11583_));
  INV_X1     g10563(.I(new_n10583_), .ZN(new_n11584_));
  NOR2_X1    g10564(.A1(new_n11584_), .A2(new_n10568_), .ZN(new_n11585_));
  OAI21_X1   g10565(.A1(new_n11585_), .A2(new_n11583_), .B(new_n11582_), .ZN(new_n11586_));
  OAI21_X1   g10566(.A1(new_n11571_), .A2(new_n10605_), .B(new_n11586_), .ZN(new_n11587_));
  INV_X1     g10567(.I(new_n11587_), .ZN(new_n11588_));
  NOR3_X1    g10568(.A1(new_n11571_), .A2(new_n10605_), .A3(new_n11586_), .ZN(new_n11589_));
  NAND3_X1   g10569(.A1(new_n11260_), .A2(new_n11340_), .A3(new_n11339_), .ZN(new_n11590_));
  INV_X1     g10570(.I(new_n11590_), .ZN(new_n11591_));
  OAI21_X1   g10571(.A1(new_n10893_), .A2(new_n10899_), .B(new_n10954_), .ZN(new_n11592_));
  NAND3_X1   g10572(.A1(new_n10975_), .A2(new_n10980_), .A3(new_n10976_), .ZN(new_n11593_));
  NAND2_X1   g10573(.A1(new_n11592_), .A2(new_n11593_), .ZN(new_n11594_));
  NOR2_X1    g10574(.A1(new_n11594_), .A2(new_n11591_), .ZN(new_n11595_));
  INV_X1     g10575(.I(new_n11595_), .ZN(new_n11596_));
  NAND2_X1   g10576(.A1(new_n11594_), .A2(new_n11591_), .ZN(new_n11597_));
  AOI21_X1   g10577(.A1(new_n11596_), .A2(new_n11597_), .B(new_n11578_), .ZN(new_n11598_));
  AND3_X2    g10578(.A1(new_n11596_), .A2(new_n11578_), .A3(new_n11597_), .Z(new_n11599_));
  NOR2_X1    g10579(.A1(new_n11599_), .A2(new_n11598_), .ZN(new_n11600_));
  OAI22_X1   g10580(.A1(new_n11588_), .A2(new_n11589_), .B1(new_n11572_), .B2(new_n11600_), .ZN(new_n11601_));
  NOR3_X1    g10581(.A1(new_n10552_), .A2(new_n10553_), .A3(new_n11400_), .ZN(new_n11602_));
  AOI21_X1   g10582(.A1(new_n11396_), .A2(new_n11397_), .B(new_n10562_), .ZN(new_n11603_));
  OAI21_X1   g10583(.A1(new_n11603_), .A2(new_n11602_), .B(new_n11402_), .ZN(new_n11604_));
  OAI21_X1   g10584(.A1(new_n11403_), .A2(new_n10563_), .B(new_n10606_), .ZN(new_n11605_));
  XNOR2_X1   g10585(.A1(new_n11446_), .A2(new_n11445_), .ZN(new_n11606_));
  AOI21_X1   g10586(.A1(new_n11604_), .A2(new_n11605_), .B(new_n11606_), .ZN(new_n11607_));
  NAND3_X1   g10587(.A1(new_n11396_), .A2(new_n11397_), .A3(new_n10562_), .ZN(new_n11608_));
  OAI21_X1   g10588(.A1(new_n10552_), .A2(new_n10553_), .B(new_n11400_), .ZN(new_n11609_));
  AOI21_X1   g10589(.A1(new_n11608_), .A2(new_n11609_), .B(new_n10606_), .ZN(new_n11610_));
  AOI21_X1   g10590(.A1(new_n11401_), .A2(new_n10607_), .B(new_n11402_), .ZN(new_n11611_));
  NOR2_X1    g10591(.A1(new_n11446_), .A2(new_n11445_), .ZN(new_n11612_));
  NOR2_X1    g10592(.A1(new_n11612_), .A2(new_n11304_), .ZN(new_n11613_));
  NOR3_X1    g10593(.A1(new_n11610_), .A2(new_n11611_), .A3(new_n11613_), .ZN(new_n11614_));
  OAI21_X1   g10594(.A1(new_n11607_), .A2(new_n11614_), .B(new_n11601_), .ZN(new_n11615_));
  INV_X1     g10595(.I(new_n11601_), .ZN(new_n11616_));
  OAI21_X1   g10596(.A1(new_n11610_), .A2(new_n11611_), .B(new_n11613_), .ZN(new_n11617_));
  NAND3_X1   g10597(.A1(new_n11604_), .A2(new_n11605_), .A3(new_n11606_), .ZN(new_n11618_));
  NAND3_X1   g10598(.A1(new_n11617_), .A2(new_n11618_), .A3(new_n11616_), .ZN(new_n11619_));
  NAND2_X1   g10599(.A1(new_n11615_), .A2(new_n11619_), .ZN(new_n11620_));
  AOI21_X1   g10600(.A1(new_n11617_), .A2(new_n11618_), .B(new_n11616_), .ZN(new_n11621_));
  NOR3_X1    g10601(.A1(new_n11607_), .A2(new_n11614_), .A3(new_n11601_), .ZN(new_n11622_));
  NOR2_X1    g10602(.A1(new_n11564_), .A2(new_n11563_), .ZN(new_n11623_));
  NOR3_X1    g10603(.A1(new_n11623_), .A2(new_n11555_), .A3(new_n11556_), .ZN(new_n11624_));
  AOI21_X1   g10604(.A1(new_n9205_), .A2(new_n9206_), .B(new_n11557_), .ZN(new_n11625_));
  OAI21_X1   g10605(.A1(new_n11625_), .A2(new_n11624_), .B(new_n11560_), .ZN(new_n11626_));
  OAI21_X1   g10606(.A1(new_n11558_), .A2(new_n9236_), .B(new_n9235_), .ZN(new_n11627_));
  NAND2_X1   g10607(.A1(new_n11626_), .A2(new_n11627_), .ZN(new_n11628_));
  INV_X1     g10608(.I(new_n11628_), .ZN(new_n11629_));
  OAI21_X1   g10609(.A1(new_n11622_), .A2(new_n11621_), .B(new_n11629_), .ZN(new_n11630_));
  NAND3_X1   g10610(.A1(new_n11615_), .A2(new_n11619_), .A3(new_n11628_), .ZN(new_n11631_));
  INV_X1     g10611(.I(new_n11589_), .ZN(new_n11632_));
  NAND3_X1   g10612(.A1(new_n11632_), .A2(new_n11587_), .A3(new_n11600_), .ZN(new_n11633_));
  INV_X1     g10613(.I(new_n11586_), .ZN(new_n11634_));
  NOR3_X1    g10614(.A1(new_n11585_), .A2(new_n11582_), .A3(new_n11583_), .ZN(new_n11635_));
  NAND2_X1   g10615(.A1(new_n9221_), .A2(new_n8423_), .ZN(new_n11636_));
  XOR2_X1    g10616(.A1(new_n9223_), .A2(new_n11636_), .Z(new_n11637_));
  NOR3_X1    g10617(.A1(new_n11634_), .A2(new_n11635_), .A3(new_n11637_), .ZN(new_n11638_));
  NAND2_X1   g10618(.A1(new_n11633_), .A2(new_n11638_), .ZN(new_n11639_));
  NOR4_X1    g10619(.A1(new_n11588_), .A2(new_n11589_), .A3(new_n11598_), .A4(new_n11599_), .ZN(new_n11640_));
  INV_X1     g10620(.I(new_n11638_), .ZN(new_n11641_));
  NAND2_X1   g10621(.A1(new_n11640_), .A2(new_n11641_), .ZN(new_n11642_));
  XOR2_X1    g10622(.A1(new_n9228_), .A2(new_n9234_), .Z(new_n11643_));
  INV_X1     g10623(.I(new_n11643_), .ZN(new_n11644_));
  AOI22_X1   g10624(.A1(new_n11642_), .A2(new_n11639_), .B1(new_n11644_), .B2(new_n11633_), .ZN(new_n11645_));
  AOI22_X1   g10625(.A1(new_n11630_), .A2(new_n11631_), .B1(new_n11620_), .B2(new_n11645_), .ZN(new_n11646_));
  AOI22_X1   g10626(.A1(new_n11646_), .A2(new_n11521_), .B1(new_n11543_), .B2(new_n11570_), .ZN(new_n11647_));
  AOI22_X1   g10627(.A1(new_n11506_), .A2(new_n11511_), .B1(new_n11495_), .B2(new_n11647_), .ZN(new_n11648_));
  NOR3_X1    g10628(.A1(new_n11425_), .A2(new_n11422_), .A3(new_n11373_), .ZN(new_n11649_));
  NOR3_X1    g10629(.A1(new_n11475_), .A2(new_n11478_), .A3(new_n11473_), .ZN(new_n11650_));
  NAND2_X1   g10630(.A1(new_n11378_), .A2(new_n10687_), .ZN(new_n11651_));
  NAND2_X1   g10631(.A1(new_n11375_), .A2(new_n10688_), .ZN(new_n11652_));
  NAND2_X1   g10632(.A1(new_n11652_), .A2(new_n11651_), .ZN(new_n11653_));
  NAND2_X1   g10633(.A1(new_n10675_), .A2(new_n11653_), .ZN(new_n11654_));
  NAND3_X1   g10634(.A1(new_n10674_), .A2(new_n11651_), .A3(new_n11652_), .ZN(new_n11655_));
  AOI21_X1   g10635(.A1(new_n11655_), .A2(new_n11420_), .B(new_n11372_), .ZN(new_n11656_));
  NOR2_X1    g10636(.A1(new_n11654_), .A2(new_n11656_), .ZN(new_n11657_));
  NOR4_X1    g10637(.A1(new_n11657_), .A2(new_n11491_), .A3(new_n11470_), .A4(new_n11650_), .ZN(new_n11658_));
  XOR2_X1    g10638(.A1(new_n11381_), .A2(new_n11372_), .Z(new_n11659_));
  OAI21_X1   g10639(.A1(new_n11658_), .A2(new_n11649_), .B(new_n11659_), .ZN(new_n11660_));
  AOI21_X1   g10640(.A1(new_n9287_), .A2(new_n9293_), .B(new_n9305_), .ZN(new_n11661_));
  NAND3_X1   g10641(.A1(new_n9287_), .A2(new_n9293_), .A3(new_n9305_), .ZN(new_n11662_));
  INV_X1     g10642(.I(new_n11662_), .ZN(new_n11663_));
  OAI21_X1   g10643(.A1(new_n11663_), .A2(new_n11661_), .B(new_n9308_), .ZN(new_n11664_));
  NAND2_X1   g10644(.A1(new_n9294_), .A2(new_n9306_), .ZN(new_n11665_));
  NAND3_X1   g10645(.A1(new_n11665_), .A2(new_n9307_), .A3(new_n11662_), .ZN(new_n11666_));
  AND2_X2    g10646(.A1(new_n11664_), .A2(new_n11666_), .Z(new_n11667_));
  NAND2_X1   g10647(.A1(new_n11660_), .A2(new_n11667_), .ZN(new_n11668_));
  OAI21_X1   g10648(.A1(new_n11424_), .A2(new_n11423_), .B(new_n10687_), .ZN(new_n11669_));
  NAND3_X1   g10649(.A1(new_n11383_), .A2(new_n11421_), .A3(new_n11375_), .ZN(new_n11670_));
  NAND3_X1   g10650(.A1(new_n11669_), .A2(new_n11670_), .A3(new_n11372_), .ZN(new_n11671_));
  NAND3_X1   g10651(.A1(new_n11459_), .A2(new_n11461_), .A3(new_n11469_), .ZN(new_n11672_));
  INV_X1     g10652(.I(new_n10664_), .ZN(new_n11673_));
  INV_X1     g10653(.I(new_n10671_), .ZN(new_n11674_));
  OAI21_X1   g10654(.A1(new_n11674_), .A2(new_n10669_), .B(new_n10624_), .ZN(new_n11675_));
  AOI22_X1   g10655(.A1(new_n10679_), .A2(new_n11414_), .B1(new_n11675_), .B2(new_n11673_), .ZN(new_n11676_));
  AOI22_X1   g10656(.A1(new_n11676_), .A2(new_n11417_), .B1(new_n10625_), .B2(new_n10662_), .ZN(new_n11677_));
  NOR3_X1    g10657(.A1(new_n11677_), .A2(new_n11376_), .A3(new_n11379_), .ZN(new_n11678_));
  OAI21_X1   g10658(.A1(new_n11678_), .A2(new_n11374_), .B(new_n11373_), .ZN(new_n11679_));
  NAND3_X1   g10659(.A1(new_n11679_), .A2(new_n10675_), .A3(new_n11653_), .ZN(new_n11680_));
  NAND4_X1   g10660(.A1(new_n11680_), .A2(new_n11456_), .A3(new_n11492_), .A4(new_n11672_), .ZN(new_n11681_));
  NAND2_X1   g10661(.A1(new_n11681_), .A2(new_n11671_), .ZN(new_n11682_));
  NAND2_X1   g10662(.A1(new_n11664_), .A2(new_n11666_), .ZN(new_n11683_));
  NAND3_X1   g10663(.A1(new_n11682_), .A2(new_n11683_), .A3(new_n11659_), .ZN(new_n11684_));
  NAND3_X1   g10664(.A1(new_n11668_), .A2(new_n11648_), .A3(new_n11684_), .ZN(new_n11685_));
  NOR2_X1    g10665(.A1(new_n11497_), .A2(new_n11496_), .ZN(new_n11686_));
  AOI21_X1   g10666(.A1(new_n11480_), .A2(new_n11494_), .B(new_n11510_), .ZN(new_n11687_));
  NOR3_X1    g10667(.A1(new_n11497_), .A2(new_n11496_), .A3(new_n11505_), .ZN(new_n11688_));
  NAND2_X1   g10668(.A1(new_n11543_), .A2(new_n11570_), .ZN(new_n11689_));
  NOR2_X1    g10669(.A1(new_n11622_), .A2(new_n11621_), .ZN(new_n11690_));
  AOI21_X1   g10670(.A1(new_n11615_), .A2(new_n11619_), .B(new_n11628_), .ZN(new_n11691_));
  NOR3_X1    g10671(.A1(new_n11622_), .A2(new_n11621_), .A3(new_n11629_), .ZN(new_n11692_));
  INV_X1     g10672(.I(new_n11639_), .ZN(new_n11693_));
  NOR2_X1    g10673(.A1(new_n11633_), .A2(new_n11638_), .ZN(new_n11694_));
  OAI22_X1   g10674(.A1(new_n11693_), .A2(new_n11694_), .B1(new_n11640_), .B2(new_n11643_), .ZN(new_n11695_));
  OAI22_X1   g10675(.A1(new_n11692_), .A2(new_n11691_), .B1(new_n11690_), .B2(new_n11695_), .ZN(new_n11696_));
  OAI21_X1   g10676(.A1(new_n11520_), .A2(new_n11696_), .B(new_n11689_), .ZN(new_n11697_));
  OAI22_X1   g10677(.A1(new_n11687_), .A2(new_n11688_), .B1(new_n11686_), .B2(new_n11697_), .ZN(new_n11698_));
  AOI21_X1   g10678(.A1(new_n11682_), .A2(new_n11659_), .B(new_n11683_), .ZN(new_n11699_));
  NOR2_X1    g10679(.A1(new_n11660_), .A2(new_n11667_), .ZN(new_n11700_));
  OAI21_X1   g10680(.A1(new_n11700_), .A2(new_n11699_), .B(new_n11698_), .ZN(new_n11701_));
  NAND2_X1   g10681(.A1(new_n11701_), .A2(new_n11685_), .ZN(new_n11702_));
  NOR2_X1    g10682(.A1(new_n7592_), .A2(new_n7619_), .ZN(new_n11703_));
  NOR2_X1    g10683(.A1(new_n11703_), .A2(new_n7718_), .ZN(new_n11704_));
  NAND2_X1   g10684(.A1(new_n4281_), .A2(new_n4276_), .ZN(new_n11705_));
  AOI21_X1   g10685(.A1(new_n11705_), .A2(new_n4320_), .B(new_n4325_), .ZN(new_n11706_));
  NOR3_X1    g10686(.A1(new_n11706_), .A2(new_n7592_), .A3(new_n7619_), .ZN(new_n11707_));
  OAI21_X1   g10687(.A1(new_n11704_), .A2(new_n11707_), .B(new_n7710_), .ZN(new_n11708_));
  NAND2_X1   g10688(.A1(new_n7707_), .A2(new_n7708_), .ZN(new_n11709_));
  NOR3_X1    g10689(.A1(new_n11709_), .A2(new_n7626_), .A3(new_n7627_), .ZN(new_n11710_));
  NOR2_X1    g10690(.A1(new_n7642_), .A2(new_n7643_), .ZN(new_n11711_));
  NOR2_X1    g10691(.A1(new_n7639_), .A2(new_n7640_), .ZN(new_n11712_));
  OAI21_X1   g10692(.A1(new_n11711_), .A2(new_n11712_), .B(new_n4316_), .ZN(new_n11713_));
  OAI21_X1   g10693(.A1(new_n4224_), .A2(new_n4302_), .B(new_n4223_), .ZN(new_n11714_));
  NOR2_X1    g10694(.A1(new_n7651_), .A2(new_n7650_), .ZN(new_n11715_));
  NOR2_X1    g10695(.A1(new_n7647_), .A2(new_n7648_), .ZN(new_n11716_));
  OAI21_X1   g10696(.A1(new_n11716_), .A2(new_n11715_), .B(new_n7522_), .ZN(new_n11717_));
  OAI21_X1   g10697(.A1(new_n7524_), .A2(new_n7612_), .B(new_n7523_), .ZN(new_n11718_));
  NAND4_X1   g10698(.A1(new_n11717_), .A2(new_n11713_), .A3(new_n11714_), .A4(new_n11718_), .ZN(new_n11719_));
  NAND2_X1   g10699(.A1(new_n7523_), .A2(new_n7656_), .ZN(new_n11720_));
  NAND2_X1   g10700(.A1(new_n7661_), .A2(new_n7662_), .ZN(new_n11721_));
  OAI21_X1   g10701(.A1(new_n4202_), .A2(new_n4203_), .B(new_n7659_), .ZN(new_n11722_));
  AOI21_X1   g10702(.A1(new_n11722_), .A2(new_n11721_), .B(new_n4314_), .ZN(new_n11723_));
  INV_X1     g10703(.I(new_n7665_), .ZN(new_n11724_));
  NOR3_X1    g10704(.A1(new_n11720_), .A2(new_n11724_), .A3(new_n11723_), .ZN(new_n11725_));
  INV_X1     g10705(.I(new_n7695_), .ZN(new_n11726_));
  AOI22_X1   g10706(.A1(new_n11726_), .A2(new_n7667_), .B1(new_n7681_), .B2(new_n7682_), .ZN(new_n11727_));
  NAND2_X1   g10707(.A1(new_n7664_), .A2(new_n7665_), .ZN(new_n11728_));
  NAND2_X1   g10708(.A1(new_n11728_), .A2(new_n11720_), .ZN(new_n11729_));
  AOI21_X1   g10709(.A1(new_n11729_), .A2(new_n11727_), .B(new_n11725_), .ZN(new_n11730_));
  AOI22_X1   g10710(.A1(new_n11717_), .A2(new_n11718_), .B1(new_n11713_), .B2(new_n11714_), .ZN(new_n11731_));
  OAI21_X1   g10711(.A1(new_n11731_), .A2(new_n11730_), .B(new_n11719_), .ZN(new_n11732_));
  OAI22_X1   g10712(.A1(new_n7626_), .A2(new_n7627_), .B1(new_n7635_), .B2(new_n7636_), .ZN(new_n11733_));
  AOI21_X1   g10713(.A1(new_n11732_), .A2(new_n11733_), .B(new_n11710_), .ZN(new_n11734_));
  AOI22_X1   g10714(.A1(new_n7721_), .A2(new_n7724_), .B1(new_n7714_), .B2(new_n7717_), .ZN(new_n11735_));
  OAI21_X1   g10715(.A1(new_n11735_), .A2(new_n7620_), .B(new_n11734_), .ZN(new_n11736_));
  NAND3_X1   g10716(.A1(new_n11708_), .A2(new_n11702_), .A3(new_n11736_), .ZN(new_n11737_));
  NOR3_X1    g10717(.A1(new_n11700_), .A2(new_n11699_), .A3(new_n11698_), .ZN(new_n11738_));
  AOI21_X1   g10718(.A1(new_n11668_), .A2(new_n11684_), .B(new_n11648_), .ZN(new_n11739_));
  NOR2_X1    g10719(.A1(new_n11738_), .A2(new_n11739_), .ZN(new_n11740_));
  NAND2_X1   g10720(.A1(new_n7725_), .A2(new_n11706_), .ZN(new_n11741_));
  NAND2_X1   g10721(.A1(new_n11703_), .A2(new_n7718_), .ZN(new_n11742_));
  AOI21_X1   g10722(.A1(new_n11742_), .A2(new_n11741_), .B(new_n11734_), .ZN(new_n11743_));
  NAND4_X1   g10723(.A1(new_n7721_), .A2(new_n7724_), .A3(new_n7714_), .A4(new_n7717_), .ZN(new_n11744_));
  AOI21_X1   g10724(.A1(new_n7726_), .A2(new_n11744_), .B(new_n7710_), .ZN(new_n11745_));
  OAI21_X1   g10725(.A1(new_n11743_), .A2(new_n11745_), .B(new_n11740_), .ZN(new_n11746_));
  NAND2_X1   g10726(.A1(new_n11492_), .A2(new_n11493_), .ZN(new_n11747_));
  NAND2_X1   g10727(.A1(new_n11520_), .A2(new_n11569_), .ZN(new_n11748_));
  NAND2_X1   g10728(.A1(new_n11689_), .A2(new_n11696_), .ZN(new_n11749_));
  NAND3_X1   g10729(.A1(new_n11749_), .A2(new_n11747_), .A3(new_n11748_), .ZN(new_n11750_));
  NOR2_X1    g10730(.A1(new_n11479_), .A2(new_n11470_), .ZN(new_n11751_));
  NAND2_X1   g10731(.A1(new_n11647_), .A2(new_n11751_), .ZN(new_n11752_));
  AOI21_X1   g10732(.A1(new_n11752_), .A2(new_n11750_), .B(new_n11510_), .ZN(new_n11753_));
  NOR2_X1    g10733(.A1(new_n11647_), .A2(new_n11751_), .ZN(new_n11754_));
  AOI21_X1   g10734(.A1(new_n11749_), .A2(new_n11748_), .B(new_n11747_), .ZN(new_n11755_));
  NOR3_X1    g10735(.A1(new_n11754_), .A2(new_n11755_), .A3(new_n11505_), .ZN(new_n11756_));
  OAI21_X1   g10736(.A1(new_n11756_), .A2(new_n11753_), .B(new_n11456_), .ZN(new_n11757_));
  OAI21_X1   g10737(.A1(new_n11754_), .A2(new_n11755_), .B(new_n11505_), .ZN(new_n11758_));
  NAND3_X1   g10738(.A1(new_n11752_), .A2(new_n11750_), .A3(new_n11510_), .ZN(new_n11759_));
  NAND3_X1   g10739(.A1(new_n11758_), .A2(new_n11759_), .A3(new_n11491_), .ZN(new_n11760_));
  NAND2_X1   g10740(.A1(new_n7703_), .A2(new_n7704_), .ZN(new_n11761_));
  NOR2_X1    g10741(.A1(new_n11761_), .A2(new_n7637_), .ZN(new_n11762_));
  NOR2_X1    g10742(.A1(new_n7628_), .A2(new_n11709_), .ZN(new_n11763_));
  OAI21_X1   g10743(.A1(new_n11762_), .A2(new_n11763_), .B(new_n11732_), .ZN(new_n11764_));
  OAI21_X1   g10744(.A1(new_n11710_), .A2(new_n7709_), .B(new_n7700_), .ZN(new_n11765_));
  NAND4_X1   g10745(.A1(new_n11757_), .A2(new_n11760_), .A3(new_n11764_), .A4(new_n11765_), .ZN(new_n11766_));
  NOR2_X1    g10746(.A1(new_n7645_), .A2(new_n7646_), .ZN(new_n11767_));
  NAND2_X1   g10747(.A1(new_n11717_), .A2(new_n11718_), .ZN(new_n11768_));
  NAND2_X1   g10748(.A1(new_n11768_), .A2(new_n11767_), .ZN(new_n11769_));
  NAND2_X1   g10749(.A1(new_n11713_), .A2(new_n11714_), .ZN(new_n11770_));
  NOR2_X1    g10750(.A1(new_n7653_), .A2(new_n7654_), .ZN(new_n11771_));
  NAND2_X1   g10751(.A1(new_n11771_), .A2(new_n11770_), .ZN(new_n11772_));
  AOI21_X1   g10752(.A1(new_n11769_), .A2(new_n11772_), .B(new_n11730_), .ZN(new_n11773_));
  AOI21_X1   g10753(.A1(new_n7699_), .A2(new_n11719_), .B(new_n7698_), .ZN(new_n11774_));
  NOR2_X1    g10754(.A1(new_n11646_), .A2(new_n11520_), .ZN(new_n11775_));
  NOR2_X1    g10755(.A1(new_n11696_), .A2(new_n11521_), .ZN(new_n11776_));
  OAI21_X1   g10756(.A1(new_n11776_), .A2(new_n11775_), .B(new_n11542_), .ZN(new_n11777_));
  NAND2_X1   g10757(.A1(new_n11696_), .A2(new_n11521_), .ZN(new_n11778_));
  NAND2_X1   g10758(.A1(new_n11646_), .A2(new_n11520_), .ZN(new_n11779_));
  NAND3_X1   g10759(.A1(new_n11778_), .A2(new_n11779_), .A3(new_n11569_), .ZN(new_n11780_));
  NAND2_X1   g10760(.A1(new_n11777_), .A2(new_n11780_), .ZN(new_n11781_));
  NOR3_X1    g10761(.A1(new_n11773_), .A2(new_n11781_), .A3(new_n11774_), .ZN(new_n11782_));
  NAND2_X1   g10762(.A1(new_n11617_), .A2(new_n11618_), .ZN(new_n11783_));
  NAND2_X1   g10763(.A1(new_n11695_), .A2(new_n11783_), .ZN(new_n11784_));
  NOR2_X1    g10764(.A1(new_n11607_), .A2(new_n11614_), .ZN(new_n11785_));
  NAND2_X1   g10765(.A1(new_n11645_), .A2(new_n11785_), .ZN(new_n11786_));
  AOI21_X1   g10766(.A1(new_n11784_), .A2(new_n11786_), .B(new_n11628_), .ZN(new_n11787_));
  NOR2_X1    g10767(.A1(new_n11645_), .A2(new_n11785_), .ZN(new_n11788_));
  INV_X1     g10768(.I(new_n11786_), .ZN(new_n11789_));
  NOR3_X1    g10769(.A1(new_n11789_), .A2(new_n11788_), .A3(new_n11629_), .ZN(new_n11790_));
  OAI21_X1   g10770(.A1(new_n11790_), .A2(new_n11787_), .B(new_n11601_), .ZN(new_n11791_));
  NOR3_X1    g10771(.A1(new_n11790_), .A2(new_n11601_), .A3(new_n11787_), .ZN(new_n11792_));
  INV_X1     g10772(.I(new_n11792_), .ZN(new_n11793_));
  NOR2_X1    g10773(.A1(new_n11724_), .A2(new_n11723_), .ZN(new_n11794_));
  NOR2_X1    g10774(.A1(new_n11794_), .A2(new_n11720_), .ZN(new_n11795_));
  NOR2_X1    g10775(.A1(new_n11728_), .A2(new_n7658_), .ZN(new_n11796_));
  OAI21_X1   g10776(.A1(new_n11795_), .A2(new_n11796_), .B(new_n11727_), .ZN(new_n11797_));
  OAI21_X1   g10777(.A1(new_n11725_), .A2(new_n7697_), .B(new_n7696_), .ZN(new_n11798_));
  NAND4_X1   g10778(.A1(new_n11793_), .A2(new_n11797_), .A3(new_n11798_), .A4(new_n11791_), .ZN(new_n11799_));
  NAND3_X1   g10779(.A1(new_n7682_), .A2(new_n7695_), .A3(new_n7681_), .ZN(new_n11800_));
  INV_X1     g10780(.I(new_n11800_), .ZN(new_n11801_));
  NAND2_X1   g10781(.A1(new_n7678_), .A2(new_n7670_), .ZN(new_n11802_));
  NAND2_X1   g10782(.A1(new_n7680_), .A2(new_n11802_), .ZN(new_n11803_));
  XOR2_X1    g10783(.A1(new_n11637_), .A2(new_n11582_), .Z(new_n11804_));
  XOR2_X1    g10784(.A1(new_n11804_), .A2(new_n11584_), .Z(new_n11805_));
  XOR2_X1    g10785(.A1(new_n11805_), .A2(new_n10568_), .Z(new_n11806_));
  NOR2_X1    g10786(.A1(new_n11803_), .A2(new_n11806_), .ZN(new_n11807_));
  XOR2_X1    g10787(.A1(new_n11800_), .A2(new_n11807_), .Z(new_n11808_));
  NAND2_X1   g10788(.A1(new_n11642_), .A2(new_n11639_), .ZN(new_n11809_));
  XOR2_X1    g10789(.A1(new_n11809_), .A2(new_n11644_), .Z(new_n11810_));
  INV_X1     g10790(.I(new_n11810_), .ZN(new_n11811_));
  OAI21_X1   g10791(.A1(new_n11801_), .A2(new_n11811_), .B(new_n11808_), .ZN(new_n11812_));
  INV_X1     g10792(.I(new_n11787_), .ZN(new_n11813_));
  NAND3_X1   g10793(.A1(new_n11784_), .A2(new_n11786_), .A3(new_n11628_), .ZN(new_n11814_));
  AOI21_X1   g10794(.A1(new_n11813_), .A2(new_n11814_), .B(new_n11616_), .ZN(new_n11815_));
  NOR2_X1    g10795(.A1(new_n11815_), .A2(new_n11792_), .ZN(new_n11816_));
  NAND2_X1   g10796(.A1(new_n11728_), .A2(new_n7658_), .ZN(new_n11817_));
  NAND2_X1   g10797(.A1(new_n11794_), .A2(new_n11720_), .ZN(new_n11818_));
  AOI21_X1   g10798(.A1(new_n11818_), .A2(new_n11817_), .B(new_n7696_), .ZN(new_n11819_));
  AOI21_X1   g10799(.A1(new_n11729_), .A2(new_n7666_), .B(new_n11727_), .ZN(new_n11820_));
  NOR2_X1    g10800(.A1(new_n11819_), .A2(new_n11820_), .ZN(new_n11821_));
  NOR2_X1    g10801(.A1(new_n11821_), .A2(new_n11816_), .ZN(new_n11822_));
  OAI21_X1   g10802(.A1(new_n11822_), .A2(new_n11812_), .B(new_n11799_), .ZN(new_n11823_));
  OAI21_X1   g10803(.A1(new_n11773_), .A2(new_n11774_), .B(new_n11781_), .ZN(new_n11824_));
  AOI21_X1   g10804(.A1(new_n11823_), .A2(new_n11824_), .B(new_n11782_), .ZN(new_n11825_));
  AOI22_X1   g10805(.A1(new_n11757_), .A2(new_n11760_), .B1(new_n11764_), .B2(new_n11765_), .ZN(new_n11826_));
  OAI21_X1   g10806(.A1(new_n11826_), .A2(new_n11825_), .B(new_n11766_), .ZN(new_n11827_));
  AOI22_X1   g10807(.A1(new_n11746_), .A2(new_n11737_), .B1(new_n11827_), .B2(new_n11702_), .ZN(new_n11828_));
  NAND2_X1   g10808(.A1(new_n11828_), .A2(new_n11432_), .ZN(new_n11829_));
  NOR2_X1    g10809(.A1(new_n11828_), .A2(new_n11432_), .ZN(new_n11830_));
  XOR2_X1    g10810(.A1(new_n11431_), .A2(new_n9309_), .Z(new_n11831_));
  NOR3_X1    g10811(.A1(new_n11743_), .A2(new_n11745_), .A3(new_n11740_), .ZN(new_n11832_));
  AOI21_X1   g10812(.A1(new_n11708_), .A2(new_n11736_), .B(new_n11702_), .ZN(new_n11833_));
  AOI21_X1   g10813(.A1(new_n11758_), .A2(new_n11759_), .B(new_n11491_), .ZN(new_n11834_));
  NOR3_X1    g10814(.A1(new_n11756_), .A2(new_n11753_), .A3(new_n11456_), .ZN(new_n11835_));
  NAND2_X1   g10815(.A1(new_n7628_), .A2(new_n11709_), .ZN(new_n11836_));
  NAND2_X1   g10816(.A1(new_n11761_), .A2(new_n7637_), .ZN(new_n11837_));
  AOI21_X1   g10817(.A1(new_n11837_), .A2(new_n11836_), .B(new_n7700_), .ZN(new_n11838_));
  AOI21_X1   g10818(.A1(new_n7638_), .A2(new_n11733_), .B(new_n11732_), .ZN(new_n11839_));
  NOR4_X1    g10819(.A1(new_n11835_), .A2(new_n11834_), .A3(new_n11838_), .A4(new_n11839_), .ZN(new_n11840_));
  NOR2_X1    g10820(.A1(new_n11771_), .A2(new_n11770_), .ZN(new_n11841_));
  NOR2_X1    g10821(.A1(new_n11768_), .A2(new_n11767_), .ZN(new_n11842_));
  OAI21_X1   g10822(.A1(new_n11842_), .A2(new_n11841_), .B(new_n7698_), .ZN(new_n11843_));
  OAI21_X1   g10823(.A1(new_n11731_), .A2(new_n7655_), .B(new_n11730_), .ZN(new_n11844_));
  AOI21_X1   g10824(.A1(new_n11778_), .A2(new_n11779_), .B(new_n11569_), .ZN(new_n11845_));
  NOR3_X1    g10825(.A1(new_n11776_), .A2(new_n11775_), .A3(new_n11542_), .ZN(new_n11846_));
  NOR2_X1    g10826(.A1(new_n11845_), .A2(new_n11846_), .ZN(new_n11847_));
  NAND3_X1   g10827(.A1(new_n11843_), .A2(new_n11847_), .A3(new_n11844_), .ZN(new_n11848_));
  NOR4_X1    g10828(.A1(new_n11819_), .A2(new_n11815_), .A3(new_n11820_), .A4(new_n11792_), .ZN(new_n11849_));
  XNOR2_X1   g10829(.A1(new_n11800_), .A2(new_n11807_), .ZN(new_n11850_));
  AOI21_X1   g10830(.A1(new_n11800_), .A2(new_n11810_), .B(new_n11850_), .ZN(new_n11851_));
  OAI22_X1   g10831(.A1(new_n11819_), .A2(new_n11820_), .B1(new_n11815_), .B2(new_n11792_), .ZN(new_n11852_));
  AOI21_X1   g10832(.A1(new_n11852_), .A2(new_n11851_), .B(new_n11849_), .ZN(new_n11853_));
  AOI21_X1   g10833(.A1(new_n11843_), .A2(new_n11844_), .B(new_n11847_), .ZN(new_n11854_));
  OAI21_X1   g10834(.A1(new_n11854_), .A2(new_n11853_), .B(new_n11848_), .ZN(new_n11855_));
  OAI22_X1   g10835(.A1(new_n11835_), .A2(new_n11834_), .B1(new_n11838_), .B2(new_n11839_), .ZN(new_n11856_));
  AOI21_X1   g10836(.A1(new_n11855_), .A2(new_n11856_), .B(new_n11840_), .ZN(new_n11857_));
  OAI22_X1   g10837(.A1(new_n11832_), .A2(new_n11833_), .B1(new_n11857_), .B2(new_n11740_), .ZN(new_n11858_));
  NOR2_X1    g10838(.A1(new_n11858_), .A2(new_n11831_), .ZN(new_n11859_));
  NAND2_X1   g10839(.A1(new_n7744_), .A2(new_n7748_), .ZN(new_n11860_));
  NAND3_X1   g10840(.A1(new_n11860_), .A2(new_n7766_), .A3(new_n7770_), .ZN(new_n11861_));
  AOI21_X1   g10841(.A1(new_n7746_), .A2(new_n7747_), .B(new_n7745_), .ZN(new_n11862_));
  NOR3_X1    g10842(.A1(new_n7743_), .A2(new_n7739_), .A3(new_n7730_), .ZN(new_n11863_));
  NOR2_X1    g10843(.A1(new_n11863_), .A2(new_n11862_), .ZN(new_n11864_));
  NAND2_X1   g10844(.A1(new_n7766_), .A2(new_n7770_), .ZN(new_n11865_));
  NAND2_X1   g10845(.A1(new_n11865_), .A2(new_n11864_), .ZN(new_n11866_));
  AOI21_X1   g10846(.A1(new_n11866_), .A2(new_n11861_), .B(new_n7727_), .ZN(new_n11867_));
  OAI21_X1   g10847(.A1(new_n11734_), .A2(new_n11735_), .B(new_n11744_), .ZN(new_n11868_));
  AOI21_X1   g10848(.A1(new_n7769_), .A2(new_n7768_), .B(new_n7767_), .ZN(new_n11869_));
  NOR3_X1    g10849(.A1(new_n7762_), .A2(new_n7765_), .A3(new_n7751_), .ZN(new_n11870_));
  OAI22_X1   g10850(.A1(new_n11869_), .A2(new_n11870_), .B1(new_n11862_), .B2(new_n11863_), .ZN(new_n11871_));
  AOI21_X1   g10851(.A1(new_n11871_), .A2(new_n7771_), .B(new_n11868_), .ZN(new_n11872_));
  NOR2_X1    g10852(.A1(new_n11867_), .A2(new_n11872_), .ZN(new_n11873_));
  OAI21_X1   g10853(.A1(new_n11859_), .A2(new_n11830_), .B(new_n11873_), .ZN(new_n11874_));
  NAND2_X1   g10854(.A1(new_n11874_), .A2(new_n11829_), .ZN(new_n11875_));
  AOI21_X1   g10855(.A1(new_n7772_), .A2(new_n7777_), .B(new_n7789_), .ZN(new_n11876_));
  INV_X1     g10856(.I(new_n11876_), .ZN(new_n11877_));
  NAND3_X1   g10857(.A1(new_n7772_), .A2(new_n7777_), .A3(new_n7789_), .ZN(new_n11878_));
  NAND3_X1   g10858(.A1(new_n11877_), .A2(new_n7788_), .A3(new_n11878_), .ZN(new_n11879_));
  NAND2_X1   g10859(.A1(new_n11431_), .A2(new_n9309_), .ZN(new_n11880_));
  NOR2_X1    g10860(.A1(new_n11428_), .A2(new_n10689_), .ZN(new_n11881_));
  NOR3_X1    g10861(.A1(new_n11431_), .A2(new_n9309_), .A3(new_n11881_), .ZN(new_n11882_));
  XOR2_X1    g10862(.A1(new_n11882_), .A2(new_n11880_), .Z(new_n11883_));
  INV_X1     g10863(.I(new_n11878_), .ZN(new_n11884_));
  OAI21_X1   g10864(.A1(new_n11884_), .A2(new_n11876_), .B(new_n7782_), .ZN(new_n11885_));
  NAND3_X1   g10865(.A1(new_n11879_), .A2(new_n11885_), .A3(new_n11883_), .ZN(new_n11886_));
  XNOR2_X1   g10866(.A1(new_n7785_), .A2(new_n7782_), .ZN(new_n11887_));
  INV_X1     g10867(.I(new_n11887_), .ZN(new_n11888_));
  NOR3_X1    g10868(.A1(new_n11888_), .A2(new_n7778_), .A3(new_n11883_), .ZN(new_n11889_));
  NAND2_X1   g10869(.A1(new_n11886_), .A2(new_n11889_), .ZN(new_n11890_));
  OAI21_X1   g10870(.A1(new_n11890_), .A2(new_n11875_), .B(new_n11429_), .ZN(new_n11891_));
  NAND2_X1   g10871(.A1(new_n11891_), .A2(new_n11430_), .ZN(new_n11892_));
  INV_X1     g10872(.I(\A[814] ), .ZN(new_n11893_));
  NOR2_X1    g10873(.A1(\A[815] ), .A2(\A[816] ), .ZN(new_n11894_));
  NAND2_X1   g10874(.A1(\A[815] ), .A2(\A[816] ), .ZN(new_n11895_));
  AOI21_X1   g10875(.A1(new_n11893_), .A2(new_n11895_), .B(new_n11894_), .ZN(new_n11896_));
  INV_X1     g10876(.I(new_n11896_), .ZN(new_n11897_));
  INV_X1     g10877(.I(\A[811] ), .ZN(new_n11898_));
  NOR2_X1    g10878(.A1(\A[812] ), .A2(\A[813] ), .ZN(new_n11899_));
  NAND2_X1   g10879(.A1(\A[812] ), .A2(\A[813] ), .ZN(new_n11900_));
  AOI21_X1   g10880(.A1(new_n11898_), .A2(new_n11900_), .B(new_n11899_), .ZN(new_n11901_));
  INV_X1     g10881(.I(new_n11901_), .ZN(new_n11902_));
  INV_X1     g10882(.I(\A[812] ), .ZN(new_n11903_));
  NAND2_X1   g10883(.A1(new_n11903_), .A2(\A[813] ), .ZN(new_n11904_));
  INV_X1     g10884(.I(\A[813] ), .ZN(new_n11905_));
  NAND2_X1   g10885(.A1(new_n11905_), .A2(\A[812] ), .ZN(new_n11906_));
  AOI21_X1   g10886(.A1(new_n11904_), .A2(new_n11906_), .B(new_n11898_), .ZN(new_n11907_));
  INV_X1     g10887(.I(new_n11899_), .ZN(new_n11908_));
  AOI21_X1   g10888(.A1(new_n11908_), .A2(new_n11900_), .B(\A[811] ), .ZN(new_n11909_));
  INV_X1     g10889(.I(\A[815] ), .ZN(new_n11910_));
  NAND2_X1   g10890(.A1(new_n11910_), .A2(\A[816] ), .ZN(new_n11911_));
  INV_X1     g10891(.I(\A[816] ), .ZN(new_n11912_));
  NAND2_X1   g10892(.A1(new_n11912_), .A2(\A[815] ), .ZN(new_n11913_));
  AOI21_X1   g10893(.A1(new_n11911_), .A2(new_n11913_), .B(new_n11893_), .ZN(new_n11914_));
  INV_X1     g10894(.I(new_n11894_), .ZN(new_n11915_));
  AOI21_X1   g10895(.A1(new_n11915_), .A2(new_n11895_), .B(\A[814] ), .ZN(new_n11916_));
  NOR4_X1    g10896(.A1(new_n11907_), .A2(new_n11909_), .A3(new_n11916_), .A4(new_n11914_), .ZN(new_n11917_));
  NOR2_X1    g10897(.A1(new_n11917_), .A2(new_n11902_), .ZN(new_n11918_));
  INV_X1     g10898(.I(new_n11918_), .ZN(new_n11919_));
  NAND2_X1   g10899(.A1(new_n11917_), .A2(new_n11902_), .ZN(new_n11920_));
  AOI21_X1   g10900(.A1(new_n11919_), .A2(new_n11920_), .B(new_n11897_), .ZN(new_n11921_));
  INV_X1     g10901(.I(new_n11920_), .ZN(new_n11922_));
  NOR3_X1    g10902(.A1(new_n11922_), .A2(new_n11896_), .A3(new_n11918_), .ZN(new_n11923_));
  NOR2_X1    g10903(.A1(new_n11921_), .A2(new_n11923_), .ZN(new_n11924_));
  INV_X1     g10904(.I(\A[820] ), .ZN(new_n11925_));
  NOR2_X1    g10905(.A1(\A[821] ), .A2(\A[822] ), .ZN(new_n11926_));
  NAND2_X1   g10906(.A1(\A[821] ), .A2(\A[822] ), .ZN(new_n11927_));
  AOI21_X1   g10907(.A1(new_n11925_), .A2(new_n11927_), .B(new_n11926_), .ZN(new_n11928_));
  INV_X1     g10908(.I(new_n11928_), .ZN(new_n11929_));
  INV_X1     g10909(.I(\A[817] ), .ZN(new_n11930_));
  NOR2_X1    g10910(.A1(\A[818] ), .A2(\A[819] ), .ZN(new_n11931_));
  NAND2_X1   g10911(.A1(\A[818] ), .A2(\A[819] ), .ZN(new_n11932_));
  AOI21_X1   g10912(.A1(new_n11930_), .A2(new_n11932_), .B(new_n11931_), .ZN(new_n11933_));
  INV_X1     g10913(.I(\A[818] ), .ZN(new_n11934_));
  NAND2_X1   g10914(.A1(new_n11934_), .A2(\A[819] ), .ZN(new_n11935_));
  INV_X1     g10915(.I(\A[819] ), .ZN(new_n11936_));
  NAND2_X1   g10916(.A1(new_n11936_), .A2(\A[818] ), .ZN(new_n11937_));
  AOI21_X1   g10917(.A1(new_n11935_), .A2(new_n11937_), .B(new_n11930_), .ZN(new_n11938_));
  INV_X1     g10918(.I(new_n11931_), .ZN(new_n11939_));
  AOI21_X1   g10919(.A1(new_n11939_), .A2(new_n11932_), .B(\A[817] ), .ZN(new_n11940_));
  NOR2_X1    g10920(.A1(new_n11940_), .A2(new_n11938_), .ZN(new_n11941_));
  INV_X1     g10921(.I(\A[821] ), .ZN(new_n11942_));
  NAND2_X1   g10922(.A1(new_n11942_), .A2(\A[822] ), .ZN(new_n11943_));
  INV_X1     g10923(.I(\A[822] ), .ZN(new_n11944_));
  NAND2_X1   g10924(.A1(new_n11944_), .A2(\A[821] ), .ZN(new_n11945_));
  AOI21_X1   g10925(.A1(new_n11943_), .A2(new_n11945_), .B(new_n11925_), .ZN(new_n11946_));
  INV_X1     g10926(.I(new_n11926_), .ZN(new_n11947_));
  AOI21_X1   g10927(.A1(new_n11947_), .A2(new_n11927_), .B(\A[820] ), .ZN(new_n11948_));
  NOR2_X1    g10928(.A1(new_n11948_), .A2(new_n11946_), .ZN(new_n11949_));
  NAND2_X1   g10929(.A1(new_n11941_), .A2(new_n11949_), .ZN(new_n11950_));
  NAND2_X1   g10930(.A1(new_n11950_), .A2(new_n11933_), .ZN(new_n11951_));
  INV_X1     g10931(.I(new_n11933_), .ZN(new_n11952_));
  NOR2_X1    g10932(.A1(new_n11936_), .A2(\A[818] ), .ZN(new_n11953_));
  NOR2_X1    g10933(.A1(new_n11934_), .A2(\A[819] ), .ZN(new_n11954_));
  OAI21_X1   g10934(.A1(new_n11953_), .A2(new_n11954_), .B(\A[817] ), .ZN(new_n11955_));
  INV_X1     g10935(.I(new_n11932_), .ZN(new_n11956_));
  OAI21_X1   g10936(.A1(new_n11956_), .A2(new_n11931_), .B(new_n11930_), .ZN(new_n11957_));
  NAND2_X1   g10937(.A1(new_n11955_), .A2(new_n11957_), .ZN(new_n11958_));
  NOR2_X1    g10938(.A1(new_n11944_), .A2(\A[821] ), .ZN(new_n11959_));
  NOR2_X1    g10939(.A1(new_n11942_), .A2(\A[822] ), .ZN(new_n11960_));
  OAI21_X1   g10940(.A1(new_n11959_), .A2(new_n11960_), .B(\A[820] ), .ZN(new_n11961_));
  INV_X1     g10941(.I(new_n11927_), .ZN(new_n11962_));
  OAI21_X1   g10942(.A1(new_n11962_), .A2(new_n11926_), .B(new_n11925_), .ZN(new_n11963_));
  NAND2_X1   g10943(.A1(new_n11961_), .A2(new_n11963_), .ZN(new_n11964_));
  NOR2_X1    g10944(.A1(new_n11958_), .A2(new_n11964_), .ZN(new_n11965_));
  NAND2_X1   g10945(.A1(new_n11965_), .A2(new_n11952_), .ZN(new_n11966_));
  AOI21_X1   g10946(.A1(new_n11966_), .A2(new_n11951_), .B(new_n11929_), .ZN(new_n11967_));
  NOR2_X1    g10947(.A1(new_n11965_), .A2(new_n11952_), .ZN(new_n11968_));
  NOR2_X1    g10948(.A1(new_n11950_), .A2(new_n11933_), .ZN(new_n11969_));
  NOR3_X1    g10949(.A1(new_n11968_), .A2(new_n11969_), .A3(new_n11928_), .ZN(new_n11970_));
  NOR2_X1    g10950(.A1(new_n11967_), .A2(new_n11970_), .ZN(new_n11971_));
  NOR2_X1    g10951(.A1(new_n11909_), .A2(new_n11907_), .ZN(new_n11972_));
  NOR2_X1    g10952(.A1(new_n11916_), .A2(new_n11914_), .ZN(new_n11973_));
  NAND2_X1   g10953(.A1(new_n11972_), .A2(new_n11973_), .ZN(new_n11974_));
  NAND2_X1   g10954(.A1(new_n11896_), .A2(new_n11901_), .ZN(new_n11975_));
  NOR2_X1    g10955(.A1(new_n11941_), .A2(new_n11949_), .ZN(new_n11976_));
  NOR4_X1    g10956(.A1(new_n11965_), .A2(new_n11976_), .A3(new_n11974_), .A4(new_n11975_), .ZN(new_n11977_));
  NOR2_X1    g10957(.A1(new_n11972_), .A2(new_n11973_), .ZN(new_n11978_));
  NOR2_X1    g10958(.A1(new_n11978_), .A2(new_n11917_), .ZN(new_n11979_));
  NAND2_X1   g10959(.A1(new_n11928_), .A2(new_n11933_), .ZN(new_n11980_));
  NOR3_X1    g10960(.A1(new_n11958_), .A2(new_n11964_), .A3(new_n11980_), .ZN(new_n11981_));
  NAND3_X1   g10961(.A1(new_n11977_), .A2(new_n11979_), .A3(new_n11981_), .ZN(new_n11982_));
  NOR2_X1    g10962(.A1(new_n11971_), .A2(new_n11982_), .ZN(new_n11983_));
  OAI21_X1   g10963(.A1(new_n11968_), .A2(new_n11969_), .B(new_n11928_), .ZN(new_n11984_));
  NAND3_X1   g10964(.A1(new_n11966_), .A2(new_n11951_), .A3(new_n11929_), .ZN(new_n11985_));
  NAND2_X1   g10965(.A1(new_n11984_), .A2(new_n11985_), .ZN(new_n11986_));
  INV_X1     g10966(.I(new_n11982_), .ZN(new_n11987_));
  NOR2_X1    g10967(.A1(new_n11987_), .A2(new_n11986_), .ZN(new_n11988_));
  OAI21_X1   g10968(.A1(new_n11988_), .A2(new_n11983_), .B(new_n11924_), .ZN(new_n11989_));
  NAND2_X1   g10969(.A1(new_n11977_), .A2(new_n11979_), .ZN(new_n11990_));
  OAI22_X1   g10970(.A1(new_n11986_), .A2(new_n11990_), .B1(new_n11976_), .B2(new_n11980_), .ZN(new_n11991_));
  NAND2_X1   g10971(.A1(new_n11987_), .A2(new_n11971_), .ZN(new_n11992_));
  NAND3_X1   g10972(.A1(new_n11991_), .A2(new_n11992_), .A3(new_n11924_), .ZN(new_n11993_));
  NAND2_X1   g10973(.A1(new_n11993_), .A2(new_n11989_), .ZN(new_n11994_));
  INV_X1     g10974(.I(new_n11924_), .ZN(new_n11995_));
  NAND2_X1   g10975(.A1(new_n11987_), .A2(new_n11986_), .ZN(new_n11996_));
  NAND2_X1   g10976(.A1(new_n11971_), .A2(new_n11982_), .ZN(new_n11997_));
  AOI21_X1   g10977(.A1(new_n11996_), .A2(new_n11997_), .B(new_n11995_), .ZN(new_n11998_));
  INV_X1     g10978(.I(new_n11990_), .ZN(new_n11999_));
  NOR2_X1    g10979(.A1(new_n11976_), .A2(new_n11980_), .ZN(new_n12000_));
  AOI21_X1   g10980(.A1(new_n11971_), .A2(new_n11999_), .B(new_n12000_), .ZN(new_n12001_));
  NOR2_X1    g10981(.A1(new_n11986_), .A2(new_n11982_), .ZN(new_n12002_));
  NOR3_X1    g10982(.A1(new_n12001_), .A2(new_n12002_), .A3(new_n11995_), .ZN(new_n12003_));
  NOR2_X1    g10983(.A1(new_n11976_), .A2(new_n11965_), .ZN(new_n12004_));
  NAND2_X1   g10984(.A1(new_n12004_), .A2(new_n11981_), .ZN(new_n12005_));
  NOR2_X1    g10985(.A1(new_n11974_), .A2(new_n11975_), .ZN(new_n12006_));
  NAND2_X1   g10986(.A1(new_n11979_), .A2(new_n12006_), .ZN(new_n12007_));
  XNOR2_X1   g10987(.A1(new_n12007_), .A2(new_n12005_), .ZN(new_n12008_));
  INV_X1     g10988(.I(\A[808] ), .ZN(new_n12009_));
  NOR2_X1    g10989(.A1(\A[809] ), .A2(\A[810] ), .ZN(new_n12010_));
  NAND2_X1   g10990(.A1(\A[809] ), .A2(\A[810] ), .ZN(new_n12011_));
  AOI21_X1   g10991(.A1(new_n12009_), .A2(new_n12011_), .B(new_n12010_), .ZN(new_n12012_));
  INV_X1     g10992(.I(new_n12012_), .ZN(new_n12013_));
  INV_X1     g10993(.I(\A[805] ), .ZN(new_n12014_));
  NOR2_X1    g10994(.A1(\A[806] ), .A2(\A[807] ), .ZN(new_n12015_));
  NAND2_X1   g10995(.A1(\A[806] ), .A2(\A[807] ), .ZN(new_n12016_));
  AOI21_X1   g10996(.A1(new_n12014_), .A2(new_n12016_), .B(new_n12015_), .ZN(new_n12017_));
  INV_X1     g10997(.I(new_n12017_), .ZN(new_n12018_));
  NOR2_X1    g10998(.A1(new_n12013_), .A2(new_n12018_), .ZN(new_n12019_));
  INV_X1     g10999(.I(new_n12019_), .ZN(new_n12020_));
  INV_X1     g11000(.I(\A[806] ), .ZN(new_n12021_));
  NAND2_X1   g11001(.A1(new_n12021_), .A2(\A[807] ), .ZN(new_n12022_));
  INV_X1     g11002(.I(\A[807] ), .ZN(new_n12023_));
  NAND2_X1   g11003(.A1(new_n12023_), .A2(\A[806] ), .ZN(new_n12024_));
  AOI21_X1   g11004(.A1(new_n12022_), .A2(new_n12024_), .B(new_n12014_), .ZN(new_n12025_));
  INV_X1     g11005(.I(new_n12015_), .ZN(new_n12026_));
  AOI21_X1   g11006(.A1(new_n12026_), .A2(new_n12016_), .B(\A[805] ), .ZN(new_n12027_));
  NOR2_X1    g11007(.A1(new_n12027_), .A2(new_n12025_), .ZN(new_n12028_));
  INV_X1     g11008(.I(\A[809] ), .ZN(new_n12029_));
  NAND2_X1   g11009(.A1(new_n12029_), .A2(\A[810] ), .ZN(new_n12030_));
  INV_X1     g11010(.I(\A[810] ), .ZN(new_n12031_));
  NAND2_X1   g11011(.A1(new_n12031_), .A2(\A[809] ), .ZN(new_n12032_));
  AOI21_X1   g11012(.A1(new_n12030_), .A2(new_n12032_), .B(new_n12009_), .ZN(new_n12033_));
  INV_X1     g11013(.I(new_n12010_), .ZN(new_n12034_));
  AOI21_X1   g11014(.A1(new_n12034_), .A2(new_n12011_), .B(\A[808] ), .ZN(new_n12035_));
  NOR2_X1    g11015(.A1(new_n12035_), .A2(new_n12033_), .ZN(new_n12036_));
  NAND2_X1   g11016(.A1(new_n12028_), .A2(new_n12036_), .ZN(new_n12037_));
  NOR2_X1    g11017(.A1(new_n12037_), .A2(new_n12020_), .ZN(new_n12038_));
  NOR2_X1    g11018(.A1(new_n12023_), .A2(\A[806] ), .ZN(new_n12039_));
  NOR2_X1    g11019(.A1(new_n12021_), .A2(\A[807] ), .ZN(new_n12040_));
  OAI21_X1   g11020(.A1(new_n12039_), .A2(new_n12040_), .B(\A[805] ), .ZN(new_n12041_));
  INV_X1     g11021(.I(new_n12016_), .ZN(new_n12042_));
  OAI21_X1   g11022(.A1(new_n12042_), .A2(new_n12015_), .B(new_n12014_), .ZN(new_n12043_));
  NAND2_X1   g11023(.A1(new_n12041_), .A2(new_n12043_), .ZN(new_n12044_));
  NOR2_X1    g11024(.A1(new_n12031_), .A2(\A[809] ), .ZN(new_n12045_));
  NOR2_X1    g11025(.A1(new_n12029_), .A2(\A[810] ), .ZN(new_n12046_));
  OAI21_X1   g11026(.A1(new_n12045_), .A2(new_n12046_), .B(\A[808] ), .ZN(new_n12047_));
  INV_X1     g11027(.I(new_n12011_), .ZN(new_n12048_));
  OAI21_X1   g11028(.A1(new_n12048_), .A2(new_n12010_), .B(new_n12009_), .ZN(new_n12049_));
  NAND2_X1   g11029(.A1(new_n12047_), .A2(new_n12049_), .ZN(new_n12050_));
  NOR2_X1    g11030(.A1(new_n12044_), .A2(new_n12050_), .ZN(new_n12051_));
  NOR2_X1    g11031(.A1(new_n12028_), .A2(new_n12036_), .ZN(new_n12052_));
  NOR2_X1    g11032(.A1(new_n12052_), .A2(new_n12051_), .ZN(new_n12053_));
  INV_X1     g11033(.I(\A[799] ), .ZN(new_n12054_));
  INV_X1     g11034(.I(\A[800] ), .ZN(new_n12055_));
  NAND2_X1   g11035(.A1(new_n12055_), .A2(\A[801] ), .ZN(new_n12056_));
  INV_X1     g11036(.I(\A[801] ), .ZN(new_n12057_));
  NAND2_X1   g11037(.A1(new_n12057_), .A2(\A[800] ), .ZN(new_n12058_));
  AOI21_X1   g11038(.A1(new_n12056_), .A2(new_n12058_), .B(new_n12054_), .ZN(new_n12059_));
  NOR2_X1    g11039(.A1(\A[800] ), .A2(\A[801] ), .ZN(new_n12060_));
  INV_X1     g11040(.I(new_n12060_), .ZN(new_n12061_));
  NAND2_X1   g11041(.A1(\A[800] ), .A2(\A[801] ), .ZN(new_n12062_));
  AOI21_X1   g11042(.A1(new_n12061_), .A2(new_n12062_), .B(\A[799] ), .ZN(new_n12063_));
  NOR2_X1    g11043(.A1(new_n12063_), .A2(new_n12059_), .ZN(new_n12064_));
  INV_X1     g11044(.I(\A[802] ), .ZN(new_n12065_));
  INV_X1     g11045(.I(\A[803] ), .ZN(new_n12066_));
  NAND2_X1   g11046(.A1(new_n12066_), .A2(\A[804] ), .ZN(new_n12067_));
  INV_X1     g11047(.I(\A[804] ), .ZN(new_n12068_));
  NAND2_X1   g11048(.A1(new_n12068_), .A2(\A[803] ), .ZN(new_n12069_));
  AOI21_X1   g11049(.A1(new_n12067_), .A2(new_n12069_), .B(new_n12065_), .ZN(new_n12070_));
  NOR2_X1    g11050(.A1(\A[803] ), .A2(\A[804] ), .ZN(new_n12071_));
  INV_X1     g11051(.I(new_n12071_), .ZN(new_n12072_));
  NAND2_X1   g11052(.A1(\A[803] ), .A2(\A[804] ), .ZN(new_n12073_));
  AOI21_X1   g11053(.A1(new_n12072_), .A2(new_n12073_), .B(\A[802] ), .ZN(new_n12074_));
  NOR2_X1    g11054(.A1(new_n12074_), .A2(new_n12070_), .ZN(new_n12075_));
  AOI21_X1   g11055(.A1(new_n12065_), .A2(new_n12073_), .B(new_n12071_), .ZN(new_n12076_));
  INV_X1     g11056(.I(new_n12076_), .ZN(new_n12077_));
  AOI21_X1   g11057(.A1(new_n12054_), .A2(new_n12062_), .B(new_n12060_), .ZN(new_n12078_));
  INV_X1     g11058(.I(new_n12078_), .ZN(new_n12079_));
  NOR2_X1    g11059(.A1(new_n12077_), .A2(new_n12079_), .ZN(new_n12080_));
  NAND2_X1   g11060(.A1(new_n12053_), .A2(new_n12038_), .ZN(new_n12081_));
  NAND2_X1   g11061(.A1(new_n12008_), .A2(new_n12081_), .ZN(new_n12082_));
  OAI21_X1   g11062(.A1(new_n12003_), .A2(new_n11998_), .B(new_n12082_), .ZN(new_n12083_));
  XOR2_X1    g11063(.A1(new_n12007_), .A2(new_n12005_), .Z(new_n12084_));
  INV_X1     g11064(.I(new_n12081_), .ZN(new_n12085_));
  NOR2_X1    g11065(.A1(new_n12084_), .A2(new_n12085_), .ZN(new_n12086_));
  NAND3_X1   g11066(.A1(new_n11989_), .A2(new_n11993_), .A3(new_n12086_), .ZN(new_n12087_));
  NAND2_X1   g11067(.A1(new_n12037_), .A2(new_n12017_), .ZN(new_n12088_));
  NAND2_X1   g11068(.A1(new_n12051_), .A2(new_n12018_), .ZN(new_n12089_));
  AOI21_X1   g11069(.A1(new_n12089_), .A2(new_n12088_), .B(new_n12013_), .ZN(new_n12090_));
  NOR2_X1    g11070(.A1(new_n12051_), .A2(new_n12018_), .ZN(new_n12091_));
  NOR2_X1    g11071(.A1(new_n12037_), .A2(new_n12017_), .ZN(new_n12092_));
  NOR3_X1    g11072(.A1(new_n12091_), .A2(new_n12092_), .A3(new_n12012_), .ZN(new_n12093_));
  NOR2_X1    g11073(.A1(new_n12090_), .A2(new_n12093_), .ZN(new_n12094_));
  INV_X1     g11074(.I(new_n12038_), .ZN(new_n12095_));
  INV_X1     g11075(.I(new_n12053_), .ZN(new_n12096_));
  NOR4_X1    g11076(.A1(new_n12059_), .A2(new_n12063_), .A3(new_n12074_), .A4(new_n12070_), .ZN(new_n12097_));
  NOR2_X1    g11077(.A1(new_n12064_), .A2(new_n12075_), .ZN(new_n12098_));
  NOR4_X1    g11078(.A1(new_n12096_), .A2(new_n12095_), .A3(new_n12097_), .A4(new_n12098_), .ZN(new_n12099_));
  NAND2_X1   g11079(.A1(new_n12064_), .A2(new_n12075_), .ZN(new_n12100_));
  INV_X1     g11080(.I(new_n12080_), .ZN(new_n12101_));
  NOR2_X1    g11081(.A1(new_n12100_), .A2(new_n12101_), .ZN(new_n12102_));
  NAND2_X1   g11082(.A1(new_n12028_), .A2(new_n12050_), .ZN(new_n12103_));
  NAND2_X1   g11083(.A1(new_n12036_), .A2(new_n12044_), .ZN(new_n12104_));
  AOI21_X1   g11084(.A1(new_n12103_), .A2(new_n12104_), .B(new_n12020_), .ZN(new_n12105_));
  INV_X1     g11085(.I(new_n12105_), .ZN(new_n12106_));
  NAND2_X1   g11086(.A1(new_n12106_), .A2(new_n12102_), .ZN(new_n12107_));
  AOI21_X1   g11087(.A1(new_n12094_), .A2(new_n12099_), .B(new_n12107_), .ZN(new_n12108_));
  NAND2_X1   g11088(.A1(new_n12100_), .A2(new_n12078_), .ZN(new_n12109_));
  NAND2_X1   g11089(.A1(new_n12097_), .A2(new_n12079_), .ZN(new_n12110_));
  AOI21_X1   g11090(.A1(new_n12109_), .A2(new_n12110_), .B(new_n12077_), .ZN(new_n12111_));
  NOR2_X1    g11091(.A1(new_n12097_), .A2(new_n12079_), .ZN(new_n12112_));
  NOR2_X1    g11092(.A1(new_n12100_), .A2(new_n12078_), .ZN(new_n12113_));
  NOR3_X1    g11093(.A1(new_n12113_), .A2(new_n12076_), .A3(new_n12112_), .ZN(new_n12114_));
  NOR2_X1    g11094(.A1(new_n12114_), .A2(new_n12111_), .ZN(new_n12115_));
  INV_X1     g11095(.I(new_n12115_), .ZN(new_n12116_));
  NAND2_X1   g11096(.A1(new_n12108_), .A2(new_n12116_), .ZN(new_n12117_));
  NOR2_X1    g11097(.A1(new_n12098_), .A2(new_n12097_), .ZN(new_n12118_));
  NAND4_X1   g11098(.A1(new_n12038_), .A2(new_n12053_), .A3(new_n12102_), .A4(new_n12118_), .ZN(new_n12119_));
  NAND2_X1   g11099(.A1(new_n12116_), .A2(new_n12119_), .ZN(new_n12120_));
  INV_X1     g11100(.I(new_n12119_), .ZN(new_n12121_));
  NOR3_X1    g11101(.A1(new_n12090_), .A2(new_n12093_), .A3(new_n12105_), .ZN(new_n12122_));
  AOI21_X1   g11102(.A1(new_n12115_), .A2(new_n12121_), .B(new_n12122_), .ZN(new_n12123_));
  OAI21_X1   g11103(.A1(new_n12091_), .A2(new_n12092_), .B(new_n12012_), .ZN(new_n12124_));
  NAND3_X1   g11104(.A1(new_n12089_), .A2(new_n12088_), .A3(new_n12013_), .ZN(new_n12125_));
  NAND3_X1   g11105(.A1(new_n12124_), .A2(new_n12125_), .A3(new_n12106_), .ZN(new_n12126_));
  NOR3_X1    g11106(.A1(new_n12116_), .A2(new_n12119_), .A3(new_n12126_), .ZN(new_n12127_));
  OAI21_X1   g11107(.A1(new_n12127_), .A2(new_n12123_), .B(new_n12120_), .ZN(new_n12128_));
  NAND2_X1   g11108(.A1(new_n12128_), .A2(new_n12117_), .ZN(new_n12129_));
  AOI22_X1   g11109(.A1(new_n12129_), .A2(new_n11994_), .B1(new_n12083_), .B2(new_n12087_), .ZN(new_n12130_));
  NOR2_X1    g11110(.A1(new_n12002_), .A2(new_n11924_), .ZN(new_n12131_));
  NOR2_X1    g11111(.A1(new_n11928_), .A2(new_n11933_), .ZN(new_n12132_));
  OAI21_X1   g11112(.A1(new_n11950_), .A2(new_n12132_), .B(new_n11980_), .ZN(new_n12133_));
  NOR2_X1    g11113(.A1(new_n11896_), .A2(new_n11901_), .ZN(new_n12134_));
  OAI21_X1   g11114(.A1(new_n11974_), .A2(new_n12134_), .B(new_n11975_), .ZN(new_n12135_));
  XNOR2_X1   g11115(.A1(new_n12133_), .A2(new_n12135_), .ZN(new_n12136_));
  INV_X1     g11116(.I(new_n12136_), .ZN(new_n12137_));
  NOR3_X1    g11117(.A1(new_n12131_), .A2(new_n12001_), .A3(new_n12137_), .ZN(new_n12138_));
  AOI21_X1   g11118(.A1(new_n12126_), .A2(new_n12121_), .B(new_n12115_), .ZN(new_n12139_));
  NOR2_X1    g11119(.A1(new_n12012_), .A2(new_n12017_), .ZN(new_n12140_));
  OAI21_X1   g11120(.A1(new_n12037_), .A2(new_n12140_), .B(new_n12020_), .ZN(new_n12141_));
  NOR2_X1    g11121(.A1(new_n12076_), .A2(new_n12078_), .ZN(new_n12142_));
  OAI21_X1   g11122(.A1(new_n12100_), .A2(new_n12142_), .B(new_n12101_), .ZN(new_n12143_));
  XOR2_X1    g11123(.A1(new_n12141_), .A2(new_n12143_), .Z(new_n12144_));
  NOR3_X1    g11124(.A1(new_n12139_), .A2(new_n12108_), .A3(new_n12144_), .ZN(new_n12145_));
  XOR2_X1    g11125(.A1(new_n12138_), .A2(new_n12145_), .Z(new_n12146_));
  NAND2_X1   g11126(.A1(new_n12146_), .A2(new_n12130_), .ZN(new_n12147_));
  NOR2_X1    g11127(.A1(new_n12003_), .A2(new_n11998_), .ZN(new_n12148_));
  AOI21_X1   g11128(.A1(new_n11993_), .A2(new_n11989_), .B(new_n12086_), .ZN(new_n12149_));
  NOR3_X1    g11129(.A1(new_n12003_), .A2(new_n12082_), .A3(new_n11998_), .ZN(new_n12150_));
  OAI21_X1   g11130(.A1(new_n12116_), .A2(new_n12119_), .B(new_n12126_), .ZN(new_n12151_));
  NAND3_X1   g11131(.A1(new_n12122_), .A2(new_n12121_), .A3(new_n12115_), .ZN(new_n12152_));
  NAND2_X1   g11132(.A1(new_n12151_), .A2(new_n12152_), .ZN(new_n12153_));
  AOI22_X1   g11133(.A1(new_n12153_), .A2(new_n12120_), .B1(new_n12108_), .B2(new_n12116_), .ZN(new_n12154_));
  OAI22_X1   g11134(.A1(new_n12154_), .A2(new_n12148_), .B1(new_n12150_), .B2(new_n12149_), .ZN(new_n12155_));
  NAND2_X1   g11135(.A1(new_n11992_), .A2(new_n11995_), .ZN(new_n12156_));
  NAND3_X1   g11136(.A1(new_n12156_), .A2(new_n11991_), .A3(new_n12136_), .ZN(new_n12157_));
  INV_X1     g11137(.I(new_n12145_), .ZN(new_n12158_));
  NAND2_X1   g11138(.A1(new_n12158_), .A2(new_n12157_), .ZN(new_n12159_));
  NAND2_X1   g11139(.A1(new_n12138_), .A2(new_n12145_), .ZN(new_n12160_));
  NAND2_X1   g11140(.A1(new_n12159_), .A2(new_n12160_), .ZN(new_n12161_));
  NAND2_X1   g11141(.A1(new_n12155_), .A2(new_n12161_), .ZN(new_n12162_));
  NAND2_X1   g11142(.A1(new_n12147_), .A2(new_n12162_), .ZN(new_n12163_));
  INV_X1     g11143(.I(\A[838] ), .ZN(new_n12164_));
  NOR2_X1    g11144(.A1(\A[839] ), .A2(\A[840] ), .ZN(new_n12165_));
  NAND2_X1   g11145(.A1(\A[839] ), .A2(\A[840] ), .ZN(new_n12166_));
  AOI21_X1   g11146(.A1(new_n12164_), .A2(new_n12166_), .B(new_n12165_), .ZN(new_n12167_));
  INV_X1     g11147(.I(\A[835] ), .ZN(new_n12168_));
  NOR2_X1    g11148(.A1(\A[836] ), .A2(\A[837] ), .ZN(new_n12169_));
  NAND2_X1   g11149(.A1(\A[836] ), .A2(\A[837] ), .ZN(new_n12170_));
  AOI21_X1   g11150(.A1(new_n12168_), .A2(new_n12170_), .B(new_n12169_), .ZN(new_n12171_));
  INV_X1     g11151(.I(new_n12171_), .ZN(new_n12172_));
  INV_X1     g11152(.I(\A[836] ), .ZN(new_n12173_));
  NAND2_X1   g11153(.A1(new_n12173_), .A2(\A[837] ), .ZN(new_n12174_));
  INV_X1     g11154(.I(\A[837] ), .ZN(new_n12175_));
  NAND2_X1   g11155(.A1(new_n12175_), .A2(\A[836] ), .ZN(new_n12176_));
  AOI21_X1   g11156(.A1(new_n12174_), .A2(new_n12176_), .B(new_n12168_), .ZN(new_n12177_));
  INV_X1     g11157(.I(new_n12169_), .ZN(new_n12178_));
  AOI21_X1   g11158(.A1(new_n12178_), .A2(new_n12170_), .B(\A[835] ), .ZN(new_n12179_));
  INV_X1     g11159(.I(\A[839] ), .ZN(new_n12180_));
  NAND2_X1   g11160(.A1(new_n12180_), .A2(\A[840] ), .ZN(new_n12181_));
  INV_X1     g11161(.I(\A[840] ), .ZN(new_n12182_));
  NAND2_X1   g11162(.A1(new_n12182_), .A2(\A[839] ), .ZN(new_n12183_));
  AOI21_X1   g11163(.A1(new_n12181_), .A2(new_n12183_), .B(new_n12164_), .ZN(new_n12184_));
  INV_X1     g11164(.I(new_n12165_), .ZN(new_n12185_));
  AOI21_X1   g11165(.A1(new_n12185_), .A2(new_n12166_), .B(\A[838] ), .ZN(new_n12186_));
  NOR4_X1    g11166(.A1(new_n12177_), .A2(new_n12179_), .A3(new_n12186_), .A4(new_n12184_), .ZN(new_n12187_));
  NOR2_X1    g11167(.A1(new_n12187_), .A2(new_n12172_), .ZN(new_n12188_));
  NAND2_X1   g11168(.A1(new_n12187_), .A2(new_n12172_), .ZN(new_n12189_));
  INV_X1     g11169(.I(new_n12189_), .ZN(new_n12190_));
  OAI21_X1   g11170(.A1(new_n12190_), .A2(new_n12188_), .B(new_n12167_), .ZN(new_n12191_));
  INV_X1     g11171(.I(new_n12167_), .ZN(new_n12192_));
  INV_X1     g11172(.I(new_n12188_), .ZN(new_n12193_));
  NAND3_X1   g11173(.A1(new_n12193_), .A2(new_n12192_), .A3(new_n12189_), .ZN(new_n12194_));
  NAND2_X1   g11174(.A1(new_n12191_), .A2(new_n12194_), .ZN(new_n12195_));
  INV_X1     g11175(.I(new_n12195_), .ZN(new_n12196_));
  INV_X1     g11176(.I(\A[844] ), .ZN(new_n12197_));
  NOR2_X1    g11177(.A1(\A[845] ), .A2(\A[846] ), .ZN(new_n12198_));
  NAND2_X1   g11178(.A1(\A[845] ), .A2(\A[846] ), .ZN(new_n12199_));
  AOI21_X1   g11179(.A1(new_n12197_), .A2(new_n12199_), .B(new_n12198_), .ZN(new_n12200_));
  INV_X1     g11180(.I(new_n12200_), .ZN(new_n12201_));
  INV_X1     g11181(.I(\A[841] ), .ZN(new_n12202_));
  NOR2_X1    g11182(.A1(\A[842] ), .A2(\A[843] ), .ZN(new_n12203_));
  NAND2_X1   g11183(.A1(\A[842] ), .A2(\A[843] ), .ZN(new_n12204_));
  AOI21_X1   g11184(.A1(new_n12202_), .A2(new_n12204_), .B(new_n12203_), .ZN(new_n12205_));
  INV_X1     g11185(.I(\A[842] ), .ZN(new_n12206_));
  NAND2_X1   g11186(.A1(new_n12206_), .A2(\A[843] ), .ZN(new_n12207_));
  INV_X1     g11187(.I(\A[843] ), .ZN(new_n12208_));
  NAND2_X1   g11188(.A1(new_n12208_), .A2(\A[842] ), .ZN(new_n12209_));
  AOI21_X1   g11189(.A1(new_n12207_), .A2(new_n12209_), .B(new_n12202_), .ZN(new_n12210_));
  INV_X1     g11190(.I(new_n12203_), .ZN(new_n12211_));
  AOI21_X1   g11191(.A1(new_n12211_), .A2(new_n12204_), .B(\A[841] ), .ZN(new_n12212_));
  NOR2_X1    g11192(.A1(new_n12212_), .A2(new_n12210_), .ZN(new_n12213_));
  INV_X1     g11193(.I(\A[845] ), .ZN(new_n12214_));
  NAND2_X1   g11194(.A1(new_n12214_), .A2(\A[846] ), .ZN(new_n12215_));
  INV_X1     g11195(.I(\A[846] ), .ZN(new_n12216_));
  NAND2_X1   g11196(.A1(new_n12216_), .A2(\A[845] ), .ZN(new_n12217_));
  AOI21_X1   g11197(.A1(new_n12215_), .A2(new_n12217_), .B(new_n12197_), .ZN(new_n12218_));
  INV_X1     g11198(.I(new_n12198_), .ZN(new_n12219_));
  AOI21_X1   g11199(.A1(new_n12219_), .A2(new_n12199_), .B(\A[844] ), .ZN(new_n12220_));
  NOR2_X1    g11200(.A1(new_n12220_), .A2(new_n12218_), .ZN(new_n12221_));
  NAND2_X1   g11201(.A1(new_n12213_), .A2(new_n12221_), .ZN(new_n12222_));
  NAND2_X1   g11202(.A1(new_n12222_), .A2(new_n12205_), .ZN(new_n12223_));
  INV_X1     g11203(.I(new_n12205_), .ZN(new_n12224_));
  NOR2_X1    g11204(.A1(new_n12208_), .A2(\A[842] ), .ZN(new_n12225_));
  NOR2_X1    g11205(.A1(new_n12206_), .A2(\A[843] ), .ZN(new_n12226_));
  OAI21_X1   g11206(.A1(new_n12225_), .A2(new_n12226_), .B(\A[841] ), .ZN(new_n12227_));
  INV_X1     g11207(.I(new_n12204_), .ZN(new_n12228_));
  OAI21_X1   g11208(.A1(new_n12228_), .A2(new_n12203_), .B(new_n12202_), .ZN(new_n12229_));
  NAND2_X1   g11209(.A1(new_n12227_), .A2(new_n12229_), .ZN(new_n12230_));
  NOR2_X1    g11210(.A1(new_n12216_), .A2(\A[845] ), .ZN(new_n12231_));
  NOR2_X1    g11211(.A1(new_n12214_), .A2(\A[846] ), .ZN(new_n12232_));
  OAI21_X1   g11212(.A1(new_n12231_), .A2(new_n12232_), .B(\A[844] ), .ZN(new_n12233_));
  INV_X1     g11213(.I(new_n12199_), .ZN(new_n12234_));
  OAI21_X1   g11214(.A1(new_n12234_), .A2(new_n12198_), .B(new_n12197_), .ZN(new_n12235_));
  NAND2_X1   g11215(.A1(new_n12233_), .A2(new_n12235_), .ZN(new_n12236_));
  NOR2_X1    g11216(.A1(new_n12230_), .A2(new_n12236_), .ZN(new_n12237_));
  NAND2_X1   g11217(.A1(new_n12237_), .A2(new_n12224_), .ZN(new_n12238_));
  AOI21_X1   g11218(.A1(new_n12238_), .A2(new_n12223_), .B(new_n12201_), .ZN(new_n12239_));
  NOR2_X1    g11219(.A1(new_n12237_), .A2(new_n12224_), .ZN(new_n12240_));
  NOR2_X1    g11220(.A1(new_n12222_), .A2(new_n12205_), .ZN(new_n12241_));
  NOR3_X1    g11221(.A1(new_n12240_), .A2(new_n12241_), .A3(new_n12200_), .ZN(new_n12242_));
  NOR2_X1    g11222(.A1(new_n12239_), .A2(new_n12242_), .ZN(new_n12243_));
  NOR2_X1    g11223(.A1(new_n12179_), .A2(new_n12177_), .ZN(new_n12244_));
  NOR2_X1    g11224(.A1(new_n12186_), .A2(new_n12184_), .ZN(new_n12245_));
  NAND2_X1   g11225(.A1(new_n12244_), .A2(new_n12245_), .ZN(new_n12246_));
  NAND2_X1   g11226(.A1(new_n12167_), .A2(new_n12171_), .ZN(new_n12247_));
  NOR2_X1    g11227(.A1(new_n12213_), .A2(new_n12221_), .ZN(new_n12248_));
  NOR4_X1    g11228(.A1(new_n12237_), .A2(new_n12248_), .A3(new_n12246_), .A4(new_n12247_), .ZN(new_n12249_));
  NOR2_X1    g11229(.A1(new_n12244_), .A2(new_n12245_), .ZN(new_n12250_));
  NOR2_X1    g11230(.A1(new_n12250_), .A2(new_n12187_), .ZN(new_n12251_));
  NAND2_X1   g11231(.A1(new_n12200_), .A2(new_n12205_), .ZN(new_n12252_));
  NOR3_X1    g11232(.A1(new_n12230_), .A2(new_n12236_), .A3(new_n12252_), .ZN(new_n12253_));
  NAND3_X1   g11233(.A1(new_n12249_), .A2(new_n12251_), .A3(new_n12253_), .ZN(new_n12254_));
  NOR2_X1    g11234(.A1(new_n12243_), .A2(new_n12254_), .ZN(new_n12255_));
  OAI21_X1   g11235(.A1(new_n12240_), .A2(new_n12241_), .B(new_n12200_), .ZN(new_n12256_));
  NAND3_X1   g11236(.A1(new_n12238_), .A2(new_n12223_), .A3(new_n12201_), .ZN(new_n12257_));
  NAND2_X1   g11237(.A1(new_n12256_), .A2(new_n12257_), .ZN(new_n12258_));
  INV_X1     g11238(.I(new_n12254_), .ZN(new_n12259_));
  NOR2_X1    g11239(.A1(new_n12259_), .A2(new_n12258_), .ZN(new_n12260_));
  OAI21_X1   g11240(.A1(new_n12260_), .A2(new_n12255_), .B(new_n12196_), .ZN(new_n12261_));
  NAND2_X1   g11241(.A1(new_n12249_), .A2(new_n12251_), .ZN(new_n12262_));
  OAI22_X1   g11242(.A1(new_n12258_), .A2(new_n12262_), .B1(new_n12248_), .B2(new_n12252_), .ZN(new_n12263_));
  NAND2_X1   g11243(.A1(new_n12259_), .A2(new_n12243_), .ZN(new_n12264_));
  NAND3_X1   g11244(.A1(new_n12263_), .A2(new_n12264_), .A3(new_n12196_), .ZN(new_n12265_));
  NAND2_X1   g11245(.A1(new_n12265_), .A2(new_n12261_), .ZN(new_n12266_));
  NAND2_X1   g11246(.A1(new_n12259_), .A2(new_n12258_), .ZN(new_n12267_));
  NAND2_X1   g11247(.A1(new_n12243_), .A2(new_n12254_), .ZN(new_n12268_));
  AOI21_X1   g11248(.A1(new_n12267_), .A2(new_n12268_), .B(new_n12195_), .ZN(new_n12269_));
  INV_X1     g11249(.I(new_n12262_), .ZN(new_n12270_));
  NOR2_X1    g11250(.A1(new_n12248_), .A2(new_n12252_), .ZN(new_n12271_));
  AOI21_X1   g11251(.A1(new_n12243_), .A2(new_n12270_), .B(new_n12271_), .ZN(new_n12272_));
  NOR2_X1    g11252(.A1(new_n12258_), .A2(new_n12254_), .ZN(new_n12273_));
  NOR3_X1    g11253(.A1(new_n12272_), .A2(new_n12273_), .A3(new_n12195_), .ZN(new_n12274_));
  NOR2_X1    g11254(.A1(new_n12248_), .A2(new_n12237_), .ZN(new_n12275_));
  NAND2_X1   g11255(.A1(new_n12275_), .A2(new_n12253_), .ZN(new_n12276_));
  NOR2_X1    g11256(.A1(new_n12246_), .A2(new_n12247_), .ZN(new_n12277_));
  NAND2_X1   g11257(.A1(new_n12251_), .A2(new_n12277_), .ZN(new_n12278_));
  XNOR2_X1   g11258(.A1(new_n12278_), .A2(new_n12276_), .ZN(new_n12279_));
  INV_X1     g11259(.I(\A[831] ), .ZN(new_n12280_));
  NOR2_X1    g11260(.A1(new_n12280_), .A2(\A[830] ), .ZN(new_n12281_));
  INV_X1     g11261(.I(\A[830] ), .ZN(new_n12282_));
  NOR2_X1    g11262(.A1(new_n12282_), .A2(\A[831] ), .ZN(new_n12283_));
  OAI21_X1   g11263(.A1(new_n12281_), .A2(new_n12283_), .B(\A[829] ), .ZN(new_n12284_));
  INV_X1     g11264(.I(\A[829] ), .ZN(new_n12285_));
  NOR2_X1    g11265(.A1(\A[830] ), .A2(\A[831] ), .ZN(new_n12286_));
  NAND2_X1   g11266(.A1(\A[830] ), .A2(\A[831] ), .ZN(new_n12287_));
  INV_X1     g11267(.I(new_n12287_), .ZN(new_n12288_));
  OAI21_X1   g11268(.A1(new_n12288_), .A2(new_n12286_), .B(new_n12285_), .ZN(new_n12289_));
  NAND2_X1   g11269(.A1(new_n12284_), .A2(new_n12289_), .ZN(new_n12290_));
  INV_X1     g11270(.I(\A[834] ), .ZN(new_n12291_));
  NOR2_X1    g11271(.A1(new_n12291_), .A2(\A[833] ), .ZN(new_n12292_));
  INV_X1     g11272(.I(\A[833] ), .ZN(new_n12293_));
  NOR2_X1    g11273(.A1(new_n12293_), .A2(\A[834] ), .ZN(new_n12294_));
  OAI21_X1   g11274(.A1(new_n12292_), .A2(new_n12294_), .B(\A[832] ), .ZN(new_n12295_));
  INV_X1     g11275(.I(\A[832] ), .ZN(new_n12296_));
  NOR2_X1    g11276(.A1(\A[833] ), .A2(\A[834] ), .ZN(new_n12297_));
  NAND2_X1   g11277(.A1(\A[833] ), .A2(\A[834] ), .ZN(new_n12298_));
  INV_X1     g11278(.I(new_n12298_), .ZN(new_n12299_));
  OAI21_X1   g11279(.A1(new_n12299_), .A2(new_n12297_), .B(new_n12296_), .ZN(new_n12300_));
  NAND2_X1   g11280(.A1(new_n12295_), .A2(new_n12300_), .ZN(new_n12301_));
  NOR2_X1    g11281(.A1(new_n12290_), .A2(new_n12301_), .ZN(new_n12302_));
  NAND2_X1   g11282(.A1(new_n12282_), .A2(\A[831] ), .ZN(new_n12303_));
  NAND2_X1   g11283(.A1(new_n12280_), .A2(\A[830] ), .ZN(new_n12304_));
  AOI21_X1   g11284(.A1(new_n12303_), .A2(new_n12304_), .B(new_n12285_), .ZN(new_n12305_));
  INV_X1     g11285(.I(new_n12286_), .ZN(new_n12306_));
  AOI21_X1   g11286(.A1(new_n12306_), .A2(new_n12287_), .B(\A[829] ), .ZN(new_n12307_));
  NOR2_X1    g11287(.A1(new_n12307_), .A2(new_n12305_), .ZN(new_n12308_));
  NAND2_X1   g11288(.A1(new_n12293_), .A2(\A[834] ), .ZN(new_n12309_));
  NAND2_X1   g11289(.A1(new_n12291_), .A2(\A[833] ), .ZN(new_n12310_));
  AOI21_X1   g11290(.A1(new_n12309_), .A2(new_n12310_), .B(new_n12296_), .ZN(new_n12311_));
  INV_X1     g11291(.I(new_n12297_), .ZN(new_n12312_));
  AOI21_X1   g11292(.A1(new_n12312_), .A2(new_n12298_), .B(\A[832] ), .ZN(new_n12313_));
  NOR2_X1    g11293(.A1(new_n12313_), .A2(new_n12311_), .ZN(new_n12314_));
  NOR2_X1    g11294(.A1(new_n12308_), .A2(new_n12314_), .ZN(new_n12315_));
  NOR2_X1    g11295(.A1(new_n12315_), .A2(new_n12302_), .ZN(new_n12316_));
  AOI21_X1   g11296(.A1(new_n12296_), .A2(new_n12298_), .B(new_n12297_), .ZN(new_n12317_));
  AOI21_X1   g11297(.A1(new_n12285_), .A2(new_n12287_), .B(new_n12286_), .ZN(new_n12318_));
  NAND2_X1   g11298(.A1(new_n12317_), .A2(new_n12318_), .ZN(new_n12319_));
  INV_X1     g11299(.I(new_n12319_), .ZN(new_n12320_));
  NAND3_X1   g11300(.A1(new_n12320_), .A2(new_n12308_), .A3(new_n12314_), .ZN(new_n12321_));
  INV_X1     g11301(.I(new_n12321_), .ZN(new_n12322_));
  INV_X1     g11302(.I(\A[826] ), .ZN(new_n12323_));
  NOR2_X1    g11303(.A1(\A[827] ), .A2(\A[828] ), .ZN(new_n12324_));
  NAND2_X1   g11304(.A1(\A[827] ), .A2(\A[828] ), .ZN(new_n12325_));
  AOI21_X1   g11305(.A1(new_n12323_), .A2(new_n12325_), .B(new_n12324_), .ZN(new_n12326_));
  INV_X1     g11306(.I(new_n12326_), .ZN(new_n12327_));
  INV_X1     g11307(.I(\A[823] ), .ZN(new_n12328_));
  NOR2_X1    g11308(.A1(\A[824] ), .A2(\A[825] ), .ZN(new_n12329_));
  NAND2_X1   g11309(.A1(\A[824] ), .A2(\A[825] ), .ZN(new_n12330_));
  AOI21_X1   g11310(.A1(new_n12328_), .A2(new_n12330_), .B(new_n12329_), .ZN(new_n12331_));
  INV_X1     g11311(.I(new_n12331_), .ZN(new_n12332_));
  NOR2_X1    g11312(.A1(new_n12327_), .A2(new_n12332_), .ZN(new_n12333_));
  INV_X1     g11313(.I(\A[824] ), .ZN(new_n12334_));
  NAND2_X1   g11314(.A1(new_n12334_), .A2(\A[825] ), .ZN(new_n12335_));
  INV_X1     g11315(.I(\A[825] ), .ZN(new_n12336_));
  NAND2_X1   g11316(.A1(new_n12336_), .A2(\A[824] ), .ZN(new_n12337_));
  AOI21_X1   g11317(.A1(new_n12335_), .A2(new_n12337_), .B(new_n12328_), .ZN(new_n12338_));
  INV_X1     g11318(.I(new_n12329_), .ZN(new_n12339_));
  AOI21_X1   g11319(.A1(new_n12339_), .A2(new_n12330_), .B(\A[823] ), .ZN(new_n12340_));
  NOR2_X1    g11320(.A1(new_n12340_), .A2(new_n12338_), .ZN(new_n12341_));
  INV_X1     g11321(.I(\A[827] ), .ZN(new_n12342_));
  NAND2_X1   g11322(.A1(new_n12342_), .A2(\A[828] ), .ZN(new_n12343_));
  INV_X1     g11323(.I(\A[828] ), .ZN(new_n12344_));
  NAND2_X1   g11324(.A1(new_n12344_), .A2(\A[827] ), .ZN(new_n12345_));
  AOI21_X1   g11325(.A1(new_n12343_), .A2(new_n12345_), .B(new_n12323_), .ZN(new_n12346_));
  INV_X1     g11326(.I(new_n12324_), .ZN(new_n12347_));
  AOI21_X1   g11327(.A1(new_n12347_), .A2(new_n12325_), .B(\A[826] ), .ZN(new_n12348_));
  NOR2_X1    g11328(.A1(new_n12348_), .A2(new_n12346_), .ZN(new_n12349_));
  NAND2_X1   g11329(.A1(new_n12316_), .A2(new_n12322_), .ZN(new_n12350_));
  NAND2_X1   g11330(.A1(new_n12279_), .A2(new_n12350_), .ZN(new_n12351_));
  OAI21_X1   g11331(.A1(new_n12274_), .A2(new_n12269_), .B(new_n12351_), .ZN(new_n12352_));
  XOR2_X1    g11332(.A1(new_n12278_), .A2(new_n12276_), .Z(new_n12353_));
  INV_X1     g11333(.I(new_n12350_), .ZN(new_n12354_));
  NOR2_X1    g11334(.A1(new_n12353_), .A2(new_n12354_), .ZN(new_n12355_));
  NAND3_X1   g11335(.A1(new_n12261_), .A2(new_n12265_), .A3(new_n12355_), .ZN(new_n12356_));
  INV_X1     g11336(.I(new_n12318_), .ZN(new_n12357_));
  NOR2_X1    g11337(.A1(new_n12302_), .A2(new_n12357_), .ZN(new_n12358_));
  NAND2_X1   g11338(.A1(new_n12308_), .A2(new_n12314_), .ZN(new_n12359_));
  NOR2_X1    g11339(.A1(new_n12359_), .A2(new_n12318_), .ZN(new_n12360_));
  OAI21_X1   g11340(.A1(new_n12358_), .A2(new_n12360_), .B(new_n12317_), .ZN(new_n12361_));
  INV_X1     g11341(.I(new_n12317_), .ZN(new_n12362_));
  NAND2_X1   g11342(.A1(new_n12359_), .A2(new_n12318_), .ZN(new_n12363_));
  NAND2_X1   g11343(.A1(new_n12302_), .A2(new_n12357_), .ZN(new_n12364_));
  NAND3_X1   g11344(.A1(new_n12364_), .A2(new_n12363_), .A3(new_n12362_), .ZN(new_n12365_));
  NAND2_X1   g11345(.A1(new_n12361_), .A2(new_n12365_), .ZN(new_n12366_));
  NOR4_X1    g11346(.A1(new_n12338_), .A2(new_n12340_), .A3(new_n12348_), .A4(new_n12346_), .ZN(new_n12367_));
  NOR2_X1    g11347(.A1(new_n12341_), .A2(new_n12349_), .ZN(new_n12368_));
  NOR2_X1    g11348(.A1(new_n12368_), .A2(new_n12367_), .ZN(new_n12369_));
  INV_X1     g11349(.I(new_n12333_), .ZN(new_n12370_));
  NAND2_X1   g11350(.A1(new_n12341_), .A2(new_n12349_), .ZN(new_n12371_));
  NOR4_X1    g11351(.A1(new_n12302_), .A2(new_n12315_), .A3(new_n12371_), .A4(new_n12370_), .ZN(new_n12372_));
  NAND2_X1   g11352(.A1(new_n12372_), .A2(new_n12369_), .ZN(new_n12373_));
  OAI21_X1   g11353(.A1(new_n12308_), .A2(new_n12314_), .B(new_n12320_), .ZN(new_n12374_));
  OAI21_X1   g11354(.A1(new_n12366_), .A2(new_n12373_), .B(new_n12374_), .ZN(new_n12375_));
  NAND2_X1   g11355(.A1(new_n12371_), .A2(new_n12331_), .ZN(new_n12376_));
  NAND2_X1   g11356(.A1(new_n12367_), .A2(new_n12332_), .ZN(new_n12377_));
  AOI21_X1   g11357(.A1(new_n12376_), .A2(new_n12377_), .B(new_n12327_), .ZN(new_n12378_));
  NOR2_X1    g11358(.A1(new_n12367_), .A2(new_n12332_), .ZN(new_n12379_));
  NOR2_X1    g11359(.A1(new_n12371_), .A2(new_n12331_), .ZN(new_n12380_));
  NOR3_X1    g11360(.A1(new_n12380_), .A2(new_n12326_), .A3(new_n12379_), .ZN(new_n12381_));
  NOR2_X1    g11361(.A1(new_n12381_), .A2(new_n12378_), .ZN(new_n12382_));
  NOR3_X1    g11362(.A1(new_n12321_), .A2(new_n12368_), .A3(new_n12367_), .ZN(new_n12383_));
  AND2_X2    g11363(.A1(new_n12372_), .A2(new_n12383_), .Z(new_n12384_));
  NOR2_X1    g11364(.A1(new_n12384_), .A2(new_n12382_), .ZN(new_n12385_));
  AOI21_X1   g11365(.A1(new_n12382_), .A2(new_n12384_), .B(new_n12366_), .ZN(new_n12386_));
  AOI21_X1   g11366(.A1(new_n12364_), .A2(new_n12363_), .B(new_n12362_), .ZN(new_n12387_));
  NOR3_X1    g11367(.A1(new_n12358_), .A2(new_n12360_), .A3(new_n12317_), .ZN(new_n12388_));
  NOR2_X1    g11368(.A1(new_n12387_), .A2(new_n12388_), .ZN(new_n12389_));
  OAI21_X1   g11369(.A1(new_n12380_), .A2(new_n12379_), .B(new_n12326_), .ZN(new_n12390_));
  NAND3_X1   g11370(.A1(new_n12376_), .A2(new_n12327_), .A3(new_n12377_), .ZN(new_n12391_));
  NAND4_X1   g11371(.A1(new_n12390_), .A2(new_n12391_), .A3(new_n12372_), .A4(new_n12383_), .ZN(new_n12392_));
  NOR2_X1    g11372(.A1(new_n12392_), .A2(new_n12389_), .ZN(new_n12393_));
  NOR2_X1    g11373(.A1(new_n12386_), .A2(new_n12393_), .ZN(new_n12394_));
  OAI22_X1   g11374(.A1(new_n12394_), .A2(new_n12385_), .B1(new_n12375_), .B2(new_n12382_), .ZN(new_n12395_));
  AOI22_X1   g11375(.A1(new_n12352_), .A2(new_n12356_), .B1(new_n12395_), .B2(new_n12266_), .ZN(new_n12396_));
  OAI21_X1   g11376(.A1(new_n12258_), .A2(new_n12254_), .B(new_n12195_), .ZN(new_n12397_));
  NOR2_X1    g11377(.A1(new_n12200_), .A2(new_n12205_), .ZN(new_n12398_));
  OAI21_X1   g11378(.A1(new_n12222_), .A2(new_n12398_), .B(new_n12252_), .ZN(new_n12399_));
  NOR2_X1    g11379(.A1(new_n12167_), .A2(new_n12171_), .ZN(new_n12400_));
  OAI21_X1   g11380(.A1(new_n12246_), .A2(new_n12400_), .B(new_n12247_), .ZN(new_n12401_));
  XNOR2_X1   g11381(.A1(new_n12399_), .A2(new_n12401_), .ZN(new_n12402_));
  NAND3_X1   g11382(.A1(new_n12397_), .A2(new_n12263_), .A3(new_n12402_), .ZN(new_n12403_));
  INV_X1     g11383(.I(new_n12382_), .ZN(new_n12404_));
  NAND2_X1   g11384(.A1(new_n12389_), .A2(new_n12384_), .ZN(new_n12405_));
  NAND2_X1   g11385(.A1(new_n12405_), .A2(new_n12404_), .ZN(new_n12406_));
  NOR2_X1    g11386(.A1(new_n12317_), .A2(new_n12318_), .ZN(new_n12407_));
  OAI21_X1   g11387(.A1(new_n12359_), .A2(new_n12407_), .B(new_n12319_), .ZN(new_n12408_));
  NOR2_X1    g11388(.A1(new_n12326_), .A2(new_n12331_), .ZN(new_n12409_));
  OAI21_X1   g11389(.A1(new_n12371_), .A2(new_n12409_), .B(new_n12370_), .ZN(new_n12410_));
  XNOR2_X1   g11390(.A1(new_n12410_), .A2(new_n12408_), .ZN(new_n12411_));
  NAND3_X1   g11391(.A1(new_n12406_), .A2(new_n12411_), .A3(new_n12375_), .ZN(new_n12412_));
  XOR2_X1    g11392(.A1(new_n12412_), .A2(new_n12403_), .Z(new_n12413_));
  NAND2_X1   g11393(.A1(new_n12413_), .A2(new_n12396_), .ZN(new_n12414_));
  NAND3_X1   g11394(.A1(new_n12261_), .A2(new_n12265_), .A3(new_n12355_), .ZN(new_n12415_));
  AOI21_X1   g11395(.A1(new_n12265_), .A2(new_n12261_), .B(new_n12355_), .ZN(new_n12416_));
  NOR3_X1    g11396(.A1(new_n12274_), .A2(new_n12351_), .A3(new_n12269_), .ZN(new_n12417_));
  NOR2_X1    g11397(.A1(new_n12375_), .A2(new_n12382_), .ZN(new_n12418_));
  INV_X1     g11398(.I(new_n12385_), .ZN(new_n12419_));
  XOR2_X1    g11399(.A1(new_n12392_), .A2(new_n12366_), .Z(new_n12420_));
  AOI21_X1   g11400(.A1(new_n12420_), .A2(new_n12419_), .B(new_n12418_), .ZN(new_n12421_));
  OAI21_X1   g11401(.A1(new_n12416_), .A2(new_n12417_), .B(new_n12421_), .ZN(new_n12422_));
  NAND2_X1   g11402(.A1(new_n12412_), .A2(new_n12403_), .ZN(new_n12423_));
  INV_X1     g11403(.I(new_n12403_), .ZN(new_n12424_));
  NAND4_X1   g11404(.A1(new_n12424_), .A2(new_n12375_), .A3(new_n12406_), .A4(new_n12411_), .ZN(new_n12425_));
  NAND2_X1   g11405(.A1(new_n12425_), .A2(new_n12423_), .ZN(new_n12426_));
  NAND3_X1   g11406(.A1(new_n12426_), .A2(new_n12415_), .A3(new_n12422_), .ZN(new_n12427_));
  NAND2_X1   g11407(.A1(new_n12427_), .A2(new_n12414_), .ZN(new_n12428_));
  NOR2_X1    g11408(.A1(new_n12428_), .A2(new_n12163_), .ZN(new_n12429_));
  NOR2_X1    g11409(.A1(new_n12417_), .A2(new_n12416_), .ZN(new_n12430_));
  NAND2_X1   g11410(.A1(new_n12353_), .A2(new_n12354_), .ZN(new_n12431_));
  NAND2_X1   g11411(.A1(new_n12084_), .A2(new_n12085_), .ZN(new_n12432_));
  NAND4_X1   g11412(.A1(new_n12082_), .A2(new_n12351_), .A3(new_n12431_), .A4(new_n12432_), .ZN(new_n12433_));
  INV_X1     g11413(.I(new_n12433_), .ZN(new_n12434_));
  AOI21_X1   g11414(.A1(new_n12430_), .A2(new_n12421_), .B(new_n12434_), .ZN(new_n12435_));
  NAND2_X1   g11415(.A1(new_n12352_), .A2(new_n12356_), .ZN(new_n12436_));
  NOR3_X1    g11416(.A1(new_n12436_), .A2(new_n12395_), .A3(new_n12433_), .ZN(new_n12437_));
  NOR2_X1    g11417(.A1(new_n12435_), .A2(new_n12437_), .ZN(new_n12438_));
  NOR2_X1    g11418(.A1(new_n12436_), .A2(new_n12395_), .ZN(new_n12439_));
  NAND2_X1   g11419(.A1(new_n12439_), .A2(new_n12434_), .ZN(new_n12440_));
  AOI21_X1   g11420(.A1(new_n12083_), .A2(new_n12087_), .B(new_n12129_), .ZN(new_n12441_));
  NOR3_X1    g11421(.A1(new_n12154_), .A2(new_n12149_), .A3(new_n12150_), .ZN(new_n12442_));
  NOR2_X1    g11422(.A1(new_n12441_), .A2(new_n12442_), .ZN(new_n12443_));
  INV_X1     g11423(.I(new_n12443_), .ZN(new_n12444_));
  OAI21_X1   g11424(.A1(new_n12444_), .A2(new_n12438_), .B(new_n12440_), .ZN(new_n12445_));
  NAND2_X1   g11425(.A1(new_n12428_), .A2(new_n12163_), .ZN(new_n12446_));
  AOI21_X1   g11426(.A1(new_n12445_), .A2(new_n12446_), .B(new_n12429_), .ZN(new_n12447_));
  NAND2_X1   g11427(.A1(new_n12133_), .A2(new_n12135_), .ZN(new_n12448_));
  NOR2_X1    g11428(.A1(new_n12131_), .A2(new_n12001_), .ZN(new_n12449_));
  OAI21_X1   g11429(.A1(new_n12133_), .A2(new_n12135_), .B(new_n12449_), .ZN(new_n12450_));
  NAND2_X1   g11430(.A1(new_n12450_), .A2(new_n12448_), .ZN(new_n12451_));
  NOR2_X1    g11431(.A1(new_n12158_), .A2(new_n12157_), .ZN(new_n12452_));
  NAND2_X1   g11432(.A1(new_n12141_), .A2(new_n12143_), .ZN(new_n12453_));
  NOR2_X1    g11433(.A1(new_n12139_), .A2(new_n12108_), .ZN(new_n12454_));
  OAI21_X1   g11434(.A1(new_n12141_), .A2(new_n12143_), .B(new_n12454_), .ZN(new_n12455_));
  NAND2_X1   g11435(.A1(new_n12455_), .A2(new_n12453_), .ZN(new_n12456_));
  INV_X1     g11436(.I(new_n12456_), .ZN(new_n12457_));
  NAND2_X1   g11437(.A1(new_n12155_), .A2(new_n12159_), .ZN(new_n12458_));
  AOI21_X1   g11438(.A1(new_n12458_), .A2(new_n12452_), .B(new_n12457_), .ZN(new_n12459_));
  NAND3_X1   g11439(.A1(new_n12130_), .A2(new_n12138_), .A3(new_n12145_), .ZN(new_n12460_));
  NOR2_X1    g11440(.A1(new_n12460_), .A2(new_n12456_), .ZN(new_n12461_));
  OAI21_X1   g11441(.A1(new_n12459_), .A2(new_n12461_), .B(new_n12451_), .ZN(new_n12462_));
  INV_X1     g11442(.I(new_n12451_), .ZN(new_n12463_));
  NAND2_X1   g11443(.A1(new_n12460_), .A2(new_n12456_), .ZN(new_n12464_));
  NAND4_X1   g11444(.A1(new_n12457_), .A2(new_n12130_), .A3(new_n12138_), .A4(new_n12145_), .ZN(new_n12465_));
  NAND3_X1   g11445(.A1(new_n12464_), .A2(new_n12463_), .A3(new_n12465_), .ZN(new_n12466_));
  NAND2_X1   g11446(.A1(new_n12397_), .A2(new_n12263_), .ZN(new_n12467_));
  NOR2_X1    g11447(.A1(new_n12399_), .A2(new_n12401_), .ZN(new_n12468_));
  NOR2_X1    g11448(.A1(new_n12467_), .A2(new_n12468_), .ZN(new_n12469_));
  AOI21_X1   g11449(.A1(new_n12399_), .A2(new_n12401_), .B(new_n12469_), .ZN(new_n12470_));
  INV_X1     g11450(.I(new_n12470_), .ZN(new_n12471_));
  INV_X1     g11451(.I(new_n12425_), .ZN(new_n12472_));
  NAND2_X1   g11452(.A1(new_n12406_), .A2(new_n12375_), .ZN(new_n12473_));
  NOR2_X1    g11453(.A1(new_n12410_), .A2(new_n12408_), .ZN(new_n12474_));
  NOR2_X1    g11454(.A1(new_n12473_), .A2(new_n12474_), .ZN(new_n12475_));
  AOI21_X1   g11455(.A1(new_n12408_), .A2(new_n12410_), .B(new_n12475_), .ZN(new_n12476_));
  NAND3_X1   g11456(.A1(new_n12422_), .A2(new_n12415_), .A3(new_n12423_), .ZN(new_n12477_));
  AOI21_X1   g11457(.A1(new_n12477_), .A2(new_n12472_), .B(new_n12476_), .ZN(new_n12478_));
  INV_X1     g11458(.I(new_n12412_), .ZN(new_n12479_));
  NAND4_X1   g11459(.A1(new_n12476_), .A2(new_n12396_), .A3(new_n12424_), .A4(new_n12479_), .ZN(new_n12480_));
  INV_X1     g11460(.I(new_n12480_), .ZN(new_n12481_));
  OAI21_X1   g11461(.A1(new_n12481_), .A2(new_n12478_), .B(new_n12471_), .ZN(new_n12482_));
  INV_X1     g11462(.I(new_n12476_), .ZN(new_n12483_));
  NAND3_X1   g11463(.A1(new_n12396_), .A2(new_n12424_), .A3(new_n12479_), .ZN(new_n12484_));
  NAND2_X1   g11464(.A1(new_n12484_), .A2(new_n12483_), .ZN(new_n12485_));
  NAND3_X1   g11465(.A1(new_n12485_), .A2(new_n12470_), .A3(new_n12480_), .ZN(new_n12486_));
  NAND4_X1   g11466(.A1(new_n12462_), .A2(new_n12482_), .A3(new_n12466_), .A4(new_n12486_), .ZN(new_n12487_));
  NAND2_X1   g11467(.A1(new_n12487_), .A2(new_n12447_), .ZN(new_n12488_));
  XOR2_X1    g11468(.A1(new_n12451_), .A2(new_n12456_), .Z(new_n12489_));
  XNOR2_X1   g11469(.A1(new_n12476_), .A2(new_n12470_), .ZN(new_n12490_));
  INV_X1     g11470(.I(new_n12490_), .ZN(new_n12491_));
  NOR4_X1    g11471(.A1(new_n12491_), .A2(new_n12460_), .A3(new_n12484_), .A4(new_n12489_), .ZN(new_n12492_));
  NAND2_X1   g11472(.A1(new_n12488_), .A2(new_n12492_), .ZN(new_n12493_));
  OAI21_X1   g11473(.A1(new_n12451_), .A2(new_n12456_), .B(new_n12460_), .ZN(new_n12494_));
  NAND2_X1   g11474(.A1(new_n12476_), .A2(new_n12470_), .ZN(new_n12495_));
  NAND2_X1   g11475(.A1(new_n12484_), .A2(new_n12495_), .ZN(new_n12496_));
  NAND2_X1   g11476(.A1(new_n12483_), .A2(new_n12471_), .ZN(new_n12497_));
  NAND2_X1   g11477(.A1(new_n12451_), .A2(new_n12456_), .ZN(new_n12498_));
  NAND4_X1   g11478(.A1(new_n12494_), .A2(new_n12496_), .A3(new_n12497_), .A4(new_n12498_), .ZN(new_n12499_));
  INV_X1     g11479(.I(new_n12499_), .ZN(new_n12500_));
  NAND2_X1   g11480(.A1(new_n12496_), .A2(new_n12497_), .ZN(new_n12501_));
  NAND2_X1   g11481(.A1(new_n12494_), .A2(new_n12498_), .ZN(new_n12502_));
  AOI22_X1   g11482(.A1(new_n12493_), .A2(new_n12500_), .B1(new_n12501_), .B2(new_n12502_), .ZN(new_n12503_));
  INV_X1     g11483(.I(new_n12503_), .ZN(new_n12504_));
  INV_X1     g11484(.I(\A[796] ), .ZN(new_n12505_));
  NOR2_X1    g11485(.A1(\A[797] ), .A2(\A[798] ), .ZN(new_n12506_));
  NAND2_X1   g11486(.A1(\A[797] ), .A2(\A[798] ), .ZN(new_n12507_));
  AOI21_X1   g11487(.A1(new_n12505_), .A2(new_n12507_), .B(new_n12506_), .ZN(new_n12508_));
  INV_X1     g11488(.I(new_n12508_), .ZN(new_n12509_));
  INV_X1     g11489(.I(\A[793] ), .ZN(new_n12510_));
  NOR2_X1    g11490(.A1(\A[794] ), .A2(\A[795] ), .ZN(new_n12511_));
  NAND2_X1   g11491(.A1(\A[794] ), .A2(\A[795] ), .ZN(new_n12512_));
  AOI21_X1   g11492(.A1(new_n12510_), .A2(new_n12512_), .B(new_n12511_), .ZN(new_n12513_));
  INV_X1     g11493(.I(new_n12513_), .ZN(new_n12514_));
  NOR2_X1    g11494(.A1(new_n12509_), .A2(new_n12514_), .ZN(new_n12515_));
  NOR2_X1    g11495(.A1(new_n12508_), .A2(new_n12513_), .ZN(new_n12516_));
  INV_X1     g11496(.I(new_n12516_), .ZN(new_n12517_));
  INV_X1     g11497(.I(\A[795] ), .ZN(new_n12518_));
  NOR2_X1    g11498(.A1(new_n12518_), .A2(\A[794] ), .ZN(new_n12519_));
  INV_X1     g11499(.I(\A[794] ), .ZN(new_n12520_));
  NOR2_X1    g11500(.A1(new_n12520_), .A2(\A[795] ), .ZN(new_n12521_));
  OAI21_X1   g11501(.A1(new_n12519_), .A2(new_n12521_), .B(\A[793] ), .ZN(new_n12522_));
  INV_X1     g11502(.I(new_n12512_), .ZN(new_n12523_));
  OAI21_X1   g11503(.A1(new_n12523_), .A2(new_n12511_), .B(new_n12510_), .ZN(new_n12524_));
  NAND2_X1   g11504(.A1(new_n12522_), .A2(new_n12524_), .ZN(new_n12525_));
  INV_X1     g11505(.I(\A[797] ), .ZN(new_n12526_));
  NAND2_X1   g11506(.A1(new_n12526_), .A2(\A[798] ), .ZN(new_n12527_));
  INV_X1     g11507(.I(\A[798] ), .ZN(new_n12528_));
  NAND2_X1   g11508(.A1(new_n12528_), .A2(\A[797] ), .ZN(new_n12529_));
  AOI21_X1   g11509(.A1(new_n12527_), .A2(new_n12529_), .B(new_n12505_), .ZN(new_n12530_));
  INV_X1     g11510(.I(new_n12506_), .ZN(new_n12531_));
  AOI21_X1   g11511(.A1(new_n12531_), .A2(new_n12507_), .B(\A[796] ), .ZN(new_n12532_));
  NOR3_X1    g11512(.A1(new_n12525_), .A2(new_n12530_), .A3(new_n12532_), .ZN(new_n12533_));
  AOI21_X1   g11513(.A1(new_n12533_), .A2(new_n12517_), .B(new_n12515_), .ZN(new_n12534_));
  INV_X1     g11514(.I(new_n12534_), .ZN(new_n12535_));
  INV_X1     g11515(.I(\A[790] ), .ZN(new_n12536_));
  NOR2_X1    g11516(.A1(\A[791] ), .A2(\A[792] ), .ZN(new_n12537_));
  NAND2_X1   g11517(.A1(\A[791] ), .A2(\A[792] ), .ZN(new_n12538_));
  AOI21_X1   g11518(.A1(new_n12536_), .A2(new_n12538_), .B(new_n12537_), .ZN(new_n12539_));
  NOR2_X1    g11519(.A1(\A[788] ), .A2(\A[789] ), .ZN(new_n12540_));
  INV_X1     g11520(.I(\A[788] ), .ZN(new_n12541_));
  INV_X1     g11521(.I(\A[789] ), .ZN(new_n12542_));
  NOR2_X1    g11522(.A1(new_n12541_), .A2(new_n12542_), .ZN(new_n12543_));
  NOR2_X1    g11523(.A1(new_n12543_), .A2(\A[787] ), .ZN(new_n12544_));
  NOR2_X1    g11524(.A1(new_n12544_), .A2(new_n12540_), .ZN(new_n12545_));
  NAND2_X1   g11525(.A1(new_n12545_), .A2(new_n12539_), .ZN(new_n12546_));
  NOR2_X1    g11526(.A1(new_n12542_), .A2(\A[788] ), .ZN(new_n12547_));
  NOR2_X1    g11527(.A1(new_n12541_), .A2(\A[789] ), .ZN(new_n12548_));
  OAI21_X1   g11528(.A1(new_n12547_), .A2(new_n12548_), .B(\A[787] ), .ZN(new_n12549_));
  INV_X1     g11529(.I(\A[787] ), .ZN(new_n12550_));
  OAI21_X1   g11530(.A1(new_n12543_), .A2(new_n12540_), .B(new_n12550_), .ZN(new_n12551_));
  NAND2_X1   g11531(.A1(new_n12551_), .A2(new_n12549_), .ZN(new_n12552_));
  INV_X1     g11532(.I(\A[792] ), .ZN(new_n12553_));
  NOR2_X1    g11533(.A1(new_n12553_), .A2(\A[791] ), .ZN(new_n12554_));
  INV_X1     g11534(.I(\A[791] ), .ZN(new_n12555_));
  NOR2_X1    g11535(.A1(new_n12555_), .A2(\A[792] ), .ZN(new_n12556_));
  OAI21_X1   g11536(.A1(new_n12554_), .A2(new_n12556_), .B(\A[790] ), .ZN(new_n12557_));
  INV_X1     g11537(.I(new_n12538_), .ZN(new_n12558_));
  OAI21_X1   g11538(.A1(new_n12558_), .A2(new_n12537_), .B(new_n12536_), .ZN(new_n12559_));
  NAND2_X1   g11539(.A1(new_n12557_), .A2(new_n12559_), .ZN(new_n12560_));
  NOR2_X1    g11540(.A1(new_n12552_), .A2(new_n12560_), .ZN(new_n12561_));
  OAI21_X1   g11541(.A1(new_n12539_), .A2(new_n12545_), .B(new_n12561_), .ZN(new_n12562_));
  NAND2_X1   g11542(.A1(new_n12562_), .A2(new_n12546_), .ZN(new_n12563_));
  NAND2_X1   g11543(.A1(new_n12563_), .A2(new_n12535_), .ZN(new_n12564_));
  NOR2_X1    g11544(.A1(new_n12563_), .A2(new_n12535_), .ZN(new_n12565_));
  INV_X1     g11545(.I(new_n12539_), .ZN(new_n12566_));
  XNOR2_X1   g11546(.A1(new_n12561_), .A2(new_n12545_), .ZN(new_n12567_));
  NOR2_X1    g11547(.A1(new_n12567_), .A2(new_n12566_), .ZN(new_n12568_));
  XOR2_X1    g11548(.A1(new_n12561_), .A2(new_n12545_), .Z(new_n12569_));
  NOR2_X1    g11549(.A1(new_n12569_), .A2(new_n12539_), .ZN(new_n12570_));
  NOR2_X1    g11550(.A1(new_n12533_), .A2(new_n12514_), .ZN(new_n12571_));
  AND2_X2    g11551(.A1(new_n12522_), .A2(new_n12524_), .Z(new_n12572_));
  NOR2_X1    g11552(.A1(new_n12532_), .A2(new_n12530_), .ZN(new_n12573_));
  NAND2_X1   g11553(.A1(new_n12572_), .A2(new_n12573_), .ZN(new_n12574_));
  NOR2_X1    g11554(.A1(new_n12574_), .A2(new_n12513_), .ZN(new_n12575_));
  OAI21_X1   g11555(.A1(new_n12575_), .A2(new_n12571_), .B(new_n12508_), .ZN(new_n12576_));
  NAND2_X1   g11556(.A1(new_n12574_), .A2(new_n12513_), .ZN(new_n12577_));
  NAND2_X1   g11557(.A1(new_n12533_), .A2(new_n12514_), .ZN(new_n12578_));
  NAND3_X1   g11558(.A1(new_n12577_), .A2(new_n12509_), .A3(new_n12578_), .ZN(new_n12579_));
  NAND2_X1   g11559(.A1(new_n12576_), .A2(new_n12579_), .ZN(new_n12580_));
  AOI22_X1   g11560(.A1(new_n12549_), .A2(new_n12551_), .B1(new_n12557_), .B2(new_n12559_), .ZN(new_n12581_));
  NOR2_X1    g11561(.A1(new_n12572_), .A2(new_n12573_), .ZN(new_n12582_));
  NOR4_X1    g11562(.A1(new_n12582_), .A2(new_n12533_), .A3(new_n12561_), .A4(new_n12581_), .ZN(new_n12583_));
  INV_X1     g11563(.I(new_n12583_), .ZN(new_n12584_));
  NAND2_X1   g11564(.A1(new_n12533_), .A2(new_n12515_), .ZN(new_n12585_));
  NOR3_X1    g11565(.A1(new_n12546_), .A2(new_n12552_), .A3(new_n12560_), .ZN(new_n12586_));
  NAND2_X1   g11566(.A1(new_n12585_), .A2(new_n12586_), .ZN(new_n12587_));
  NOR2_X1    g11567(.A1(new_n12584_), .A2(new_n12587_), .ZN(new_n12588_));
  OAI22_X1   g11568(.A1(new_n12580_), .A2(new_n12588_), .B1(new_n12568_), .B2(new_n12570_), .ZN(new_n12589_));
  INV_X1     g11569(.I(new_n12515_), .ZN(new_n12590_));
  OAI21_X1   g11570(.A1(new_n12582_), .A2(new_n12590_), .B(new_n12586_), .ZN(new_n12591_));
  XNOR2_X1   g11571(.A1(new_n12508_), .A2(new_n12513_), .ZN(new_n12592_));
  NOR2_X1    g11572(.A1(new_n12574_), .A2(new_n12592_), .ZN(new_n12593_));
  AOI21_X1   g11573(.A1(new_n12590_), .A2(new_n12517_), .B(new_n12533_), .ZN(new_n12594_));
  NOR3_X1    g11574(.A1(new_n12591_), .A2(new_n12594_), .A3(new_n12593_), .ZN(new_n12595_));
  NAND2_X1   g11575(.A1(new_n12595_), .A2(new_n12583_), .ZN(new_n12596_));
  NAND2_X1   g11576(.A1(new_n12589_), .A2(new_n12596_), .ZN(new_n12597_));
  OAI21_X1   g11577(.A1(new_n12597_), .A2(new_n12565_), .B(new_n12564_), .ZN(new_n12598_));
  INV_X1     g11578(.I(\A[784] ), .ZN(new_n12599_));
  NOR2_X1    g11579(.A1(\A[785] ), .A2(\A[786] ), .ZN(new_n12600_));
  NAND2_X1   g11580(.A1(\A[785] ), .A2(\A[786] ), .ZN(new_n12601_));
  AOI21_X1   g11581(.A1(new_n12599_), .A2(new_n12601_), .B(new_n12600_), .ZN(new_n12602_));
  INV_X1     g11582(.I(new_n12602_), .ZN(new_n12603_));
  INV_X1     g11583(.I(\A[781] ), .ZN(new_n12604_));
  NOR2_X1    g11584(.A1(\A[782] ), .A2(\A[783] ), .ZN(new_n12605_));
  NAND2_X1   g11585(.A1(\A[782] ), .A2(\A[783] ), .ZN(new_n12606_));
  AOI21_X1   g11586(.A1(new_n12604_), .A2(new_n12606_), .B(new_n12605_), .ZN(new_n12607_));
  INV_X1     g11587(.I(new_n12607_), .ZN(new_n12608_));
  NOR2_X1    g11588(.A1(new_n12603_), .A2(new_n12608_), .ZN(new_n12609_));
  NAND2_X1   g11589(.A1(new_n12603_), .A2(new_n12608_), .ZN(new_n12610_));
  INV_X1     g11590(.I(\A[782] ), .ZN(new_n12611_));
  NAND2_X1   g11591(.A1(new_n12611_), .A2(\A[783] ), .ZN(new_n12612_));
  INV_X1     g11592(.I(\A[783] ), .ZN(new_n12613_));
  NAND2_X1   g11593(.A1(new_n12613_), .A2(\A[782] ), .ZN(new_n12614_));
  AOI21_X1   g11594(.A1(new_n12612_), .A2(new_n12614_), .B(new_n12604_), .ZN(new_n12615_));
  INV_X1     g11595(.I(new_n12605_), .ZN(new_n12616_));
  AOI21_X1   g11596(.A1(new_n12616_), .A2(new_n12606_), .B(\A[781] ), .ZN(new_n12617_));
  INV_X1     g11597(.I(\A[785] ), .ZN(new_n12618_));
  NAND2_X1   g11598(.A1(new_n12618_), .A2(\A[786] ), .ZN(new_n12619_));
  INV_X1     g11599(.I(\A[786] ), .ZN(new_n12620_));
  NAND2_X1   g11600(.A1(new_n12620_), .A2(\A[785] ), .ZN(new_n12621_));
  AOI21_X1   g11601(.A1(new_n12619_), .A2(new_n12621_), .B(new_n12599_), .ZN(new_n12622_));
  INV_X1     g11602(.I(new_n12600_), .ZN(new_n12623_));
  AOI21_X1   g11603(.A1(new_n12623_), .A2(new_n12601_), .B(\A[784] ), .ZN(new_n12624_));
  NOR4_X1    g11604(.A1(new_n12615_), .A2(new_n12617_), .A3(new_n12624_), .A4(new_n12622_), .ZN(new_n12625_));
  AOI21_X1   g11605(.A1(new_n12625_), .A2(new_n12610_), .B(new_n12609_), .ZN(new_n12626_));
  INV_X1     g11606(.I(\A[778] ), .ZN(new_n12627_));
  NOR2_X1    g11607(.A1(\A[779] ), .A2(\A[780] ), .ZN(new_n12628_));
  NAND2_X1   g11608(.A1(\A[779] ), .A2(\A[780] ), .ZN(new_n12629_));
  AOI21_X1   g11609(.A1(new_n12627_), .A2(new_n12629_), .B(new_n12628_), .ZN(new_n12630_));
  INV_X1     g11610(.I(\A[775] ), .ZN(new_n12631_));
  NOR2_X1    g11611(.A1(\A[776] ), .A2(\A[777] ), .ZN(new_n12632_));
  NAND2_X1   g11612(.A1(\A[776] ), .A2(\A[777] ), .ZN(new_n12633_));
  AOI21_X1   g11613(.A1(new_n12631_), .A2(new_n12633_), .B(new_n12632_), .ZN(new_n12634_));
  NAND2_X1   g11614(.A1(new_n12630_), .A2(new_n12634_), .ZN(new_n12635_));
  INV_X1     g11615(.I(\A[776] ), .ZN(new_n12636_));
  NAND2_X1   g11616(.A1(new_n12636_), .A2(\A[777] ), .ZN(new_n12637_));
  INV_X1     g11617(.I(\A[777] ), .ZN(new_n12638_));
  NAND2_X1   g11618(.A1(new_n12638_), .A2(\A[776] ), .ZN(new_n12639_));
  AOI21_X1   g11619(.A1(new_n12637_), .A2(new_n12639_), .B(new_n12631_), .ZN(new_n12640_));
  INV_X1     g11620(.I(new_n12632_), .ZN(new_n12641_));
  AOI21_X1   g11621(.A1(new_n12641_), .A2(new_n12633_), .B(\A[775] ), .ZN(new_n12642_));
  INV_X1     g11622(.I(\A[779] ), .ZN(new_n12643_));
  NAND2_X1   g11623(.A1(new_n12643_), .A2(\A[780] ), .ZN(new_n12644_));
  INV_X1     g11624(.I(\A[780] ), .ZN(new_n12645_));
  NAND2_X1   g11625(.A1(new_n12645_), .A2(\A[779] ), .ZN(new_n12646_));
  AOI21_X1   g11626(.A1(new_n12644_), .A2(new_n12646_), .B(new_n12627_), .ZN(new_n12647_));
  INV_X1     g11627(.I(new_n12628_), .ZN(new_n12648_));
  AOI21_X1   g11628(.A1(new_n12648_), .A2(new_n12629_), .B(\A[778] ), .ZN(new_n12649_));
  NOR4_X1    g11629(.A1(new_n12640_), .A2(new_n12642_), .A3(new_n12649_), .A4(new_n12647_), .ZN(new_n12650_));
  OAI21_X1   g11630(.A1(new_n12630_), .A2(new_n12634_), .B(new_n12650_), .ZN(new_n12651_));
  NAND2_X1   g11631(.A1(new_n12651_), .A2(new_n12635_), .ZN(new_n12652_));
  INV_X1     g11632(.I(new_n12652_), .ZN(new_n12653_));
  NOR2_X1    g11633(.A1(new_n12653_), .A2(new_n12626_), .ZN(new_n12654_));
  INV_X1     g11634(.I(new_n12630_), .ZN(new_n12655_));
  INV_X1     g11635(.I(new_n12634_), .ZN(new_n12656_));
  NOR2_X1    g11636(.A1(new_n12650_), .A2(new_n12656_), .ZN(new_n12657_));
  INV_X1     g11637(.I(new_n12657_), .ZN(new_n12658_));
  NAND2_X1   g11638(.A1(new_n12650_), .A2(new_n12656_), .ZN(new_n12659_));
  AOI21_X1   g11639(.A1(new_n12658_), .A2(new_n12659_), .B(new_n12655_), .ZN(new_n12660_));
  INV_X1     g11640(.I(new_n12659_), .ZN(new_n12661_));
  NOR3_X1    g11641(.A1(new_n12661_), .A2(new_n12630_), .A3(new_n12657_), .ZN(new_n12662_));
  NOR2_X1    g11642(.A1(new_n12625_), .A2(new_n12608_), .ZN(new_n12663_));
  NAND2_X1   g11643(.A1(new_n12625_), .A2(new_n12608_), .ZN(new_n12664_));
  INV_X1     g11644(.I(new_n12664_), .ZN(new_n12665_));
  OAI21_X1   g11645(.A1(new_n12665_), .A2(new_n12663_), .B(new_n12602_), .ZN(new_n12666_));
  NOR2_X1    g11646(.A1(new_n12617_), .A2(new_n12615_), .ZN(new_n12667_));
  NOR2_X1    g11647(.A1(new_n12624_), .A2(new_n12622_), .ZN(new_n12668_));
  NAND2_X1   g11648(.A1(new_n12667_), .A2(new_n12668_), .ZN(new_n12669_));
  NAND2_X1   g11649(.A1(new_n12669_), .A2(new_n12607_), .ZN(new_n12670_));
  NAND3_X1   g11650(.A1(new_n12670_), .A2(new_n12603_), .A3(new_n12664_), .ZN(new_n12671_));
  NAND2_X1   g11651(.A1(new_n12666_), .A2(new_n12671_), .ZN(new_n12672_));
  NOR2_X1    g11652(.A1(new_n12642_), .A2(new_n12640_), .ZN(new_n12673_));
  NOR2_X1    g11653(.A1(new_n12649_), .A2(new_n12647_), .ZN(new_n12674_));
  NOR2_X1    g11654(.A1(new_n12673_), .A2(new_n12674_), .ZN(new_n12675_));
  NOR2_X1    g11655(.A1(new_n12675_), .A2(new_n12650_), .ZN(new_n12676_));
  NOR2_X1    g11656(.A1(new_n12667_), .A2(new_n12668_), .ZN(new_n12677_));
  NOR2_X1    g11657(.A1(new_n12677_), .A2(new_n12625_), .ZN(new_n12678_));
  NAND2_X1   g11658(.A1(new_n12676_), .A2(new_n12678_), .ZN(new_n12679_));
  NAND2_X1   g11659(.A1(new_n12625_), .A2(new_n12609_), .ZN(new_n12680_));
  NAND2_X1   g11660(.A1(new_n12673_), .A2(new_n12674_), .ZN(new_n12681_));
  NOR2_X1    g11661(.A1(new_n12681_), .A2(new_n12635_), .ZN(new_n12682_));
  NAND2_X1   g11662(.A1(new_n12682_), .A2(new_n12680_), .ZN(new_n12683_));
  NOR2_X1    g11663(.A1(new_n12679_), .A2(new_n12683_), .ZN(new_n12684_));
  OAI22_X1   g11664(.A1(new_n12672_), .A2(new_n12684_), .B1(new_n12660_), .B2(new_n12662_), .ZN(new_n12685_));
  INV_X1     g11665(.I(new_n12609_), .ZN(new_n12686_));
  OAI21_X1   g11666(.A1(new_n12686_), .A2(new_n12677_), .B(new_n12682_), .ZN(new_n12687_));
  XNOR2_X1   g11667(.A1(new_n12602_), .A2(new_n12607_), .ZN(new_n12688_));
  NOR2_X1    g11668(.A1(new_n12669_), .A2(new_n12688_), .ZN(new_n12689_));
  AOI21_X1   g11669(.A1(new_n12686_), .A2(new_n12610_), .B(new_n12625_), .ZN(new_n12690_));
  NOR4_X1    g11670(.A1(new_n12687_), .A2(new_n12679_), .A3(new_n12689_), .A4(new_n12690_), .ZN(new_n12691_));
  INV_X1     g11671(.I(new_n12691_), .ZN(new_n12692_));
  NAND2_X1   g11672(.A1(new_n12685_), .A2(new_n12692_), .ZN(new_n12693_));
  AOI21_X1   g11673(.A1(new_n12626_), .A2(new_n12653_), .B(new_n12693_), .ZN(new_n12694_));
  NOR2_X1    g11674(.A1(new_n12694_), .A2(new_n12654_), .ZN(new_n12695_));
  INV_X1     g11675(.I(new_n12695_), .ZN(new_n12696_));
  NOR2_X1    g11676(.A1(new_n12568_), .A2(new_n12570_), .ZN(new_n12697_));
  AOI21_X1   g11677(.A1(new_n12577_), .A2(new_n12578_), .B(new_n12509_), .ZN(new_n12698_));
  NOR3_X1    g11678(.A1(new_n12575_), .A2(new_n12508_), .A3(new_n12571_), .ZN(new_n12699_));
  NOR2_X1    g11679(.A1(new_n12699_), .A2(new_n12698_), .ZN(new_n12700_));
  NAND3_X1   g11680(.A1(new_n12583_), .A2(new_n12585_), .A3(new_n12586_), .ZN(new_n12701_));
  NAND2_X1   g11681(.A1(new_n12700_), .A2(new_n12701_), .ZN(new_n12702_));
  NAND3_X1   g11682(.A1(new_n12702_), .A2(new_n12697_), .A3(new_n12596_), .ZN(new_n12703_));
  NOR2_X1    g11683(.A1(new_n12700_), .A2(new_n12588_), .ZN(new_n12704_));
  NOR2_X1    g11684(.A1(new_n12580_), .A2(new_n12701_), .ZN(new_n12705_));
  OAI21_X1   g11685(.A1(new_n12704_), .A2(new_n12705_), .B(new_n12697_), .ZN(new_n12706_));
  NAND2_X1   g11686(.A1(new_n12706_), .A2(new_n12703_), .ZN(new_n12707_));
  NOR2_X1    g11687(.A1(new_n12582_), .A2(new_n12533_), .ZN(new_n12708_));
  NAND2_X1   g11688(.A1(new_n12708_), .A2(new_n12585_), .ZN(new_n12709_));
  NOR2_X1    g11689(.A1(new_n12561_), .A2(new_n12581_), .ZN(new_n12710_));
  NAND2_X1   g11690(.A1(new_n12710_), .A2(new_n12586_), .ZN(new_n12711_));
  XNOR2_X1   g11691(.A1(new_n12709_), .A2(new_n12711_), .ZN(new_n12712_));
  NAND2_X1   g11692(.A1(new_n12678_), .A2(new_n12680_), .ZN(new_n12713_));
  NAND2_X1   g11693(.A1(new_n12676_), .A2(new_n12682_), .ZN(new_n12714_));
  XNOR2_X1   g11694(.A1(new_n12714_), .A2(new_n12713_), .ZN(new_n12715_));
  NOR2_X1    g11695(.A1(new_n12712_), .A2(new_n12715_), .ZN(new_n12716_));
  AOI21_X1   g11696(.A1(new_n12706_), .A2(new_n12703_), .B(new_n12716_), .ZN(new_n12717_));
  INV_X1     g11697(.I(new_n12717_), .ZN(new_n12718_));
  NAND3_X1   g11698(.A1(new_n12706_), .A2(new_n12716_), .A3(new_n12703_), .ZN(new_n12719_));
  NOR2_X1    g11699(.A1(new_n12660_), .A2(new_n12662_), .ZN(new_n12720_));
  INV_X1     g11700(.I(new_n12720_), .ZN(new_n12721_));
  NAND2_X1   g11701(.A1(new_n12721_), .A2(new_n12684_), .ZN(new_n12722_));
  INV_X1     g11702(.I(new_n12684_), .ZN(new_n12723_));
  AOI21_X1   g11703(.A1(new_n12723_), .A2(new_n12720_), .B(new_n12672_), .ZN(new_n12724_));
  INV_X1     g11704(.I(new_n12672_), .ZN(new_n12725_));
  NOR3_X1    g11705(.A1(new_n12721_), .A2(new_n12725_), .A3(new_n12684_), .ZN(new_n12726_));
  OAI21_X1   g11706(.A1(new_n12726_), .A2(new_n12724_), .B(new_n12722_), .ZN(new_n12727_));
  OAI21_X1   g11707(.A1(new_n12720_), .A2(new_n12692_), .B(new_n12727_), .ZN(new_n12728_));
  AOI22_X1   g11708(.A1(new_n12718_), .A2(new_n12719_), .B1(new_n12728_), .B2(new_n12707_), .ZN(new_n12729_));
  INV_X1     g11709(.I(new_n12563_), .ZN(new_n12730_));
  AOI21_X1   g11710(.A1(new_n12589_), .A2(new_n12596_), .B(new_n12730_), .ZN(new_n12731_));
  NAND2_X1   g11711(.A1(new_n12569_), .A2(new_n12539_), .ZN(new_n12732_));
  NAND2_X1   g11712(.A1(new_n12567_), .A2(new_n12566_), .ZN(new_n12733_));
  AOI22_X1   g11713(.A1(new_n12700_), .A2(new_n12701_), .B1(new_n12733_), .B2(new_n12732_), .ZN(new_n12734_));
  INV_X1     g11714(.I(new_n12596_), .ZN(new_n12735_));
  NOR3_X1    g11715(.A1(new_n12734_), .A2(new_n12735_), .A3(new_n12563_), .ZN(new_n12736_));
  OAI21_X1   g11716(.A1(new_n12731_), .A2(new_n12736_), .B(new_n12535_), .ZN(new_n12737_));
  OAI21_X1   g11717(.A1(new_n12734_), .A2(new_n12735_), .B(new_n12563_), .ZN(new_n12738_));
  NAND3_X1   g11718(.A1(new_n12589_), .A2(new_n12730_), .A3(new_n12596_), .ZN(new_n12739_));
  NAND3_X1   g11719(.A1(new_n12738_), .A2(new_n12739_), .A3(new_n12534_), .ZN(new_n12740_));
  NAND2_X1   g11720(.A1(new_n12737_), .A2(new_n12740_), .ZN(new_n12741_));
  INV_X1     g11721(.I(new_n12626_), .ZN(new_n12742_));
  AOI21_X1   g11722(.A1(new_n12685_), .A2(new_n12692_), .B(new_n12653_), .ZN(new_n12743_));
  NAND3_X1   g11723(.A1(new_n12685_), .A2(new_n12692_), .A3(new_n12653_), .ZN(new_n12744_));
  INV_X1     g11724(.I(new_n12744_), .ZN(new_n12745_));
  OAI21_X1   g11725(.A1(new_n12745_), .A2(new_n12743_), .B(new_n12742_), .ZN(new_n12746_));
  INV_X1     g11726(.I(new_n12743_), .ZN(new_n12747_));
  NAND3_X1   g11727(.A1(new_n12747_), .A2(new_n12626_), .A3(new_n12744_), .ZN(new_n12748_));
  NAND2_X1   g11728(.A1(new_n12748_), .A2(new_n12746_), .ZN(new_n12749_));
  NOR2_X1    g11729(.A1(new_n12749_), .A2(new_n12741_), .ZN(new_n12750_));
  XOR2_X1    g11730(.A1(new_n12563_), .A2(new_n12534_), .Z(new_n12751_));
  INV_X1     g11731(.I(new_n12751_), .ZN(new_n12752_));
  XOR2_X1    g11732(.A1(new_n12652_), .A2(new_n12742_), .Z(new_n12753_));
  NOR4_X1    g11733(.A1(new_n12597_), .A2(new_n12693_), .A3(new_n12752_), .A4(new_n12753_), .ZN(new_n12754_));
  OAI21_X1   g11734(.A1(new_n12750_), .A2(new_n12729_), .B(new_n12754_), .ZN(new_n12755_));
  OAI21_X1   g11735(.A1(new_n12598_), .A2(new_n12696_), .B(new_n12755_), .ZN(new_n12756_));
  NAND2_X1   g11736(.A1(new_n12696_), .A2(new_n12598_), .ZN(new_n12757_));
  NAND2_X1   g11737(.A1(new_n12756_), .A2(new_n12757_), .ZN(new_n12758_));
  INV_X1     g11738(.I(new_n12758_), .ZN(new_n12759_));
  INV_X1     g11739(.I(\A[772] ), .ZN(new_n12760_));
  NOR2_X1    g11740(.A1(\A[773] ), .A2(\A[774] ), .ZN(new_n12761_));
  NAND2_X1   g11741(.A1(\A[773] ), .A2(\A[774] ), .ZN(new_n12762_));
  AOI21_X1   g11742(.A1(new_n12760_), .A2(new_n12762_), .B(new_n12761_), .ZN(new_n12763_));
  INV_X1     g11743(.I(new_n12763_), .ZN(new_n12764_));
  INV_X1     g11744(.I(\A[769] ), .ZN(new_n12765_));
  NOR2_X1    g11745(.A1(\A[770] ), .A2(\A[771] ), .ZN(new_n12766_));
  NAND2_X1   g11746(.A1(\A[770] ), .A2(\A[771] ), .ZN(new_n12767_));
  AOI21_X1   g11747(.A1(new_n12765_), .A2(new_n12767_), .B(new_n12766_), .ZN(new_n12768_));
  INV_X1     g11748(.I(new_n12768_), .ZN(new_n12769_));
  NOR2_X1    g11749(.A1(new_n12764_), .A2(new_n12769_), .ZN(new_n12770_));
  INV_X1     g11750(.I(new_n12770_), .ZN(new_n12771_));
  NOR2_X1    g11751(.A1(new_n12763_), .A2(new_n12768_), .ZN(new_n12772_));
  INV_X1     g11752(.I(\A[770] ), .ZN(new_n12773_));
  NAND2_X1   g11753(.A1(new_n12773_), .A2(\A[771] ), .ZN(new_n12774_));
  INV_X1     g11754(.I(\A[771] ), .ZN(new_n12775_));
  NAND2_X1   g11755(.A1(new_n12775_), .A2(\A[770] ), .ZN(new_n12776_));
  AOI21_X1   g11756(.A1(new_n12774_), .A2(new_n12776_), .B(new_n12765_), .ZN(new_n12777_));
  INV_X1     g11757(.I(new_n12766_), .ZN(new_n12778_));
  AOI21_X1   g11758(.A1(new_n12778_), .A2(new_n12767_), .B(\A[769] ), .ZN(new_n12779_));
  NOR2_X1    g11759(.A1(new_n12779_), .A2(new_n12777_), .ZN(new_n12780_));
  INV_X1     g11760(.I(\A[773] ), .ZN(new_n12781_));
  NAND2_X1   g11761(.A1(new_n12781_), .A2(\A[774] ), .ZN(new_n12782_));
  INV_X1     g11762(.I(\A[774] ), .ZN(new_n12783_));
  NAND2_X1   g11763(.A1(new_n12783_), .A2(\A[773] ), .ZN(new_n12784_));
  AOI21_X1   g11764(.A1(new_n12782_), .A2(new_n12784_), .B(new_n12760_), .ZN(new_n12785_));
  INV_X1     g11765(.I(new_n12761_), .ZN(new_n12786_));
  AOI21_X1   g11766(.A1(new_n12786_), .A2(new_n12762_), .B(\A[772] ), .ZN(new_n12787_));
  NOR2_X1    g11767(.A1(new_n12787_), .A2(new_n12785_), .ZN(new_n12788_));
  NAND2_X1   g11768(.A1(new_n12780_), .A2(new_n12788_), .ZN(new_n12789_));
  OAI21_X1   g11769(.A1(new_n12789_), .A2(new_n12772_), .B(new_n12771_), .ZN(new_n12790_));
  INV_X1     g11770(.I(\A[766] ), .ZN(new_n12791_));
  NOR2_X1    g11771(.A1(\A[767] ), .A2(\A[768] ), .ZN(new_n12792_));
  NAND2_X1   g11772(.A1(\A[767] ), .A2(\A[768] ), .ZN(new_n12793_));
  AOI21_X1   g11773(.A1(new_n12791_), .A2(new_n12793_), .B(new_n12792_), .ZN(new_n12794_));
  INV_X1     g11774(.I(\A[763] ), .ZN(new_n12795_));
  NOR2_X1    g11775(.A1(\A[764] ), .A2(\A[765] ), .ZN(new_n12796_));
  NAND2_X1   g11776(.A1(\A[764] ), .A2(\A[765] ), .ZN(new_n12797_));
  AOI21_X1   g11777(.A1(new_n12795_), .A2(new_n12797_), .B(new_n12796_), .ZN(new_n12798_));
  NAND2_X1   g11778(.A1(new_n12794_), .A2(new_n12798_), .ZN(new_n12799_));
  NOR2_X1    g11779(.A1(new_n12794_), .A2(new_n12798_), .ZN(new_n12800_));
  INV_X1     g11780(.I(\A[764] ), .ZN(new_n12801_));
  NAND2_X1   g11781(.A1(new_n12801_), .A2(\A[765] ), .ZN(new_n12802_));
  INV_X1     g11782(.I(\A[765] ), .ZN(new_n12803_));
  NAND2_X1   g11783(.A1(new_n12803_), .A2(\A[764] ), .ZN(new_n12804_));
  AOI21_X1   g11784(.A1(new_n12802_), .A2(new_n12804_), .B(new_n12795_), .ZN(new_n12805_));
  INV_X1     g11785(.I(new_n12796_), .ZN(new_n12806_));
  AOI21_X1   g11786(.A1(new_n12806_), .A2(new_n12797_), .B(\A[763] ), .ZN(new_n12807_));
  NOR2_X1    g11787(.A1(new_n12807_), .A2(new_n12805_), .ZN(new_n12808_));
  INV_X1     g11788(.I(\A[767] ), .ZN(new_n12809_));
  NAND2_X1   g11789(.A1(new_n12809_), .A2(\A[768] ), .ZN(new_n12810_));
  INV_X1     g11790(.I(\A[768] ), .ZN(new_n12811_));
  NAND2_X1   g11791(.A1(new_n12811_), .A2(\A[767] ), .ZN(new_n12812_));
  AOI21_X1   g11792(.A1(new_n12810_), .A2(new_n12812_), .B(new_n12791_), .ZN(new_n12813_));
  INV_X1     g11793(.I(new_n12792_), .ZN(new_n12814_));
  AOI21_X1   g11794(.A1(new_n12814_), .A2(new_n12793_), .B(\A[766] ), .ZN(new_n12815_));
  NOR2_X1    g11795(.A1(new_n12815_), .A2(new_n12813_), .ZN(new_n12816_));
  NAND2_X1   g11796(.A1(new_n12808_), .A2(new_n12816_), .ZN(new_n12817_));
  OAI21_X1   g11797(.A1(new_n12817_), .A2(new_n12800_), .B(new_n12799_), .ZN(new_n12818_));
  NAND2_X1   g11798(.A1(new_n12790_), .A2(new_n12818_), .ZN(new_n12819_));
  NAND2_X1   g11799(.A1(new_n12789_), .A2(new_n12768_), .ZN(new_n12820_));
  NOR2_X1    g11800(.A1(new_n12775_), .A2(\A[770] ), .ZN(new_n12821_));
  NOR2_X1    g11801(.A1(new_n12773_), .A2(\A[771] ), .ZN(new_n12822_));
  OAI21_X1   g11802(.A1(new_n12821_), .A2(new_n12822_), .B(\A[769] ), .ZN(new_n12823_));
  INV_X1     g11803(.I(new_n12767_), .ZN(new_n12824_));
  OAI21_X1   g11804(.A1(new_n12824_), .A2(new_n12766_), .B(new_n12765_), .ZN(new_n12825_));
  NAND2_X1   g11805(.A1(new_n12823_), .A2(new_n12825_), .ZN(new_n12826_));
  NOR2_X1    g11806(.A1(new_n12783_), .A2(\A[773] ), .ZN(new_n12827_));
  NOR2_X1    g11807(.A1(new_n12781_), .A2(\A[774] ), .ZN(new_n12828_));
  OAI21_X1   g11808(.A1(new_n12827_), .A2(new_n12828_), .B(\A[772] ), .ZN(new_n12829_));
  INV_X1     g11809(.I(new_n12762_), .ZN(new_n12830_));
  OAI21_X1   g11810(.A1(new_n12830_), .A2(new_n12761_), .B(new_n12760_), .ZN(new_n12831_));
  NAND2_X1   g11811(.A1(new_n12829_), .A2(new_n12831_), .ZN(new_n12832_));
  NOR2_X1    g11812(.A1(new_n12826_), .A2(new_n12832_), .ZN(new_n12833_));
  NAND2_X1   g11813(.A1(new_n12833_), .A2(new_n12769_), .ZN(new_n12834_));
  AOI21_X1   g11814(.A1(new_n12834_), .A2(new_n12820_), .B(new_n12764_), .ZN(new_n12835_));
  NOR2_X1    g11815(.A1(new_n12833_), .A2(new_n12769_), .ZN(new_n12836_));
  NOR2_X1    g11816(.A1(new_n12789_), .A2(new_n12768_), .ZN(new_n12837_));
  NOR3_X1    g11817(.A1(new_n12836_), .A2(new_n12837_), .A3(new_n12763_), .ZN(new_n12838_));
  NOR2_X1    g11818(.A1(new_n12835_), .A2(new_n12838_), .ZN(new_n12839_));
  NOR4_X1    g11819(.A1(new_n12805_), .A2(new_n12807_), .A3(new_n12815_), .A4(new_n12813_), .ZN(new_n12840_));
  NAND2_X1   g11820(.A1(new_n12826_), .A2(new_n12832_), .ZN(new_n12841_));
  NAND2_X1   g11821(.A1(new_n12789_), .A2(new_n12841_), .ZN(new_n12842_));
  NAND2_X1   g11822(.A1(new_n12833_), .A2(new_n12770_), .ZN(new_n12843_));
  NOR2_X1    g11823(.A1(new_n12808_), .A2(new_n12816_), .ZN(new_n12844_));
  NOR4_X1    g11824(.A1(new_n12842_), .A2(new_n12843_), .A3(new_n12840_), .A4(new_n12844_), .ZN(new_n12845_));
  NAND2_X1   g11825(.A1(new_n12780_), .A2(new_n12832_), .ZN(new_n12846_));
  NAND2_X1   g11826(.A1(new_n12788_), .A2(new_n12826_), .ZN(new_n12847_));
  AOI21_X1   g11827(.A1(new_n12846_), .A2(new_n12847_), .B(new_n12771_), .ZN(new_n12848_));
  NOR3_X1    g11828(.A1(new_n12848_), .A2(new_n12799_), .A3(new_n12817_), .ZN(new_n12849_));
  INV_X1     g11829(.I(new_n12849_), .ZN(new_n12850_));
  AOI21_X1   g11830(.A1(new_n12839_), .A2(new_n12845_), .B(new_n12850_), .ZN(new_n12851_));
  INV_X1     g11831(.I(new_n12794_), .ZN(new_n12852_));
  INV_X1     g11832(.I(new_n12798_), .ZN(new_n12853_));
  NOR2_X1    g11833(.A1(new_n12840_), .A2(new_n12853_), .ZN(new_n12854_));
  INV_X1     g11834(.I(new_n12854_), .ZN(new_n12855_));
  NAND2_X1   g11835(.A1(new_n12840_), .A2(new_n12853_), .ZN(new_n12856_));
  AOI21_X1   g11836(.A1(new_n12855_), .A2(new_n12856_), .B(new_n12852_), .ZN(new_n12857_));
  INV_X1     g11837(.I(new_n12856_), .ZN(new_n12858_));
  NOR3_X1    g11838(.A1(new_n12858_), .A2(new_n12794_), .A3(new_n12854_), .ZN(new_n12859_));
  NOR2_X1    g11839(.A1(new_n12857_), .A2(new_n12859_), .ZN(new_n12860_));
  NOR3_X1    g11840(.A1(new_n12835_), .A2(new_n12838_), .A3(new_n12848_), .ZN(new_n12861_));
  NOR2_X1    g11841(.A1(new_n12842_), .A2(new_n12843_), .ZN(new_n12862_));
  NOR2_X1    g11842(.A1(new_n12844_), .A2(new_n12840_), .ZN(new_n12863_));
  NOR2_X1    g11843(.A1(new_n12817_), .A2(new_n12799_), .ZN(new_n12864_));
  NAND2_X1   g11844(.A1(new_n12863_), .A2(new_n12864_), .ZN(new_n12865_));
  INV_X1     g11845(.I(new_n12865_), .ZN(new_n12866_));
  NAND2_X1   g11846(.A1(new_n12866_), .A2(new_n12862_), .ZN(new_n12867_));
  NOR2_X1    g11847(.A1(new_n12867_), .A2(new_n12861_), .ZN(new_n12868_));
  NOR2_X1    g11848(.A1(new_n12868_), .A2(new_n12860_), .ZN(new_n12869_));
  NOR2_X1    g11849(.A1(new_n12869_), .A2(new_n12851_), .ZN(new_n12870_));
  OAI21_X1   g11850(.A1(new_n12790_), .A2(new_n12818_), .B(new_n12870_), .ZN(new_n12871_));
  NAND2_X1   g11851(.A1(new_n12871_), .A2(new_n12819_), .ZN(new_n12872_));
  INV_X1     g11852(.I(\A[760] ), .ZN(new_n12873_));
  NOR2_X1    g11853(.A1(\A[761] ), .A2(\A[762] ), .ZN(new_n12874_));
  NAND2_X1   g11854(.A1(\A[761] ), .A2(\A[762] ), .ZN(new_n12875_));
  AOI21_X1   g11855(.A1(new_n12873_), .A2(new_n12875_), .B(new_n12874_), .ZN(new_n12876_));
  INV_X1     g11856(.I(new_n12876_), .ZN(new_n12877_));
  INV_X1     g11857(.I(\A[757] ), .ZN(new_n12878_));
  NOR2_X1    g11858(.A1(\A[758] ), .A2(\A[759] ), .ZN(new_n12879_));
  NAND2_X1   g11859(.A1(\A[758] ), .A2(\A[759] ), .ZN(new_n12880_));
  AOI21_X1   g11860(.A1(new_n12878_), .A2(new_n12880_), .B(new_n12879_), .ZN(new_n12881_));
  INV_X1     g11861(.I(new_n12881_), .ZN(new_n12882_));
  NOR2_X1    g11862(.A1(new_n12877_), .A2(new_n12882_), .ZN(new_n12883_));
  INV_X1     g11863(.I(new_n12883_), .ZN(new_n12884_));
  NOR2_X1    g11864(.A1(new_n12876_), .A2(new_n12881_), .ZN(new_n12885_));
  INV_X1     g11865(.I(\A[758] ), .ZN(new_n12886_));
  NAND2_X1   g11866(.A1(new_n12886_), .A2(\A[759] ), .ZN(new_n12887_));
  INV_X1     g11867(.I(\A[759] ), .ZN(new_n12888_));
  NAND2_X1   g11868(.A1(new_n12888_), .A2(\A[758] ), .ZN(new_n12889_));
  AOI21_X1   g11869(.A1(new_n12887_), .A2(new_n12889_), .B(new_n12878_), .ZN(new_n12890_));
  INV_X1     g11870(.I(new_n12879_), .ZN(new_n12891_));
  AOI21_X1   g11871(.A1(new_n12891_), .A2(new_n12880_), .B(\A[757] ), .ZN(new_n12892_));
  NOR2_X1    g11872(.A1(new_n12892_), .A2(new_n12890_), .ZN(new_n12893_));
  INV_X1     g11873(.I(\A[761] ), .ZN(new_n12894_));
  NAND2_X1   g11874(.A1(new_n12894_), .A2(\A[762] ), .ZN(new_n12895_));
  INV_X1     g11875(.I(\A[762] ), .ZN(new_n12896_));
  NAND2_X1   g11876(.A1(new_n12896_), .A2(\A[761] ), .ZN(new_n12897_));
  AOI21_X1   g11877(.A1(new_n12895_), .A2(new_n12897_), .B(new_n12873_), .ZN(new_n12898_));
  INV_X1     g11878(.I(new_n12874_), .ZN(new_n12899_));
  AOI21_X1   g11879(.A1(new_n12899_), .A2(new_n12875_), .B(\A[760] ), .ZN(new_n12900_));
  NOR2_X1    g11880(.A1(new_n12900_), .A2(new_n12898_), .ZN(new_n12901_));
  NAND2_X1   g11881(.A1(new_n12893_), .A2(new_n12901_), .ZN(new_n12902_));
  OAI21_X1   g11882(.A1(new_n12902_), .A2(new_n12885_), .B(new_n12884_), .ZN(new_n12903_));
  INV_X1     g11883(.I(\A[754] ), .ZN(new_n12904_));
  NOR2_X1    g11884(.A1(\A[755] ), .A2(\A[756] ), .ZN(new_n12905_));
  NAND2_X1   g11885(.A1(\A[755] ), .A2(\A[756] ), .ZN(new_n12906_));
  AOI21_X1   g11886(.A1(new_n12904_), .A2(new_n12906_), .B(new_n12905_), .ZN(new_n12907_));
  INV_X1     g11887(.I(\A[751] ), .ZN(new_n12908_));
  NOR2_X1    g11888(.A1(\A[752] ), .A2(\A[753] ), .ZN(new_n12909_));
  NAND2_X1   g11889(.A1(\A[752] ), .A2(\A[753] ), .ZN(new_n12910_));
  AOI21_X1   g11890(.A1(new_n12908_), .A2(new_n12910_), .B(new_n12909_), .ZN(new_n12911_));
  NAND2_X1   g11891(.A1(new_n12907_), .A2(new_n12911_), .ZN(new_n12912_));
  NOR2_X1    g11892(.A1(new_n12907_), .A2(new_n12911_), .ZN(new_n12913_));
  INV_X1     g11893(.I(\A[752] ), .ZN(new_n12914_));
  NAND2_X1   g11894(.A1(new_n12914_), .A2(\A[753] ), .ZN(new_n12915_));
  INV_X1     g11895(.I(\A[753] ), .ZN(new_n12916_));
  NAND2_X1   g11896(.A1(new_n12916_), .A2(\A[752] ), .ZN(new_n12917_));
  AOI21_X1   g11897(.A1(new_n12915_), .A2(new_n12917_), .B(new_n12908_), .ZN(new_n12918_));
  INV_X1     g11898(.I(new_n12909_), .ZN(new_n12919_));
  AOI21_X1   g11899(.A1(new_n12919_), .A2(new_n12910_), .B(\A[751] ), .ZN(new_n12920_));
  NOR2_X1    g11900(.A1(new_n12920_), .A2(new_n12918_), .ZN(new_n12921_));
  INV_X1     g11901(.I(\A[755] ), .ZN(new_n12922_));
  NAND2_X1   g11902(.A1(new_n12922_), .A2(\A[756] ), .ZN(new_n12923_));
  INV_X1     g11903(.I(\A[756] ), .ZN(new_n12924_));
  NAND2_X1   g11904(.A1(new_n12924_), .A2(\A[755] ), .ZN(new_n12925_));
  AOI21_X1   g11905(.A1(new_n12923_), .A2(new_n12925_), .B(new_n12904_), .ZN(new_n12926_));
  INV_X1     g11906(.I(new_n12905_), .ZN(new_n12927_));
  AOI21_X1   g11907(.A1(new_n12927_), .A2(new_n12906_), .B(\A[754] ), .ZN(new_n12928_));
  NOR2_X1    g11908(.A1(new_n12928_), .A2(new_n12926_), .ZN(new_n12929_));
  NAND2_X1   g11909(.A1(new_n12921_), .A2(new_n12929_), .ZN(new_n12930_));
  OAI21_X1   g11910(.A1(new_n12930_), .A2(new_n12913_), .B(new_n12912_), .ZN(new_n12931_));
  NAND2_X1   g11911(.A1(new_n12903_), .A2(new_n12931_), .ZN(new_n12932_));
  NOR2_X1    g11912(.A1(new_n12888_), .A2(\A[758] ), .ZN(new_n12933_));
  NOR2_X1    g11913(.A1(new_n12886_), .A2(\A[759] ), .ZN(new_n12934_));
  OAI21_X1   g11914(.A1(new_n12933_), .A2(new_n12934_), .B(\A[757] ), .ZN(new_n12935_));
  INV_X1     g11915(.I(new_n12880_), .ZN(new_n12936_));
  OAI21_X1   g11916(.A1(new_n12936_), .A2(new_n12879_), .B(new_n12878_), .ZN(new_n12937_));
  NAND2_X1   g11917(.A1(new_n12935_), .A2(new_n12937_), .ZN(new_n12938_));
  NOR2_X1    g11918(.A1(new_n12896_), .A2(\A[761] ), .ZN(new_n12939_));
  NOR2_X1    g11919(.A1(new_n12894_), .A2(\A[762] ), .ZN(new_n12940_));
  OAI21_X1   g11920(.A1(new_n12939_), .A2(new_n12940_), .B(\A[760] ), .ZN(new_n12941_));
  INV_X1     g11921(.I(new_n12875_), .ZN(new_n12942_));
  OAI21_X1   g11922(.A1(new_n12942_), .A2(new_n12874_), .B(new_n12873_), .ZN(new_n12943_));
  NAND2_X1   g11923(.A1(new_n12941_), .A2(new_n12943_), .ZN(new_n12944_));
  NOR2_X1    g11924(.A1(new_n12938_), .A2(new_n12944_), .ZN(new_n12945_));
  NOR2_X1    g11925(.A1(new_n12945_), .A2(new_n12882_), .ZN(new_n12946_));
  NOR2_X1    g11926(.A1(new_n12902_), .A2(new_n12881_), .ZN(new_n12947_));
  OAI21_X1   g11927(.A1(new_n12946_), .A2(new_n12947_), .B(new_n12876_), .ZN(new_n12948_));
  NAND2_X1   g11928(.A1(new_n12902_), .A2(new_n12881_), .ZN(new_n12949_));
  NAND2_X1   g11929(.A1(new_n12945_), .A2(new_n12882_), .ZN(new_n12950_));
  NAND3_X1   g11930(.A1(new_n12950_), .A2(new_n12949_), .A3(new_n12877_), .ZN(new_n12951_));
  NAND2_X1   g11931(.A1(new_n12948_), .A2(new_n12951_), .ZN(new_n12952_));
  NAND2_X1   g11932(.A1(new_n12938_), .A2(new_n12944_), .ZN(new_n12953_));
  NAND2_X1   g11933(.A1(new_n12902_), .A2(new_n12953_), .ZN(new_n12954_));
  NAND2_X1   g11934(.A1(new_n12945_), .A2(new_n12883_), .ZN(new_n12955_));
  NOR2_X1    g11935(.A1(new_n12916_), .A2(\A[752] ), .ZN(new_n12956_));
  NOR2_X1    g11936(.A1(new_n12914_), .A2(\A[753] ), .ZN(new_n12957_));
  OAI21_X1   g11937(.A1(new_n12956_), .A2(new_n12957_), .B(\A[751] ), .ZN(new_n12958_));
  INV_X1     g11938(.I(new_n12910_), .ZN(new_n12959_));
  OAI21_X1   g11939(.A1(new_n12959_), .A2(new_n12909_), .B(new_n12908_), .ZN(new_n12960_));
  NAND2_X1   g11940(.A1(new_n12958_), .A2(new_n12960_), .ZN(new_n12961_));
  NOR2_X1    g11941(.A1(new_n12924_), .A2(\A[755] ), .ZN(new_n12962_));
  NOR2_X1    g11942(.A1(new_n12922_), .A2(\A[756] ), .ZN(new_n12963_));
  OAI21_X1   g11943(.A1(new_n12962_), .A2(new_n12963_), .B(\A[754] ), .ZN(new_n12964_));
  INV_X1     g11944(.I(new_n12906_), .ZN(new_n12965_));
  OAI21_X1   g11945(.A1(new_n12965_), .A2(new_n12905_), .B(new_n12904_), .ZN(new_n12966_));
  NAND2_X1   g11946(.A1(new_n12964_), .A2(new_n12966_), .ZN(new_n12967_));
  NAND2_X1   g11947(.A1(new_n12961_), .A2(new_n12967_), .ZN(new_n12968_));
  NAND2_X1   g11948(.A1(new_n12930_), .A2(new_n12968_), .ZN(new_n12969_));
  NOR3_X1    g11949(.A1(new_n12954_), .A2(new_n12969_), .A3(new_n12955_), .ZN(new_n12970_));
  INV_X1     g11950(.I(new_n12970_), .ZN(new_n12971_));
  NAND4_X1   g11951(.A1(new_n12921_), .A2(new_n12929_), .A3(new_n12907_), .A4(new_n12911_), .ZN(new_n12972_));
  NAND2_X1   g11952(.A1(new_n12893_), .A2(new_n12944_), .ZN(new_n12973_));
  NAND2_X1   g11953(.A1(new_n12901_), .A2(new_n12938_), .ZN(new_n12974_));
  AOI21_X1   g11954(.A1(new_n12973_), .A2(new_n12974_), .B(new_n12884_), .ZN(new_n12975_));
  NOR2_X1    g11955(.A1(new_n12975_), .A2(new_n12972_), .ZN(new_n12976_));
  OAI21_X1   g11956(.A1(new_n12952_), .A2(new_n12971_), .B(new_n12976_), .ZN(new_n12977_));
  INV_X1     g11957(.I(new_n12911_), .ZN(new_n12978_));
  NOR2_X1    g11958(.A1(new_n12961_), .A2(new_n12967_), .ZN(new_n12979_));
  NOR2_X1    g11959(.A1(new_n12979_), .A2(new_n12978_), .ZN(new_n12980_));
  NOR2_X1    g11960(.A1(new_n12930_), .A2(new_n12911_), .ZN(new_n12981_));
  OAI21_X1   g11961(.A1(new_n12980_), .A2(new_n12981_), .B(new_n12907_), .ZN(new_n12982_));
  INV_X1     g11962(.I(new_n12907_), .ZN(new_n12983_));
  NAND2_X1   g11963(.A1(new_n12930_), .A2(new_n12911_), .ZN(new_n12984_));
  NAND2_X1   g11964(.A1(new_n12979_), .A2(new_n12978_), .ZN(new_n12985_));
  NAND3_X1   g11965(.A1(new_n12985_), .A2(new_n12984_), .A3(new_n12983_), .ZN(new_n12986_));
  NAND2_X1   g11966(.A1(new_n12982_), .A2(new_n12986_), .ZN(new_n12987_));
  AOI21_X1   g11967(.A1(new_n12950_), .A2(new_n12949_), .B(new_n12877_), .ZN(new_n12988_));
  NOR3_X1    g11968(.A1(new_n12946_), .A2(new_n12947_), .A3(new_n12876_), .ZN(new_n12989_));
  NOR3_X1    g11969(.A1(new_n12988_), .A2(new_n12989_), .A3(new_n12975_), .ZN(new_n12990_));
  NOR2_X1    g11970(.A1(new_n12954_), .A2(new_n12955_), .ZN(new_n12991_));
  NOR2_X1    g11971(.A1(new_n12969_), .A2(new_n12972_), .ZN(new_n12992_));
  NAND2_X1   g11972(.A1(new_n12991_), .A2(new_n12992_), .ZN(new_n12993_));
  OAI21_X1   g11973(.A1(new_n12990_), .A2(new_n12993_), .B(new_n12987_), .ZN(new_n12994_));
  AND2_X2    g11974(.A1(new_n12994_), .A2(new_n12977_), .Z(new_n12995_));
  OAI21_X1   g11975(.A1(new_n12903_), .A2(new_n12931_), .B(new_n12995_), .ZN(new_n12996_));
  NAND2_X1   g11976(.A1(new_n12996_), .A2(new_n12932_), .ZN(new_n12997_));
  NAND2_X1   g11977(.A1(new_n12872_), .A2(new_n12997_), .ZN(new_n12998_));
  OAI21_X1   g11978(.A1(new_n12836_), .A2(new_n12837_), .B(new_n12763_), .ZN(new_n12999_));
  NAND3_X1   g11979(.A1(new_n12834_), .A2(new_n12820_), .A3(new_n12764_), .ZN(new_n13000_));
  INV_X1     g11980(.I(new_n12848_), .ZN(new_n13001_));
  NAND3_X1   g11981(.A1(new_n12999_), .A2(new_n13000_), .A3(new_n13001_), .ZN(new_n13002_));
  NOR2_X1    g11982(.A1(new_n12867_), .A2(new_n13002_), .ZN(new_n13003_));
  OR2_X2     g11983(.A1(new_n12842_), .A2(new_n12843_), .Z(new_n13004_));
  NOR2_X1    g11984(.A1(new_n13004_), .A2(new_n12865_), .ZN(new_n13005_));
  NOR2_X1    g11985(.A1(new_n13005_), .A2(new_n12861_), .ZN(new_n13006_));
  OAI21_X1   g11986(.A1(new_n13003_), .A2(new_n13006_), .B(new_n12860_), .ZN(new_n13007_));
  NAND2_X1   g11987(.A1(new_n12999_), .A2(new_n13000_), .ZN(new_n13008_));
  INV_X1     g11988(.I(new_n12845_), .ZN(new_n13009_));
  OAI21_X1   g11989(.A1(new_n13008_), .A2(new_n13009_), .B(new_n12849_), .ZN(new_n13010_));
  NAND2_X1   g11990(.A1(new_n13005_), .A2(new_n13002_), .ZN(new_n13011_));
  NAND3_X1   g11991(.A1(new_n13011_), .A2(new_n13010_), .A3(new_n12860_), .ZN(new_n13012_));
  NAND2_X1   g11992(.A1(new_n13007_), .A2(new_n13012_), .ZN(new_n13013_));
  INV_X1     g11993(.I(new_n12860_), .ZN(new_n13014_));
  NAND2_X1   g11994(.A1(new_n13005_), .A2(new_n12861_), .ZN(new_n13015_));
  NAND2_X1   g11995(.A1(new_n12867_), .A2(new_n13002_), .ZN(new_n13016_));
  AOI21_X1   g11996(.A1(new_n13016_), .A2(new_n13015_), .B(new_n13014_), .ZN(new_n13017_));
  NOR3_X1    g11997(.A1(new_n12868_), .A2(new_n12851_), .A3(new_n13014_), .ZN(new_n13018_));
  NOR2_X1    g11998(.A1(new_n12865_), .A2(new_n12862_), .ZN(new_n13019_));
  INV_X1     g11999(.I(new_n13019_), .ZN(new_n13020_));
  NAND2_X1   g12000(.A1(new_n12865_), .A2(new_n12862_), .ZN(new_n13021_));
  INV_X1     g12001(.I(new_n12991_), .ZN(new_n13022_));
  NAND2_X1   g12002(.A1(new_n13022_), .A2(new_n12992_), .ZN(new_n13023_));
  INV_X1     g12003(.I(new_n12972_), .ZN(new_n13024_));
  NAND3_X1   g12004(.A1(new_n13024_), .A2(new_n12930_), .A3(new_n12968_), .ZN(new_n13025_));
  NAND2_X1   g12005(.A1(new_n13025_), .A2(new_n12991_), .ZN(new_n13026_));
  NAND4_X1   g12006(.A1(new_n13020_), .A2(new_n13023_), .A3(new_n13026_), .A4(new_n13021_), .ZN(new_n13027_));
  OAI21_X1   g12007(.A1(new_n13017_), .A2(new_n13018_), .B(new_n13027_), .ZN(new_n13028_));
  INV_X1     g12008(.I(new_n13027_), .ZN(new_n13029_));
  NAND3_X1   g12009(.A1(new_n13007_), .A2(new_n13029_), .A3(new_n13012_), .ZN(new_n13030_));
  NOR2_X1    g12010(.A1(new_n12988_), .A2(new_n12989_), .ZN(new_n13031_));
  NAND2_X1   g12011(.A1(new_n13031_), .A2(new_n12970_), .ZN(new_n13032_));
  NAND3_X1   g12012(.A1(new_n13032_), .A2(new_n12976_), .A3(new_n12987_), .ZN(new_n13033_));
  NAND2_X1   g12013(.A1(new_n12987_), .A2(new_n12993_), .ZN(new_n13034_));
  AND2_X2    g12014(.A1(new_n12982_), .A2(new_n12986_), .Z(new_n13035_));
  NOR2_X1    g12015(.A1(new_n13022_), .A2(new_n13025_), .ZN(new_n13036_));
  AOI21_X1   g12016(.A1(new_n13035_), .A2(new_n13036_), .B(new_n12990_), .ZN(new_n13037_));
  NAND4_X1   g12017(.A1(new_n12982_), .A2(new_n12986_), .A3(new_n12991_), .A4(new_n12992_), .ZN(new_n13038_));
  NOR3_X1    g12018(.A1(new_n13038_), .A2(new_n12952_), .A3(new_n12975_), .ZN(new_n13039_));
  OAI21_X1   g12019(.A1(new_n13037_), .A2(new_n13039_), .B(new_n13034_), .ZN(new_n13040_));
  NAND2_X1   g12020(.A1(new_n13040_), .A2(new_n13033_), .ZN(new_n13041_));
  AOI22_X1   g12021(.A1(new_n13028_), .A2(new_n13030_), .B1(new_n13041_), .B2(new_n13013_), .ZN(new_n13042_));
  XNOR2_X1   g12022(.A1(new_n12790_), .A2(new_n12818_), .ZN(new_n13043_));
  INV_X1     g12023(.I(new_n13043_), .ZN(new_n13044_));
  NOR3_X1    g12024(.A1(new_n12869_), .A2(new_n12851_), .A3(new_n13044_), .ZN(new_n13045_));
  XNOR2_X1   g12025(.A1(new_n12903_), .A2(new_n12931_), .ZN(new_n13046_));
  NAND3_X1   g12026(.A1(new_n12994_), .A2(new_n12977_), .A3(new_n13046_), .ZN(new_n13047_));
  INV_X1     g12027(.I(new_n13047_), .ZN(new_n13048_));
  NAND3_X1   g12028(.A1(new_n13042_), .A2(new_n13045_), .A3(new_n13048_), .ZN(new_n13049_));
  OAI21_X1   g12029(.A1(new_n12872_), .A2(new_n12997_), .B(new_n13049_), .ZN(new_n13050_));
  NAND2_X1   g12030(.A1(new_n13050_), .A2(new_n12998_), .ZN(new_n13051_));
  INV_X1     g12031(.I(new_n13051_), .ZN(new_n13052_));
  NOR2_X1    g12032(.A1(new_n12759_), .A2(new_n13052_), .ZN(new_n13053_));
  NOR2_X1    g12033(.A1(new_n13017_), .A2(new_n13018_), .ZN(new_n13054_));
  AOI21_X1   g12034(.A1(new_n13007_), .A2(new_n13012_), .B(new_n13029_), .ZN(new_n13055_));
  NOR3_X1    g12035(.A1(new_n13017_), .A2(new_n13018_), .A3(new_n13027_), .ZN(new_n13056_));
  NOR2_X1    g12036(.A1(new_n12977_), .A2(new_n13035_), .ZN(new_n13057_));
  XOR2_X1    g12037(.A1(new_n13038_), .A2(new_n12990_), .Z(new_n13058_));
  AOI21_X1   g12038(.A1(new_n13058_), .A2(new_n13034_), .B(new_n13057_), .ZN(new_n13059_));
  OAI22_X1   g12039(.A1(new_n13055_), .A2(new_n13056_), .B1(new_n13059_), .B2(new_n13054_), .ZN(new_n13060_));
  NAND2_X1   g12040(.A1(new_n13011_), .A2(new_n13014_), .ZN(new_n13061_));
  NAND3_X1   g12041(.A1(new_n13061_), .A2(new_n13010_), .A3(new_n13043_), .ZN(new_n13062_));
  XOR2_X1    g12042(.A1(new_n13062_), .A2(new_n13048_), .Z(new_n13063_));
  NAND2_X1   g12043(.A1(new_n13062_), .A2(new_n13047_), .ZN(new_n13064_));
  NAND2_X1   g12044(.A1(new_n13045_), .A2(new_n13048_), .ZN(new_n13065_));
  NAND2_X1   g12045(.A1(new_n13065_), .A2(new_n13064_), .ZN(new_n13066_));
  NAND2_X1   g12046(.A1(new_n13060_), .A2(new_n13066_), .ZN(new_n13067_));
  OAI21_X1   g12047(.A1(new_n13060_), .A2(new_n13063_), .B(new_n13067_), .ZN(new_n13068_));
  INV_X1     g12048(.I(new_n12707_), .ZN(new_n13069_));
  INV_X1     g12049(.I(new_n12719_), .ZN(new_n13070_));
  NAND2_X1   g12050(.A1(new_n12721_), .A2(new_n12691_), .ZN(new_n13071_));
  AND2_X2    g12051(.A1(new_n12727_), .A2(new_n13071_), .Z(new_n13072_));
  OAI22_X1   g12052(.A1(new_n13072_), .A2(new_n13069_), .B1(new_n13070_), .B2(new_n12717_), .ZN(new_n13073_));
  AOI21_X1   g12053(.A1(new_n12747_), .A2(new_n12744_), .B(new_n12626_), .ZN(new_n13074_));
  NOR3_X1    g12054(.A1(new_n12745_), .A2(new_n12742_), .A3(new_n12743_), .ZN(new_n13075_));
  NOR2_X1    g12055(.A1(new_n13074_), .A2(new_n13075_), .ZN(new_n13076_));
  NAND2_X1   g12056(.A1(new_n13076_), .A2(new_n12741_), .ZN(new_n13077_));
  AOI21_X1   g12057(.A1(new_n12738_), .A2(new_n12739_), .B(new_n12534_), .ZN(new_n13078_));
  NOR3_X1    g12058(.A1(new_n12731_), .A2(new_n12736_), .A3(new_n12535_), .ZN(new_n13079_));
  NOR2_X1    g12059(.A1(new_n13078_), .A2(new_n13079_), .ZN(new_n13080_));
  NAND2_X1   g12060(.A1(new_n12749_), .A2(new_n13080_), .ZN(new_n13081_));
  AOI21_X1   g12061(.A1(new_n13081_), .A2(new_n13077_), .B(new_n13073_), .ZN(new_n13082_));
  NAND2_X1   g12062(.A1(new_n13076_), .A2(new_n13080_), .ZN(new_n13083_));
  NAND2_X1   g12063(.A1(new_n12749_), .A2(new_n12741_), .ZN(new_n13084_));
  AOI21_X1   g12064(.A1(new_n13083_), .A2(new_n13084_), .B(new_n12729_), .ZN(new_n13085_));
  NOR3_X1    g12065(.A1(new_n13068_), .A2(new_n13082_), .A3(new_n13085_), .ZN(new_n13086_));
  INV_X1     g12066(.I(new_n12872_), .ZN(new_n13087_));
  NAND2_X1   g12067(.A1(new_n13049_), .A2(new_n12997_), .ZN(new_n13088_));
  INV_X1     g12068(.I(new_n12997_), .ZN(new_n13089_));
  NAND4_X1   g12069(.A1(new_n13089_), .A2(new_n13042_), .A3(new_n13045_), .A4(new_n13048_), .ZN(new_n13090_));
  AOI21_X1   g12070(.A1(new_n13088_), .A2(new_n13090_), .B(new_n13087_), .ZN(new_n13091_));
  NAND2_X1   g12071(.A1(new_n13060_), .A2(new_n13064_), .ZN(new_n13092_));
  INV_X1     g12072(.I(new_n13065_), .ZN(new_n13093_));
  AOI21_X1   g12073(.A1(new_n13092_), .A2(new_n13093_), .B(new_n13089_), .ZN(new_n13094_));
  NOR2_X1    g12074(.A1(new_n13049_), .A2(new_n12997_), .ZN(new_n13095_));
  NOR3_X1    g12075(.A1(new_n13094_), .A2(new_n13095_), .A3(new_n12872_), .ZN(new_n13096_));
  XNOR2_X1   g12076(.A1(new_n12695_), .A2(new_n12598_), .ZN(new_n13097_));
  NOR2_X1    g12077(.A1(new_n12755_), .A2(new_n13097_), .ZN(new_n13098_));
  NOR3_X1    g12078(.A1(new_n13096_), .A2(new_n13091_), .A3(new_n13098_), .ZN(new_n13099_));
  NAND2_X1   g12079(.A1(new_n13083_), .A2(new_n13073_), .ZN(new_n13100_));
  XOR2_X1    g12080(.A1(new_n12695_), .A2(new_n12598_), .Z(new_n13101_));
  NAND3_X1   g12081(.A1(new_n13100_), .A2(new_n12754_), .A3(new_n13101_), .ZN(new_n13102_));
  XOR2_X1    g12082(.A1(new_n12872_), .A2(new_n12997_), .Z(new_n13103_));
  NOR3_X1    g12083(.A1(new_n13102_), .A2(new_n13049_), .A3(new_n13103_), .ZN(new_n13104_));
  OAI21_X1   g12084(.A1(new_n13099_), .A2(new_n13086_), .B(new_n13104_), .ZN(new_n13105_));
  INV_X1     g12085(.I(new_n13105_), .ZN(new_n13106_));
  NAND4_X1   g12086(.A1(new_n12756_), .A2(new_n12757_), .A3(new_n12998_), .A4(new_n13050_), .ZN(new_n13107_));
  NOR2_X1    g12087(.A1(new_n13106_), .A2(new_n13107_), .ZN(new_n13108_));
  NOR2_X1    g12088(.A1(new_n13108_), .A2(new_n13053_), .ZN(new_n13109_));
  NAND2_X1   g12089(.A1(new_n12504_), .A2(new_n13109_), .ZN(new_n13110_));
  OAI21_X1   g12090(.A1(new_n12504_), .A2(new_n13053_), .B(new_n13108_), .ZN(new_n13111_));
  NAND4_X1   g12091(.A1(new_n12147_), .A2(new_n12427_), .A3(new_n12414_), .A4(new_n12162_), .ZN(new_n13112_));
  OAI21_X1   g12092(.A1(new_n12436_), .A2(new_n12395_), .B(new_n12433_), .ZN(new_n13113_));
  NAND3_X1   g12093(.A1(new_n12430_), .A2(new_n12434_), .A3(new_n12421_), .ZN(new_n13114_));
  NAND2_X1   g12094(.A1(new_n13114_), .A2(new_n13113_), .ZN(new_n13115_));
  OAI21_X1   g12095(.A1(new_n12439_), .A2(new_n12443_), .B(new_n13115_), .ZN(new_n13116_));
  XNOR2_X1   g12096(.A1(new_n12138_), .A2(new_n12145_), .ZN(new_n13117_));
  NOR2_X1    g12097(.A1(new_n13117_), .A2(new_n12155_), .ZN(new_n13118_));
  NOR2_X1    g12098(.A1(new_n12138_), .A2(new_n12145_), .ZN(new_n13119_));
  NOR2_X1    g12099(.A1(new_n12452_), .A2(new_n13119_), .ZN(new_n13120_));
  NOR2_X1    g12100(.A1(new_n12130_), .A2(new_n13120_), .ZN(new_n13121_));
  NOR2_X1    g12101(.A1(new_n13118_), .A2(new_n13121_), .ZN(new_n13122_));
  NAND2_X1   g12102(.A1(new_n12424_), .A2(new_n12412_), .ZN(new_n13123_));
  NAND2_X1   g12103(.A1(new_n12479_), .A2(new_n12403_), .ZN(new_n13124_));
  AOI22_X1   g12104(.A1(new_n12422_), .A2(new_n12415_), .B1(new_n13124_), .B2(new_n13123_), .ZN(new_n13125_));
  AOI21_X1   g12105(.A1(new_n12423_), .A2(new_n12425_), .B(new_n12396_), .ZN(new_n13126_));
  NOR2_X1    g12106(.A1(new_n13126_), .A2(new_n13125_), .ZN(new_n13127_));
  NOR2_X1    g12107(.A1(new_n13127_), .A2(new_n13122_), .ZN(new_n13128_));
  OAI21_X1   g12108(.A1(new_n13128_), .A2(new_n13116_), .B(new_n13112_), .ZN(new_n13129_));
  AOI21_X1   g12109(.A1(new_n12464_), .A2(new_n12465_), .B(new_n12463_), .ZN(new_n13130_));
  NOR3_X1    g12110(.A1(new_n12459_), .A2(new_n12461_), .A3(new_n12451_), .ZN(new_n13131_));
  NOR2_X1    g12111(.A1(new_n13131_), .A2(new_n13130_), .ZN(new_n13132_));
  NAND2_X1   g12112(.A1(new_n12482_), .A2(new_n12486_), .ZN(new_n13133_));
  NOR2_X1    g12113(.A1(new_n13132_), .A2(new_n13133_), .ZN(new_n13134_));
  NAND2_X1   g12114(.A1(new_n12462_), .A2(new_n12466_), .ZN(new_n13135_));
  AOI21_X1   g12115(.A1(new_n12485_), .A2(new_n12480_), .B(new_n12470_), .ZN(new_n13136_));
  NOR3_X1    g12116(.A1(new_n12481_), .A2(new_n12478_), .A3(new_n12471_), .ZN(new_n13137_));
  NOR2_X1    g12117(.A1(new_n13137_), .A2(new_n13136_), .ZN(new_n13138_));
  NOR2_X1    g12118(.A1(new_n13135_), .A2(new_n13138_), .ZN(new_n13139_));
  OAI21_X1   g12119(.A1(new_n13139_), .A2(new_n13134_), .B(new_n13129_), .ZN(new_n13140_));
  NOR2_X1    g12120(.A1(new_n13135_), .A2(new_n13133_), .ZN(new_n13141_));
  AOI22_X1   g12121(.A1(new_n12462_), .A2(new_n12466_), .B1(new_n12482_), .B2(new_n12486_), .ZN(new_n13142_));
  OAI21_X1   g12122(.A1(new_n13141_), .A2(new_n13142_), .B(new_n12447_), .ZN(new_n13143_));
  NAND2_X1   g12123(.A1(new_n13140_), .A2(new_n13143_), .ZN(new_n13144_));
  NOR2_X1    g12124(.A1(new_n13063_), .A2(new_n13060_), .ZN(new_n13145_));
  AOI21_X1   g12125(.A1(new_n13064_), .A2(new_n13065_), .B(new_n13042_), .ZN(new_n13146_));
  NOR2_X1    g12126(.A1(new_n13146_), .A2(new_n13145_), .ZN(new_n13147_));
  NOR2_X1    g12127(.A1(new_n12749_), .A2(new_n13080_), .ZN(new_n13148_));
  NOR2_X1    g12128(.A1(new_n13076_), .A2(new_n12741_), .ZN(new_n13149_));
  OAI21_X1   g12129(.A1(new_n13148_), .A2(new_n13149_), .B(new_n12729_), .ZN(new_n13150_));
  NOR2_X1    g12130(.A1(new_n13076_), .A2(new_n13080_), .ZN(new_n13151_));
  OAI21_X1   g12131(.A1(new_n13151_), .A2(new_n12750_), .B(new_n13073_), .ZN(new_n13152_));
  NAND3_X1   g12132(.A1(new_n13147_), .A2(new_n13150_), .A3(new_n13152_), .ZN(new_n13153_));
  OAI21_X1   g12133(.A1(new_n13082_), .A2(new_n13085_), .B(new_n13068_), .ZN(new_n13154_));
  NAND2_X1   g12134(.A1(new_n13154_), .A2(new_n13153_), .ZN(new_n13155_));
  NAND2_X1   g12135(.A1(new_n12428_), .A2(new_n13122_), .ZN(new_n13156_));
  NAND2_X1   g12136(.A1(new_n13127_), .A2(new_n12163_), .ZN(new_n13157_));
  AOI21_X1   g12137(.A1(new_n13156_), .A2(new_n13157_), .B(new_n13116_), .ZN(new_n13158_));
  AOI21_X1   g12138(.A1(new_n12446_), .A2(new_n13112_), .B(new_n12445_), .ZN(new_n13159_));
  NOR3_X1    g12139(.A1(new_n13155_), .A2(new_n13158_), .A3(new_n13159_), .ZN(new_n13160_));
  NAND2_X1   g12140(.A1(new_n12438_), .A2(new_n12443_), .ZN(new_n13161_));
  INV_X1     g12141(.I(new_n12714_), .ZN(new_n13162_));
  XNOR2_X1   g12142(.A1(new_n12709_), .A2(new_n12713_), .ZN(new_n13163_));
  NOR2_X1    g12143(.A1(new_n13163_), .A2(new_n13162_), .ZN(new_n13164_));
  XOR2_X1    g12144(.A1(new_n12709_), .A2(new_n12713_), .Z(new_n13165_));
  NOR2_X1    g12145(.A1(new_n13165_), .A2(new_n12714_), .ZN(new_n13166_));
  OAI21_X1   g12146(.A1(new_n13164_), .A2(new_n13166_), .B(new_n12711_), .ZN(new_n13167_));
  NOR3_X1    g12147(.A1(new_n13164_), .A2(new_n13166_), .A3(new_n12711_), .ZN(new_n13168_));
  INV_X1     g12148(.I(new_n13168_), .ZN(new_n13169_));
  NAND2_X1   g12149(.A1(new_n13020_), .A2(new_n13021_), .ZN(new_n13170_));
  NAND2_X1   g12150(.A1(new_n13023_), .A2(new_n13026_), .ZN(new_n13171_));
  NAND2_X1   g12151(.A1(new_n13170_), .A2(new_n13171_), .ZN(new_n13172_));
  NAND2_X1   g12152(.A1(new_n13172_), .A2(new_n13027_), .ZN(new_n13173_));
  INV_X1     g12153(.I(new_n13173_), .ZN(new_n13174_));
  NAND3_X1   g12154(.A1(new_n13169_), .A2(new_n13174_), .A3(new_n13167_), .ZN(new_n13175_));
  AOI21_X1   g12155(.A1(new_n13169_), .A2(new_n13167_), .B(new_n13174_), .ZN(new_n13176_));
  INV_X1     g12156(.I(new_n13176_), .ZN(new_n13177_));
  AOI22_X1   g12157(.A1(new_n12082_), .A2(new_n12432_), .B1(new_n12351_), .B2(new_n12431_), .ZN(new_n13178_));
  NOR2_X1    g12158(.A1(new_n12434_), .A2(new_n13178_), .ZN(new_n13179_));
  NAND3_X1   g12159(.A1(new_n13177_), .A2(new_n13179_), .A3(new_n13175_), .ZN(new_n13180_));
  NAND2_X1   g12160(.A1(new_n13161_), .A2(new_n13180_), .ZN(new_n13181_));
  AND3_X2    g12161(.A1(new_n13169_), .A2(new_n13167_), .A3(new_n13174_), .Z(new_n13182_));
  OR2_X2     g12162(.A1(new_n12434_), .A2(new_n13178_), .Z(new_n13183_));
  NOR3_X1    g12163(.A1(new_n13183_), .A2(new_n13182_), .A3(new_n13176_), .ZN(new_n13184_));
  NAND3_X1   g12164(.A1(new_n13184_), .A2(new_n12438_), .A3(new_n12443_), .ZN(new_n13185_));
  NAND2_X1   g12165(.A1(new_n13181_), .A2(new_n13185_), .ZN(new_n13186_));
  NOR2_X1    g12166(.A1(new_n13161_), .A2(new_n13180_), .ZN(new_n13187_));
  AOI21_X1   g12167(.A1(new_n13028_), .A2(new_n13030_), .B(new_n13041_), .ZN(new_n13188_));
  INV_X1     g12168(.I(new_n13188_), .ZN(new_n13189_));
  NAND3_X1   g12169(.A1(new_n13072_), .A2(new_n12718_), .A3(new_n12719_), .ZN(new_n13190_));
  NOR3_X1    g12170(.A1(new_n13055_), .A2(new_n13059_), .A3(new_n13056_), .ZN(new_n13191_));
  INV_X1     g12171(.I(new_n13191_), .ZN(new_n13192_));
  NAND3_X1   g12172(.A1(new_n13189_), .A2(new_n13192_), .A3(new_n13190_), .ZN(new_n13193_));
  NOR3_X1    g12173(.A1(new_n12728_), .A2(new_n13070_), .A3(new_n12717_), .ZN(new_n13194_));
  OAI21_X1   g12174(.A1(new_n13188_), .A2(new_n13191_), .B(new_n13194_), .ZN(new_n13195_));
  AOI21_X1   g12175(.A1(new_n13193_), .A2(new_n13195_), .B(new_n13182_), .ZN(new_n13196_));
  NOR3_X1    g12176(.A1(new_n13194_), .A2(new_n13191_), .A3(new_n13188_), .ZN(new_n13197_));
  AOI21_X1   g12177(.A1(new_n13192_), .A2(new_n13189_), .B(new_n13190_), .ZN(new_n13198_));
  NOR3_X1    g12178(.A1(new_n13198_), .A2(new_n13197_), .A3(new_n13175_), .ZN(new_n13199_));
  NOR2_X1    g12179(.A1(new_n13196_), .A2(new_n13199_), .ZN(new_n13200_));
  AOI21_X1   g12180(.A1(new_n13186_), .A2(new_n13200_), .B(new_n13187_), .ZN(new_n13201_));
  INV_X1     g12181(.I(new_n13201_), .ZN(new_n13202_));
  OAI21_X1   g12182(.A1(new_n13158_), .A2(new_n13159_), .B(new_n13155_), .ZN(new_n13203_));
  AOI21_X1   g12183(.A1(new_n13202_), .A2(new_n13203_), .B(new_n13160_), .ZN(new_n13204_));
  NOR2_X1    g12184(.A1(new_n13204_), .A2(new_n13144_), .ZN(new_n13205_));
  OAI21_X1   g12185(.A1(new_n13094_), .A2(new_n13095_), .B(new_n12872_), .ZN(new_n13206_));
  NAND3_X1   g12186(.A1(new_n13088_), .A2(new_n13090_), .A3(new_n13087_), .ZN(new_n13207_));
  AOI21_X1   g12187(.A1(new_n13206_), .A2(new_n13207_), .B(new_n13086_), .ZN(new_n13208_));
  NOR3_X1    g12188(.A1(new_n13153_), .A2(new_n13096_), .A3(new_n13091_), .ZN(new_n13209_));
  OAI21_X1   g12189(.A1(new_n13208_), .A2(new_n13209_), .B(new_n13098_), .ZN(new_n13210_));
  AOI21_X1   g12190(.A1(new_n13206_), .A2(new_n13207_), .B(new_n13153_), .ZN(new_n13211_));
  NOR3_X1    g12191(.A1(new_n13086_), .A2(new_n13096_), .A3(new_n13091_), .ZN(new_n13212_));
  OAI21_X1   g12192(.A1(new_n13211_), .A2(new_n13212_), .B(new_n13102_), .ZN(new_n13213_));
  NAND2_X1   g12193(.A1(new_n13210_), .A2(new_n13213_), .ZN(new_n13214_));
  AOI21_X1   g12194(.A1(new_n13204_), .A2(new_n13144_), .B(new_n13214_), .ZN(new_n13215_));
  XNOR2_X1   g12195(.A1(new_n12502_), .A2(new_n12501_), .ZN(new_n13216_));
  AND3_X2    g12196(.A1(new_n13216_), .A2(new_n12488_), .A3(new_n12492_), .Z(new_n13217_));
  NAND2_X1   g12197(.A1(new_n13105_), .A2(new_n12758_), .ZN(new_n13218_));
  NAND2_X1   g12198(.A1(new_n13206_), .A2(new_n13207_), .ZN(new_n13219_));
  OAI21_X1   g12199(.A1(new_n13219_), .A2(new_n13098_), .B(new_n13153_), .ZN(new_n13220_));
  NAND3_X1   g12200(.A1(new_n13220_), .A2(new_n12759_), .A3(new_n13104_), .ZN(new_n13221_));
  AOI21_X1   g12201(.A1(new_n13218_), .A2(new_n13221_), .B(new_n13052_), .ZN(new_n13222_));
  AOI21_X1   g12202(.A1(new_n13220_), .A2(new_n13104_), .B(new_n12759_), .ZN(new_n13223_));
  NOR2_X1    g12203(.A1(new_n13105_), .A2(new_n12758_), .ZN(new_n13224_));
  NOR3_X1    g12204(.A1(new_n13224_), .A2(new_n13223_), .A3(new_n13051_), .ZN(new_n13225_));
  NOR3_X1    g12205(.A1(new_n13225_), .A2(new_n13222_), .A3(new_n13217_), .ZN(new_n13226_));
  NOR3_X1    g12206(.A1(new_n13226_), .A2(new_n13205_), .A3(new_n13215_), .ZN(new_n13227_));
  XOR2_X1    g12207(.A1(new_n12758_), .A2(new_n13052_), .Z(new_n13228_));
  NAND3_X1   g12208(.A1(new_n13217_), .A2(new_n13228_), .A3(new_n13106_), .ZN(new_n13229_));
  OAI21_X1   g12209(.A1(new_n13227_), .A2(new_n13229_), .B(new_n13111_), .ZN(new_n13230_));
  NAND2_X1   g12210(.A1(new_n13230_), .A2(new_n13110_), .ZN(new_n13231_));
  INV_X1     g12211(.I(\A[718] ), .ZN(new_n13232_));
  NOR2_X1    g12212(.A1(\A[719] ), .A2(\A[720] ), .ZN(new_n13233_));
  NAND2_X1   g12213(.A1(\A[719] ), .A2(\A[720] ), .ZN(new_n13234_));
  AOI21_X1   g12214(.A1(new_n13232_), .A2(new_n13234_), .B(new_n13233_), .ZN(new_n13235_));
  INV_X1     g12215(.I(\A[715] ), .ZN(new_n13236_));
  NOR2_X1    g12216(.A1(\A[716] ), .A2(\A[717] ), .ZN(new_n13237_));
  NAND2_X1   g12217(.A1(\A[716] ), .A2(\A[717] ), .ZN(new_n13238_));
  AOI21_X1   g12218(.A1(new_n13236_), .A2(new_n13238_), .B(new_n13237_), .ZN(new_n13239_));
  INV_X1     g12219(.I(\A[716] ), .ZN(new_n13240_));
  NAND2_X1   g12220(.A1(new_n13240_), .A2(\A[717] ), .ZN(new_n13241_));
  INV_X1     g12221(.I(\A[717] ), .ZN(new_n13242_));
  NAND2_X1   g12222(.A1(new_n13242_), .A2(\A[716] ), .ZN(new_n13243_));
  AOI21_X1   g12223(.A1(new_n13241_), .A2(new_n13243_), .B(new_n13236_), .ZN(new_n13244_));
  INV_X1     g12224(.I(new_n13237_), .ZN(new_n13245_));
  AOI21_X1   g12225(.A1(new_n13245_), .A2(new_n13238_), .B(\A[715] ), .ZN(new_n13246_));
  INV_X1     g12226(.I(\A[719] ), .ZN(new_n13247_));
  NAND2_X1   g12227(.A1(new_n13247_), .A2(\A[720] ), .ZN(new_n13248_));
  INV_X1     g12228(.I(\A[720] ), .ZN(new_n13249_));
  NAND2_X1   g12229(.A1(new_n13249_), .A2(\A[719] ), .ZN(new_n13250_));
  AOI21_X1   g12230(.A1(new_n13248_), .A2(new_n13250_), .B(new_n13232_), .ZN(new_n13251_));
  INV_X1     g12231(.I(new_n13233_), .ZN(new_n13252_));
  AOI21_X1   g12232(.A1(new_n13252_), .A2(new_n13234_), .B(\A[718] ), .ZN(new_n13253_));
  NOR4_X1    g12233(.A1(new_n13244_), .A2(new_n13246_), .A3(new_n13253_), .A4(new_n13251_), .ZN(new_n13254_));
  XNOR2_X1   g12234(.A1(new_n13254_), .A2(new_n13239_), .ZN(new_n13255_));
  XOR2_X1    g12235(.A1(new_n13255_), .A2(new_n13235_), .Z(new_n13256_));
  INV_X1     g12236(.I(\A[724] ), .ZN(new_n13257_));
  NOR2_X1    g12237(.A1(\A[725] ), .A2(\A[726] ), .ZN(new_n13258_));
  NAND2_X1   g12238(.A1(\A[725] ), .A2(\A[726] ), .ZN(new_n13259_));
  AOI21_X1   g12239(.A1(new_n13257_), .A2(new_n13259_), .B(new_n13258_), .ZN(new_n13260_));
  INV_X1     g12240(.I(\A[721] ), .ZN(new_n13261_));
  NOR2_X1    g12241(.A1(\A[722] ), .A2(\A[723] ), .ZN(new_n13262_));
  NAND2_X1   g12242(.A1(\A[722] ), .A2(\A[723] ), .ZN(new_n13263_));
  AOI21_X1   g12243(.A1(new_n13261_), .A2(new_n13263_), .B(new_n13262_), .ZN(new_n13264_));
  INV_X1     g12244(.I(new_n13264_), .ZN(new_n13265_));
  INV_X1     g12245(.I(\A[723] ), .ZN(new_n13266_));
  NOR2_X1    g12246(.A1(new_n13266_), .A2(\A[722] ), .ZN(new_n13267_));
  INV_X1     g12247(.I(\A[722] ), .ZN(new_n13268_));
  NOR2_X1    g12248(.A1(new_n13268_), .A2(\A[723] ), .ZN(new_n13269_));
  OAI21_X1   g12249(.A1(new_n13267_), .A2(new_n13269_), .B(\A[721] ), .ZN(new_n13270_));
  INV_X1     g12250(.I(new_n13263_), .ZN(new_n13271_));
  OAI21_X1   g12251(.A1(new_n13271_), .A2(new_n13262_), .B(new_n13261_), .ZN(new_n13272_));
  NAND2_X1   g12252(.A1(new_n13270_), .A2(new_n13272_), .ZN(new_n13273_));
  INV_X1     g12253(.I(\A[726] ), .ZN(new_n13274_));
  NOR2_X1    g12254(.A1(new_n13274_), .A2(\A[725] ), .ZN(new_n13275_));
  INV_X1     g12255(.I(\A[725] ), .ZN(new_n13276_));
  NOR2_X1    g12256(.A1(new_n13276_), .A2(\A[726] ), .ZN(new_n13277_));
  OAI21_X1   g12257(.A1(new_n13275_), .A2(new_n13277_), .B(\A[724] ), .ZN(new_n13278_));
  INV_X1     g12258(.I(new_n13259_), .ZN(new_n13279_));
  OAI21_X1   g12259(.A1(new_n13279_), .A2(new_n13258_), .B(new_n13257_), .ZN(new_n13280_));
  NAND2_X1   g12260(.A1(new_n13278_), .A2(new_n13280_), .ZN(new_n13281_));
  NOR2_X1    g12261(.A1(new_n13273_), .A2(new_n13281_), .ZN(new_n13282_));
  NOR2_X1    g12262(.A1(new_n13282_), .A2(new_n13265_), .ZN(new_n13283_));
  NAND2_X1   g12263(.A1(new_n13268_), .A2(\A[723] ), .ZN(new_n13284_));
  NAND2_X1   g12264(.A1(new_n13266_), .A2(\A[722] ), .ZN(new_n13285_));
  AOI21_X1   g12265(.A1(new_n13284_), .A2(new_n13285_), .B(new_n13261_), .ZN(new_n13286_));
  INV_X1     g12266(.I(new_n13262_), .ZN(new_n13287_));
  AOI21_X1   g12267(.A1(new_n13287_), .A2(new_n13263_), .B(\A[721] ), .ZN(new_n13288_));
  NOR2_X1    g12268(.A1(new_n13288_), .A2(new_n13286_), .ZN(new_n13289_));
  NAND2_X1   g12269(.A1(new_n13276_), .A2(\A[726] ), .ZN(new_n13290_));
  NAND2_X1   g12270(.A1(new_n13274_), .A2(\A[725] ), .ZN(new_n13291_));
  AOI21_X1   g12271(.A1(new_n13290_), .A2(new_n13291_), .B(new_n13257_), .ZN(new_n13292_));
  INV_X1     g12272(.I(new_n13258_), .ZN(new_n13293_));
  AOI21_X1   g12273(.A1(new_n13293_), .A2(new_n13259_), .B(\A[724] ), .ZN(new_n13294_));
  NOR2_X1    g12274(.A1(new_n13294_), .A2(new_n13292_), .ZN(new_n13295_));
  NAND2_X1   g12275(.A1(new_n13289_), .A2(new_n13295_), .ZN(new_n13296_));
  NOR2_X1    g12276(.A1(new_n13296_), .A2(new_n13264_), .ZN(new_n13297_));
  OAI21_X1   g12277(.A1(new_n13283_), .A2(new_n13297_), .B(new_n13260_), .ZN(new_n13298_));
  INV_X1     g12278(.I(new_n13260_), .ZN(new_n13299_));
  NAND2_X1   g12279(.A1(new_n13296_), .A2(new_n13264_), .ZN(new_n13300_));
  NAND2_X1   g12280(.A1(new_n13282_), .A2(new_n13265_), .ZN(new_n13301_));
  NAND3_X1   g12281(.A1(new_n13301_), .A2(new_n13300_), .A3(new_n13299_), .ZN(new_n13302_));
  NAND2_X1   g12282(.A1(new_n13298_), .A2(new_n13302_), .ZN(new_n13303_));
  NOR2_X1    g12283(.A1(new_n13246_), .A2(new_n13244_), .ZN(new_n13304_));
  NOR2_X1    g12284(.A1(new_n13253_), .A2(new_n13251_), .ZN(new_n13305_));
  NAND2_X1   g12285(.A1(new_n13304_), .A2(new_n13305_), .ZN(new_n13306_));
  NAND2_X1   g12286(.A1(new_n13235_), .A2(new_n13239_), .ZN(new_n13307_));
  NOR2_X1    g12287(.A1(new_n13289_), .A2(new_n13295_), .ZN(new_n13308_));
  NOR4_X1    g12288(.A1(new_n13282_), .A2(new_n13308_), .A3(new_n13306_), .A4(new_n13307_), .ZN(new_n13309_));
  NOR2_X1    g12289(.A1(new_n13304_), .A2(new_n13305_), .ZN(new_n13310_));
  NOR2_X1    g12290(.A1(new_n13310_), .A2(new_n13254_), .ZN(new_n13311_));
  NAND2_X1   g12291(.A1(new_n13260_), .A2(new_n13264_), .ZN(new_n13312_));
  NOR3_X1    g12292(.A1(new_n13273_), .A2(new_n13281_), .A3(new_n13312_), .ZN(new_n13313_));
  NAND3_X1   g12293(.A1(new_n13309_), .A2(new_n13311_), .A3(new_n13313_), .ZN(new_n13314_));
  INV_X1     g12294(.I(new_n13314_), .ZN(new_n13315_));
  NAND2_X1   g12295(.A1(new_n13315_), .A2(new_n13303_), .ZN(new_n13316_));
  AOI21_X1   g12296(.A1(new_n13301_), .A2(new_n13300_), .B(new_n13299_), .ZN(new_n13317_));
  NOR3_X1    g12297(.A1(new_n13283_), .A2(new_n13297_), .A3(new_n13260_), .ZN(new_n13318_));
  NOR2_X1    g12298(.A1(new_n13317_), .A2(new_n13318_), .ZN(new_n13319_));
  NAND2_X1   g12299(.A1(new_n13319_), .A2(new_n13314_), .ZN(new_n13320_));
  AOI21_X1   g12300(.A1(new_n13316_), .A2(new_n13320_), .B(new_n13256_), .ZN(new_n13321_));
  NAND2_X1   g12301(.A1(new_n13309_), .A2(new_n13311_), .ZN(new_n13322_));
  INV_X1     g12302(.I(new_n13322_), .ZN(new_n13323_));
  NOR2_X1    g12303(.A1(new_n13308_), .A2(new_n13312_), .ZN(new_n13324_));
  AOI21_X1   g12304(.A1(new_n13319_), .A2(new_n13323_), .B(new_n13324_), .ZN(new_n13325_));
  NOR2_X1    g12305(.A1(new_n13303_), .A2(new_n13314_), .ZN(new_n13326_));
  NOR3_X1    g12306(.A1(new_n13325_), .A2(new_n13256_), .A3(new_n13326_), .ZN(new_n13327_));
  NOR2_X1    g12307(.A1(new_n13321_), .A2(new_n13327_), .ZN(new_n13328_));
  XNOR2_X1   g12308(.A1(new_n13255_), .A2(new_n13235_), .ZN(new_n13329_));
  NOR2_X1    g12309(.A1(new_n13319_), .A2(new_n13314_), .ZN(new_n13330_));
  NOR2_X1    g12310(.A1(new_n13315_), .A2(new_n13303_), .ZN(new_n13331_));
  OAI21_X1   g12311(.A1(new_n13331_), .A2(new_n13330_), .B(new_n13329_), .ZN(new_n13332_));
  OAI22_X1   g12312(.A1(new_n13303_), .A2(new_n13322_), .B1(new_n13308_), .B2(new_n13312_), .ZN(new_n13333_));
  NAND2_X1   g12313(.A1(new_n13315_), .A2(new_n13319_), .ZN(new_n13334_));
  NAND3_X1   g12314(.A1(new_n13329_), .A2(new_n13333_), .A3(new_n13334_), .ZN(new_n13335_));
  NOR2_X1    g12315(.A1(new_n13308_), .A2(new_n13282_), .ZN(new_n13336_));
  NAND2_X1   g12316(.A1(new_n13336_), .A2(new_n13313_), .ZN(new_n13337_));
  NOR2_X1    g12317(.A1(new_n13306_), .A2(new_n13307_), .ZN(new_n13338_));
  NAND2_X1   g12318(.A1(new_n13311_), .A2(new_n13338_), .ZN(new_n13339_));
  XOR2_X1    g12319(.A1(new_n13339_), .A2(new_n13337_), .Z(new_n13340_));
  NOR2_X1    g12320(.A1(\A[713] ), .A2(\A[714] ), .ZN(new_n13341_));
  INV_X1     g12321(.I(new_n13341_), .ZN(new_n13342_));
  INV_X1     g12322(.I(\A[713] ), .ZN(new_n13343_));
  INV_X1     g12323(.I(\A[714] ), .ZN(new_n13344_));
  NOR2_X1    g12324(.A1(new_n13343_), .A2(new_n13344_), .ZN(new_n13345_));
  OAI21_X1   g12325(.A1(\A[712] ), .A2(new_n13345_), .B(new_n13342_), .ZN(new_n13346_));
  NOR2_X1    g12326(.A1(\A[710] ), .A2(\A[711] ), .ZN(new_n13347_));
  INV_X1     g12327(.I(new_n13347_), .ZN(new_n13348_));
  INV_X1     g12328(.I(\A[710] ), .ZN(new_n13349_));
  INV_X1     g12329(.I(\A[711] ), .ZN(new_n13350_));
  NOR2_X1    g12330(.A1(new_n13349_), .A2(new_n13350_), .ZN(new_n13351_));
  OAI21_X1   g12331(.A1(\A[709] ), .A2(new_n13351_), .B(new_n13348_), .ZN(new_n13352_));
  NOR2_X1    g12332(.A1(new_n13346_), .A2(new_n13352_), .ZN(new_n13353_));
  INV_X1     g12333(.I(new_n13353_), .ZN(new_n13354_));
  NOR2_X1    g12334(.A1(new_n13350_), .A2(\A[710] ), .ZN(new_n13355_));
  NOR2_X1    g12335(.A1(new_n13349_), .A2(\A[711] ), .ZN(new_n13356_));
  OAI21_X1   g12336(.A1(new_n13355_), .A2(new_n13356_), .B(\A[709] ), .ZN(new_n13357_));
  INV_X1     g12337(.I(\A[709] ), .ZN(new_n13358_));
  OAI21_X1   g12338(.A1(new_n13351_), .A2(new_n13347_), .B(new_n13358_), .ZN(new_n13359_));
  NOR2_X1    g12339(.A1(new_n13344_), .A2(\A[713] ), .ZN(new_n13360_));
  NOR2_X1    g12340(.A1(new_n13343_), .A2(\A[714] ), .ZN(new_n13361_));
  OAI21_X1   g12341(.A1(new_n13360_), .A2(new_n13361_), .B(\A[712] ), .ZN(new_n13362_));
  INV_X1     g12342(.I(\A[712] ), .ZN(new_n13363_));
  OAI21_X1   g12343(.A1(new_n13345_), .A2(new_n13341_), .B(new_n13363_), .ZN(new_n13364_));
  NAND4_X1   g12344(.A1(new_n13357_), .A2(new_n13359_), .A3(new_n13364_), .A4(new_n13362_), .ZN(new_n13365_));
  NOR2_X1    g12345(.A1(new_n13354_), .A2(new_n13365_), .ZN(new_n13366_));
  NAND2_X1   g12346(.A1(new_n13359_), .A2(new_n13357_), .ZN(new_n13367_));
  NAND2_X1   g12347(.A1(new_n13364_), .A2(new_n13362_), .ZN(new_n13368_));
  NAND2_X1   g12348(.A1(new_n13367_), .A2(new_n13368_), .ZN(new_n13369_));
  AND2_X2    g12349(.A1(new_n13369_), .A2(new_n13365_), .Z(new_n13370_));
  INV_X1     g12350(.I(\A[703] ), .ZN(new_n13371_));
  INV_X1     g12351(.I(\A[704] ), .ZN(new_n13372_));
  NAND2_X1   g12352(.A1(new_n13372_), .A2(\A[705] ), .ZN(new_n13373_));
  INV_X1     g12353(.I(\A[705] ), .ZN(new_n13374_));
  NAND2_X1   g12354(.A1(new_n13374_), .A2(\A[704] ), .ZN(new_n13375_));
  AOI21_X1   g12355(.A1(new_n13373_), .A2(new_n13375_), .B(new_n13371_), .ZN(new_n13376_));
  NOR2_X1    g12356(.A1(\A[704] ), .A2(\A[705] ), .ZN(new_n13377_));
  INV_X1     g12357(.I(new_n13377_), .ZN(new_n13378_));
  NAND2_X1   g12358(.A1(\A[704] ), .A2(\A[705] ), .ZN(new_n13379_));
  AOI21_X1   g12359(.A1(new_n13378_), .A2(new_n13379_), .B(\A[703] ), .ZN(new_n13380_));
  NOR2_X1    g12360(.A1(new_n13380_), .A2(new_n13376_), .ZN(new_n13381_));
  INV_X1     g12361(.I(\A[706] ), .ZN(new_n13382_));
  INV_X1     g12362(.I(\A[707] ), .ZN(new_n13383_));
  NAND2_X1   g12363(.A1(new_n13383_), .A2(\A[708] ), .ZN(new_n13384_));
  INV_X1     g12364(.I(\A[708] ), .ZN(new_n13385_));
  NAND2_X1   g12365(.A1(new_n13385_), .A2(\A[707] ), .ZN(new_n13386_));
  AOI21_X1   g12366(.A1(new_n13384_), .A2(new_n13386_), .B(new_n13382_), .ZN(new_n13387_));
  NOR2_X1    g12367(.A1(\A[707] ), .A2(\A[708] ), .ZN(new_n13388_));
  INV_X1     g12368(.I(new_n13388_), .ZN(new_n13389_));
  NAND2_X1   g12369(.A1(\A[707] ), .A2(\A[708] ), .ZN(new_n13390_));
  AOI21_X1   g12370(.A1(new_n13389_), .A2(new_n13390_), .B(\A[706] ), .ZN(new_n13391_));
  NOR2_X1    g12371(.A1(new_n13391_), .A2(new_n13387_), .ZN(new_n13392_));
  AOI21_X1   g12372(.A1(new_n13382_), .A2(new_n13390_), .B(new_n13388_), .ZN(new_n13393_));
  INV_X1     g12373(.I(new_n13393_), .ZN(new_n13394_));
  AOI21_X1   g12374(.A1(new_n13371_), .A2(new_n13379_), .B(new_n13377_), .ZN(new_n13395_));
  INV_X1     g12375(.I(new_n13395_), .ZN(new_n13396_));
  NOR2_X1    g12376(.A1(new_n13394_), .A2(new_n13396_), .ZN(new_n13397_));
  NAND2_X1   g12377(.A1(new_n13370_), .A2(new_n13366_), .ZN(new_n13398_));
  INV_X1     g12378(.I(new_n13398_), .ZN(new_n13399_));
  NOR2_X1    g12379(.A1(new_n13340_), .A2(new_n13399_), .ZN(new_n13400_));
  AOI21_X1   g12380(.A1(new_n13332_), .A2(new_n13335_), .B(new_n13400_), .ZN(new_n13401_));
  XNOR2_X1   g12381(.A1(new_n13339_), .A2(new_n13337_), .ZN(new_n13402_));
  NAND2_X1   g12382(.A1(new_n13402_), .A2(new_n13398_), .ZN(new_n13403_));
  NOR3_X1    g12383(.A1(new_n13321_), .A2(new_n13327_), .A3(new_n13403_), .ZN(new_n13404_));
  NAND2_X1   g12384(.A1(new_n13381_), .A2(new_n13392_), .ZN(new_n13405_));
  INV_X1     g12385(.I(new_n13397_), .ZN(new_n13406_));
  NOR2_X1    g12386(.A1(new_n13405_), .A2(new_n13406_), .ZN(new_n13407_));
  INV_X1     g12387(.I(new_n13346_), .ZN(new_n13408_));
  INV_X1     g12388(.I(new_n13352_), .ZN(new_n13409_));
  NAND2_X1   g12389(.A1(new_n13365_), .A2(new_n13409_), .ZN(new_n13410_));
  INV_X1     g12390(.I(new_n13410_), .ZN(new_n13411_));
  NOR2_X1    g12391(.A1(new_n13365_), .A2(new_n13409_), .ZN(new_n13412_));
  OAI21_X1   g12392(.A1(new_n13411_), .A2(new_n13412_), .B(new_n13408_), .ZN(new_n13413_));
  INV_X1     g12393(.I(new_n13412_), .ZN(new_n13414_));
  NAND3_X1   g12394(.A1(new_n13414_), .A2(new_n13410_), .A3(new_n13346_), .ZN(new_n13415_));
  INV_X1     g12395(.I(new_n13365_), .ZN(new_n13416_));
  NAND2_X1   g12396(.A1(new_n13416_), .A2(new_n13353_), .ZN(new_n13417_));
  NOR2_X1    g12397(.A1(new_n13374_), .A2(\A[704] ), .ZN(new_n13418_));
  NOR2_X1    g12398(.A1(new_n13372_), .A2(\A[705] ), .ZN(new_n13419_));
  OAI21_X1   g12399(.A1(new_n13418_), .A2(new_n13419_), .B(\A[703] ), .ZN(new_n13420_));
  INV_X1     g12400(.I(new_n13379_), .ZN(new_n13421_));
  OAI21_X1   g12401(.A1(new_n13421_), .A2(new_n13377_), .B(new_n13371_), .ZN(new_n13422_));
  NAND2_X1   g12402(.A1(new_n13420_), .A2(new_n13422_), .ZN(new_n13423_));
  NOR2_X1    g12403(.A1(new_n13385_), .A2(\A[707] ), .ZN(new_n13424_));
  NOR2_X1    g12404(.A1(new_n13383_), .A2(\A[708] ), .ZN(new_n13425_));
  OAI21_X1   g12405(.A1(new_n13424_), .A2(new_n13425_), .B(\A[706] ), .ZN(new_n13426_));
  INV_X1     g12406(.I(new_n13390_), .ZN(new_n13427_));
  OAI21_X1   g12407(.A1(new_n13427_), .A2(new_n13388_), .B(new_n13382_), .ZN(new_n13428_));
  NAND2_X1   g12408(.A1(new_n13426_), .A2(new_n13428_), .ZN(new_n13429_));
  NOR2_X1    g12409(.A1(new_n13423_), .A2(new_n13429_), .ZN(new_n13430_));
  NOR2_X1    g12410(.A1(new_n13381_), .A2(new_n13392_), .ZN(new_n13431_));
  NOR3_X1    g12411(.A1(new_n13417_), .A2(new_n13430_), .A3(new_n13431_), .ZN(new_n13432_));
  NAND4_X1   g12412(.A1(new_n13413_), .A2(new_n13432_), .A3(new_n13415_), .A4(new_n13370_), .ZN(new_n13433_));
  XOR2_X1    g12413(.A1(new_n13367_), .A2(new_n13368_), .Z(new_n13434_));
  NAND2_X1   g12414(.A1(new_n13434_), .A2(new_n13353_), .ZN(new_n13435_));
  NAND3_X1   g12415(.A1(new_n13433_), .A2(new_n13407_), .A3(new_n13435_), .ZN(new_n13436_));
  NAND2_X1   g12416(.A1(new_n13405_), .A2(new_n13395_), .ZN(new_n13437_));
  NAND2_X1   g12417(.A1(new_n13430_), .A2(new_n13396_), .ZN(new_n13438_));
  AOI21_X1   g12418(.A1(new_n13438_), .A2(new_n13437_), .B(new_n13394_), .ZN(new_n13439_));
  NOR2_X1    g12419(.A1(new_n13430_), .A2(new_n13396_), .ZN(new_n13440_));
  NOR2_X1    g12420(.A1(new_n13405_), .A2(new_n13395_), .ZN(new_n13441_));
  NOR3_X1    g12421(.A1(new_n13440_), .A2(new_n13441_), .A3(new_n13393_), .ZN(new_n13442_));
  NOR2_X1    g12422(.A1(new_n13439_), .A2(new_n13442_), .ZN(new_n13443_));
  NOR2_X1    g12423(.A1(new_n13436_), .A2(new_n13443_), .ZN(new_n13444_));
  OR2_X2     g12424(.A1(new_n13439_), .A2(new_n13442_), .Z(new_n13445_));
  NOR2_X1    g12425(.A1(new_n13431_), .A2(new_n13430_), .ZN(new_n13446_));
  NAND4_X1   g12426(.A1(new_n13370_), .A2(new_n13366_), .A3(new_n13446_), .A4(new_n13407_), .ZN(new_n13447_));
  NAND2_X1   g12427(.A1(new_n13445_), .A2(new_n13447_), .ZN(new_n13448_));
  NAND3_X1   g12428(.A1(new_n13435_), .A2(new_n13413_), .A3(new_n13415_), .ZN(new_n13449_));
  NOR3_X1    g12429(.A1(new_n13447_), .A2(new_n13439_), .A3(new_n13442_), .ZN(new_n13450_));
  XOR2_X1    g12430(.A1(new_n13450_), .A2(new_n13449_), .Z(new_n13451_));
  AOI21_X1   g12431(.A1(new_n13451_), .A2(new_n13448_), .B(new_n13444_), .ZN(new_n13452_));
  OAI22_X1   g12432(.A1(new_n13452_), .A2(new_n13328_), .B1(new_n13401_), .B2(new_n13404_), .ZN(new_n13453_));
  NOR2_X1    g12433(.A1(new_n13329_), .A2(new_n13326_), .ZN(new_n13454_));
  NOR2_X1    g12434(.A1(new_n13260_), .A2(new_n13264_), .ZN(new_n13455_));
  OAI21_X1   g12435(.A1(new_n13296_), .A2(new_n13455_), .B(new_n13312_), .ZN(new_n13456_));
  NOR2_X1    g12436(.A1(new_n13235_), .A2(new_n13239_), .ZN(new_n13457_));
  OAI21_X1   g12437(.A1(new_n13306_), .A2(new_n13457_), .B(new_n13307_), .ZN(new_n13458_));
  XNOR2_X1   g12438(.A1(new_n13456_), .A2(new_n13458_), .ZN(new_n13459_));
  INV_X1     g12439(.I(new_n13459_), .ZN(new_n13460_));
  NOR3_X1    g12440(.A1(new_n13454_), .A2(new_n13325_), .A3(new_n13460_), .ZN(new_n13461_));
  AND3_X2    g12441(.A1(new_n13435_), .A2(new_n13413_), .A3(new_n13415_), .Z(new_n13462_));
  OAI21_X1   g12442(.A1(new_n13462_), .A2(new_n13447_), .B(new_n13445_), .ZN(new_n13463_));
  NOR2_X1    g12443(.A1(new_n13408_), .A2(new_n13409_), .ZN(new_n13464_));
  OAI21_X1   g12444(.A1(new_n13365_), .A2(new_n13464_), .B(new_n13354_), .ZN(new_n13465_));
  NOR2_X1    g12445(.A1(new_n13393_), .A2(new_n13395_), .ZN(new_n13466_));
  OAI21_X1   g12446(.A1(new_n13405_), .A2(new_n13466_), .B(new_n13406_), .ZN(new_n13467_));
  XNOR2_X1   g12447(.A1(new_n13467_), .A2(new_n13465_), .ZN(new_n13468_));
  NAND3_X1   g12448(.A1(new_n13463_), .A2(new_n13436_), .A3(new_n13468_), .ZN(new_n13469_));
  XOR2_X1    g12449(.A1(new_n13461_), .A2(new_n13469_), .Z(new_n13470_));
  NOR2_X1    g12450(.A1(new_n13470_), .A2(new_n13453_), .ZN(new_n13471_));
  NAND2_X1   g12451(.A1(new_n13332_), .A2(new_n13335_), .ZN(new_n13472_));
  OAI21_X1   g12452(.A1(new_n13321_), .A2(new_n13327_), .B(new_n13403_), .ZN(new_n13473_));
  NAND3_X1   g12453(.A1(new_n13332_), .A2(new_n13335_), .A3(new_n13400_), .ZN(new_n13474_));
  AND4_X2    g12454(.A1(new_n13370_), .A2(new_n13413_), .A3(new_n13432_), .A4(new_n13415_), .Z(new_n13475_));
  NAND2_X1   g12455(.A1(new_n13435_), .A2(new_n13407_), .ZN(new_n13476_));
  NOR2_X1    g12456(.A1(new_n13475_), .A2(new_n13476_), .ZN(new_n13477_));
  NAND2_X1   g12457(.A1(new_n13477_), .A2(new_n13445_), .ZN(new_n13478_));
  NOR2_X1    g12458(.A1(new_n13462_), .A2(new_n13450_), .ZN(new_n13479_));
  NOR3_X1    g12459(.A1(new_n13445_), .A2(new_n13447_), .A3(new_n13449_), .ZN(new_n13480_));
  OAI21_X1   g12460(.A1(new_n13479_), .A2(new_n13480_), .B(new_n13448_), .ZN(new_n13481_));
  NAND2_X1   g12461(.A1(new_n13481_), .A2(new_n13478_), .ZN(new_n13482_));
  AOI22_X1   g12462(.A1(new_n13482_), .A2(new_n13472_), .B1(new_n13474_), .B2(new_n13473_), .ZN(new_n13483_));
  INV_X1     g12463(.I(new_n13447_), .ZN(new_n13484_));
  AOI21_X1   g12464(.A1(new_n13484_), .A2(new_n13449_), .B(new_n13443_), .ZN(new_n13485_));
  INV_X1     g12465(.I(new_n13468_), .ZN(new_n13486_));
  NOR3_X1    g12466(.A1(new_n13477_), .A2(new_n13485_), .A3(new_n13486_), .ZN(new_n13487_));
  NOR2_X1    g12467(.A1(new_n13461_), .A2(new_n13487_), .ZN(new_n13488_));
  NAND2_X1   g12468(.A1(new_n13334_), .A2(new_n13256_), .ZN(new_n13489_));
  NAND3_X1   g12469(.A1(new_n13489_), .A2(new_n13333_), .A3(new_n13459_), .ZN(new_n13490_));
  NOR2_X1    g12470(.A1(new_n13490_), .A2(new_n13469_), .ZN(new_n13491_));
  NOR2_X1    g12471(.A1(new_n13488_), .A2(new_n13491_), .ZN(new_n13492_));
  NOR2_X1    g12472(.A1(new_n13483_), .A2(new_n13492_), .ZN(new_n13493_));
  NOR2_X1    g12473(.A1(new_n13471_), .A2(new_n13493_), .ZN(new_n13494_));
  INV_X1     g12474(.I(\A[742] ), .ZN(new_n13495_));
  NOR2_X1    g12475(.A1(\A[743] ), .A2(\A[744] ), .ZN(new_n13496_));
  NAND2_X1   g12476(.A1(\A[743] ), .A2(\A[744] ), .ZN(new_n13497_));
  AOI21_X1   g12477(.A1(new_n13495_), .A2(new_n13497_), .B(new_n13496_), .ZN(new_n13498_));
  INV_X1     g12478(.I(\A[739] ), .ZN(new_n13499_));
  NOR2_X1    g12479(.A1(\A[740] ), .A2(\A[741] ), .ZN(new_n13500_));
  NAND2_X1   g12480(.A1(\A[740] ), .A2(\A[741] ), .ZN(new_n13501_));
  AOI21_X1   g12481(.A1(new_n13499_), .A2(new_n13501_), .B(new_n13500_), .ZN(new_n13502_));
  INV_X1     g12482(.I(new_n13502_), .ZN(new_n13503_));
  INV_X1     g12483(.I(\A[740] ), .ZN(new_n13504_));
  NAND2_X1   g12484(.A1(new_n13504_), .A2(\A[741] ), .ZN(new_n13505_));
  INV_X1     g12485(.I(\A[741] ), .ZN(new_n13506_));
  NAND2_X1   g12486(.A1(new_n13506_), .A2(\A[740] ), .ZN(new_n13507_));
  AOI21_X1   g12487(.A1(new_n13505_), .A2(new_n13507_), .B(new_n13499_), .ZN(new_n13508_));
  INV_X1     g12488(.I(new_n13500_), .ZN(new_n13509_));
  AOI21_X1   g12489(.A1(new_n13509_), .A2(new_n13501_), .B(\A[739] ), .ZN(new_n13510_));
  INV_X1     g12490(.I(\A[743] ), .ZN(new_n13511_));
  NAND2_X1   g12491(.A1(new_n13511_), .A2(\A[744] ), .ZN(new_n13512_));
  INV_X1     g12492(.I(\A[744] ), .ZN(new_n13513_));
  NAND2_X1   g12493(.A1(new_n13513_), .A2(\A[743] ), .ZN(new_n13514_));
  AOI21_X1   g12494(.A1(new_n13512_), .A2(new_n13514_), .B(new_n13495_), .ZN(new_n13515_));
  INV_X1     g12495(.I(new_n13496_), .ZN(new_n13516_));
  AOI21_X1   g12496(.A1(new_n13516_), .A2(new_n13497_), .B(\A[742] ), .ZN(new_n13517_));
  NOR4_X1    g12497(.A1(new_n13508_), .A2(new_n13510_), .A3(new_n13517_), .A4(new_n13515_), .ZN(new_n13518_));
  NOR2_X1    g12498(.A1(new_n13518_), .A2(new_n13503_), .ZN(new_n13519_));
  NAND2_X1   g12499(.A1(new_n13518_), .A2(new_n13503_), .ZN(new_n13520_));
  INV_X1     g12500(.I(new_n13520_), .ZN(new_n13521_));
  OAI21_X1   g12501(.A1(new_n13521_), .A2(new_n13519_), .B(new_n13498_), .ZN(new_n13522_));
  INV_X1     g12502(.I(new_n13498_), .ZN(new_n13523_));
  INV_X1     g12503(.I(new_n13519_), .ZN(new_n13524_));
  NAND3_X1   g12504(.A1(new_n13524_), .A2(new_n13523_), .A3(new_n13520_), .ZN(new_n13525_));
  NAND2_X1   g12505(.A1(new_n13522_), .A2(new_n13525_), .ZN(new_n13526_));
  INV_X1     g12506(.I(\A[748] ), .ZN(new_n13527_));
  NOR2_X1    g12507(.A1(\A[749] ), .A2(\A[750] ), .ZN(new_n13528_));
  NAND2_X1   g12508(.A1(\A[749] ), .A2(\A[750] ), .ZN(new_n13529_));
  AOI21_X1   g12509(.A1(new_n13527_), .A2(new_n13529_), .B(new_n13528_), .ZN(new_n13530_));
  INV_X1     g12510(.I(\A[745] ), .ZN(new_n13531_));
  NOR2_X1    g12511(.A1(\A[746] ), .A2(\A[747] ), .ZN(new_n13532_));
  NAND2_X1   g12512(.A1(\A[746] ), .A2(\A[747] ), .ZN(new_n13533_));
  AOI21_X1   g12513(.A1(new_n13531_), .A2(new_n13533_), .B(new_n13532_), .ZN(new_n13534_));
  INV_X1     g12514(.I(new_n13534_), .ZN(new_n13535_));
  INV_X1     g12515(.I(\A[747] ), .ZN(new_n13536_));
  NOR2_X1    g12516(.A1(new_n13536_), .A2(\A[746] ), .ZN(new_n13537_));
  INV_X1     g12517(.I(\A[746] ), .ZN(new_n13538_));
  NOR2_X1    g12518(.A1(new_n13538_), .A2(\A[747] ), .ZN(new_n13539_));
  OAI21_X1   g12519(.A1(new_n13537_), .A2(new_n13539_), .B(\A[745] ), .ZN(new_n13540_));
  INV_X1     g12520(.I(new_n13533_), .ZN(new_n13541_));
  OAI21_X1   g12521(.A1(new_n13541_), .A2(new_n13532_), .B(new_n13531_), .ZN(new_n13542_));
  NAND2_X1   g12522(.A1(new_n13540_), .A2(new_n13542_), .ZN(new_n13543_));
  INV_X1     g12523(.I(\A[750] ), .ZN(new_n13544_));
  NOR2_X1    g12524(.A1(new_n13544_), .A2(\A[749] ), .ZN(new_n13545_));
  INV_X1     g12525(.I(\A[749] ), .ZN(new_n13546_));
  NOR2_X1    g12526(.A1(new_n13546_), .A2(\A[750] ), .ZN(new_n13547_));
  OAI21_X1   g12527(.A1(new_n13545_), .A2(new_n13547_), .B(\A[748] ), .ZN(new_n13548_));
  INV_X1     g12528(.I(new_n13529_), .ZN(new_n13549_));
  OAI21_X1   g12529(.A1(new_n13549_), .A2(new_n13528_), .B(new_n13527_), .ZN(new_n13550_));
  NAND2_X1   g12530(.A1(new_n13548_), .A2(new_n13550_), .ZN(new_n13551_));
  NOR2_X1    g12531(.A1(new_n13543_), .A2(new_n13551_), .ZN(new_n13552_));
  NOR2_X1    g12532(.A1(new_n13552_), .A2(new_n13535_), .ZN(new_n13553_));
  NAND2_X1   g12533(.A1(new_n13538_), .A2(\A[747] ), .ZN(new_n13554_));
  NAND2_X1   g12534(.A1(new_n13536_), .A2(\A[746] ), .ZN(new_n13555_));
  AOI21_X1   g12535(.A1(new_n13554_), .A2(new_n13555_), .B(new_n13531_), .ZN(new_n13556_));
  INV_X1     g12536(.I(new_n13532_), .ZN(new_n13557_));
  AOI21_X1   g12537(.A1(new_n13557_), .A2(new_n13533_), .B(\A[745] ), .ZN(new_n13558_));
  NOR2_X1    g12538(.A1(new_n13558_), .A2(new_n13556_), .ZN(new_n13559_));
  NAND2_X1   g12539(.A1(new_n13546_), .A2(\A[750] ), .ZN(new_n13560_));
  NAND2_X1   g12540(.A1(new_n13544_), .A2(\A[749] ), .ZN(new_n13561_));
  AOI21_X1   g12541(.A1(new_n13560_), .A2(new_n13561_), .B(new_n13527_), .ZN(new_n13562_));
  INV_X1     g12542(.I(new_n13528_), .ZN(new_n13563_));
  AOI21_X1   g12543(.A1(new_n13563_), .A2(new_n13529_), .B(\A[748] ), .ZN(new_n13564_));
  NOR2_X1    g12544(.A1(new_n13564_), .A2(new_n13562_), .ZN(new_n13565_));
  NAND2_X1   g12545(.A1(new_n13559_), .A2(new_n13565_), .ZN(new_n13566_));
  NOR2_X1    g12546(.A1(new_n13566_), .A2(new_n13534_), .ZN(new_n13567_));
  OAI21_X1   g12547(.A1(new_n13553_), .A2(new_n13567_), .B(new_n13530_), .ZN(new_n13568_));
  INV_X1     g12548(.I(new_n13530_), .ZN(new_n13569_));
  NAND2_X1   g12549(.A1(new_n13566_), .A2(new_n13534_), .ZN(new_n13570_));
  NAND2_X1   g12550(.A1(new_n13552_), .A2(new_n13535_), .ZN(new_n13571_));
  NAND3_X1   g12551(.A1(new_n13571_), .A2(new_n13570_), .A3(new_n13569_), .ZN(new_n13572_));
  NAND2_X1   g12552(.A1(new_n13568_), .A2(new_n13572_), .ZN(new_n13573_));
  NOR2_X1    g12553(.A1(new_n13510_), .A2(new_n13508_), .ZN(new_n13574_));
  NOR2_X1    g12554(.A1(new_n13517_), .A2(new_n13515_), .ZN(new_n13575_));
  NAND2_X1   g12555(.A1(new_n13574_), .A2(new_n13575_), .ZN(new_n13576_));
  NAND2_X1   g12556(.A1(new_n13498_), .A2(new_n13502_), .ZN(new_n13577_));
  NOR2_X1    g12557(.A1(new_n13559_), .A2(new_n13565_), .ZN(new_n13578_));
  NOR4_X1    g12558(.A1(new_n13552_), .A2(new_n13578_), .A3(new_n13576_), .A4(new_n13577_), .ZN(new_n13579_));
  NOR2_X1    g12559(.A1(new_n13574_), .A2(new_n13575_), .ZN(new_n13580_));
  NOR2_X1    g12560(.A1(new_n13580_), .A2(new_n13518_), .ZN(new_n13581_));
  NAND2_X1   g12561(.A1(new_n13530_), .A2(new_n13534_), .ZN(new_n13582_));
  NOR3_X1    g12562(.A1(new_n13543_), .A2(new_n13551_), .A3(new_n13582_), .ZN(new_n13583_));
  NAND3_X1   g12563(.A1(new_n13579_), .A2(new_n13581_), .A3(new_n13583_), .ZN(new_n13584_));
  INV_X1     g12564(.I(new_n13584_), .ZN(new_n13585_));
  NAND2_X1   g12565(.A1(new_n13585_), .A2(new_n13573_), .ZN(new_n13586_));
  AOI21_X1   g12566(.A1(new_n13571_), .A2(new_n13570_), .B(new_n13569_), .ZN(new_n13587_));
  NOR3_X1    g12567(.A1(new_n13553_), .A2(new_n13567_), .A3(new_n13530_), .ZN(new_n13588_));
  NOR2_X1    g12568(.A1(new_n13587_), .A2(new_n13588_), .ZN(new_n13589_));
  NAND2_X1   g12569(.A1(new_n13589_), .A2(new_n13584_), .ZN(new_n13590_));
  AOI21_X1   g12570(.A1(new_n13586_), .A2(new_n13590_), .B(new_n13526_), .ZN(new_n13591_));
  NAND2_X1   g12571(.A1(new_n13579_), .A2(new_n13581_), .ZN(new_n13592_));
  INV_X1     g12572(.I(new_n13592_), .ZN(new_n13593_));
  NOR2_X1    g12573(.A1(new_n13578_), .A2(new_n13582_), .ZN(new_n13594_));
  AOI21_X1   g12574(.A1(new_n13589_), .A2(new_n13593_), .B(new_n13594_), .ZN(new_n13595_));
  NOR2_X1    g12575(.A1(new_n13573_), .A2(new_n13584_), .ZN(new_n13596_));
  NOR3_X1    g12576(.A1(new_n13595_), .A2(new_n13596_), .A3(new_n13526_), .ZN(new_n13597_));
  NOR2_X1    g12577(.A1(new_n13597_), .A2(new_n13591_), .ZN(new_n13598_));
  INV_X1     g12578(.I(new_n13526_), .ZN(new_n13599_));
  NOR2_X1    g12579(.A1(new_n13589_), .A2(new_n13584_), .ZN(new_n13600_));
  NOR2_X1    g12580(.A1(new_n13585_), .A2(new_n13573_), .ZN(new_n13601_));
  OAI21_X1   g12581(.A1(new_n13601_), .A2(new_n13600_), .B(new_n13599_), .ZN(new_n13602_));
  OAI22_X1   g12582(.A1(new_n13573_), .A2(new_n13592_), .B1(new_n13578_), .B2(new_n13582_), .ZN(new_n13603_));
  NAND2_X1   g12583(.A1(new_n13585_), .A2(new_n13589_), .ZN(new_n13604_));
  NAND3_X1   g12584(.A1(new_n13603_), .A2(new_n13604_), .A3(new_n13599_), .ZN(new_n13605_));
  NOR2_X1    g12585(.A1(new_n13578_), .A2(new_n13552_), .ZN(new_n13606_));
  NAND2_X1   g12586(.A1(new_n13606_), .A2(new_n13583_), .ZN(new_n13607_));
  NOR2_X1    g12587(.A1(new_n13576_), .A2(new_n13577_), .ZN(new_n13608_));
  NAND2_X1   g12588(.A1(new_n13581_), .A2(new_n13608_), .ZN(new_n13609_));
  XOR2_X1    g12589(.A1(new_n13609_), .A2(new_n13607_), .Z(new_n13610_));
  INV_X1     g12590(.I(\A[735] ), .ZN(new_n13611_));
  NOR2_X1    g12591(.A1(new_n13611_), .A2(\A[734] ), .ZN(new_n13612_));
  INV_X1     g12592(.I(\A[734] ), .ZN(new_n13613_));
  NOR2_X1    g12593(.A1(new_n13613_), .A2(\A[735] ), .ZN(new_n13614_));
  OAI21_X1   g12594(.A1(new_n13612_), .A2(new_n13614_), .B(\A[733] ), .ZN(new_n13615_));
  INV_X1     g12595(.I(\A[733] ), .ZN(new_n13616_));
  NOR2_X1    g12596(.A1(\A[734] ), .A2(\A[735] ), .ZN(new_n13617_));
  NAND2_X1   g12597(.A1(\A[734] ), .A2(\A[735] ), .ZN(new_n13618_));
  INV_X1     g12598(.I(new_n13618_), .ZN(new_n13619_));
  OAI21_X1   g12599(.A1(new_n13619_), .A2(new_n13617_), .B(new_n13616_), .ZN(new_n13620_));
  NAND2_X1   g12600(.A1(new_n13615_), .A2(new_n13620_), .ZN(new_n13621_));
  INV_X1     g12601(.I(\A[738] ), .ZN(new_n13622_));
  NOR2_X1    g12602(.A1(new_n13622_), .A2(\A[737] ), .ZN(new_n13623_));
  INV_X1     g12603(.I(\A[737] ), .ZN(new_n13624_));
  NOR2_X1    g12604(.A1(new_n13624_), .A2(\A[738] ), .ZN(new_n13625_));
  OAI21_X1   g12605(.A1(new_n13623_), .A2(new_n13625_), .B(\A[736] ), .ZN(new_n13626_));
  INV_X1     g12606(.I(\A[736] ), .ZN(new_n13627_));
  NOR2_X1    g12607(.A1(\A[737] ), .A2(\A[738] ), .ZN(new_n13628_));
  NAND2_X1   g12608(.A1(\A[737] ), .A2(\A[738] ), .ZN(new_n13629_));
  INV_X1     g12609(.I(new_n13629_), .ZN(new_n13630_));
  OAI21_X1   g12610(.A1(new_n13630_), .A2(new_n13628_), .B(new_n13627_), .ZN(new_n13631_));
  NAND2_X1   g12611(.A1(new_n13626_), .A2(new_n13631_), .ZN(new_n13632_));
  NOR2_X1    g12612(.A1(new_n13621_), .A2(new_n13632_), .ZN(new_n13633_));
  NAND2_X1   g12613(.A1(new_n13613_), .A2(\A[735] ), .ZN(new_n13634_));
  NAND2_X1   g12614(.A1(new_n13611_), .A2(\A[734] ), .ZN(new_n13635_));
  AOI21_X1   g12615(.A1(new_n13634_), .A2(new_n13635_), .B(new_n13616_), .ZN(new_n13636_));
  INV_X1     g12616(.I(new_n13617_), .ZN(new_n13637_));
  AOI21_X1   g12617(.A1(new_n13637_), .A2(new_n13618_), .B(\A[733] ), .ZN(new_n13638_));
  NOR2_X1    g12618(.A1(new_n13638_), .A2(new_n13636_), .ZN(new_n13639_));
  NAND2_X1   g12619(.A1(new_n13624_), .A2(\A[738] ), .ZN(new_n13640_));
  NAND2_X1   g12620(.A1(new_n13622_), .A2(\A[737] ), .ZN(new_n13641_));
  AOI21_X1   g12621(.A1(new_n13640_), .A2(new_n13641_), .B(new_n13627_), .ZN(new_n13642_));
  INV_X1     g12622(.I(new_n13628_), .ZN(new_n13643_));
  AOI21_X1   g12623(.A1(new_n13643_), .A2(new_n13629_), .B(\A[736] ), .ZN(new_n13644_));
  NOR2_X1    g12624(.A1(new_n13644_), .A2(new_n13642_), .ZN(new_n13645_));
  NOR2_X1    g12625(.A1(new_n13639_), .A2(new_n13645_), .ZN(new_n13646_));
  NOR2_X1    g12626(.A1(new_n13646_), .A2(new_n13633_), .ZN(new_n13647_));
  AOI21_X1   g12627(.A1(new_n13627_), .A2(new_n13629_), .B(new_n13628_), .ZN(new_n13648_));
  AOI21_X1   g12628(.A1(new_n13616_), .A2(new_n13618_), .B(new_n13617_), .ZN(new_n13649_));
  NAND2_X1   g12629(.A1(new_n13648_), .A2(new_n13649_), .ZN(new_n13650_));
  NOR3_X1    g12630(.A1(new_n13621_), .A2(new_n13632_), .A3(new_n13650_), .ZN(new_n13651_));
  INV_X1     g12631(.I(\A[730] ), .ZN(new_n13652_));
  NOR2_X1    g12632(.A1(\A[731] ), .A2(\A[732] ), .ZN(new_n13653_));
  NAND2_X1   g12633(.A1(\A[731] ), .A2(\A[732] ), .ZN(new_n13654_));
  AOI21_X1   g12634(.A1(new_n13652_), .A2(new_n13654_), .B(new_n13653_), .ZN(new_n13655_));
  INV_X1     g12635(.I(new_n13655_), .ZN(new_n13656_));
  INV_X1     g12636(.I(\A[727] ), .ZN(new_n13657_));
  NOR2_X1    g12637(.A1(\A[728] ), .A2(\A[729] ), .ZN(new_n13658_));
  NAND2_X1   g12638(.A1(\A[728] ), .A2(\A[729] ), .ZN(new_n13659_));
  AOI21_X1   g12639(.A1(new_n13657_), .A2(new_n13659_), .B(new_n13658_), .ZN(new_n13660_));
  INV_X1     g12640(.I(new_n13660_), .ZN(new_n13661_));
  NOR2_X1    g12641(.A1(new_n13656_), .A2(new_n13661_), .ZN(new_n13662_));
  INV_X1     g12642(.I(\A[728] ), .ZN(new_n13663_));
  NAND2_X1   g12643(.A1(new_n13663_), .A2(\A[729] ), .ZN(new_n13664_));
  INV_X1     g12644(.I(\A[729] ), .ZN(new_n13665_));
  NAND2_X1   g12645(.A1(new_n13665_), .A2(\A[728] ), .ZN(new_n13666_));
  AOI21_X1   g12646(.A1(new_n13664_), .A2(new_n13666_), .B(new_n13657_), .ZN(new_n13667_));
  INV_X1     g12647(.I(new_n13658_), .ZN(new_n13668_));
  AOI21_X1   g12648(.A1(new_n13668_), .A2(new_n13659_), .B(\A[727] ), .ZN(new_n13669_));
  NOR2_X1    g12649(.A1(new_n13669_), .A2(new_n13667_), .ZN(new_n13670_));
  INV_X1     g12650(.I(\A[731] ), .ZN(new_n13671_));
  NAND2_X1   g12651(.A1(new_n13671_), .A2(\A[732] ), .ZN(new_n13672_));
  INV_X1     g12652(.I(\A[732] ), .ZN(new_n13673_));
  NAND2_X1   g12653(.A1(new_n13673_), .A2(\A[731] ), .ZN(new_n13674_));
  AOI21_X1   g12654(.A1(new_n13672_), .A2(new_n13674_), .B(new_n13652_), .ZN(new_n13675_));
  INV_X1     g12655(.I(new_n13653_), .ZN(new_n13676_));
  AOI21_X1   g12656(.A1(new_n13676_), .A2(new_n13654_), .B(\A[730] ), .ZN(new_n13677_));
  NOR2_X1    g12657(.A1(new_n13677_), .A2(new_n13675_), .ZN(new_n13678_));
  NAND2_X1   g12658(.A1(new_n13647_), .A2(new_n13651_), .ZN(new_n13679_));
  INV_X1     g12659(.I(new_n13679_), .ZN(new_n13680_));
  NOR2_X1    g12660(.A1(new_n13610_), .A2(new_n13680_), .ZN(new_n13681_));
  AOI21_X1   g12661(.A1(new_n13605_), .A2(new_n13602_), .B(new_n13681_), .ZN(new_n13682_));
  XNOR2_X1   g12662(.A1(new_n13609_), .A2(new_n13607_), .ZN(new_n13683_));
  NAND2_X1   g12663(.A1(new_n13683_), .A2(new_n13679_), .ZN(new_n13684_));
  NOR3_X1    g12664(.A1(new_n13597_), .A2(new_n13684_), .A3(new_n13591_), .ZN(new_n13685_));
  INV_X1     g12665(.I(new_n13649_), .ZN(new_n13686_));
  NOR2_X1    g12666(.A1(new_n13633_), .A2(new_n13686_), .ZN(new_n13687_));
  NAND2_X1   g12667(.A1(new_n13639_), .A2(new_n13645_), .ZN(new_n13688_));
  NOR2_X1    g12668(.A1(new_n13688_), .A2(new_n13649_), .ZN(new_n13689_));
  OAI21_X1   g12669(.A1(new_n13687_), .A2(new_n13689_), .B(new_n13648_), .ZN(new_n13690_));
  INV_X1     g12670(.I(new_n13648_), .ZN(new_n13691_));
  NAND2_X1   g12671(.A1(new_n13688_), .A2(new_n13649_), .ZN(new_n13692_));
  NAND2_X1   g12672(.A1(new_n13633_), .A2(new_n13686_), .ZN(new_n13693_));
  NAND3_X1   g12673(.A1(new_n13693_), .A2(new_n13692_), .A3(new_n13691_), .ZN(new_n13694_));
  NAND2_X1   g12674(.A1(new_n13690_), .A2(new_n13694_), .ZN(new_n13695_));
  NOR4_X1    g12675(.A1(new_n13667_), .A2(new_n13669_), .A3(new_n13677_), .A4(new_n13675_), .ZN(new_n13696_));
  NOR2_X1    g12676(.A1(new_n13670_), .A2(new_n13678_), .ZN(new_n13697_));
  NOR2_X1    g12677(.A1(new_n13697_), .A2(new_n13696_), .ZN(new_n13698_));
  INV_X1     g12678(.I(new_n13662_), .ZN(new_n13699_));
  NAND2_X1   g12679(.A1(new_n13670_), .A2(new_n13678_), .ZN(new_n13700_));
  NOR4_X1    g12680(.A1(new_n13633_), .A2(new_n13646_), .A3(new_n13700_), .A4(new_n13699_), .ZN(new_n13701_));
  NAND2_X1   g12681(.A1(new_n13701_), .A2(new_n13698_), .ZN(new_n13702_));
  INV_X1     g12682(.I(new_n13650_), .ZN(new_n13703_));
  OAI21_X1   g12683(.A1(new_n13639_), .A2(new_n13645_), .B(new_n13703_), .ZN(new_n13704_));
  OAI21_X1   g12684(.A1(new_n13695_), .A2(new_n13702_), .B(new_n13704_), .ZN(new_n13705_));
  NAND2_X1   g12685(.A1(new_n13700_), .A2(new_n13660_), .ZN(new_n13706_));
  NAND2_X1   g12686(.A1(new_n13696_), .A2(new_n13661_), .ZN(new_n13707_));
  AOI21_X1   g12687(.A1(new_n13706_), .A2(new_n13707_), .B(new_n13656_), .ZN(new_n13708_));
  NOR2_X1    g12688(.A1(new_n13696_), .A2(new_n13661_), .ZN(new_n13709_));
  NOR2_X1    g12689(.A1(new_n13700_), .A2(new_n13660_), .ZN(new_n13710_));
  NOR3_X1    g12690(.A1(new_n13710_), .A2(new_n13655_), .A3(new_n13709_), .ZN(new_n13711_));
  NOR2_X1    g12691(.A1(new_n13711_), .A2(new_n13708_), .ZN(new_n13712_));
  NOR2_X1    g12692(.A1(new_n13705_), .A2(new_n13712_), .ZN(new_n13713_));
  NAND3_X1   g12693(.A1(new_n13647_), .A2(new_n13662_), .A3(new_n13696_), .ZN(new_n13714_));
  NAND2_X1   g12694(.A1(new_n13698_), .A2(new_n13651_), .ZN(new_n13715_));
  NOR2_X1    g12695(.A1(new_n13714_), .A2(new_n13715_), .ZN(new_n13716_));
  NOR2_X1    g12696(.A1(new_n13712_), .A2(new_n13716_), .ZN(new_n13717_));
  INV_X1     g12697(.I(new_n13717_), .ZN(new_n13718_));
  OAI21_X1   g12698(.A1(new_n13710_), .A2(new_n13709_), .B(new_n13655_), .ZN(new_n13719_));
  NAND3_X1   g12699(.A1(new_n13706_), .A2(new_n13656_), .A3(new_n13707_), .ZN(new_n13720_));
  NAND2_X1   g12700(.A1(new_n13703_), .A2(new_n13639_), .ZN(new_n13721_));
  NOR4_X1    g12701(.A1(new_n13721_), .A2(new_n13697_), .A3(new_n13632_), .A4(new_n13696_), .ZN(new_n13722_));
  NAND4_X1   g12702(.A1(new_n13719_), .A2(new_n13720_), .A3(new_n13701_), .A4(new_n13722_), .ZN(new_n13723_));
  XOR2_X1    g12703(.A1(new_n13723_), .A2(new_n13695_), .Z(new_n13724_));
  AOI21_X1   g12704(.A1(new_n13724_), .A2(new_n13718_), .B(new_n13713_), .ZN(new_n13725_));
  OAI22_X1   g12705(.A1(new_n13682_), .A2(new_n13685_), .B1(new_n13725_), .B2(new_n13598_), .ZN(new_n13726_));
  OAI21_X1   g12706(.A1(new_n13573_), .A2(new_n13584_), .B(new_n13526_), .ZN(new_n13727_));
  NOR2_X1    g12707(.A1(new_n13530_), .A2(new_n13534_), .ZN(new_n13728_));
  OAI21_X1   g12708(.A1(new_n13566_), .A2(new_n13728_), .B(new_n13582_), .ZN(new_n13729_));
  NOR2_X1    g12709(.A1(new_n13498_), .A2(new_n13502_), .ZN(new_n13730_));
  OAI21_X1   g12710(.A1(new_n13576_), .A2(new_n13730_), .B(new_n13577_), .ZN(new_n13731_));
  XNOR2_X1   g12711(.A1(new_n13729_), .A2(new_n13731_), .ZN(new_n13732_));
  NAND3_X1   g12712(.A1(new_n13727_), .A2(new_n13603_), .A3(new_n13732_), .ZN(new_n13733_));
  INV_X1     g12713(.I(new_n13712_), .ZN(new_n13734_));
  AOI21_X1   g12714(.A1(new_n13693_), .A2(new_n13692_), .B(new_n13691_), .ZN(new_n13735_));
  NOR3_X1    g12715(.A1(new_n13687_), .A2(new_n13689_), .A3(new_n13648_), .ZN(new_n13736_));
  NOR2_X1    g12716(.A1(new_n13735_), .A2(new_n13736_), .ZN(new_n13737_));
  NAND2_X1   g12717(.A1(new_n13737_), .A2(new_n13716_), .ZN(new_n13738_));
  NAND2_X1   g12718(.A1(new_n13738_), .A2(new_n13734_), .ZN(new_n13739_));
  NOR2_X1    g12719(.A1(new_n13648_), .A2(new_n13649_), .ZN(new_n13740_));
  OAI21_X1   g12720(.A1(new_n13688_), .A2(new_n13740_), .B(new_n13650_), .ZN(new_n13741_));
  NOR2_X1    g12721(.A1(new_n13655_), .A2(new_n13660_), .ZN(new_n13742_));
  OAI21_X1   g12722(.A1(new_n13700_), .A2(new_n13742_), .B(new_n13699_), .ZN(new_n13743_));
  XNOR2_X1   g12723(.A1(new_n13743_), .A2(new_n13741_), .ZN(new_n13744_));
  NAND3_X1   g12724(.A1(new_n13739_), .A2(new_n13744_), .A3(new_n13705_), .ZN(new_n13745_));
  XNOR2_X1   g12725(.A1(new_n13745_), .A2(new_n13733_), .ZN(new_n13746_));
  NOR2_X1    g12726(.A1(new_n13746_), .A2(new_n13726_), .ZN(new_n13747_));
  NAND2_X1   g12727(.A1(new_n13605_), .A2(new_n13602_), .ZN(new_n13748_));
  OAI21_X1   g12728(.A1(new_n13597_), .A2(new_n13591_), .B(new_n13684_), .ZN(new_n13749_));
  NAND3_X1   g12729(.A1(new_n13602_), .A2(new_n13605_), .A3(new_n13681_), .ZN(new_n13750_));
  AOI21_X1   g12730(.A1(new_n13712_), .A2(new_n13716_), .B(new_n13695_), .ZN(new_n13751_));
  NOR2_X1    g12731(.A1(new_n13723_), .A2(new_n13737_), .ZN(new_n13752_));
  NOR2_X1    g12732(.A1(new_n13751_), .A2(new_n13752_), .ZN(new_n13753_));
  OAI22_X1   g12733(.A1(new_n13753_), .A2(new_n13717_), .B1(new_n13705_), .B2(new_n13712_), .ZN(new_n13754_));
  AOI22_X1   g12734(.A1(new_n13749_), .A2(new_n13750_), .B1(new_n13754_), .B2(new_n13748_), .ZN(new_n13755_));
  NAND2_X1   g12735(.A1(new_n13745_), .A2(new_n13733_), .ZN(new_n13756_));
  AOI21_X1   g12736(.A1(new_n13526_), .A2(new_n13604_), .B(new_n13595_), .ZN(new_n13757_));
  NAND3_X1   g12737(.A1(new_n13737_), .A2(new_n13698_), .A3(new_n13701_), .ZN(new_n13758_));
  AOI22_X1   g12738(.A1(new_n13758_), .A2(new_n13704_), .B1(new_n13738_), .B2(new_n13734_), .ZN(new_n13759_));
  NAND4_X1   g12739(.A1(new_n13757_), .A2(new_n13759_), .A3(new_n13732_), .A4(new_n13744_), .ZN(new_n13760_));
  AOI21_X1   g12740(.A1(new_n13756_), .A2(new_n13760_), .B(new_n13755_), .ZN(new_n13761_));
  NOR2_X1    g12741(.A1(new_n13761_), .A2(new_n13747_), .ZN(new_n13762_));
  NAND2_X1   g12742(.A1(new_n13494_), .A2(new_n13762_), .ZN(new_n13763_));
  NOR3_X1    g12743(.A1(new_n13685_), .A2(new_n13754_), .A3(new_n13682_), .ZN(new_n13764_));
  NOR2_X1    g12744(.A1(new_n13683_), .A2(new_n13679_), .ZN(new_n13765_));
  NOR2_X1    g12745(.A1(new_n13765_), .A2(new_n13681_), .ZN(new_n13766_));
  NOR2_X1    g12746(.A1(new_n13402_), .A2(new_n13398_), .ZN(new_n13767_));
  NOR2_X1    g12747(.A1(new_n13767_), .A2(new_n13400_), .ZN(new_n13768_));
  NAND2_X1   g12748(.A1(new_n13766_), .A2(new_n13768_), .ZN(new_n13769_));
  INV_X1     g12749(.I(new_n13769_), .ZN(new_n13770_));
  NOR2_X1    g12750(.A1(new_n13770_), .A2(new_n13764_), .ZN(new_n13771_));
  NAND2_X1   g12751(.A1(new_n13770_), .A2(new_n13764_), .ZN(new_n13772_));
  INV_X1     g12752(.I(new_n13772_), .ZN(new_n13773_));
  AOI21_X1   g12753(.A1(new_n13473_), .A2(new_n13474_), .B(new_n13482_), .ZN(new_n13774_));
  NOR3_X1    g12754(.A1(new_n13452_), .A2(new_n13401_), .A3(new_n13404_), .ZN(new_n13775_));
  NOR2_X1    g12755(.A1(new_n13774_), .A2(new_n13775_), .ZN(new_n13776_));
  OAI22_X1   g12756(.A1(new_n13773_), .A2(new_n13771_), .B1(new_n13776_), .B2(new_n13764_), .ZN(new_n13777_));
  XOR2_X1    g12757(.A1(new_n13490_), .A2(new_n13469_), .Z(new_n13778_));
  NAND2_X1   g12758(.A1(new_n13778_), .A2(new_n13483_), .ZN(new_n13779_));
  NAND2_X1   g12759(.A1(new_n13490_), .A2(new_n13469_), .ZN(new_n13780_));
  NAND2_X1   g12760(.A1(new_n13461_), .A2(new_n13487_), .ZN(new_n13781_));
  NAND2_X1   g12761(.A1(new_n13781_), .A2(new_n13780_), .ZN(new_n13782_));
  NAND2_X1   g12762(.A1(new_n13453_), .A2(new_n13782_), .ZN(new_n13783_));
  XOR2_X1    g12763(.A1(new_n13745_), .A2(new_n13733_), .Z(new_n13784_));
  NAND2_X1   g12764(.A1(new_n13784_), .A2(new_n13755_), .ZN(new_n13785_));
  NAND2_X1   g12765(.A1(new_n13760_), .A2(new_n13756_), .ZN(new_n13786_));
  NAND2_X1   g12766(.A1(new_n13726_), .A2(new_n13786_), .ZN(new_n13787_));
  AOI22_X1   g12767(.A1(new_n13779_), .A2(new_n13783_), .B1(new_n13785_), .B2(new_n13787_), .ZN(new_n13788_));
  OAI21_X1   g12768(.A1(new_n13777_), .A2(new_n13788_), .B(new_n13763_), .ZN(new_n13789_));
  NAND2_X1   g12769(.A1(new_n13456_), .A2(new_n13458_), .ZN(new_n13790_));
  NOR2_X1    g12770(.A1(new_n13454_), .A2(new_n13325_), .ZN(new_n13791_));
  OAI21_X1   g12771(.A1(new_n13456_), .A2(new_n13458_), .B(new_n13791_), .ZN(new_n13792_));
  NAND2_X1   g12772(.A1(new_n13792_), .A2(new_n13790_), .ZN(new_n13793_));
  NAND2_X1   g12773(.A1(new_n13467_), .A2(new_n13465_), .ZN(new_n13794_));
  OR2_X2     g12774(.A1(new_n13467_), .A2(new_n13465_), .Z(new_n13795_));
  NAND3_X1   g12775(.A1(new_n13463_), .A2(new_n13436_), .A3(new_n13795_), .ZN(new_n13796_));
  NAND2_X1   g12776(.A1(new_n13796_), .A2(new_n13794_), .ZN(new_n13797_));
  INV_X1     g12777(.I(new_n13797_), .ZN(new_n13798_));
  NAND2_X1   g12778(.A1(new_n13453_), .A2(new_n13780_), .ZN(new_n13799_));
  AOI21_X1   g12779(.A1(new_n13799_), .A2(new_n13491_), .B(new_n13798_), .ZN(new_n13800_));
  NAND4_X1   g12780(.A1(new_n13483_), .A2(new_n13798_), .A3(new_n13461_), .A4(new_n13487_), .ZN(new_n13801_));
  INV_X1     g12781(.I(new_n13801_), .ZN(new_n13802_));
  OAI21_X1   g12782(.A1(new_n13800_), .A2(new_n13802_), .B(new_n13793_), .ZN(new_n13803_));
  INV_X1     g12783(.I(new_n13793_), .ZN(new_n13804_));
  NAND3_X1   g12784(.A1(new_n13483_), .A2(new_n13461_), .A3(new_n13487_), .ZN(new_n13805_));
  NAND2_X1   g12785(.A1(new_n13805_), .A2(new_n13797_), .ZN(new_n13806_));
  NAND3_X1   g12786(.A1(new_n13806_), .A2(new_n13804_), .A3(new_n13801_), .ZN(new_n13807_));
  NAND2_X1   g12787(.A1(new_n13803_), .A2(new_n13807_), .ZN(new_n13808_));
  INV_X1     g12788(.I(new_n13757_), .ZN(new_n13809_));
  NAND2_X1   g12789(.A1(new_n13729_), .A2(new_n13731_), .ZN(new_n13810_));
  NOR2_X1    g12790(.A1(new_n13729_), .A2(new_n13731_), .ZN(new_n13811_));
  OAI21_X1   g12791(.A1(new_n13809_), .A2(new_n13811_), .B(new_n13810_), .ZN(new_n13812_));
  NAND2_X1   g12792(.A1(new_n13743_), .A2(new_n13741_), .ZN(new_n13813_));
  OAI21_X1   g12793(.A1(new_n13741_), .A2(new_n13743_), .B(new_n13759_), .ZN(new_n13814_));
  NAND2_X1   g12794(.A1(new_n13814_), .A2(new_n13813_), .ZN(new_n13815_));
  INV_X1     g12795(.I(new_n13815_), .ZN(new_n13816_));
  AOI21_X1   g12796(.A1(new_n13726_), .A2(new_n13756_), .B(new_n13760_), .ZN(new_n13817_));
  NOR2_X1    g12797(.A1(new_n13817_), .A2(new_n13816_), .ZN(new_n13818_));
  INV_X1     g12798(.I(new_n13733_), .ZN(new_n13819_));
  INV_X1     g12799(.I(new_n13745_), .ZN(new_n13820_));
  NAND3_X1   g12800(.A1(new_n13755_), .A2(new_n13819_), .A3(new_n13820_), .ZN(new_n13821_));
  NOR2_X1    g12801(.A1(new_n13821_), .A2(new_n13815_), .ZN(new_n13822_));
  OAI21_X1   g12802(.A1(new_n13818_), .A2(new_n13822_), .B(new_n13812_), .ZN(new_n13823_));
  INV_X1     g12803(.I(new_n13812_), .ZN(new_n13824_));
  NAND2_X1   g12804(.A1(new_n13821_), .A2(new_n13815_), .ZN(new_n13825_));
  NAND4_X1   g12805(.A1(new_n13816_), .A2(new_n13755_), .A3(new_n13819_), .A4(new_n13820_), .ZN(new_n13826_));
  NAND3_X1   g12806(.A1(new_n13825_), .A2(new_n13824_), .A3(new_n13826_), .ZN(new_n13827_));
  NAND2_X1   g12807(.A1(new_n13823_), .A2(new_n13827_), .ZN(new_n13828_));
  NOR2_X1    g12808(.A1(new_n13808_), .A2(new_n13828_), .ZN(new_n13829_));
  NOR2_X1    g12809(.A1(new_n13829_), .A2(new_n13789_), .ZN(new_n13830_));
  XOR2_X1    g12810(.A1(new_n13793_), .A2(new_n13797_), .Z(new_n13831_));
  XNOR2_X1   g12811(.A1(new_n13815_), .A2(new_n13812_), .ZN(new_n13832_));
  INV_X1     g12812(.I(new_n13832_), .ZN(new_n13833_));
  NOR4_X1    g12813(.A1(new_n13833_), .A2(new_n13831_), .A3(new_n13805_), .A4(new_n13821_), .ZN(new_n13834_));
  INV_X1     g12814(.I(new_n13834_), .ZN(new_n13835_));
  NOR2_X1    g12815(.A1(new_n13830_), .A2(new_n13835_), .ZN(new_n13836_));
  OAI21_X1   g12816(.A1(new_n13793_), .A2(new_n13797_), .B(new_n13805_), .ZN(new_n13837_));
  OAI21_X1   g12817(.A1(new_n13812_), .A2(new_n13815_), .B(new_n13821_), .ZN(new_n13838_));
  NAND2_X1   g12818(.A1(new_n13815_), .A2(new_n13812_), .ZN(new_n13839_));
  NAND2_X1   g12819(.A1(new_n13793_), .A2(new_n13797_), .ZN(new_n13840_));
  NAND4_X1   g12820(.A1(new_n13837_), .A2(new_n13838_), .A3(new_n13839_), .A4(new_n13840_), .ZN(new_n13841_));
  NAND2_X1   g12821(.A1(new_n13838_), .A2(new_n13839_), .ZN(new_n13842_));
  NAND2_X1   g12822(.A1(new_n13837_), .A2(new_n13840_), .ZN(new_n13843_));
  NAND2_X1   g12823(.A1(new_n13843_), .A2(new_n13842_), .ZN(new_n13844_));
  OAI21_X1   g12824(.A1(new_n13836_), .A2(new_n13841_), .B(new_n13844_), .ZN(new_n13845_));
  INV_X1     g12825(.I(new_n13845_), .ZN(new_n13846_));
  INV_X1     g12826(.I(\A[694] ), .ZN(new_n13847_));
  NOR2_X1    g12827(.A1(\A[695] ), .A2(\A[696] ), .ZN(new_n13848_));
  NAND2_X1   g12828(.A1(\A[695] ), .A2(\A[696] ), .ZN(new_n13849_));
  AOI21_X1   g12829(.A1(new_n13847_), .A2(new_n13849_), .B(new_n13848_), .ZN(new_n13850_));
  INV_X1     g12830(.I(new_n13850_), .ZN(new_n13851_));
  INV_X1     g12831(.I(\A[691] ), .ZN(new_n13852_));
  NOR2_X1    g12832(.A1(\A[692] ), .A2(\A[693] ), .ZN(new_n13853_));
  NAND2_X1   g12833(.A1(\A[692] ), .A2(\A[693] ), .ZN(new_n13854_));
  AOI21_X1   g12834(.A1(new_n13852_), .A2(new_n13854_), .B(new_n13853_), .ZN(new_n13855_));
  INV_X1     g12835(.I(new_n13855_), .ZN(new_n13856_));
  INV_X1     g12836(.I(\A[692] ), .ZN(new_n13857_));
  NAND2_X1   g12837(.A1(new_n13857_), .A2(\A[693] ), .ZN(new_n13858_));
  INV_X1     g12838(.I(\A[693] ), .ZN(new_n13859_));
  NAND2_X1   g12839(.A1(new_n13859_), .A2(\A[692] ), .ZN(new_n13860_));
  AOI21_X1   g12840(.A1(new_n13858_), .A2(new_n13860_), .B(new_n13852_), .ZN(new_n13861_));
  INV_X1     g12841(.I(new_n13853_), .ZN(new_n13862_));
  AOI21_X1   g12842(.A1(new_n13862_), .A2(new_n13854_), .B(\A[691] ), .ZN(new_n13863_));
  INV_X1     g12843(.I(\A[695] ), .ZN(new_n13864_));
  NAND2_X1   g12844(.A1(new_n13864_), .A2(\A[696] ), .ZN(new_n13865_));
  INV_X1     g12845(.I(\A[696] ), .ZN(new_n13866_));
  NAND2_X1   g12846(.A1(new_n13866_), .A2(\A[695] ), .ZN(new_n13867_));
  AOI21_X1   g12847(.A1(new_n13865_), .A2(new_n13867_), .B(new_n13847_), .ZN(new_n13868_));
  INV_X1     g12848(.I(new_n13848_), .ZN(new_n13869_));
  AOI21_X1   g12849(.A1(new_n13869_), .A2(new_n13849_), .B(\A[694] ), .ZN(new_n13870_));
  NOR4_X1    g12850(.A1(new_n13861_), .A2(new_n13863_), .A3(new_n13870_), .A4(new_n13868_), .ZN(new_n13871_));
  NOR2_X1    g12851(.A1(new_n13871_), .A2(new_n13856_), .ZN(new_n13872_));
  INV_X1     g12852(.I(new_n13872_), .ZN(new_n13873_));
  NAND2_X1   g12853(.A1(new_n13871_), .A2(new_n13856_), .ZN(new_n13874_));
  AOI21_X1   g12854(.A1(new_n13873_), .A2(new_n13874_), .B(new_n13851_), .ZN(new_n13875_));
  INV_X1     g12855(.I(new_n13874_), .ZN(new_n13876_));
  NOR3_X1    g12856(.A1(new_n13876_), .A2(new_n13850_), .A3(new_n13872_), .ZN(new_n13877_));
  NOR2_X1    g12857(.A1(new_n13875_), .A2(new_n13877_), .ZN(new_n13878_));
  INV_X1     g12858(.I(\A[700] ), .ZN(new_n13879_));
  NOR2_X1    g12859(.A1(\A[701] ), .A2(\A[702] ), .ZN(new_n13880_));
  NAND2_X1   g12860(.A1(\A[701] ), .A2(\A[702] ), .ZN(new_n13881_));
  AOI21_X1   g12861(.A1(new_n13879_), .A2(new_n13881_), .B(new_n13880_), .ZN(new_n13882_));
  INV_X1     g12862(.I(new_n13882_), .ZN(new_n13883_));
  INV_X1     g12863(.I(\A[697] ), .ZN(new_n13884_));
  NOR2_X1    g12864(.A1(\A[698] ), .A2(\A[699] ), .ZN(new_n13885_));
  NAND2_X1   g12865(.A1(\A[698] ), .A2(\A[699] ), .ZN(new_n13886_));
  AOI21_X1   g12866(.A1(new_n13884_), .A2(new_n13886_), .B(new_n13885_), .ZN(new_n13887_));
  INV_X1     g12867(.I(new_n13887_), .ZN(new_n13888_));
  NOR2_X1    g12868(.A1(new_n13883_), .A2(new_n13888_), .ZN(new_n13889_));
  INV_X1     g12869(.I(new_n13889_), .ZN(new_n13890_));
  INV_X1     g12870(.I(\A[698] ), .ZN(new_n13891_));
  NAND2_X1   g12871(.A1(new_n13891_), .A2(\A[699] ), .ZN(new_n13892_));
  INV_X1     g12872(.I(\A[699] ), .ZN(new_n13893_));
  NAND2_X1   g12873(.A1(new_n13893_), .A2(\A[698] ), .ZN(new_n13894_));
  AOI21_X1   g12874(.A1(new_n13892_), .A2(new_n13894_), .B(new_n13884_), .ZN(new_n13895_));
  INV_X1     g12875(.I(new_n13885_), .ZN(new_n13896_));
  AOI21_X1   g12876(.A1(new_n13896_), .A2(new_n13886_), .B(\A[697] ), .ZN(new_n13897_));
  NOR2_X1    g12877(.A1(new_n13897_), .A2(new_n13895_), .ZN(new_n13898_));
  INV_X1     g12878(.I(\A[702] ), .ZN(new_n13899_));
  NOR2_X1    g12879(.A1(new_n13899_), .A2(\A[701] ), .ZN(new_n13900_));
  INV_X1     g12880(.I(\A[701] ), .ZN(new_n13901_));
  NOR2_X1    g12881(.A1(new_n13901_), .A2(\A[702] ), .ZN(new_n13902_));
  OAI21_X1   g12882(.A1(new_n13900_), .A2(new_n13902_), .B(\A[700] ), .ZN(new_n13903_));
  INV_X1     g12883(.I(new_n13881_), .ZN(new_n13904_));
  OAI21_X1   g12884(.A1(new_n13904_), .A2(new_n13880_), .B(new_n13879_), .ZN(new_n13905_));
  NAND2_X1   g12885(.A1(new_n13903_), .A2(new_n13905_), .ZN(new_n13906_));
  NAND2_X1   g12886(.A1(new_n13898_), .A2(new_n13906_), .ZN(new_n13907_));
  NOR2_X1    g12887(.A1(new_n13893_), .A2(\A[698] ), .ZN(new_n13908_));
  NOR2_X1    g12888(.A1(new_n13891_), .A2(\A[699] ), .ZN(new_n13909_));
  OAI21_X1   g12889(.A1(new_n13908_), .A2(new_n13909_), .B(\A[697] ), .ZN(new_n13910_));
  INV_X1     g12890(.I(new_n13886_), .ZN(new_n13911_));
  OAI21_X1   g12891(.A1(new_n13911_), .A2(new_n13885_), .B(new_n13884_), .ZN(new_n13912_));
  NAND2_X1   g12892(.A1(new_n13910_), .A2(new_n13912_), .ZN(new_n13913_));
  NAND2_X1   g12893(.A1(new_n13901_), .A2(\A[702] ), .ZN(new_n13914_));
  NAND2_X1   g12894(.A1(new_n13899_), .A2(\A[701] ), .ZN(new_n13915_));
  AOI21_X1   g12895(.A1(new_n13914_), .A2(new_n13915_), .B(new_n13879_), .ZN(new_n13916_));
  INV_X1     g12896(.I(new_n13880_), .ZN(new_n13917_));
  AOI21_X1   g12897(.A1(new_n13917_), .A2(new_n13881_), .B(\A[700] ), .ZN(new_n13918_));
  NOR2_X1    g12898(.A1(new_n13918_), .A2(new_n13916_), .ZN(new_n13919_));
  NAND2_X1   g12899(.A1(new_n13919_), .A2(new_n13913_), .ZN(new_n13920_));
  AOI21_X1   g12900(.A1(new_n13907_), .A2(new_n13920_), .B(new_n13890_), .ZN(new_n13921_));
  INV_X1     g12901(.I(new_n13921_), .ZN(new_n13922_));
  NOR2_X1    g12902(.A1(new_n13913_), .A2(new_n13906_), .ZN(new_n13923_));
  NOR2_X1    g12903(.A1(new_n13923_), .A2(new_n13888_), .ZN(new_n13924_));
  NAND2_X1   g12904(.A1(new_n13898_), .A2(new_n13919_), .ZN(new_n13925_));
  NOR2_X1    g12905(.A1(new_n13925_), .A2(new_n13887_), .ZN(new_n13926_));
  OAI21_X1   g12906(.A1(new_n13924_), .A2(new_n13926_), .B(new_n13882_), .ZN(new_n13927_));
  NAND2_X1   g12907(.A1(new_n13925_), .A2(new_n13887_), .ZN(new_n13928_));
  NAND2_X1   g12908(.A1(new_n13923_), .A2(new_n13888_), .ZN(new_n13929_));
  NAND3_X1   g12909(.A1(new_n13929_), .A2(new_n13928_), .A3(new_n13883_), .ZN(new_n13930_));
  NAND3_X1   g12910(.A1(new_n13927_), .A2(new_n13930_), .A3(new_n13922_), .ZN(new_n13931_));
  NOR2_X1    g12911(.A1(new_n13925_), .A2(new_n13890_), .ZN(new_n13932_));
  NOR2_X1    g12912(.A1(new_n13898_), .A2(new_n13919_), .ZN(new_n13933_));
  NOR2_X1    g12913(.A1(new_n13933_), .A2(new_n13923_), .ZN(new_n13934_));
  NOR2_X1    g12914(.A1(new_n13863_), .A2(new_n13861_), .ZN(new_n13935_));
  NOR2_X1    g12915(.A1(new_n13870_), .A2(new_n13868_), .ZN(new_n13936_));
  NOR2_X1    g12916(.A1(new_n13935_), .A2(new_n13936_), .ZN(new_n13937_));
  NOR2_X1    g12917(.A1(new_n13937_), .A2(new_n13871_), .ZN(new_n13938_));
  NAND2_X1   g12918(.A1(new_n13935_), .A2(new_n13936_), .ZN(new_n13939_));
  NAND2_X1   g12919(.A1(new_n13850_), .A2(new_n13855_), .ZN(new_n13940_));
  NOR2_X1    g12920(.A1(new_n13939_), .A2(new_n13940_), .ZN(new_n13941_));
  NAND4_X1   g12921(.A1(new_n13932_), .A2(new_n13934_), .A3(new_n13938_), .A4(new_n13941_), .ZN(new_n13942_));
  NOR2_X1    g12922(.A1(new_n13931_), .A2(new_n13942_), .ZN(new_n13943_));
  AOI21_X1   g12923(.A1(new_n13929_), .A2(new_n13928_), .B(new_n13883_), .ZN(new_n13944_));
  NOR3_X1    g12924(.A1(new_n13924_), .A2(new_n13926_), .A3(new_n13882_), .ZN(new_n13945_));
  NOR3_X1    g12925(.A1(new_n13944_), .A2(new_n13945_), .A3(new_n13921_), .ZN(new_n13946_));
  INV_X1     g12926(.I(new_n13942_), .ZN(new_n13947_));
  NOR2_X1    g12927(.A1(new_n13946_), .A2(new_n13947_), .ZN(new_n13948_));
  OAI21_X1   g12928(.A1(new_n13948_), .A2(new_n13943_), .B(new_n13878_), .ZN(new_n13949_));
  NAND2_X1   g12929(.A1(new_n13931_), .A2(new_n13947_), .ZN(new_n13950_));
  NAND2_X1   g12930(.A1(new_n13927_), .A2(new_n13930_), .ZN(new_n13951_));
  NAND3_X1   g12931(.A1(new_n13934_), .A2(new_n13932_), .A3(new_n13938_), .ZN(new_n13952_));
  NOR3_X1    g12932(.A1(new_n13921_), .A2(new_n13939_), .A3(new_n13940_), .ZN(new_n13953_));
  OAI21_X1   g12933(.A1(new_n13951_), .A2(new_n13952_), .B(new_n13953_), .ZN(new_n13954_));
  NAND3_X1   g12934(.A1(new_n13950_), .A2(new_n13954_), .A3(new_n13878_), .ZN(new_n13955_));
  NAND2_X1   g12935(.A1(new_n13949_), .A2(new_n13955_), .ZN(new_n13956_));
  INV_X1     g12936(.I(new_n13878_), .ZN(new_n13957_));
  NAND2_X1   g12937(.A1(new_n13946_), .A2(new_n13947_), .ZN(new_n13958_));
  NAND2_X1   g12938(.A1(new_n13931_), .A2(new_n13942_), .ZN(new_n13959_));
  AOI21_X1   g12939(.A1(new_n13958_), .A2(new_n13959_), .B(new_n13957_), .ZN(new_n13960_));
  NOR2_X1    g12940(.A1(new_n13946_), .A2(new_n13942_), .ZN(new_n13961_));
  NOR2_X1    g12941(.A1(new_n13944_), .A2(new_n13945_), .ZN(new_n13962_));
  INV_X1     g12942(.I(new_n13952_), .ZN(new_n13963_));
  INV_X1     g12943(.I(new_n13953_), .ZN(new_n13964_));
  AOI21_X1   g12944(.A1(new_n13962_), .A2(new_n13963_), .B(new_n13964_), .ZN(new_n13965_));
  NOR3_X1    g12945(.A1(new_n13965_), .A2(new_n13961_), .A3(new_n13957_), .ZN(new_n13966_));
  NAND2_X1   g12946(.A1(new_n13934_), .A2(new_n13932_), .ZN(new_n13967_));
  NAND2_X1   g12947(.A1(new_n13938_), .A2(new_n13941_), .ZN(new_n13968_));
  XNOR2_X1   g12948(.A1(new_n13967_), .A2(new_n13968_), .ZN(new_n13969_));
  INV_X1     g12949(.I(\A[685] ), .ZN(new_n13970_));
  INV_X1     g12950(.I(\A[686] ), .ZN(new_n13971_));
  NAND2_X1   g12951(.A1(new_n13971_), .A2(\A[687] ), .ZN(new_n13972_));
  INV_X1     g12952(.I(\A[687] ), .ZN(new_n13973_));
  NAND2_X1   g12953(.A1(new_n13973_), .A2(\A[686] ), .ZN(new_n13974_));
  AOI21_X1   g12954(.A1(new_n13972_), .A2(new_n13974_), .B(new_n13970_), .ZN(new_n13975_));
  NOR2_X1    g12955(.A1(\A[686] ), .A2(\A[687] ), .ZN(new_n13976_));
  INV_X1     g12956(.I(new_n13976_), .ZN(new_n13977_));
  NAND2_X1   g12957(.A1(\A[686] ), .A2(\A[687] ), .ZN(new_n13978_));
  AOI21_X1   g12958(.A1(new_n13977_), .A2(new_n13978_), .B(\A[685] ), .ZN(new_n13979_));
  NOR2_X1    g12959(.A1(new_n13979_), .A2(new_n13975_), .ZN(new_n13980_));
  INV_X1     g12960(.I(\A[688] ), .ZN(new_n13981_));
  INV_X1     g12961(.I(\A[689] ), .ZN(new_n13982_));
  NAND2_X1   g12962(.A1(new_n13982_), .A2(\A[690] ), .ZN(new_n13983_));
  INV_X1     g12963(.I(\A[690] ), .ZN(new_n13984_));
  NAND2_X1   g12964(.A1(new_n13984_), .A2(\A[689] ), .ZN(new_n13985_));
  AOI21_X1   g12965(.A1(new_n13983_), .A2(new_n13985_), .B(new_n13981_), .ZN(new_n13986_));
  NOR2_X1    g12966(.A1(\A[689] ), .A2(\A[690] ), .ZN(new_n13987_));
  INV_X1     g12967(.I(new_n13987_), .ZN(new_n13988_));
  NAND2_X1   g12968(.A1(\A[689] ), .A2(\A[690] ), .ZN(new_n13989_));
  AOI21_X1   g12969(.A1(new_n13988_), .A2(new_n13989_), .B(\A[688] ), .ZN(new_n13990_));
  NOR2_X1    g12970(.A1(new_n13990_), .A2(new_n13986_), .ZN(new_n13991_));
  NAND2_X1   g12971(.A1(new_n13980_), .A2(new_n13991_), .ZN(new_n13992_));
  AOI21_X1   g12972(.A1(new_n13981_), .A2(new_n13989_), .B(new_n13987_), .ZN(new_n13993_));
  INV_X1     g12973(.I(new_n13993_), .ZN(new_n13994_));
  AOI21_X1   g12974(.A1(new_n13970_), .A2(new_n13978_), .B(new_n13976_), .ZN(new_n13995_));
  INV_X1     g12975(.I(new_n13995_), .ZN(new_n13996_));
  NOR2_X1    g12976(.A1(new_n13994_), .A2(new_n13996_), .ZN(new_n13997_));
  INV_X1     g12977(.I(new_n13997_), .ZN(new_n13998_));
  NOR2_X1    g12978(.A1(new_n13992_), .A2(new_n13998_), .ZN(new_n13999_));
  NOR2_X1    g12979(.A1(new_n13973_), .A2(\A[686] ), .ZN(new_n14000_));
  NOR2_X1    g12980(.A1(new_n13971_), .A2(\A[687] ), .ZN(new_n14001_));
  OAI21_X1   g12981(.A1(new_n14000_), .A2(new_n14001_), .B(\A[685] ), .ZN(new_n14002_));
  INV_X1     g12982(.I(new_n13978_), .ZN(new_n14003_));
  OAI21_X1   g12983(.A1(new_n14003_), .A2(new_n13976_), .B(new_n13970_), .ZN(new_n14004_));
  NAND2_X1   g12984(.A1(new_n14002_), .A2(new_n14004_), .ZN(new_n14005_));
  NOR2_X1    g12985(.A1(new_n13984_), .A2(\A[689] ), .ZN(new_n14006_));
  NOR2_X1    g12986(.A1(new_n13982_), .A2(\A[690] ), .ZN(new_n14007_));
  OAI21_X1   g12987(.A1(new_n14006_), .A2(new_n14007_), .B(\A[688] ), .ZN(new_n14008_));
  INV_X1     g12988(.I(new_n13989_), .ZN(new_n14009_));
  OAI21_X1   g12989(.A1(new_n14009_), .A2(new_n13987_), .B(new_n13981_), .ZN(new_n14010_));
  NAND2_X1   g12990(.A1(new_n14008_), .A2(new_n14010_), .ZN(new_n14011_));
  NAND2_X1   g12991(.A1(new_n14005_), .A2(new_n14011_), .ZN(new_n14012_));
  NAND3_X1   g12992(.A1(new_n13999_), .A2(new_n13992_), .A3(new_n14012_), .ZN(new_n14013_));
  INV_X1     g12993(.I(\A[679] ), .ZN(new_n14014_));
  INV_X1     g12994(.I(\A[680] ), .ZN(new_n14015_));
  NAND2_X1   g12995(.A1(new_n14015_), .A2(\A[681] ), .ZN(new_n14016_));
  INV_X1     g12996(.I(\A[681] ), .ZN(new_n14017_));
  NAND2_X1   g12997(.A1(new_n14017_), .A2(\A[680] ), .ZN(new_n14018_));
  AOI21_X1   g12998(.A1(new_n14016_), .A2(new_n14018_), .B(new_n14014_), .ZN(new_n14019_));
  NAND2_X1   g12999(.A1(new_n14015_), .A2(new_n14017_), .ZN(new_n14020_));
  NAND2_X1   g13000(.A1(\A[680] ), .A2(\A[681] ), .ZN(new_n14021_));
  AOI21_X1   g13001(.A1(new_n14020_), .A2(new_n14021_), .B(\A[679] ), .ZN(new_n14022_));
  INV_X1     g13002(.I(\A[682] ), .ZN(new_n14023_));
  INV_X1     g13003(.I(\A[683] ), .ZN(new_n14024_));
  NAND2_X1   g13004(.A1(new_n14024_), .A2(\A[684] ), .ZN(new_n14025_));
  INV_X1     g13005(.I(\A[684] ), .ZN(new_n14026_));
  NAND2_X1   g13006(.A1(new_n14026_), .A2(\A[683] ), .ZN(new_n14027_));
  AOI21_X1   g13007(.A1(new_n14025_), .A2(new_n14027_), .B(new_n14023_), .ZN(new_n14028_));
  NAND2_X1   g13008(.A1(new_n14024_), .A2(new_n14026_), .ZN(new_n14029_));
  NAND2_X1   g13009(.A1(\A[683] ), .A2(\A[684] ), .ZN(new_n14030_));
  AOI21_X1   g13010(.A1(new_n14029_), .A2(new_n14030_), .B(\A[682] ), .ZN(new_n14031_));
  NOR4_X1    g13011(.A1(new_n14019_), .A2(new_n14022_), .A3(new_n14031_), .A4(new_n14028_), .ZN(new_n14032_));
  NAND2_X1   g13012(.A1(new_n14030_), .A2(new_n14023_), .ZN(new_n14033_));
  NAND2_X1   g13013(.A1(new_n14033_), .A2(new_n14029_), .ZN(new_n14034_));
  NAND2_X1   g13014(.A1(new_n14021_), .A2(new_n14014_), .ZN(new_n14035_));
  NAND2_X1   g13015(.A1(new_n14035_), .A2(new_n14020_), .ZN(new_n14036_));
  NOR2_X1    g13016(.A1(new_n14034_), .A2(new_n14036_), .ZN(new_n14037_));
  NOR2_X1    g13017(.A1(new_n14022_), .A2(new_n14019_), .ZN(new_n14038_));
  NOR2_X1    g13018(.A1(new_n14031_), .A2(new_n14028_), .ZN(new_n14039_));
  NOR2_X1    g13019(.A1(new_n14038_), .A2(new_n14039_), .ZN(new_n14040_));
  NAND2_X1   g13020(.A1(new_n13969_), .A2(new_n14013_), .ZN(new_n14041_));
  OAI21_X1   g13021(.A1(new_n13966_), .A2(new_n13960_), .B(new_n14041_), .ZN(new_n14042_));
  XOR2_X1    g13022(.A1(new_n13967_), .A2(new_n13968_), .Z(new_n14043_));
  NOR2_X1    g13023(.A1(new_n14005_), .A2(new_n14011_), .ZN(new_n14044_));
  NAND2_X1   g13024(.A1(new_n14044_), .A2(new_n13997_), .ZN(new_n14045_));
  NAND2_X1   g13025(.A1(new_n13992_), .A2(new_n14012_), .ZN(new_n14046_));
  NOR2_X1    g13026(.A1(new_n14046_), .A2(new_n14045_), .ZN(new_n14047_));
  NOR2_X1    g13027(.A1(new_n14043_), .A2(new_n14047_), .ZN(new_n14048_));
  NAND3_X1   g13028(.A1(new_n13949_), .A2(new_n13955_), .A3(new_n14048_), .ZN(new_n14049_));
  NOR2_X1    g13029(.A1(new_n14044_), .A2(new_n13996_), .ZN(new_n14050_));
  NOR2_X1    g13030(.A1(new_n13992_), .A2(new_n13995_), .ZN(new_n14051_));
  OAI21_X1   g13031(.A1(new_n14050_), .A2(new_n14051_), .B(new_n13993_), .ZN(new_n14052_));
  NAND2_X1   g13032(.A1(new_n13992_), .A2(new_n13995_), .ZN(new_n14053_));
  NAND2_X1   g13033(.A1(new_n14044_), .A2(new_n13996_), .ZN(new_n14054_));
  NAND3_X1   g13034(.A1(new_n14054_), .A2(new_n14053_), .A3(new_n13994_), .ZN(new_n14055_));
  NAND2_X1   g13035(.A1(new_n14052_), .A2(new_n14055_), .ZN(new_n14056_));
  NOR2_X1    g13036(.A1(new_n14046_), .A2(new_n14045_), .ZN(new_n14057_));
  NOR2_X1    g13037(.A1(new_n14040_), .A2(new_n14032_), .ZN(new_n14058_));
  NAND2_X1   g13038(.A1(new_n14057_), .A2(new_n14058_), .ZN(new_n14059_));
  NAND2_X1   g13039(.A1(new_n14032_), .A2(new_n14037_), .ZN(new_n14060_));
  NAND2_X1   g13040(.A1(new_n13980_), .A2(new_n14011_), .ZN(new_n14061_));
  NAND2_X1   g13041(.A1(new_n13991_), .A2(new_n14005_), .ZN(new_n14062_));
  AOI21_X1   g13042(.A1(new_n14061_), .A2(new_n14062_), .B(new_n13998_), .ZN(new_n14063_));
  NOR2_X1    g13043(.A1(new_n14063_), .A2(new_n14060_), .ZN(new_n14064_));
  OAI21_X1   g13044(.A1(new_n14056_), .A2(new_n14059_), .B(new_n14064_), .ZN(new_n14065_));
  INV_X1     g13045(.I(new_n14034_), .ZN(new_n14066_));
  NOR2_X1    g13046(.A1(new_n14032_), .A2(new_n14036_), .ZN(new_n14067_));
  NAND2_X1   g13047(.A1(new_n14032_), .A2(new_n14036_), .ZN(new_n14068_));
  INV_X1     g13048(.I(new_n14068_), .ZN(new_n14069_));
  OAI21_X1   g13049(.A1(new_n14069_), .A2(new_n14067_), .B(new_n14066_), .ZN(new_n14070_));
  INV_X1     g13050(.I(new_n14067_), .ZN(new_n14071_));
  NAND3_X1   g13051(.A1(new_n14071_), .A2(new_n14034_), .A3(new_n14068_), .ZN(new_n14072_));
  AND2_X2    g13052(.A1(new_n14070_), .A2(new_n14072_), .Z(new_n14073_));
  NOR2_X1    g13053(.A1(new_n14065_), .A2(new_n14073_), .ZN(new_n14074_));
  INV_X1     g13054(.I(new_n14074_), .ZN(new_n14075_));
  NAND2_X1   g13055(.A1(new_n14070_), .A2(new_n14072_), .ZN(new_n14076_));
  INV_X1     g13056(.I(new_n14058_), .ZN(new_n14077_));
  NOR2_X1    g13057(.A1(new_n14077_), .A2(new_n14060_), .ZN(new_n14078_));
  NAND2_X1   g13058(.A1(new_n14078_), .A2(new_n14057_), .ZN(new_n14079_));
  NAND2_X1   g13059(.A1(new_n14079_), .A2(new_n14076_), .ZN(new_n14080_));
  NOR3_X1    g13060(.A1(new_n14013_), .A2(new_n14060_), .A3(new_n14077_), .ZN(new_n14081_));
  AOI21_X1   g13061(.A1(new_n14054_), .A2(new_n14053_), .B(new_n13994_), .ZN(new_n14082_));
  NOR3_X1    g13062(.A1(new_n14050_), .A2(new_n14051_), .A3(new_n13993_), .ZN(new_n14083_));
  NOR3_X1    g13063(.A1(new_n14082_), .A2(new_n14083_), .A3(new_n14063_), .ZN(new_n14084_));
  AOI21_X1   g13064(.A1(new_n14073_), .A2(new_n14081_), .B(new_n14084_), .ZN(new_n14085_));
  NOR4_X1    g13065(.A1(new_n14079_), .A2(new_n14056_), .A3(new_n14076_), .A4(new_n14063_), .ZN(new_n14086_));
  OAI21_X1   g13066(.A1(new_n14085_), .A2(new_n14086_), .B(new_n14080_), .ZN(new_n14087_));
  NAND2_X1   g13067(.A1(new_n14087_), .A2(new_n14075_), .ZN(new_n14088_));
  AOI22_X1   g13068(.A1(new_n14088_), .A2(new_n13956_), .B1(new_n14042_), .B2(new_n14049_), .ZN(new_n14089_));
  NOR2_X1    g13069(.A1(new_n13961_), .A2(new_n13878_), .ZN(new_n14090_));
  NOR2_X1    g13070(.A1(new_n13882_), .A2(new_n13887_), .ZN(new_n14091_));
  OAI21_X1   g13071(.A1(new_n13925_), .A2(new_n14091_), .B(new_n13890_), .ZN(new_n14092_));
  NOR2_X1    g13072(.A1(new_n13850_), .A2(new_n13855_), .ZN(new_n14093_));
  OAI21_X1   g13073(.A1(new_n13939_), .A2(new_n14093_), .B(new_n13940_), .ZN(new_n14094_));
  XNOR2_X1   g13074(.A1(new_n14092_), .A2(new_n14094_), .ZN(new_n14095_));
  INV_X1     g13075(.I(new_n14095_), .ZN(new_n14096_));
  NOR3_X1    g13076(.A1(new_n14090_), .A2(new_n13965_), .A3(new_n14096_), .ZN(new_n14097_));
  OAI21_X1   g13077(.A1(new_n14079_), .A2(new_n14084_), .B(new_n14076_), .ZN(new_n14098_));
  NOR2_X1    g13078(.A1(new_n13993_), .A2(new_n13995_), .ZN(new_n14099_));
  OAI21_X1   g13079(.A1(new_n13992_), .A2(new_n14099_), .B(new_n13998_), .ZN(new_n14100_));
  INV_X1     g13080(.I(new_n14032_), .ZN(new_n14101_));
  INV_X1     g13081(.I(new_n14037_), .ZN(new_n14102_));
  AOI21_X1   g13082(.A1(new_n14020_), .A2(new_n14035_), .B(new_n14066_), .ZN(new_n14103_));
  OAI21_X1   g13083(.A1(new_n14101_), .A2(new_n14103_), .B(new_n14102_), .ZN(new_n14104_));
  XNOR2_X1   g13084(.A1(new_n14104_), .A2(new_n14100_), .ZN(new_n14105_));
  NAND3_X1   g13085(.A1(new_n14098_), .A2(new_n14065_), .A3(new_n14105_), .ZN(new_n14106_));
  INV_X1     g13086(.I(new_n14106_), .ZN(new_n14107_));
  NAND3_X1   g13087(.A1(new_n14089_), .A2(new_n14097_), .A3(new_n14107_), .ZN(new_n14108_));
  NAND2_X1   g13088(.A1(new_n14104_), .A2(new_n14100_), .ZN(new_n14109_));
  OR2_X2     g13089(.A1(new_n14104_), .A2(new_n14100_), .Z(new_n14110_));
  NAND3_X1   g13090(.A1(new_n14098_), .A2(new_n14065_), .A3(new_n14110_), .ZN(new_n14111_));
  NAND2_X1   g13091(.A1(new_n14111_), .A2(new_n14109_), .ZN(new_n14112_));
  NAND2_X1   g13092(.A1(new_n14092_), .A2(new_n14094_), .ZN(new_n14113_));
  NOR2_X1    g13093(.A1(new_n14090_), .A2(new_n13965_), .ZN(new_n14114_));
  OAI21_X1   g13094(.A1(new_n14092_), .A2(new_n14094_), .B(new_n14114_), .ZN(new_n14115_));
  NAND2_X1   g13095(.A1(new_n14115_), .A2(new_n14113_), .ZN(new_n14116_));
  OAI21_X1   g13096(.A1(new_n14112_), .A2(new_n14116_), .B(new_n14108_), .ZN(new_n14117_));
  NAND2_X1   g13097(.A1(new_n14116_), .A2(new_n14112_), .ZN(new_n14118_));
  NAND2_X1   g13098(.A1(new_n14117_), .A2(new_n14118_), .ZN(new_n14119_));
  INV_X1     g13099(.I(\A[670] ), .ZN(new_n14120_));
  NOR2_X1    g13100(.A1(\A[671] ), .A2(\A[672] ), .ZN(new_n14121_));
  NAND2_X1   g13101(.A1(\A[671] ), .A2(\A[672] ), .ZN(new_n14122_));
  AOI21_X1   g13102(.A1(new_n14120_), .A2(new_n14122_), .B(new_n14121_), .ZN(new_n14123_));
  INV_X1     g13103(.I(new_n14123_), .ZN(new_n14124_));
  INV_X1     g13104(.I(\A[667] ), .ZN(new_n14125_));
  NOR2_X1    g13105(.A1(\A[668] ), .A2(\A[669] ), .ZN(new_n14126_));
  NAND2_X1   g13106(.A1(\A[668] ), .A2(\A[669] ), .ZN(new_n14127_));
  AOI21_X1   g13107(.A1(new_n14125_), .A2(new_n14127_), .B(new_n14126_), .ZN(new_n14128_));
  INV_X1     g13108(.I(new_n14128_), .ZN(new_n14129_));
  INV_X1     g13109(.I(\A[668] ), .ZN(new_n14130_));
  NAND2_X1   g13110(.A1(new_n14130_), .A2(\A[669] ), .ZN(new_n14131_));
  INV_X1     g13111(.I(\A[669] ), .ZN(new_n14132_));
  NAND2_X1   g13112(.A1(new_n14132_), .A2(\A[668] ), .ZN(new_n14133_));
  AOI21_X1   g13113(.A1(new_n14131_), .A2(new_n14133_), .B(new_n14125_), .ZN(new_n14134_));
  INV_X1     g13114(.I(new_n14126_), .ZN(new_n14135_));
  AOI21_X1   g13115(.A1(new_n14135_), .A2(new_n14127_), .B(\A[667] ), .ZN(new_n14136_));
  INV_X1     g13116(.I(\A[671] ), .ZN(new_n14137_));
  NAND2_X1   g13117(.A1(new_n14137_), .A2(\A[672] ), .ZN(new_n14138_));
  INV_X1     g13118(.I(\A[672] ), .ZN(new_n14139_));
  NAND2_X1   g13119(.A1(new_n14139_), .A2(\A[671] ), .ZN(new_n14140_));
  AOI21_X1   g13120(.A1(new_n14138_), .A2(new_n14140_), .B(new_n14120_), .ZN(new_n14141_));
  INV_X1     g13121(.I(new_n14121_), .ZN(new_n14142_));
  AOI21_X1   g13122(.A1(new_n14142_), .A2(new_n14122_), .B(\A[670] ), .ZN(new_n14143_));
  NOR4_X1    g13123(.A1(new_n14134_), .A2(new_n14136_), .A3(new_n14143_), .A4(new_n14141_), .ZN(new_n14144_));
  NOR2_X1    g13124(.A1(new_n14144_), .A2(new_n14129_), .ZN(new_n14145_));
  INV_X1     g13125(.I(new_n14145_), .ZN(new_n14146_));
  NAND2_X1   g13126(.A1(new_n14144_), .A2(new_n14129_), .ZN(new_n14147_));
  AOI21_X1   g13127(.A1(new_n14146_), .A2(new_n14147_), .B(new_n14124_), .ZN(new_n14148_));
  AND3_X2    g13128(.A1(new_n14146_), .A2(new_n14124_), .A3(new_n14147_), .Z(new_n14149_));
  NOR2_X1    g13129(.A1(new_n14149_), .A2(new_n14148_), .ZN(new_n14150_));
  INV_X1     g13130(.I(\A[676] ), .ZN(new_n14151_));
  NOR2_X1    g13131(.A1(\A[677] ), .A2(\A[678] ), .ZN(new_n14152_));
  NAND2_X1   g13132(.A1(\A[677] ), .A2(\A[678] ), .ZN(new_n14153_));
  AOI21_X1   g13133(.A1(new_n14151_), .A2(new_n14153_), .B(new_n14152_), .ZN(new_n14154_));
  INV_X1     g13134(.I(new_n14154_), .ZN(new_n14155_));
  INV_X1     g13135(.I(\A[673] ), .ZN(new_n14156_));
  NOR2_X1    g13136(.A1(\A[674] ), .A2(\A[675] ), .ZN(new_n14157_));
  NAND2_X1   g13137(.A1(\A[674] ), .A2(\A[675] ), .ZN(new_n14158_));
  AOI21_X1   g13138(.A1(new_n14156_), .A2(new_n14158_), .B(new_n14157_), .ZN(new_n14159_));
  INV_X1     g13139(.I(new_n14159_), .ZN(new_n14160_));
  NOR2_X1    g13140(.A1(new_n14155_), .A2(new_n14160_), .ZN(new_n14161_));
  INV_X1     g13141(.I(\A[674] ), .ZN(new_n14162_));
  NAND2_X1   g13142(.A1(new_n14162_), .A2(\A[675] ), .ZN(new_n14163_));
  INV_X1     g13143(.I(\A[675] ), .ZN(new_n14164_));
  NAND2_X1   g13144(.A1(new_n14164_), .A2(\A[674] ), .ZN(new_n14165_));
  AOI21_X1   g13145(.A1(new_n14163_), .A2(new_n14165_), .B(new_n14156_), .ZN(new_n14166_));
  INV_X1     g13146(.I(new_n14157_), .ZN(new_n14167_));
  AOI21_X1   g13147(.A1(new_n14167_), .A2(new_n14158_), .B(\A[673] ), .ZN(new_n14168_));
  NOR2_X1    g13148(.A1(new_n14168_), .A2(new_n14166_), .ZN(new_n14169_));
  INV_X1     g13149(.I(\A[678] ), .ZN(new_n14170_));
  NOR2_X1    g13150(.A1(new_n14170_), .A2(\A[677] ), .ZN(new_n14171_));
  INV_X1     g13151(.I(\A[677] ), .ZN(new_n14172_));
  NOR2_X1    g13152(.A1(new_n14172_), .A2(\A[678] ), .ZN(new_n14173_));
  OAI21_X1   g13153(.A1(new_n14171_), .A2(new_n14173_), .B(\A[676] ), .ZN(new_n14174_));
  INV_X1     g13154(.I(new_n14153_), .ZN(new_n14175_));
  OAI21_X1   g13155(.A1(new_n14175_), .A2(new_n14152_), .B(new_n14151_), .ZN(new_n14176_));
  NAND2_X1   g13156(.A1(new_n14174_), .A2(new_n14176_), .ZN(new_n14177_));
  NAND2_X1   g13157(.A1(new_n14169_), .A2(new_n14177_), .ZN(new_n14178_));
  NOR2_X1    g13158(.A1(new_n14164_), .A2(\A[674] ), .ZN(new_n14179_));
  NOR2_X1    g13159(.A1(new_n14162_), .A2(\A[675] ), .ZN(new_n14180_));
  OAI21_X1   g13160(.A1(new_n14179_), .A2(new_n14180_), .B(\A[673] ), .ZN(new_n14181_));
  INV_X1     g13161(.I(new_n14158_), .ZN(new_n14182_));
  OAI21_X1   g13162(.A1(new_n14182_), .A2(new_n14157_), .B(new_n14156_), .ZN(new_n14183_));
  NAND2_X1   g13163(.A1(new_n14181_), .A2(new_n14183_), .ZN(new_n14184_));
  NAND2_X1   g13164(.A1(new_n14172_), .A2(\A[678] ), .ZN(new_n14185_));
  NAND2_X1   g13165(.A1(new_n14170_), .A2(\A[677] ), .ZN(new_n14186_));
  AOI21_X1   g13166(.A1(new_n14185_), .A2(new_n14186_), .B(new_n14151_), .ZN(new_n14187_));
  INV_X1     g13167(.I(new_n14152_), .ZN(new_n14188_));
  AOI21_X1   g13168(.A1(new_n14188_), .A2(new_n14153_), .B(\A[676] ), .ZN(new_n14189_));
  NOR2_X1    g13169(.A1(new_n14189_), .A2(new_n14187_), .ZN(new_n14190_));
  NAND2_X1   g13170(.A1(new_n14190_), .A2(new_n14184_), .ZN(new_n14191_));
  NAND2_X1   g13171(.A1(new_n14178_), .A2(new_n14191_), .ZN(new_n14192_));
  NAND2_X1   g13172(.A1(new_n14192_), .A2(new_n14161_), .ZN(new_n14193_));
  NOR2_X1    g13173(.A1(new_n14184_), .A2(new_n14177_), .ZN(new_n14194_));
  NOR2_X1    g13174(.A1(new_n14194_), .A2(new_n14160_), .ZN(new_n14195_));
  NAND2_X1   g13175(.A1(new_n14169_), .A2(new_n14190_), .ZN(new_n14196_));
  NOR2_X1    g13176(.A1(new_n14196_), .A2(new_n14159_), .ZN(new_n14197_));
  OAI21_X1   g13177(.A1(new_n14195_), .A2(new_n14197_), .B(new_n14154_), .ZN(new_n14198_));
  NAND2_X1   g13178(.A1(new_n14196_), .A2(new_n14159_), .ZN(new_n14199_));
  NAND2_X1   g13179(.A1(new_n14194_), .A2(new_n14160_), .ZN(new_n14200_));
  NAND3_X1   g13180(.A1(new_n14200_), .A2(new_n14199_), .A3(new_n14155_), .ZN(new_n14201_));
  NAND3_X1   g13181(.A1(new_n14198_), .A2(new_n14201_), .A3(new_n14193_), .ZN(new_n14202_));
  INV_X1     g13182(.I(new_n14161_), .ZN(new_n14203_));
  NOR2_X1    g13183(.A1(new_n14196_), .A2(new_n14203_), .ZN(new_n14204_));
  NOR2_X1    g13184(.A1(new_n14169_), .A2(new_n14190_), .ZN(new_n14205_));
  NOR2_X1    g13185(.A1(new_n14205_), .A2(new_n14194_), .ZN(new_n14206_));
  NOR2_X1    g13186(.A1(new_n14136_), .A2(new_n14134_), .ZN(new_n14207_));
  NOR2_X1    g13187(.A1(new_n14143_), .A2(new_n14141_), .ZN(new_n14208_));
  NOR2_X1    g13188(.A1(new_n14207_), .A2(new_n14208_), .ZN(new_n14209_));
  NOR2_X1    g13189(.A1(new_n14209_), .A2(new_n14144_), .ZN(new_n14210_));
  INV_X1     g13190(.I(new_n14144_), .ZN(new_n14211_));
  NAND2_X1   g13191(.A1(new_n14123_), .A2(new_n14128_), .ZN(new_n14212_));
  NOR2_X1    g13192(.A1(new_n14211_), .A2(new_n14212_), .ZN(new_n14213_));
  NAND4_X1   g13193(.A1(new_n14206_), .A2(new_n14213_), .A3(new_n14204_), .A4(new_n14210_), .ZN(new_n14214_));
  NOR2_X1    g13194(.A1(new_n14202_), .A2(new_n14214_), .ZN(new_n14215_));
  AOI21_X1   g13195(.A1(new_n14178_), .A2(new_n14191_), .B(new_n14203_), .ZN(new_n14216_));
  AOI21_X1   g13196(.A1(new_n14200_), .A2(new_n14199_), .B(new_n14155_), .ZN(new_n14217_));
  NOR3_X1    g13197(.A1(new_n14195_), .A2(new_n14197_), .A3(new_n14154_), .ZN(new_n14218_));
  NOR3_X1    g13198(.A1(new_n14217_), .A2(new_n14218_), .A3(new_n14216_), .ZN(new_n14219_));
  INV_X1     g13199(.I(new_n14214_), .ZN(new_n14220_));
  NOR2_X1    g13200(.A1(new_n14219_), .A2(new_n14220_), .ZN(new_n14221_));
  OAI21_X1   g13201(.A1(new_n14221_), .A2(new_n14215_), .B(new_n14150_), .ZN(new_n14222_));
  NAND2_X1   g13202(.A1(new_n14202_), .A2(new_n14220_), .ZN(new_n14223_));
  NAND2_X1   g13203(.A1(new_n14198_), .A2(new_n14201_), .ZN(new_n14224_));
  NAND3_X1   g13204(.A1(new_n14206_), .A2(new_n14204_), .A3(new_n14210_), .ZN(new_n14225_));
  NOR3_X1    g13205(.A1(new_n14216_), .A2(new_n14211_), .A3(new_n14212_), .ZN(new_n14226_));
  OAI21_X1   g13206(.A1(new_n14224_), .A2(new_n14225_), .B(new_n14226_), .ZN(new_n14227_));
  NAND3_X1   g13207(.A1(new_n14223_), .A2(new_n14227_), .A3(new_n14150_), .ZN(new_n14228_));
  NAND2_X1   g13208(.A1(new_n14222_), .A2(new_n14228_), .ZN(new_n14229_));
  INV_X1     g13209(.I(new_n14229_), .ZN(new_n14230_));
  NAND2_X1   g13210(.A1(new_n14206_), .A2(new_n14204_), .ZN(new_n14231_));
  NAND2_X1   g13211(.A1(new_n14213_), .A2(new_n14210_), .ZN(new_n14232_));
  XOR2_X1    g13212(.A1(new_n14231_), .A2(new_n14232_), .Z(new_n14233_));
  INV_X1     g13213(.I(\A[663] ), .ZN(new_n14234_));
  NOR2_X1    g13214(.A1(new_n14234_), .A2(\A[662] ), .ZN(new_n14235_));
  INV_X1     g13215(.I(\A[662] ), .ZN(new_n14236_));
  NOR2_X1    g13216(.A1(new_n14236_), .A2(\A[663] ), .ZN(new_n14237_));
  OAI21_X1   g13217(.A1(new_n14235_), .A2(new_n14237_), .B(\A[661] ), .ZN(new_n14238_));
  INV_X1     g13218(.I(\A[661] ), .ZN(new_n14239_));
  NOR2_X1    g13219(.A1(\A[662] ), .A2(\A[663] ), .ZN(new_n14240_));
  NAND2_X1   g13220(.A1(\A[662] ), .A2(\A[663] ), .ZN(new_n14241_));
  INV_X1     g13221(.I(new_n14241_), .ZN(new_n14242_));
  OAI21_X1   g13222(.A1(new_n14242_), .A2(new_n14240_), .B(new_n14239_), .ZN(new_n14243_));
  NAND2_X1   g13223(.A1(new_n14238_), .A2(new_n14243_), .ZN(new_n14244_));
  INV_X1     g13224(.I(\A[666] ), .ZN(new_n14245_));
  NOR2_X1    g13225(.A1(new_n14245_), .A2(\A[665] ), .ZN(new_n14246_));
  INV_X1     g13226(.I(\A[665] ), .ZN(new_n14247_));
  NOR2_X1    g13227(.A1(new_n14247_), .A2(\A[666] ), .ZN(new_n14248_));
  OAI21_X1   g13228(.A1(new_n14246_), .A2(new_n14248_), .B(\A[664] ), .ZN(new_n14249_));
  INV_X1     g13229(.I(\A[664] ), .ZN(new_n14250_));
  NOR2_X1    g13230(.A1(\A[665] ), .A2(\A[666] ), .ZN(new_n14251_));
  NAND2_X1   g13231(.A1(\A[665] ), .A2(\A[666] ), .ZN(new_n14252_));
  INV_X1     g13232(.I(new_n14252_), .ZN(new_n14253_));
  OAI21_X1   g13233(.A1(new_n14253_), .A2(new_n14251_), .B(new_n14250_), .ZN(new_n14254_));
  NAND2_X1   g13234(.A1(new_n14249_), .A2(new_n14254_), .ZN(new_n14255_));
  NOR2_X1    g13235(.A1(new_n14244_), .A2(new_n14255_), .ZN(new_n14256_));
  AOI21_X1   g13236(.A1(new_n14250_), .A2(new_n14252_), .B(new_n14251_), .ZN(new_n14257_));
  INV_X1     g13237(.I(new_n14257_), .ZN(new_n14258_));
  AOI21_X1   g13238(.A1(new_n14239_), .A2(new_n14241_), .B(new_n14240_), .ZN(new_n14259_));
  INV_X1     g13239(.I(new_n14259_), .ZN(new_n14260_));
  NOR2_X1    g13240(.A1(new_n14258_), .A2(new_n14260_), .ZN(new_n14261_));
  NAND2_X1   g13241(.A1(new_n14256_), .A2(new_n14261_), .ZN(new_n14262_));
  NAND2_X1   g13242(.A1(new_n14236_), .A2(\A[663] ), .ZN(new_n14263_));
  NAND2_X1   g13243(.A1(new_n14234_), .A2(\A[662] ), .ZN(new_n14264_));
  AOI21_X1   g13244(.A1(new_n14263_), .A2(new_n14264_), .B(new_n14239_), .ZN(new_n14265_));
  INV_X1     g13245(.I(new_n14240_), .ZN(new_n14266_));
  AOI21_X1   g13246(.A1(new_n14266_), .A2(new_n14241_), .B(\A[661] ), .ZN(new_n14267_));
  NOR2_X1    g13247(.A1(new_n14267_), .A2(new_n14265_), .ZN(new_n14268_));
  NAND2_X1   g13248(.A1(new_n14247_), .A2(\A[666] ), .ZN(new_n14269_));
  NAND2_X1   g13249(.A1(new_n14245_), .A2(\A[665] ), .ZN(new_n14270_));
  AOI21_X1   g13250(.A1(new_n14269_), .A2(new_n14270_), .B(new_n14250_), .ZN(new_n14271_));
  INV_X1     g13251(.I(new_n14251_), .ZN(new_n14272_));
  AOI21_X1   g13252(.A1(new_n14272_), .A2(new_n14252_), .B(\A[664] ), .ZN(new_n14273_));
  NOR2_X1    g13253(.A1(new_n14273_), .A2(new_n14271_), .ZN(new_n14274_));
  NAND2_X1   g13254(.A1(new_n14268_), .A2(new_n14274_), .ZN(new_n14275_));
  NAND2_X1   g13255(.A1(new_n14244_), .A2(new_n14255_), .ZN(new_n14276_));
  NAND2_X1   g13256(.A1(new_n14275_), .A2(new_n14276_), .ZN(new_n14277_));
  INV_X1     g13257(.I(\A[655] ), .ZN(new_n14278_));
  INV_X1     g13258(.I(\A[656] ), .ZN(new_n14279_));
  NAND2_X1   g13259(.A1(new_n14279_), .A2(\A[657] ), .ZN(new_n14280_));
  INV_X1     g13260(.I(\A[657] ), .ZN(new_n14281_));
  NAND2_X1   g13261(.A1(new_n14281_), .A2(\A[656] ), .ZN(new_n14282_));
  AOI21_X1   g13262(.A1(new_n14280_), .A2(new_n14282_), .B(new_n14278_), .ZN(new_n14283_));
  NAND2_X1   g13263(.A1(new_n14279_), .A2(new_n14281_), .ZN(new_n14284_));
  NAND2_X1   g13264(.A1(\A[656] ), .A2(\A[657] ), .ZN(new_n14285_));
  AOI21_X1   g13265(.A1(new_n14284_), .A2(new_n14285_), .B(\A[655] ), .ZN(new_n14286_));
  NOR2_X1    g13266(.A1(new_n14286_), .A2(new_n14283_), .ZN(new_n14287_));
  INV_X1     g13267(.I(\A[658] ), .ZN(new_n14288_));
  INV_X1     g13268(.I(\A[659] ), .ZN(new_n14289_));
  NAND2_X1   g13269(.A1(new_n14289_), .A2(\A[660] ), .ZN(new_n14290_));
  INV_X1     g13270(.I(\A[660] ), .ZN(new_n14291_));
  NAND2_X1   g13271(.A1(new_n14291_), .A2(\A[659] ), .ZN(new_n14292_));
  AOI21_X1   g13272(.A1(new_n14290_), .A2(new_n14292_), .B(new_n14288_), .ZN(new_n14293_));
  NAND2_X1   g13273(.A1(new_n14289_), .A2(new_n14291_), .ZN(new_n14294_));
  NAND2_X1   g13274(.A1(\A[659] ), .A2(\A[660] ), .ZN(new_n14295_));
  AOI21_X1   g13275(.A1(new_n14294_), .A2(new_n14295_), .B(\A[658] ), .ZN(new_n14296_));
  NOR2_X1    g13276(.A1(new_n14296_), .A2(new_n14293_), .ZN(new_n14297_));
  NAND2_X1   g13277(.A1(new_n14295_), .A2(new_n14288_), .ZN(new_n14298_));
  NAND2_X1   g13278(.A1(new_n14298_), .A2(new_n14294_), .ZN(new_n14299_));
  NAND2_X1   g13279(.A1(new_n14285_), .A2(new_n14278_), .ZN(new_n14300_));
  NAND2_X1   g13280(.A1(new_n14300_), .A2(new_n14284_), .ZN(new_n14301_));
  NOR2_X1    g13281(.A1(new_n14299_), .A2(new_n14301_), .ZN(new_n14302_));
  NOR2_X1    g13282(.A1(new_n14277_), .A2(new_n14262_), .ZN(new_n14303_));
  NOR2_X1    g13283(.A1(new_n14233_), .A2(new_n14303_), .ZN(new_n14304_));
  AOI21_X1   g13284(.A1(new_n14222_), .A2(new_n14228_), .B(new_n14304_), .ZN(new_n14305_));
  AND3_X2    g13285(.A1(new_n14222_), .A2(new_n14228_), .A3(new_n14304_), .Z(new_n14306_));
  NOR2_X1    g13286(.A1(new_n14256_), .A2(new_n14260_), .ZN(new_n14307_));
  NOR2_X1    g13287(.A1(new_n14275_), .A2(new_n14259_), .ZN(new_n14308_));
  OAI21_X1   g13288(.A1(new_n14307_), .A2(new_n14308_), .B(new_n14257_), .ZN(new_n14309_));
  NAND2_X1   g13289(.A1(new_n14275_), .A2(new_n14259_), .ZN(new_n14310_));
  NAND2_X1   g13290(.A1(new_n14256_), .A2(new_n14260_), .ZN(new_n14311_));
  NAND3_X1   g13291(.A1(new_n14311_), .A2(new_n14310_), .A3(new_n14258_), .ZN(new_n14312_));
  NAND2_X1   g13292(.A1(new_n14309_), .A2(new_n14312_), .ZN(new_n14313_));
  NOR2_X1    g13293(.A1(new_n14277_), .A2(new_n14262_), .ZN(new_n14314_));
  NOR4_X1    g13294(.A1(new_n14283_), .A2(new_n14286_), .A3(new_n14296_), .A4(new_n14293_), .ZN(new_n14315_));
  NOR2_X1    g13295(.A1(new_n14287_), .A2(new_n14297_), .ZN(new_n14316_));
  NOR2_X1    g13296(.A1(new_n14316_), .A2(new_n14315_), .ZN(new_n14317_));
  NAND2_X1   g13297(.A1(new_n14314_), .A2(new_n14317_), .ZN(new_n14318_));
  NAND2_X1   g13298(.A1(new_n14315_), .A2(new_n14302_), .ZN(new_n14319_));
  INV_X1     g13299(.I(new_n14261_), .ZN(new_n14320_));
  NAND2_X1   g13300(.A1(new_n14268_), .A2(new_n14255_), .ZN(new_n14321_));
  NAND2_X1   g13301(.A1(new_n14274_), .A2(new_n14244_), .ZN(new_n14322_));
  AOI21_X1   g13302(.A1(new_n14321_), .A2(new_n14322_), .B(new_n14320_), .ZN(new_n14323_));
  NOR2_X1    g13303(.A1(new_n14323_), .A2(new_n14319_), .ZN(new_n14324_));
  OAI21_X1   g13304(.A1(new_n14313_), .A2(new_n14318_), .B(new_n14324_), .ZN(new_n14325_));
  INV_X1     g13305(.I(new_n14325_), .ZN(new_n14326_));
  INV_X1     g13306(.I(new_n14299_), .ZN(new_n14327_));
  NOR2_X1    g13307(.A1(new_n14315_), .A2(new_n14301_), .ZN(new_n14328_));
  NAND2_X1   g13308(.A1(new_n14315_), .A2(new_n14301_), .ZN(new_n14329_));
  INV_X1     g13309(.I(new_n14329_), .ZN(new_n14330_));
  OAI21_X1   g13310(.A1(new_n14330_), .A2(new_n14328_), .B(new_n14327_), .ZN(new_n14331_));
  INV_X1     g13311(.I(new_n14328_), .ZN(new_n14332_));
  NAND3_X1   g13312(.A1(new_n14332_), .A2(new_n14299_), .A3(new_n14329_), .ZN(new_n14333_));
  NAND2_X1   g13313(.A1(new_n14331_), .A2(new_n14333_), .ZN(new_n14334_));
  OR2_X2     g13314(.A1(new_n14316_), .A2(new_n14315_), .Z(new_n14335_));
  NOR2_X1    g13315(.A1(new_n14335_), .A2(new_n14319_), .ZN(new_n14336_));
  NAND2_X1   g13316(.A1(new_n14336_), .A2(new_n14314_), .ZN(new_n14337_));
  NAND2_X1   g13317(.A1(new_n14337_), .A2(new_n14334_), .ZN(new_n14338_));
  AOI21_X1   g13318(.A1(new_n14311_), .A2(new_n14310_), .B(new_n14258_), .ZN(new_n14339_));
  NOR3_X1    g13319(.A1(new_n14307_), .A2(new_n14308_), .A3(new_n14257_), .ZN(new_n14340_));
  NOR3_X1    g13320(.A1(new_n14339_), .A2(new_n14340_), .A3(new_n14323_), .ZN(new_n14341_));
  NAND4_X1   g13321(.A1(new_n14336_), .A2(new_n14331_), .A3(new_n14333_), .A4(new_n14314_), .ZN(new_n14342_));
  XOR2_X1    g13322(.A1(new_n14342_), .A2(new_n14341_), .Z(new_n14343_));
  AOI22_X1   g13323(.A1(new_n14343_), .A2(new_n14338_), .B1(new_n14326_), .B2(new_n14334_), .ZN(new_n14344_));
  OAI22_X1   g13324(.A1(new_n14344_), .A2(new_n14230_), .B1(new_n14306_), .B2(new_n14305_), .ZN(new_n14345_));
  OAI22_X1   g13325(.A1(new_n14219_), .A2(new_n14214_), .B1(new_n14148_), .B2(new_n14149_), .ZN(new_n14346_));
  NOR2_X1    g13326(.A1(new_n14154_), .A2(new_n14159_), .ZN(new_n14347_));
  OAI21_X1   g13327(.A1(new_n14196_), .A2(new_n14347_), .B(new_n14203_), .ZN(new_n14348_));
  NOR2_X1    g13328(.A1(new_n14123_), .A2(new_n14128_), .ZN(new_n14349_));
  OAI21_X1   g13329(.A1(new_n14211_), .A2(new_n14349_), .B(new_n14212_), .ZN(new_n14350_));
  XNOR2_X1   g13330(.A1(new_n14350_), .A2(new_n14348_), .ZN(new_n14351_));
  NAND3_X1   g13331(.A1(new_n14346_), .A2(new_n14227_), .A3(new_n14351_), .ZN(new_n14352_));
  OAI21_X1   g13332(.A1(new_n14337_), .A2(new_n14341_), .B(new_n14334_), .ZN(new_n14353_));
  NOR2_X1    g13333(.A1(new_n14257_), .A2(new_n14259_), .ZN(new_n14354_));
  OAI21_X1   g13334(.A1(new_n14275_), .A2(new_n14354_), .B(new_n14320_), .ZN(new_n14355_));
  INV_X1     g13335(.I(new_n14315_), .ZN(new_n14356_));
  INV_X1     g13336(.I(new_n14302_), .ZN(new_n14357_));
  AOI21_X1   g13337(.A1(new_n14284_), .A2(new_n14300_), .B(new_n14327_), .ZN(new_n14358_));
  OAI21_X1   g13338(.A1(new_n14356_), .A2(new_n14358_), .B(new_n14357_), .ZN(new_n14359_));
  XNOR2_X1   g13339(.A1(new_n14359_), .A2(new_n14355_), .ZN(new_n14360_));
  NAND3_X1   g13340(.A1(new_n14353_), .A2(new_n14325_), .A3(new_n14360_), .ZN(new_n14361_));
  NAND2_X1   g13341(.A1(new_n14352_), .A2(new_n14361_), .ZN(new_n14362_));
  NOR2_X1    g13342(.A1(new_n14352_), .A2(new_n14361_), .ZN(new_n14363_));
  INV_X1     g13343(.I(new_n14363_), .ZN(new_n14364_));
  AOI21_X1   g13344(.A1(new_n14345_), .A2(new_n14362_), .B(new_n14364_), .ZN(new_n14365_));
  NAND2_X1   g13345(.A1(new_n14359_), .A2(new_n14355_), .ZN(new_n14366_));
  OR2_X2     g13346(.A1(new_n14359_), .A2(new_n14355_), .Z(new_n14367_));
  NAND3_X1   g13347(.A1(new_n14353_), .A2(new_n14325_), .A3(new_n14367_), .ZN(new_n14368_));
  NAND2_X1   g13348(.A1(new_n14368_), .A2(new_n14366_), .ZN(new_n14369_));
  INV_X1     g13349(.I(new_n14369_), .ZN(new_n14370_));
  NAND2_X1   g13350(.A1(new_n14350_), .A2(new_n14348_), .ZN(new_n14371_));
  INV_X1     g13351(.I(new_n14227_), .ZN(new_n14372_));
  AOI21_X1   g13352(.A1(new_n14220_), .A2(new_n14202_), .B(new_n14150_), .ZN(new_n14373_));
  NOR2_X1    g13353(.A1(new_n14373_), .A2(new_n14372_), .ZN(new_n14374_));
  OAI21_X1   g13354(.A1(new_n14348_), .A2(new_n14350_), .B(new_n14374_), .ZN(new_n14375_));
  NAND2_X1   g13355(.A1(new_n14375_), .A2(new_n14371_), .ZN(new_n14376_));
  INV_X1     g13356(.I(new_n14376_), .ZN(new_n14377_));
  AOI21_X1   g13357(.A1(new_n14370_), .A2(new_n14377_), .B(new_n14365_), .ZN(new_n14378_));
  NAND2_X1   g13358(.A1(new_n14376_), .A2(new_n14369_), .ZN(new_n14379_));
  INV_X1     g13359(.I(new_n14379_), .ZN(new_n14380_));
  NOR2_X1    g13360(.A1(new_n14378_), .A2(new_n14380_), .ZN(new_n14381_));
  INV_X1     g13361(.I(new_n14381_), .ZN(new_n14382_));
  NAND2_X1   g13362(.A1(new_n14382_), .A2(new_n14119_), .ZN(new_n14383_));
  XNOR2_X1   g13363(.A1(new_n14231_), .A2(new_n14232_), .ZN(new_n14384_));
  INV_X1     g13364(.I(new_n14314_), .ZN(new_n14385_));
  NAND2_X1   g13365(.A1(new_n14384_), .A2(new_n14385_), .ZN(new_n14386_));
  NAND2_X1   g13366(.A1(new_n14229_), .A2(new_n14386_), .ZN(new_n14387_));
  NAND3_X1   g13367(.A1(new_n14222_), .A2(new_n14228_), .A3(new_n14304_), .ZN(new_n14388_));
  NAND2_X1   g13368(.A1(new_n14326_), .A2(new_n14334_), .ZN(new_n14389_));
  AND2_X2    g13369(.A1(new_n14331_), .A2(new_n14333_), .Z(new_n14390_));
  NOR3_X1    g13370(.A1(new_n14385_), .A2(new_n14319_), .A3(new_n14335_), .ZN(new_n14391_));
  AOI21_X1   g13371(.A1(new_n14390_), .A2(new_n14391_), .B(new_n14341_), .ZN(new_n14392_));
  NOR3_X1    g13372(.A1(new_n14342_), .A2(new_n14313_), .A3(new_n14323_), .ZN(new_n14393_));
  OAI21_X1   g13373(.A1(new_n14392_), .A2(new_n14393_), .B(new_n14338_), .ZN(new_n14394_));
  NAND2_X1   g13374(.A1(new_n14394_), .A2(new_n14389_), .ZN(new_n14395_));
  AOI22_X1   g13375(.A1(new_n14387_), .A2(new_n14388_), .B1(new_n14395_), .B2(new_n14229_), .ZN(new_n14396_));
  XNOR2_X1   g13376(.A1(new_n14352_), .A2(new_n14361_), .ZN(new_n14397_));
  INV_X1     g13377(.I(new_n14397_), .ZN(new_n14398_));
  NAND2_X1   g13378(.A1(new_n14398_), .A2(new_n14396_), .ZN(new_n14399_));
  NAND2_X1   g13379(.A1(new_n14364_), .A2(new_n14362_), .ZN(new_n14400_));
  NAND2_X1   g13380(.A1(new_n14345_), .A2(new_n14400_), .ZN(new_n14401_));
  NAND2_X1   g13381(.A1(new_n13950_), .A2(new_n13957_), .ZN(new_n14402_));
  NAND3_X1   g13382(.A1(new_n14402_), .A2(new_n13954_), .A3(new_n14095_), .ZN(new_n14403_));
  XOR2_X1    g13383(.A1(new_n14403_), .A2(new_n14106_), .Z(new_n14404_));
  NAND2_X1   g13384(.A1(new_n14404_), .A2(new_n14089_), .ZN(new_n14405_));
  NOR2_X1    g13385(.A1(new_n13966_), .A2(new_n13960_), .ZN(new_n14406_));
  AOI21_X1   g13386(.A1(new_n13949_), .A2(new_n13955_), .B(new_n14048_), .ZN(new_n14407_));
  NOR3_X1    g13387(.A1(new_n13966_), .A2(new_n13960_), .A3(new_n14041_), .ZN(new_n14408_));
  NAND4_X1   g13388(.A1(new_n14078_), .A2(new_n14070_), .A3(new_n14072_), .A4(new_n14057_), .ZN(new_n14409_));
  XOR2_X1    g13389(.A1(new_n14409_), .A2(new_n14084_), .Z(new_n14410_));
  AOI21_X1   g13390(.A1(new_n14410_), .A2(new_n14080_), .B(new_n14074_), .ZN(new_n14411_));
  OAI22_X1   g13391(.A1(new_n14411_), .A2(new_n14406_), .B1(new_n14408_), .B2(new_n14407_), .ZN(new_n14412_));
  NAND2_X1   g13392(.A1(new_n14403_), .A2(new_n14106_), .ZN(new_n14413_));
  NAND2_X1   g13393(.A1(new_n14107_), .A2(new_n14097_), .ZN(new_n14414_));
  NAND2_X1   g13394(.A1(new_n14414_), .A2(new_n14413_), .ZN(new_n14415_));
  NAND2_X1   g13395(.A1(new_n14412_), .A2(new_n14415_), .ZN(new_n14416_));
  NAND4_X1   g13396(.A1(new_n14399_), .A2(new_n14401_), .A3(new_n14405_), .A4(new_n14416_), .ZN(new_n14417_));
  NOR3_X1    g13397(.A1(new_n14088_), .A2(new_n14408_), .A3(new_n14407_), .ZN(new_n14418_));
  NAND2_X1   g13398(.A1(new_n14043_), .A2(new_n14047_), .ZN(new_n14419_));
  NAND2_X1   g13399(.A1(new_n14041_), .A2(new_n14419_), .ZN(new_n14420_));
  NAND2_X1   g13400(.A1(new_n14233_), .A2(new_n14303_), .ZN(new_n14421_));
  NAND2_X1   g13401(.A1(new_n14386_), .A2(new_n14421_), .ZN(new_n14422_));
  NOR2_X1    g13402(.A1(new_n14422_), .A2(new_n14420_), .ZN(new_n14423_));
  NOR2_X1    g13403(.A1(new_n14418_), .A2(new_n14423_), .ZN(new_n14424_));
  NAND2_X1   g13404(.A1(new_n14418_), .A2(new_n14423_), .ZN(new_n14425_));
  INV_X1     g13405(.I(new_n14425_), .ZN(new_n14426_));
  AOI21_X1   g13406(.A1(new_n14387_), .A2(new_n14388_), .B(new_n14395_), .ZN(new_n14427_));
  NOR3_X1    g13407(.A1(new_n14344_), .A2(new_n14306_), .A3(new_n14305_), .ZN(new_n14428_));
  NOR2_X1    g13408(.A1(new_n14427_), .A2(new_n14428_), .ZN(new_n14429_));
  OAI22_X1   g13409(.A1(new_n14426_), .A2(new_n14424_), .B1(new_n14429_), .B2(new_n14418_), .ZN(new_n14430_));
  AOI22_X1   g13410(.A1(new_n14399_), .A2(new_n14401_), .B1(new_n14405_), .B2(new_n14416_), .ZN(new_n14431_));
  OAI21_X1   g13411(.A1(new_n14431_), .A2(new_n14430_), .B(new_n14417_), .ZN(new_n14432_));
  INV_X1     g13412(.I(new_n14352_), .ZN(new_n14433_));
  INV_X1     g13413(.I(new_n14361_), .ZN(new_n14434_));
  NAND3_X1   g13414(.A1(new_n14396_), .A2(new_n14433_), .A3(new_n14434_), .ZN(new_n14435_));
  NAND2_X1   g13415(.A1(new_n14435_), .A2(new_n14369_), .ZN(new_n14436_));
  NAND4_X1   g13416(.A1(new_n14396_), .A2(new_n14433_), .A3(new_n14434_), .A4(new_n14370_), .ZN(new_n14437_));
  AOI21_X1   g13417(.A1(new_n14436_), .A2(new_n14437_), .B(new_n14377_), .ZN(new_n14438_));
  NOR2_X1    g13418(.A1(new_n14365_), .A2(new_n14370_), .ZN(new_n14439_));
  INV_X1     g13419(.I(new_n14437_), .ZN(new_n14440_));
  NOR3_X1    g13420(.A1(new_n14439_), .A2(new_n14440_), .A3(new_n14376_), .ZN(new_n14441_));
  NOR2_X1    g13421(.A1(new_n14441_), .A2(new_n14438_), .ZN(new_n14442_));
  INV_X1     g13422(.I(new_n14116_), .ZN(new_n14443_));
  NAND2_X1   g13423(.A1(new_n14108_), .A2(new_n14112_), .ZN(new_n14444_));
  INV_X1     g13424(.I(new_n14112_), .ZN(new_n14445_));
  NAND4_X1   g13425(.A1(new_n14089_), .A2(new_n14097_), .A3(new_n14107_), .A4(new_n14445_), .ZN(new_n14446_));
  AOI21_X1   g13426(.A1(new_n14444_), .A2(new_n14446_), .B(new_n14443_), .ZN(new_n14447_));
  NAND2_X1   g13427(.A1(new_n14412_), .A2(new_n14413_), .ZN(new_n14448_));
  NOR2_X1    g13428(.A1(new_n14403_), .A2(new_n14106_), .ZN(new_n14449_));
  AOI21_X1   g13429(.A1(new_n14448_), .A2(new_n14449_), .B(new_n14445_), .ZN(new_n14450_));
  INV_X1     g13430(.I(new_n14446_), .ZN(new_n14451_));
  NOR3_X1    g13431(.A1(new_n14450_), .A2(new_n14451_), .A3(new_n14116_), .ZN(new_n14452_));
  NOR2_X1    g13432(.A1(new_n14452_), .A2(new_n14447_), .ZN(new_n14453_));
  AOI21_X1   g13433(.A1(new_n14442_), .A2(new_n14453_), .B(new_n14432_), .ZN(new_n14454_));
  XOR2_X1    g13434(.A1(new_n14116_), .A2(new_n14112_), .Z(new_n14455_));
  XOR2_X1    g13435(.A1(new_n14376_), .A2(new_n14369_), .Z(new_n14456_));
  NOR4_X1    g13436(.A1(new_n14455_), .A2(new_n14456_), .A3(new_n14108_), .A4(new_n14435_), .ZN(new_n14457_));
  INV_X1     g13437(.I(new_n14457_), .ZN(new_n14458_));
  NOR2_X1    g13438(.A1(new_n14454_), .A2(new_n14458_), .ZN(new_n14459_));
  NAND3_X1   g13439(.A1(new_n14117_), .A2(new_n14118_), .A3(new_n14379_), .ZN(new_n14460_));
  OR3_X2     g13440(.A1(new_n14459_), .A2(new_n14378_), .A3(new_n14460_), .Z(new_n14461_));
  NAND2_X1   g13441(.A1(new_n14461_), .A2(new_n14383_), .ZN(new_n14462_));
  NOR2_X1    g13442(.A1(new_n14462_), .A2(new_n13846_), .ZN(new_n14463_));
  INV_X1     g13443(.I(new_n14463_), .ZN(new_n14464_));
  AOI21_X1   g13444(.A1(new_n14119_), .A2(new_n14382_), .B(new_n13845_), .ZN(new_n14465_));
  AOI21_X1   g13445(.A1(new_n13806_), .A2(new_n13801_), .B(new_n13804_), .ZN(new_n14466_));
  NOR3_X1    g13446(.A1(new_n13800_), .A2(new_n13802_), .A3(new_n13793_), .ZN(new_n14467_));
  NOR2_X1    g13447(.A1(new_n14467_), .A2(new_n14466_), .ZN(new_n14468_));
  NOR2_X1    g13448(.A1(new_n14468_), .A2(new_n13828_), .ZN(new_n14469_));
  AOI21_X1   g13449(.A1(new_n13825_), .A2(new_n13826_), .B(new_n13824_), .ZN(new_n14470_));
  NOR3_X1    g13450(.A1(new_n13818_), .A2(new_n13822_), .A3(new_n13812_), .ZN(new_n14471_));
  NOR2_X1    g13451(.A1(new_n14471_), .A2(new_n14470_), .ZN(new_n14472_));
  NOR2_X1    g13452(.A1(new_n13808_), .A2(new_n14472_), .ZN(new_n14473_));
  OAI21_X1   g13453(.A1(new_n14469_), .A2(new_n14473_), .B(new_n13789_), .ZN(new_n14474_));
  NAND2_X1   g13454(.A1(new_n13779_), .A2(new_n13783_), .ZN(new_n14475_));
  NAND2_X1   g13455(.A1(new_n13785_), .A2(new_n13787_), .ZN(new_n14476_));
  NOR2_X1    g13456(.A1(new_n14475_), .A2(new_n14476_), .ZN(new_n14477_));
  INV_X1     g13457(.I(new_n13764_), .ZN(new_n14478_));
  INV_X1     g13458(.I(new_n13771_), .ZN(new_n14479_));
  OAI21_X1   g13459(.A1(new_n13401_), .A2(new_n13404_), .B(new_n13452_), .ZN(new_n14480_));
  NAND3_X1   g13460(.A1(new_n13482_), .A2(new_n13474_), .A3(new_n13473_), .ZN(new_n14481_));
  NAND2_X1   g13461(.A1(new_n14480_), .A2(new_n14481_), .ZN(new_n14482_));
  AOI22_X1   g13462(.A1(new_n14479_), .A2(new_n13772_), .B1(new_n14482_), .B2(new_n14478_), .ZN(new_n14483_));
  INV_X1     g13463(.I(new_n13788_), .ZN(new_n14484_));
  AOI21_X1   g13464(.A1(new_n14484_), .A2(new_n14483_), .B(new_n14477_), .ZN(new_n14485_));
  NOR2_X1    g13465(.A1(new_n14468_), .A2(new_n14472_), .ZN(new_n14486_));
  OAI21_X1   g13466(.A1(new_n14486_), .A2(new_n13829_), .B(new_n14485_), .ZN(new_n14487_));
  OAI21_X1   g13467(.A1(new_n14450_), .A2(new_n14451_), .B(new_n14116_), .ZN(new_n14488_));
  NAND3_X1   g13468(.A1(new_n14444_), .A2(new_n14443_), .A3(new_n14446_), .ZN(new_n14489_));
  NAND2_X1   g13469(.A1(new_n14488_), .A2(new_n14489_), .ZN(new_n14490_));
  NOR2_X1    g13470(.A1(new_n14442_), .A2(new_n14490_), .ZN(new_n14491_));
  OAI21_X1   g13471(.A1(new_n14439_), .A2(new_n14440_), .B(new_n14376_), .ZN(new_n14492_));
  NAND3_X1   g13472(.A1(new_n14436_), .A2(new_n14377_), .A3(new_n14437_), .ZN(new_n14493_));
  NAND2_X1   g13473(.A1(new_n14492_), .A2(new_n14493_), .ZN(new_n14494_));
  NOR2_X1    g13474(.A1(new_n14494_), .A2(new_n14453_), .ZN(new_n14495_));
  OAI21_X1   g13475(.A1(new_n14491_), .A2(new_n14495_), .B(new_n14432_), .ZN(new_n14496_));
  NOR2_X1    g13476(.A1(new_n14345_), .A2(new_n14397_), .ZN(new_n14497_));
  INV_X1     g13477(.I(new_n14362_), .ZN(new_n14498_));
  NOR2_X1    g13478(.A1(new_n14498_), .A2(new_n14363_), .ZN(new_n14499_));
  NOR2_X1    g13479(.A1(new_n14396_), .A2(new_n14499_), .ZN(new_n14500_));
  XOR2_X1    g13480(.A1(new_n14097_), .A2(new_n14106_), .Z(new_n14501_));
  NOR2_X1    g13481(.A1(new_n14501_), .A2(new_n14412_), .ZN(new_n14502_));
  NOR2_X1    g13482(.A1(new_n14107_), .A2(new_n14097_), .ZN(new_n14503_));
  NOR2_X1    g13483(.A1(new_n14503_), .A2(new_n14449_), .ZN(new_n14504_));
  NOR2_X1    g13484(.A1(new_n14089_), .A2(new_n14504_), .ZN(new_n14505_));
  NOR4_X1    g13485(.A1(new_n14497_), .A2(new_n14500_), .A3(new_n14502_), .A4(new_n14505_), .ZN(new_n14506_));
  INV_X1     g13486(.I(new_n14418_), .ZN(new_n14507_));
  INV_X1     g13487(.I(new_n14424_), .ZN(new_n14508_));
  OAI21_X1   g13488(.A1(new_n14305_), .A2(new_n14306_), .B(new_n14344_), .ZN(new_n14509_));
  NAND3_X1   g13489(.A1(new_n14387_), .A2(new_n14388_), .A3(new_n14395_), .ZN(new_n14510_));
  NAND2_X1   g13490(.A1(new_n14509_), .A2(new_n14510_), .ZN(new_n14511_));
  AOI22_X1   g13491(.A1(new_n14508_), .A2(new_n14425_), .B1(new_n14511_), .B2(new_n14507_), .ZN(new_n14512_));
  OAI22_X1   g13492(.A1(new_n14497_), .A2(new_n14500_), .B1(new_n14502_), .B2(new_n14505_), .ZN(new_n14513_));
  AOI21_X1   g13493(.A1(new_n14512_), .A2(new_n14513_), .B(new_n14506_), .ZN(new_n14514_));
  NOR4_X1    g13494(.A1(new_n14441_), .A2(new_n14438_), .A3(new_n14452_), .A4(new_n14447_), .ZN(new_n14515_));
  AOI22_X1   g13495(.A1(new_n14492_), .A2(new_n14493_), .B1(new_n14488_), .B2(new_n14489_), .ZN(new_n14516_));
  OAI21_X1   g13496(.A1(new_n14516_), .A2(new_n14515_), .B(new_n14514_), .ZN(new_n14517_));
  NAND4_X1   g13497(.A1(new_n14496_), .A2(new_n14474_), .A3(new_n14487_), .A4(new_n14517_), .ZN(new_n14518_));
  NOR2_X1    g13498(.A1(new_n14497_), .A2(new_n14500_), .ZN(new_n14519_));
  NAND2_X1   g13499(.A1(new_n14405_), .A2(new_n14416_), .ZN(new_n14520_));
  NAND2_X1   g13500(.A1(new_n14519_), .A2(new_n14520_), .ZN(new_n14521_));
  NAND2_X1   g13501(.A1(new_n14399_), .A2(new_n14401_), .ZN(new_n14522_));
  NOR2_X1    g13502(.A1(new_n14502_), .A2(new_n14505_), .ZN(new_n14523_));
  NAND2_X1   g13503(.A1(new_n14522_), .A2(new_n14523_), .ZN(new_n14524_));
  AOI21_X1   g13504(.A1(new_n14524_), .A2(new_n14521_), .B(new_n14430_), .ZN(new_n14525_));
  AOI21_X1   g13505(.A1(new_n14417_), .A2(new_n14513_), .B(new_n14512_), .ZN(new_n14526_));
  NAND2_X1   g13506(.A1(new_n13494_), .A2(new_n14476_), .ZN(new_n14527_));
  NAND2_X1   g13507(.A1(new_n14475_), .A2(new_n13762_), .ZN(new_n14528_));
  AOI21_X1   g13508(.A1(new_n14528_), .A2(new_n14527_), .B(new_n13777_), .ZN(new_n14529_));
  AOI21_X1   g13509(.A1(new_n14484_), .A2(new_n13763_), .B(new_n14483_), .ZN(new_n14530_));
  NOR4_X1    g13510(.A1(new_n14525_), .A2(new_n14530_), .A3(new_n14529_), .A4(new_n14526_), .ZN(new_n14531_));
  NOR2_X1    g13511(.A1(new_n13773_), .A2(new_n13771_), .ZN(new_n14532_));
  NAND2_X1   g13512(.A1(new_n14532_), .A2(new_n13776_), .ZN(new_n14533_));
  NAND2_X1   g13513(.A1(new_n14479_), .A2(new_n13772_), .ZN(new_n14534_));
  XNOR2_X1   g13514(.A1(new_n13766_), .A2(new_n13768_), .ZN(new_n14535_));
  XNOR2_X1   g13515(.A1(new_n14422_), .A2(new_n14420_), .ZN(new_n14536_));
  NOR2_X1    g13516(.A1(new_n14535_), .A2(new_n14536_), .ZN(new_n14537_));
  INV_X1     g13517(.I(new_n14537_), .ZN(new_n14538_));
  OAI21_X1   g13518(.A1(new_n14534_), .A2(new_n14482_), .B(new_n14538_), .ZN(new_n14539_));
  NAND3_X1   g13519(.A1(new_n14532_), .A2(new_n13776_), .A3(new_n14537_), .ZN(new_n14540_));
  AOI21_X1   g13520(.A1(new_n14508_), .A2(new_n14425_), .B(new_n14511_), .ZN(new_n14541_));
  NOR3_X1    g13521(.A1(new_n14426_), .A2(new_n14429_), .A3(new_n14424_), .ZN(new_n14542_));
  NOR2_X1    g13522(.A1(new_n14541_), .A2(new_n14542_), .ZN(new_n14543_));
  INV_X1     g13523(.I(new_n14543_), .ZN(new_n14544_));
  AOI22_X1   g13524(.A1(new_n14544_), .A2(new_n14533_), .B1(new_n14539_), .B2(new_n14540_), .ZN(new_n14545_));
  NOR2_X1    g13525(.A1(new_n14522_), .A2(new_n14523_), .ZN(new_n14546_));
  NOR2_X1    g13526(.A1(new_n14519_), .A2(new_n14520_), .ZN(new_n14547_));
  OAI21_X1   g13527(.A1(new_n14546_), .A2(new_n14547_), .B(new_n14512_), .ZN(new_n14548_));
  OAI21_X1   g13528(.A1(new_n14506_), .A2(new_n14431_), .B(new_n14430_), .ZN(new_n14549_));
  NAND2_X1   g13529(.A1(new_n14548_), .A2(new_n14549_), .ZN(new_n14550_));
  NOR2_X1    g13530(.A1(new_n14475_), .A2(new_n13762_), .ZN(new_n14551_));
  NOR2_X1    g13531(.A1(new_n13494_), .A2(new_n14476_), .ZN(new_n14552_));
  OAI21_X1   g13532(.A1(new_n14551_), .A2(new_n14552_), .B(new_n14483_), .ZN(new_n14553_));
  OAI21_X1   g13533(.A1(new_n14477_), .A2(new_n13788_), .B(new_n13777_), .ZN(new_n14554_));
  NAND2_X1   g13534(.A1(new_n14553_), .A2(new_n14554_), .ZN(new_n14555_));
  NAND2_X1   g13535(.A1(new_n14550_), .A2(new_n14555_), .ZN(new_n14556_));
  AOI21_X1   g13536(.A1(new_n14556_), .A2(new_n14545_), .B(new_n14531_), .ZN(new_n14557_));
  AOI22_X1   g13537(.A1(new_n14496_), .A2(new_n14517_), .B1(new_n14474_), .B2(new_n14487_), .ZN(new_n14558_));
  OAI21_X1   g13538(.A1(new_n14558_), .A2(new_n14557_), .B(new_n14518_), .ZN(new_n14559_));
  XOR2_X1    g13539(.A1(new_n13843_), .A2(new_n13842_), .Z(new_n14560_));
  NOR3_X1    g13540(.A1(new_n13830_), .A2(new_n13835_), .A3(new_n14560_), .ZN(new_n14561_));
  INV_X1     g13541(.I(new_n14119_), .ZN(new_n14562_));
  OAI21_X1   g13542(.A1(new_n14454_), .A2(new_n14458_), .B(new_n14382_), .ZN(new_n14563_));
  OAI21_X1   g13543(.A1(new_n14494_), .A2(new_n14490_), .B(new_n14514_), .ZN(new_n14564_));
  NAND3_X1   g13544(.A1(new_n14564_), .A2(new_n14381_), .A3(new_n14457_), .ZN(new_n14565_));
  AOI21_X1   g13545(.A1(new_n14563_), .A2(new_n14565_), .B(new_n14562_), .ZN(new_n14566_));
  AOI21_X1   g13546(.A1(new_n14564_), .A2(new_n14457_), .B(new_n14381_), .ZN(new_n14567_));
  NOR3_X1    g13547(.A1(new_n14454_), .A2(new_n14382_), .A3(new_n14458_), .ZN(new_n14568_));
  NOR3_X1    g13548(.A1(new_n14568_), .A2(new_n14567_), .A3(new_n14119_), .ZN(new_n14569_));
  NOR3_X1    g13549(.A1(new_n14569_), .A2(new_n14566_), .A3(new_n14561_), .ZN(new_n14570_));
  NAND3_X1   g13550(.A1(new_n14472_), .A2(new_n13803_), .A3(new_n13807_), .ZN(new_n14571_));
  NAND2_X1   g13551(.A1(new_n14571_), .A2(new_n14485_), .ZN(new_n14572_));
  INV_X1     g13552(.I(new_n14560_), .ZN(new_n14573_));
  NAND3_X1   g13553(.A1(new_n14573_), .A2(new_n14572_), .A3(new_n13834_), .ZN(new_n14574_));
  XNOR2_X1   g13554(.A1(new_n14381_), .A2(new_n14119_), .ZN(new_n14575_));
  NOR4_X1    g13555(.A1(new_n14574_), .A2(new_n14454_), .A3(new_n14458_), .A4(new_n14575_), .ZN(new_n14576_));
  OAI21_X1   g13556(.A1(new_n14559_), .A2(new_n14570_), .B(new_n14576_), .ZN(new_n14577_));
  OAI21_X1   g13557(.A1(new_n14461_), .A2(new_n14465_), .B(new_n14577_), .ZN(new_n14578_));
  NAND2_X1   g13558(.A1(new_n14578_), .A2(new_n14464_), .ZN(new_n14579_));
  NOR2_X1    g13559(.A1(new_n14579_), .A2(new_n13231_), .ZN(new_n14580_));
  NOR2_X1    g13560(.A1(new_n14569_), .A2(new_n14566_), .ZN(new_n14581_));
  INV_X1     g13561(.I(new_n14581_), .ZN(new_n14582_));
  NAND2_X1   g13562(.A1(new_n13808_), .A2(new_n14472_), .ZN(new_n14583_));
  NAND2_X1   g13563(.A1(new_n14468_), .A2(new_n13828_), .ZN(new_n14584_));
  AOI21_X1   g13564(.A1(new_n14584_), .A2(new_n14583_), .B(new_n14485_), .ZN(new_n14585_));
  NAND2_X1   g13565(.A1(new_n13808_), .A2(new_n13828_), .ZN(new_n14586_));
  AOI21_X1   g13566(.A1(new_n14586_), .A2(new_n14571_), .B(new_n13789_), .ZN(new_n14587_));
  NOR2_X1    g13567(.A1(new_n14585_), .A2(new_n14587_), .ZN(new_n14588_));
  NAND2_X1   g13568(.A1(new_n14494_), .A2(new_n14453_), .ZN(new_n14589_));
  NAND2_X1   g13569(.A1(new_n14442_), .A2(new_n14490_), .ZN(new_n14590_));
  AOI21_X1   g13570(.A1(new_n14590_), .A2(new_n14589_), .B(new_n14514_), .ZN(new_n14591_));
  NAND3_X1   g13571(.A1(new_n14453_), .A2(new_n14492_), .A3(new_n14493_), .ZN(new_n14592_));
  NAND2_X1   g13572(.A1(new_n14494_), .A2(new_n14490_), .ZN(new_n14593_));
  AOI21_X1   g13573(.A1(new_n14593_), .A2(new_n14592_), .B(new_n14432_), .ZN(new_n14594_));
  NOR2_X1    g13574(.A1(new_n14591_), .A2(new_n14594_), .ZN(new_n14595_));
  NAND4_X1   g13575(.A1(new_n14548_), .A2(new_n14553_), .A3(new_n14554_), .A4(new_n14549_), .ZN(new_n14596_));
  NAND2_X1   g13576(.A1(new_n14539_), .A2(new_n14540_), .ZN(new_n14597_));
  NOR2_X1    g13577(.A1(new_n14533_), .A2(new_n14538_), .ZN(new_n14598_));
  AOI21_X1   g13578(.A1(new_n14597_), .A2(new_n14543_), .B(new_n14598_), .ZN(new_n14599_));
  AOI22_X1   g13579(.A1(new_n14548_), .A2(new_n14549_), .B1(new_n14553_), .B2(new_n14554_), .ZN(new_n14600_));
  OAI21_X1   g13580(.A1(new_n14600_), .A2(new_n14599_), .B(new_n14596_), .ZN(new_n14601_));
  OAI21_X1   g13581(.A1(new_n14595_), .A2(new_n14588_), .B(new_n14601_), .ZN(new_n14602_));
  AOI21_X1   g13582(.A1(new_n14602_), .A2(new_n14518_), .B(new_n14561_), .ZN(new_n14603_));
  NOR2_X1    g13583(.A1(new_n14559_), .A2(new_n14574_), .ZN(new_n14604_));
  OAI21_X1   g13584(.A1(new_n14604_), .A2(new_n14603_), .B(new_n14582_), .ZN(new_n14605_));
  AOI21_X1   g13585(.A1(new_n14602_), .A2(new_n14518_), .B(new_n14574_), .ZN(new_n14606_));
  NOR2_X1    g13586(.A1(new_n14559_), .A2(new_n14561_), .ZN(new_n14607_));
  OAI21_X1   g13587(.A1(new_n14607_), .A2(new_n14606_), .B(new_n14581_), .ZN(new_n14608_));
  NAND3_X1   g13588(.A1(new_n13216_), .A2(new_n12488_), .A3(new_n12492_), .ZN(new_n14609_));
  NOR3_X1    g13589(.A1(new_n13225_), .A2(new_n13222_), .A3(new_n14609_), .ZN(new_n14610_));
  OAI21_X1   g13590(.A1(new_n13224_), .A2(new_n13223_), .B(new_n13051_), .ZN(new_n14611_));
  NAND3_X1   g13591(.A1(new_n13218_), .A2(new_n13221_), .A3(new_n13052_), .ZN(new_n14612_));
  AOI21_X1   g13592(.A1(new_n14611_), .A2(new_n14612_), .B(new_n13217_), .ZN(new_n14613_));
  OAI22_X1   g13593(.A1(new_n14610_), .A2(new_n14613_), .B1(new_n13205_), .B2(new_n13215_), .ZN(new_n14614_));
  NOR2_X1    g13594(.A1(new_n13215_), .A2(new_n13205_), .ZN(new_n14615_));
  NAND3_X1   g13595(.A1(new_n14611_), .A2(new_n14612_), .A3(new_n14609_), .ZN(new_n14616_));
  OAI21_X1   g13596(.A1(new_n13225_), .A2(new_n13222_), .B(new_n13217_), .ZN(new_n14617_));
  NAND2_X1   g13597(.A1(new_n14617_), .A2(new_n14616_), .ZN(new_n14618_));
  NAND2_X1   g13598(.A1(new_n14618_), .A2(new_n14615_), .ZN(new_n14619_));
  NAND4_X1   g13599(.A1(new_n14605_), .A2(new_n14608_), .A3(new_n14614_), .A4(new_n14619_), .ZN(new_n14620_));
  NAND2_X1   g13600(.A1(new_n14559_), .A2(new_n14574_), .ZN(new_n14621_));
  NAND3_X1   g13601(.A1(new_n14602_), .A2(new_n14518_), .A3(new_n14561_), .ZN(new_n14622_));
  AOI21_X1   g13602(.A1(new_n14621_), .A2(new_n14622_), .B(new_n14581_), .ZN(new_n14623_));
  NOR4_X1    g13603(.A1(new_n14591_), .A2(new_n14585_), .A3(new_n14594_), .A4(new_n14587_), .ZN(new_n14624_));
  NAND2_X1   g13604(.A1(new_n14474_), .A2(new_n14487_), .ZN(new_n14625_));
  NAND2_X1   g13605(.A1(new_n14496_), .A2(new_n14517_), .ZN(new_n14626_));
  AOI21_X1   g13606(.A1(new_n14626_), .A2(new_n14625_), .B(new_n14557_), .ZN(new_n14627_));
  OAI21_X1   g13607(.A1(new_n14627_), .A2(new_n14624_), .B(new_n14561_), .ZN(new_n14628_));
  NAND3_X1   g13608(.A1(new_n14602_), .A2(new_n14518_), .A3(new_n14574_), .ZN(new_n14629_));
  AOI21_X1   g13609(.A1(new_n14628_), .A2(new_n14629_), .B(new_n14582_), .ZN(new_n14630_));
  NOR2_X1    g13610(.A1(new_n14623_), .A2(new_n14630_), .ZN(new_n14631_));
  NOR2_X1    g13611(.A1(new_n14610_), .A2(new_n14613_), .ZN(new_n14632_));
  NOR2_X1    g13612(.A1(new_n14632_), .A2(new_n14615_), .ZN(new_n14633_));
  NAND2_X1   g13613(.A1(new_n13135_), .A2(new_n13138_), .ZN(new_n14634_));
  NAND2_X1   g13614(.A1(new_n13132_), .A2(new_n13133_), .ZN(new_n14635_));
  AOI21_X1   g13615(.A1(new_n14634_), .A2(new_n14635_), .B(new_n12447_), .ZN(new_n14636_));
  NAND2_X1   g13616(.A1(new_n13135_), .A2(new_n13133_), .ZN(new_n14637_));
  AOI21_X1   g13617(.A1(new_n14637_), .A2(new_n12487_), .B(new_n13129_), .ZN(new_n14638_));
  NOR2_X1    g13618(.A1(new_n14636_), .A2(new_n14638_), .ZN(new_n14639_));
  AOI21_X1   g13619(.A1(new_n13150_), .A2(new_n13152_), .B(new_n13147_), .ZN(new_n14640_));
  NOR2_X1    g13620(.A1(new_n14640_), .A2(new_n13086_), .ZN(new_n14641_));
  NOR2_X1    g13621(.A1(new_n13127_), .A2(new_n12163_), .ZN(new_n14642_));
  NOR2_X1    g13622(.A1(new_n12428_), .A2(new_n13122_), .ZN(new_n14643_));
  OAI21_X1   g13623(.A1(new_n14643_), .A2(new_n14642_), .B(new_n12445_), .ZN(new_n14644_));
  OAI21_X1   g13624(.A1(new_n13128_), .A2(new_n12429_), .B(new_n13116_), .ZN(new_n14645_));
  NAND3_X1   g13625(.A1(new_n14641_), .A2(new_n14644_), .A3(new_n14645_), .ZN(new_n14646_));
  AOI21_X1   g13626(.A1(new_n14644_), .A2(new_n14645_), .B(new_n14641_), .ZN(new_n14647_));
  OAI21_X1   g13627(.A1(new_n14647_), .A2(new_n13201_), .B(new_n14646_), .ZN(new_n14648_));
  NAND2_X1   g13628(.A1(new_n14639_), .A2(new_n14648_), .ZN(new_n14649_));
  NAND2_X1   g13629(.A1(new_n13219_), .A2(new_n13153_), .ZN(new_n14650_));
  NAND3_X1   g13630(.A1(new_n13086_), .A2(new_n13206_), .A3(new_n13207_), .ZN(new_n14651_));
  AOI21_X1   g13631(.A1(new_n14650_), .A2(new_n14651_), .B(new_n13102_), .ZN(new_n14652_));
  NAND2_X1   g13632(.A1(new_n13219_), .A2(new_n13086_), .ZN(new_n14653_));
  NAND3_X1   g13633(.A1(new_n13153_), .A2(new_n13206_), .A3(new_n13207_), .ZN(new_n14654_));
  AOI21_X1   g13634(.A1(new_n14653_), .A2(new_n14654_), .B(new_n13098_), .ZN(new_n14655_));
  NOR2_X1    g13635(.A1(new_n14655_), .A2(new_n14652_), .ZN(new_n14656_));
  OAI21_X1   g13636(.A1(new_n14639_), .A2(new_n14648_), .B(new_n14656_), .ZN(new_n14657_));
  NAND2_X1   g13637(.A1(new_n14657_), .A2(new_n14649_), .ZN(new_n14658_));
  AOI21_X1   g13638(.A1(new_n14616_), .A2(new_n14617_), .B(new_n14658_), .ZN(new_n14659_));
  NOR2_X1    g13639(.A1(new_n14659_), .A2(new_n14633_), .ZN(new_n14660_));
  NOR2_X1    g13640(.A1(new_n14595_), .A2(new_n14625_), .ZN(new_n14661_));
  NOR2_X1    g13641(.A1(new_n14626_), .A2(new_n14588_), .ZN(new_n14662_));
  OAI21_X1   g13642(.A1(new_n14661_), .A2(new_n14662_), .B(new_n14601_), .ZN(new_n14663_));
  OAI21_X1   g13643(.A1(new_n14558_), .A2(new_n14624_), .B(new_n14557_), .ZN(new_n14664_));
  NAND2_X1   g13644(.A1(new_n14663_), .A2(new_n14664_), .ZN(new_n14665_));
  NOR2_X1    g13645(.A1(new_n14525_), .A2(new_n14526_), .ZN(new_n14666_));
  NAND2_X1   g13646(.A1(new_n14666_), .A2(new_n14555_), .ZN(new_n14667_));
  NOR2_X1    g13647(.A1(new_n14530_), .A2(new_n14529_), .ZN(new_n14668_));
  NAND2_X1   g13648(.A1(new_n14668_), .A2(new_n14550_), .ZN(new_n14669_));
  AOI21_X1   g13649(.A1(new_n14669_), .A2(new_n14667_), .B(new_n14599_), .ZN(new_n14670_));
  AOI21_X1   g13650(.A1(new_n14556_), .A2(new_n14596_), .B(new_n14545_), .ZN(new_n14671_));
  NAND2_X1   g13651(.A1(new_n14644_), .A2(new_n14645_), .ZN(new_n14672_));
  NAND2_X1   g13652(.A1(new_n14672_), .A2(new_n14641_), .ZN(new_n14673_));
  NOR2_X1    g13653(.A1(new_n13158_), .A2(new_n13159_), .ZN(new_n14674_));
  NAND2_X1   g13654(.A1(new_n14674_), .A2(new_n13155_), .ZN(new_n14675_));
  AOI21_X1   g13655(.A1(new_n14673_), .A2(new_n14675_), .B(new_n13201_), .ZN(new_n14676_));
  AOI21_X1   g13656(.A1(new_n13203_), .A2(new_n14646_), .B(new_n13202_), .ZN(new_n14677_));
  NOR4_X1    g13657(.A1(new_n14670_), .A2(new_n14671_), .A3(new_n14677_), .A4(new_n14676_), .ZN(new_n14678_));
  NOR3_X1    g13658(.A1(new_n13186_), .A2(new_n13196_), .A3(new_n13199_), .ZN(new_n14679_));
  AOI21_X1   g13659(.A1(new_n13177_), .A2(new_n13175_), .B(new_n13179_), .ZN(new_n14680_));
  OR2_X2     g13660(.A1(new_n13184_), .A2(new_n14680_), .Z(new_n14681_));
  NAND2_X1   g13661(.A1(new_n14535_), .A2(new_n14536_), .ZN(new_n14682_));
  NAND2_X1   g13662(.A1(new_n14538_), .A2(new_n14682_), .ZN(new_n14683_));
  NOR2_X1    g13663(.A1(new_n14681_), .A2(new_n14683_), .ZN(new_n14684_));
  NOR2_X1    g13664(.A1(new_n14679_), .A2(new_n14684_), .ZN(new_n14685_));
  INV_X1     g13665(.I(new_n14684_), .ZN(new_n14686_));
  NOR4_X1    g13666(.A1(new_n14686_), .A2(new_n13186_), .A3(new_n13196_), .A4(new_n13199_), .ZN(new_n14687_));
  XOR2_X1    g13667(.A1(new_n14597_), .A2(new_n14543_), .Z(new_n14688_));
  OAI22_X1   g13668(.A1(new_n14688_), .A2(new_n14679_), .B1(new_n14687_), .B2(new_n14685_), .ZN(new_n14689_));
  INV_X1     g13669(.I(new_n14689_), .ZN(new_n14690_));
  OAI22_X1   g13670(.A1(new_n14670_), .A2(new_n14671_), .B1(new_n14677_), .B2(new_n14676_), .ZN(new_n14691_));
  AOI21_X1   g13671(.A1(new_n14690_), .A2(new_n14691_), .B(new_n14678_), .ZN(new_n14692_));
  NOR2_X1    g13672(.A1(new_n14665_), .A2(new_n14692_), .ZN(new_n14693_));
  NOR2_X1    g13673(.A1(new_n14639_), .A2(new_n14648_), .ZN(new_n14694_));
  OAI21_X1   g13674(.A1(new_n13205_), .A2(new_n14694_), .B(new_n13214_), .ZN(new_n14695_));
  NOR2_X1    g13675(.A1(new_n13204_), .A2(new_n14639_), .ZN(new_n14696_));
  AOI21_X1   g13676(.A1(new_n14672_), .A2(new_n13155_), .B(new_n13201_), .ZN(new_n14697_));
  NOR4_X1    g13677(.A1(new_n14697_), .A2(new_n14636_), .A3(new_n14638_), .A4(new_n13160_), .ZN(new_n14698_));
  OAI21_X1   g13678(.A1(new_n14696_), .A2(new_n14698_), .B(new_n14656_), .ZN(new_n14699_));
  NAND2_X1   g13679(.A1(new_n14695_), .A2(new_n14699_), .ZN(new_n14700_));
  AOI21_X1   g13680(.A1(new_n14665_), .A2(new_n14692_), .B(new_n14700_), .ZN(new_n14701_));
  OAI22_X1   g13681(.A1(new_n14631_), .A2(new_n14660_), .B1(new_n14701_), .B2(new_n14693_), .ZN(new_n14702_));
  OAI21_X1   g13682(.A1(new_n14568_), .A2(new_n14567_), .B(new_n14119_), .ZN(new_n14703_));
  NAND3_X1   g13683(.A1(new_n14563_), .A2(new_n14565_), .A3(new_n14562_), .ZN(new_n14704_));
  NAND3_X1   g13684(.A1(new_n14703_), .A2(new_n14704_), .A3(new_n14574_), .ZN(new_n14705_));
  NAND3_X1   g13685(.A1(new_n14705_), .A2(new_n14602_), .A3(new_n14518_), .ZN(new_n14706_));
  AOI21_X1   g13686(.A1(new_n14706_), .A2(new_n14576_), .B(new_n14462_), .ZN(new_n14707_));
  INV_X1     g13687(.I(new_n14462_), .ZN(new_n14708_));
  NOR2_X1    g13688(.A1(new_n14577_), .A2(new_n14708_), .ZN(new_n14709_));
  OAI21_X1   g13689(.A1(new_n14709_), .A2(new_n14707_), .B(new_n13845_), .ZN(new_n14710_));
  NAND2_X1   g13690(.A1(new_n14577_), .A2(new_n14708_), .ZN(new_n14711_));
  NAND3_X1   g13691(.A1(new_n14706_), .A2(new_n14462_), .A3(new_n14576_), .ZN(new_n14712_));
  NAND3_X1   g13692(.A1(new_n14711_), .A2(new_n14712_), .A3(new_n13846_), .ZN(new_n14713_));
  INV_X1     g13693(.I(new_n13109_), .ZN(new_n14714_));
  NAND3_X1   g13694(.A1(new_n14616_), .A2(new_n14657_), .A3(new_n14649_), .ZN(new_n14715_));
  INV_X1     g13695(.I(new_n13229_), .ZN(new_n14716_));
  AOI21_X1   g13696(.A1(new_n14715_), .A2(new_n14716_), .B(new_n14714_), .ZN(new_n14717_));
  NOR3_X1    g13697(.A1(new_n13227_), .A2(new_n13109_), .A3(new_n13229_), .ZN(new_n14718_));
  OAI21_X1   g13698(.A1(new_n14718_), .A2(new_n14717_), .B(new_n12504_), .ZN(new_n14719_));
  OAI21_X1   g13699(.A1(new_n13227_), .A2(new_n13229_), .B(new_n13109_), .ZN(new_n14720_));
  NAND3_X1   g13700(.A1(new_n14715_), .A2(new_n14714_), .A3(new_n14716_), .ZN(new_n14721_));
  NAND3_X1   g13701(.A1(new_n14720_), .A2(new_n14721_), .A3(new_n12503_), .ZN(new_n14722_));
  NAND4_X1   g13702(.A1(new_n14710_), .A2(new_n14713_), .A3(new_n14719_), .A4(new_n14722_), .ZN(new_n14723_));
  NAND3_X1   g13703(.A1(new_n14723_), .A2(new_n14620_), .A3(new_n14702_), .ZN(new_n14724_));
  NAND2_X1   g13704(.A1(new_n14715_), .A2(new_n14716_), .ZN(new_n14725_));
  XOR2_X1    g13705(.A1(new_n14462_), .A2(new_n13846_), .Z(new_n14726_));
  XNOR2_X1   g13706(.A1(new_n13109_), .A2(new_n12503_), .ZN(new_n14727_));
  NOR4_X1    g13707(.A1(new_n14726_), .A2(new_n14725_), .A3(new_n14577_), .A4(new_n14727_), .ZN(new_n14728_));
  NAND4_X1   g13708(.A1(new_n14578_), .A2(new_n13110_), .A3(new_n13230_), .A4(new_n14464_), .ZN(new_n14729_));
  AOI21_X1   g13709(.A1(new_n14724_), .A2(new_n14728_), .B(new_n14729_), .ZN(new_n14730_));
  INV_X1     g13710(.I(\A[646] ), .ZN(new_n14731_));
  NOR2_X1    g13711(.A1(\A[647] ), .A2(\A[648] ), .ZN(new_n14732_));
  NAND2_X1   g13712(.A1(\A[647] ), .A2(\A[648] ), .ZN(new_n14733_));
  AOI21_X1   g13713(.A1(new_n14731_), .A2(new_n14733_), .B(new_n14732_), .ZN(new_n14734_));
  INV_X1     g13714(.I(new_n14734_), .ZN(new_n14735_));
  INV_X1     g13715(.I(\A[643] ), .ZN(new_n14736_));
  NOR2_X1    g13716(.A1(\A[644] ), .A2(\A[645] ), .ZN(new_n14737_));
  NAND2_X1   g13717(.A1(\A[644] ), .A2(\A[645] ), .ZN(new_n14738_));
  AOI21_X1   g13718(.A1(new_n14736_), .A2(new_n14738_), .B(new_n14737_), .ZN(new_n14739_));
  INV_X1     g13719(.I(\A[644] ), .ZN(new_n14740_));
  NAND2_X1   g13720(.A1(new_n14740_), .A2(\A[645] ), .ZN(new_n14741_));
  INV_X1     g13721(.I(\A[645] ), .ZN(new_n14742_));
  NAND2_X1   g13722(.A1(new_n14742_), .A2(\A[644] ), .ZN(new_n14743_));
  AOI21_X1   g13723(.A1(new_n14741_), .A2(new_n14743_), .B(new_n14736_), .ZN(new_n14744_));
  INV_X1     g13724(.I(new_n14737_), .ZN(new_n14745_));
  AOI21_X1   g13725(.A1(new_n14745_), .A2(new_n14738_), .B(\A[643] ), .ZN(new_n14746_));
  NOR2_X1    g13726(.A1(new_n14746_), .A2(new_n14744_), .ZN(new_n14747_));
  INV_X1     g13727(.I(\A[647] ), .ZN(new_n14748_));
  NAND2_X1   g13728(.A1(new_n14748_), .A2(\A[648] ), .ZN(new_n14749_));
  INV_X1     g13729(.I(\A[648] ), .ZN(new_n14750_));
  NAND2_X1   g13730(.A1(new_n14750_), .A2(\A[647] ), .ZN(new_n14751_));
  AOI21_X1   g13731(.A1(new_n14749_), .A2(new_n14751_), .B(new_n14731_), .ZN(new_n14752_));
  INV_X1     g13732(.I(new_n14732_), .ZN(new_n14753_));
  AOI21_X1   g13733(.A1(new_n14753_), .A2(new_n14733_), .B(\A[646] ), .ZN(new_n14754_));
  NOR2_X1    g13734(.A1(new_n14754_), .A2(new_n14752_), .ZN(new_n14755_));
  NAND2_X1   g13735(.A1(new_n14747_), .A2(new_n14755_), .ZN(new_n14756_));
  NAND2_X1   g13736(.A1(new_n14756_), .A2(new_n14739_), .ZN(new_n14757_));
  INV_X1     g13737(.I(new_n14739_), .ZN(new_n14758_));
  NOR4_X1    g13738(.A1(new_n14744_), .A2(new_n14746_), .A3(new_n14754_), .A4(new_n14752_), .ZN(new_n14759_));
  NAND2_X1   g13739(.A1(new_n14759_), .A2(new_n14758_), .ZN(new_n14760_));
  AOI21_X1   g13740(.A1(new_n14757_), .A2(new_n14760_), .B(new_n14735_), .ZN(new_n14761_));
  AND3_X2    g13741(.A1(new_n14757_), .A2(new_n14735_), .A3(new_n14760_), .Z(new_n14762_));
  NOR2_X1    g13742(.A1(new_n14762_), .A2(new_n14761_), .ZN(new_n14763_));
  INV_X1     g13743(.I(new_n14763_), .ZN(new_n14764_));
  INV_X1     g13744(.I(\A[652] ), .ZN(new_n14765_));
  NOR2_X1    g13745(.A1(\A[653] ), .A2(\A[654] ), .ZN(new_n14766_));
  NAND2_X1   g13746(.A1(\A[653] ), .A2(\A[654] ), .ZN(new_n14767_));
  AOI21_X1   g13747(.A1(new_n14765_), .A2(new_n14767_), .B(new_n14766_), .ZN(new_n14768_));
  INV_X1     g13748(.I(new_n14768_), .ZN(new_n14769_));
  INV_X1     g13749(.I(\A[649] ), .ZN(new_n14770_));
  NOR2_X1    g13750(.A1(\A[650] ), .A2(\A[651] ), .ZN(new_n14771_));
  NAND2_X1   g13751(.A1(\A[650] ), .A2(\A[651] ), .ZN(new_n14772_));
  AOI21_X1   g13752(.A1(new_n14770_), .A2(new_n14772_), .B(new_n14771_), .ZN(new_n14773_));
  INV_X1     g13753(.I(new_n14773_), .ZN(new_n14774_));
  NOR2_X1    g13754(.A1(new_n14769_), .A2(new_n14774_), .ZN(new_n14775_));
  INV_X1     g13755(.I(new_n14775_), .ZN(new_n14776_));
  INV_X1     g13756(.I(\A[650] ), .ZN(new_n14777_));
  NAND2_X1   g13757(.A1(new_n14777_), .A2(\A[651] ), .ZN(new_n14778_));
  INV_X1     g13758(.I(\A[651] ), .ZN(new_n14779_));
  NAND2_X1   g13759(.A1(new_n14779_), .A2(\A[650] ), .ZN(new_n14780_));
  AOI21_X1   g13760(.A1(new_n14778_), .A2(new_n14780_), .B(new_n14770_), .ZN(new_n14781_));
  INV_X1     g13761(.I(new_n14771_), .ZN(new_n14782_));
  AOI21_X1   g13762(.A1(new_n14782_), .A2(new_n14772_), .B(\A[649] ), .ZN(new_n14783_));
  NOR2_X1    g13763(.A1(new_n14783_), .A2(new_n14781_), .ZN(new_n14784_));
  INV_X1     g13764(.I(\A[654] ), .ZN(new_n14785_));
  NOR2_X1    g13765(.A1(new_n14785_), .A2(\A[653] ), .ZN(new_n14786_));
  INV_X1     g13766(.I(\A[653] ), .ZN(new_n14787_));
  NOR2_X1    g13767(.A1(new_n14787_), .A2(\A[654] ), .ZN(new_n14788_));
  OAI21_X1   g13768(.A1(new_n14786_), .A2(new_n14788_), .B(\A[652] ), .ZN(new_n14789_));
  INV_X1     g13769(.I(new_n14767_), .ZN(new_n14790_));
  OAI21_X1   g13770(.A1(new_n14790_), .A2(new_n14766_), .B(new_n14765_), .ZN(new_n14791_));
  NAND2_X1   g13771(.A1(new_n14789_), .A2(new_n14791_), .ZN(new_n14792_));
  NAND2_X1   g13772(.A1(new_n14784_), .A2(new_n14792_), .ZN(new_n14793_));
  NOR2_X1    g13773(.A1(new_n14779_), .A2(\A[650] ), .ZN(new_n14794_));
  NOR2_X1    g13774(.A1(new_n14777_), .A2(\A[651] ), .ZN(new_n14795_));
  OAI21_X1   g13775(.A1(new_n14794_), .A2(new_n14795_), .B(\A[649] ), .ZN(new_n14796_));
  INV_X1     g13776(.I(new_n14772_), .ZN(new_n14797_));
  OAI21_X1   g13777(.A1(new_n14797_), .A2(new_n14771_), .B(new_n14770_), .ZN(new_n14798_));
  NAND2_X1   g13778(.A1(new_n14796_), .A2(new_n14798_), .ZN(new_n14799_));
  NAND2_X1   g13779(.A1(new_n14787_), .A2(\A[654] ), .ZN(new_n14800_));
  NAND2_X1   g13780(.A1(new_n14785_), .A2(\A[653] ), .ZN(new_n14801_));
  AOI21_X1   g13781(.A1(new_n14800_), .A2(new_n14801_), .B(new_n14765_), .ZN(new_n14802_));
  INV_X1     g13782(.I(new_n14766_), .ZN(new_n14803_));
  AOI21_X1   g13783(.A1(new_n14803_), .A2(new_n14767_), .B(\A[652] ), .ZN(new_n14804_));
  NOR2_X1    g13784(.A1(new_n14804_), .A2(new_n14802_), .ZN(new_n14805_));
  NAND2_X1   g13785(.A1(new_n14805_), .A2(new_n14799_), .ZN(new_n14806_));
  AOI21_X1   g13786(.A1(new_n14793_), .A2(new_n14806_), .B(new_n14776_), .ZN(new_n14807_));
  INV_X1     g13787(.I(new_n14807_), .ZN(new_n14808_));
  NOR2_X1    g13788(.A1(new_n14799_), .A2(new_n14792_), .ZN(new_n14809_));
  NOR2_X1    g13789(.A1(new_n14809_), .A2(new_n14774_), .ZN(new_n14810_));
  NAND2_X1   g13790(.A1(new_n14784_), .A2(new_n14805_), .ZN(new_n14811_));
  NOR2_X1    g13791(.A1(new_n14811_), .A2(new_n14773_), .ZN(new_n14812_));
  OAI21_X1   g13792(.A1(new_n14810_), .A2(new_n14812_), .B(new_n14768_), .ZN(new_n14813_));
  NAND2_X1   g13793(.A1(new_n14811_), .A2(new_n14773_), .ZN(new_n14814_));
  NAND2_X1   g13794(.A1(new_n14809_), .A2(new_n14774_), .ZN(new_n14815_));
  NAND3_X1   g13795(.A1(new_n14815_), .A2(new_n14814_), .A3(new_n14769_), .ZN(new_n14816_));
  NAND3_X1   g13796(.A1(new_n14813_), .A2(new_n14816_), .A3(new_n14808_), .ZN(new_n14817_));
  NOR2_X1    g13797(.A1(new_n14811_), .A2(new_n14776_), .ZN(new_n14818_));
  NOR2_X1    g13798(.A1(new_n14784_), .A2(new_n14805_), .ZN(new_n14819_));
  NOR2_X1    g13799(.A1(new_n14819_), .A2(new_n14809_), .ZN(new_n14820_));
  NOR2_X1    g13800(.A1(new_n14747_), .A2(new_n14755_), .ZN(new_n14821_));
  NOR2_X1    g13801(.A1(new_n14821_), .A2(new_n14759_), .ZN(new_n14822_));
  NAND2_X1   g13802(.A1(new_n14734_), .A2(new_n14739_), .ZN(new_n14823_));
  NOR2_X1    g13803(.A1(new_n14756_), .A2(new_n14823_), .ZN(new_n14824_));
  NAND4_X1   g13804(.A1(new_n14818_), .A2(new_n14820_), .A3(new_n14822_), .A4(new_n14824_), .ZN(new_n14825_));
  NOR2_X1    g13805(.A1(new_n14817_), .A2(new_n14825_), .ZN(new_n14826_));
  INV_X1     g13806(.I(new_n14826_), .ZN(new_n14827_));
  NAND2_X1   g13807(.A1(new_n14817_), .A2(new_n14825_), .ZN(new_n14828_));
  AOI21_X1   g13808(.A1(new_n14827_), .A2(new_n14828_), .B(new_n14764_), .ZN(new_n14829_));
  NAND2_X1   g13809(.A1(new_n14820_), .A2(new_n14818_), .ZN(new_n14830_));
  NAND2_X1   g13810(.A1(new_n14822_), .A2(new_n14824_), .ZN(new_n14831_));
  NOR2_X1    g13811(.A1(new_n14830_), .A2(new_n14831_), .ZN(new_n14832_));
  NAND2_X1   g13812(.A1(new_n14817_), .A2(new_n14832_), .ZN(new_n14833_));
  NAND2_X1   g13813(.A1(new_n14813_), .A2(new_n14816_), .ZN(new_n14834_));
  NAND3_X1   g13814(.A1(new_n14820_), .A2(new_n14818_), .A3(new_n14822_), .ZN(new_n14835_));
  NOR3_X1    g13815(.A1(new_n14807_), .A2(new_n14756_), .A3(new_n14823_), .ZN(new_n14836_));
  OAI21_X1   g13816(.A1(new_n14834_), .A2(new_n14835_), .B(new_n14836_), .ZN(new_n14837_));
  AND3_X2    g13817(.A1(new_n14833_), .A2(new_n14837_), .A3(new_n14763_), .Z(new_n14838_));
  NOR2_X1    g13818(.A1(new_n14829_), .A2(new_n14838_), .ZN(new_n14839_));
  INV_X1     g13819(.I(new_n14828_), .ZN(new_n14840_));
  OAI21_X1   g13820(.A1(new_n14840_), .A2(new_n14826_), .B(new_n14763_), .ZN(new_n14841_));
  NAND3_X1   g13821(.A1(new_n14833_), .A2(new_n14837_), .A3(new_n14763_), .ZN(new_n14842_));
  XOR2_X1    g13822(.A1(new_n14830_), .A2(new_n14831_), .Z(new_n14843_));
  INV_X1     g13823(.I(\A[637] ), .ZN(new_n14844_));
  INV_X1     g13824(.I(\A[638] ), .ZN(new_n14845_));
  NAND2_X1   g13825(.A1(new_n14845_), .A2(\A[639] ), .ZN(new_n14846_));
  INV_X1     g13826(.I(\A[639] ), .ZN(new_n14847_));
  NAND2_X1   g13827(.A1(new_n14847_), .A2(\A[638] ), .ZN(new_n14848_));
  AOI21_X1   g13828(.A1(new_n14846_), .A2(new_n14848_), .B(new_n14844_), .ZN(new_n14849_));
  NOR2_X1    g13829(.A1(\A[638] ), .A2(\A[639] ), .ZN(new_n14850_));
  INV_X1     g13830(.I(new_n14850_), .ZN(new_n14851_));
  NAND2_X1   g13831(.A1(\A[638] ), .A2(\A[639] ), .ZN(new_n14852_));
  AOI21_X1   g13832(.A1(new_n14851_), .A2(new_n14852_), .B(\A[637] ), .ZN(new_n14853_));
  NOR2_X1    g13833(.A1(new_n14853_), .A2(new_n14849_), .ZN(new_n14854_));
  INV_X1     g13834(.I(\A[640] ), .ZN(new_n14855_));
  INV_X1     g13835(.I(\A[641] ), .ZN(new_n14856_));
  NAND2_X1   g13836(.A1(new_n14856_), .A2(\A[642] ), .ZN(new_n14857_));
  INV_X1     g13837(.I(\A[642] ), .ZN(new_n14858_));
  NAND2_X1   g13838(.A1(new_n14858_), .A2(\A[641] ), .ZN(new_n14859_));
  AOI21_X1   g13839(.A1(new_n14857_), .A2(new_n14859_), .B(new_n14855_), .ZN(new_n14860_));
  NOR2_X1    g13840(.A1(\A[641] ), .A2(\A[642] ), .ZN(new_n14861_));
  INV_X1     g13841(.I(new_n14861_), .ZN(new_n14862_));
  NAND2_X1   g13842(.A1(\A[641] ), .A2(\A[642] ), .ZN(new_n14863_));
  AOI21_X1   g13843(.A1(new_n14862_), .A2(new_n14863_), .B(\A[640] ), .ZN(new_n14864_));
  NOR2_X1    g13844(.A1(new_n14864_), .A2(new_n14860_), .ZN(new_n14865_));
  NAND2_X1   g13845(.A1(new_n14854_), .A2(new_n14865_), .ZN(new_n14866_));
  AOI21_X1   g13846(.A1(new_n14855_), .A2(new_n14863_), .B(new_n14861_), .ZN(new_n14867_));
  AOI21_X1   g13847(.A1(new_n14844_), .A2(new_n14852_), .B(new_n14850_), .ZN(new_n14868_));
  NAND2_X1   g13848(.A1(new_n14867_), .A2(new_n14868_), .ZN(new_n14869_));
  NOR2_X1    g13849(.A1(new_n14866_), .A2(new_n14869_), .ZN(new_n14870_));
  INV_X1     g13850(.I(new_n14870_), .ZN(new_n14871_));
  NOR2_X1    g13851(.A1(new_n14847_), .A2(\A[638] ), .ZN(new_n14872_));
  NOR2_X1    g13852(.A1(new_n14845_), .A2(\A[639] ), .ZN(new_n14873_));
  OAI21_X1   g13853(.A1(new_n14872_), .A2(new_n14873_), .B(\A[637] ), .ZN(new_n14874_));
  INV_X1     g13854(.I(new_n14852_), .ZN(new_n14875_));
  OAI21_X1   g13855(.A1(new_n14875_), .A2(new_n14850_), .B(new_n14844_), .ZN(new_n14876_));
  NAND2_X1   g13856(.A1(new_n14874_), .A2(new_n14876_), .ZN(new_n14877_));
  NOR2_X1    g13857(.A1(new_n14858_), .A2(\A[641] ), .ZN(new_n14878_));
  NOR2_X1    g13858(.A1(new_n14856_), .A2(\A[642] ), .ZN(new_n14879_));
  OAI21_X1   g13859(.A1(new_n14878_), .A2(new_n14879_), .B(\A[640] ), .ZN(new_n14880_));
  INV_X1     g13860(.I(new_n14863_), .ZN(new_n14881_));
  OAI21_X1   g13861(.A1(new_n14881_), .A2(new_n14861_), .B(new_n14855_), .ZN(new_n14882_));
  NAND2_X1   g13862(.A1(new_n14880_), .A2(new_n14882_), .ZN(new_n14883_));
  NAND2_X1   g13863(.A1(new_n14877_), .A2(new_n14883_), .ZN(new_n14884_));
  NAND2_X1   g13864(.A1(new_n14866_), .A2(new_n14884_), .ZN(new_n14885_));
  INV_X1     g13865(.I(\A[631] ), .ZN(new_n14886_));
  INV_X1     g13866(.I(\A[632] ), .ZN(new_n14887_));
  NAND2_X1   g13867(.A1(new_n14887_), .A2(\A[633] ), .ZN(new_n14888_));
  INV_X1     g13868(.I(\A[633] ), .ZN(new_n14889_));
  NAND2_X1   g13869(.A1(new_n14889_), .A2(\A[632] ), .ZN(new_n14890_));
  AOI21_X1   g13870(.A1(new_n14888_), .A2(new_n14890_), .B(new_n14886_), .ZN(new_n14891_));
  NAND2_X1   g13871(.A1(new_n14887_), .A2(new_n14889_), .ZN(new_n14892_));
  NAND2_X1   g13872(.A1(\A[632] ), .A2(\A[633] ), .ZN(new_n14893_));
  AOI21_X1   g13873(.A1(new_n14892_), .A2(new_n14893_), .B(\A[631] ), .ZN(new_n14894_));
  NOR2_X1    g13874(.A1(new_n14894_), .A2(new_n14891_), .ZN(new_n14895_));
  INV_X1     g13875(.I(\A[634] ), .ZN(new_n14896_));
  INV_X1     g13876(.I(\A[635] ), .ZN(new_n14897_));
  NAND2_X1   g13877(.A1(new_n14897_), .A2(\A[636] ), .ZN(new_n14898_));
  INV_X1     g13878(.I(\A[636] ), .ZN(new_n14899_));
  NAND2_X1   g13879(.A1(new_n14899_), .A2(\A[635] ), .ZN(new_n14900_));
  AOI21_X1   g13880(.A1(new_n14898_), .A2(new_n14900_), .B(new_n14896_), .ZN(new_n14901_));
  NAND2_X1   g13881(.A1(new_n14897_), .A2(new_n14899_), .ZN(new_n14902_));
  NAND2_X1   g13882(.A1(\A[635] ), .A2(\A[636] ), .ZN(new_n14903_));
  AOI21_X1   g13883(.A1(new_n14902_), .A2(new_n14903_), .B(\A[634] ), .ZN(new_n14904_));
  NOR2_X1    g13884(.A1(new_n14904_), .A2(new_n14901_), .ZN(new_n14905_));
  NAND2_X1   g13885(.A1(new_n14903_), .A2(new_n14896_), .ZN(new_n14906_));
  NAND2_X1   g13886(.A1(new_n14906_), .A2(new_n14902_), .ZN(new_n14907_));
  NAND2_X1   g13887(.A1(new_n14893_), .A2(new_n14886_), .ZN(new_n14908_));
  NAND2_X1   g13888(.A1(new_n14908_), .A2(new_n14892_), .ZN(new_n14909_));
  NOR2_X1    g13889(.A1(new_n14907_), .A2(new_n14909_), .ZN(new_n14910_));
  NOR2_X1    g13890(.A1(new_n14871_), .A2(new_n14885_), .ZN(new_n14911_));
  NOR2_X1    g13891(.A1(new_n14843_), .A2(new_n14911_), .ZN(new_n14912_));
  AOI21_X1   g13892(.A1(new_n14841_), .A2(new_n14842_), .B(new_n14912_), .ZN(new_n14913_));
  XNOR2_X1   g13893(.A1(new_n14830_), .A2(new_n14831_), .ZN(new_n14914_));
  NAND3_X1   g13894(.A1(new_n14870_), .A2(new_n14866_), .A3(new_n14884_), .ZN(new_n14915_));
  NOR4_X1    g13895(.A1(new_n14891_), .A2(new_n14894_), .A3(new_n14904_), .A4(new_n14901_), .ZN(new_n14916_));
  NOR2_X1    g13896(.A1(new_n14895_), .A2(new_n14905_), .ZN(new_n14917_));
  NAND2_X1   g13897(.A1(new_n14914_), .A2(new_n14915_), .ZN(new_n14918_));
  NOR3_X1    g13898(.A1(new_n14829_), .A2(new_n14838_), .A3(new_n14918_), .ZN(new_n14919_));
  NOR2_X1    g13899(.A1(new_n14877_), .A2(new_n14883_), .ZN(new_n14920_));
  INV_X1     g13900(.I(new_n14868_), .ZN(new_n14921_));
  NOR2_X1    g13901(.A1(new_n14920_), .A2(new_n14921_), .ZN(new_n14922_));
  NOR2_X1    g13902(.A1(new_n14866_), .A2(new_n14868_), .ZN(new_n14923_));
  OAI21_X1   g13903(.A1(new_n14922_), .A2(new_n14923_), .B(new_n14867_), .ZN(new_n14924_));
  INV_X1     g13904(.I(new_n14867_), .ZN(new_n14925_));
  NAND2_X1   g13905(.A1(new_n14866_), .A2(new_n14868_), .ZN(new_n14926_));
  NAND2_X1   g13906(.A1(new_n14920_), .A2(new_n14921_), .ZN(new_n14927_));
  NAND3_X1   g13907(.A1(new_n14927_), .A2(new_n14926_), .A3(new_n14925_), .ZN(new_n14928_));
  AND2_X2    g13908(.A1(new_n14924_), .A2(new_n14928_), .Z(new_n14929_));
  NOR3_X1    g13909(.A1(new_n14915_), .A2(new_n14916_), .A3(new_n14917_), .ZN(new_n14930_));
  INV_X1     g13910(.I(new_n14869_), .ZN(new_n14931_));
  NOR2_X1    g13911(.A1(new_n14865_), .A2(new_n14877_), .ZN(new_n14932_));
  NOR2_X1    g13912(.A1(new_n14854_), .A2(new_n14883_), .ZN(new_n14933_));
  OAI21_X1   g13913(.A1(new_n14932_), .A2(new_n14933_), .B(new_n14931_), .ZN(new_n14934_));
  NAND3_X1   g13914(.A1(new_n14934_), .A2(new_n14916_), .A3(new_n14910_), .ZN(new_n14935_));
  AOI21_X1   g13915(.A1(new_n14929_), .A2(new_n14930_), .B(new_n14935_), .ZN(new_n14936_));
  NAND2_X1   g13916(.A1(new_n14895_), .A2(new_n14905_), .ZN(new_n14937_));
  INV_X1     g13917(.I(new_n14909_), .ZN(new_n14938_));
  NAND2_X1   g13918(.A1(new_n14937_), .A2(new_n14938_), .ZN(new_n14939_));
  NAND2_X1   g13919(.A1(new_n14916_), .A2(new_n14909_), .ZN(new_n14940_));
  AOI21_X1   g13920(.A1(new_n14939_), .A2(new_n14940_), .B(new_n14907_), .ZN(new_n14941_));
  INV_X1     g13921(.I(new_n14907_), .ZN(new_n14942_));
  NOR2_X1    g13922(.A1(new_n14916_), .A2(new_n14909_), .ZN(new_n14943_));
  NOR2_X1    g13923(.A1(new_n14937_), .A2(new_n14938_), .ZN(new_n14944_));
  NOR3_X1    g13924(.A1(new_n14944_), .A2(new_n14942_), .A3(new_n14943_), .ZN(new_n14945_));
  OR2_X2     g13925(.A1(new_n14945_), .A2(new_n14941_), .Z(new_n14946_));
  NOR2_X1    g13926(.A1(new_n14917_), .A2(new_n14916_), .ZN(new_n14947_));
  NAND3_X1   g13927(.A1(new_n14947_), .A2(new_n14916_), .A3(new_n14910_), .ZN(new_n14948_));
  NOR2_X1    g13928(.A1(new_n14948_), .A2(new_n14915_), .ZN(new_n14949_));
  INV_X1     g13929(.I(new_n14949_), .ZN(new_n14950_));
  NAND2_X1   g13930(.A1(new_n14950_), .A2(new_n14946_), .ZN(new_n14951_));
  NAND3_X1   g13931(.A1(new_n14924_), .A2(new_n14928_), .A3(new_n14934_), .ZN(new_n14952_));
  NOR4_X1    g13932(.A1(new_n14948_), .A2(new_n14941_), .A3(new_n14945_), .A4(new_n14915_), .ZN(new_n14953_));
  XOR2_X1    g13933(.A1(new_n14953_), .A2(new_n14952_), .Z(new_n14954_));
  AOI22_X1   g13934(.A1(new_n14954_), .A2(new_n14951_), .B1(new_n14936_), .B2(new_n14946_), .ZN(new_n14955_));
  OAI22_X1   g13935(.A1(new_n14913_), .A2(new_n14919_), .B1(new_n14955_), .B2(new_n14839_), .ZN(new_n14956_));
  AOI21_X1   g13936(.A1(new_n14817_), .A2(new_n14832_), .B(new_n14763_), .ZN(new_n14957_));
  INV_X1     g13937(.I(new_n14957_), .ZN(new_n14958_));
  NOR2_X1    g13938(.A1(new_n14768_), .A2(new_n14773_), .ZN(new_n14959_));
  OAI21_X1   g13939(.A1(new_n14811_), .A2(new_n14959_), .B(new_n14776_), .ZN(new_n14960_));
  NOR2_X1    g13940(.A1(new_n14734_), .A2(new_n14739_), .ZN(new_n14961_));
  OAI21_X1   g13941(.A1(new_n14756_), .A2(new_n14961_), .B(new_n14823_), .ZN(new_n14962_));
  XNOR2_X1   g13942(.A1(new_n14960_), .A2(new_n14962_), .ZN(new_n14963_));
  NAND3_X1   g13943(.A1(new_n14958_), .A2(new_n14837_), .A3(new_n14963_), .ZN(new_n14964_));
  NOR2_X1    g13944(.A1(new_n14945_), .A2(new_n14941_), .ZN(new_n14965_));
  AOI21_X1   g13945(.A1(new_n14952_), .A2(new_n14949_), .B(new_n14965_), .ZN(new_n14966_));
  NOR2_X1    g13946(.A1(new_n14867_), .A2(new_n14868_), .ZN(new_n14967_));
  OAI21_X1   g13947(.A1(new_n14866_), .A2(new_n14967_), .B(new_n14869_), .ZN(new_n14968_));
  OAI21_X1   g13948(.A1(new_n14942_), .A2(new_n14938_), .B(new_n14916_), .ZN(new_n14969_));
  OAI21_X1   g13949(.A1(new_n14907_), .A2(new_n14909_), .B(new_n14969_), .ZN(new_n14970_));
  XOR2_X1    g13950(.A1(new_n14970_), .A2(new_n14968_), .Z(new_n14971_));
  NOR3_X1    g13951(.A1(new_n14936_), .A2(new_n14966_), .A3(new_n14971_), .ZN(new_n14972_));
  INV_X1     g13952(.I(new_n14972_), .ZN(new_n14973_));
  NAND2_X1   g13953(.A1(new_n14964_), .A2(new_n14973_), .ZN(new_n14974_));
  INV_X1     g13954(.I(new_n14837_), .ZN(new_n14975_));
  INV_X1     g13955(.I(new_n14963_), .ZN(new_n14976_));
  NOR3_X1    g13956(.A1(new_n14975_), .A2(new_n14957_), .A3(new_n14976_), .ZN(new_n14977_));
  NAND2_X1   g13957(.A1(new_n14977_), .A2(new_n14972_), .ZN(new_n14978_));
  AOI21_X1   g13958(.A1(new_n14956_), .A2(new_n14974_), .B(new_n14978_), .ZN(new_n14979_));
  NAND2_X1   g13959(.A1(new_n14970_), .A2(new_n14968_), .ZN(new_n14980_));
  NOR2_X1    g13960(.A1(new_n14936_), .A2(new_n14966_), .ZN(new_n14981_));
  OAI21_X1   g13961(.A1(new_n14968_), .A2(new_n14970_), .B(new_n14981_), .ZN(new_n14982_));
  NAND2_X1   g13962(.A1(new_n14982_), .A2(new_n14980_), .ZN(new_n14983_));
  INV_X1     g13963(.I(new_n14983_), .ZN(new_n14984_));
  NAND2_X1   g13964(.A1(new_n14960_), .A2(new_n14962_), .ZN(new_n14985_));
  NOR2_X1    g13965(.A1(new_n14975_), .A2(new_n14957_), .ZN(new_n14986_));
  OAI21_X1   g13966(.A1(new_n14960_), .A2(new_n14962_), .B(new_n14986_), .ZN(new_n14987_));
  NAND2_X1   g13967(.A1(new_n14987_), .A2(new_n14985_), .ZN(new_n14988_));
  INV_X1     g13968(.I(new_n14988_), .ZN(new_n14989_));
  AOI21_X1   g13969(.A1(new_n14984_), .A2(new_n14989_), .B(new_n14979_), .ZN(new_n14990_));
  NOR2_X1    g13970(.A1(new_n14989_), .A2(new_n14984_), .ZN(new_n14991_));
  NOR2_X1    g13971(.A1(new_n14990_), .A2(new_n14991_), .ZN(new_n14992_));
  INV_X1     g13972(.I(new_n14992_), .ZN(new_n14993_));
  INV_X1     g13973(.I(\A[622] ), .ZN(new_n14994_));
  NOR2_X1    g13974(.A1(\A[623] ), .A2(\A[624] ), .ZN(new_n14995_));
  NAND2_X1   g13975(.A1(\A[623] ), .A2(\A[624] ), .ZN(new_n14996_));
  AOI21_X1   g13976(.A1(new_n14994_), .A2(new_n14996_), .B(new_n14995_), .ZN(new_n14997_));
  INV_X1     g13977(.I(new_n14997_), .ZN(new_n14998_));
  INV_X1     g13978(.I(\A[619] ), .ZN(new_n14999_));
  NOR2_X1    g13979(.A1(\A[620] ), .A2(\A[621] ), .ZN(new_n15000_));
  INV_X1     g13980(.I(\A[620] ), .ZN(new_n15001_));
  INV_X1     g13981(.I(\A[621] ), .ZN(new_n15002_));
  NOR2_X1    g13982(.A1(new_n15001_), .A2(new_n15002_), .ZN(new_n15003_));
  INV_X1     g13983(.I(new_n15003_), .ZN(new_n15004_));
  AOI21_X1   g13984(.A1(new_n15004_), .A2(new_n14999_), .B(new_n15000_), .ZN(new_n15005_));
  INV_X1     g13985(.I(new_n15005_), .ZN(new_n15006_));
  NAND2_X1   g13986(.A1(new_n15001_), .A2(\A[621] ), .ZN(new_n15007_));
  NAND2_X1   g13987(.A1(new_n15002_), .A2(\A[620] ), .ZN(new_n15008_));
  AOI21_X1   g13988(.A1(new_n15007_), .A2(new_n15008_), .B(new_n14999_), .ZN(new_n15009_));
  NOR2_X1    g13989(.A1(new_n15003_), .A2(new_n15000_), .ZN(new_n15010_));
  NOR2_X1    g13990(.A1(new_n15010_), .A2(\A[619] ), .ZN(new_n15011_));
  INV_X1     g13991(.I(\A[623] ), .ZN(new_n15012_));
  NAND2_X1   g13992(.A1(new_n15012_), .A2(\A[624] ), .ZN(new_n15013_));
  INV_X1     g13993(.I(\A[624] ), .ZN(new_n15014_));
  NAND2_X1   g13994(.A1(new_n15014_), .A2(\A[623] ), .ZN(new_n15015_));
  AOI21_X1   g13995(.A1(new_n15013_), .A2(new_n15015_), .B(new_n14994_), .ZN(new_n15016_));
  INV_X1     g13996(.I(new_n14995_), .ZN(new_n15017_));
  AOI21_X1   g13997(.A1(new_n15017_), .A2(new_n14996_), .B(\A[622] ), .ZN(new_n15018_));
  NOR4_X1    g13998(.A1(new_n15011_), .A2(new_n15009_), .A3(new_n15016_), .A4(new_n15018_), .ZN(new_n15019_));
  NOR2_X1    g13999(.A1(new_n15019_), .A2(new_n15006_), .ZN(new_n15020_));
  INV_X1     g14000(.I(new_n15020_), .ZN(new_n15021_));
  NAND2_X1   g14001(.A1(new_n15019_), .A2(new_n15006_), .ZN(new_n15022_));
  AOI21_X1   g14002(.A1(new_n15021_), .A2(new_n15022_), .B(new_n14998_), .ZN(new_n15023_));
  INV_X1     g14003(.I(new_n15022_), .ZN(new_n15024_));
  NOR3_X1    g14004(.A1(new_n15024_), .A2(new_n14997_), .A3(new_n15020_), .ZN(new_n15025_));
  NOR2_X1    g14005(.A1(new_n15023_), .A2(new_n15025_), .ZN(new_n15026_));
  INV_X1     g14006(.I(new_n15026_), .ZN(new_n15027_));
  INV_X1     g14007(.I(\A[628] ), .ZN(new_n15028_));
  NOR2_X1    g14008(.A1(\A[629] ), .A2(\A[630] ), .ZN(new_n15029_));
  NAND2_X1   g14009(.A1(\A[629] ), .A2(\A[630] ), .ZN(new_n15030_));
  AOI21_X1   g14010(.A1(new_n15028_), .A2(new_n15030_), .B(new_n15029_), .ZN(new_n15031_));
  INV_X1     g14011(.I(new_n15031_), .ZN(new_n15032_));
  INV_X1     g14012(.I(\A[625] ), .ZN(new_n15033_));
  NOR2_X1    g14013(.A1(\A[626] ), .A2(\A[627] ), .ZN(new_n15034_));
  NAND2_X1   g14014(.A1(\A[626] ), .A2(\A[627] ), .ZN(new_n15035_));
  AOI21_X1   g14015(.A1(new_n15033_), .A2(new_n15035_), .B(new_n15034_), .ZN(new_n15036_));
  INV_X1     g14016(.I(new_n15036_), .ZN(new_n15037_));
  NOR2_X1    g14017(.A1(new_n15032_), .A2(new_n15037_), .ZN(new_n15038_));
  INV_X1     g14018(.I(new_n15038_), .ZN(new_n15039_));
  INV_X1     g14019(.I(\A[626] ), .ZN(new_n15040_));
  NAND2_X1   g14020(.A1(new_n15040_), .A2(\A[627] ), .ZN(new_n15041_));
  INV_X1     g14021(.I(\A[627] ), .ZN(new_n15042_));
  NAND2_X1   g14022(.A1(new_n15042_), .A2(\A[626] ), .ZN(new_n15043_));
  AOI21_X1   g14023(.A1(new_n15041_), .A2(new_n15043_), .B(new_n15033_), .ZN(new_n15044_));
  INV_X1     g14024(.I(new_n15034_), .ZN(new_n15045_));
  AOI21_X1   g14025(.A1(new_n15045_), .A2(new_n15035_), .B(\A[625] ), .ZN(new_n15046_));
  NOR2_X1    g14026(.A1(new_n15046_), .A2(new_n15044_), .ZN(new_n15047_));
  INV_X1     g14027(.I(\A[630] ), .ZN(new_n15048_));
  NOR2_X1    g14028(.A1(new_n15048_), .A2(\A[629] ), .ZN(new_n15049_));
  INV_X1     g14029(.I(\A[629] ), .ZN(new_n15050_));
  NOR2_X1    g14030(.A1(new_n15050_), .A2(\A[630] ), .ZN(new_n15051_));
  OAI21_X1   g14031(.A1(new_n15049_), .A2(new_n15051_), .B(\A[628] ), .ZN(new_n15052_));
  INV_X1     g14032(.I(new_n15030_), .ZN(new_n15053_));
  OAI21_X1   g14033(.A1(new_n15053_), .A2(new_n15029_), .B(new_n15028_), .ZN(new_n15054_));
  NAND2_X1   g14034(.A1(new_n15052_), .A2(new_n15054_), .ZN(new_n15055_));
  NAND2_X1   g14035(.A1(new_n15047_), .A2(new_n15055_), .ZN(new_n15056_));
  NOR2_X1    g14036(.A1(new_n15042_), .A2(\A[626] ), .ZN(new_n15057_));
  NOR2_X1    g14037(.A1(new_n15040_), .A2(\A[627] ), .ZN(new_n15058_));
  OAI21_X1   g14038(.A1(new_n15057_), .A2(new_n15058_), .B(\A[625] ), .ZN(new_n15059_));
  INV_X1     g14039(.I(new_n15035_), .ZN(new_n15060_));
  OAI21_X1   g14040(.A1(new_n15060_), .A2(new_n15034_), .B(new_n15033_), .ZN(new_n15061_));
  NAND2_X1   g14041(.A1(new_n15059_), .A2(new_n15061_), .ZN(new_n15062_));
  NAND2_X1   g14042(.A1(new_n15050_), .A2(\A[630] ), .ZN(new_n15063_));
  NAND2_X1   g14043(.A1(new_n15048_), .A2(\A[629] ), .ZN(new_n15064_));
  AOI21_X1   g14044(.A1(new_n15063_), .A2(new_n15064_), .B(new_n15028_), .ZN(new_n15065_));
  INV_X1     g14045(.I(new_n15029_), .ZN(new_n15066_));
  AOI21_X1   g14046(.A1(new_n15066_), .A2(new_n15030_), .B(\A[628] ), .ZN(new_n15067_));
  NOR2_X1    g14047(.A1(new_n15067_), .A2(new_n15065_), .ZN(new_n15068_));
  NAND2_X1   g14048(.A1(new_n15068_), .A2(new_n15062_), .ZN(new_n15069_));
  AOI21_X1   g14049(.A1(new_n15056_), .A2(new_n15069_), .B(new_n15039_), .ZN(new_n15070_));
  INV_X1     g14050(.I(new_n15070_), .ZN(new_n15071_));
  NOR2_X1    g14051(.A1(new_n15062_), .A2(new_n15055_), .ZN(new_n15072_));
  NOR2_X1    g14052(.A1(new_n15072_), .A2(new_n15037_), .ZN(new_n15073_));
  NAND2_X1   g14053(.A1(new_n15047_), .A2(new_n15068_), .ZN(new_n15074_));
  NOR2_X1    g14054(.A1(new_n15074_), .A2(new_n15036_), .ZN(new_n15075_));
  OAI21_X1   g14055(.A1(new_n15073_), .A2(new_n15075_), .B(new_n15031_), .ZN(new_n15076_));
  NAND2_X1   g14056(.A1(new_n15074_), .A2(new_n15036_), .ZN(new_n15077_));
  NAND2_X1   g14057(.A1(new_n15072_), .A2(new_n15037_), .ZN(new_n15078_));
  NAND3_X1   g14058(.A1(new_n15078_), .A2(new_n15077_), .A3(new_n15032_), .ZN(new_n15079_));
  NAND3_X1   g14059(.A1(new_n15076_), .A2(new_n15079_), .A3(new_n15071_), .ZN(new_n15080_));
  NOR2_X1    g14060(.A1(new_n15074_), .A2(new_n15039_), .ZN(new_n15081_));
  NOR2_X1    g14061(.A1(new_n15047_), .A2(new_n15068_), .ZN(new_n15082_));
  NOR2_X1    g14062(.A1(new_n15082_), .A2(new_n15072_), .ZN(new_n15083_));
  NOR2_X1    g14063(.A1(new_n15011_), .A2(new_n15009_), .ZN(new_n15084_));
  NOR2_X1    g14064(.A1(new_n15018_), .A2(new_n15016_), .ZN(new_n15085_));
  NOR2_X1    g14065(.A1(new_n15084_), .A2(new_n15085_), .ZN(new_n15086_));
  NOR2_X1    g14066(.A1(new_n15086_), .A2(new_n15019_), .ZN(new_n15087_));
  INV_X1     g14067(.I(new_n15019_), .ZN(new_n15088_));
  NAND2_X1   g14068(.A1(new_n15005_), .A2(new_n14997_), .ZN(new_n15089_));
  NOR2_X1    g14069(.A1(new_n15088_), .A2(new_n15089_), .ZN(new_n15090_));
  NAND4_X1   g14070(.A1(new_n15090_), .A2(new_n15087_), .A3(new_n15081_), .A4(new_n15083_), .ZN(new_n15091_));
  NOR2_X1    g14071(.A1(new_n15080_), .A2(new_n15091_), .ZN(new_n15092_));
  INV_X1     g14072(.I(new_n15092_), .ZN(new_n15093_));
  NAND2_X1   g14073(.A1(new_n15080_), .A2(new_n15091_), .ZN(new_n15094_));
  AOI21_X1   g14074(.A1(new_n15093_), .A2(new_n15094_), .B(new_n15027_), .ZN(new_n15095_));
  INV_X1     g14075(.I(new_n15091_), .ZN(new_n15096_));
  NAND2_X1   g14076(.A1(new_n15096_), .A2(new_n15080_), .ZN(new_n15097_));
  NAND2_X1   g14077(.A1(new_n15076_), .A2(new_n15079_), .ZN(new_n15098_));
  NAND3_X1   g14078(.A1(new_n15087_), .A2(new_n15081_), .A3(new_n15083_), .ZN(new_n15099_));
  NOR3_X1    g14079(.A1(new_n15070_), .A2(new_n15088_), .A3(new_n15089_), .ZN(new_n15100_));
  OAI21_X1   g14080(.A1(new_n15098_), .A2(new_n15099_), .B(new_n15100_), .ZN(new_n15101_));
  NAND3_X1   g14081(.A1(new_n15097_), .A2(new_n15101_), .A3(new_n15026_), .ZN(new_n15102_));
  INV_X1     g14082(.I(new_n15102_), .ZN(new_n15103_));
  NOR2_X1    g14083(.A1(new_n15103_), .A2(new_n15095_), .ZN(new_n15104_));
  INV_X1     g14084(.I(new_n15094_), .ZN(new_n15105_));
  OAI21_X1   g14085(.A1(new_n15105_), .A2(new_n15092_), .B(new_n15026_), .ZN(new_n15106_));
  NAND2_X1   g14086(.A1(new_n15083_), .A2(new_n15081_), .ZN(new_n15107_));
  NAND2_X1   g14087(.A1(new_n15090_), .A2(new_n15087_), .ZN(new_n15108_));
  XOR2_X1    g14088(.A1(new_n15108_), .A2(new_n15107_), .Z(new_n15109_));
  INV_X1     g14089(.I(\A[613] ), .ZN(new_n15110_));
  INV_X1     g14090(.I(\A[614] ), .ZN(new_n15111_));
  NAND2_X1   g14091(.A1(new_n15111_), .A2(\A[615] ), .ZN(new_n15112_));
  INV_X1     g14092(.I(\A[615] ), .ZN(new_n15113_));
  NAND2_X1   g14093(.A1(new_n15113_), .A2(\A[614] ), .ZN(new_n15114_));
  AOI21_X1   g14094(.A1(new_n15112_), .A2(new_n15114_), .B(new_n15110_), .ZN(new_n15115_));
  NOR2_X1    g14095(.A1(\A[614] ), .A2(\A[615] ), .ZN(new_n15116_));
  INV_X1     g14096(.I(new_n15116_), .ZN(new_n15117_));
  NAND2_X1   g14097(.A1(\A[614] ), .A2(\A[615] ), .ZN(new_n15118_));
  AOI21_X1   g14098(.A1(new_n15117_), .A2(new_n15118_), .B(\A[613] ), .ZN(new_n15119_));
  NOR2_X1    g14099(.A1(new_n15119_), .A2(new_n15115_), .ZN(new_n15120_));
  INV_X1     g14100(.I(\A[616] ), .ZN(new_n15121_));
  INV_X1     g14101(.I(\A[617] ), .ZN(new_n15122_));
  NAND2_X1   g14102(.A1(new_n15122_), .A2(\A[618] ), .ZN(new_n15123_));
  INV_X1     g14103(.I(\A[618] ), .ZN(new_n15124_));
  NAND2_X1   g14104(.A1(new_n15124_), .A2(\A[617] ), .ZN(new_n15125_));
  AOI21_X1   g14105(.A1(new_n15123_), .A2(new_n15125_), .B(new_n15121_), .ZN(new_n15126_));
  NOR2_X1    g14106(.A1(\A[617] ), .A2(\A[618] ), .ZN(new_n15127_));
  INV_X1     g14107(.I(new_n15127_), .ZN(new_n15128_));
  NAND2_X1   g14108(.A1(\A[617] ), .A2(\A[618] ), .ZN(new_n15129_));
  AOI21_X1   g14109(.A1(new_n15128_), .A2(new_n15129_), .B(\A[616] ), .ZN(new_n15130_));
  NOR2_X1    g14110(.A1(new_n15130_), .A2(new_n15126_), .ZN(new_n15131_));
  NAND2_X1   g14111(.A1(new_n15120_), .A2(new_n15131_), .ZN(new_n15132_));
  AOI21_X1   g14112(.A1(new_n15121_), .A2(new_n15129_), .B(new_n15127_), .ZN(new_n15133_));
  INV_X1     g14113(.I(new_n15133_), .ZN(new_n15134_));
  AOI21_X1   g14114(.A1(new_n15110_), .A2(new_n15118_), .B(new_n15116_), .ZN(new_n15135_));
  INV_X1     g14115(.I(new_n15135_), .ZN(new_n15136_));
  NOR2_X1    g14116(.A1(new_n15134_), .A2(new_n15136_), .ZN(new_n15137_));
  INV_X1     g14117(.I(new_n15137_), .ZN(new_n15138_));
  NOR2_X1    g14118(.A1(new_n15132_), .A2(new_n15138_), .ZN(new_n15139_));
  INV_X1     g14119(.I(new_n15139_), .ZN(new_n15140_));
  NOR2_X1    g14120(.A1(new_n15113_), .A2(\A[614] ), .ZN(new_n15141_));
  NOR2_X1    g14121(.A1(new_n15111_), .A2(\A[615] ), .ZN(new_n15142_));
  OAI21_X1   g14122(.A1(new_n15141_), .A2(new_n15142_), .B(\A[613] ), .ZN(new_n15143_));
  INV_X1     g14123(.I(new_n15118_), .ZN(new_n15144_));
  OAI21_X1   g14124(.A1(new_n15144_), .A2(new_n15116_), .B(new_n15110_), .ZN(new_n15145_));
  NAND2_X1   g14125(.A1(new_n15143_), .A2(new_n15145_), .ZN(new_n15146_));
  NOR2_X1    g14126(.A1(new_n15124_), .A2(\A[617] ), .ZN(new_n15147_));
  NOR2_X1    g14127(.A1(new_n15122_), .A2(\A[618] ), .ZN(new_n15148_));
  OAI21_X1   g14128(.A1(new_n15147_), .A2(new_n15148_), .B(\A[616] ), .ZN(new_n15149_));
  INV_X1     g14129(.I(new_n15129_), .ZN(new_n15150_));
  OAI21_X1   g14130(.A1(new_n15150_), .A2(new_n15127_), .B(new_n15121_), .ZN(new_n15151_));
  NAND2_X1   g14131(.A1(new_n15149_), .A2(new_n15151_), .ZN(new_n15152_));
  NAND2_X1   g14132(.A1(new_n15146_), .A2(new_n15152_), .ZN(new_n15153_));
  NAND2_X1   g14133(.A1(new_n15132_), .A2(new_n15153_), .ZN(new_n15154_));
  INV_X1     g14134(.I(\A[607] ), .ZN(new_n15155_));
  INV_X1     g14135(.I(\A[608] ), .ZN(new_n15156_));
  NAND2_X1   g14136(.A1(new_n15156_), .A2(\A[609] ), .ZN(new_n15157_));
  INV_X1     g14137(.I(\A[609] ), .ZN(new_n15158_));
  NAND2_X1   g14138(.A1(new_n15158_), .A2(\A[608] ), .ZN(new_n15159_));
  AOI21_X1   g14139(.A1(new_n15157_), .A2(new_n15159_), .B(new_n15155_), .ZN(new_n15160_));
  NAND2_X1   g14140(.A1(new_n15156_), .A2(new_n15158_), .ZN(new_n15161_));
  NAND2_X1   g14141(.A1(\A[608] ), .A2(\A[609] ), .ZN(new_n15162_));
  AOI21_X1   g14142(.A1(new_n15161_), .A2(new_n15162_), .B(\A[607] ), .ZN(new_n15163_));
  NOR2_X1    g14143(.A1(new_n15163_), .A2(new_n15160_), .ZN(new_n15164_));
  INV_X1     g14144(.I(\A[610] ), .ZN(new_n15165_));
  INV_X1     g14145(.I(\A[611] ), .ZN(new_n15166_));
  NAND2_X1   g14146(.A1(new_n15166_), .A2(\A[612] ), .ZN(new_n15167_));
  INV_X1     g14147(.I(\A[612] ), .ZN(new_n15168_));
  NAND2_X1   g14148(.A1(new_n15168_), .A2(\A[611] ), .ZN(new_n15169_));
  AOI21_X1   g14149(.A1(new_n15167_), .A2(new_n15169_), .B(new_n15165_), .ZN(new_n15170_));
  NAND2_X1   g14150(.A1(new_n15166_), .A2(new_n15168_), .ZN(new_n15171_));
  NAND2_X1   g14151(.A1(\A[611] ), .A2(\A[612] ), .ZN(new_n15172_));
  AOI21_X1   g14152(.A1(new_n15171_), .A2(new_n15172_), .B(\A[610] ), .ZN(new_n15173_));
  NOR2_X1    g14153(.A1(new_n15173_), .A2(new_n15170_), .ZN(new_n15174_));
  NAND2_X1   g14154(.A1(new_n15172_), .A2(new_n15165_), .ZN(new_n15175_));
  NAND2_X1   g14155(.A1(new_n15175_), .A2(new_n15171_), .ZN(new_n15176_));
  NAND2_X1   g14156(.A1(new_n15162_), .A2(new_n15155_), .ZN(new_n15177_));
  NAND2_X1   g14157(.A1(new_n15177_), .A2(new_n15161_), .ZN(new_n15178_));
  NOR2_X1    g14158(.A1(new_n15176_), .A2(new_n15178_), .ZN(new_n15179_));
  NOR2_X1    g14159(.A1(new_n15140_), .A2(new_n15154_), .ZN(new_n15180_));
  NOR2_X1    g14160(.A1(new_n15109_), .A2(new_n15180_), .ZN(new_n15181_));
  AOI21_X1   g14161(.A1(new_n15106_), .A2(new_n15102_), .B(new_n15181_), .ZN(new_n15182_));
  XNOR2_X1   g14162(.A1(new_n15108_), .A2(new_n15107_), .ZN(new_n15183_));
  NAND3_X1   g14163(.A1(new_n15139_), .A2(new_n15132_), .A3(new_n15153_), .ZN(new_n15184_));
  NOR4_X1    g14164(.A1(new_n15160_), .A2(new_n15163_), .A3(new_n15173_), .A4(new_n15170_), .ZN(new_n15185_));
  NOR2_X1    g14165(.A1(new_n15164_), .A2(new_n15174_), .ZN(new_n15186_));
  NAND2_X1   g14166(.A1(new_n15183_), .A2(new_n15184_), .ZN(new_n15187_));
  NOR3_X1    g14167(.A1(new_n15103_), .A2(new_n15095_), .A3(new_n15187_), .ZN(new_n15188_));
  NOR2_X1    g14168(.A1(new_n15146_), .A2(new_n15152_), .ZN(new_n15189_));
  NOR2_X1    g14169(.A1(new_n15189_), .A2(new_n15136_), .ZN(new_n15190_));
  NOR2_X1    g14170(.A1(new_n15132_), .A2(new_n15135_), .ZN(new_n15191_));
  OAI21_X1   g14171(.A1(new_n15190_), .A2(new_n15191_), .B(new_n15133_), .ZN(new_n15192_));
  NAND2_X1   g14172(.A1(new_n15132_), .A2(new_n15135_), .ZN(new_n15193_));
  NAND2_X1   g14173(.A1(new_n15189_), .A2(new_n15136_), .ZN(new_n15194_));
  NAND3_X1   g14174(.A1(new_n15194_), .A2(new_n15193_), .A3(new_n15134_), .ZN(new_n15195_));
  AND2_X2    g14175(.A1(new_n15192_), .A2(new_n15195_), .Z(new_n15196_));
  NOR3_X1    g14176(.A1(new_n15184_), .A2(new_n15185_), .A3(new_n15186_), .ZN(new_n15197_));
  NAND2_X1   g14177(.A1(new_n15164_), .A2(new_n15174_), .ZN(new_n15198_));
  INV_X1     g14178(.I(new_n15179_), .ZN(new_n15199_));
  NOR2_X1    g14179(.A1(new_n15198_), .A2(new_n15199_), .ZN(new_n15200_));
  NOR2_X1    g14180(.A1(new_n15131_), .A2(new_n15146_), .ZN(new_n15201_));
  NOR2_X1    g14181(.A1(new_n15120_), .A2(new_n15152_), .ZN(new_n15202_));
  OAI21_X1   g14182(.A1(new_n15201_), .A2(new_n15202_), .B(new_n15137_), .ZN(new_n15203_));
  NAND2_X1   g14183(.A1(new_n15203_), .A2(new_n15200_), .ZN(new_n15204_));
  AOI21_X1   g14184(.A1(new_n15196_), .A2(new_n15197_), .B(new_n15204_), .ZN(new_n15205_));
  NOR2_X1    g14185(.A1(new_n15185_), .A2(new_n15178_), .ZN(new_n15206_));
  INV_X1     g14186(.I(new_n15206_), .ZN(new_n15207_));
  NAND2_X1   g14187(.A1(new_n15185_), .A2(new_n15178_), .ZN(new_n15208_));
  AOI21_X1   g14188(.A1(new_n15207_), .A2(new_n15208_), .B(new_n15176_), .ZN(new_n15209_));
  INV_X1     g14189(.I(new_n15176_), .ZN(new_n15210_));
  INV_X1     g14190(.I(new_n15208_), .ZN(new_n15211_));
  NOR3_X1    g14191(.A1(new_n15211_), .A2(new_n15210_), .A3(new_n15206_), .ZN(new_n15212_));
  NOR2_X1    g14192(.A1(new_n15209_), .A2(new_n15212_), .ZN(new_n15213_));
  INV_X1     g14193(.I(new_n15213_), .ZN(new_n15214_));
  NOR2_X1    g14194(.A1(new_n15186_), .A2(new_n15185_), .ZN(new_n15215_));
  NAND2_X1   g14195(.A1(new_n15215_), .A2(new_n15200_), .ZN(new_n15216_));
  NOR2_X1    g14196(.A1(new_n15184_), .A2(new_n15216_), .ZN(new_n15217_));
  INV_X1     g14197(.I(new_n15217_), .ZN(new_n15218_));
  NAND2_X1   g14198(.A1(new_n15214_), .A2(new_n15218_), .ZN(new_n15219_));
  NAND3_X1   g14199(.A1(new_n15192_), .A2(new_n15195_), .A3(new_n15203_), .ZN(new_n15220_));
  NOR4_X1    g14200(.A1(new_n15209_), .A2(new_n15212_), .A3(new_n15184_), .A4(new_n15216_), .ZN(new_n15221_));
  XOR2_X1    g14201(.A1(new_n15221_), .A2(new_n15220_), .Z(new_n15222_));
  AOI22_X1   g14202(.A1(new_n15222_), .A2(new_n15219_), .B1(new_n15205_), .B2(new_n15214_), .ZN(new_n15223_));
  OAI22_X1   g14203(.A1(new_n15182_), .A2(new_n15188_), .B1(new_n15223_), .B2(new_n15104_), .ZN(new_n15224_));
  NAND2_X1   g14204(.A1(new_n15027_), .A2(new_n15097_), .ZN(new_n15225_));
  NOR2_X1    g14205(.A1(new_n15031_), .A2(new_n15036_), .ZN(new_n15226_));
  OAI21_X1   g14206(.A1(new_n15074_), .A2(new_n15226_), .B(new_n15039_), .ZN(new_n15227_));
  NOR2_X1    g14207(.A1(new_n15005_), .A2(new_n14997_), .ZN(new_n15228_));
  OAI21_X1   g14208(.A1(new_n15088_), .A2(new_n15228_), .B(new_n15089_), .ZN(new_n15229_));
  XNOR2_X1   g14209(.A1(new_n15229_), .A2(new_n15227_), .ZN(new_n15230_));
  NAND3_X1   g14210(.A1(new_n15225_), .A2(new_n15101_), .A3(new_n15230_), .ZN(new_n15231_));
  AOI21_X1   g14211(.A1(new_n15220_), .A2(new_n15217_), .B(new_n15213_), .ZN(new_n15232_));
  NOR2_X1    g14212(.A1(new_n15133_), .A2(new_n15135_), .ZN(new_n15233_));
  OAI21_X1   g14213(.A1(new_n15132_), .A2(new_n15233_), .B(new_n15138_), .ZN(new_n15234_));
  AOI21_X1   g14214(.A1(new_n15161_), .A2(new_n15177_), .B(new_n15210_), .ZN(new_n15235_));
  OAI21_X1   g14215(.A1(new_n15198_), .A2(new_n15235_), .B(new_n15199_), .ZN(new_n15236_));
  XOR2_X1    g14216(.A1(new_n15234_), .A2(new_n15236_), .Z(new_n15237_));
  NOR3_X1    g14217(.A1(new_n15205_), .A2(new_n15232_), .A3(new_n15237_), .ZN(new_n15238_));
  INV_X1     g14218(.I(new_n15238_), .ZN(new_n15239_));
  NAND2_X1   g14219(.A1(new_n15239_), .A2(new_n15231_), .ZN(new_n15240_));
  INV_X1     g14220(.I(new_n15231_), .ZN(new_n15241_));
  NAND2_X1   g14221(.A1(new_n15241_), .A2(new_n15238_), .ZN(new_n15242_));
  AOI21_X1   g14222(.A1(new_n15224_), .A2(new_n15240_), .B(new_n15242_), .ZN(new_n15243_));
  NAND2_X1   g14223(.A1(new_n15234_), .A2(new_n15236_), .ZN(new_n15244_));
  NOR2_X1    g14224(.A1(new_n15205_), .A2(new_n15232_), .ZN(new_n15245_));
  OAI21_X1   g14225(.A1(new_n15234_), .A2(new_n15236_), .B(new_n15245_), .ZN(new_n15246_));
  NAND2_X1   g14226(.A1(new_n15246_), .A2(new_n15244_), .ZN(new_n15247_));
  INV_X1     g14227(.I(new_n15247_), .ZN(new_n15248_));
  NAND2_X1   g14228(.A1(new_n15229_), .A2(new_n15227_), .ZN(new_n15249_));
  OR2_X2     g14229(.A1(new_n15229_), .A2(new_n15227_), .Z(new_n15250_));
  NAND3_X1   g14230(.A1(new_n15225_), .A2(new_n15101_), .A3(new_n15250_), .ZN(new_n15251_));
  NAND2_X1   g14231(.A1(new_n15251_), .A2(new_n15249_), .ZN(new_n15252_));
  INV_X1     g14232(.I(new_n15252_), .ZN(new_n15253_));
  AOI21_X1   g14233(.A1(new_n15248_), .A2(new_n15253_), .B(new_n15243_), .ZN(new_n15254_));
  NOR2_X1    g14234(.A1(new_n15248_), .A2(new_n15253_), .ZN(new_n15255_));
  NOR2_X1    g14235(.A1(new_n15254_), .A2(new_n15255_), .ZN(new_n15256_));
  INV_X1     g14236(.I(new_n15256_), .ZN(new_n15257_));
  NAND2_X1   g14237(.A1(new_n15257_), .A2(new_n14993_), .ZN(new_n15258_));
  XOR2_X1    g14238(.A1(new_n15231_), .A2(new_n15238_), .Z(new_n15259_));
  NOR2_X1    g14239(.A1(new_n15259_), .A2(new_n15224_), .ZN(new_n15260_));
  NAND2_X1   g14240(.A1(new_n15106_), .A2(new_n15102_), .ZN(new_n15261_));
  OAI21_X1   g14241(.A1(new_n15103_), .A2(new_n15095_), .B(new_n15187_), .ZN(new_n15262_));
  NAND3_X1   g14242(.A1(new_n15106_), .A2(new_n15102_), .A3(new_n15181_), .ZN(new_n15263_));
  NAND2_X1   g14243(.A1(new_n15205_), .A2(new_n15214_), .ZN(new_n15264_));
  AOI21_X1   g14244(.A1(new_n15196_), .A2(new_n15203_), .B(new_n15221_), .ZN(new_n15265_));
  NOR3_X1    g14245(.A1(new_n15214_), .A2(new_n15218_), .A3(new_n15220_), .ZN(new_n15266_));
  OAI21_X1   g14246(.A1(new_n15266_), .A2(new_n15265_), .B(new_n15219_), .ZN(new_n15267_));
  NAND2_X1   g14247(.A1(new_n15267_), .A2(new_n15264_), .ZN(new_n15268_));
  AOI22_X1   g14248(.A1(new_n15262_), .A2(new_n15263_), .B1(new_n15268_), .B2(new_n15261_), .ZN(new_n15269_));
  AOI21_X1   g14249(.A1(new_n15240_), .A2(new_n15242_), .B(new_n15269_), .ZN(new_n15270_));
  NAND2_X1   g14250(.A1(new_n14841_), .A2(new_n14842_), .ZN(new_n15271_));
  OAI21_X1   g14251(.A1(new_n14829_), .A2(new_n14838_), .B(new_n14918_), .ZN(new_n15272_));
  NAND3_X1   g14252(.A1(new_n14841_), .A2(new_n14842_), .A3(new_n14912_), .ZN(new_n15273_));
  NAND2_X1   g14253(.A1(new_n14936_), .A2(new_n14946_), .ZN(new_n15274_));
  AOI21_X1   g14254(.A1(new_n14929_), .A2(new_n14934_), .B(new_n14953_), .ZN(new_n15275_));
  NOR3_X1    g14255(.A1(new_n14950_), .A2(new_n14946_), .A3(new_n14952_), .ZN(new_n15276_));
  OAI21_X1   g14256(.A1(new_n15275_), .A2(new_n15276_), .B(new_n14951_), .ZN(new_n15277_));
  NAND2_X1   g14257(.A1(new_n15277_), .A2(new_n15274_), .ZN(new_n15278_));
  AOI22_X1   g14258(.A1(new_n15272_), .A2(new_n15273_), .B1(new_n15278_), .B2(new_n15271_), .ZN(new_n15279_));
  XOR2_X1    g14259(.A1(new_n14977_), .A2(new_n14972_), .Z(new_n15280_));
  NAND2_X1   g14260(.A1(new_n15279_), .A2(new_n15280_), .ZN(new_n15281_));
  NAND2_X1   g14261(.A1(new_n14974_), .A2(new_n14978_), .ZN(new_n15282_));
  NAND2_X1   g14262(.A1(new_n14956_), .A2(new_n15282_), .ZN(new_n15283_));
  NAND2_X1   g14263(.A1(new_n15283_), .A2(new_n15281_), .ZN(new_n15284_));
  NOR3_X1    g14264(.A1(new_n15284_), .A2(new_n15260_), .A3(new_n15270_), .ZN(new_n15285_));
  NOR3_X1    g14265(.A1(new_n14919_), .A2(new_n14913_), .A3(new_n15278_), .ZN(new_n15286_));
  INV_X1     g14266(.I(new_n15286_), .ZN(new_n15287_));
  NAND2_X1   g14267(.A1(new_n14843_), .A2(new_n14911_), .ZN(new_n15288_));
  NAND2_X1   g14268(.A1(new_n14918_), .A2(new_n15288_), .ZN(new_n15289_));
  NAND2_X1   g14269(.A1(new_n15109_), .A2(new_n15180_), .ZN(new_n15290_));
  NAND2_X1   g14270(.A1(new_n15187_), .A2(new_n15290_), .ZN(new_n15291_));
  NOR2_X1    g14271(.A1(new_n15291_), .A2(new_n15289_), .ZN(new_n15292_));
  NOR2_X1    g14272(.A1(new_n15286_), .A2(new_n15292_), .ZN(new_n15293_));
  INV_X1     g14273(.I(new_n15293_), .ZN(new_n15294_));
  NAND2_X1   g14274(.A1(new_n15286_), .A2(new_n15292_), .ZN(new_n15295_));
  OAI21_X1   g14275(.A1(new_n15188_), .A2(new_n15182_), .B(new_n15223_), .ZN(new_n15296_));
  NAND3_X1   g14276(.A1(new_n15262_), .A2(new_n15268_), .A3(new_n15263_), .ZN(new_n15297_));
  NAND2_X1   g14277(.A1(new_n15296_), .A2(new_n15297_), .ZN(new_n15298_));
  AOI22_X1   g14278(.A1(new_n15294_), .A2(new_n15295_), .B1(new_n15287_), .B2(new_n15298_), .ZN(new_n15299_));
  XNOR2_X1   g14279(.A1(new_n15231_), .A2(new_n15238_), .ZN(new_n15300_));
  NAND2_X1   g14280(.A1(new_n15300_), .A2(new_n15269_), .ZN(new_n15301_));
  NAND2_X1   g14281(.A1(new_n15242_), .A2(new_n15240_), .ZN(new_n15302_));
  NAND2_X1   g14282(.A1(new_n15302_), .A2(new_n15224_), .ZN(new_n15303_));
  NAND2_X1   g14283(.A1(new_n15303_), .A2(new_n15301_), .ZN(new_n15304_));
  NAND2_X1   g14284(.A1(new_n15304_), .A2(new_n15284_), .ZN(new_n15305_));
  AOI21_X1   g14285(.A1(new_n15305_), .A2(new_n15299_), .B(new_n15285_), .ZN(new_n15306_));
  NOR2_X1    g14286(.A1(new_n15243_), .A2(new_n15248_), .ZN(new_n15307_));
  NAND4_X1   g14287(.A1(new_n15248_), .A2(new_n15269_), .A3(new_n15241_), .A4(new_n15238_), .ZN(new_n15308_));
  INV_X1     g14288(.I(new_n15308_), .ZN(new_n15309_));
  OAI21_X1   g14289(.A1(new_n15307_), .A2(new_n15309_), .B(new_n15252_), .ZN(new_n15310_));
  NAND3_X1   g14290(.A1(new_n15269_), .A2(new_n15241_), .A3(new_n15238_), .ZN(new_n15311_));
  NAND2_X1   g14291(.A1(new_n15311_), .A2(new_n15247_), .ZN(new_n15312_));
  NAND3_X1   g14292(.A1(new_n15312_), .A2(new_n15253_), .A3(new_n15308_), .ZN(new_n15313_));
  NOR2_X1    g14293(.A1(new_n14979_), .A2(new_n14984_), .ZN(new_n15314_));
  NAND4_X1   g14294(.A1(new_n14984_), .A2(new_n15279_), .A3(new_n14977_), .A4(new_n14972_), .ZN(new_n15315_));
  INV_X1     g14295(.I(new_n15315_), .ZN(new_n15316_));
  OAI21_X1   g14296(.A1(new_n15314_), .A2(new_n15316_), .B(new_n14988_), .ZN(new_n15317_));
  NAND3_X1   g14297(.A1(new_n15279_), .A2(new_n14977_), .A3(new_n14972_), .ZN(new_n15318_));
  NAND2_X1   g14298(.A1(new_n15318_), .A2(new_n14983_), .ZN(new_n15319_));
  NAND3_X1   g14299(.A1(new_n15319_), .A2(new_n14989_), .A3(new_n15315_), .ZN(new_n15320_));
  NAND4_X1   g14300(.A1(new_n15310_), .A2(new_n15317_), .A3(new_n15313_), .A4(new_n15320_), .ZN(new_n15321_));
  NAND2_X1   g14301(.A1(new_n15321_), .A2(new_n15306_), .ZN(new_n15322_));
  XOR2_X1    g14302(.A1(new_n14988_), .A2(new_n14983_), .Z(new_n15323_));
  XOR2_X1    g14303(.A1(new_n15247_), .A2(new_n15252_), .Z(new_n15324_));
  NOR4_X1    g14304(.A1(new_n15323_), .A2(new_n15324_), .A3(new_n15318_), .A4(new_n15311_), .ZN(new_n15325_));
  NAND2_X1   g14305(.A1(new_n15322_), .A2(new_n15325_), .ZN(new_n15326_));
  NOR4_X1    g14306(.A1(new_n15254_), .A2(new_n14990_), .A3(new_n14991_), .A4(new_n15255_), .ZN(new_n15327_));
  NAND2_X1   g14307(.A1(new_n15326_), .A2(new_n15327_), .ZN(new_n15328_));
  NAND2_X1   g14308(.A1(new_n15328_), .A2(new_n15258_), .ZN(new_n15329_));
  INV_X1     g14309(.I(\A[598] ), .ZN(new_n15330_));
  NOR2_X1    g14310(.A1(\A[599] ), .A2(\A[600] ), .ZN(new_n15331_));
  NAND2_X1   g14311(.A1(\A[599] ), .A2(\A[600] ), .ZN(new_n15332_));
  AOI21_X1   g14312(.A1(new_n15330_), .A2(new_n15332_), .B(new_n15331_), .ZN(new_n15333_));
  INV_X1     g14313(.I(new_n15333_), .ZN(new_n15334_));
  INV_X1     g14314(.I(\A[595] ), .ZN(new_n15335_));
  NOR2_X1    g14315(.A1(\A[596] ), .A2(\A[597] ), .ZN(new_n15336_));
  NAND2_X1   g14316(.A1(\A[596] ), .A2(\A[597] ), .ZN(new_n15337_));
  AOI21_X1   g14317(.A1(new_n15335_), .A2(new_n15337_), .B(new_n15336_), .ZN(new_n15338_));
  INV_X1     g14318(.I(new_n15338_), .ZN(new_n15339_));
  INV_X1     g14319(.I(\A[596] ), .ZN(new_n15340_));
  NAND2_X1   g14320(.A1(new_n15340_), .A2(\A[597] ), .ZN(new_n15341_));
  INV_X1     g14321(.I(\A[597] ), .ZN(new_n15342_));
  NAND2_X1   g14322(.A1(new_n15342_), .A2(\A[596] ), .ZN(new_n15343_));
  AOI21_X1   g14323(.A1(new_n15341_), .A2(new_n15343_), .B(new_n15335_), .ZN(new_n15344_));
  INV_X1     g14324(.I(new_n15336_), .ZN(new_n15345_));
  AOI21_X1   g14325(.A1(new_n15345_), .A2(new_n15337_), .B(\A[595] ), .ZN(new_n15346_));
  INV_X1     g14326(.I(\A[599] ), .ZN(new_n15347_));
  NAND2_X1   g14327(.A1(new_n15347_), .A2(\A[600] ), .ZN(new_n15348_));
  INV_X1     g14328(.I(\A[600] ), .ZN(new_n15349_));
  NAND2_X1   g14329(.A1(new_n15349_), .A2(\A[599] ), .ZN(new_n15350_));
  AOI21_X1   g14330(.A1(new_n15348_), .A2(new_n15350_), .B(new_n15330_), .ZN(new_n15351_));
  INV_X1     g14331(.I(new_n15331_), .ZN(new_n15352_));
  AOI21_X1   g14332(.A1(new_n15352_), .A2(new_n15332_), .B(\A[598] ), .ZN(new_n15353_));
  NOR4_X1    g14333(.A1(new_n15344_), .A2(new_n15346_), .A3(new_n15353_), .A4(new_n15351_), .ZN(new_n15354_));
  NOR2_X1    g14334(.A1(new_n15354_), .A2(new_n15339_), .ZN(new_n15355_));
  INV_X1     g14335(.I(new_n15355_), .ZN(new_n15356_));
  NAND2_X1   g14336(.A1(new_n15354_), .A2(new_n15339_), .ZN(new_n15357_));
  AOI21_X1   g14337(.A1(new_n15356_), .A2(new_n15357_), .B(new_n15334_), .ZN(new_n15358_));
  INV_X1     g14338(.I(new_n15357_), .ZN(new_n15359_));
  NOR3_X1    g14339(.A1(new_n15359_), .A2(new_n15333_), .A3(new_n15355_), .ZN(new_n15360_));
  NOR2_X1    g14340(.A1(new_n15358_), .A2(new_n15360_), .ZN(new_n15361_));
  INV_X1     g14341(.I(\A[604] ), .ZN(new_n15362_));
  NOR2_X1    g14342(.A1(\A[605] ), .A2(\A[606] ), .ZN(new_n15363_));
  NAND2_X1   g14343(.A1(\A[605] ), .A2(\A[606] ), .ZN(new_n15364_));
  AOI21_X1   g14344(.A1(new_n15362_), .A2(new_n15364_), .B(new_n15363_), .ZN(new_n15365_));
  INV_X1     g14345(.I(new_n15365_), .ZN(new_n15366_));
  INV_X1     g14346(.I(\A[601] ), .ZN(new_n15367_));
  NOR2_X1    g14347(.A1(\A[602] ), .A2(\A[603] ), .ZN(new_n15368_));
  NAND2_X1   g14348(.A1(\A[602] ), .A2(\A[603] ), .ZN(new_n15369_));
  AOI21_X1   g14349(.A1(new_n15367_), .A2(new_n15369_), .B(new_n15368_), .ZN(new_n15370_));
  INV_X1     g14350(.I(new_n15370_), .ZN(new_n15371_));
  NOR2_X1    g14351(.A1(new_n15366_), .A2(new_n15371_), .ZN(new_n15372_));
  INV_X1     g14352(.I(new_n15372_), .ZN(new_n15373_));
  INV_X1     g14353(.I(\A[602] ), .ZN(new_n15374_));
  NAND2_X1   g14354(.A1(new_n15374_), .A2(\A[603] ), .ZN(new_n15375_));
  INV_X1     g14355(.I(\A[603] ), .ZN(new_n15376_));
  NAND2_X1   g14356(.A1(new_n15376_), .A2(\A[602] ), .ZN(new_n15377_));
  AOI21_X1   g14357(.A1(new_n15375_), .A2(new_n15377_), .B(new_n15367_), .ZN(new_n15378_));
  INV_X1     g14358(.I(new_n15368_), .ZN(new_n15379_));
  AOI21_X1   g14359(.A1(new_n15379_), .A2(new_n15369_), .B(\A[601] ), .ZN(new_n15380_));
  NOR2_X1    g14360(.A1(new_n15380_), .A2(new_n15378_), .ZN(new_n15381_));
  INV_X1     g14361(.I(\A[606] ), .ZN(new_n15382_));
  NOR2_X1    g14362(.A1(new_n15382_), .A2(\A[605] ), .ZN(new_n15383_));
  INV_X1     g14363(.I(\A[605] ), .ZN(new_n15384_));
  NOR2_X1    g14364(.A1(new_n15384_), .A2(\A[606] ), .ZN(new_n15385_));
  OAI21_X1   g14365(.A1(new_n15383_), .A2(new_n15385_), .B(\A[604] ), .ZN(new_n15386_));
  INV_X1     g14366(.I(new_n15364_), .ZN(new_n15387_));
  OAI21_X1   g14367(.A1(new_n15387_), .A2(new_n15363_), .B(new_n15362_), .ZN(new_n15388_));
  NAND2_X1   g14368(.A1(new_n15386_), .A2(new_n15388_), .ZN(new_n15389_));
  NAND2_X1   g14369(.A1(new_n15381_), .A2(new_n15389_), .ZN(new_n15390_));
  NOR2_X1    g14370(.A1(new_n15376_), .A2(\A[602] ), .ZN(new_n15391_));
  NOR2_X1    g14371(.A1(new_n15374_), .A2(\A[603] ), .ZN(new_n15392_));
  OAI21_X1   g14372(.A1(new_n15391_), .A2(new_n15392_), .B(\A[601] ), .ZN(new_n15393_));
  INV_X1     g14373(.I(new_n15369_), .ZN(new_n15394_));
  OAI21_X1   g14374(.A1(new_n15394_), .A2(new_n15368_), .B(new_n15367_), .ZN(new_n15395_));
  NAND2_X1   g14375(.A1(new_n15393_), .A2(new_n15395_), .ZN(new_n15396_));
  NAND2_X1   g14376(.A1(new_n15384_), .A2(\A[606] ), .ZN(new_n15397_));
  NAND2_X1   g14377(.A1(new_n15382_), .A2(\A[605] ), .ZN(new_n15398_));
  AOI21_X1   g14378(.A1(new_n15397_), .A2(new_n15398_), .B(new_n15362_), .ZN(new_n15399_));
  INV_X1     g14379(.I(new_n15363_), .ZN(new_n15400_));
  AOI21_X1   g14380(.A1(new_n15400_), .A2(new_n15364_), .B(\A[604] ), .ZN(new_n15401_));
  NOR2_X1    g14381(.A1(new_n15401_), .A2(new_n15399_), .ZN(new_n15402_));
  NAND2_X1   g14382(.A1(new_n15402_), .A2(new_n15396_), .ZN(new_n15403_));
  AOI21_X1   g14383(.A1(new_n15390_), .A2(new_n15403_), .B(new_n15373_), .ZN(new_n15404_));
  INV_X1     g14384(.I(new_n15404_), .ZN(new_n15405_));
  NOR2_X1    g14385(.A1(new_n15396_), .A2(new_n15389_), .ZN(new_n15406_));
  NOR2_X1    g14386(.A1(new_n15406_), .A2(new_n15371_), .ZN(new_n15407_));
  NAND2_X1   g14387(.A1(new_n15381_), .A2(new_n15402_), .ZN(new_n15408_));
  NOR2_X1    g14388(.A1(new_n15408_), .A2(new_n15370_), .ZN(new_n15409_));
  OAI21_X1   g14389(.A1(new_n15407_), .A2(new_n15409_), .B(new_n15365_), .ZN(new_n15410_));
  NAND2_X1   g14390(.A1(new_n15408_), .A2(new_n15370_), .ZN(new_n15411_));
  NAND2_X1   g14391(.A1(new_n15406_), .A2(new_n15371_), .ZN(new_n15412_));
  NAND3_X1   g14392(.A1(new_n15412_), .A2(new_n15411_), .A3(new_n15366_), .ZN(new_n15413_));
  NAND3_X1   g14393(.A1(new_n15410_), .A2(new_n15413_), .A3(new_n15405_), .ZN(new_n15414_));
  NOR2_X1    g14394(.A1(new_n15408_), .A2(new_n15373_), .ZN(new_n15415_));
  NOR2_X1    g14395(.A1(new_n15381_), .A2(new_n15402_), .ZN(new_n15416_));
  NOR2_X1    g14396(.A1(new_n15416_), .A2(new_n15406_), .ZN(new_n15417_));
  NOR2_X1    g14397(.A1(new_n15346_), .A2(new_n15344_), .ZN(new_n15418_));
  NOR2_X1    g14398(.A1(new_n15353_), .A2(new_n15351_), .ZN(new_n15419_));
  NOR2_X1    g14399(.A1(new_n15418_), .A2(new_n15419_), .ZN(new_n15420_));
  NOR2_X1    g14400(.A1(new_n15420_), .A2(new_n15354_), .ZN(new_n15421_));
  NAND2_X1   g14401(.A1(new_n15418_), .A2(new_n15419_), .ZN(new_n15422_));
  NAND2_X1   g14402(.A1(new_n15333_), .A2(new_n15338_), .ZN(new_n15423_));
  NOR2_X1    g14403(.A1(new_n15422_), .A2(new_n15423_), .ZN(new_n15424_));
  NAND4_X1   g14404(.A1(new_n15415_), .A2(new_n15417_), .A3(new_n15421_), .A4(new_n15424_), .ZN(new_n15425_));
  NOR2_X1    g14405(.A1(new_n15414_), .A2(new_n15425_), .ZN(new_n15426_));
  AOI21_X1   g14406(.A1(new_n15412_), .A2(new_n15411_), .B(new_n15366_), .ZN(new_n15427_));
  NOR3_X1    g14407(.A1(new_n15407_), .A2(new_n15409_), .A3(new_n15365_), .ZN(new_n15428_));
  NOR3_X1    g14408(.A1(new_n15427_), .A2(new_n15428_), .A3(new_n15404_), .ZN(new_n15429_));
  NAND2_X1   g14409(.A1(new_n15417_), .A2(new_n15415_), .ZN(new_n15430_));
  NAND2_X1   g14410(.A1(new_n15421_), .A2(new_n15424_), .ZN(new_n15431_));
  NOR2_X1    g14411(.A1(new_n15430_), .A2(new_n15431_), .ZN(new_n15432_));
  NOR2_X1    g14412(.A1(new_n15429_), .A2(new_n15432_), .ZN(new_n15433_));
  OAI21_X1   g14413(.A1(new_n15433_), .A2(new_n15426_), .B(new_n15361_), .ZN(new_n15434_));
  NAND2_X1   g14414(.A1(new_n15414_), .A2(new_n15432_), .ZN(new_n15435_));
  NAND2_X1   g14415(.A1(new_n15410_), .A2(new_n15413_), .ZN(new_n15436_));
  NAND3_X1   g14416(.A1(new_n15417_), .A2(new_n15415_), .A3(new_n15421_), .ZN(new_n15437_));
  NOR3_X1    g14417(.A1(new_n15404_), .A2(new_n15422_), .A3(new_n15423_), .ZN(new_n15438_));
  OAI21_X1   g14418(.A1(new_n15436_), .A2(new_n15437_), .B(new_n15438_), .ZN(new_n15439_));
  NAND3_X1   g14419(.A1(new_n15435_), .A2(new_n15439_), .A3(new_n15361_), .ZN(new_n15440_));
  NAND2_X1   g14420(.A1(new_n15434_), .A2(new_n15440_), .ZN(new_n15441_));
  INV_X1     g14421(.I(new_n15361_), .ZN(new_n15442_));
  NAND2_X1   g14422(.A1(new_n15429_), .A2(new_n15432_), .ZN(new_n15443_));
  NAND2_X1   g14423(.A1(new_n15414_), .A2(new_n15425_), .ZN(new_n15444_));
  AOI21_X1   g14424(.A1(new_n15443_), .A2(new_n15444_), .B(new_n15442_), .ZN(new_n15445_));
  INV_X1     g14425(.I(new_n15440_), .ZN(new_n15446_));
  XNOR2_X1   g14426(.A1(new_n15430_), .A2(new_n15431_), .ZN(new_n15447_));
  INV_X1     g14427(.I(\A[591] ), .ZN(new_n15448_));
  NOR2_X1    g14428(.A1(new_n15448_), .A2(\A[590] ), .ZN(new_n15449_));
  INV_X1     g14429(.I(\A[590] ), .ZN(new_n15450_));
  NOR2_X1    g14430(.A1(new_n15450_), .A2(\A[591] ), .ZN(new_n15451_));
  OAI21_X1   g14431(.A1(new_n15449_), .A2(new_n15451_), .B(\A[589] ), .ZN(new_n15452_));
  INV_X1     g14432(.I(\A[589] ), .ZN(new_n15453_));
  NOR2_X1    g14433(.A1(\A[590] ), .A2(\A[591] ), .ZN(new_n15454_));
  NOR2_X1    g14434(.A1(new_n15450_), .A2(new_n15448_), .ZN(new_n15455_));
  OAI21_X1   g14435(.A1(new_n15455_), .A2(new_n15454_), .B(new_n15453_), .ZN(new_n15456_));
  INV_X1     g14436(.I(\A[594] ), .ZN(new_n15457_));
  NOR2_X1    g14437(.A1(new_n15457_), .A2(\A[593] ), .ZN(new_n15458_));
  INV_X1     g14438(.I(\A[593] ), .ZN(new_n15459_));
  NOR2_X1    g14439(.A1(new_n15459_), .A2(\A[594] ), .ZN(new_n15460_));
  OAI21_X1   g14440(.A1(new_n15458_), .A2(new_n15460_), .B(\A[592] ), .ZN(new_n15461_));
  INV_X1     g14441(.I(\A[592] ), .ZN(new_n15462_));
  NOR2_X1    g14442(.A1(\A[593] ), .A2(\A[594] ), .ZN(new_n15463_));
  NOR2_X1    g14443(.A1(new_n15459_), .A2(new_n15457_), .ZN(new_n15464_));
  OAI21_X1   g14444(.A1(new_n15464_), .A2(new_n15463_), .B(new_n15462_), .ZN(new_n15465_));
  NAND4_X1   g14445(.A1(new_n15452_), .A2(new_n15456_), .A3(new_n15465_), .A4(new_n15461_), .ZN(new_n15466_));
  NOR2_X1    g14446(.A1(new_n15464_), .A2(\A[592] ), .ZN(new_n15467_));
  NOR2_X1    g14447(.A1(new_n15467_), .A2(new_n15463_), .ZN(new_n15468_));
  NOR2_X1    g14448(.A1(new_n15455_), .A2(\A[589] ), .ZN(new_n15469_));
  NOR2_X1    g14449(.A1(new_n15469_), .A2(new_n15454_), .ZN(new_n15470_));
  NAND2_X1   g14450(.A1(new_n15468_), .A2(new_n15470_), .ZN(new_n15471_));
  NOR2_X1    g14451(.A1(new_n15471_), .A2(new_n15466_), .ZN(new_n15472_));
  NAND2_X1   g14452(.A1(new_n15456_), .A2(new_n15452_), .ZN(new_n15473_));
  NAND2_X1   g14453(.A1(new_n15465_), .A2(new_n15461_), .ZN(new_n15474_));
  NAND2_X1   g14454(.A1(new_n15473_), .A2(new_n15474_), .ZN(new_n15475_));
  NAND3_X1   g14455(.A1(new_n15472_), .A2(new_n15466_), .A3(new_n15475_), .ZN(new_n15476_));
  INV_X1     g14456(.I(\A[583] ), .ZN(new_n15477_));
  INV_X1     g14457(.I(\A[584] ), .ZN(new_n15478_));
  NAND2_X1   g14458(.A1(new_n15478_), .A2(\A[585] ), .ZN(new_n15479_));
  INV_X1     g14459(.I(\A[585] ), .ZN(new_n15480_));
  NAND2_X1   g14460(.A1(new_n15480_), .A2(\A[584] ), .ZN(new_n15481_));
  AOI21_X1   g14461(.A1(new_n15479_), .A2(new_n15481_), .B(new_n15477_), .ZN(new_n15482_));
  NAND2_X1   g14462(.A1(new_n15478_), .A2(new_n15480_), .ZN(new_n15483_));
  NAND2_X1   g14463(.A1(\A[584] ), .A2(\A[585] ), .ZN(new_n15484_));
  AOI21_X1   g14464(.A1(new_n15483_), .A2(new_n15484_), .B(\A[583] ), .ZN(new_n15485_));
  INV_X1     g14465(.I(\A[586] ), .ZN(new_n15486_));
  INV_X1     g14466(.I(\A[587] ), .ZN(new_n15487_));
  NAND2_X1   g14467(.A1(new_n15487_), .A2(\A[588] ), .ZN(new_n15488_));
  INV_X1     g14468(.I(\A[588] ), .ZN(new_n15489_));
  NAND2_X1   g14469(.A1(new_n15489_), .A2(\A[587] ), .ZN(new_n15490_));
  AOI21_X1   g14470(.A1(new_n15488_), .A2(new_n15490_), .B(new_n15486_), .ZN(new_n15491_));
  NAND2_X1   g14471(.A1(new_n15487_), .A2(new_n15489_), .ZN(new_n15492_));
  NAND2_X1   g14472(.A1(\A[587] ), .A2(\A[588] ), .ZN(new_n15493_));
  AOI21_X1   g14473(.A1(new_n15492_), .A2(new_n15493_), .B(\A[586] ), .ZN(new_n15494_));
  NOR4_X1    g14474(.A1(new_n15482_), .A2(new_n15485_), .A3(new_n15494_), .A4(new_n15491_), .ZN(new_n15495_));
  NAND2_X1   g14475(.A1(new_n15493_), .A2(new_n15486_), .ZN(new_n15496_));
  NAND2_X1   g14476(.A1(new_n15496_), .A2(new_n15492_), .ZN(new_n15497_));
  NAND2_X1   g14477(.A1(new_n15484_), .A2(new_n15477_), .ZN(new_n15498_));
  NAND2_X1   g14478(.A1(new_n15498_), .A2(new_n15483_), .ZN(new_n15499_));
  NOR2_X1    g14479(.A1(new_n15497_), .A2(new_n15499_), .ZN(new_n15500_));
  NOR2_X1    g14480(.A1(new_n15485_), .A2(new_n15482_), .ZN(new_n15501_));
  NOR2_X1    g14481(.A1(new_n15494_), .A2(new_n15491_), .ZN(new_n15502_));
  NOR2_X1    g14482(.A1(new_n15501_), .A2(new_n15502_), .ZN(new_n15503_));
  NAND2_X1   g14483(.A1(new_n15447_), .A2(new_n15476_), .ZN(new_n15504_));
  OAI21_X1   g14484(.A1(new_n15446_), .A2(new_n15445_), .B(new_n15504_), .ZN(new_n15505_));
  XOR2_X1    g14485(.A1(new_n15430_), .A2(new_n15431_), .Z(new_n15506_));
  INV_X1     g14486(.I(new_n15476_), .ZN(new_n15507_));
  NOR2_X1    g14487(.A1(new_n15506_), .A2(new_n15507_), .ZN(new_n15508_));
  NAND3_X1   g14488(.A1(new_n15434_), .A2(new_n15440_), .A3(new_n15508_), .ZN(new_n15509_));
  NAND2_X1   g14489(.A1(new_n15466_), .A2(new_n15470_), .ZN(new_n15510_));
  INV_X1     g14490(.I(new_n15510_), .ZN(new_n15511_));
  NOR2_X1    g14491(.A1(new_n15466_), .A2(new_n15470_), .ZN(new_n15512_));
  OAI21_X1   g14492(.A1(new_n15511_), .A2(new_n15512_), .B(new_n15468_), .ZN(new_n15513_));
  INV_X1     g14493(.I(new_n15468_), .ZN(new_n15514_));
  OR3_X2     g14494(.A1(new_n15473_), .A2(new_n15474_), .A3(new_n15470_), .Z(new_n15515_));
  NAND3_X1   g14495(.A1(new_n15515_), .A2(new_n15510_), .A3(new_n15514_), .ZN(new_n15516_));
  AND2_X2    g14496(.A1(new_n15513_), .A2(new_n15516_), .Z(new_n15517_));
  NOR3_X1    g14497(.A1(new_n15476_), .A2(new_n15495_), .A3(new_n15503_), .ZN(new_n15518_));
  NAND2_X1   g14498(.A1(new_n15501_), .A2(new_n15502_), .ZN(new_n15519_));
  INV_X1     g14499(.I(new_n15500_), .ZN(new_n15520_));
  NOR2_X1    g14500(.A1(new_n15519_), .A2(new_n15520_), .ZN(new_n15521_));
  INV_X1     g14501(.I(new_n15471_), .ZN(new_n15522_));
  XOR2_X1    g14502(.A1(new_n15473_), .A2(new_n15474_), .Z(new_n15523_));
  NAND2_X1   g14503(.A1(new_n15523_), .A2(new_n15522_), .ZN(new_n15524_));
  NAND2_X1   g14504(.A1(new_n15524_), .A2(new_n15521_), .ZN(new_n15525_));
  AOI21_X1   g14505(.A1(new_n15517_), .A2(new_n15518_), .B(new_n15525_), .ZN(new_n15526_));
  INV_X1     g14506(.I(new_n15497_), .ZN(new_n15527_));
  NOR2_X1    g14507(.A1(new_n15495_), .A2(new_n15499_), .ZN(new_n15528_));
  INV_X1     g14508(.I(new_n15499_), .ZN(new_n15529_));
  NOR2_X1    g14509(.A1(new_n15519_), .A2(new_n15529_), .ZN(new_n15530_));
  OAI21_X1   g14510(.A1(new_n15530_), .A2(new_n15528_), .B(new_n15527_), .ZN(new_n15531_));
  INV_X1     g14511(.I(new_n15528_), .ZN(new_n15532_));
  NAND2_X1   g14512(.A1(new_n15495_), .A2(new_n15499_), .ZN(new_n15533_));
  NAND3_X1   g14513(.A1(new_n15532_), .A2(new_n15497_), .A3(new_n15533_), .ZN(new_n15534_));
  NAND2_X1   g14514(.A1(new_n15534_), .A2(new_n15531_), .ZN(new_n15535_));
  NAND2_X1   g14515(.A1(new_n15526_), .A2(new_n15535_), .ZN(new_n15536_));
  NOR2_X1    g14516(.A1(new_n15503_), .A2(new_n15495_), .ZN(new_n15537_));
  NAND2_X1   g14517(.A1(new_n15537_), .A2(new_n15521_), .ZN(new_n15538_));
  NOR2_X1    g14518(.A1(new_n15538_), .A2(new_n15476_), .ZN(new_n15539_));
  INV_X1     g14519(.I(new_n15539_), .ZN(new_n15540_));
  NAND2_X1   g14520(.A1(new_n15540_), .A2(new_n15535_), .ZN(new_n15541_));
  AOI21_X1   g14521(.A1(new_n15532_), .A2(new_n15533_), .B(new_n15497_), .ZN(new_n15542_));
  NOR3_X1    g14522(.A1(new_n15530_), .A2(new_n15527_), .A3(new_n15528_), .ZN(new_n15543_));
  NOR4_X1    g14523(.A1(new_n15542_), .A2(new_n15543_), .A3(new_n15538_), .A4(new_n15476_), .ZN(new_n15544_));
  AOI21_X1   g14524(.A1(new_n15517_), .A2(new_n15524_), .B(new_n15544_), .ZN(new_n15545_));
  NAND3_X1   g14525(.A1(new_n15524_), .A2(new_n15513_), .A3(new_n15516_), .ZN(new_n15546_));
  NOR3_X1    g14526(.A1(new_n15540_), .A2(new_n15535_), .A3(new_n15546_), .ZN(new_n15547_));
  OAI21_X1   g14527(.A1(new_n15545_), .A2(new_n15547_), .B(new_n15541_), .ZN(new_n15548_));
  NAND2_X1   g14528(.A1(new_n15548_), .A2(new_n15536_), .ZN(new_n15549_));
  AOI22_X1   g14529(.A1(new_n15505_), .A2(new_n15509_), .B1(new_n15549_), .B2(new_n15441_), .ZN(new_n15550_));
  INV_X1     g14530(.I(new_n15439_), .ZN(new_n15551_));
  AOI21_X1   g14531(.A1(new_n15414_), .A2(new_n15432_), .B(new_n15361_), .ZN(new_n15552_));
  NOR2_X1    g14532(.A1(new_n15365_), .A2(new_n15370_), .ZN(new_n15553_));
  OAI21_X1   g14533(.A1(new_n15408_), .A2(new_n15553_), .B(new_n15373_), .ZN(new_n15554_));
  NOR2_X1    g14534(.A1(new_n15333_), .A2(new_n15338_), .ZN(new_n15555_));
  OAI21_X1   g14535(.A1(new_n15422_), .A2(new_n15555_), .B(new_n15423_), .ZN(new_n15556_));
  XNOR2_X1   g14536(.A1(new_n15554_), .A2(new_n15556_), .ZN(new_n15557_));
  INV_X1     g14537(.I(new_n15557_), .ZN(new_n15558_));
  NOR3_X1    g14538(.A1(new_n15551_), .A2(new_n15552_), .A3(new_n15558_), .ZN(new_n15559_));
  AOI22_X1   g14539(.A1(new_n15546_), .A2(new_n15539_), .B1(new_n15531_), .B2(new_n15534_), .ZN(new_n15560_));
  NOR2_X1    g14540(.A1(new_n15468_), .A2(new_n15470_), .ZN(new_n15561_));
  OAI21_X1   g14541(.A1(new_n15466_), .A2(new_n15561_), .B(new_n15471_), .ZN(new_n15562_));
  NOR2_X1    g14542(.A1(new_n15527_), .A2(new_n15529_), .ZN(new_n15563_));
  OAI21_X1   g14543(.A1(new_n15519_), .A2(new_n15563_), .B(new_n15520_), .ZN(new_n15564_));
  XOR2_X1    g14544(.A1(new_n15564_), .A2(new_n15562_), .Z(new_n15565_));
  NOR3_X1    g14545(.A1(new_n15526_), .A2(new_n15560_), .A3(new_n15565_), .ZN(new_n15566_));
  NAND3_X1   g14546(.A1(new_n15550_), .A2(new_n15559_), .A3(new_n15566_), .ZN(new_n15567_));
  NAND2_X1   g14547(.A1(new_n15564_), .A2(new_n15562_), .ZN(new_n15568_));
  NOR2_X1    g14548(.A1(new_n15526_), .A2(new_n15560_), .ZN(new_n15569_));
  OAI21_X1   g14549(.A1(new_n15562_), .A2(new_n15564_), .B(new_n15569_), .ZN(new_n15570_));
  NAND2_X1   g14550(.A1(new_n15570_), .A2(new_n15568_), .ZN(new_n15571_));
  NAND2_X1   g14551(.A1(new_n15554_), .A2(new_n15556_), .ZN(new_n15572_));
  NOR2_X1    g14552(.A1(new_n15551_), .A2(new_n15552_), .ZN(new_n15573_));
  OAI21_X1   g14553(.A1(new_n15554_), .A2(new_n15556_), .B(new_n15573_), .ZN(new_n15574_));
  NAND2_X1   g14554(.A1(new_n15574_), .A2(new_n15572_), .ZN(new_n15575_));
  OAI21_X1   g14555(.A1(new_n15571_), .A2(new_n15575_), .B(new_n15567_), .ZN(new_n15576_));
  NAND2_X1   g14556(.A1(new_n15575_), .A2(new_n15571_), .ZN(new_n15577_));
  NAND2_X1   g14557(.A1(new_n15576_), .A2(new_n15577_), .ZN(new_n15578_));
  INV_X1     g14558(.I(\A[574] ), .ZN(new_n15579_));
  NOR2_X1    g14559(.A1(\A[575] ), .A2(\A[576] ), .ZN(new_n15580_));
  NAND2_X1   g14560(.A1(\A[575] ), .A2(\A[576] ), .ZN(new_n15581_));
  AOI21_X1   g14561(.A1(new_n15579_), .A2(new_n15581_), .B(new_n15580_), .ZN(new_n15582_));
  INV_X1     g14562(.I(new_n15582_), .ZN(new_n15583_));
  INV_X1     g14563(.I(\A[571] ), .ZN(new_n15584_));
  NOR2_X1    g14564(.A1(\A[572] ), .A2(\A[573] ), .ZN(new_n15585_));
  NAND2_X1   g14565(.A1(\A[572] ), .A2(\A[573] ), .ZN(new_n15586_));
  AOI21_X1   g14566(.A1(new_n15584_), .A2(new_n15586_), .B(new_n15585_), .ZN(new_n15587_));
  INV_X1     g14567(.I(\A[572] ), .ZN(new_n15588_));
  NAND2_X1   g14568(.A1(new_n15588_), .A2(\A[573] ), .ZN(new_n15589_));
  INV_X1     g14569(.I(\A[573] ), .ZN(new_n15590_));
  NAND2_X1   g14570(.A1(new_n15590_), .A2(\A[572] ), .ZN(new_n15591_));
  AOI21_X1   g14571(.A1(new_n15589_), .A2(new_n15591_), .B(new_n15584_), .ZN(new_n15592_));
  INV_X1     g14572(.I(new_n15585_), .ZN(new_n15593_));
  AOI21_X1   g14573(.A1(new_n15593_), .A2(new_n15586_), .B(\A[571] ), .ZN(new_n15594_));
  NOR2_X1    g14574(.A1(new_n15594_), .A2(new_n15592_), .ZN(new_n15595_));
  INV_X1     g14575(.I(\A[575] ), .ZN(new_n15596_));
  NAND2_X1   g14576(.A1(new_n15596_), .A2(\A[576] ), .ZN(new_n15597_));
  INV_X1     g14577(.I(\A[576] ), .ZN(new_n15598_));
  NAND2_X1   g14578(.A1(new_n15598_), .A2(\A[575] ), .ZN(new_n15599_));
  AOI21_X1   g14579(.A1(new_n15597_), .A2(new_n15599_), .B(new_n15579_), .ZN(new_n15600_));
  INV_X1     g14580(.I(new_n15580_), .ZN(new_n15601_));
  AOI21_X1   g14581(.A1(new_n15601_), .A2(new_n15581_), .B(\A[574] ), .ZN(new_n15602_));
  NOR2_X1    g14582(.A1(new_n15602_), .A2(new_n15600_), .ZN(new_n15603_));
  NAND2_X1   g14583(.A1(new_n15595_), .A2(new_n15603_), .ZN(new_n15604_));
  NAND2_X1   g14584(.A1(new_n15604_), .A2(new_n15587_), .ZN(new_n15605_));
  INV_X1     g14585(.I(new_n15587_), .ZN(new_n15606_));
  NOR4_X1    g14586(.A1(new_n15592_), .A2(new_n15594_), .A3(new_n15602_), .A4(new_n15600_), .ZN(new_n15607_));
  NAND2_X1   g14587(.A1(new_n15607_), .A2(new_n15606_), .ZN(new_n15608_));
  AOI21_X1   g14588(.A1(new_n15605_), .A2(new_n15608_), .B(new_n15583_), .ZN(new_n15609_));
  AND3_X2    g14589(.A1(new_n15605_), .A2(new_n15583_), .A3(new_n15608_), .Z(new_n15610_));
  NOR2_X1    g14590(.A1(new_n15610_), .A2(new_n15609_), .ZN(new_n15611_));
  INV_X1     g14591(.I(\A[580] ), .ZN(new_n15612_));
  NOR2_X1    g14592(.A1(\A[581] ), .A2(\A[582] ), .ZN(new_n15613_));
  NAND2_X1   g14593(.A1(\A[581] ), .A2(\A[582] ), .ZN(new_n15614_));
  AOI21_X1   g14594(.A1(new_n15612_), .A2(new_n15614_), .B(new_n15613_), .ZN(new_n15615_));
  INV_X1     g14595(.I(new_n15615_), .ZN(new_n15616_));
  INV_X1     g14596(.I(\A[577] ), .ZN(new_n15617_));
  NOR2_X1    g14597(.A1(\A[578] ), .A2(\A[579] ), .ZN(new_n15618_));
  NAND2_X1   g14598(.A1(\A[578] ), .A2(\A[579] ), .ZN(new_n15619_));
  AOI21_X1   g14599(.A1(new_n15617_), .A2(new_n15619_), .B(new_n15618_), .ZN(new_n15620_));
  INV_X1     g14600(.I(new_n15620_), .ZN(new_n15621_));
  NOR2_X1    g14601(.A1(new_n15616_), .A2(new_n15621_), .ZN(new_n15622_));
  INV_X1     g14602(.I(new_n15622_), .ZN(new_n15623_));
  INV_X1     g14603(.I(\A[578] ), .ZN(new_n15624_));
  NAND2_X1   g14604(.A1(new_n15624_), .A2(\A[579] ), .ZN(new_n15625_));
  INV_X1     g14605(.I(\A[579] ), .ZN(new_n15626_));
  NAND2_X1   g14606(.A1(new_n15626_), .A2(\A[578] ), .ZN(new_n15627_));
  AOI21_X1   g14607(.A1(new_n15625_), .A2(new_n15627_), .B(new_n15617_), .ZN(new_n15628_));
  INV_X1     g14608(.I(new_n15618_), .ZN(new_n15629_));
  AOI21_X1   g14609(.A1(new_n15629_), .A2(new_n15619_), .B(\A[577] ), .ZN(new_n15630_));
  NOR2_X1    g14610(.A1(new_n15630_), .A2(new_n15628_), .ZN(new_n15631_));
  INV_X1     g14611(.I(\A[582] ), .ZN(new_n15632_));
  NOR2_X1    g14612(.A1(new_n15632_), .A2(\A[581] ), .ZN(new_n15633_));
  INV_X1     g14613(.I(\A[581] ), .ZN(new_n15634_));
  NOR2_X1    g14614(.A1(new_n15634_), .A2(\A[582] ), .ZN(new_n15635_));
  OAI21_X1   g14615(.A1(new_n15633_), .A2(new_n15635_), .B(\A[580] ), .ZN(new_n15636_));
  INV_X1     g14616(.I(new_n15614_), .ZN(new_n15637_));
  OAI21_X1   g14617(.A1(new_n15637_), .A2(new_n15613_), .B(new_n15612_), .ZN(new_n15638_));
  NAND2_X1   g14618(.A1(new_n15636_), .A2(new_n15638_), .ZN(new_n15639_));
  NAND2_X1   g14619(.A1(new_n15631_), .A2(new_n15639_), .ZN(new_n15640_));
  NOR2_X1    g14620(.A1(new_n15626_), .A2(\A[578] ), .ZN(new_n15641_));
  NOR2_X1    g14621(.A1(new_n15624_), .A2(\A[579] ), .ZN(new_n15642_));
  OAI21_X1   g14622(.A1(new_n15641_), .A2(new_n15642_), .B(\A[577] ), .ZN(new_n15643_));
  INV_X1     g14623(.I(new_n15619_), .ZN(new_n15644_));
  OAI21_X1   g14624(.A1(new_n15644_), .A2(new_n15618_), .B(new_n15617_), .ZN(new_n15645_));
  NAND2_X1   g14625(.A1(new_n15643_), .A2(new_n15645_), .ZN(new_n15646_));
  NAND2_X1   g14626(.A1(new_n15634_), .A2(\A[582] ), .ZN(new_n15647_));
  NAND2_X1   g14627(.A1(new_n15632_), .A2(\A[581] ), .ZN(new_n15648_));
  AOI21_X1   g14628(.A1(new_n15647_), .A2(new_n15648_), .B(new_n15612_), .ZN(new_n15649_));
  INV_X1     g14629(.I(new_n15613_), .ZN(new_n15650_));
  AOI21_X1   g14630(.A1(new_n15650_), .A2(new_n15614_), .B(\A[580] ), .ZN(new_n15651_));
  NOR2_X1    g14631(.A1(new_n15651_), .A2(new_n15649_), .ZN(new_n15652_));
  NAND2_X1   g14632(.A1(new_n15652_), .A2(new_n15646_), .ZN(new_n15653_));
  AOI21_X1   g14633(.A1(new_n15640_), .A2(new_n15653_), .B(new_n15623_), .ZN(new_n15654_));
  INV_X1     g14634(.I(new_n15654_), .ZN(new_n15655_));
  NOR2_X1    g14635(.A1(new_n15646_), .A2(new_n15639_), .ZN(new_n15656_));
  NOR2_X1    g14636(.A1(new_n15656_), .A2(new_n15621_), .ZN(new_n15657_));
  NAND2_X1   g14637(.A1(new_n15631_), .A2(new_n15652_), .ZN(new_n15658_));
  NOR2_X1    g14638(.A1(new_n15658_), .A2(new_n15620_), .ZN(new_n15659_));
  OAI21_X1   g14639(.A1(new_n15657_), .A2(new_n15659_), .B(new_n15615_), .ZN(new_n15660_));
  NAND2_X1   g14640(.A1(new_n15658_), .A2(new_n15620_), .ZN(new_n15661_));
  NAND2_X1   g14641(.A1(new_n15656_), .A2(new_n15621_), .ZN(new_n15662_));
  NAND3_X1   g14642(.A1(new_n15662_), .A2(new_n15661_), .A3(new_n15616_), .ZN(new_n15663_));
  NAND3_X1   g14643(.A1(new_n15660_), .A2(new_n15663_), .A3(new_n15655_), .ZN(new_n15664_));
  NOR2_X1    g14644(.A1(new_n15658_), .A2(new_n15623_), .ZN(new_n15665_));
  NOR2_X1    g14645(.A1(new_n15631_), .A2(new_n15652_), .ZN(new_n15666_));
  NOR2_X1    g14646(.A1(new_n15666_), .A2(new_n15656_), .ZN(new_n15667_));
  NOR2_X1    g14647(.A1(new_n15595_), .A2(new_n15603_), .ZN(new_n15668_));
  NOR2_X1    g14648(.A1(new_n15668_), .A2(new_n15607_), .ZN(new_n15669_));
  NAND2_X1   g14649(.A1(new_n15582_), .A2(new_n15587_), .ZN(new_n15670_));
  NOR2_X1    g14650(.A1(new_n15604_), .A2(new_n15670_), .ZN(new_n15671_));
  NAND4_X1   g14651(.A1(new_n15665_), .A2(new_n15667_), .A3(new_n15669_), .A4(new_n15671_), .ZN(new_n15672_));
  NOR2_X1    g14652(.A1(new_n15664_), .A2(new_n15672_), .ZN(new_n15673_));
  AOI21_X1   g14653(.A1(new_n15662_), .A2(new_n15661_), .B(new_n15616_), .ZN(new_n15674_));
  NOR3_X1    g14654(.A1(new_n15657_), .A2(new_n15659_), .A3(new_n15615_), .ZN(new_n15675_));
  NOR3_X1    g14655(.A1(new_n15674_), .A2(new_n15675_), .A3(new_n15654_), .ZN(new_n15676_));
  NAND2_X1   g14656(.A1(new_n15667_), .A2(new_n15665_), .ZN(new_n15677_));
  NAND2_X1   g14657(.A1(new_n15669_), .A2(new_n15671_), .ZN(new_n15678_));
  NOR2_X1    g14658(.A1(new_n15677_), .A2(new_n15678_), .ZN(new_n15679_));
  NOR2_X1    g14659(.A1(new_n15676_), .A2(new_n15679_), .ZN(new_n15680_));
  OAI21_X1   g14660(.A1(new_n15680_), .A2(new_n15673_), .B(new_n15611_), .ZN(new_n15681_));
  NAND2_X1   g14661(.A1(new_n15664_), .A2(new_n15679_), .ZN(new_n15682_));
  NAND2_X1   g14662(.A1(new_n15660_), .A2(new_n15663_), .ZN(new_n15683_));
  NAND3_X1   g14663(.A1(new_n15667_), .A2(new_n15665_), .A3(new_n15669_), .ZN(new_n15684_));
  NOR3_X1    g14664(.A1(new_n15654_), .A2(new_n15604_), .A3(new_n15670_), .ZN(new_n15685_));
  OAI21_X1   g14665(.A1(new_n15683_), .A2(new_n15684_), .B(new_n15685_), .ZN(new_n15686_));
  NAND3_X1   g14666(.A1(new_n15682_), .A2(new_n15686_), .A3(new_n15611_), .ZN(new_n15687_));
  NAND2_X1   g14667(.A1(new_n15681_), .A2(new_n15687_), .ZN(new_n15688_));
  XOR2_X1    g14668(.A1(new_n15677_), .A2(new_n15678_), .Z(new_n15689_));
  INV_X1     g14669(.I(\A[567] ), .ZN(new_n15690_));
  NOR2_X1    g14670(.A1(new_n15690_), .A2(\A[566] ), .ZN(new_n15691_));
  INV_X1     g14671(.I(\A[566] ), .ZN(new_n15692_));
  NOR2_X1    g14672(.A1(new_n15692_), .A2(\A[567] ), .ZN(new_n15693_));
  OAI21_X1   g14673(.A1(new_n15691_), .A2(new_n15693_), .B(\A[565] ), .ZN(new_n15694_));
  INV_X1     g14674(.I(\A[565] ), .ZN(new_n15695_));
  NOR2_X1    g14675(.A1(\A[566] ), .A2(\A[567] ), .ZN(new_n15696_));
  NAND2_X1   g14676(.A1(\A[566] ), .A2(\A[567] ), .ZN(new_n15697_));
  INV_X1     g14677(.I(new_n15697_), .ZN(new_n15698_));
  OAI21_X1   g14678(.A1(new_n15698_), .A2(new_n15696_), .B(new_n15695_), .ZN(new_n15699_));
  NAND2_X1   g14679(.A1(new_n15694_), .A2(new_n15699_), .ZN(new_n15700_));
  INV_X1     g14680(.I(\A[570] ), .ZN(new_n15701_));
  NOR2_X1    g14681(.A1(new_n15701_), .A2(\A[569] ), .ZN(new_n15702_));
  INV_X1     g14682(.I(\A[569] ), .ZN(new_n15703_));
  NOR2_X1    g14683(.A1(new_n15703_), .A2(\A[570] ), .ZN(new_n15704_));
  OAI21_X1   g14684(.A1(new_n15702_), .A2(new_n15704_), .B(\A[568] ), .ZN(new_n15705_));
  INV_X1     g14685(.I(\A[568] ), .ZN(new_n15706_));
  NOR2_X1    g14686(.A1(\A[569] ), .A2(\A[570] ), .ZN(new_n15707_));
  NAND2_X1   g14687(.A1(\A[569] ), .A2(\A[570] ), .ZN(new_n15708_));
  INV_X1     g14688(.I(new_n15708_), .ZN(new_n15709_));
  OAI21_X1   g14689(.A1(new_n15709_), .A2(new_n15707_), .B(new_n15706_), .ZN(new_n15710_));
  NAND2_X1   g14690(.A1(new_n15705_), .A2(new_n15710_), .ZN(new_n15711_));
  NOR2_X1    g14691(.A1(new_n15700_), .A2(new_n15711_), .ZN(new_n15712_));
  AOI21_X1   g14692(.A1(new_n15706_), .A2(new_n15708_), .B(new_n15707_), .ZN(new_n15713_));
  INV_X1     g14693(.I(new_n15713_), .ZN(new_n15714_));
  AOI21_X1   g14694(.A1(new_n15695_), .A2(new_n15697_), .B(new_n15696_), .ZN(new_n15715_));
  INV_X1     g14695(.I(new_n15715_), .ZN(new_n15716_));
  NOR2_X1    g14696(.A1(new_n15714_), .A2(new_n15716_), .ZN(new_n15717_));
  NAND2_X1   g14697(.A1(new_n15712_), .A2(new_n15717_), .ZN(new_n15718_));
  NAND2_X1   g14698(.A1(new_n15692_), .A2(\A[567] ), .ZN(new_n15719_));
  NAND2_X1   g14699(.A1(new_n15690_), .A2(\A[566] ), .ZN(new_n15720_));
  AOI21_X1   g14700(.A1(new_n15719_), .A2(new_n15720_), .B(new_n15695_), .ZN(new_n15721_));
  INV_X1     g14701(.I(new_n15696_), .ZN(new_n15722_));
  AOI21_X1   g14702(.A1(new_n15722_), .A2(new_n15697_), .B(\A[565] ), .ZN(new_n15723_));
  NOR2_X1    g14703(.A1(new_n15723_), .A2(new_n15721_), .ZN(new_n15724_));
  NAND2_X1   g14704(.A1(new_n15703_), .A2(\A[570] ), .ZN(new_n15725_));
  NAND2_X1   g14705(.A1(new_n15701_), .A2(\A[569] ), .ZN(new_n15726_));
  AOI21_X1   g14706(.A1(new_n15725_), .A2(new_n15726_), .B(new_n15706_), .ZN(new_n15727_));
  INV_X1     g14707(.I(new_n15707_), .ZN(new_n15728_));
  AOI21_X1   g14708(.A1(new_n15728_), .A2(new_n15708_), .B(\A[568] ), .ZN(new_n15729_));
  NOR2_X1    g14709(.A1(new_n15729_), .A2(new_n15727_), .ZN(new_n15730_));
  NAND2_X1   g14710(.A1(new_n15724_), .A2(new_n15730_), .ZN(new_n15731_));
  NAND2_X1   g14711(.A1(new_n15700_), .A2(new_n15711_), .ZN(new_n15732_));
  NAND2_X1   g14712(.A1(new_n15731_), .A2(new_n15732_), .ZN(new_n15733_));
  INV_X1     g14713(.I(\A[559] ), .ZN(new_n15734_));
  INV_X1     g14714(.I(\A[560] ), .ZN(new_n15735_));
  NAND2_X1   g14715(.A1(new_n15735_), .A2(\A[561] ), .ZN(new_n15736_));
  INV_X1     g14716(.I(\A[561] ), .ZN(new_n15737_));
  NAND2_X1   g14717(.A1(new_n15737_), .A2(\A[560] ), .ZN(new_n15738_));
  AOI21_X1   g14718(.A1(new_n15736_), .A2(new_n15738_), .B(new_n15734_), .ZN(new_n15739_));
  NAND2_X1   g14719(.A1(new_n15735_), .A2(new_n15737_), .ZN(new_n15740_));
  NAND2_X1   g14720(.A1(\A[560] ), .A2(\A[561] ), .ZN(new_n15741_));
  AOI21_X1   g14721(.A1(new_n15740_), .A2(new_n15741_), .B(\A[559] ), .ZN(new_n15742_));
  NOR2_X1    g14722(.A1(new_n15742_), .A2(new_n15739_), .ZN(new_n15743_));
  INV_X1     g14723(.I(\A[562] ), .ZN(new_n15744_));
  INV_X1     g14724(.I(\A[563] ), .ZN(new_n15745_));
  NAND2_X1   g14725(.A1(new_n15745_), .A2(\A[564] ), .ZN(new_n15746_));
  INV_X1     g14726(.I(\A[564] ), .ZN(new_n15747_));
  NAND2_X1   g14727(.A1(new_n15747_), .A2(\A[563] ), .ZN(new_n15748_));
  AOI21_X1   g14728(.A1(new_n15746_), .A2(new_n15748_), .B(new_n15744_), .ZN(new_n15749_));
  NAND2_X1   g14729(.A1(new_n15745_), .A2(new_n15747_), .ZN(new_n15750_));
  NAND2_X1   g14730(.A1(\A[563] ), .A2(\A[564] ), .ZN(new_n15751_));
  AOI21_X1   g14731(.A1(new_n15750_), .A2(new_n15751_), .B(\A[562] ), .ZN(new_n15752_));
  NOR2_X1    g14732(.A1(new_n15752_), .A2(new_n15749_), .ZN(new_n15753_));
  NAND2_X1   g14733(.A1(new_n15751_), .A2(new_n15744_), .ZN(new_n15754_));
  NAND2_X1   g14734(.A1(new_n15754_), .A2(new_n15750_), .ZN(new_n15755_));
  NAND2_X1   g14735(.A1(new_n15741_), .A2(new_n15734_), .ZN(new_n15756_));
  NAND2_X1   g14736(.A1(new_n15756_), .A2(new_n15740_), .ZN(new_n15757_));
  NOR2_X1    g14737(.A1(new_n15755_), .A2(new_n15757_), .ZN(new_n15758_));
  NOR2_X1    g14738(.A1(new_n15733_), .A2(new_n15718_), .ZN(new_n15759_));
  NOR2_X1    g14739(.A1(new_n15689_), .A2(new_n15759_), .ZN(new_n15760_));
  AOI21_X1   g14740(.A1(new_n15681_), .A2(new_n15687_), .B(new_n15760_), .ZN(new_n15761_));
  INV_X1     g14741(.I(new_n15761_), .ZN(new_n15762_));
  NAND3_X1   g14742(.A1(new_n15681_), .A2(new_n15687_), .A3(new_n15760_), .ZN(new_n15763_));
  NOR2_X1    g14743(.A1(new_n15712_), .A2(new_n15716_), .ZN(new_n15764_));
  NOR2_X1    g14744(.A1(new_n15731_), .A2(new_n15715_), .ZN(new_n15765_));
  OAI21_X1   g14745(.A1(new_n15764_), .A2(new_n15765_), .B(new_n15713_), .ZN(new_n15766_));
  NAND2_X1   g14746(.A1(new_n15731_), .A2(new_n15715_), .ZN(new_n15767_));
  NAND2_X1   g14747(.A1(new_n15712_), .A2(new_n15716_), .ZN(new_n15768_));
  NAND3_X1   g14748(.A1(new_n15768_), .A2(new_n15767_), .A3(new_n15714_), .ZN(new_n15769_));
  AND2_X2    g14749(.A1(new_n15766_), .A2(new_n15769_), .Z(new_n15770_));
  INV_X1     g14750(.I(new_n15717_), .ZN(new_n15771_));
  NOR2_X1    g14751(.A1(new_n15731_), .A2(new_n15771_), .ZN(new_n15772_));
  NAND3_X1   g14752(.A1(new_n15772_), .A2(new_n15731_), .A3(new_n15732_), .ZN(new_n15773_));
  XNOR2_X1   g14753(.A1(new_n15743_), .A2(new_n15753_), .ZN(new_n15774_));
  NOR2_X1    g14754(.A1(new_n15773_), .A2(new_n15774_), .ZN(new_n15775_));
  NOR4_X1    g14755(.A1(new_n15739_), .A2(new_n15742_), .A3(new_n15752_), .A4(new_n15749_), .ZN(new_n15776_));
  XOR2_X1    g14756(.A1(new_n15700_), .A2(new_n15711_), .Z(new_n15777_));
  NAND2_X1   g14757(.A1(new_n15777_), .A2(new_n15717_), .ZN(new_n15778_));
  NAND3_X1   g14758(.A1(new_n15778_), .A2(new_n15776_), .A3(new_n15758_), .ZN(new_n15779_));
  AOI21_X1   g14759(.A1(new_n15770_), .A2(new_n15775_), .B(new_n15779_), .ZN(new_n15780_));
  INV_X1     g14760(.I(new_n15755_), .ZN(new_n15781_));
  NOR2_X1    g14761(.A1(new_n15776_), .A2(new_n15757_), .ZN(new_n15782_));
  NAND2_X1   g14762(.A1(new_n15776_), .A2(new_n15757_), .ZN(new_n15783_));
  INV_X1     g14763(.I(new_n15783_), .ZN(new_n15784_));
  OAI21_X1   g14764(.A1(new_n15784_), .A2(new_n15782_), .B(new_n15781_), .ZN(new_n15785_));
  NAND2_X1   g14765(.A1(new_n15743_), .A2(new_n15753_), .ZN(new_n15786_));
  INV_X1     g14766(.I(new_n15757_), .ZN(new_n15787_));
  NAND2_X1   g14767(.A1(new_n15786_), .A2(new_n15787_), .ZN(new_n15788_));
  NAND3_X1   g14768(.A1(new_n15788_), .A2(new_n15755_), .A3(new_n15783_), .ZN(new_n15789_));
  NAND2_X1   g14769(.A1(new_n15785_), .A2(new_n15789_), .ZN(new_n15790_));
  NAND2_X1   g14770(.A1(new_n15780_), .A2(new_n15790_), .ZN(new_n15791_));
  NOR2_X1    g14771(.A1(new_n15733_), .A2(new_n15718_), .ZN(new_n15792_));
  NAND2_X1   g14772(.A1(new_n15776_), .A2(new_n15758_), .ZN(new_n15793_));
  NOR2_X1    g14773(.A1(new_n15774_), .A2(new_n15793_), .ZN(new_n15794_));
  NAND2_X1   g14774(.A1(new_n15794_), .A2(new_n15792_), .ZN(new_n15795_));
  NAND2_X1   g14775(.A1(new_n15795_), .A2(new_n15790_), .ZN(new_n15796_));
  AND3_X2    g14776(.A1(new_n15778_), .A2(new_n15766_), .A3(new_n15769_), .Z(new_n15797_));
  NOR2_X1    g14777(.A1(new_n15795_), .A2(new_n15790_), .ZN(new_n15798_));
  NOR2_X1    g14778(.A1(new_n15798_), .A2(new_n15797_), .ZN(new_n15799_));
  NAND3_X1   g14779(.A1(new_n15778_), .A2(new_n15766_), .A3(new_n15769_), .ZN(new_n15800_));
  NOR3_X1    g14780(.A1(new_n15800_), .A2(new_n15795_), .A3(new_n15790_), .ZN(new_n15801_));
  OAI21_X1   g14781(.A1(new_n15799_), .A2(new_n15801_), .B(new_n15796_), .ZN(new_n15802_));
  NAND2_X1   g14782(.A1(new_n15802_), .A2(new_n15791_), .ZN(new_n15803_));
  AOI22_X1   g14783(.A1(new_n15762_), .A2(new_n15763_), .B1(new_n15803_), .B2(new_n15688_), .ZN(new_n15804_));
  OAI22_X1   g14784(.A1(new_n15676_), .A2(new_n15672_), .B1(new_n15609_), .B2(new_n15610_), .ZN(new_n15805_));
  NOR2_X1    g14785(.A1(new_n15615_), .A2(new_n15620_), .ZN(new_n15806_));
  OAI21_X1   g14786(.A1(new_n15658_), .A2(new_n15806_), .B(new_n15623_), .ZN(new_n15807_));
  NOR2_X1    g14787(.A1(new_n15582_), .A2(new_n15587_), .ZN(new_n15808_));
  OAI21_X1   g14788(.A1(new_n15604_), .A2(new_n15808_), .B(new_n15670_), .ZN(new_n15809_));
  XNOR2_X1   g14789(.A1(new_n15807_), .A2(new_n15809_), .ZN(new_n15810_));
  NAND3_X1   g14790(.A1(new_n15805_), .A2(new_n15686_), .A3(new_n15810_), .ZN(new_n15811_));
  INV_X1     g14791(.I(new_n15811_), .ZN(new_n15812_));
  NOR3_X1    g14792(.A1(new_n15773_), .A2(new_n15793_), .A3(new_n15774_), .ZN(new_n15813_));
  AOI22_X1   g14793(.A1(new_n15800_), .A2(new_n15813_), .B1(new_n15785_), .B2(new_n15789_), .ZN(new_n15814_));
  NOR2_X1    g14794(.A1(new_n15713_), .A2(new_n15715_), .ZN(new_n15815_));
  OAI21_X1   g14795(.A1(new_n15731_), .A2(new_n15815_), .B(new_n15771_), .ZN(new_n15816_));
  OAI21_X1   g14796(.A1(new_n15781_), .A2(new_n15787_), .B(new_n15776_), .ZN(new_n15817_));
  OAI21_X1   g14797(.A1(new_n15755_), .A2(new_n15757_), .B(new_n15817_), .ZN(new_n15818_));
  XOR2_X1    g14798(.A1(new_n15818_), .A2(new_n15816_), .Z(new_n15819_));
  NOR3_X1    g14799(.A1(new_n15780_), .A2(new_n15814_), .A3(new_n15819_), .ZN(new_n15820_));
  NAND3_X1   g14800(.A1(new_n15804_), .A2(new_n15812_), .A3(new_n15820_), .ZN(new_n15821_));
  NAND2_X1   g14801(.A1(new_n15818_), .A2(new_n15816_), .ZN(new_n15822_));
  NOR2_X1    g14802(.A1(new_n15780_), .A2(new_n15814_), .ZN(new_n15823_));
  OAI21_X1   g14803(.A1(new_n15816_), .A2(new_n15818_), .B(new_n15823_), .ZN(new_n15824_));
  NAND2_X1   g14804(.A1(new_n15824_), .A2(new_n15822_), .ZN(new_n15825_));
  NAND2_X1   g14805(.A1(new_n15807_), .A2(new_n15809_), .ZN(new_n15826_));
  INV_X1     g14806(.I(new_n15686_), .ZN(new_n15827_));
  INV_X1     g14807(.I(new_n15805_), .ZN(new_n15828_));
  NOR2_X1    g14808(.A1(new_n15828_), .A2(new_n15827_), .ZN(new_n15829_));
  OAI21_X1   g14809(.A1(new_n15807_), .A2(new_n15809_), .B(new_n15829_), .ZN(new_n15830_));
  NAND2_X1   g14810(.A1(new_n15830_), .A2(new_n15826_), .ZN(new_n15831_));
  OAI21_X1   g14811(.A1(new_n15825_), .A2(new_n15831_), .B(new_n15821_), .ZN(new_n15832_));
  NAND2_X1   g14812(.A1(new_n15831_), .A2(new_n15825_), .ZN(new_n15833_));
  NAND2_X1   g14813(.A1(new_n15832_), .A2(new_n15833_), .ZN(new_n15834_));
  NAND2_X1   g14814(.A1(new_n15834_), .A2(new_n15578_), .ZN(new_n15835_));
  INV_X1     g14815(.I(new_n15688_), .ZN(new_n15836_));
  INV_X1     g14816(.I(new_n15763_), .ZN(new_n15837_));
  OAI21_X1   g14817(.A1(new_n15790_), .A2(new_n15795_), .B(new_n15800_), .ZN(new_n15838_));
  NAND2_X1   g14818(.A1(new_n15798_), .A2(new_n15797_), .ZN(new_n15839_));
  NAND2_X1   g14819(.A1(new_n15839_), .A2(new_n15838_), .ZN(new_n15840_));
  AOI22_X1   g14820(.A1(new_n15840_), .A2(new_n15796_), .B1(new_n15780_), .B2(new_n15790_), .ZN(new_n15841_));
  OAI22_X1   g14821(.A1(new_n15761_), .A2(new_n15837_), .B1(new_n15841_), .B2(new_n15836_), .ZN(new_n15842_));
  XOR2_X1    g14822(.A1(new_n15820_), .A2(new_n15811_), .Z(new_n15843_));
  NOR2_X1    g14823(.A1(new_n15842_), .A2(new_n15843_), .ZN(new_n15844_));
  NOR2_X1    g14824(.A1(new_n15812_), .A2(new_n15820_), .ZN(new_n15845_));
  NOR4_X1    g14825(.A1(new_n15811_), .A2(new_n15780_), .A3(new_n15814_), .A4(new_n15819_), .ZN(new_n15846_));
  NOR2_X1    g14826(.A1(new_n15845_), .A2(new_n15846_), .ZN(new_n15847_));
  NOR2_X1    g14827(.A1(new_n15804_), .A2(new_n15847_), .ZN(new_n15848_));
  NOR2_X1    g14828(.A1(new_n15446_), .A2(new_n15445_), .ZN(new_n15849_));
  AOI21_X1   g14829(.A1(new_n15434_), .A2(new_n15440_), .B(new_n15508_), .ZN(new_n15850_));
  INV_X1     g14830(.I(new_n15509_), .ZN(new_n15851_));
  XOR2_X1    g14831(.A1(new_n15544_), .A2(new_n15546_), .Z(new_n15852_));
  AOI22_X1   g14832(.A1(new_n15852_), .A2(new_n15541_), .B1(new_n15526_), .B2(new_n15535_), .ZN(new_n15853_));
  OAI22_X1   g14833(.A1(new_n15851_), .A2(new_n15850_), .B1(new_n15853_), .B2(new_n15849_), .ZN(new_n15854_));
  XNOR2_X1   g14834(.A1(new_n15559_), .A2(new_n15566_), .ZN(new_n15855_));
  NOR2_X1    g14835(.A1(new_n15854_), .A2(new_n15855_), .ZN(new_n15856_));
  NOR2_X1    g14836(.A1(new_n15559_), .A2(new_n15566_), .ZN(new_n15857_));
  INV_X1     g14837(.I(new_n15552_), .ZN(new_n15858_));
  NAND3_X1   g14838(.A1(new_n15858_), .A2(new_n15439_), .A3(new_n15557_), .ZN(new_n15859_));
  INV_X1     g14839(.I(new_n15566_), .ZN(new_n15860_));
  NOR2_X1    g14840(.A1(new_n15860_), .A2(new_n15859_), .ZN(new_n15861_));
  NOR2_X1    g14841(.A1(new_n15861_), .A2(new_n15857_), .ZN(new_n15862_));
  NOR2_X1    g14842(.A1(new_n15550_), .A2(new_n15862_), .ZN(new_n15863_));
  NOR4_X1    g14843(.A1(new_n15844_), .A2(new_n15856_), .A3(new_n15848_), .A4(new_n15863_), .ZN(new_n15864_));
  NOR3_X1    g14844(.A1(new_n15851_), .A2(new_n15850_), .A3(new_n15549_), .ZN(new_n15865_));
  INV_X1     g14845(.I(new_n15865_), .ZN(new_n15866_));
  NAND2_X1   g14846(.A1(new_n15506_), .A2(new_n15507_), .ZN(new_n15867_));
  NAND2_X1   g14847(.A1(new_n15504_), .A2(new_n15867_), .ZN(new_n15868_));
  INV_X1     g14848(.I(new_n15760_), .ZN(new_n15869_));
  NAND2_X1   g14849(.A1(new_n15689_), .A2(new_n15759_), .ZN(new_n15870_));
  NAND2_X1   g14850(.A1(new_n15869_), .A2(new_n15870_), .ZN(new_n15871_));
  NOR2_X1    g14851(.A1(new_n15871_), .A2(new_n15868_), .ZN(new_n15872_));
  NOR2_X1    g14852(.A1(new_n15865_), .A2(new_n15872_), .ZN(new_n15873_));
  INV_X1     g14853(.I(new_n15873_), .ZN(new_n15874_));
  NAND2_X1   g14854(.A1(new_n15865_), .A2(new_n15872_), .ZN(new_n15875_));
  OAI21_X1   g14855(.A1(new_n15837_), .A2(new_n15761_), .B(new_n15841_), .ZN(new_n15876_));
  NAND3_X1   g14856(.A1(new_n15762_), .A2(new_n15803_), .A3(new_n15763_), .ZN(new_n15877_));
  NAND2_X1   g14857(.A1(new_n15876_), .A2(new_n15877_), .ZN(new_n15878_));
  AOI22_X1   g14858(.A1(new_n15874_), .A2(new_n15875_), .B1(new_n15866_), .B2(new_n15878_), .ZN(new_n15879_));
  OAI22_X1   g14859(.A1(new_n15844_), .A2(new_n15848_), .B1(new_n15856_), .B2(new_n15863_), .ZN(new_n15880_));
  AOI21_X1   g14860(.A1(new_n15879_), .A2(new_n15880_), .B(new_n15864_), .ZN(new_n15881_));
  INV_X1     g14861(.I(new_n15845_), .ZN(new_n15882_));
  NAND2_X1   g14862(.A1(new_n15842_), .A2(new_n15882_), .ZN(new_n15883_));
  INV_X1     g14863(.I(new_n15825_), .ZN(new_n15884_));
  AOI21_X1   g14864(.A1(new_n15883_), .A2(new_n15846_), .B(new_n15884_), .ZN(new_n15885_));
  NOR2_X1    g14865(.A1(new_n15821_), .A2(new_n15825_), .ZN(new_n15886_));
  OAI21_X1   g14866(.A1(new_n15885_), .A2(new_n15886_), .B(new_n15831_), .ZN(new_n15887_));
  INV_X1     g14867(.I(new_n15831_), .ZN(new_n15888_));
  NAND2_X1   g14868(.A1(new_n15821_), .A2(new_n15825_), .ZN(new_n15889_));
  NAND4_X1   g14869(.A1(new_n15884_), .A2(new_n15804_), .A3(new_n15812_), .A4(new_n15820_), .ZN(new_n15890_));
  NAND3_X1   g14870(.A1(new_n15889_), .A2(new_n15888_), .A3(new_n15890_), .ZN(new_n15891_));
  NAND2_X1   g14871(.A1(new_n15887_), .A2(new_n15891_), .ZN(new_n15892_));
  INV_X1     g14872(.I(new_n15857_), .ZN(new_n15893_));
  NAND2_X1   g14873(.A1(new_n15854_), .A2(new_n15893_), .ZN(new_n15894_));
  INV_X1     g14874(.I(new_n15571_), .ZN(new_n15895_));
  AOI21_X1   g14875(.A1(new_n15894_), .A2(new_n15861_), .B(new_n15895_), .ZN(new_n15896_));
  NOR2_X1    g14876(.A1(new_n15567_), .A2(new_n15571_), .ZN(new_n15897_));
  OAI21_X1   g14877(.A1(new_n15896_), .A2(new_n15897_), .B(new_n15575_), .ZN(new_n15898_));
  INV_X1     g14878(.I(new_n15575_), .ZN(new_n15899_));
  NAND2_X1   g14879(.A1(new_n15567_), .A2(new_n15571_), .ZN(new_n15900_));
  NAND4_X1   g14880(.A1(new_n15895_), .A2(new_n15550_), .A3(new_n15559_), .A4(new_n15566_), .ZN(new_n15901_));
  NAND3_X1   g14881(.A1(new_n15900_), .A2(new_n15899_), .A3(new_n15901_), .ZN(new_n15902_));
  NAND2_X1   g14882(.A1(new_n15898_), .A2(new_n15902_), .ZN(new_n15903_));
  OAI21_X1   g14883(.A1(new_n15892_), .A2(new_n15903_), .B(new_n15881_), .ZN(new_n15904_));
  XOR2_X1    g14884(.A1(new_n15575_), .A2(new_n15571_), .Z(new_n15905_));
  XOR2_X1    g14885(.A1(new_n15831_), .A2(new_n15825_), .Z(new_n15906_));
  NOR4_X1    g14886(.A1(new_n15906_), .A2(new_n15905_), .A3(new_n15567_), .A4(new_n15821_), .ZN(new_n15907_));
  NAND2_X1   g14887(.A1(new_n15904_), .A2(new_n15907_), .ZN(new_n15908_));
  AND3_X2    g14888(.A1(new_n15576_), .A2(new_n15577_), .A3(new_n15833_), .Z(new_n15909_));
  NAND3_X1   g14889(.A1(new_n15908_), .A2(new_n15832_), .A3(new_n15909_), .ZN(new_n15910_));
  NAND2_X1   g14890(.A1(new_n15910_), .A2(new_n15835_), .ZN(new_n15911_));
  NOR2_X1    g14891(.A1(new_n15329_), .A2(new_n15911_), .ZN(new_n15912_));
  NAND4_X1   g14892(.A1(new_n15303_), .A2(new_n15301_), .A3(new_n15283_), .A4(new_n15281_), .ZN(new_n15913_));
  INV_X1     g14893(.I(new_n15295_), .ZN(new_n15914_));
  INV_X1     g14894(.I(new_n15298_), .ZN(new_n15915_));
  OAI22_X1   g14895(.A1(new_n15915_), .A2(new_n15286_), .B1(new_n15914_), .B2(new_n15293_), .ZN(new_n15916_));
  AOI22_X1   g14896(.A1(new_n15303_), .A2(new_n15301_), .B1(new_n15283_), .B2(new_n15281_), .ZN(new_n15917_));
  OAI21_X1   g14897(.A1(new_n15916_), .A2(new_n15917_), .B(new_n15913_), .ZN(new_n15918_));
  AOI21_X1   g14898(.A1(new_n15312_), .A2(new_n15308_), .B(new_n15253_), .ZN(new_n15919_));
  NOR3_X1    g14899(.A1(new_n15307_), .A2(new_n15309_), .A3(new_n15252_), .ZN(new_n15920_));
  NOR2_X1    g14900(.A1(new_n15920_), .A2(new_n15919_), .ZN(new_n15921_));
  NAND2_X1   g14901(.A1(new_n15317_), .A2(new_n15320_), .ZN(new_n15922_));
  NOR2_X1    g14902(.A1(new_n15921_), .A2(new_n15922_), .ZN(new_n15923_));
  NAND2_X1   g14903(.A1(new_n15310_), .A2(new_n15313_), .ZN(new_n15924_));
  AOI21_X1   g14904(.A1(new_n15319_), .A2(new_n15315_), .B(new_n14989_), .ZN(new_n15925_));
  NOR3_X1    g14905(.A1(new_n15314_), .A2(new_n15316_), .A3(new_n14988_), .ZN(new_n15926_));
  NOR2_X1    g14906(.A1(new_n15926_), .A2(new_n15925_), .ZN(new_n15927_));
  NOR2_X1    g14907(.A1(new_n15924_), .A2(new_n15927_), .ZN(new_n15928_));
  OAI21_X1   g14908(.A1(new_n15928_), .A2(new_n15923_), .B(new_n15918_), .ZN(new_n15929_));
  NOR2_X1    g14909(.A1(new_n15924_), .A2(new_n15922_), .ZN(new_n15930_));
  AOI22_X1   g14910(.A1(new_n15310_), .A2(new_n15313_), .B1(new_n15317_), .B2(new_n15320_), .ZN(new_n15931_));
  OAI21_X1   g14911(.A1(new_n15930_), .A2(new_n15931_), .B(new_n15306_), .ZN(new_n15932_));
  INV_X1     g14912(.I(new_n15843_), .ZN(new_n15933_));
  NAND2_X1   g14913(.A1(new_n15933_), .A2(new_n15804_), .ZN(new_n15934_));
  INV_X1     g14914(.I(new_n15847_), .ZN(new_n15935_));
  NAND2_X1   g14915(.A1(new_n15935_), .A2(new_n15842_), .ZN(new_n15936_));
  XOR2_X1    g14916(.A1(new_n15559_), .A2(new_n15566_), .Z(new_n15937_));
  NAND2_X1   g14917(.A1(new_n15550_), .A2(new_n15937_), .ZN(new_n15938_));
  NAND2_X1   g14918(.A1(new_n15559_), .A2(new_n15566_), .ZN(new_n15939_));
  NAND2_X1   g14919(.A1(new_n15893_), .A2(new_n15939_), .ZN(new_n15940_));
  NAND2_X1   g14920(.A1(new_n15854_), .A2(new_n15940_), .ZN(new_n15941_));
  NAND4_X1   g14921(.A1(new_n15936_), .A2(new_n15934_), .A3(new_n15941_), .A4(new_n15938_), .ZN(new_n15942_));
  INV_X1     g14922(.I(new_n15875_), .ZN(new_n15943_));
  INV_X1     g14923(.I(new_n15878_), .ZN(new_n15944_));
  OAI22_X1   g14924(.A1(new_n15944_), .A2(new_n15865_), .B1(new_n15943_), .B2(new_n15873_), .ZN(new_n15945_));
  AOI22_X1   g14925(.A1(new_n15936_), .A2(new_n15934_), .B1(new_n15941_), .B2(new_n15938_), .ZN(new_n15946_));
  OAI21_X1   g14926(.A1(new_n15945_), .A2(new_n15946_), .B(new_n15942_), .ZN(new_n15947_));
  AOI21_X1   g14927(.A1(new_n15889_), .A2(new_n15890_), .B(new_n15888_), .ZN(new_n15948_));
  NOR3_X1    g14928(.A1(new_n15885_), .A2(new_n15886_), .A3(new_n15831_), .ZN(new_n15949_));
  NOR2_X1    g14929(.A1(new_n15949_), .A2(new_n15948_), .ZN(new_n15950_));
  NOR2_X1    g14930(.A1(new_n15950_), .A2(new_n15903_), .ZN(new_n15951_));
  AOI21_X1   g14931(.A1(new_n15900_), .A2(new_n15901_), .B(new_n15899_), .ZN(new_n15952_));
  NOR3_X1    g14932(.A1(new_n15896_), .A2(new_n15897_), .A3(new_n15575_), .ZN(new_n15953_));
  NOR2_X1    g14933(.A1(new_n15953_), .A2(new_n15952_), .ZN(new_n15954_));
  NOR2_X1    g14934(.A1(new_n15892_), .A2(new_n15954_), .ZN(new_n15955_));
  OAI21_X1   g14935(.A1(new_n15955_), .A2(new_n15951_), .B(new_n15947_), .ZN(new_n15956_));
  NOR2_X1    g14936(.A1(new_n15892_), .A2(new_n15903_), .ZN(new_n15957_));
  AOI22_X1   g14937(.A1(new_n15887_), .A2(new_n15891_), .B1(new_n15898_), .B2(new_n15902_), .ZN(new_n15958_));
  OAI21_X1   g14938(.A1(new_n15957_), .A2(new_n15958_), .B(new_n15881_), .ZN(new_n15959_));
  NAND4_X1   g14939(.A1(new_n15929_), .A2(new_n15956_), .A3(new_n15932_), .A4(new_n15959_), .ZN(new_n15960_));
  NOR2_X1    g14940(.A1(new_n15844_), .A2(new_n15848_), .ZN(new_n15961_));
  NAND2_X1   g14941(.A1(new_n15941_), .A2(new_n15938_), .ZN(new_n15962_));
  NAND2_X1   g14942(.A1(new_n15961_), .A2(new_n15962_), .ZN(new_n15963_));
  NAND2_X1   g14943(.A1(new_n15936_), .A2(new_n15934_), .ZN(new_n15964_));
  NAND3_X1   g14944(.A1(new_n15964_), .A2(new_n15938_), .A3(new_n15941_), .ZN(new_n15965_));
  AOI21_X1   g14945(.A1(new_n15965_), .A2(new_n15963_), .B(new_n15945_), .ZN(new_n15966_));
  AOI21_X1   g14946(.A1(new_n15942_), .A2(new_n15880_), .B(new_n15879_), .ZN(new_n15967_));
  NOR2_X1    g14947(.A1(new_n15270_), .A2(new_n15260_), .ZN(new_n15968_));
  NAND2_X1   g14948(.A1(new_n15968_), .A2(new_n15284_), .ZN(new_n15969_));
  INV_X1     g14949(.I(new_n15284_), .ZN(new_n15970_));
  NAND2_X1   g14950(.A1(new_n15970_), .A2(new_n15304_), .ZN(new_n15971_));
  AOI21_X1   g14951(.A1(new_n15971_), .A2(new_n15969_), .B(new_n15916_), .ZN(new_n15972_));
  AOI21_X1   g14952(.A1(new_n15305_), .A2(new_n15913_), .B(new_n15299_), .ZN(new_n15973_));
  NOR4_X1    g14953(.A1(new_n15972_), .A2(new_n15966_), .A3(new_n15967_), .A4(new_n15973_), .ZN(new_n15974_));
  NOR3_X1    g14954(.A1(new_n15914_), .A2(new_n15293_), .A3(new_n15298_), .ZN(new_n15975_));
  INV_X1     g14955(.I(new_n15975_), .ZN(new_n15976_));
  XOR2_X1    g14956(.A1(new_n15291_), .A2(new_n15289_), .Z(new_n15977_));
  XOR2_X1    g14957(.A1(new_n15868_), .A2(new_n15871_), .Z(new_n15978_));
  NAND2_X1   g14958(.A1(new_n15978_), .A2(new_n15977_), .ZN(new_n15979_));
  INV_X1     g14959(.I(new_n15979_), .ZN(new_n15980_));
  NOR2_X1    g14960(.A1(new_n15975_), .A2(new_n15980_), .ZN(new_n15981_));
  INV_X1     g14961(.I(new_n15981_), .ZN(new_n15982_));
  NAND2_X1   g14962(.A1(new_n15975_), .A2(new_n15980_), .ZN(new_n15983_));
  OAI21_X1   g14963(.A1(new_n15873_), .A2(new_n15943_), .B(new_n15944_), .ZN(new_n15984_));
  NAND3_X1   g14964(.A1(new_n15874_), .A2(new_n15875_), .A3(new_n15878_), .ZN(new_n15985_));
  NAND2_X1   g14965(.A1(new_n15984_), .A2(new_n15985_), .ZN(new_n15986_));
  AOI22_X1   g14966(.A1(new_n15982_), .A2(new_n15983_), .B1(new_n15976_), .B2(new_n15986_), .ZN(new_n15987_));
  OAI22_X1   g14967(.A1(new_n15972_), .A2(new_n15973_), .B1(new_n15966_), .B2(new_n15967_), .ZN(new_n15988_));
  AOI21_X1   g14968(.A1(new_n15988_), .A2(new_n15987_), .B(new_n15974_), .ZN(new_n15989_));
  AOI22_X1   g14969(.A1(new_n15929_), .A2(new_n15932_), .B1(new_n15956_), .B2(new_n15959_), .ZN(new_n15990_));
  OAI21_X1   g14970(.A1(new_n15990_), .A2(new_n15989_), .B(new_n15960_), .ZN(new_n15991_));
  AOI21_X1   g14971(.A1(new_n15921_), .A2(new_n15927_), .B(new_n15918_), .ZN(new_n15992_));
  INV_X1     g14972(.I(new_n15325_), .ZN(new_n15993_));
  OAI21_X1   g14973(.A1(new_n15992_), .A2(new_n15993_), .B(new_n15257_), .ZN(new_n15994_));
  NAND3_X1   g14974(.A1(new_n15322_), .A2(new_n15256_), .A3(new_n15325_), .ZN(new_n15995_));
  AOI21_X1   g14975(.A1(new_n15995_), .A2(new_n15994_), .B(new_n14992_), .ZN(new_n15996_));
  AOI21_X1   g14976(.A1(new_n15322_), .A2(new_n15325_), .B(new_n15256_), .ZN(new_n15997_));
  NOR3_X1    g14977(.A1(new_n15992_), .A2(new_n15257_), .A3(new_n15993_), .ZN(new_n15998_));
  NOR3_X1    g14978(.A1(new_n15997_), .A2(new_n15998_), .A3(new_n14993_), .ZN(new_n15999_));
  INV_X1     g14979(.I(new_n15578_), .ZN(new_n16000_));
  AOI21_X1   g14980(.A1(new_n15950_), .A2(new_n15954_), .B(new_n15947_), .ZN(new_n16001_));
  INV_X1     g14981(.I(new_n15907_), .ZN(new_n16002_));
  OAI21_X1   g14982(.A1(new_n16001_), .A2(new_n16002_), .B(new_n15834_), .ZN(new_n16003_));
  INV_X1     g14983(.I(new_n15834_), .ZN(new_n16004_));
  NAND3_X1   g14984(.A1(new_n15904_), .A2(new_n16004_), .A3(new_n15907_), .ZN(new_n16005_));
  AOI21_X1   g14985(.A1(new_n16003_), .A2(new_n16005_), .B(new_n16000_), .ZN(new_n16006_));
  AOI21_X1   g14986(.A1(new_n15904_), .A2(new_n15907_), .B(new_n16004_), .ZN(new_n16007_));
  NOR3_X1    g14987(.A1(new_n16001_), .A2(new_n15834_), .A3(new_n16002_), .ZN(new_n16008_));
  NOR3_X1    g14988(.A1(new_n16008_), .A2(new_n16007_), .A3(new_n15578_), .ZN(new_n16009_));
  NOR4_X1    g14989(.A1(new_n15996_), .A2(new_n15999_), .A3(new_n16009_), .A4(new_n16006_), .ZN(new_n16010_));
  XOR2_X1    g14990(.A1(new_n15256_), .A2(new_n14992_), .Z(new_n16011_));
  XOR2_X1    g14991(.A1(new_n15834_), .A2(new_n15578_), .Z(new_n16012_));
  NOR4_X1    g14992(.A1(new_n15326_), .A2(new_n15908_), .A3(new_n16011_), .A4(new_n16012_), .ZN(new_n16013_));
  OAI21_X1   g14993(.A1(new_n16010_), .A2(new_n15991_), .B(new_n16013_), .ZN(new_n16014_));
  INV_X1     g14994(.I(new_n16014_), .ZN(new_n16015_));
  NAND4_X1   g14995(.A1(new_n15328_), .A2(new_n15910_), .A3(new_n15258_), .A4(new_n15835_), .ZN(new_n16016_));
  NOR2_X1    g14996(.A1(new_n16015_), .A2(new_n16016_), .ZN(new_n16017_));
  NOR2_X1    g14997(.A1(new_n16017_), .A2(new_n15912_), .ZN(new_n16018_));
  INV_X1     g14998(.I(new_n16018_), .ZN(new_n16019_));
  INV_X1     g14999(.I(\A[550] ), .ZN(new_n16020_));
  NOR2_X1    g15000(.A1(\A[551] ), .A2(\A[552] ), .ZN(new_n16021_));
  NAND2_X1   g15001(.A1(\A[551] ), .A2(\A[552] ), .ZN(new_n16022_));
  AOI21_X1   g15002(.A1(new_n16020_), .A2(new_n16022_), .B(new_n16021_), .ZN(new_n16023_));
  INV_X1     g15003(.I(new_n16023_), .ZN(new_n16024_));
  INV_X1     g15004(.I(\A[547] ), .ZN(new_n16025_));
  NOR2_X1    g15005(.A1(\A[548] ), .A2(\A[549] ), .ZN(new_n16026_));
  NAND2_X1   g15006(.A1(\A[548] ), .A2(\A[549] ), .ZN(new_n16027_));
  AOI21_X1   g15007(.A1(new_n16025_), .A2(new_n16027_), .B(new_n16026_), .ZN(new_n16028_));
  INV_X1     g15008(.I(new_n16028_), .ZN(new_n16029_));
  INV_X1     g15009(.I(\A[548] ), .ZN(new_n16030_));
  NAND2_X1   g15010(.A1(new_n16030_), .A2(\A[549] ), .ZN(new_n16031_));
  INV_X1     g15011(.I(\A[549] ), .ZN(new_n16032_));
  NAND2_X1   g15012(.A1(new_n16032_), .A2(\A[548] ), .ZN(new_n16033_));
  AOI21_X1   g15013(.A1(new_n16031_), .A2(new_n16033_), .B(new_n16025_), .ZN(new_n16034_));
  INV_X1     g15014(.I(new_n16026_), .ZN(new_n16035_));
  AOI21_X1   g15015(.A1(new_n16035_), .A2(new_n16027_), .B(\A[547] ), .ZN(new_n16036_));
  INV_X1     g15016(.I(\A[551] ), .ZN(new_n16037_));
  NAND2_X1   g15017(.A1(new_n16037_), .A2(\A[552] ), .ZN(new_n16038_));
  INV_X1     g15018(.I(\A[552] ), .ZN(new_n16039_));
  NAND2_X1   g15019(.A1(new_n16039_), .A2(\A[551] ), .ZN(new_n16040_));
  AOI21_X1   g15020(.A1(new_n16038_), .A2(new_n16040_), .B(new_n16020_), .ZN(new_n16041_));
  INV_X1     g15021(.I(new_n16021_), .ZN(new_n16042_));
  AOI21_X1   g15022(.A1(new_n16042_), .A2(new_n16022_), .B(\A[550] ), .ZN(new_n16043_));
  NOR4_X1    g15023(.A1(new_n16034_), .A2(new_n16036_), .A3(new_n16043_), .A4(new_n16041_), .ZN(new_n16044_));
  NOR2_X1    g15024(.A1(new_n16044_), .A2(new_n16029_), .ZN(new_n16045_));
  INV_X1     g15025(.I(new_n16045_), .ZN(new_n16046_));
  NAND2_X1   g15026(.A1(new_n16044_), .A2(new_n16029_), .ZN(new_n16047_));
  AOI21_X1   g15027(.A1(new_n16046_), .A2(new_n16047_), .B(new_n16024_), .ZN(new_n16048_));
  INV_X1     g15028(.I(new_n16047_), .ZN(new_n16049_));
  NOR3_X1    g15029(.A1(new_n16049_), .A2(new_n16023_), .A3(new_n16045_), .ZN(new_n16050_));
  NOR2_X1    g15030(.A1(new_n16048_), .A2(new_n16050_), .ZN(new_n16051_));
  INV_X1     g15031(.I(\A[556] ), .ZN(new_n16052_));
  NOR2_X1    g15032(.A1(\A[557] ), .A2(\A[558] ), .ZN(new_n16053_));
  NAND2_X1   g15033(.A1(\A[557] ), .A2(\A[558] ), .ZN(new_n16054_));
  AOI21_X1   g15034(.A1(new_n16052_), .A2(new_n16054_), .B(new_n16053_), .ZN(new_n16055_));
  INV_X1     g15035(.I(new_n16055_), .ZN(new_n16056_));
  INV_X1     g15036(.I(\A[553] ), .ZN(new_n16057_));
  NOR2_X1    g15037(.A1(\A[554] ), .A2(\A[555] ), .ZN(new_n16058_));
  NAND2_X1   g15038(.A1(\A[554] ), .A2(\A[555] ), .ZN(new_n16059_));
  AOI21_X1   g15039(.A1(new_n16057_), .A2(new_n16059_), .B(new_n16058_), .ZN(new_n16060_));
  INV_X1     g15040(.I(new_n16060_), .ZN(new_n16061_));
  NOR2_X1    g15041(.A1(new_n16056_), .A2(new_n16061_), .ZN(new_n16062_));
  INV_X1     g15042(.I(\A[554] ), .ZN(new_n16063_));
  NAND2_X1   g15043(.A1(new_n16063_), .A2(\A[555] ), .ZN(new_n16064_));
  INV_X1     g15044(.I(\A[555] ), .ZN(new_n16065_));
  NAND2_X1   g15045(.A1(new_n16065_), .A2(\A[554] ), .ZN(new_n16066_));
  AOI21_X1   g15046(.A1(new_n16064_), .A2(new_n16066_), .B(new_n16057_), .ZN(new_n16067_));
  INV_X1     g15047(.I(new_n16058_), .ZN(new_n16068_));
  AOI21_X1   g15048(.A1(new_n16068_), .A2(new_n16059_), .B(\A[553] ), .ZN(new_n16069_));
  NOR2_X1    g15049(.A1(new_n16069_), .A2(new_n16067_), .ZN(new_n16070_));
  INV_X1     g15050(.I(\A[558] ), .ZN(new_n16071_));
  NOR2_X1    g15051(.A1(new_n16071_), .A2(\A[557] ), .ZN(new_n16072_));
  INV_X1     g15052(.I(\A[557] ), .ZN(new_n16073_));
  NOR2_X1    g15053(.A1(new_n16073_), .A2(\A[558] ), .ZN(new_n16074_));
  OAI21_X1   g15054(.A1(new_n16072_), .A2(new_n16074_), .B(\A[556] ), .ZN(new_n16075_));
  INV_X1     g15055(.I(new_n16054_), .ZN(new_n16076_));
  OAI21_X1   g15056(.A1(new_n16076_), .A2(new_n16053_), .B(new_n16052_), .ZN(new_n16077_));
  NAND2_X1   g15057(.A1(new_n16075_), .A2(new_n16077_), .ZN(new_n16078_));
  NAND2_X1   g15058(.A1(new_n16070_), .A2(new_n16078_), .ZN(new_n16079_));
  NOR2_X1    g15059(.A1(new_n16065_), .A2(\A[554] ), .ZN(new_n16080_));
  NOR2_X1    g15060(.A1(new_n16063_), .A2(\A[555] ), .ZN(new_n16081_));
  OAI21_X1   g15061(.A1(new_n16080_), .A2(new_n16081_), .B(\A[553] ), .ZN(new_n16082_));
  INV_X1     g15062(.I(new_n16059_), .ZN(new_n16083_));
  OAI21_X1   g15063(.A1(new_n16083_), .A2(new_n16058_), .B(new_n16057_), .ZN(new_n16084_));
  NAND2_X1   g15064(.A1(new_n16082_), .A2(new_n16084_), .ZN(new_n16085_));
  NAND2_X1   g15065(.A1(new_n16073_), .A2(\A[558] ), .ZN(new_n16086_));
  NAND2_X1   g15066(.A1(new_n16071_), .A2(\A[557] ), .ZN(new_n16087_));
  AOI21_X1   g15067(.A1(new_n16086_), .A2(new_n16087_), .B(new_n16052_), .ZN(new_n16088_));
  INV_X1     g15068(.I(new_n16053_), .ZN(new_n16089_));
  AOI21_X1   g15069(.A1(new_n16089_), .A2(new_n16054_), .B(\A[556] ), .ZN(new_n16090_));
  NOR2_X1    g15070(.A1(new_n16090_), .A2(new_n16088_), .ZN(new_n16091_));
  NAND2_X1   g15071(.A1(new_n16091_), .A2(new_n16085_), .ZN(new_n16092_));
  NAND2_X1   g15072(.A1(new_n16079_), .A2(new_n16092_), .ZN(new_n16093_));
  NAND2_X1   g15073(.A1(new_n16093_), .A2(new_n16062_), .ZN(new_n16094_));
  NOR2_X1    g15074(.A1(new_n16085_), .A2(new_n16078_), .ZN(new_n16095_));
  NOR2_X1    g15075(.A1(new_n16095_), .A2(new_n16061_), .ZN(new_n16096_));
  NAND2_X1   g15076(.A1(new_n16070_), .A2(new_n16091_), .ZN(new_n16097_));
  NOR2_X1    g15077(.A1(new_n16097_), .A2(new_n16060_), .ZN(new_n16098_));
  OAI21_X1   g15078(.A1(new_n16096_), .A2(new_n16098_), .B(new_n16055_), .ZN(new_n16099_));
  NAND2_X1   g15079(.A1(new_n16097_), .A2(new_n16060_), .ZN(new_n16100_));
  NAND2_X1   g15080(.A1(new_n16095_), .A2(new_n16061_), .ZN(new_n16101_));
  NAND3_X1   g15081(.A1(new_n16101_), .A2(new_n16100_), .A3(new_n16056_), .ZN(new_n16102_));
  NAND3_X1   g15082(.A1(new_n16099_), .A2(new_n16102_), .A3(new_n16094_), .ZN(new_n16103_));
  INV_X1     g15083(.I(new_n16062_), .ZN(new_n16104_));
  NOR2_X1    g15084(.A1(new_n16097_), .A2(new_n16104_), .ZN(new_n16105_));
  NOR2_X1    g15085(.A1(new_n16070_), .A2(new_n16091_), .ZN(new_n16106_));
  NOR2_X1    g15086(.A1(new_n16106_), .A2(new_n16095_), .ZN(new_n16107_));
  NOR2_X1    g15087(.A1(new_n16036_), .A2(new_n16034_), .ZN(new_n16108_));
  NOR2_X1    g15088(.A1(new_n16043_), .A2(new_n16041_), .ZN(new_n16109_));
  NOR2_X1    g15089(.A1(new_n16108_), .A2(new_n16109_), .ZN(new_n16110_));
  NOR2_X1    g15090(.A1(new_n16110_), .A2(new_n16044_), .ZN(new_n16111_));
  NAND2_X1   g15091(.A1(new_n16108_), .A2(new_n16109_), .ZN(new_n16112_));
  NAND2_X1   g15092(.A1(new_n16023_), .A2(new_n16028_), .ZN(new_n16113_));
  NOR2_X1    g15093(.A1(new_n16112_), .A2(new_n16113_), .ZN(new_n16114_));
  NAND4_X1   g15094(.A1(new_n16105_), .A2(new_n16107_), .A3(new_n16111_), .A4(new_n16114_), .ZN(new_n16115_));
  NOR2_X1    g15095(.A1(new_n16103_), .A2(new_n16115_), .ZN(new_n16116_));
  AOI21_X1   g15096(.A1(new_n16079_), .A2(new_n16092_), .B(new_n16104_), .ZN(new_n16117_));
  AOI21_X1   g15097(.A1(new_n16101_), .A2(new_n16100_), .B(new_n16056_), .ZN(new_n16118_));
  NOR3_X1    g15098(.A1(new_n16096_), .A2(new_n16098_), .A3(new_n16055_), .ZN(new_n16119_));
  NOR3_X1    g15099(.A1(new_n16118_), .A2(new_n16119_), .A3(new_n16117_), .ZN(new_n16120_));
  NAND2_X1   g15100(.A1(new_n16107_), .A2(new_n16105_), .ZN(new_n16121_));
  NAND2_X1   g15101(.A1(new_n16111_), .A2(new_n16114_), .ZN(new_n16122_));
  NOR2_X1    g15102(.A1(new_n16121_), .A2(new_n16122_), .ZN(new_n16123_));
  NOR2_X1    g15103(.A1(new_n16120_), .A2(new_n16123_), .ZN(new_n16124_));
  OAI21_X1   g15104(.A1(new_n16124_), .A2(new_n16116_), .B(new_n16051_), .ZN(new_n16125_));
  NAND2_X1   g15105(.A1(new_n16103_), .A2(new_n16123_), .ZN(new_n16126_));
  NAND2_X1   g15106(.A1(new_n16099_), .A2(new_n16102_), .ZN(new_n16127_));
  NAND3_X1   g15107(.A1(new_n16107_), .A2(new_n16105_), .A3(new_n16111_), .ZN(new_n16128_));
  NOR3_X1    g15108(.A1(new_n16117_), .A2(new_n16112_), .A3(new_n16113_), .ZN(new_n16129_));
  OAI21_X1   g15109(.A1(new_n16127_), .A2(new_n16128_), .B(new_n16129_), .ZN(new_n16130_));
  NAND3_X1   g15110(.A1(new_n16130_), .A2(new_n16126_), .A3(new_n16051_), .ZN(new_n16131_));
  NAND2_X1   g15111(.A1(new_n16125_), .A2(new_n16131_), .ZN(new_n16132_));
  XNOR2_X1   g15112(.A1(new_n16121_), .A2(new_n16122_), .ZN(new_n16133_));
  INV_X1     g15113(.I(\A[541] ), .ZN(new_n16134_));
  INV_X1     g15114(.I(\A[542] ), .ZN(new_n16135_));
  NAND2_X1   g15115(.A1(new_n16135_), .A2(\A[543] ), .ZN(new_n16136_));
  INV_X1     g15116(.I(\A[543] ), .ZN(new_n16137_));
  NAND2_X1   g15117(.A1(new_n16137_), .A2(\A[542] ), .ZN(new_n16138_));
  AOI21_X1   g15118(.A1(new_n16136_), .A2(new_n16138_), .B(new_n16134_), .ZN(new_n16139_));
  NOR2_X1    g15119(.A1(\A[542] ), .A2(\A[543] ), .ZN(new_n16140_));
  INV_X1     g15120(.I(new_n16140_), .ZN(new_n16141_));
  NAND2_X1   g15121(.A1(\A[542] ), .A2(\A[543] ), .ZN(new_n16142_));
  AOI21_X1   g15122(.A1(new_n16141_), .A2(new_n16142_), .B(\A[541] ), .ZN(new_n16143_));
  NOR2_X1    g15123(.A1(new_n16143_), .A2(new_n16139_), .ZN(new_n16144_));
  INV_X1     g15124(.I(\A[544] ), .ZN(new_n16145_));
  INV_X1     g15125(.I(\A[545] ), .ZN(new_n16146_));
  NAND2_X1   g15126(.A1(new_n16146_), .A2(\A[546] ), .ZN(new_n16147_));
  INV_X1     g15127(.I(\A[546] ), .ZN(new_n16148_));
  NAND2_X1   g15128(.A1(new_n16148_), .A2(\A[545] ), .ZN(new_n16149_));
  AOI21_X1   g15129(.A1(new_n16147_), .A2(new_n16149_), .B(new_n16145_), .ZN(new_n16150_));
  NOR2_X1    g15130(.A1(\A[545] ), .A2(\A[546] ), .ZN(new_n16151_));
  INV_X1     g15131(.I(new_n16151_), .ZN(new_n16152_));
  NAND2_X1   g15132(.A1(\A[545] ), .A2(\A[546] ), .ZN(new_n16153_));
  AOI21_X1   g15133(.A1(new_n16152_), .A2(new_n16153_), .B(\A[544] ), .ZN(new_n16154_));
  NOR2_X1    g15134(.A1(new_n16154_), .A2(new_n16150_), .ZN(new_n16155_));
  NAND2_X1   g15135(.A1(new_n16144_), .A2(new_n16155_), .ZN(new_n16156_));
  AOI21_X1   g15136(.A1(new_n16145_), .A2(new_n16153_), .B(new_n16151_), .ZN(new_n16157_));
  INV_X1     g15137(.I(new_n16157_), .ZN(new_n16158_));
  AOI21_X1   g15138(.A1(new_n16134_), .A2(new_n16142_), .B(new_n16140_), .ZN(new_n16159_));
  INV_X1     g15139(.I(new_n16159_), .ZN(new_n16160_));
  NOR2_X1    g15140(.A1(new_n16158_), .A2(new_n16160_), .ZN(new_n16161_));
  INV_X1     g15141(.I(new_n16161_), .ZN(new_n16162_));
  NOR2_X1    g15142(.A1(new_n16156_), .A2(new_n16162_), .ZN(new_n16163_));
  NOR2_X1    g15143(.A1(new_n16137_), .A2(\A[542] ), .ZN(new_n16164_));
  NOR2_X1    g15144(.A1(new_n16135_), .A2(\A[543] ), .ZN(new_n16165_));
  OAI21_X1   g15145(.A1(new_n16164_), .A2(new_n16165_), .B(\A[541] ), .ZN(new_n16166_));
  INV_X1     g15146(.I(new_n16142_), .ZN(new_n16167_));
  OAI21_X1   g15147(.A1(new_n16167_), .A2(new_n16140_), .B(new_n16134_), .ZN(new_n16168_));
  NAND2_X1   g15148(.A1(new_n16166_), .A2(new_n16168_), .ZN(new_n16169_));
  NOR2_X1    g15149(.A1(new_n16148_), .A2(\A[545] ), .ZN(new_n16170_));
  NOR2_X1    g15150(.A1(new_n16146_), .A2(\A[546] ), .ZN(new_n16171_));
  OAI21_X1   g15151(.A1(new_n16170_), .A2(new_n16171_), .B(\A[544] ), .ZN(new_n16172_));
  INV_X1     g15152(.I(new_n16153_), .ZN(new_n16173_));
  OAI21_X1   g15153(.A1(new_n16173_), .A2(new_n16151_), .B(new_n16145_), .ZN(new_n16174_));
  NAND2_X1   g15154(.A1(new_n16172_), .A2(new_n16174_), .ZN(new_n16175_));
  NAND2_X1   g15155(.A1(new_n16169_), .A2(new_n16175_), .ZN(new_n16176_));
  NAND3_X1   g15156(.A1(new_n16163_), .A2(new_n16156_), .A3(new_n16176_), .ZN(new_n16177_));
  INV_X1     g15157(.I(\A[535] ), .ZN(new_n16178_));
  INV_X1     g15158(.I(\A[536] ), .ZN(new_n16179_));
  NAND2_X1   g15159(.A1(new_n16179_), .A2(\A[537] ), .ZN(new_n16180_));
  INV_X1     g15160(.I(\A[537] ), .ZN(new_n16181_));
  NAND2_X1   g15161(.A1(new_n16181_), .A2(\A[536] ), .ZN(new_n16182_));
  AOI21_X1   g15162(.A1(new_n16180_), .A2(new_n16182_), .B(new_n16178_), .ZN(new_n16183_));
  NAND2_X1   g15163(.A1(new_n16179_), .A2(new_n16181_), .ZN(new_n16184_));
  NAND2_X1   g15164(.A1(\A[536] ), .A2(\A[537] ), .ZN(new_n16185_));
  AOI21_X1   g15165(.A1(new_n16184_), .A2(new_n16185_), .B(\A[535] ), .ZN(new_n16186_));
  INV_X1     g15166(.I(\A[538] ), .ZN(new_n16187_));
  INV_X1     g15167(.I(\A[539] ), .ZN(new_n16188_));
  NAND2_X1   g15168(.A1(new_n16188_), .A2(\A[540] ), .ZN(new_n16189_));
  INV_X1     g15169(.I(\A[540] ), .ZN(new_n16190_));
  NAND2_X1   g15170(.A1(new_n16190_), .A2(\A[539] ), .ZN(new_n16191_));
  AOI21_X1   g15171(.A1(new_n16189_), .A2(new_n16191_), .B(new_n16187_), .ZN(new_n16192_));
  NAND2_X1   g15172(.A1(new_n16188_), .A2(new_n16190_), .ZN(new_n16193_));
  NAND2_X1   g15173(.A1(\A[539] ), .A2(\A[540] ), .ZN(new_n16194_));
  AOI21_X1   g15174(.A1(new_n16193_), .A2(new_n16194_), .B(\A[538] ), .ZN(new_n16195_));
  NOR4_X1    g15175(.A1(new_n16183_), .A2(new_n16186_), .A3(new_n16195_), .A4(new_n16192_), .ZN(new_n16196_));
  NAND2_X1   g15176(.A1(new_n16194_), .A2(new_n16187_), .ZN(new_n16197_));
  NAND2_X1   g15177(.A1(new_n16197_), .A2(new_n16193_), .ZN(new_n16198_));
  NAND2_X1   g15178(.A1(new_n16185_), .A2(new_n16178_), .ZN(new_n16199_));
  NAND2_X1   g15179(.A1(new_n16199_), .A2(new_n16184_), .ZN(new_n16200_));
  NOR2_X1    g15180(.A1(new_n16198_), .A2(new_n16200_), .ZN(new_n16201_));
  NOR2_X1    g15181(.A1(new_n16186_), .A2(new_n16183_), .ZN(new_n16202_));
  NOR2_X1    g15182(.A1(new_n16195_), .A2(new_n16192_), .ZN(new_n16203_));
  NOR2_X1    g15183(.A1(new_n16202_), .A2(new_n16203_), .ZN(new_n16204_));
  NAND2_X1   g15184(.A1(new_n16133_), .A2(new_n16177_), .ZN(new_n16205_));
  NAND2_X1   g15185(.A1(new_n16132_), .A2(new_n16205_), .ZN(new_n16206_));
  XOR2_X1    g15186(.A1(new_n16121_), .A2(new_n16122_), .Z(new_n16207_));
  NOR2_X1    g15187(.A1(new_n16169_), .A2(new_n16175_), .ZN(new_n16208_));
  NAND2_X1   g15188(.A1(new_n16208_), .A2(new_n16161_), .ZN(new_n16209_));
  NAND2_X1   g15189(.A1(new_n16156_), .A2(new_n16176_), .ZN(new_n16210_));
  NOR2_X1    g15190(.A1(new_n16210_), .A2(new_n16209_), .ZN(new_n16211_));
  NOR2_X1    g15191(.A1(new_n16207_), .A2(new_n16211_), .ZN(new_n16212_));
  NAND3_X1   g15192(.A1(new_n16125_), .A2(new_n16212_), .A3(new_n16131_), .ZN(new_n16213_));
  NOR2_X1    g15193(.A1(new_n16204_), .A2(new_n16196_), .ZN(new_n16214_));
  INV_X1     g15194(.I(new_n16214_), .ZN(new_n16215_));
  NAND2_X1   g15195(.A1(new_n16156_), .A2(new_n16159_), .ZN(new_n16216_));
  NAND2_X1   g15196(.A1(new_n16208_), .A2(new_n16160_), .ZN(new_n16217_));
  AOI21_X1   g15197(.A1(new_n16217_), .A2(new_n16216_), .B(new_n16158_), .ZN(new_n16218_));
  NOR2_X1    g15198(.A1(new_n16208_), .A2(new_n16160_), .ZN(new_n16219_));
  NOR2_X1    g15199(.A1(new_n16156_), .A2(new_n16159_), .ZN(new_n16220_));
  NOR3_X1    g15200(.A1(new_n16219_), .A2(new_n16220_), .A3(new_n16157_), .ZN(new_n16221_));
  NOR4_X1    g15201(.A1(new_n16218_), .A2(new_n16221_), .A3(new_n16177_), .A4(new_n16215_), .ZN(new_n16222_));
  NAND2_X1   g15202(.A1(new_n16202_), .A2(new_n16203_), .ZN(new_n16223_));
  INV_X1     g15203(.I(new_n16201_), .ZN(new_n16224_));
  NOR2_X1    g15204(.A1(new_n16223_), .A2(new_n16224_), .ZN(new_n16225_));
  NOR2_X1    g15205(.A1(new_n16155_), .A2(new_n16169_), .ZN(new_n16226_));
  NOR2_X1    g15206(.A1(new_n16144_), .A2(new_n16175_), .ZN(new_n16227_));
  OAI21_X1   g15207(.A1(new_n16226_), .A2(new_n16227_), .B(new_n16161_), .ZN(new_n16228_));
  NAND2_X1   g15208(.A1(new_n16228_), .A2(new_n16225_), .ZN(new_n16229_));
  NOR2_X1    g15209(.A1(new_n16222_), .A2(new_n16229_), .ZN(new_n16230_));
  INV_X1     g15210(.I(new_n16198_), .ZN(new_n16231_));
  NOR2_X1    g15211(.A1(new_n16196_), .A2(new_n16200_), .ZN(new_n16232_));
  INV_X1     g15212(.I(new_n16200_), .ZN(new_n16233_));
  NOR2_X1    g15213(.A1(new_n16223_), .A2(new_n16233_), .ZN(new_n16234_));
  OAI21_X1   g15214(.A1(new_n16234_), .A2(new_n16232_), .B(new_n16231_), .ZN(new_n16235_));
  NAND2_X1   g15215(.A1(new_n16223_), .A2(new_n16233_), .ZN(new_n16236_));
  NAND2_X1   g15216(.A1(new_n16196_), .A2(new_n16200_), .ZN(new_n16237_));
  NAND3_X1   g15217(.A1(new_n16236_), .A2(new_n16198_), .A3(new_n16237_), .ZN(new_n16238_));
  NAND2_X1   g15218(.A1(new_n16235_), .A2(new_n16238_), .ZN(new_n16239_));
  NAND2_X1   g15219(.A1(new_n16230_), .A2(new_n16239_), .ZN(new_n16240_));
  NOR2_X1    g15220(.A1(new_n16210_), .A2(new_n16209_), .ZN(new_n16241_));
  NAND3_X1   g15221(.A1(new_n16241_), .A2(new_n16225_), .A3(new_n16214_), .ZN(new_n16242_));
  NAND2_X1   g15222(.A1(new_n16242_), .A2(new_n16239_), .ZN(new_n16243_));
  OAI21_X1   g15223(.A1(new_n16219_), .A2(new_n16220_), .B(new_n16157_), .ZN(new_n16244_));
  NAND3_X1   g15224(.A1(new_n16217_), .A2(new_n16216_), .A3(new_n16158_), .ZN(new_n16245_));
  AND3_X2    g15225(.A1(new_n16244_), .A2(new_n16245_), .A3(new_n16228_), .Z(new_n16246_));
  NOR2_X1    g15226(.A1(new_n16242_), .A2(new_n16239_), .ZN(new_n16247_));
  NOR2_X1    g15227(.A1(new_n16247_), .A2(new_n16246_), .ZN(new_n16248_));
  NAND3_X1   g15228(.A1(new_n16244_), .A2(new_n16245_), .A3(new_n16228_), .ZN(new_n16249_));
  NOR3_X1    g15229(.A1(new_n16249_), .A2(new_n16242_), .A3(new_n16239_), .ZN(new_n16250_));
  OAI21_X1   g15230(.A1(new_n16248_), .A2(new_n16250_), .B(new_n16243_), .ZN(new_n16251_));
  NAND2_X1   g15231(.A1(new_n16251_), .A2(new_n16240_), .ZN(new_n16252_));
  AOI22_X1   g15232(.A1(new_n16206_), .A2(new_n16213_), .B1(new_n16252_), .B2(new_n16132_), .ZN(new_n16253_));
  INV_X1     g15233(.I(new_n16130_), .ZN(new_n16254_));
  AOI21_X1   g15234(.A1(new_n16103_), .A2(new_n16123_), .B(new_n16051_), .ZN(new_n16255_));
  NOR2_X1    g15235(.A1(new_n16055_), .A2(new_n16060_), .ZN(new_n16256_));
  OAI21_X1   g15236(.A1(new_n16097_), .A2(new_n16256_), .B(new_n16104_), .ZN(new_n16257_));
  NOR2_X1    g15237(.A1(new_n16023_), .A2(new_n16028_), .ZN(new_n16258_));
  OAI21_X1   g15238(.A1(new_n16112_), .A2(new_n16258_), .B(new_n16113_), .ZN(new_n16259_));
  XOR2_X1    g15239(.A1(new_n16257_), .A2(new_n16259_), .Z(new_n16260_));
  NOR3_X1    g15240(.A1(new_n16254_), .A2(new_n16255_), .A3(new_n16260_), .ZN(new_n16261_));
  NOR4_X1    g15241(.A1(new_n16177_), .A2(new_n16223_), .A3(new_n16224_), .A4(new_n16215_), .ZN(new_n16262_));
  AOI22_X1   g15242(.A1(new_n16262_), .A2(new_n16249_), .B1(new_n16235_), .B2(new_n16238_), .ZN(new_n16263_));
  NOR2_X1    g15243(.A1(new_n16157_), .A2(new_n16159_), .ZN(new_n16264_));
  OAI21_X1   g15244(.A1(new_n16156_), .A2(new_n16264_), .B(new_n16162_), .ZN(new_n16265_));
  NOR2_X1    g15245(.A1(new_n16231_), .A2(new_n16233_), .ZN(new_n16266_));
  OAI21_X1   g15246(.A1(new_n16223_), .A2(new_n16266_), .B(new_n16224_), .ZN(new_n16267_));
  XOR2_X1    g15247(.A1(new_n16265_), .A2(new_n16267_), .Z(new_n16268_));
  NOR3_X1    g15248(.A1(new_n16263_), .A2(new_n16230_), .A3(new_n16268_), .ZN(new_n16269_));
  NAND3_X1   g15249(.A1(new_n16253_), .A2(new_n16261_), .A3(new_n16269_), .ZN(new_n16270_));
  NAND2_X1   g15250(.A1(new_n16265_), .A2(new_n16267_), .ZN(new_n16271_));
  NOR2_X1    g15251(.A1(new_n16263_), .A2(new_n16230_), .ZN(new_n16272_));
  OAI21_X1   g15252(.A1(new_n16265_), .A2(new_n16267_), .B(new_n16272_), .ZN(new_n16273_));
  NAND2_X1   g15253(.A1(new_n16273_), .A2(new_n16271_), .ZN(new_n16274_));
  NAND2_X1   g15254(.A1(new_n16257_), .A2(new_n16259_), .ZN(new_n16275_));
  NOR2_X1    g15255(.A1(new_n16254_), .A2(new_n16255_), .ZN(new_n16276_));
  OAI21_X1   g15256(.A1(new_n16257_), .A2(new_n16259_), .B(new_n16276_), .ZN(new_n16277_));
  NAND2_X1   g15257(.A1(new_n16277_), .A2(new_n16275_), .ZN(new_n16278_));
  OAI21_X1   g15258(.A1(new_n16274_), .A2(new_n16278_), .B(new_n16270_), .ZN(new_n16279_));
  INV_X1     g15259(.I(new_n16279_), .ZN(new_n16280_));
  INV_X1     g15260(.I(new_n16274_), .ZN(new_n16281_));
  INV_X1     g15261(.I(new_n16278_), .ZN(new_n16282_));
  NOR2_X1    g15262(.A1(new_n16282_), .A2(new_n16281_), .ZN(new_n16283_));
  NOR2_X1    g15263(.A1(new_n16280_), .A2(new_n16283_), .ZN(new_n16284_));
  INV_X1     g15264(.I(new_n16284_), .ZN(new_n16285_));
  INV_X1     g15265(.I(\A[526] ), .ZN(new_n16286_));
  NOR2_X1    g15266(.A1(\A[527] ), .A2(\A[528] ), .ZN(new_n16287_));
  NAND2_X1   g15267(.A1(\A[527] ), .A2(\A[528] ), .ZN(new_n16288_));
  AOI21_X1   g15268(.A1(new_n16286_), .A2(new_n16288_), .B(new_n16287_), .ZN(new_n16289_));
  INV_X1     g15269(.I(new_n16289_), .ZN(new_n16290_));
  INV_X1     g15270(.I(\A[523] ), .ZN(new_n16291_));
  NOR2_X1    g15271(.A1(\A[524] ), .A2(\A[525] ), .ZN(new_n16292_));
  NAND2_X1   g15272(.A1(\A[524] ), .A2(\A[525] ), .ZN(new_n16293_));
  AOI21_X1   g15273(.A1(new_n16291_), .A2(new_n16293_), .B(new_n16292_), .ZN(new_n16294_));
  INV_X1     g15274(.I(new_n16294_), .ZN(new_n16295_));
  INV_X1     g15275(.I(\A[524] ), .ZN(new_n16296_));
  NAND2_X1   g15276(.A1(new_n16296_), .A2(\A[525] ), .ZN(new_n16297_));
  INV_X1     g15277(.I(\A[525] ), .ZN(new_n16298_));
  NAND2_X1   g15278(.A1(new_n16298_), .A2(\A[524] ), .ZN(new_n16299_));
  AOI21_X1   g15279(.A1(new_n16297_), .A2(new_n16299_), .B(new_n16291_), .ZN(new_n16300_));
  INV_X1     g15280(.I(new_n16292_), .ZN(new_n16301_));
  AOI21_X1   g15281(.A1(new_n16301_), .A2(new_n16293_), .B(\A[523] ), .ZN(new_n16302_));
  INV_X1     g15282(.I(\A[527] ), .ZN(new_n16303_));
  NAND2_X1   g15283(.A1(new_n16303_), .A2(\A[528] ), .ZN(new_n16304_));
  INV_X1     g15284(.I(\A[528] ), .ZN(new_n16305_));
  NAND2_X1   g15285(.A1(new_n16305_), .A2(\A[527] ), .ZN(new_n16306_));
  AOI21_X1   g15286(.A1(new_n16304_), .A2(new_n16306_), .B(new_n16286_), .ZN(new_n16307_));
  INV_X1     g15287(.I(new_n16287_), .ZN(new_n16308_));
  AOI21_X1   g15288(.A1(new_n16308_), .A2(new_n16288_), .B(\A[526] ), .ZN(new_n16309_));
  NOR4_X1    g15289(.A1(new_n16300_), .A2(new_n16302_), .A3(new_n16309_), .A4(new_n16307_), .ZN(new_n16310_));
  NOR2_X1    g15290(.A1(new_n16310_), .A2(new_n16295_), .ZN(new_n16311_));
  INV_X1     g15291(.I(new_n16311_), .ZN(new_n16312_));
  NAND2_X1   g15292(.A1(new_n16310_), .A2(new_n16295_), .ZN(new_n16313_));
  AOI21_X1   g15293(.A1(new_n16312_), .A2(new_n16313_), .B(new_n16290_), .ZN(new_n16314_));
  INV_X1     g15294(.I(new_n16313_), .ZN(new_n16315_));
  NOR3_X1    g15295(.A1(new_n16315_), .A2(new_n16289_), .A3(new_n16311_), .ZN(new_n16316_));
  NOR2_X1    g15296(.A1(new_n16314_), .A2(new_n16316_), .ZN(new_n16317_));
  INV_X1     g15297(.I(new_n16317_), .ZN(new_n16318_));
  INV_X1     g15298(.I(\A[532] ), .ZN(new_n16319_));
  NOR2_X1    g15299(.A1(\A[533] ), .A2(\A[534] ), .ZN(new_n16320_));
  NAND2_X1   g15300(.A1(\A[533] ), .A2(\A[534] ), .ZN(new_n16321_));
  AOI21_X1   g15301(.A1(new_n16319_), .A2(new_n16321_), .B(new_n16320_), .ZN(new_n16322_));
  INV_X1     g15302(.I(new_n16322_), .ZN(new_n16323_));
  INV_X1     g15303(.I(\A[529] ), .ZN(new_n16324_));
  NOR2_X1    g15304(.A1(\A[530] ), .A2(\A[531] ), .ZN(new_n16325_));
  NAND2_X1   g15305(.A1(\A[530] ), .A2(\A[531] ), .ZN(new_n16326_));
  AOI21_X1   g15306(.A1(new_n16324_), .A2(new_n16326_), .B(new_n16325_), .ZN(new_n16327_));
  INV_X1     g15307(.I(new_n16327_), .ZN(new_n16328_));
  NOR2_X1    g15308(.A1(new_n16323_), .A2(new_n16328_), .ZN(new_n16329_));
  INV_X1     g15309(.I(\A[530] ), .ZN(new_n16330_));
  NAND2_X1   g15310(.A1(new_n16330_), .A2(\A[531] ), .ZN(new_n16331_));
  INV_X1     g15311(.I(\A[531] ), .ZN(new_n16332_));
  NAND2_X1   g15312(.A1(new_n16332_), .A2(\A[530] ), .ZN(new_n16333_));
  AOI21_X1   g15313(.A1(new_n16331_), .A2(new_n16333_), .B(new_n16324_), .ZN(new_n16334_));
  INV_X1     g15314(.I(new_n16325_), .ZN(new_n16335_));
  AOI21_X1   g15315(.A1(new_n16335_), .A2(new_n16326_), .B(\A[529] ), .ZN(new_n16336_));
  NOR2_X1    g15316(.A1(new_n16336_), .A2(new_n16334_), .ZN(new_n16337_));
  INV_X1     g15317(.I(\A[534] ), .ZN(new_n16338_));
  NOR2_X1    g15318(.A1(new_n16338_), .A2(\A[533] ), .ZN(new_n16339_));
  INV_X1     g15319(.I(\A[533] ), .ZN(new_n16340_));
  NOR2_X1    g15320(.A1(new_n16340_), .A2(\A[534] ), .ZN(new_n16341_));
  OAI21_X1   g15321(.A1(new_n16339_), .A2(new_n16341_), .B(\A[532] ), .ZN(new_n16342_));
  INV_X1     g15322(.I(new_n16321_), .ZN(new_n16343_));
  OAI21_X1   g15323(.A1(new_n16343_), .A2(new_n16320_), .B(new_n16319_), .ZN(new_n16344_));
  NAND2_X1   g15324(.A1(new_n16342_), .A2(new_n16344_), .ZN(new_n16345_));
  NAND2_X1   g15325(.A1(new_n16337_), .A2(new_n16345_), .ZN(new_n16346_));
  NOR2_X1    g15326(.A1(new_n16332_), .A2(\A[530] ), .ZN(new_n16347_));
  NOR2_X1    g15327(.A1(new_n16330_), .A2(\A[531] ), .ZN(new_n16348_));
  OAI21_X1   g15328(.A1(new_n16347_), .A2(new_n16348_), .B(\A[529] ), .ZN(new_n16349_));
  INV_X1     g15329(.I(new_n16326_), .ZN(new_n16350_));
  OAI21_X1   g15330(.A1(new_n16350_), .A2(new_n16325_), .B(new_n16324_), .ZN(new_n16351_));
  NAND2_X1   g15331(.A1(new_n16349_), .A2(new_n16351_), .ZN(new_n16352_));
  NAND2_X1   g15332(.A1(new_n16340_), .A2(\A[534] ), .ZN(new_n16353_));
  NAND2_X1   g15333(.A1(new_n16338_), .A2(\A[533] ), .ZN(new_n16354_));
  AOI21_X1   g15334(.A1(new_n16353_), .A2(new_n16354_), .B(new_n16319_), .ZN(new_n16355_));
  INV_X1     g15335(.I(new_n16320_), .ZN(new_n16356_));
  AOI21_X1   g15336(.A1(new_n16356_), .A2(new_n16321_), .B(\A[532] ), .ZN(new_n16357_));
  NOR2_X1    g15337(.A1(new_n16357_), .A2(new_n16355_), .ZN(new_n16358_));
  NAND2_X1   g15338(.A1(new_n16358_), .A2(new_n16352_), .ZN(new_n16359_));
  NAND2_X1   g15339(.A1(new_n16346_), .A2(new_n16359_), .ZN(new_n16360_));
  NAND2_X1   g15340(.A1(new_n16360_), .A2(new_n16329_), .ZN(new_n16361_));
  NOR2_X1    g15341(.A1(new_n16352_), .A2(new_n16345_), .ZN(new_n16362_));
  NOR2_X1    g15342(.A1(new_n16362_), .A2(new_n16328_), .ZN(new_n16363_));
  NAND2_X1   g15343(.A1(new_n16337_), .A2(new_n16358_), .ZN(new_n16364_));
  NOR2_X1    g15344(.A1(new_n16364_), .A2(new_n16327_), .ZN(new_n16365_));
  OAI21_X1   g15345(.A1(new_n16363_), .A2(new_n16365_), .B(new_n16322_), .ZN(new_n16366_));
  NAND2_X1   g15346(.A1(new_n16364_), .A2(new_n16327_), .ZN(new_n16367_));
  NAND2_X1   g15347(.A1(new_n16362_), .A2(new_n16328_), .ZN(new_n16368_));
  NAND3_X1   g15348(.A1(new_n16368_), .A2(new_n16367_), .A3(new_n16323_), .ZN(new_n16369_));
  NAND3_X1   g15349(.A1(new_n16366_), .A2(new_n16369_), .A3(new_n16361_), .ZN(new_n16370_));
  INV_X1     g15350(.I(new_n16329_), .ZN(new_n16371_));
  NOR2_X1    g15351(.A1(new_n16364_), .A2(new_n16371_), .ZN(new_n16372_));
  NOR2_X1    g15352(.A1(new_n16337_), .A2(new_n16358_), .ZN(new_n16373_));
  NOR2_X1    g15353(.A1(new_n16373_), .A2(new_n16362_), .ZN(new_n16374_));
  NOR2_X1    g15354(.A1(new_n16302_), .A2(new_n16300_), .ZN(new_n16375_));
  NOR2_X1    g15355(.A1(new_n16309_), .A2(new_n16307_), .ZN(new_n16376_));
  NOR2_X1    g15356(.A1(new_n16375_), .A2(new_n16376_), .ZN(new_n16377_));
  NOR2_X1    g15357(.A1(new_n16377_), .A2(new_n16310_), .ZN(new_n16378_));
  NAND2_X1   g15358(.A1(new_n16375_), .A2(new_n16376_), .ZN(new_n16379_));
  NAND2_X1   g15359(.A1(new_n16289_), .A2(new_n16294_), .ZN(new_n16380_));
  NOR2_X1    g15360(.A1(new_n16379_), .A2(new_n16380_), .ZN(new_n16381_));
  NAND4_X1   g15361(.A1(new_n16372_), .A2(new_n16374_), .A3(new_n16378_), .A4(new_n16381_), .ZN(new_n16382_));
  NOR2_X1    g15362(.A1(new_n16370_), .A2(new_n16382_), .ZN(new_n16383_));
  INV_X1     g15363(.I(new_n16383_), .ZN(new_n16384_));
  NAND2_X1   g15364(.A1(new_n16370_), .A2(new_n16382_), .ZN(new_n16385_));
  AOI21_X1   g15365(.A1(new_n16384_), .A2(new_n16385_), .B(new_n16318_), .ZN(new_n16386_));
  NAND2_X1   g15366(.A1(new_n16374_), .A2(new_n16372_), .ZN(new_n16387_));
  NAND2_X1   g15367(.A1(new_n16378_), .A2(new_n16381_), .ZN(new_n16388_));
  NOR2_X1    g15368(.A1(new_n16387_), .A2(new_n16388_), .ZN(new_n16389_));
  NAND2_X1   g15369(.A1(new_n16370_), .A2(new_n16389_), .ZN(new_n16390_));
  NAND2_X1   g15370(.A1(new_n16366_), .A2(new_n16369_), .ZN(new_n16391_));
  NAND3_X1   g15371(.A1(new_n16374_), .A2(new_n16372_), .A3(new_n16378_), .ZN(new_n16392_));
  NAND3_X1   g15372(.A1(new_n16310_), .A2(new_n16289_), .A3(new_n16294_), .ZN(new_n16393_));
  AOI21_X1   g15373(.A1(new_n16360_), .A2(new_n16329_), .B(new_n16393_), .ZN(new_n16394_));
  OAI21_X1   g15374(.A1(new_n16391_), .A2(new_n16392_), .B(new_n16394_), .ZN(new_n16395_));
  AND3_X2    g15375(.A1(new_n16395_), .A2(new_n16390_), .A3(new_n16317_), .Z(new_n16396_));
  NOR2_X1    g15376(.A1(new_n16386_), .A2(new_n16396_), .ZN(new_n16397_));
  INV_X1     g15377(.I(new_n16385_), .ZN(new_n16398_));
  OAI21_X1   g15378(.A1(new_n16398_), .A2(new_n16383_), .B(new_n16317_), .ZN(new_n16399_));
  NAND3_X1   g15379(.A1(new_n16395_), .A2(new_n16390_), .A3(new_n16317_), .ZN(new_n16400_));
  XOR2_X1    g15380(.A1(new_n16387_), .A2(new_n16388_), .Z(new_n16401_));
  INV_X1     g15381(.I(\A[519] ), .ZN(new_n16402_));
  NOR2_X1    g15382(.A1(new_n16402_), .A2(\A[518] ), .ZN(new_n16403_));
  INV_X1     g15383(.I(\A[518] ), .ZN(new_n16404_));
  NOR2_X1    g15384(.A1(new_n16404_), .A2(\A[519] ), .ZN(new_n16405_));
  OAI21_X1   g15385(.A1(new_n16403_), .A2(new_n16405_), .B(\A[517] ), .ZN(new_n16406_));
  INV_X1     g15386(.I(\A[517] ), .ZN(new_n16407_));
  NOR2_X1    g15387(.A1(\A[518] ), .A2(\A[519] ), .ZN(new_n16408_));
  NAND2_X1   g15388(.A1(\A[518] ), .A2(\A[519] ), .ZN(new_n16409_));
  INV_X1     g15389(.I(new_n16409_), .ZN(new_n16410_));
  OAI21_X1   g15390(.A1(new_n16410_), .A2(new_n16408_), .B(new_n16407_), .ZN(new_n16411_));
  NAND2_X1   g15391(.A1(new_n16406_), .A2(new_n16411_), .ZN(new_n16412_));
  INV_X1     g15392(.I(\A[522] ), .ZN(new_n16413_));
  NOR2_X1    g15393(.A1(new_n16413_), .A2(\A[521] ), .ZN(new_n16414_));
  INV_X1     g15394(.I(\A[521] ), .ZN(new_n16415_));
  NOR2_X1    g15395(.A1(new_n16415_), .A2(\A[522] ), .ZN(new_n16416_));
  OAI21_X1   g15396(.A1(new_n16414_), .A2(new_n16416_), .B(\A[520] ), .ZN(new_n16417_));
  INV_X1     g15397(.I(\A[520] ), .ZN(new_n16418_));
  NOR2_X1    g15398(.A1(\A[521] ), .A2(\A[522] ), .ZN(new_n16419_));
  NAND2_X1   g15399(.A1(\A[521] ), .A2(\A[522] ), .ZN(new_n16420_));
  INV_X1     g15400(.I(new_n16420_), .ZN(new_n16421_));
  OAI21_X1   g15401(.A1(new_n16421_), .A2(new_n16419_), .B(new_n16418_), .ZN(new_n16422_));
  NAND2_X1   g15402(.A1(new_n16417_), .A2(new_n16422_), .ZN(new_n16423_));
  NOR2_X1    g15403(.A1(new_n16412_), .A2(new_n16423_), .ZN(new_n16424_));
  AOI21_X1   g15404(.A1(new_n16418_), .A2(new_n16420_), .B(new_n16419_), .ZN(new_n16425_));
  INV_X1     g15405(.I(new_n16425_), .ZN(new_n16426_));
  AOI21_X1   g15406(.A1(new_n16407_), .A2(new_n16409_), .B(new_n16408_), .ZN(new_n16427_));
  INV_X1     g15407(.I(new_n16427_), .ZN(new_n16428_));
  NOR2_X1    g15408(.A1(new_n16426_), .A2(new_n16428_), .ZN(new_n16429_));
  NAND2_X1   g15409(.A1(new_n16424_), .A2(new_n16429_), .ZN(new_n16430_));
  NAND2_X1   g15410(.A1(new_n16404_), .A2(\A[519] ), .ZN(new_n16431_));
  NAND2_X1   g15411(.A1(new_n16402_), .A2(\A[518] ), .ZN(new_n16432_));
  AOI21_X1   g15412(.A1(new_n16431_), .A2(new_n16432_), .B(new_n16407_), .ZN(new_n16433_));
  INV_X1     g15413(.I(new_n16408_), .ZN(new_n16434_));
  AOI21_X1   g15414(.A1(new_n16434_), .A2(new_n16409_), .B(\A[517] ), .ZN(new_n16435_));
  NOR2_X1    g15415(.A1(new_n16435_), .A2(new_n16433_), .ZN(new_n16436_));
  NAND2_X1   g15416(.A1(new_n16415_), .A2(\A[522] ), .ZN(new_n16437_));
  NAND2_X1   g15417(.A1(new_n16413_), .A2(\A[521] ), .ZN(new_n16438_));
  AOI21_X1   g15418(.A1(new_n16437_), .A2(new_n16438_), .B(new_n16418_), .ZN(new_n16439_));
  INV_X1     g15419(.I(new_n16419_), .ZN(new_n16440_));
  AOI21_X1   g15420(.A1(new_n16440_), .A2(new_n16420_), .B(\A[520] ), .ZN(new_n16441_));
  NOR2_X1    g15421(.A1(new_n16441_), .A2(new_n16439_), .ZN(new_n16442_));
  NAND2_X1   g15422(.A1(new_n16436_), .A2(new_n16442_), .ZN(new_n16443_));
  NAND2_X1   g15423(.A1(new_n16412_), .A2(new_n16423_), .ZN(new_n16444_));
  NAND2_X1   g15424(.A1(new_n16443_), .A2(new_n16444_), .ZN(new_n16445_));
  INV_X1     g15425(.I(\A[511] ), .ZN(new_n16446_));
  INV_X1     g15426(.I(\A[512] ), .ZN(new_n16447_));
  NAND2_X1   g15427(.A1(new_n16447_), .A2(\A[513] ), .ZN(new_n16448_));
  INV_X1     g15428(.I(\A[513] ), .ZN(new_n16449_));
  NAND2_X1   g15429(.A1(new_n16449_), .A2(\A[512] ), .ZN(new_n16450_));
  AOI21_X1   g15430(.A1(new_n16448_), .A2(new_n16450_), .B(new_n16446_), .ZN(new_n16451_));
  NAND2_X1   g15431(.A1(new_n16447_), .A2(new_n16449_), .ZN(new_n16452_));
  NAND2_X1   g15432(.A1(\A[512] ), .A2(\A[513] ), .ZN(new_n16453_));
  AOI21_X1   g15433(.A1(new_n16452_), .A2(new_n16453_), .B(\A[511] ), .ZN(new_n16454_));
  NOR2_X1    g15434(.A1(new_n16454_), .A2(new_n16451_), .ZN(new_n16455_));
  INV_X1     g15435(.I(\A[514] ), .ZN(new_n16456_));
  INV_X1     g15436(.I(\A[515] ), .ZN(new_n16457_));
  NAND2_X1   g15437(.A1(new_n16457_), .A2(\A[516] ), .ZN(new_n16458_));
  INV_X1     g15438(.I(\A[516] ), .ZN(new_n16459_));
  NAND2_X1   g15439(.A1(new_n16459_), .A2(\A[515] ), .ZN(new_n16460_));
  AOI21_X1   g15440(.A1(new_n16458_), .A2(new_n16460_), .B(new_n16456_), .ZN(new_n16461_));
  NAND2_X1   g15441(.A1(new_n16457_), .A2(new_n16459_), .ZN(new_n16462_));
  NAND2_X1   g15442(.A1(\A[515] ), .A2(\A[516] ), .ZN(new_n16463_));
  AOI21_X1   g15443(.A1(new_n16462_), .A2(new_n16463_), .B(\A[514] ), .ZN(new_n16464_));
  NOR2_X1    g15444(.A1(new_n16464_), .A2(new_n16461_), .ZN(new_n16465_));
  NAND2_X1   g15445(.A1(new_n16463_), .A2(new_n16456_), .ZN(new_n16466_));
  NAND2_X1   g15446(.A1(new_n16466_), .A2(new_n16462_), .ZN(new_n16467_));
  NAND2_X1   g15447(.A1(new_n16453_), .A2(new_n16446_), .ZN(new_n16468_));
  NAND2_X1   g15448(.A1(new_n16468_), .A2(new_n16452_), .ZN(new_n16469_));
  NOR2_X1    g15449(.A1(new_n16467_), .A2(new_n16469_), .ZN(new_n16470_));
  NOR2_X1    g15450(.A1(new_n16445_), .A2(new_n16430_), .ZN(new_n16471_));
  NOR2_X1    g15451(.A1(new_n16401_), .A2(new_n16471_), .ZN(new_n16472_));
  AOI21_X1   g15452(.A1(new_n16399_), .A2(new_n16400_), .B(new_n16472_), .ZN(new_n16473_));
  INV_X1     g15453(.I(new_n16472_), .ZN(new_n16474_));
  NOR3_X1    g15454(.A1(new_n16386_), .A2(new_n16474_), .A3(new_n16396_), .ZN(new_n16475_));
  NOR2_X1    g15455(.A1(new_n16424_), .A2(new_n16428_), .ZN(new_n16476_));
  NOR2_X1    g15456(.A1(new_n16443_), .A2(new_n16427_), .ZN(new_n16477_));
  OAI21_X1   g15457(.A1(new_n16476_), .A2(new_n16477_), .B(new_n16425_), .ZN(new_n16478_));
  NAND2_X1   g15458(.A1(new_n16443_), .A2(new_n16427_), .ZN(new_n16479_));
  NAND2_X1   g15459(.A1(new_n16424_), .A2(new_n16428_), .ZN(new_n16480_));
  NAND3_X1   g15460(.A1(new_n16480_), .A2(new_n16479_), .A3(new_n16426_), .ZN(new_n16481_));
  AND2_X2    g15461(.A1(new_n16478_), .A2(new_n16481_), .Z(new_n16482_));
  NOR4_X1    g15462(.A1(new_n16451_), .A2(new_n16454_), .A3(new_n16464_), .A4(new_n16461_), .ZN(new_n16483_));
  NOR2_X1    g15463(.A1(new_n16455_), .A2(new_n16465_), .ZN(new_n16484_));
  NOR4_X1    g15464(.A1(new_n16445_), .A2(new_n16430_), .A3(new_n16483_), .A4(new_n16484_), .ZN(new_n16485_));
  NAND2_X1   g15465(.A1(new_n16455_), .A2(new_n16465_), .ZN(new_n16486_));
  INV_X1     g15466(.I(new_n16470_), .ZN(new_n16487_));
  NOR2_X1    g15467(.A1(new_n16486_), .A2(new_n16487_), .ZN(new_n16488_));
  NOR2_X1    g15468(.A1(new_n16442_), .A2(new_n16412_), .ZN(new_n16489_));
  NOR2_X1    g15469(.A1(new_n16436_), .A2(new_n16423_), .ZN(new_n16490_));
  OAI21_X1   g15470(.A1(new_n16489_), .A2(new_n16490_), .B(new_n16429_), .ZN(new_n16491_));
  NAND2_X1   g15471(.A1(new_n16491_), .A2(new_n16488_), .ZN(new_n16492_));
  AOI21_X1   g15472(.A1(new_n16482_), .A2(new_n16485_), .B(new_n16492_), .ZN(new_n16493_));
  INV_X1     g15473(.I(new_n16469_), .ZN(new_n16494_));
  NAND2_X1   g15474(.A1(new_n16486_), .A2(new_n16494_), .ZN(new_n16495_));
  NAND2_X1   g15475(.A1(new_n16483_), .A2(new_n16469_), .ZN(new_n16496_));
  AOI21_X1   g15476(.A1(new_n16495_), .A2(new_n16496_), .B(new_n16467_), .ZN(new_n16497_));
  INV_X1     g15477(.I(new_n16467_), .ZN(new_n16498_));
  NOR2_X1    g15478(.A1(new_n16483_), .A2(new_n16469_), .ZN(new_n16499_));
  NOR2_X1    g15479(.A1(new_n16486_), .A2(new_n16494_), .ZN(new_n16500_));
  NOR3_X1    g15480(.A1(new_n16500_), .A2(new_n16498_), .A3(new_n16499_), .ZN(new_n16501_));
  OR2_X2     g15481(.A1(new_n16501_), .A2(new_n16497_), .Z(new_n16502_));
  NOR2_X1    g15482(.A1(new_n16445_), .A2(new_n16430_), .ZN(new_n16503_));
  NOR2_X1    g15483(.A1(new_n16484_), .A2(new_n16483_), .ZN(new_n16504_));
  NAND3_X1   g15484(.A1(new_n16503_), .A2(new_n16488_), .A3(new_n16504_), .ZN(new_n16505_));
  NAND2_X1   g15485(.A1(new_n16502_), .A2(new_n16505_), .ZN(new_n16506_));
  NAND3_X1   g15486(.A1(new_n16478_), .A2(new_n16481_), .A3(new_n16491_), .ZN(new_n16507_));
  OAI21_X1   g15487(.A1(new_n16502_), .A2(new_n16505_), .B(new_n16507_), .ZN(new_n16508_));
  NOR2_X1    g15488(.A1(new_n16501_), .A2(new_n16497_), .ZN(new_n16509_));
  INV_X1     g15489(.I(new_n16505_), .ZN(new_n16510_));
  AND3_X2    g15490(.A1(new_n16478_), .A2(new_n16481_), .A3(new_n16491_), .Z(new_n16511_));
  NAND3_X1   g15491(.A1(new_n16511_), .A2(new_n16510_), .A3(new_n16509_), .ZN(new_n16512_));
  NAND2_X1   g15492(.A1(new_n16512_), .A2(new_n16508_), .ZN(new_n16513_));
  AOI22_X1   g15493(.A1(new_n16513_), .A2(new_n16506_), .B1(new_n16493_), .B2(new_n16502_), .ZN(new_n16514_));
  OAI22_X1   g15494(.A1(new_n16475_), .A2(new_n16473_), .B1(new_n16514_), .B2(new_n16397_), .ZN(new_n16515_));
  NAND2_X1   g15495(.A1(new_n16390_), .A2(new_n16318_), .ZN(new_n16516_));
  NOR2_X1    g15496(.A1(new_n16322_), .A2(new_n16327_), .ZN(new_n16517_));
  OAI21_X1   g15497(.A1(new_n16364_), .A2(new_n16517_), .B(new_n16371_), .ZN(new_n16518_));
  NOR2_X1    g15498(.A1(new_n16289_), .A2(new_n16294_), .ZN(new_n16519_));
  OAI21_X1   g15499(.A1(new_n16379_), .A2(new_n16519_), .B(new_n16380_), .ZN(new_n16520_));
  XNOR2_X1   g15500(.A1(new_n16518_), .A2(new_n16520_), .ZN(new_n16521_));
  NAND3_X1   g15501(.A1(new_n16516_), .A2(new_n16395_), .A3(new_n16521_), .ZN(new_n16522_));
  AOI21_X1   g15502(.A1(new_n16510_), .A2(new_n16507_), .B(new_n16509_), .ZN(new_n16523_));
  OAI21_X1   g15503(.A1(new_n16425_), .A2(new_n16427_), .B(new_n16424_), .ZN(new_n16524_));
  OAI21_X1   g15504(.A1(new_n16426_), .A2(new_n16428_), .B(new_n16524_), .ZN(new_n16525_));
  NOR2_X1    g15505(.A1(new_n16498_), .A2(new_n16494_), .ZN(new_n16526_));
  OAI21_X1   g15506(.A1(new_n16486_), .A2(new_n16526_), .B(new_n16487_), .ZN(new_n16527_));
  XOR2_X1    g15507(.A1(new_n16525_), .A2(new_n16527_), .Z(new_n16528_));
  NOR3_X1    g15508(.A1(new_n16523_), .A2(new_n16528_), .A3(new_n16493_), .ZN(new_n16529_));
  INV_X1     g15509(.I(new_n16529_), .ZN(new_n16530_));
  NAND2_X1   g15510(.A1(new_n16530_), .A2(new_n16522_), .ZN(new_n16531_));
  NAND2_X1   g15511(.A1(new_n16515_), .A2(new_n16531_), .ZN(new_n16532_));
  NOR2_X1    g15512(.A1(new_n16530_), .A2(new_n16522_), .ZN(new_n16533_));
  NAND2_X1   g15513(.A1(new_n16525_), .A2(new_n16527_), .ZN(new_n16534_));
  NOR2_X1    g15514(.A1(new_n16523_), .A2(new_n16493_), .ZN(new_n16535_));
  OAI21_X1   g15515(.A1(new_n16525_), .A2(new_n16527_), .B(new_n16535_), .ZN(new_n16536_));
  NAND2_X1   g15516(.A1(new_n16536_), .A2(new_n16534_), .ZN(new_n16537_));
  INV_X1     g15517(.I(new_n16537_), .ZN(new_n16538_));
  NAND2_X1   g15518(.A1(new_n16518_), .A2(new_n16520_), .ZN(new_n16539_));
  OR2_X2     g15519(.A1(new_n16518_), .A2(new_n16520_), .Z(new_n16540_));
  NAND3_X1   g15520(.A1(new_n16516_), .A2(new_n16395_), .A3(new_n16540_), .ZN(new_n16541_));
  NAND2_X1   g15521(.A1(new_n16541_), .A2(new_n16539_), .ZN(new_n16542_));
  INV_X1     g15522(.I(new_n16542_), .ZN(new_n16543_));
  AOI22_X1   g15523(.A1(new_n16532_), .A2(new_n16533_), .B1(new_n16543_), .B2(new_n16538_), .ZN(new_n16544_));
  NAND2_X1   g15524(.A1(new_n16537_), .A2(new_n16542_), .ZN(new_n16545_));
  INV_X1     g15525(.I(new_n16545_), .ZN(new_n16546_));
  NOR2_X1    g15526(.A1(new_n16544_), .A2(new_n16546_), .ZN(new_n16547_));
  INV_X1     g15527(.I(new_n16547_), .ZN(new_n16548_));
  NAND2_X1   g15528(.A1(new_n16285_), .A2(new_n16548_), .ZN(new_n16549_));
  XOR2_X1    g15529(.A1(new_n16529_), .A2(new_n16522_), .Z(new_n16550_));
  NOR2_X1    g15530(.A1(new_n16515_), .A2(new_n16550_), .ZN(new_n16551_));
  NAND2_X1   g15531(.A1(new_n16399_), .A2(new_n16400_), .ZN(new_n16552_));
  OAI21_X1   g15532(.A1(new_n16396_), .A2(new_n16386_), .B(new_n16474_), .ZN(new_n16553_));
  NAND3_X1   g15533(.A1(new_n16399_), .A2(new_n16400_), .A3(new_n16472_), .ZN(new_n16554_));
  NAND2_X1   g15534(.A1(new_n16493_), .A2(new_n16502_), .ZN(new_n16555_));
  AOI21_X1   g15535(.A1(new_n16509_), .A2(new_n16510_), .B(new_n16511_), .ZN(new_n16556_));
  NOR3_X1    g15536(.A1(new_n16502_), .A2(new_n16505_), .A3(new_n16507_), .ZN(new_n16557_));
  OAI21_X1   g15537(.A1(new_n16556_), .A2(new_n16557_), .B(new_n16506_), .ZN(new_n16558_));
  NAND2_X1   g15538(.A1(new_n16558_), .A2(new_n16555_), .ZN(new_n16559_));
  AOI22_X1   g15539(.A1(new_n16553_), .A2(new_n16554_), .B1(new_n16559_), .B2(new_n16552_), .ZN(new_n16560_));
  XNOR2_X1   g15540(.A1(new_n16529_), .A2(new_n16522_), .ZN(new_n16561_));
  NOR2_X1    g15541(.A1(new_n16560_), .A2(new_n16561_), .ZN(new_n16562_));
  AND2_X2    g15542(.A1(new_n16125_), .A2(new_n16131_), .Z(new_n16563_));
  AOI21_X1   g15543(.A1(new_n16125_), .A2(new_n16131_), .B(new_n16212_), .ZN(new_n16564_));
  INV_X1     g15544(.I(new_n16213_), .ZN(new_n16565_));
  OAI21_X1   g15545(.A1(new_n16239_), .A2(new_n16242_), .B(new_n16249_), .ZN(new_n16566_));
  NAND2_X1   g15546(.A1(new_n16247_), .A2(new_n16246_), .ZN(new_n16567_));
  NAND2_X1   g15547(.A1(new_n16567_), .A2(new_n16566_), .ZN(new_n16568_));
  AOI22_X1   g15548(.A1(new_n16568_), .A2(new_n16243_), .B1(new_n16230_), .B2(new_n16239_), .ZN(new_n16569_));
  OAI22_X1   g15549(.A1(new_n16565_), .A2(new_n16564_), .B1(new_n16569_), .B2(new_n16563_), .ZN(new_n16570_));
  XNOR2_X1   g15550(.A1(new_n16261_), .A2(new_n16269_), .ZN(new_n16571_));
  NOR2_X1    g15551(.A1(new_n16570_), .A2(new_n16571_), .ZN(new_n16572_));
  NOR2_X1    g15552(.A1(new_n16261_), .A2(new_n16269_), .ZN(new_n16573_));
  AND2_X2    g15553(.A1(new_n16261_), .A2(new_n16269_), .Z(new_n16574_));
  NOR2_X1    g15554(.A1(new_n16574_), .A2(new_n16573_), .ZN(new_n16575_));
  NOR2_X1    g15555(.A1(new_n16253_), .A2(new_n16575_), .ZN(new_n16576_));
  NOR4_X1    g15556(.A1(new_n16551_), .A2(new_n16562_), .A3(new_n16572_), .A4(new_n16576_), .ZN(new_n16577_));
  NOR3_X1    g15557(.A1(new_n16565_), .A2(new_n16564_), .A3(new_n16252_), .ZN(new_n16578_));
  INV_X1     g15558(.I(new_n16578_), .ZN(new_n16579_));
  NOR2_X1    g15559(.A1(new_n16133_), .A2(new_n16177_), .ZN(new_n16580_));
  NOR2_X1    g15560(.A1(new_n16580_), .A2(new_n16212_), .ZN(new_n16581_));
  XOR2_X1    g15561(.A1(new_n16401_), .A2(new_n16471_), .Z(new_n16582_));
  NAND2_X1   g15562(.A1(new_n16582_), .A2(new_n16581_), .ZN(new_n16583_));
  INV_X1     g15563(.I(new_n16583_), .ZN(new_n16584_));
  NOR2_X1    g15564(.A1(new_n16578_), .A2(new_n16584_), .ZN(new_n16585_));
  INV_X1     g15565(.I(new_n16585_), .ZN(new_n16586_));
  NAND2_X1   g15566(.A1(new_n16578_), .A2(new_n16584_), .ZN(new_n16587_));
  OAI21_X1   g15567(.A1(new_n16475_), .A2(new_n16473_), .B(new_n16514_), .ZN(new_n16588_));
  NAND3_X1   g15568(.A1(new_n16553_), .A2(new_n16559_), .A3(new_n16554_), .ZN(new_n16589_));
  NAND2_X1   g15569(.A1(new_n16588_), .A2(new_n16589_), .ZN(new_n16590_));
  AOI22_X1   g15570(.A1(new_n16586_), .A2(new_n16587_), .B1(new_n16579_), .B2(new_n16590_), .ZN(new_n16591_));
  OAI22_X1   g15571(.A1(new_n16551_), .A2(new_n16562_), .B1(new_n16572_), .B2(new_n16576_), .ZN(new_n16592_));
  AOI21_X1   g15572(.A1(new_n16591_), .A2(new_n16592_), .B(new_n16577_), .ZN(new_n16593_));
  AOI21_X1   g15573(.A1(new_n16532_), .A2(new_n16533_), .B(new_n16538_), .ZN(new_n16594_));
  INV_X1     g15574(.I(new_n16522_), .ZN(new_n16595_));
  NAND3_X1   g15575(.A1(new_n16560_), .A2(new_n16595_), .A3(new_n16529_), .ZN(new_n16596_));
  NOR2_X1    g15576(.A1(new_n16596_), .A2(new_n16537_), .ZN(new_n16597_));
  OAI21_X1   g15577(.A1(new_n16597_), .A2(new_n16594_), .B(new_n16542_), .ZN(new_n16598_));
  NAND2_X1   g15578(.A1(new_n16596_), .A2(new_n16537_), .ZN(new_n16599_));
  NAND3_X1   g15579(.A1(new_n16532_), .A2(new_n16533_), .A3(new_n16538_), .ZN(new_n16600_));
  NAND3_X1   g15580(.A1(new_n16599_), .A2(new_n16600_), .A3(new_n16543_), .ZN(new_n16601_));
  NAND2_X1   g15581(.A1(new_n16598_), .A2(new_n16601_), .ZN(new_n16602_));
  INV_X1     g15582(.I(new_n16573_), .ZN(new_n16603_));
  NAND2_X1   g15583(.A1(new_n16570_), .A2(new_n16603_), .ZN(new_n16604_));
  AOI21_X1   g15584(.A1(new_n16604_), .A2(new_n16574_), .B(new_n16281_), .ZN(new_n16605_));
  NOR2_X1    g15585(.A1(new_n16270_), .A2(new_n16274_), .ZN(new_n16606_));
  OAI21_X1   g15586(.A1(new_n16605_), .A2(new_n16606_), .B(new_n16278_), .ZN(new_n16607_));
  NAND2_X1   g15587(.A1(new_n16270_), .A2(new_n16274_), .ZN(new_n16608_));
  NAND4_X1   g15588(.A1(new_n16253_), .A2(new_n16281_), .A3(new_n16261_), .A4(new_n16269_), .ZN(new_n16609_));
  NAND3_X1   g15589(.A1(new_n16608_), .A2(new_n16282_), .A3(new_n16609_), .ZN(new_n16610_));
  NAND2_X1   g15590(.A1(new_n16607_), .A2(new_n16610_), .ZN(new_n16611_));
  OAI21_X1   g15591(.A1(new_n16602_), .A2(new_n16611_), .B(new_n16593_), .ZN(new_n16612_));
  XOR2_X1    g15592(.A1(new_n16278_), .A2(new_n16274_), .Z(new_n16613_));
  XOR2_X1    g15593(.A1(new_n16537_), .A2(new_n16542_), .Z(new_n16614_));
  NOR4_X1    g15594(.A1(new_n16614_), .A2(new_n16613_), .A3(new_n16270_), .A4(new_n16596_), .ZN(new_n16615_));
  NAND2_X1   g15595(.A1(new_n16612_), .A2(new_n16615_), .ZN(new_n16616_));
  NOR4_X1    g15596(.A1(new_n16280_), .A2(new_n16283_), .A3(new_n16544_), .A4(new_n16546_), .ZN(new_n16617_));
  NAND2_X1   g15597(.A1(new_n16616_), .A2(new_n16617_), .ZN(new_n16618_));
  NAND2_X1   g15598(.A1(new_n16618_), .A2(new_n16549_), .ZN(new_n16619_));
  INV_X1     g15599(.I(\A[502] ), .ZN(new_n16620_));
  NOR2_X1    g15600(.A1(\A[503] ), .A2(\A[504] ), .ZN(new_n16621_));
  NAND2_X1   g15601(.A1(\A[503] ), .A2(\A[504] ), .ZN(new_n16622_));
  AOI21_X1   g15602(.A1(new_n16620_), .A2(new_n16622_), .B(new_n16621_), .ZN(new_n16623_));
  INV_X1     g15603(.I(new_n16623_), .ZN(new_n16624_));
  INV_X1     g15604(.I(\A[499] ), .ZN(new_n16625_));
  NOR2_X1    g15605(.A1(\A[500] ), .A2(\A[501] ), .ZN(new_n16626_));
  NAND2_X1   g15606(.A1(\A[500] ), .A2(\A[501] ), .ZN(new_n16627_));
  AOI21_X1   g15607(.A1(new_n16625_), .A2(new_n16627_), .B(new_n16626_), .ZN(new_n16628_));
  INV_X1     g15608(.I(\A[500] ), .ZN(new_n16629_));
  NAND2_X1   g15609(.A1(new_n16629_), .A2(\A[501] ), .ZN(new_n16630_));
  INV_X1     g15610(.I(\A[501] ), .ZN(new_n16631_));
  NAND2_X1   g15611(.A1(new_n16631_), .A2(\A[500] ), .ZN(new_n16632_));
  AOI21_X1   g15612(.A1(new_n16630_), .A2(new_n16632_), .B(new_n16625_), .ZN(new_n16633_));
  INV_X1     g15613(.I(new_n16626_), .ZN(new_n16634_));
  AOI21_X1   g15614(.A1(new_n16634_), .A2(new_n16627_), .B(\A[499] ), .ZN(new_n16635_));
  INV_X1     g15615(.I(\A[503] ), .ZN(new_n16636_));
  NAND2_X1   g15616(.A1(new_n16636_), .A2(\A[504] ), .ZN(new_n16637_));
  INV_X1     g15617(.I(\A[504] ), .ZN(new_n16638_));
  NAND2_X1   g15618(.A1(new_n16638_), .A2(\A[503] ), .ZN(new_n16639_));
  AOI21_X1   g15619(.A1(new_n16637_), .A2(new_n16639_), .B(new_n16620_), .ZN(new_n16640_));
  INV_X1     g15620(.I(new_n16621_), .ZN(new_n16641_));
  AOI21_X1   g15621(.A1(new_n16641_), .A2(new_n16622_), .B(\A[502] ), .ZN(new_n16642_));
  NOR4_X1    g15622(.A1(new_n16633_), .A2(new_n16635_), .A3(new_n16642_), .A4(new_n16640_), .ZN(new_n16643_));
  INV_X1     g15623(.I(new_n16643_), .ZN(new_n16644_));
  NAND2_X1   g15624(.A1(new_n16644_), .A2(new_n16628_), .ZN(new_n16645_));
  INV_X1     g15625(.I(new_n16628_), .ZN(new_n16646_));
  NAND2_X1   g15626(.A1(new_n16643_), .A2(new_n16646_), .ZN(new_n16647_));
  AOI21_X1   g15627(.A1(new_n16645_), .A2(new_n16647_), .B(new_n16624_), .ZN(new_n16648_));
  AND3_X2    g15628(.A1(new_n16645_), .A2(new_n16624_), .A3(new_n16647_), .Z(new_n16649_));
  NOR2_X1    g15629(.A1(new_n16649_), .A2(new_n16648_), .ZN(new_n16650_));
  INV_X1     g15630(.I(\A[508] ), .ZN(new_n16651_));
  NOR2_X1    g15631(.A1(\A[509] ), .A2(\A[510] ), .ZN(new_n16652_));
  NAND2_X1   g15632(.A1(\A[509] ), .A2(\A[510] ), .ZN(new_n16653_));
  AOI21_X1   g15633(.A1(new_n16651_), .A2(new_n16653_), .B(new_n16652_), .ZN(new_n16654_));
  INV_X1     g15634(.I(new_n16654_), .ZN(new_n16655_));
  INV_X1     g15635(.I(\A[505] ), .ZN(new_n16656_));
  NOR2_X1    g15636(.A1(\A[506] ), .A2(\A[507] ), .ZN(new_n16657_));
  NAND2_X1   g15637(.A1(\A[506] ), .A2(\A[507] ), .ZN(new_n16658_));
  AOI21_X1   g15638(.A1(new_n16656_), .A2(new_n16658_), .B(new_n16657_), .ZN(new_n16659_));
  INV_X1     g15639(.I(new_n16659_), .ZN(new_n16660_));
  NOR2_X1    g15640(.A1(new_n16655_), .A2(new_n16660_), .ZN(new_n16661_));
  INV_X1     g15641(.I(new_n16661_), .ZN(new_n16662_));
  INV_X1     g15642(.I(\A[506] ), .ZN(new_n16663_));
  NAND2_X1   g15643(.A1(new_n16663_), .A2(\A[507] ), .ZN(new_n16664_));
  INV_X1     g15644(.I(\A[507] ), .ZN(new_n16665_));
  NAND2_X1   g15645(.A1(new_n16665_), .A2(\A[506] ), .ZN(new_n16666_));
  AOI21_X1   g15646(.A1(new_n16664_), .A2(new_n16666_), .B(new_n16656_), .ZN(new_n16667_));
  INV_X1     g15647(.I(new_n16657_), .ZN(new_n16668_));
  AOI21_X1   g15648(.A1(new_n16668_), .A2(new_n16658_), .B(\A[505] ), .ZN(new_n16669_));
  NOR2_X1    g15649(.A1(new_n16669_), .A2(new_n16667_), .ZN(new_n16670_));
  INV_X1     g15650(.I(\A[510] ), .ZN(new_n16671_));
  NOR2_X1    g15651(.A1(new_n16671_), .A2(\A[509] ), .ZN(new_n16672_));
  INV_X1     g15652(.I(\A[509] ), .ZN(new_n16673_));
  NOR2_X1    g15653(.A1(new_n16673_), .A2(\A[510] ), .ZN(new_n16674_));
  OAI21_X1   g15654(.A1(new_n16672_), .A2(new_n16674_), .B(\A[508] ), .ZN(new_n16675_));
  INV_X1     g15655(.I(new_n16653_), .ZN(new_n16676_));
  OAI21_X1   g15656(.A1(new_n16676_), .A2(new_n16652_), .B(new_n16651_), .ZN(new_n16677_));
  NAND2_X1   g15657(.A1(new_n16675_), .A2(new_n16677_), .ZN(new_n16678_));
  NAND2_X1   g15658(.A1(new_n16670_), .A2(new_n16678_), .ZN(new_n16679_));
  NOR2_X1    g15659(.A1(new_n16665_), .A2(\A[506] ), .ZN(new_n16680_));
  NOR2_X1    g15660(.A1(new_n16663_), .A2(\A[507] ), .ZN(new_n16681_));
  OAI21_X1   g15661(.A1(new_n16680_), .A2(new_n16681_), .B(\A[505] ), .ZN(new_n16682_));
  INV_X1     g15662(.I(new_n16658_), .ZN(new_n16683_));
  OAI21_X1   g15663(.A1(new_n16683_), .A2(new_n16657_), .B(new_n16656_), .ZN(new_n16684_));
  NAND2_X1   g15664(.A1(new_n16682_), .A2(new_n16684_), .ZN(new_n16685_));
  NAND2_X1   g15665(.A1(new_n16673_), .A2(\A[510] ), .ZN(new_n16686_));
  NAND2_X1   g15666(.A1(new_n16671_), .A2(\A[509] ), .ZN(new_n16687_));
  AOI21_X1   g15667(.A1(new_n16686_), .A2(new_n16687_), .B(new_n16651_), .ZN(new_n16688_));
  INV_X1     g15668(.I(new_n16652_), .ZN(new_n16689_));
  AOI21_X1   g15669(.A1(new_n16689_), .A2(new_n16653_), .B(\A[508] ), .ZN(new_n16690_));
  NOR2_X1    g15670(.A1(new_n16690_), .A2(new_n16688_), .ZN(new_n16691_));
  NAND2_X1   g15671(.A1(new_n16691_), .A2(new_n16685_), .ZN(new_n16692_));
  AOI21_X1   g15672(.A1(new_n16679_), .A2(new_n16692_), .B(new_n16662_), .ZN(new_n16693_));
  INV_X1     g15673(.I(new_n16693_), .ZN(new_n16694_));
  NOR2_X1    g15674(.A1(new_n16685_), .A2(new_n16678_), .ZN(new_n16695_));
  NOR2_X1    g15675(.A1(new_n16695_), .A2(new_n16660_), .ZN(new_n16696_));
  NAND2_X1   g15676(.A1(new_n16670_), .A2(new_n16691_), .ZN(new_n16697_));
  NOR2_X1    g15677(.A1(new_n16697_), .A2(new_n16659_), .ZN(new_n16698_));
  OAI21_X1   g15678(.A1(new_n16696_), .A2(new_n16698_), .B(new_n16654_), .ZN(new_n16699_));
  NAND2_X1   g15679(.A1(new_n16697_), .A2(new_n16659_), .ZN(new_n16700_));
  NAND2_X1   g15680(.A1(new_n16695_), .A2(new_n16660_), .ZN(new_n16701_));
  NAND3_X1   g15681(.A1(new_n16701_), .A2(new_n16700_), .A3(new_n16655_), .ZN(new_n16702_));
  NAND3_X1   g15682(.A1(new_n16699_), .A2(new_n16702_), .A3(new_n16694_), .ZN(new_n16703_));
  NOR2_X1    g15683(.A1(new_n16697_), .A2(new_n16662_), .ZN(new_n16704_));
  NOR2_X1    g15684(.A1(new_n16670_), .A2(new_n16691_), .ZN(new_n16705_));
  NOR2_X1    g15685(.A1(new_n16705_), .A2(new_n16695_), .ZN(new_n16706_));
  NOR2_X1    g15686(.A1(new_n16635_), .A2(new_n16633_), .ZN(new_n16707_));
  NOR2_X1    g15687(.A1(new_n16642_), .A2(new_n16640_), .ZN(new_n16708_));
  NOR2_X1    g15688(.A1(new_n16707_), .A2(new_n16708_), .ZN(new_n16709_));
  NOR2_X1    g15689(.A1(new_n16709_), .A2(new_n16643_), .ZN(new_n16710_));
  NAND2_X1   g15690(.A1(new_n16623_), .A2(new_n16628_), .ZN(new_n16711_));
  NOR2_X1    g15691(.A1(new_n16644_), .A2(new_n16711_), .ZN(new_n16712_));
  NAND4_X1   g15692(.A1(new_n16706_), .A2(new_n16712_), .A3(new_n16704_), .A4(new_n16710_), .ZN(new_n16713_));
  NOR2_X1    g15693(.A1(new_n16703_), .A2(new_n16713_), .ZN(new_n16714_));
  AOI21_X1   g15694(.A1(new_n16701_), .A2(new_n16700_), .B(new_n16655_), .ZN(new_n16715_));
  NOR3_X1    g15695(.A1(new_n16696_), .A2(new_n16698_), .A3(new_n16654_), .ZN(new_n16716_));
  NOR3_X1    g15696(.A1(new_n16715_), .A2(new_n16716_), .A3(new_n16693_), .ZN(new_n16717_));
  INV_X1     g15697(.I(new_n16713_), .ZN(new_n16718_));
  NOR2_X1    g15698(.A1(new_n16717_), .A2(new_n16718_), .ZN(new_n16719_));
  OAI21_X1   g15699(.A1(new_n16719_), .A2(new_n16714_), .B(new_n16650_), .ZN(new_n16720_));
  NAND2_X1   g15700(.A1(new_n16703_), .A2(new_n16718_), .ZN(new_n16721_));
  NAND2_X1   g15701(.A1(new_n16699_), .A2(new_n16702_), .ZN(new_n16722_));
  NAND3_X1   g15702(.A1(new_n16706_), .A2(new_n16704_), .A3(new_n16710_), .ZN(new_n16723_));
  NOR3_X1    g15703(.A1(new_n16693_), .A2(new_n16644_), .A3(new_n16711_), .ZN(new_n16724_));
  OAI21_X1   g15704(.A1(new_n16722_), .A2(new_n16723_), .B(new_n16724_), .ZN(new_n16725_));
  NAND3_X1   g15705(.A1(new_n16721_), .A2(new_n16725_), .A3(new_n16650_), .ZN(new_n16726_));
  NAND2_X1   g15706(.A1(new_n16720_), .A2(new_n16726_), .ZN(new_n16727_));
  NAND2_X1   g15707(.A1(new_n16706_), .A2(new_n16704_), .ZN(new_n16728_));
  NAND2_X1   g15708(.A1(new_n16712_), .A2(new_n16710_), .ZN(new_n16729_));
  XOR2_X1    g15709(.A1(new_n16728_), .A2(new_n16729_), .Z(new_n16730_));
  INV_X1     g15710(.I(\A[495] ), .ZN(new_n16731_));
  NOR2_X1    g15711(.A1(new_n16731_), .A2(\A[494] ), .ZN(new_n16732_));
  INV_X1     g15712(.I(\A[494] ), .ZN(new_n16733_));
  NOR2_X1    g15713(.A1(new_n16733_), .A2(\A[495] ), .ZN(new_n16734_));
  OAI21_X1   g15714(.A1(new_n16732_), .A2(new_n16734_), .B(\A[493] ), .ZN(new_n16735_));
  INV_X1     g15715(.I(\A[493] ), .ZN(new_n16736_));
  NOR2_X1    g15716(.A1(\A[494] ), .A2(\A[495] ), .ZN(new_n16737_));
  NOR2_X1    g15717(.A1(new_n16733_), .A2(new_n16731_), .ZN(new_n16738_));
  OAI21_X1   g15718(.A1(new_n16738_), .A2(new_n16737_), .B(new_n16736_), .ZN(new_n16739_));
  INV_X1     g15719(.I(\A[498] ), .ZN(new_n16740_));
  NOR2_X1    g15720(.A1(new_n16740_), .A2(\A[497] ), .ZN(new_n16741_));
  INV_X1     g15721(.I(\A[497] ), .ZN(new_n16742_));
  NOR2_X1    g15722(.A1(new_n16742_), .A2(\A[498] ), .ZN(new_n16743_));
  OAI21_X1   g15723(.A1(new_n16741_), .A2(new_n16743_), .B(\A[496] ), .ZN(new_n16744_));
  INV_X1     g15724(.I(\A[496] ), .ZN(new_n16745_));
  NOR2_X1    g15725(.A1(\A[497] ), .A2(\A[498] ), .ZN(new_n16746_));
  NOR2_X1    g15726(.A1(new_n16742_), .A2(new_n16740_), .ZN(new_n16747_));
  OAI21_X1   g15727(.A1(new_n16747_), .A2(new_n16746_), .B(new_n16745_), .ZN(new_n16748_));
  NAND4_X1   g15728(.A1(new_n16735_), .A2(new_n16739_), .A3(new_n16748_), .A4(new_n16744_), .ZN(new_n16749_));
  INV_X1     g15729(.I(new_n16749_), .ZN(new_n16750_));
  INV_X1     g15730(.I(new_n16746_), .ZN(new_n16751_));
  OAI21_X1   g15731(.A1(\A[496] ), .A2(new_n16747_), .B(new_n16751_), .ZN(new_n16752_));
  INV_X1     g15732(.I(new_n16737_), .ZN(new_n16753_));
  OAI21_X1   g15733(.A1(\A[493] ), .A2(new_n16738_), .B(new_n16753_), .ZN(new_n16754_));
  NOR2_X1    g15734(.A1(new_n16752_), .A2(new_n16754_), .ZN(new_n16755_));
  NAND2_X1   g15735(.A1(new_n16750_), .A2(new_n16755_), .ZN(new_n16756_));
  NAND2_X1   g15736(.A1(new_n16739_), .A2(new_n16735_), .ZN(new_n16757_));
  NAND2_X1   g15737(.A1(new_n16748_), .A2(new_n16744_), .ZN(new_n16758_));
  NAND2_X1   g15738(.A1(new_n16757_), .A2(new_n16758_), .ZN(new_n16759_));
  NAND2_X1   g15739(.A1(new_n16759_), .A2(new_n16749_), .ZN(new_n16760_));
  INV_X1     g15740(.I(\A[487] ), .ZN(new_n16761_));
  INV_X1     g15741(.I(\A[488] ), .ZN(new_n16762_));
  NAND2_X1   g15742(.A1(new_n16762_), .A2(\A[489] ), .ZN(new_n16763_));
  INV_X1     g15743(.I(\A[489] ), .ZN(new_n16764_));
  NAND2_X1   g15744(.A1(new_n16764_), .A2(\A[488] ), .ZN(new_n16765_));
  AOI21_X1   g15745(.A1(new_n16763_), .A2(new_n16765_), .B(new_n16761_), .ZN(new_n16766_));
  NAND2_X1   g15746(.A1(new_n16762_), .A2(new_n16764_), .ZN(new_n16767_));
  NAND2_X1   g15747(.A1(\A[488] ), .A2(\A[489] ), .ZN(new_n16768_));
  AOI21_X1   g15748(.A1(new_n16767_), .A2(new_n16768_), .B(\A[487] ), .ZN(new_n16769_));
  NOR2_X1    g15749(.A1(new_n16769_), .A2(new_n16766_), .ZN(new_n16770_));
  INV_X1     g15750(.I(\A[490] ), .ZN(new_n16771_));
  INV_X1     g15751(.I(\A[491] ), .ZN(new_n16772_));
  NAND2_X1   g15752(.A1(new_n16772_), .A2(\A[492] ), .ZN(new_n16773_));
  INV_X1     g15753(.I(\A[492] ), .ZN(new_n16774_));
  NAND2_X1   g15754(.A1(new_n16774_), .A2(\A[491] ), .ZN(new_n16775_));
  AOI21_X1   g15755(.A1(new_n16773_), .A2(new_n16775_), .B(new_n16771_), .ZN(new_n16776_));
  NAND2_X1   g15756(.A1(new_n16772_), .A2(new_n16774_), .ZN(new_n16777_));
  NAND2_X1   g15757(.A1(\A[491] ), .A2(\A[492] ), .ZN(new_n16778_));
  AOI21_X1   g15758(.A1(new_n16777_), .A2(new_n16778_), .B(\A[490] ), .ZN(new_n16779_));
  NOR2_X1    g15759(.A1(new_n16779_), .A2(new_n16776_), .ZN(new_n16780_));
  NAND2_X1   g15760(.A1(new_n16778_), .A2(new_n16771_), .ZN(new_n16781_));
  NAND2_X1   g15761(.A1(new_n16781_), .A2(new_n16777_), .ZN(new_n16782_));
  NAND2_X1   g15762(.A1(new_n16768_), .A2(new_n16761_), .ZN(new_n16783_));
  NAND2_X1   g15763(.A1(new_n16783_), .A2(new_n16767_), .ZN(new_n16784_));
  NOR2_X1    g15764(.A1(new_n16782_), .A2(new_n16784_), .ZN(new_n16785_));
  NOR2_X1    g15765(.A1(new_n16756_), .A2(new_n16760_), .ZN(new_n16786_));
  NOR2_X1    g15766(.A1(new_n16730_), .A2(new_n16786_), .ZN(new_n16787_));
  AOI21_X1   g15767(.A1(new_n16720_), .A2(new_n16726_), .B(new_n16787_), .ZN(new_n16788_));
  INV_X1     g15768(.I(new_n16788_), .ZN(new_n16789_));
  NAND3_X1   g15769(.A1(new_n16720_), .A2(new_n16726_), .A3(new_n16787_), .ZN(new_n16790_));
  INV_X1     g15770(.I(new_n16752_), .ZN(new_n16791_));
  INV_X1     g15771(.I(new_n16754_), .ZN(new_n16792_));
  NAND2_X1   g15772(.A1(new_n16749_), .A2(new_n16792_), .ZN(new_n16793_));
  INV_X1     g15773(.I(new_n16793_), .ZN(new_n16794_));
  NOR2_X1    g15774(.A1(new_n16749_), .A2(new_n16792_), .ZN(new_n16795_));
  OAI21_X1   g15775(.A1(new_n16794_), .A2(new_n16795_), .B(new_n16791_), .ZN(new_n16796_));
  INV_X1     g15776(.I(new_n16795_), .ZN(new_n16797_));
  NAND3_X1   g15777(.A1(new_n16797_), .A2(new_n16793_), .A3(new_n16752_), .ZN(new_n16798_));
  AND2_X2    g15778(.A1(new_n16796_), .A2(new_n16798_), .Z(new_n16799_));
  OR2_X2     g15779(.A1(new_n16756_), .A2(new_n16760_), .Z(new_n16800_));
  NOR4_X1    g15780(.A1(new_n16766_), .A2(new_n16769_), .A3(new_n16779_), .A4(new_n16776_), .ZN(new_n16801_));
  NOR2_X1    g15781(.A1(new_n16770_), .A2(new_n16780_), .ZN(new_n16802_));
  OR2_X2     g15782(.A1(new_n16802_), .A2(new_n16801_), .Z(new_n16803_));
  NOR2_X1    g15783(.A1(new_n16800_), .A2(new_n16803_), .ZN(new_n16804_));
  XOR2_X1    g15784(.A1(new_n16757_), .A2(new_n16758_), .Z(new_n16805_));
  NAND2_X1   g15785(.A1(new_n16805_), .A2(new_n16755_), .ZN(new_n16806_));
  NAND3_X1   g15786(.A1(new_n16806_), .A2(new_n16801_), .A3(new_n16785_), .ZN(new_n16807_));
  AOI21_X1   g15787(.A1(new_n16799_), .A2(new_n16804_), .B(new_n16807_), .ZN(new_n16808_));
  INV_X1     g15788(.I(new_n16782_), .ZN(new_n16809_));
  NOR2_X1    g15789(.A1(new_n16801_), .A2(new_n16784_), .ZN(new_n16810_));
  NAND2_X1   g15790(.A1(new_n16801_), .A2(new_n16784_), .ZN(new_n16811_));
  INV_X1     g15791(.I(new_n16811_), .ZN(new_n16812_));
  OAI21_X1   g15792(.A1(new_n16812_), .A2(new_n16810_), .B(new_n16809_), .ZN(new_n16813_));
  INV_X1     g15793(.I(new_n16810_), .ZN(new_n16814_));
  NAND3_X1   g15794(.A1(new_n16814_), .A2(new_n16782_), .A3(new_n16811_), .ZN(new_n16815_));
  NAND2_X1   g15795(.A1(new_n16813_), .A2(new_n16815_), .ZN(new_n16816_));
  NAND2_X1   g15796(.A1(new_n16808_), .A2(new_n16816_), .ZN(new_n16817_));
  NAND2_X1   g15797(.A1(new_n16801_), .A2(new_n16785_), .ZN(new_n16818_));
  OR4_X2     g15798(.A1(new_n16756_), .A2(new_n16803_), .A3(new_n16760_), .A4(new_n16818_), .Z(new_n16819_));
  NAND2_X1   g15799(.A1(new_n16819_), .A2(new_n16816_), .ZN(new_n16820_));
  AOI21_X1   g15800(.A1(new_n16814_), .A2(new_n16811_), .B(new_n16782_), .ZN(new_n16821_));
  NOR3_X1    g15801(.A1(new_n16812_), .A2(new_n16809_), .A3(new_n16810_), .ZN(new_n16822_));
  NOR2_X1    g15802(.A1(new_n16821_), .A2(new_n16822_), .ZN(new_n16823_));
  OR3_X2     g15803(.A1(new_n16818_), .A2(new_n16801_), .A3(new_n16802_), .Z(new_n16824_));
  NOR2_X1    g15804(.A1(new_n16800_), .A2(new_n16824_), .ZN(new_n16825_));
  AOI22_X1   g15805(.A1(new_n16799_), .A2(new_n16806_), .B1(new_n16825_), .B2(new_n16823_), .ZN(new_n16826_));
  NAND3_X1   g15806(.A1(new_n16806_), .A2(new_n16796_), .A3(new_n16798_), .ZN(new_n16827_));
  NOR3_X1    g15807(.A1(new_n16819_), .A2(new_n16827_), .A3(new_n16816_), .ZN(new_n16828_));
  OAI21_X1   g15808(.A1(new_n16826_), .A2(new_n16828_), .B(new_n16820_), .ZN(new_n16829_));
  NAND2_X1   g15809(.A1(new_n16829_), .A2(new_n16817_), .ZN(new_n16830_));
  AOI22_X1   g15810(.A1(new_n16789_), .A2(new_n16790_), .B1(new_n16727_), .B2(new_n16830_), .ZN(new_n16831_));
  INV_X1     g15811(.I(new_n16725_), .ZN(new_n16832_));
  AOI21_X1   g15812(.A1(new_n16703_), .A2(new_n16718_), .B(new_n16650_), .ZN(new_n16833_));
  NOR2_X1    g15813(.A1(new_n16654_), .A2(new_n16659_), .ZN(new_n16834_));
  OAI21_X1   g15814(.A1(new_n16697_), .A2(new_n16834_), .B(new_n16662_), .ZN(new_n16835_));
  NOR2_X1    g15815(.A1(new_n16623_), .A2(new_n16628_), .ZN(new_n16836_));
  OAI21_X1   g15816(.A1(new_n16644_), .A2(new_n16836_), .B(new_n16711_), .ZN(new_n16837_));
  XNOR2_X1   g15817(.A1(new_n16837_), .A2(new_n16835_), .ZN(new_n16838_));
  INV_X1     g15818(.I(new_n16838_), .ZN(new_n16839_));
  NOR3_X1    g15819(.A1(new_n16833_), .A2(new_n16832_), .A3(new_n16839_), .ZN(new_n16840_));
  AOI21_X1   g15820(.A1(new_n16825_), .A2(new_n16827_), .B(new_n16823_), .ZN(new_n16841_));
  OAI21_X1   g15821(.A1(new_n16791_), .A2(new_n16792_), .B(new_n16750_), .ZN(new_n16842_));
  OAI21_X1   g15822(.A1(new_n16752_), .A2(new_n16754_), .B(new_n16842_), .ZN(new_n16843_));
  NAND2_X1   g15823(.A1(new_n16782_), .A2(new_n16784_), .ZN(new_n16844_));
  NAND2_X1   g15824(.A1(new_n16801_), .A2(new_n16844_), .ZN(new_n16845_));
  OAI21_X1   g15825(.A1(new_n16782_), .A2(new_n16784_), .B(new_n16845_), .ZN(new_n16846_));
  XOR2_X1    g15826(.A1(new_n16843_), .A2(new_n16846_), .Z(new_n16847_));
  NOR3_X1    g15827(.A1(new_n16847_), .A2(new_n16808_), .A3(new_n16841_), .ZN(new_n16848_));
  NAND3_X1   g15828(.A1(new_n16831_), .A2(new_n16840_), .A3(new_n16848_), .ZN(new_n16849_));
  NAND2_X1   g15829(.A1(new_n16843_), .A2(new_n16846_), .ZN(new_n16850_));
  NOR2_X1    g15830(.A1(new_n16808_), .A2(new_n16841_), .ZN(new_n16851_));
  OAI21_X1   g15831(.A1(new_n16843_), .A2(new_n16846_), .B(new_n16851_), .ZN(new_n16852_));
  NAND2_X1   g15832(.A1(new_n16852_), .A2(new_n16850_), .ZN(new_n16853_));
  NAND2_X1   g15833(.A1(new_n16837_), .A2(new_n16835_), .ZN(new_n16854_));
  NOR2_X1    g15834(.A1(new_n16833_), .A2(new_n16832_), .ZN(new_n16855_));
  OAI21_X1   g15835(.A1(new_n16835_), .A2(new_n16837_), .B(new_n16855_), .ZN(new_n16856_));
  NAND2_X1   g15836(.A1(new_n16856_), .A2(new_n16854_), .ZN(new_n16857_));
  OAI21_X1   g15837(.A1(new_n16853_), .A2(new_n16857_), .B(new_n16849_), .ZN(new_n16858_));
  NAND2_X1   g15838(.A1(new_n16857_), .A2(new_n16853_), .ZN(new_n16859_));
  NAND2_X1   g15839(.A1(new_n16858_), .A2(new_n16859_), .ZN(new_n16860_));
  INV_X1     g15840(.I(\A[478] ), .ZN(new_n16861_));
  NOR2_X1    g15841(.A1(\A[479] ), .A2(\A[480] ), .ZN(new_n16862_));
  NAND2_X1   g15842(.A1(\A[479] ), .A2(\A[480] ), .ZN(new_n16863_));
  AOI21_X1   g15843(.A1(new_n16861_), .A2(new_n16863_), .B(new_n16862_), .ZN(new_n16864_));
  NOR2_X1    g15844(.A1(\A[476] ), .A2(\A[477] ), .ZN(new_n16865_));
  INV_X1     g15845(.I(\A[476] ), .ZN(new_n16866_));
  INV_X1     g15846(.I(\A[477] ), .ZN(new_n16867_));
  NOR2_X1    g15847(.A1(new_n16866_), .A2(new_n16867_), .ZN(new_n16868_));
  NOR2_X1    g15848(.A1(new_n16868_), .A2(\A[475] ), .ZN(new_n16869_));
  NOR2_X1    g15849(.A1(new_n16869_), .A2(new_n16865_), .ZN(new_n16870_));
  NOR2_X1    g15850(.A1(new_n16867_), .A2(\A[476] ), .ZN(new_n16871_));
  NOR2_X1    g15851(.A1(new_n16866_), .A2(\A[477] ), .ZN(new_n16872_));
  OAI21_X1   g15852(.A1(new_n16871_), .A2(new_n16872_), .B(\A[475] ), .ZN(new_n16873_));
  INV_X1     g15853(.I(\A[475] ), .ZN(new_n16874_));
  OAI21_X1   g15854(.A1(new_n16868_), .A2(new_n16865_), .B(new_n16874_), .ZN(new_n16875_));
  NAND2_X1   g15855(.A1(new_n16875_), .A2(new_n16873_), .ZN(new_n16876_));
  INV_X1     g15856(.I(\A[479] ), .ZN(new_n16877_));
  NAND2_X1   g15857(.A1(new_n16877_), .A2(\A[480] ), .ZN(new_n16878_));
  INV_X1     g15858(.I(\A[480] ), .ZN(new_n16879_));
  NAND2_X1   g15859(.A1(new_n16879_), .A2(\A[479] ), .ZN(new_n16880_));
  AOI21_X1   g15860(.A1(new_n16878_), .A2(new_n16880_), .B(new_n16861_), .ZN(new_n16881_));
  INV_X1     g15861(.I(new_n16862_), .ZN(new_n16882_));
  AOI21_X1   g15862(.A1(new_n16882_), .A2(new_n16863_), .B(\A[478] ), .ZN(new_n16883_));
  NOR3_X1    g15863(.A1(new_n16876_), .A2(new_n16881_), .A3(new_n16883_), .ZN(new_n16884_));
  XOR2_X1    g15864(.A1(new_n16884_), .A2(new_n16870_), .Z(new_n16885_));
  XOR2_X1    g15865(.A1(new_n16885_), .A2(new_n16864_), .Z(new_n16886_));
  INV_X1     g15866(.I(\A[484] ), .ZN(new_n16887_));
  NOR2_X1    g15867(.A1(\A[485] ), .A2(\A[486] ), .ZN(new_n16888_));
  NAND2_X1   g15868(.A1(\A[485] ), .A2(\A[486] ), .ZN(new_n16889_));
  AOI21_X1   g15869(.A1(new_n16887_), .A2(new_n16889_), .B(new_n16888_), .ZN(new_n16890_));
  INV_X1     g15870(.I(new_n16890_), .ZN(new_n16891_));
  INV_X1     g15871(.I(\A[481] ), .ZN(new_n16892_));
  NOR2_X1    g15872(.A1(\A[482] ), .A2(\A[483] ), .ZN(new_n16893_));
  NAND2_X1   g15873(.A1(\A[482] ), .A2(\A[483] ), .ZN(new_n16894_));
  AOI21_X1   g15874(.A1(new_n16892_), .A2(new_n16894_), .B(new_n16893_), .ZN(new_n16895_));
  INV_X1     g15875(.I(new_n16895_), .ZN(new_n16896_));
  NOR2_X1    g15876(.A1(new_n16891_), .A2(new_n16896_), .ZN(new_n16897_));
  INV_X1     g15877(.I(new_n16897_), .ZN(new_n16898_));
  INV_X1     g15878(.I(\A[482] ), .ZN(new_n16899_));
  NAND2_X1   g15879(.A1(new_n16899_), .A2(\A[483] ), .ZN(new_n16900_));
  INV_X1     g15880(.I(\A[483] ), .ZN(new_n16901_));
  NAND2_X1   g15881(.A1(new_n16901_), .A2(\A[482] ), .ZN(new_n16902_));
  AOI21_X1   g15882(.A1(new_n16900_), .A2(new_n16902_), .B(new_n16892_), .ZN(new_n16903_));
  INV_X1     g15883(.I(new_n16893_), .ZN(new_n16904_));
  AOI21_X1   g15884(.A1(new_n16904_), .A2(new_n16894_), .B(\A[481] ), .ZN(new_n16905_));
  NOR2_X1    g15885(.A1(new_n16905_), .A2(new_n16903_), .ZN(new_n16906_));
  INV_X1     g15886(.I(\A[486] ), .ZN(new_n16907_));
  NOR2_X1    g15887(.A1(new_n16907_), .A2(\A[485] ), .ZN(new_n16908_));
  INV_X1     g15888(.I(\A[485] ), .ZN(new_n16909_));
  NOR2_X1    g15889(.A1(new_n16909_), .A2(\A[486] ), .ZN(new_n16910_));
  OAI21_X1   g15890(.A1(new_n16908_), .A2(new_n16910_), .B(\A[484] ), .ZN(new_n16911_));
  INV_X1     g15891(.I(new_n16889_), .ZN(new_n16912_));
  OAI21_X1   g15892(.A1(new_n16912_), .A2(new_n16888_), .B(new_n16887_), .ZN(new_n16913_));
  NAND2_X1   g15893(.A1(new_n16911_), .A2(new_n16913_), .ZN(new_n16914_));
  NAND2_X1   g15894(.A1(new_n16906_), .A2(new_n16914_), .ZN(new_n16915_));
  NOR2_X1    g15895(.A1(new_n16901_), .A2(\A[482] ), .ZN(new_n16916_));
  NOR2_X1    g15896(.A1(new_n16899_), .A2(\A[483] ), .ZN(new_n16917_));
  OAI21_X1   g15897(.A1(new_n16916_), .A2(new_n16917_), .B(\A[481] ), .ZN(new_n16918_));
  INV_X1     g15898(.I(new_n16894_), .ZN(new_n16919_));
  OAI21_X1   g15899(.A1(new_n16919_), .A2(new_n16893_), .B(new_n16892_), .ZN(new_n16920_));
  NAND2_X1   g15900(.A1(new_n16918_), .A2(new_n16920_), .ZN(new_n16921_));
  NAND2_X1   g15901(.A1(new_n16909_), .A2(\A[486] ), .ZN(new_n16922_));
  NAND2_X1   g15902(.A1(new_n16907_), .A2(\A[485] ), .ZN(new_n16923_));
  AOI21_X1   g15903(.A1(new_n16922_), .A2(new_n16923_), .B(new_n16887_), .ZN(new_n16924_));
  INV_X1     g15904(.I(new_n16888_), .ZN(new_n16925_));
  AOI21_X1   g15905(.A1(new_n16925_), .A2(new_n16889_), .B(\A[484] ), .ZN(new_n16926_));
  NOR2_X1    g15906(.A1(new_n16926_), .A2(new_n16924_), .ZN(new_n16927_));
  NAND2_X1   g15907(.A1(new_n16927_), .A2(new_n16921_), .ZN(new_n16928_));
  AOI21_X1   g15908(.A1(new_n16915_), .A2(new_n16928_), .B(new_n16898_), .ZN(new_n16929_));
  INV_X1     g15909(.I(new_n16929_), .ZN(new_n16930_));
  NOR2_X1    g15910(.A1(new_n16921_), .A2(new_n16914_), .ZN(new_n16931_));
  NOR2_X1    g15911(.A1(new_n16931_), .A2(new_n16896_), .ZN(new_n16932_));
  NAND2_X1   g15912(.A1(new_n16906_), .A2(new_n16927_), .ZN(new_n16933_));
  NOR2_X1    g15913(.A1(new_n16933_), .A2(new_n16895_), .ZN(new_n16934_));
  OAI21_X1   g15914(.A1(new_n16932_), .A2(new_n16934_), .B(new_n16890_), .ZN(new_n16935_));
  NAND2_X1   g15915(.A1(new_n16933_), .A2(new_n16895_), .ZN(new_n16936_));
  NAND2_X1   g15916(.A1(new_n16931_), .A2(new_n16896_), .ZN(new_n16937_));
  NAND3_X1   g15917(.A1(new_n16937_), .A2(new_n16936_), .A3(new_n16891_), .ZN(new_n16938_));
  NAND3_X1   g15918(.A1(new_n16935_), .A2(new_n16938_), .A3(new_n16930_), .ZN(new_n16939_));
  NOR2_X1    g15919(.A1(new_n16933_), .A2(new_n16898_), .ZN(new_n16940_));
  NOR2_X1    g15920(.A1(new_n16906_), .A2(new_n16927_), .ZN(new_n16941_));
  NOR2_X1    g15921(.A1(new_n16941_), .A2(new_n16931_), .ZN(new_n16942_));
  INV_X1     g15922(.I(new_n16876_), .ZN(new_n16943_));
  NOR2_X1    g15923(.A1(new_n16883_), .A2(new_n16881_), .ZN(new_n16944_));
  NOR2_X1    g15924(.A1(new_n16943_), .A2(new_n16944_), .ZN(new_n16945_));
  NOR2_X1    g15925(.A1(new_n16945_), .A2(new_n16884_), .ZN(new_n16946_));
  NAND2_X1   g15926(.A1(new_n16943_), .A2(new_n16944_), .ZN(new_n16947_));
  NAND2_X1   g15927(.A1(new_n16870_), .A2(new_n16864_), .ZN(new_n16948_));
  NOR2_X1    g15928(.A1(new_n16947_), .A2(new_n16948_), .ZN(new_n16949_));
  NAND4_X1   g15929(.A1(new_n16946_), .A2(new_n16949_), .A3(new_n16940_), .A4(new_n16942_), .ZN(new_n16950_));
  NOR2_X1    g15930(.A1(new_n16939_), .A2(new_n16950_), .ZN(new_n16951_));
  AOI21_X1   g15931(.A1(new_n16937_), .A2(new_n16936_), .B(new_n16891_), .ZN(new_n16952_));
  NOR3_X1    g15932(.A1(new_n16932_), .A2(new_n16934_), .A3(new_n16890_), .ZN(new_n16953_));
  NOR3_X1    g15933(.A1(new_n16952_), .A2(new_n16953_), .A3(new_n16929_), .ZN(new_n16954_));
  INV_X1     g15934(.I(new_n16950_), .ZN(new_n16955_));
  NOR2_X1    g15935(.A1(new_n16955_), .A2(new_n16954_), .ZN(new_n16956_));
  OAI21_X1   g15936(.A1(new_n16951_), .A2(new_n16956_), .B(new_n16886_), .ZN(new_n16957_));
  NAND2_X1   g15937(.A1(new_n16955_), .A2(new_n16939_), .ZN(new_n16958_));
  NAND2_X1   g15938(.A1(new_n16935_), .A2(new_n16938_), .ZN(new_n16959_));
  NAND3_X1   g15939(.A1(new_n16946_), .A2(new_n16940_), .A3(new_n16942_), .ZN(new_n16960_));
  NOR3_X1    g15940(.A1(new_n16929_), .A2(new_n16947_), .A3(new_n16948_), .ZN(new_n16961_));
  OAI21_X1   g15941(.A1(new_n16959_), .A2(new_n16960_), .B(new_n16961_), .ZN(new_n16962_));
  NAND3_X1   g15942(.A1(new_n16886_), .A2(new_n16958_), .A3(new_n16962_), .ZN(new_n16963_));
  NAND2_X1   g15943(.A1(new_n16957_), .A2(new_n16963_), .ZN(new_n16964_));
  INV_X1     g15944(.I(new_n16964_), .ZN(new_n16965_));
  INV_X1     g15945(.I(\A[471] ), .ZN(new_n16966_));
  NOR2_X1    g15946(.A1(new_n16966_), .A2(\A[470] ), .ZN(new_n16967_));
  INV_X1     g15947(.I(\A[470] ), .ZN(new_n16968_));
  NOR2_X1    g15948(.A1(new_n16968_), .A2(\A[471] ), .ZN(new_n16969_));
  OAI21_X1   g15949(.A1(new_n16967_), .A2(new_n16969_), .B(\A[469] ), .ZN(new_n16970_));
  INV_X1     g15950(.I(\A[469] ), .ZN(new_n16971_));
  NOR2_X1    g15951(.A1(\A[470] ), .A2(\A[471] ), .ZN(new_n16972_));
  NAND2_X1   g15952(.A1(\A[470] ), .A2(\A[471] ), .ZN(new_n16973_));
  INV_X1     g15953(.I(new_n16973_), .ZN(new_n16974_));
  OAI21_X1   g15954(.A1(new_n16974_), .A2(new_n16972_), .B(new_n16971_), .ZN(new_n16975_));
  NAND2_X1   g15955(.A1(new_n16970_), .A2(new_n16975_), .ZN(new_n16976_));
  INV_X1     g15956(.I(\A[474] ), .ZN(new_n16977_));
  NOR2_X1    g15957(.A1(new_n16977_), .A2(\A[473] ), .ZN(new_n16978_));
  INV_X1     g15958(.I(\A[473] ), .ZN(new_n16979_));
  NOR2_X1    g15959(.A1(new_n16979_), .A2(\A[474] ), .ZN(new_n16980_));
  OAI21_X1   g15960(.A1(new_n16978_), .A2(new_n16980_), .B(\A[472] ), .ZN(new_n16981_));
  INV_X1     g15961(.I(\A[472] ), .ZN(new_n16982_));
  NOR2_X1    g15962(.A1(\A[473] ), .A2(\A[474] ), .ZN(new_n16983_));
  NAND2_X1   g15963(.A1(\A[473] ), .A2(\A[474] ), .ZN(new_n16984_));
  INV_X1     g15964(.I(new_n16984_), .ZN(new_n16985_));
  OAI21_X1   g15965(.A1(new_n16985_), .A2(new_n16983_), .B(new_n16982_), .ZN(new_n16986_));
  NAND2_X1   g15966(.A1(new_n16981_), .A2(new_n16986_), .ZN(new_n16987_));
  NOR2_X1    g15967(.A1(new_n16976_), .A2(new_n16987_), .ZN(new_n16988_));
  AOI21_X1   g15968(.A1(new_n16982_), .A2(new_n16984_), .B(new_n16983_), .ZN(new_n16989_));
  INV_X1     g15969(.I(new_n16989_), .ZN(new_n16990_));
  AOI21_X1   g15970(.A1(new_n16971_), .A2(new_n16973_), .B(new_n16972_), .ZN(new_n16991_));
  INV_X1     g15971(.I(new_n16991_), .ZN(new_n16992_));
  NOR2_X1    g15972(.A1(new_n16990_), .A2(new_n16992_), .ZN(new_n16993_));
  NAND2_X1   g15973(.A1(new_n16988_), .A2(new_n16993_), .ZN(new_n16994_));
  NAND2_X1   g15974(.A1(new_n16968_), .A2(\A[471] ), .ZN(new_n16995_));
  NAND2_X1   g15975(.A1(new_n16966_), .A2(\A[470] ), .ZN(new_n16996_));
  AOI21_X1   g15976(.A1(new_n16995_), .A2(new_n16996_), .B(new_n16971_), .ZN(new_n16997_));
  INV_X1     g15977(.I(new_n16972_), .ZN(new_n16998_));
  AOI21_X1   g15978(.A1(new_n16998_), .A2(new_n16973_), .B(\A[469] ), .ZN(new_n16999_));
  NOR2_X1    g15979(.A1(new_n16999_), .A2(new_n16997_), .ZN(new_n17000_));
  NAND2_X1   g15980(.A1(new_n16979_), .A2(\A[474] ), .ZN(new_n17001_));
  NAND2_X1   g15981(.A1(new_n16977_), .A2(\A[473] ), .ZN(new_n17002_));
  AOI21_X1   g15982(.A1(new_n17001_), .A2(new_n17002_), .B(new_n16982_), .ZN(new_n17003_));
  INV_X1     g15983(.I(new_n16983_), .ZN(new_n17004_));
  AOI21_X1   g15984(.A1(new_n17004_), .A2(new_n16984_), .B(\A[472] ), .ZN(new_n17005_));
  NOR2_X1    g15985(.A1(new_n17005_), .A2(new_n17003_), .ZN(new_n17006_));
  NAND2_X1   g15986(.A1(new_n17000_), .A2(new_n17006_), .ZN(new_n17007_));
  NAND2_X1   g15987(.A1(new_n16976_), .A2(new_n16987_), .ZN(new_n17008_));
  NAND2_X1   g15988(.A1(new_n17007_), .A2(new_n17008_), .ZN(new_n17009_));
  INV_X1     g15989(.I(\A[466] ), .ZN(new_n17010_));
  INV_X1     g15990(.I(\A[467] ), .ZN(new_n17011_));
  NAND2_X1   g15991(.A1(new_n17011_), .A2(\A[468] ), .ZN(new_n17012_));
  INV_X1     g15992(.I(\A[468] ), .ZN(new_n17013_));
  NAND2_X1   g15993(.A1(new_n17013_), .A2(\A[467] ), .ZN(new_n17014_));
  AOI21_X1   g15994(.A1(new_n17012_), .A2(new_n17014_), .B(new_n17010_), .ZN(new_n17015_));
  NAND2_X1   g15995(.A1(new_n17011_), .A2(new_n17013_), .ZN(new_n17016_));
  NAND2_X1   g15996(.A1(\A[467] ), .A2(\A[468] ), .ZN(new_n17017_));
  AOI21_X1   g15997(.A1(new_n17016_), .A2(new_n17017_), .B(\A[466] ), .ZN(new_n17018_));
  NOR2_X1    g15998(.A1(new_n17018_), .A2(new_n17015_), .ZN(new_n17019_));
  INV_X1     g15999(.I(\A[463] ), .ZN(new_n17020_));
  INV_X1     g16000(.I(\A[464] ), .ZN(new_n17021_));
  NAND2_X1   g16001(.A1(new_n17021_), .A2(\A[465] ), .ZN(new_n17022_));
  INV_X1     g16002(.I(\A[465] ), .ZN(new_n17023_));
  NAND2_X1   g16003(.A1(new_n17023_), .A2(\A[464] ), .ZN(new_n17024_));
  AOI21_X1   g16004(.A1(new_n17022_), .A2(new_n17024_), .B(new_n17020_), .ZN(new_n17025_));
  NAND2_X1   g16005(.A1(new_n17021_), .A2(new_n17023_), .ZN(new_n17026_));
  NAND2_X1   g16006(.A1(\A[464] ), .A2(\A[465] ), .ZN(new_n17027_));
  AOI21_X1   g16007(.A1(new_n17026_), .A2(new_n17027_), .B(\A[463] ), .ZN(new_n17028_));
  NOR2_X1    g16008(.A1(new_n17028_), .A2(new_n17025_), .ZN(new_n17029_));
  NAND2_X1   g16009(.A1(new_n17017_), .A2(new_n17010_), .ZN(new_n17030_));
  NAND2_X1   g16010(.A1(new_n17030_), .A2(new_n17016_), .ZN(new_n17031_));
  NAND2_X1   g16011(.A1(new_n17027_), .A2(new_n17020_), .ZN(new_n17032_));
  NAND2_X1   g16012(.A1(new_n17032_), .A2(new_n17026_), .ZN(new_n17033_));
  NOR2_X1    g16013(.A1(new_n17031_), .A2(new_n17033_), .ZN(new_n17034_));
  NOR2_X1    g16014(.A1(new_n17009_), .A2(new_n16994_), .ZN(new_n17035_));
  NAND2_X1   g16015(.A1(new_n16942_), .A2(new_n16940_), .ZN(new_n17036_));
  NAND2_X1   g16016(.A1(new_n16946_), .A2(new_n16949_), .ZN(new_n17037_));
  XOR2_X1    g16017(.A1(new_n17037_), .A2(new_n17036_), .Z(new_n17038_));
  NOR2_X1    g16018(.A1(new_n17038_), .A2(new_n17035_), .ZN(new_n17039_));
  NAND2_X1   g16019(.A1(new_n16965_), .A2(new_n17039_), .ZN(new_n17040_));
  AOI21_X1   g16020(.A1(new_n16957_), .A2(new_n16963_), .B(new_n17039_), .ZN(new_n17041_));
  NAND3_X1   g16021(.A1(new_n16957_), .A2(new_n17039_), .A3(new_n16963_), .ZN(new_n17042_));
  INV_X1     g16022(.I(new_n17042_), .ZN(new_n17043_));
  INV_X1     g16023(.I(new_n16993_), .ZN(new_n17044_));
  NOR2_X1    g16024(.A1(new_n17007_), .A2(new_n17044_), .ZN(new_n17045_));
  NAND3_X1   g16025(.A1(new_n17045_), .A2(new_n17007_), .A3(new_n17008_), .ZN(new_n17046_));
  XNOR2_X1   g16026(.A1(new_n17019_), .A2(new_n17029_), .ZN(new_n17047_));
  NAND2_X1   g16027(.A1(new_n17007_), .A2(new_n16991_), .ZN(new_n17048_));
  NAND2_X1   g16028(.A1(new_n16988_), .A2(new_n16992_), .ZN(new_n17049_));
  AOI21_X1   g16029(.A1(new_n17049_), .A2(new_n17048_), .B(new_n16990_), .ZN(new_n17050_));
  NOR2_X1    g16030(.A1(new_n16988_), .A2(new_n16992_), .ZN(new_n17051_));
  NOR2_X1    g16031(.A1(new_n17007_), .A2(new_n16991_), .ZN(new_n17052_));
  NOR3_X1    g16032(.A1(new_n17051_), .A2(new_n17052_), .A3(new_n16989_), .ZN(new_n17053_));
  NOR4_X1    g16033(.A1(new_n17050_), .A2(new_n17053_), .A3(new_n17046_), .A4(new_n17047_), .ZN(new_n17054_));
  NOR4_X1    g16034(.A1(new_n17015_), .A2(new_n17018_), .A3(new_n17028_), .A4(new_n17025_), .ZN(new_n17055_));
  NOR2_X1    g16035(.A1(new_n17006_), .A2(new_n16976_), .ZN(new_n17056_));
  NOR2_X1    g16036(.A1(new_n17000_), .A2(new_n16987_), .ZN(new_n17057_));
  OAI21_X1   g16037(.A1(new_n17056_), .A2(new_n17057_), .B(new_n16993_), .ZN(new_n17058_));
  NAND3_X1   g16038(.A1(new_n17058_), .A2(new_n17055_), .A3(new_n17034_), .ZN(new_n17059_));
  NOR2_X1    g16039(.A1(new_n17054_), .A2(new_n17059_), .ZN(new_n17060_));
  INV_X1     g16040(.I(new_n17031_), .ZN(new_n17061_));
  NOR2_X1    g16041(.A1(new_n17055_), .A2(new_n17033_), .ZN(new_n17062_));
  NAND2_X1   g16042(.A1(new_n17055_), .A2(new_n17033_), .ZN(new_n17063_));
  INV_X1     g16043(.I(new_n17063_), .ZN(new_n17064_));
  OAI21_X1   g16044(.A1(new_n17064_), .A2(new_n17062_), .B(new_n17061_), .ZN(new_n17065_));
  INV_X1     g16045(.I(new_n17062_), .ZN(new_n17066_));
  NAND3_X1   g16046(.A1(new_n17066_), .A2(new_n17031_), .A3(new_n17063_), .ZN(new_n17067_));
  NAND2_X1   g16047(.A1(new_n17065_), .A2(new_n17067_), .ZN(new_n17068_));
  NAND2_X1   g16048(.A1(new_n17055_), .A2(new_n17034_), .ZN(new_n17069_));
  OR4_X2     g16049(.A1(new_n16994_), .A2(new_n17047_), .A3(new_n17009_), .A4(new_n17069_), .Z(new_n17070_));
  NAND2_X1   g16050(.A1(new_n17070_), .A2(new_n17068_), .ZN(new_n17071_));
  OAI21_X1   g16051(.A1(new_n17051_), .A2(new_n17052_), .B(new_n16989_), .ZN(new_n17072_));
  NAND3_X1   g16052(.A1(new_n17049_), .A2(new_n17048_), .A3(new_n16990_), .ZN(new_n17073_));
  NAND3_X1   g16053(.A1(new_n17072_), .A2(new_n17073_), .A3(new_n17058_), .ZN(new_n17074_));
  OAI21_X1   g16054(.A1(new_n17070_), .A2(new_n17068_), .B(new_n17074_), .ZN(new_n17075_));
  NOR3_X1    g16055(.A1(new_n17070_), .A2(new_n17074_), .A3(new_n17068_), .ZN(new_n17076_));
  INV_X1     g16056(.I(new_n17076_), .ZN(new_n17077_));
  NAND2_X1   g16057(.A1(new_n17077_), .A2(new_n17075_), .ZN(new_n17078_));
  AOI22_X1   g16058(.A1(new_n17078_), .A2(new_n17071_), .B1(new_n17060_), .B2(new_n17068_), .ZN(new_n17079_));
  OAI21_X1   g16059(.A1(new_n17043_), .A2(new_n17041_), .B(new_n17079_), .ZN(new_n17080_));
  XNOR2_X1   g16060(.A1(new_n16885_), .A2(new_n16864_), .ZN(new_n17081_));
  NAND2_X1   g16061(.A1(new_n17081_), .A2(new_n16958_), .ZN(new_n17082_));
  NOR2_X1    g16062(.A1(new_n16890_), .A2(new_n16895_), .ZN(new_n17083_));
  OAI21_X1   g16063(.A1(new_n16933_), .A2(new_n17083_), .B(new_n16898_), .ZN(new_n17084_));
  NOR2_X1    g16064(.A1(new_n16870_), .A2(new_n16864_), .ZN(new_n17085_));
  OAI21_X1   g16065(.A1(new_n16947_), .A2(new_n17085_), .B(new_n16948_), .ZN(new_n17086_));
  XNOR2_X1   g16066(.A1(new_n17086_), .A2(new_n17084_), .ZN(new_n17087_));
  NAND3_X1   g16067(.A1(new_n17082_), .A2(new_n16962_), .A3(new_n17087_), .ZN(new_n17088_));
  NOR3_X1    g16068(.A1(new_n17046_), .A2(new_n17069_), .A3(new_n17047_), .ZN(new_n17089_));
  AOI22_X1   g16069(.A1(new_n17074_), .A2(new_n17089_), .B1(new_n17065_), .B2(new_n17067_), .ZN(new_n17090_));
  NOR2_X1    g16070(.A1(new_n16989_), .A2(new_n16991_), .ZN(new_n17091_));
  OAI21_X1   g16071(.A1(new_n17007_), .A2(new_n17091_), .B(new_n17044_), .ZN(new_n17092_));
  NAND2_X1   g16072(.A1(new_n17031_), .A2(new_n17033_), .ZN(new_n17093_));
  NAND2_X1   g16073(.A1(new_n17055_), .A2(new_n17093_), .ZN(new_n17094_));
  OAI21_X1   g16074(.A1(new_n17031_), .A2(new_n17033_), .B(new_n17094_), .ZN(new_n17095_));
  XOR2_X1    g16075(.A1(new_n17095_), .A2(new_n17092_), .Z(new_n17096_));
  NOR3_X1    g16076(.A1(new_n17090_), .A2(new_n17060_), .A3(new_n17096_), .ZN(new_n17097_));
  INV_X1     g16077(.I(new_n17097_), .ZN(new_n17098_));
  NAND2_X1   g16078(.A1(new_n17088_), .A2(new_n17098_), .ZN(new_n17099_));
  NAND3_X1   g16079(.A1(new_n17080_), .A2(new_n17040_), .A3(new_n17099_), .ZN(new_n17100_));
  INV_X1     g16080(.I(new_n16962_), .ZN(new_n17101_));
  AOI21_X1   g16081(.A1(new_n16939_), .A2(new_n16955_), .B(new_n16886_), .ZN(new_n17102_));
  INV_X1     g16082(.I(new_n17087_), .ZN(new_n17103_));
  NOR3_X1    g16083(.A1(new_n17102_), .A2(new_n17101_), .A3(new_n17103_), .ZN(new_n17104_));
  NAND2_X1   g16084(.A1(new_n17104_), .A2(new_n17097_), .ZN(new_n17105_));
  INV_X1     g16085(.I(new_n17105_), .ZN(new_n17106_));
  NAND2_X1   g16086(.A1(new_n17095_), .A2(new_n17092_), .ZN(new_n17107_));
  NOR2_X1    g16087(.A1(new_n17090_), .A2(new_n17060_), .ZN(new_n17108_));
  OAI21_X1   g16088(.A1(new_n17092_), .A2(new_n17095_), .B(new_n17108_), .ZN(new_n17109_));
  NAND2_X1   g16089(.A1(new_n17109_), .A2(new_n17107_), .ZN(new_n17110_));
  INV_X1     g16090(.I(new_n17110_), .ZN(new_n17111_));
  NAND2_X1   g16091(.A1(new_n17086_), .A2(new_n17084_), .ZN(new_n17112_));
  NOR2_X1    g16092(.A1(new_n17102_), .A2(new_n17101_), .ZN(new_n17113_));
  OAI21_X1   g16093(.A1(new_n17084_), .A2(new_n17086_), .B(new_n17113_), .ZN(new_n17114_));
  NAND2_X1   g16094(.A1(new_n17114_), .A2(new_n17112_), .ZN(new_n17115_));
  INV_X1     g16095(.I(new_n17115_), .ZN(new_n17116_));
  AOI22_X1   g16096(.A1(new_n17100_), .A2(new_n17106_), .B1(new_n17111_), .B2(new_n17116_), .ZN(new_n17117_));
  NAND2_X1   g16097(.A1(new_n17115_), .A2(new_n17110_), .ZN(new_n17118_));
  INV_X1     g16098(.I(new_n17118_), .ZN(new_n17119_));
  NOR2_X1    g16099(.A1(new_n17117_), .A2(new_n17119_), .ZN(new_n17120_));
  INV_X1     g16100(.I(new_n17120_), .ZN(new_n17121_));
  NAND2_X1   g16101(.A1(new_n17121_), .A2(new_n16860_), .ZN(new_n17122_));
  OAI22_X1   g16102(.A1(new_n17041_), .A2(new_n17043_), .B1(new_n16965_), .B2(new_n17079_), .ZN(new_n17123_));
  XOR2_X1    g16103(.A1(new_n17088_), .A2(new_n17097_), .Z(new_n17124_));
  NOR2_X1    g16104(.A1(new_n17123_), .A2(new_n17124_), .ZN(new_n17125_));
  INV_X1     g16105(.I(new_n17035_), .ZN(new_n17126_));
  XNOR2_X1   g16106(.A1(new_n17037_), .A2(new_n17036_), .ZN(new_n17127_));
  NAND2_X1   g16107(.A1(new_n17127_), .A2(new_n17126_), .ZN(new_n17128_));
  NAND2_X1   g16108(.A1(new_n16964_), .A2(new_n17128_), .ZN(new_n17129_));
  NAND2_X1   g16109(.A1(new_n17060_), .A2(new_n17068_), .ZN(new_n17130_));
  INV_X1     g16110(.I(new_n17075_), .ZN(new_n17131_));
  OAI21_X1   g16111(.A1(new_n17131_), .A2(new_n17076_), .B(new_n17071_), .ZN(new_n17132_));
  NAND2_X1   g16112(.A1(new_n17132_), .A2(new_n17130_), .ZN(new_n17133_));
  AOI22_X1   g16113(.A1(new_n17129_), .A2(new_n17042_), .B1(new_n17133_), .B2(new_n16964_), .ZN(new_n17134_));
  AOI21_X1   g16114(.A1(new_n17099_), .A2(new_n17105_), .B(new_n17134_), .ZN(new_n17135_));
  INV_X1     g16115(.I(new_n16727_), .ZN(new_n17136_));
  INV_X1     g16116(.I(new_n16790_), .ZN(new_n17137_));
  NAND2_X1   g16117(.A1(new_n16796_), .A2(new_n16798_), .ZN(new_n17138_));
  NOR3_X1    g16118(.A1(new_n17138_), .A2(new_n16800_), .A3(new_n16803_), .ZN(new_n17139_));
  NOR3_X1    g16119(.A1(new_n17139_), .A2(new_n16807_), .A3(new_n16823_), .ZN(new_n17140_));
  NOR4_X1    g16120(.A1(new_n16800_), .A2(new_n16824_), .A3(new_n16821_), .A4(new_n16822_), .ZN(new_n17141_));
  XOR2_X1    g16121(.A1(new_n17141_), .A2(new_n16827_), .Z(new_n17142_));
  AOI21_X1   g16122(.A1(new_n17142_), .A2(new_n16820_), .B(new_n17140_), .ZN(new_n17143_));
  OAI22_X1   g16123(.A1(new_n17137_), .A2(new_n16788_), .B1(new_n17143_), .B2(new_n17136_), .ZN(new_n17144_));
  XNOR2_X1   g16124(.A1(new_n16848_), .A2(new_n16840_), .ZN(new_n17145_));
  NOR2_X1    g16125(.A1(new_n17144_), .A2(new_n17145_), .ZN(new_n17146_));
  NOR2_X1    g16126(.A1(new_n16848_), .A2(new_n16840_), .ZN(new_n17147_));
  AND2_X2    g16127(.A1(new_n16848_), .A2(new_n16840_), .Z(new_n17148_));
  NOR2_X1    g16128(.A1(new_n17148_), .A2(new_n17147_), .ZN(new_n17149_));
  NOR2_X1    g16129(.A1(new_n17149_), .A2(new_n16831_), .ZN(new_n17150_));
  NOR4_X1    g16130(.A1(new_n17135_), .A2(new_n17125_), .A3(new_n17146_), .A4(new_n17150_), .ZN(new_n17151_));
  NOR3_X1    g16131(.A1(new_n17137_), .A2(new_n16788_), .A3(new_n16830_), .ZN(new_n17152_));
  INV_X1     g16132(.I(new_n17152_), .ZN(new_n17153_));
  NAND2_X1   g16133(.A1(new_n17038_), .A2(new_n17035_), .ZN(new_n17154_));
  NAND2_X1   g16134(.A1(new_n17128_), .A2(new_n17154_), .ZN(new_n17155_));
  INV_X1     g16135(.I(new_n16787_), .ZN(new_n17156_));
  NAND2_X1   g16136(.A1(new_n16730_), .A2(new_n16786_), .ZN(new_n17157_));
  NAND2_X1   g16137(.A1(new_n17156_), .A2(new_n17157_), .ZN(new_n17158_));
  NOR2_X1    g16138(.A1(new_n17158_), .A2(new_n17155_), .ZN(new_n17159_));
  NOR2_X1    g16139(.A1(new_n17152_), .A2(new_n17159_), .ZN(new_n17160_));
  INV_X1     g16140(.I(new_n17160_), .ZN(new_n17161_));
  NAND2_X1   g16141(.A1(new_n17152_), .A2(new_n17159_), .ZN(new_n17162_));
  AOI21_X1   g16142(.A1(new_n17129_), .A2(new_n17042_), .B(new_n17133_), .ZN(new_n17163_));
  NOR3_X1    g16143(.A1(new_n17043_), .A2(new_n17079_), .A3(new_n17041_), .ZN(new_n17164_));
  OR2_X2     g16144(.A1(new_n17164_), .A2(new_n17163_), .Z(new_n17165_));
  AOI22_X1   g16145(.A1(new_n17165_), .A2(new_n17153_), .B1(new_n17161_), .B2(new_n17162_), .ZN(new_n17166_));
  OAI22_X1   g16146(.A1(new_n17135_), .A2(new_n17125_), .B1(new_n17146_), .B2(new_n17150_), .ZN(new_n17167_));
  AOI21_X1   g16147(.A1(new_n17166_), .A2(new_n17167_), .B(new_n17151_), .ZN(new_n17168_));
  AOI21_X1   g16148(.A1(new_n17100_), .A2(new_n17106_), .B(new_n17111_), .ZN(new_n17169_));
  NOR4_X1    g16149(.A1(new_n17123_), .A2(new_n17088_), .A3(new_n17098_), .A4(new_n17110_), .ZN(new_n17170_));
  OAI21_X1   g16150(.A1(new_n17169_), .A2(new_n17170_), .B(new_n17115_), .ZN(new_n17171_));
  NAND3_X1   g16151(.A1(new_n17134_), .A2(new_n17104_), .A3(new_n17097_), .ZN(new_n17172_));
  NAND2_X1   g16152(.A1(new_n17172_), .A2(new_n17110_), .ZN(new_n17173_));
  NAND4_X1   g16153(.A1(new_n17134_), .A2(new_n17111_), .A3(new_n17104_), .A4(new_n17097_), .ZN(new_n17174_));
  NAND3_X1   g16154(.A1(new_n17173_), .A2(new_n17116_), .A3(new_n17174_), .ZN(new_n17175_));
  INV_X1     g16155(.I(new_n17147_), .ZN(new_n17176_));
  NAND2_X1   g16156(.A1(new_n17144_), .A2(new_n17176_), .ZN(new_n17177_));
  INV_X1     g16157(.I(new_n16853_), .ZN(new_n17178_));
  AOI21_X1   g16158(.A1(new_n17177_), .A2(new_n17148_), .B(new_n17178_), .ZN(new_n17179_));
  NOR2_X1    g16159(.A1(new_n16849_), .A2(new_n16853_), .ZN(new_n17180_));
  OAI21_X1   g16160(.A1(new_n17179_), .A2(new_n17180_), .B(new_n16857_), .ZN(new_n17181_));
  INV_X1     g16161(.I(new_n16857_), .ZN(new_n17182_));
  NAND2_X1   g16162(.A1(new_n16849_), .A2(new_n16853_), .ZN(new_n17183_));
  NAND4_X1   g16163(.A1(new_n17178_), .A2(new_n16831_), .A3(new_n16840_), .A4(new_n16848_), .ZN(new_n17184_));
  NAND3_X1   g16164(.A1(new_n17183_), .A2(new_n17182_), .A3(new_n17184_), .ZN(new_n17185_));
  NAND4_X1   g16165(.A1(new_n17171_), .A2(new_n17175_), .A3(new_n17181_), .A4(new_n17185_), .ZN(new_n17186_));
  NAND2_X1   g16166(.A1(new_n17186_), .A2(new_n17168_), .ZN(new_n17187_));
  XOR2_X1    g16167(.A1(new_n16857_), .A2(new_n16853_), .Z(new_n17188_));
  XOR2_X1    g16168(.A1(new_n17115_), .A2(new_n17110_), .Z(new_n17189_));
  NOR4_X1    g16169(.A1(new_n17189_), .A2(new_n17188_), .A3(new_n16849_), .A4(new_n17172_), .ZN(new_n17190_));
  NAND2_X1   g16170(.A1(new_n17187_), .A2(new_n17190_), .ZN(new_n17191_));
  NAND3_X1   g16171(.A1(new_n16858_), .A2(new_n16859_), .A3(new_n17118_), .ZN(new_n17192_));
  NOR2_X1    g16172(.A1(new_n17192_), .A2(new_n17117_), .ZN(new_n17193_));
  NAND2_X1   g16173(.A1(new_n17191_), .A2(new_n17193_), .ZN(new_n17194_));
  NAND2_X1   g16174(.A1(new_n17194_), .A2(new_n17122_), .ZN(new_n17195_));
  NOR2_X1    g16175(.A1(new_n17195_), .A2(new_n16619_), .ZN(new_n17196_));
  XNOR2_X1   g16176(.A1(new_n16529_), .A2(new_n16522_), .ZN(new_n17197_));
  NAND2_X1   g16177(.A1(new_n16560_), .A2(new_n17197_), .ZN(new_n17198_));
  XOR2_X1    g16178(.A1(new_n16529_), .A2(new_n16522_), .Z(new_n17199_));
  NAND2_X1   g16179(.A1(new_n16515_), .A2(new_n17199_), .ZN(new_n17200_));
  XOR2_X1    g16180(.A1(new_n16261_), .A2(new_n16269_), .Z(new_n17201_));
  NAND2_X1   g16181(.A1(new_n16253_), .A2(new_n17201_), .ZN(new_n17202_));
  OAI21_X1   g16182(.A1(new_n16573_), .A2(new_n16574_), .B(new_n16570_), .ZN(new_n17203_));
  NAND4_X1   g16183(.A1(new_n17203_), .A2(new_n17198_), .A3(new_n17200_), .A4(new_n17202_), .ZN(new_n17204_));
  INV_X1     g16184(.I(new_n16587_), .ZN(new_n17205_));
  AND2_X2    g16185(.A1(new_n16588_), .A2(new_n16589_), .Z(new_n17206_));
  OAI22_X1   g16186(.A1(new_n16585_), .A2(new_n17205_), .B1(new_n17206_), .B2(new_n16578_), .ZN(new_n17207_));
  AOI22_X1   g16187(.A1(new_n17203_), .A2(new_n17202_), .B1(new_n17198_), .B2(new_n17200_), .ZN(new_n17208_));
  OAI21_X1   g16188(.A1(new_n17207_), .A2(new_n17208_), .B(new_n17204_), .ZN(new_n17209_));
  AOI21_X1   g16189(.A1(new_n16599_), .A2(new_n16600_), .B(new_n16543_), .ZN(new_n17210_));
  NOR3_X1    g16190(.A1(new_n16597_), .A2(new_n16594_), .A3(new_n16542_), .ZN(new_n17211_));
  NOR2_X1    g16191(.A1(new_n17211_), .A2(new_n17210_), .ZN(new_n17212_));
  NOR2_X1    g16192(.A1(new_n17212_), .A2(new_n16611_), .ZN(new_n17213_));
  AOI21_X1   g16193(.A1(new_n16608_), .A2(new_n16609_), .B(new_n16282_), .ZN(new_n17214_));
  NOR3_X1    g16194(.A1(new_n16605_), .A2(new_n16606_), .A3(new_n16278_), .ZN(new_n17215_));
  NOR2_X1    g16195(.A1(new_n17215_), .A2(new_n17214_), .ZN(new_n17216_));
  NOR2_X1    g16196(.A1(new_n16602_), .A2(new_n17216_), .ZN(new_n17217_));
  OAI21_X1   g16197(.A1(new_n17213_), .A2(new_n17217_), .B(new_n17209_), .ZN(new_n17218_));
  NOR2_X1    g16198(.A1(new_n16602_), .A2(new_n16611_), .ZN(new_n17219_));
  AOI22_X1   g16199(.A1(new_n16598_), .A2(new_n16601_), .B1(new_n16607_), .B2(new_n16610_), .ZN(new_n17220_));
  OAI21_X1   g16200(.A1(new_n17219_), .A2(new_n17220_), .B(new_n16593_), .ZN(new_n17221_));
  XOR2_X1    g16201(.A1(new_n17088_), .A2(new_n17098_), .Z(new_n17222_));
  NAND2_X1   g16202(.A1(new_n17134_), .A2(new_n17222_), .ZN(new_n17223_));
  NAND2_X1   g16203(.A1(new_n17105_), .A2(new_n17099_), .ZN(new_n17224_));
  NAND2_X1   g16204(.A1(new_n17123_), .A2(new_n17224_), .ZN(new_n17225_));
  XOR2_X1    g16205(.A1(new_n16848_), .A2(new_n16840_), .Z(new_n17226_));
  NAND2_X1   g16206(.A1(new_n16831_), .A2(new_n17226_), .ZN(new_n17227_));
  OAI21_X1   g16207(.A1(new_n17147_), .A2(new_n17148_), .B(new_n17144_), .ZN(new_n17228_));
  NAND4_X1   g16208(.A1(new_n17228_), .A2(new_n17225_), .A3(new_n17223_), .A4(new_n17227_), .ZN(new_n17229_));
  INV_X1     g16209(.I(new_n17162_), .ZN(new_n17230_));
  NOR2_X1    g16210(.A1(new_n17164_), .A2(new_n17163_), .ZN(new_n17231_));
  OAI22_X1   g16211(.A1(new_n17230_), .A2(new_n17160_), .B1(new_n17231_), .B2(new_n17152_), .ZN(new_n17232_));
  AOI22_X1   g16212(.A1(new_n17228_), .A2(new_n17227_), .B1(new_n17225_), .B2(new_n17223_), .ZN(new_n17233_));
  OAI21_X1   g16213(.A1(new_n17233_), .A2(new_n17232_), .B(new_n17229_), .ZN(new_n17234_));
  AOI21_X1   g16214(.A1(new_n17173_), .A2(new_n17174_), .B(new_n17116_), .ZN(new_n17235_));
  NOR3_X1    g16215(.A1(new_n17169_), .A2(new_n17115_), .A3(new_n17170_), .ZN(new_n17236_));
  NOR2_X1    g16216(.A1(new_n17236_), .A2(new_n17235_), .ZN(new_n17237_));
  NAND2_X1   g16217(.A1(new_n17181_), .A2(new_n17185_), .ZN(new_n17238_));
  NOR2_X1    g16218(.A1(new_n17237_), .A2(new_n17238_), .ZN(new_n17239_));
  NAND2_X1   g16219(.A1(new_n17171_), .A2(new_n17175_), .ZN(new_n17240_));
  AOI21_X1   g16220(.A1(new_n17183_), .A2(new_n17184_), .B(new_n17182_), .ZN(new_n17241_));
  NOR3_X1    g16221(.A1(new_n17179_), .A2(new_n17180_), .A3(new_n16857_), .ZN(new_n17242_));
  NOR2_X1    g16222(.A1(new_n17242_), .A2(new_n17241_), .ZN(new_n17243_));
  NOR2_X1    g16223(.A1(new_n17240_), .A2(new_n17243_), .ZN(new_n17244_));
  OAI21_X1   g16224(.A1(new_n17239_), .A2(new_n17244_), .B(new_n17234_), .ZN(new_n17245_));
  NOR2_X1    g16225(.A1(new_n17240_), .A2(new_n17238_), .ZN(new_n17246_));
  AOI22_X1   g16226(.A1(new_n17171_), .A2(new_n17175_), .B1(new_n17181_), .B2(new_n17185_), .ZN(new_n17247_));
  OAI21_X1   g16227(.A1(new_n17246_), .A2(new_n17247_), .B(new_n17168_), .ZN(new_n17248_));
  NAND4_X1   g16228(.A1(new_n17245_), .A2(new_n17248_), .A3(new_n17218_), .A4(new_n17221_), .ZN(new_n17249_));
  NOR2_X1    g16229(.A1(new_n17135_), .A2(new_n17125_), .ZN(new_n17250_));
  NAND2_X1   g16230(.A1(new_n17228_), .A2(new_n17227_), .ZN(new_n17251_));
  NAND2_X1   g16231(.A1(new_n17250_), .A2(new_n17251_), .ZN(new_n17252_));
  NAND2_X1   g16232(.A1(new_n17225_), .A2(new_n17223_), .ZN(new_n17253_));
  NOR2_X1    g16233(.A1(new_n17150_), .A2(new_n17146_), .ZN(new_n17254_));
  NAND2_X1   g16234(.A1(new_n17253_), .A2(new_n17254_), .ZN(new_n17255_));
  AOI21_X1   g16235(.A1(new_n17252_), .A2(new_n17255_), .B(new_n17232_), .ZN(new_n17256_));
  AOI21_X1   g16236(.A1(new_n17229_), .A2(new_n17167_), .B(new_n17166_), .ZN(new_n17257_));
  NOR2_X1    g16237(.A1(new_n16562_), .A2(new_n16551_), .ZN(new_n17258_));
  NAND2_X1   g16238(.A1(new_n17203_), .A2(new_n17202_), .ZN(new_n17259_));
  NAND2_X1   g16239(.A1(new_n17259_), .A2(new_n17258_), .ZN(new_n17260_));
  NAND2_X1   g16240(.A1(new_n17198_), .A2(new_n17200_), .ZN(new_n17261_));
  NOR2_X1    g16241(.A1(new_n16572_), .A2(new_n16576_), .ZN(new_n17262_));
  NAND2_X1   g16242(.A1(new_n17262_), .A2(new_n17261_), .ZN(new_n17263_));
  AOI21_X1   g16243(.A1(new_n17260_), .A2(new_n17263_), .B(new_n17207_), .ZN(new_n17264_));
  AOI21_X1   g16244(.A1(new_n17204_), .A2(new_n16592_), .B(new_n16591_), .ZN(new_n17265_));
  NOR4_X1    g16245(.A1(new_n17256_), .A2(new_n17257_), .A3(new_n17264_), .A4(new_n17265_), .ZN(new_n17266_));
  NOR3_X1    g16246(.A1(new_n17205_), .A2(new_n16585_), .A3(new_n16590_), .ZN(new_n17267_));
  INV_X1     g16247(.I(new_n17267_), .ZN(new_n17268_));
  INV_X1     g16248(.I(new_n17159_), .ZN(new_n17269_));
  NAND2_X1   g16249(.A1(new_n17158_), .A2(new_n17155_), .ZN(new_n17270_));
  NAND2_X1   g16250(.A1(new_n17269_), .A2(new_n17270_), .ZN(new_n17271_));
  INV_X1     g16251(.I(new_n17271_), .ZN(new_n17272_));
  NOR2_X1    g16252(.A1(new_n16582_), .A2(new_n16581_), .ZN(new_n17273_));
  NOR2_X1    g16253(.A1(new_n16584_), .A2(new_n17273_), .ZN(new_n17274_));
  NAND2_X1   g16254(.A1(new_n17272_), .A2(new_n17274_), .ZN(new_n17275_));
  NAND2_X1   g16255(.A1(new_n17268_), .A2(new_n17275_), .ZN(new_n17276_));
  INV_X1     g16256(.I(new_n17275_), .ZN(new_n17277_));
  NAND2_X1   g16257(.A1(new_n17277_), .A2(new_n17267_), .ZN(new_n17278_));
  OAI21_X1   g16258(.A1(new_n17230_), .A2(new_n17160_), .B(new_n17231_), .ZN(new_n17279_));
  NAND3_X1   g16259(.A1(new_n17165_), .A2(new_n17161_), .A3(new_n17162_), .ZN(new_n17280_));
  NAND2_X1   g16260(.A1(new_n17280_), .A2(new_n17279_), .ZN(new_n17281_));
  AOI22_X1   g16261(.A1(new_n17276_), .A2(new_n17278_), .B1(new_n17281_), .B2(new_n17268_), .ZN(new_n17282_));
  OAI22_X1   g16262(.A1(new_n17256_), .A2(new_n17257_), .B1(new_n17264_), .B2(new_n17265_), .ZN(new_n17283_));
  AOI21_X1   g16263(.A1(new_n17283_), .A2(new_n17282_), .B(new_n17266_), .ZN(new_n17284_));
  AOI22_X1   g16264(.A1(new_n17245_), .A2(new_n17248_), .B1(new_n17218_), .B2(new_n17221_), .ZN(new_n17285_));
  OAI21_X1   g16265(.A1(new_n17285_), .A2(new_n17284_), .B(new_n17249_), .ZN(new_n17286_));
  AOI21_X1   g16266(.A1(new_n17212_), .A2(new_n17216_), .B(new_n17209_), .ZN(new_n17287_));
  INV_X1     g16267(.I(new_n16615_), .ZN(new_n17288_));
  OAI21_X1   g16268(.A1(new_n17287_), .A2(new_n17288_), .B(new_n16548_), .ZN(new_n17289_));
  NAND3_X1   g16269(.A1(new_n16612_), .A2(new_n16547_), .A3(new_n16615_), .ZN(new_n17290_));
  AOI21_X1   g16270(.A1(new_n17289_), .A2(new_n17290_), .B(new_n16284_), .ZN(new_n17291_));
  AOI21_X1   g16271(.A1(new_n16612_), .A2(new_n16615_), .B(new_n16547_), .ZN(new_n17292_));
  NOR3_X1    g16272(.A1(new_n17287_), .A2(new_n16548_), .A3(new_n17288_), .ZN(new_n17293_));
  NOR3_X1    g16273(.A1(new_n17293_), .A2(new_n17292_), .A3(new_n16285_), .ZN(new_n17294_));
  INV_X1     g16274(.I(new_n16860_), .ZN(new_n17295_));
  AOI21_X1   g16275(.A1(new_n17237_), .A2(new_n17243_), .B(new_n17234_), .ZN(new_n17296_));
  INV_X1     g16276(.I(new_n17190_), .ZN(new_n17297_));
  OAI21_X1   g16277(.A1(new_n17296_), .A2(new_n17297_), .B(new_n17121_), .ZN(new_n17298_));
  NAND3_X1   g16278(.A1(new_n17187_), .A2(new_n17120_), .A3(new_n17190_), .ZN(new_n17299_));
  AOI21_X1   g16279(.A1(new_n17299_), .A2(new_n17298_), .B(new_n17295_), .ZN(new_n17300_));
  AOI21_X1   g16280(.A1(new_n17187_), .A2(new_n17190_), .B(new_n17120_), .ZN(new_n17301_));
  NOR3_X1    g16281(.A1(new_n17296_), .A2(new_n17121_), .A3(new_n17297_), .ZN(new_n17302_));
  NOR3_X1    g16282(.A1(new_n17301_), .A2(new_n17302_), .A3(new_n16860_), .ZN(new_n17303_));
  NOR4_X1    g16283(.A1(new_n17300_), .A2(new_n17303_), .A3(new_n17294_), .A4(new_n17291_), .ZN(new_n17304_));
  XOR2_X1    g16284(.A1(new_n16284_), .A2(new_n16547_), .Z(new_n17305_));
  XNOR2_X1   g16285(.A1(new_n17120_), .A2(new_n16860_), .ZN(new_n17306_));
  NOR4_X1    g16286(.A1(new_n17191_), .A2(new_n16616_), .A3(new_n17305_), .A4(new_n17306_), .ZN(new_n17307_));
  OAI21_X1   g16287(.A1(new_n17304_), .A2(new_n17286_), .B(new_n17307_), .ZN(new_n17308_));
  INV_X1     g16288(.I(new_n17308_), .ZN(new_n17309_));
  NAND4_X1   g16289(.A1(new_n17194_), .A2(new_n16618_), .A3(new_n16549_), .A4(new_n17122_), .ZN(new_n17310_));
  NOR2_X1    g16290(.A1(new_n17309_), .A2(new_n17310_), .ZN(new_n17311_));
  NOR2_X1    g16291(.A1(new_n17311_), .A2(new_n17196_), .ZN(new_n17312_));
  INV_X1     g16292(.I(new_n17312_), .ZN(new_n17313_));
  NOR2_X1    g16293(.A1(new_n17313_), .A2(new_n16019_), .ZN(new_n17314_));
  NOR2_X1    g16294(.A1(new_n16009_), .A2(new_n16006_), .ZN(new_n17315_));
  NOR2_X1    g16295(.A1(new_n15996_), .A2(new_n15999_), .ZN(new_n17316_));
  NAND2_X1   g16296(.A1(new_n15991_), .A2(new_n17316_), .ZN(new_n17317_));
  NAND2_X1   g16297(.A1(new_n15924_), .A2(new_n15927_), .ZN(new_n17318_));
  NAND2_X1   g16298(.A1(new_n15921_), .A2(new_n15922_), .ZN(new_n17319_));
  AOI21_X1   g16299(.A1(new_n17318_), .A2(new_n17319_), .B(new_n15306_), .ZN(new_n17320_));
  NAND2_X1   g16300(.A1(new_n15924_), .A2(new_n15922_), .ZN(new_n17321_));
  AOI21_X1   g16301(.A1(new_n17321_), .A2(new_n15321_), .B(new_n15918_), .ZN(new_n17322_));
  NOR2_X1    g16302(.A1(new_n17320_), .A2(new_n17322_), .ZN(new_n17323_));
  NAND2_X1   g16303(.A1(new_n15892_), .A2(new_n15954_), .ZN(new_n17324_));
  NAND2_X1   g16304(.A1(new_n15950_), .A2(new_n15903_), .ZN(new_n17325_));
  AOI21_X1   g16305(.A1(new_n17324_), .A2(new_n17325_), .B(new_n15881_), .ZN(new_n17326_));
  NAND2_X1   g16306(.A1(new_n15950_), .A2(new_n15954_), .ZN(new_n17327_));
  NAND2_X1   g16307(.A1(new_n15892_), .A2(new_n15903_), .ZN(new_n17328_));
  AOI21_X1   g16308(.A1(new_n17327_), .A2(new_n17328_), .B(new_n15947_), .ZN(new_n17329_));
  NOR2_X1    g16309(.A1(new_n17326_), .A2(new_n17329_), .ZN(new_n17330_));
  AOI21_X1   g16310(.A1(new_n15938_), .A2(new_n15941_), .B(new_n15964_), .ZN(new_n17331_));
  NOR2_X1    g16311(.A1(new_n15961_), .A2(new_n15962_), .ZN(new_n17332_));
  OAI21_X1   g16312(.A1(new_n17331_), .A2(new_n17332_), .B(new_n15879_), .ZN(new_n17333_));
  OAI21_X1   g16313(.A1(new_n15864_), .A2(new_n15946_), .B(new_n15945_), .ZN(new_n17334_));
  NOR2_X1    g16314(.A1(new_n15970_), .A2(new_n15304_), .ZN(new_n17335_));
  NOR2_X1    g16315(.A1(new_n15968_), .A2(new_n15284_), .ZN(new_n17336_));
  OAI21_X1   g16316(.A1(new_n17335_), .A2(new_n17336_), .B(new_n15299_), .ZN(new_n17337_));
  OAI21_X1   g16317(.A1(new_n15285_), .A2(new_n15917_), .B(new_n15916_), .ZN(new_n17338_));
  NAND4_X1   g16318(.A1(new_n17333_), .A2(new_n17337_), .A3(new_n17338_), .A4(new_n17334_), .ZN(new_n17339_));
  INV_X1     g16319(.I(new_n15983_), .ZN(new_n17340_));
  INV_X1     g16320(.I(new_n15986_), .ZN(new_n17341_));
  OAI22_X1   g16321(.A1(new_n17341_), .A2(new_n15975_), .B1(new_n17340_), .B2(new_n15981_), .ZN(new_n17342_));
  AOI22_X1   g16322(.A1(new_n17333_), .A2(new_n17334_), .B1(new_n17337_), .B2(new_n17338_), .ZN(new_n17343_));
  OAI21_X1   g16323(.A1(new_n17343_), .A2(new_n17342_), .B(new_n17339_), .ZN(new_n17344_));
  OAI21_X1   g16324(.A1(new_n17330_), .A2(new_n17323_), .B(new_n17344_), .ZN(new_n17345_));
  OAI21_X1   g16325(.A1(new_n15997_), .A2(new_n15998_), .B(new_n14993_), .ZN(new_n17346_));
  NAND3_X1   g16326(.A1(new_n15995_), .A2(new_n15994_), .A3(new_n14992_), .ZN(new_n17347_));
  NAND2_X1   g16327(.A1(new_n17346_), .A2(new_n17347_), .ZN(new_n17348_));
  NAND3_X1   g16328(.A1(new_n17348_), .A2(new_n17345_), .A3(new_n15960_), .ZN(new_n17349_));
  AOI21_X1   g16329(.A1(new_n17317_), .A2(new_n17349_), .B(new_n17315_), .ZN(new_n17350_));
  INV_X1     g16330(.I(new_n17315_), .ZN(new_n17351_));
  NAND2_X1   g16331(.A1(new_n15991_), .A2(new_n17348_), .ZN(new_n17352_));
  NAND3_X1   g16332(.A1(new_n17316_), .A2(new_n17345_), .A3(new_n15960_), .ZN(new_n17353_));
  AOI21_X1   g16333(.A1(new_n17352_), .A2(new_n17353_), .B(new_n17351_), .ZN(new_n17354_));
  NOR2_X1    g16334(.A1(new_n17354_), .A2(new_n17350_), .ZN(new_n17355_));
  NAND2_X1   g16335(.A1(new_n15929_), .A2(new_n15932_), .ZN(new_n17356_));
  NOR2_X1    g16336(.A1(new_n17330_), .A2(new_n17356_), .ZN(new_n17357_));
  NAND2_X1   g16337(.A1(new_n15956_), .A2(new_n15959_), .ZN(new_n17358_));
  NOR2_X1    g16338(.A1(new_n17323_), .A2(new_n17358_), .ZN(new_n17359_));
  OAI21_X1   g16339(.A1(new_n17357_), .A2(new_n17359_), .B(new_n17344_), .ZN(new_n17360_));
  NOR2_X1    g16340(.A1(new_n17356_), .A2(new_n17358_), .ZN(new_n17361_));
  OAI21_X1   g16341(.A1(new_n17361_), .A2(new_n15990_), .B(new_n15989_), .ZN(new_n17362_));
  NOR2_X1    g16342(.A1(new_n17253_), .A2(new_n17254_), .ZN(new_n17363_));
  NOR2_X1    g16343(.A1(new_n17250_), .A2(new_n17251_), .ZN(new_n17364_));
  OAI21_X1   g16344(.A1(new_n17364_), .A2(new_n17363_), .B(new_n17166_), .ZN(new_n17365_));
  OAI21_X1   g16345(.A1(new_n17233_), .A2(new_n17151_), .B(new_n17232_), .ZN(new_n17366_));
  NOR2_X1    g16346(.A1(new_n17262_), .A2(new_n17261_), .ZN(new_n17367_));
  NOR2_X1    g16347(.A1(new_n17259_), .A2(new_n17258_), .ZN(new_n17368_));
  OAI21_X1   g16348(.A1(new_n17368_), .A2(new_n17367_), .B(new_n16591_), .ZN(new_n17369_));
  OAI21_X1   g16349(.A1(new_n16577_), .A2(new_n17208_), .B(new_n17207_), .ZN(new_n17370_));
  NAND4_X1   g16350(.A1(new_n17365_), .A2(new_n17369_), .A3(new_n17370_), .A4(new_n17366_), .ZN(new_n17371_));
  NOR2_X1    g16351(.A1(new_n17277_), .A2(new_n17267_), .ZN(new_n17372_));
  NOR2_X1    g16352(.A1(new_n17268_), .A2(new_n17275_), .ZN(new_n17373_));
  INV_X1     g16353(.I(new_n17281_), .ZN(new_n17374_));
  OAI22_X1   g16354(.A1(new_n17374_), .A2(new_n17267_), .B1(new_n17373_), .B2(new_n17372_), .ZN(new_n17375_));
  AOI22_X1   g16355(.A1(new_n17365_), .A2(new_n17366_), .B1(new_n17369_), .B2(new_n17370_), .ZN(new_n17376_));
  OAI21_X1   g16356(.A1(new_n17376_), .A2(new_n17375_), .B(new_n17371_), .ZN(new_n17377_));
  NAND2_X1   g16357(.A1(new_n17218_), .A2(new_n17221_), .ZN(new_n17378_));
  NAND2_X1   g16358(.A1(new_n17240_), .A2(new_n17243_), .ZN(new_n17379_));
  NAND2_X1   g16359(.A1(new_n17237_), .A2(new_n17238_), .ZN(new_n17380_));
  AOI21_X1   g16360(.A1(new_n17380_), .A2(new_n17379_), .B(new_n17168_), .ZN(new_n17381_));
  OAI22_X1   g16361(.A1(new_n17236_), .A2(new_n17235_), .B1(new_n17242_), .B2(new_n17241_), .ZN(new_n17382_));
  AOI21_X1   g16362(.A1(new_n17382_), .A2(new_n17186_), .B(new_n17234_), .ZN(new_n17383_));
  NOR2_X1    g16363(.A1(new_n17381_), .A2(new_n17383_), .ZN(new_n17384_));
  NOR2_X1    g16364(.A1(new_n17384_), .A2(new_n17378_), .ZN(new_n17385_));
  NAND2_X1   g16365(.A1(new_n16602_), .A2(new_n17216_), .ZN(new_n17386_));
  NAND2_X1   g16366(.A1(new_n17212_), .A2(new_n16611_), .ZN(new_n17387_));
  AOI21_X1   g16367(.A1(new_n17387_), .A2(new_n17386_), .B(new_n16593_), .ZN(new_n17388_));
  NAND4_X1   g16368(.A1(new_n16598_), .A2(new_n16601_), .A3(new_n16607_), .A4(new_n16610_), .ZN(new_n17389_));
  NAND2_X1   g16369(.A1(new_n16602_), .A2(new_n16611_), .ZN(new_n17390_));
  AOI21_X1   g16370(.A1(new_n17390_), .A2(new_n17389_), .B(new_n17209_), .ZN(new_n17391_));
  NOR2_X1    g16371(.A1(new_n17388_), .A2(new_n17391_), .ZN(new_n17392_));
  NAND2_X1   g16372(.A1(new_n17245_), .A2(new_n17248_), .ZN(new_n17393_));
  NOR2_X1    g16373(.A1(new_n17393_), .A2(new_n17392_), .ZN(new_n17394_));
  OAI21_X1   g16374(.A1(new_n17394_), .A2(new_n17385_), .B(new_n17377_), .ZN(new_n17395_));
  NOR4_X1    g16375(.A1(new_n17381_), .A2(new_n17388_), .A3(new_n17391_), .A4(new_n17383_), .ZN(new_n17396_));
  OAI21_X1   g16376(.A1(new_n17285_), .A2(new_n17396_), .B(new_n17284_), .ZN(new_n17397_));
  NAND4_X1   g16377(.A1(new_n17395_), .A2(new_n17360_), .A3(new_n17362_), .A4(new_n17397_), .ZN(new_n17398_));
  NAND2_X1   g16378(.A1(new_n17365_), .A2(new_n17366_), .ZN(new_n17399_));
  NOR2_X1    g16379(.A1(new_n17264_), .A2(new_n17265_), .ZN(new_n17400_));
  NOR2_X1    g16380(.A1(new_n17399_), .A2(new_n17400_), .ZN(new_n17401_));
  NOR2_X1    g16381(.A1(new_n17256_), .A2(new_n17257_), .ZN(new_n17402_));
  NAND2_X1   g16382(.A1(new_n17369_), .A2(new_n17370_), .ZN(new_n17403_));
  NOR2_X1    g16383(.A1(new_n17402_), .A2(new_n17403_), .ZN(new_n17404_));
  OAI21_X1   g16384(.A1(new_n17404_), .A2(new_n17401_), .B(new_n17282_), .ZN(new_n17405_));
  AOI21_X1   g16385(.A1(new_n17283_), .A2(new_n17371_), .B(new_n17282_), .ZN(new_n17406_));
  INV_X1     g16386(.I(new_n17406_), .ZN(new_n17407_));
  NAND2_X1   g16387(.A1(new_n17407_), .A2(new_n17405_), .ZN(new_n17408_));
  NAND2_X1   g16388(.A1(new_n17333_), .A2(new_n17334_), .ZN(new_n17409_));
  NOR2_X1    g16389(.A1(new_n15972_), .A2(new_n15973_), .ZN(new_n17410_));
  NOR2_X1    g16390(.A1(new_n17409_), .A2(new_n17410_), .ZN(new_n17411_));
  NOR2_X1    g16391(.A1(new_n15966_), .A2(new_n15967_), .ZN(new_n17412_));
  NAND2_X1   g16392(.A1(new_n17337_), .A2(new_n17338_), .ZN(new_n17413_));
  NOR2_X1    g16393(.A1(new_n17413_), .A2(new_n17412_), .ZN(new_n17414_));
  OAI21_X1   g16394(.A1(new_n17411_), .A2(new_n17414_), .B(new_n15987_), .ZN(new_n17415_));
  OAI21_X1   g16395(.A1(new_n17343_), .A2(new_n15974_), .B(new_n17342_), .ZN(new_n17416_));
  NAND2_X1   g16396(.A1(new_n17415_), .A2(new_n17416_), .ZN(new_n17417_));
  NOR2_X1    g16397(.A1(new_n17408_), .A2(new_n17417_), .ZN(new_n17418_));
  NOR2_X1    g16398(.A1(new_n17340_), .A2(new_n15981_), .ZN(new_n17419_));
  NAND2_X1   g16399(.A1(new_n17419_), .A2(new_n17341_), .ZN(new_n17420_));
  NOR2_X1    g16400(.A1(new_n17272_), .A2(new_n17274_), .ZN(new_n17421_));
  NOR2_X1    g16401(.A1(new_n17277_), .A2(new_n17421_), .ZN(new_n17422_));
  NOR2_X1    g16402(.A1(new_n15978_), .A2(new_n15977_), .ZN(new_n17423_));
  NOR2_X1    g16403(.A1(new_n15980_), .A2(new_n17423_), .ZN(new_n17424_));
  NAND2_X1   g16404(.A1(new_n17422_), .A2(new_n17424_), .ZN(new_n17425_));
  NAND2_X1   g16405(.A1(new_n17420_), .A2(new_n17425_), .ZN(new_n17426_));
  NAND4_X1   g16406(.A1(new_n17419_), .A2(new_n17341_), .A3(new_n17422_), .A4(new_n17424_), .ZN(new_n17427_));
  AOI21_X1   g16407(.A1(new_n17276_), .A2(new_n17278_), .B(new_n17281_), .ZN(new_n17428_));
  NOR3_X1    g16408(.A1(new_n17374_), .A2(new_n17372_), .A3(new_n17373_), .ZN(new_n17429_));
  NOR2_X1    g16409(.A1(new_n17429_), .A2(new_n17428_), .ZN(new_n17430_));
  INV_X1     g16410(.I(new_n17430_), .ZN(new_n17431_));
  AOI22_X1   g16411(.A1(new_n17431_), .A2(new_n17420_), .B1(new_n17426_), .B2(new_n17427_), .ZN(new_n17432_));
  AOI22_X1   g16412(.A1(new_n17407_), .A2(new_n17405_), .B1(new_n17415_), .B2(new_n17416_), .ZN(new_n17433_));
  INV_X1     g16413(.I(new_n17433_), .ZN(new_n17434_));
  AOI21_X1   g16414(.A1(new_n17434_), .A2(new_n17432_), .B(new_n17418_), .ZN(new_n17435_));
  AOI22_X1   g16415(.A1(new_n17395_), .A2(new_n17397_), .B1(new_n17360_), .B2(new_n17362_), .ZN(new_n17436_));
  OAI21_X1   g16416(.A1(new_n17436_), .A2(new_n17435_), .B(new_n17398_), .ZN(new_n17437_));
  NAND2_X1   g16417(.A1(new_n17437_), .A2(new_n17355_), .ZN(new_n17438_));
  NOR2_X1    g16418(.A1(new_n17300_), .A2(new_n17303_), .ZN(new_n17439_));
  NOR2_X1    g16419(.A1(new_n17294_), .A2(new_n17291_), .ZN(new_n17440_));
  NAND2_X1   g16420(.A1(new_n17286_), .A2(new_n17440_), .ZN(new_n17441_));
  OAI21_X1   g16421(.A1(new_n17384_), .A2(new_n17392_), .B(new_n17377_), .ZN(new_n17442_));
  OAI21_X1   g16422(.A1(new_n17293_), .A2(new_n17292_), .B(new_n16285_), .ZN(new_n17443_));
  NAND3_X1   g16423(.A1(new_n17289_), .A2(new_n17290_), .A3(new_n16284_), .ZN(new_n17444_));
  NAND2_X1   g16424(.A1(new_n17443_), .A2(new_n17444_), .ZN(new_n17445_));
  NAND3_X1   g16425(.A1(new_n17445_), .A2(new_n17442_), .A3(new_n17249_), .ZN(new_n17446_));
  AOI21_X1   g16426(.A1(new_n17441_), .A2(new_n17446_), .B(new_n17439_), .ZN(new_n17447_));
  INV_X1     g16427(.I(new_n17439_), .ZN(new_n17448_));
  AOI21_X1   g16428(.A1(new_n17393_), .A2(new_n17378_), .B(new_n17284_), .ZN(new_n17449_));
  OAI21_X1   g16429(.A1(new_n17396_), .A2(new_n17449_), .B(new_n17445_), .ZN(new_n17450_));
  NAND3_X1   g16430(.A1(new_n17440_), .A2(new_n17442_), .A3(new_n17249_), .ZN(new_n17451_));
  AOI21_X1   g16431(.A1(new_n17450_), .A2(new_n17451_), .B(new_n17448_), .ZN(new_n17452_));
  NOR2_X1    g16432(.A1(new_n17447_), .A2(new_n17452_), .ZN(new_n17453_));
  OAI21_X1   g16433(.A1(new_n17437_), .A2(new_n17355_), .B(new_n17453_), .ZN(new_n17454_));
  NAND2_X1   g16434(.A1(new_n17454_), .A2(new_n17438_), .ZN(new_n17455_));
  INV_X1     g16435(.I(new_n17195_), .ZN(new_n17456_));
  NAND2_X1   g16436(.A1(new_n17308_), .A2(new_n17456_), .ZN(new_n17457_));
  OAI21_X1   g16437(.A1(new_n17301_), .A2(new_n17302_), .B(new_n16860_), .ZN(new_n17458_));
  NAND3_X1   g16438(.A1(new_n17299_), .A2(new_n17298_), .A3(new_n17295_), .ZN(new_n17459_));
  NAND4_X1   g16439(.A1(new_n17458_), .A2(new_n17459_), .A3(new_n17443_), .A4(new_n17444_), .ZN(new_n17460_));
  NAND3_X1   g16440(.A1(new_n17460_), .A2(new_n17249_), .A3(new_n17442_), .ZN(new_n17461_));
  NAND3_X1   g16441(.A1(new_n17461_), .A2(new_n17195_), .A3(new_n17307_), .ZN(new_n17462_));
  AOI21_X1   g16442(.A1(new_n17457_), .A2(new_n17462_), .B(new_n16619_), .ZN(new_n17463_));
  INV_X1     g16443(.I(new_n16619_), .ZN(new_n17464_));
  AOI21_X1   g16444(.A1(new_n17461_), .A2(new_n17307_), .B(new_n17195_), .ZN(new_n17465_));
  NOR2_X1    g16445(.A1(new_n17308_), .A2(new_n17456_), .ZN(new_n17466_));
  NOR3_X1    g16446(.A1(new_n17466_), .A2(new_n17465_), .A3(new_n17464_), .ZN(new_n17467_));
  INV_X1     g16447(.I(new_n15911_), .ZN(new_n17468_));
  NAND2_X1   g16448(.A1(new_n16014_), .A2(new_n17468_), .ZN(new_n17469_));
  OAI21_X1   g16449(.A1(new_n16008_), .A2(new_n16007_), .B(new_n15578_), .ZN(new_n17470_));
  NAND3_X1   g16450(.A1(new_n16003_), .A2(new_n16005_), .A3(new_n16000_), .ZN(new_n17471_));
  NAND4_X1   g16451(.A1(new_n17346_), .A2(new_n17347_), .A3(new_n17470_), .A4(new_n17471_), .ZN(new_n17472_));
  NAND3_X1   g16452(.A1(new_n17472_), .A2(new_n15960_), .A3(new_n17345_), .ZN(new_n17473_));
  NAND3_X1   g16453(.A1(new_n17473_), .A2(new_n15911_), .A3(new_n16013_), .ZN(new_n17474_));
  AOI21_X1   g16454(.A1(new_n17474_), .A2(new_n17469_), .B(new_n15329_), .ZN(new_n17475_));
  INV_X1     g16455(.I(new_n15329_), .ZN(new_n17476_));
  AOI21_X1   g16456(.A1(new_n17473_), .A2(new_n16013_), .B(new_n15911_), .ZN(new_n17477_));
  NOR2_X1    g16457(.A1(new_n16014_), .A2(new_n17468_), .ZN(new_n17478_));
  NOR3_X1    g16458(.A1(new_n17477_), .A2(new_n17478_), .A3(new_n17476_), .ZN(new_n17479_));
  NOR4_X1    g16459(.A1(new_n17463_), .A2(new_n17467_), .A3(new_n17475_), .A4(new_n17479_), .ZN(new_n17480_));
  XOR2_X1    g16460(.A1(new_n17195_), .A2(new_n16619_), .Z(new_n17481_));
  XOR2_X1    g16461(.A1(new_n15329_), .A2(new_n15911_), .Z(new_n17482_));
  NOR4_X1    g16462(.A1(new_n17481_), .A2(new_n17482_), .A3(new_n17308_), .A4(new_n16014_), .ZN(new_n17483_));
  OAI21_X1   g16463(.A1(new_n17455_), .A2(new_n17480_), .B(new_n17483_), .ZN(new_n17484_));
  NOR4_X1    g16464(.A1(new_n17311_), .A2(new_n16017_), .A3(new_n15912_), .A4(new_n17196_), .ZN(new_n17485_));
  NAND2_X1   g16465(.A1(new_n17484_), .A2(new_n17485_), .ZN(new_n17486_));
  INV_X1     g16466(.I(new_n17486_), .ZN(new_n17487_));
  NOR2_X1    g16467(.A1(new_n14701_), .A2(new_n14693_), .ZN(new_n17488_));
  AOI22_X1   g16468(.A1(new_n14605_), .A2(new_n14608_), .B1(new_n14614_), .B2(new_n14619_), .ZN(new_n17489_));
  OAI21_X1   g16469(.A1(new_n17488_), .A2(new_n17489_), .B(new_n14620_), .ZN(new_n17490_));
  AOI21_X1   g16470(.A1(new_n14711_), .A2(new_n14712_), .B(new_n13846_), .ZN(new_n17491_));
  NOR3_X1    g16471(.A1(new_n14709_), .A2(new_n14707_), .A3(new_n13845_), .ZN(new_n17492_));
  NOR2_X1    g16472(.A1(new_n17492_), .A2(new_n17491_), .ZN(new_n17493_));
  NAND2_X1   g16473(.A1(new_n14719_), .A2(new_n14722_), .ZN(new_n17494_));
  NOR2_X1    g16474(.A1(new_n17493_), .A2(new_n17494_), .ZN(new_n17495_));
  NAND2_X1   g16475(.A1(new_n14710_), .A2(new_n14713_), .ZN(new_n17496_));
  AOI21_X1   g16476(.A1(new_n14720_), .A2(new_n14721_), .B(new_n12503_), .ZN(new_n17497_));
  NOR3_X1    g16477(.A1(new_n14718_), .A2(new_n14717_), .A3(new_n12504_), .ZN(new_n17498_));
  NOR2_X1    g16478(.A1(new_n17498_), .A2(new_n17497_), .ZN(new_n17499_));
  NOR2_X1    g16479(.A1(new_n17496_), .A2(new_n17499_), .ZN(new_n17500_));
  OAI21_X1   g16480(.A1(new_n17495_), .A2(new_n17500_), .B(new_n17490_), .ZN(new_n17501_));
  NAND2_X1   g16481(.A1(new_n14619_), .A2(new_n14614_), .ZN(new_n17502_));
  NOR3_X1    g16482(.A1(new_n17502_), .A2(new_n14623_), .A3(new_n14630_), .ZN(new_n17503_));
  NOR2_X1    g16483(.A1(new_n14668_), .A2(new_n14550_), .ZN(new_n17504_));
  NOR2_X1    g16484(.A1(new_n14666_), .A2(new_n14555_), .ZN(new_n17505_));
  OAI21_X1   g16485(.A1(new_n17504_), .A2(new_n17505_), .B(new_n14545_), .ZN(new_n17506_));
  OAI21_X1   g16486(.A1(new_n14600_), .A2(new_n14531_), .B(new_n14599_), .ZN(new_n17507_));
  NOR2_X1    g16487(.A1(new_n14674_), .A2(new_n13155_), .ZN(new_n17508_));
  NOR2_X1    g16488(.A1(new_n14672_), .A2(new_n14641_), .ZN(new_n17509_));
  OAI21_X1   g16489(.A1(new_n17509_), .A2(new_n17508_), .B(new_n13202_), .ZN(new_n17510_));
  OAI21_X1   g16490(.A1(new_n14647_), .A2(new_n13160_), .B(new_n13201_), .ZN(new_n17511_));
  NAND4_X1   g16491(.A1(new_n17506_), .A2(new_n17510_), .A3(new_n17507_), .A4(new_n17511_), .ZN(new_n17512_));
  AOI22_X1   g16492(.A1(new_n17506_), .A2(new_n17507_), .B1(new_n17510_), .B2(new_n17511_), .ZN(new_n17513_));
  OAI21_X1   g16493(.A1(new_n17513_), .A2(new_n14689_), .B(new_n17512_), .ZN(new_n17514_));
  NAND3_X1   g16494(.A1(new_n17514_), .A2(new_n14663_), .A3(new_n14664_), .ZN(new_n17515_));
  AOI21_X1   g16495(.A1(new_n14663_), .A2(new_n14664_), .B(new_n17514_), .ZN(new_n17516_));
  OAI21_X1   g16496(.A1(new_n17516_), .A2(new_n14700_), .B(new_n17515_), .ZN(new_n17517_));
  OAI21_X1   g16497(.A1(new_n14623_), .A2(new_n14630_), .B(new_n17502_), .ZN(new_n17518_));
  AOI21_X1   g16498(.A1(new_n17518_), .A2(new_n17517_), .B(new_n17503_), .ZN(new_n17519_));
  NOR4_X1    g16499(.A1(new_n17492_), .A2(new_n17491_), .A3(new_n17498_), .A4(new_n17497_), .ZN(new_n17520_));
  NOR2_X1    g16500(.A1(new_n17493_), .A2(new_n17499_), .ZN(new_n17521_));
  OAI21_X1   g16501(.A1(new_n17521_), .A2(new_n17520_), .B(new_n17519_), .ZN(new_n17522_));
  NAND2_X1   g16502(.A1(new_n17501_), .A2(new_n17522_), .ZN(new_n17523_));
  AOI21_X1   g16503(.A1(new_n15960_), .A2(new_n17345_), .B(new_n17348_), .ZN(new_n17524_));
  NOR2_X1    g16504(.A1(new_n15991_), .A2(new_n17316_), .ZN(new_n17525_));
  OAI21_X1   g16505(.A1(new_n17524_), .A2(new_n17525_), .B(new_n17351_), .ZN(new_n17526_));
  AOI22_X1   g16506(.A1(new_n17345_), .A2(new_n15960_), .B1(new_n17346_), .B2(new_n17347_), .ZN(new_n17527_));
  AOI21_X1   g16507(.A1(new_n17356_), .A2(new_n17358_), .B(new_n15989_), .ZN(new_n17528_));
  NOR3_X1    g16508(.A1(new_n17348_), .A2(new_n17528_), .A3(new_n17361_), .ZN(new_n17529_));
  OAI21_X1   g16509(.A1(new_n17527_), .A2(new_n17529_), .B(new_n17315_), .ZN(new_n17530_));
  NAND2_X1   g16510(.A1(new_n17526_), .A2(new_n17530_), .ZN(new_n17531_));
  NAND2_X1   g16511(.A1(new_n17323_), .A2(new_n17358_), .ZN(new_n17532_));
  NAND2_X1   g16512(.A1(new_n17330_), .A2(new_n17356_), .ZN(new_n17533_));
  AOI21_X1   g16513(.A1(new_n17533_), .A2(new_n17532_), .B(new_n15989_), .ZN(new_n17534_));
  NAND2_X1   g16514(.A1(new_n17356_), .A2(new_n17358_), .ZN(new_n17535_));
  AOI21_X1   g16515(.A1(new_n17535_), .A2(new_n15960_), .B(new_n17344_), .ZN(new_n17536_));
  NAND2_X1   g16516(.A1(new_n17393_), .A2(new_n17392_), .ZN(new_n17537_));
  NAND2_X1   g16517(.A1(new_n17384_), .A2(new_n17378_), .ZN(new_n17538_));
  AOI21_X1   g16518(.A1(new_n17537_), .A2(new_n17538_), .B(new_n17284_), .ZN(new_n17539_));
  OAI22_X1   g16519(.A1(new_n17381_), .A2(new_n17383_), .B1(new_n17388_), .B2(new_n17391_), .ZN(new_n17540_));
  AOI21_X1   g16520(.A1(new_n17540_), .A2(new_n17249_), .B(new_n17377_), .ZN(new_n17541_));
  NOR4_X1    g16521(.A1(new_n17539_), .A2(new_n17534_), .A3(new_n17536_), .A4(new_n17541_), .ZN(new_n17542_));
  NAND4_X1   g16522(.A1(new_n17407_), .A2(new_n17415_), .A3(new_n17405_), .A4(new_n17416_), .ZN(new_n17543_));
  INV_X1     g16523(.I(new_n17432_), .ZN(new_n17544_));
  OAI21_X1   g16524(.A1(new_n17433_), .A2(new_n17544_), .B(new_n17543_), .ZN(new_n17545_));
  OAI22_X1   g16525(.A1(new_n17539_), .A2(new_n17541_), .B1(new_n17534_), .B2(new_n17536_), .ZN(new_n17546_));
  AOI21_X1   g16526(.A1(new_n17546_), .A2(new_n17545_), .B(new_n17542_), .ZN(new_n17547_));
  NOR2_X1    g16527(.A1(new_n17547_), .A2(new_n17531_), .ZN(new_n17548_));
  NAND2_X1   g16528(.A1(new_n17547_), .A2(new_n17531_), .ZN(new_n17549_));
  AOI21_X1   g16529(.A1(new_n17453_), .A2(new_n17549_), .B(new_n17548_), .ZN(new_n17550_));
  OAI21_X1   g16530(.A1(new_n17466_), .A2(new_n17465_), .B(new_n17464_), .ZN(new_n17551_));
  NAND3_X1   g16531(.A1(new_n17457_), .A2(new_n17462_), .A3(new_n16619_), .ZN(new_n17552_));
  NAND2_X1   g16532(.A1(new_n17551_), .A2(new_n17552_), .ZN(new_n17553_));
  NOR2_X1    g16533(.A1(new_n17475_), .A2(new_n17479_), .ZN(new_n17554_));
  NAND2_X1   g16534(.A1(new_n17554_), .A2(new_n17553_), .ZN(new_n17555_));
  NOR2_X1    g16535(.A1(new_n17467_), .A2(new_n17463_), .ZN(new_n17556_));
  OAI21_X1   g16536(.A1(new_n17477_), .A2(new_n17478_), .B(new_n17476_), .ZN(new_n17557_));
  NAND3_X1   g16537(.A1(new_n17474_), .A2(new_n17469_), .A3(new_n15329_), .ZN(new_n17558_));
  NAND2_X1   g16538(.A1(new_n17557_), .A2(new_n17558_), .ZN(new_n17559_));
  NAND2_X1   g16539(.A1(new_n17556_), .A2(new_n17559_), .ZN(new_n17560_));
  AOI21_X1   g16540(.A1(new_n17555_), .A2(new_n17560_), .B(new_n17550_), .ZN(new_n17561_));
  NAND4_X1   g16541(.A1(new_n17551_), .A2(new_n17552_), .A3(new_n17557_), .A4(new_n17558_), .ZN(new_n17562_));
  NAND2_X1   g16542(.A1(new_n17553_), .A2(new_n17559_), .ZN(new_n17563_));
  AOI21_X1   g16543(.A1(new_n17563_), .A2(new_n17562_), .B(new_n17455_), .ZN(new_n17564_));
  NOR3_X1    g16544(.A1(new_n17523_), .A2(new_n17561_), .A3(new_n17564_), .ZN(new_n17565_));
  INV_X1     g16545(.I(new_n17453_), .ZN(new_n17566_));
  NOR2_X1    g16546(.A1(new_n17437_), .A2(new_n17355_), .ZN(new_n17567_));
  OAI21_X1   g16547(.A1(new_n17567_), .A2(new_n17548_), .B(new_n17566_), .ZN(new_n17568_));
  NOR2_X1    g16548(.A1(new_n17547_), .A2(new_n17355_), .ZN(new_n17569_));
  NOR2_X1    g16549(.A1(new_n17437_), .A2(new_n17531_), .ZN(new_n17570_));
  OAI21_X1   g16550(.A1(new_n17569_), .A2(new_n17570_), .B(new_n17453_), .ZN(new_n17571_));
  NAND2_X1   g16551(.A1(new_n14631_), .A2(new_n17502_), .ZN(new_n17572_));
  OAI21_X1   g16552(.A1(new_n14623_), .A2(new_n14630_), .B(new_n14660_), .ZN(new_n17573_));
  AOI21_X1   g16553(.A1(new_n17573_), .A2(new_n17572_), .B(new_n17488_), .ZN(new_n17574_));
  AOI21_X1   g16554(.A1(new_n17518_), .A2(new_n14620_), .B(new_n17517_), .ZN(new_n17575_));
  NOR2_X1    g16555(.A1(new_n17574_), .A2(new_n17575_), .ZN(new_n17576_));
  NAND3_X1   g16556(.A1(new_n17576_), .A2(new_n17568_), .A3(new_n17571_), .ZN(new_n17577_));
  NOR2_X1    g16557(.A1(new_n17534_), .A2(new_n17536_), .ZN(new_n17578_));
  NAND2_X1   g16558(.A1(new_n17395_), .A2(new_n17397_), .ZN(new_n17579_));
  NAND2_X1   g16559(.A1(new_n17579_), .A2(new_n17578_), .ZN(new_n17580_));
  NAND2_X1   g16560(.A1(new_n17360_), .A2(new_n17362_), .ZN(new_n17581_));
  NOR2_X1    g16561(.A1(new_n17539_), .A2(new_n17541_), .ZN(new_n17582_));
  NAND2_X1   g16562(.A1(new_n17582_), .A2(new_n17581_), .ZN(new_n17583_));
  AOI21_X1   g16563(.A1(new_n17580_), .A2(new_n17583_), .B(new_n17435_), .ZN(new_n17584_));
  AOI21_X1   g16564(.A1(new_n17546_), .A2(new_n17398_), .B(new_n17545_), .ZN(new_n17585_));
  NAND2_X1   g16565(.A1(new_n17413_), .A2(new_n17412_), .ZN(new_n17586_));
  NAND2_X1   g16566(.A1(new_n17409_), .A2(new_n17410_), .ZN(new_n17587_));
  AOI21_X1   g16567(.A1(new_n17587_), .A2(new_n17586_), .B(new_n17342_), .ZN(new_n17588_));
  AOI21_X1   g16568(.A1(new_n17339_), .A2(new_n15988_), .B(new_n15987_), .ZN(new_n17589_));
  NOR2_X1    g16569(.A1(new_n17588_), .A2(new_n17589_), .ZN(new_n17590_));
  NOR2_X1    g16570(.A1(new_n17408_), .A2(new_n17590_), .ZN(new_n17591_));
  NAND2_X1   g16571(.A1(new_n17402_), .A2(new_n17403_), .ZN(new_n17592_));
  NAND2_X1   g16572(.A1(new_n17399_), .A2(new_n17400_), .ZN(new_n17593_));
  AOI21_X1   g16573(.A1(new_n17592_), .A2(new_n17593_), .B(new_n17375_), .ZN(new_n17594_));
  NOR2_X1    g16574(.A1(new_n17594_), .A2(new_n17406_), .ZN(new_n17595_));
  NOR2_X1    g16575(.A1(new_n17417_), .A2(new_n17595_), .ZN(new_n17596_));
  OAI21_X1   g16576(.A1(new_n17591_), .A2(new_n17596_), .B(new_n17432_), .ZN(new_n17597_));
  AOI21_X1   g16577(.A1(new_n17434_), .A2(new_n17543_), .B(new_n17432_), .ZN(new_n17598_));
  INV_X1     g16578(.I(new_n17598_), .ZN(new_n17599_));
  NOR2_X1    g16579(.A1(new_n14670_), .A2(new_n14671_), .ZN(new_n17600_));
  NAND2_X1   g16580(.A1(new_n17510_), .A2(new_n17511_), .ZN(new_n17601_));
  NAND2_X1   g16581(.A1(new_n17600_), .A2(new_n17601_), .ZN(new_n17602_));
  NOR2_X1    g16582(.A1(new_n14677_), .A2(new_n14676_), .ZN(new_n17603_));
  OAI21_X1   g16583(.A1(new_n14670_), .A2(new_n14671_), .B(new_n17603_), .ZN(new_n17604_));
  AOI21_X1   g16584(.A1(new_n17604_), .A2(new_n17602_), .B(new_n14689_), .ZN(new_n17605_));
  AOI21_X1   g16585(.A1(new_n14691_), .A2(new_n17512_), .B(new_n14690_), .ZN(new_n17606_));
  NOR2_X1    g16586(.A1(new_n17605_), .A2(new_n17606_), .ZN(new_n17607_));
  NAND3_X1   g16587(.A1(new_n17599_), .A2(new_n17607_), .A3(new_n17597_), .ZN(new_n17608_));
  NOR3_X1    g16588(.A1(new_n17608_), .A2(new_n17584_), .A3(new_n17585_), .ZN(new_n17609_));
  INV_X1     g16589(.I(new_n14700_), .ZN(new_n17610_));
  OAI21_X1   g16590(.A1(new_n14693_), .A2(new_n17516_), .B(new_n14700_), .ZN(new_n17611_));
  INV_X1     g16591(.I(new_n17611_), .ZN(new_n17612_));
  XOR2_X1    g16592(.A1(new_n14665_), .A2(new_n14692_), .Z(new_n17613_));
  AOI21_X1   g16593(.A1(new_n17610_), .A2(new_n17613_), .B(new_n17612_), .ZN(new_n17614_));
  OAI21_X1   g16594(.A1(new_n17584_), .A2(new_n17585_), .B(new_n17608_), .ZN(new_n17615_));
  AOI21_X1   g16595(.A1(new_n17614_), .A2(new_n17615_), .B(new_n17609_), .ZN(new_n17616_));
  NOR3_X1    g16596(.A1(new_n14660_), .A2(new_n14623_), .A3(new_n14630_), .ZN(new_n17617_));
  NOR2_X1    g16597(.A1(new_n14631_), .A2(new_n17502_), .ZN(new_n17618_));
  OAI21_X1   g16598(.A1(new_n17618_), .A2(new_n17617_), .B(new_n17517_), .ZN(new_n17619_));
  OAI21_X1   g16599(.A1(new_n17503_), .A2(new_n17489_), .B(new_n17488_), .ZN(new_n17620_));
  AOI22_X1   g16600(.A1(new_n17568_), .A2(new_n17571_), .B1(new_n17619_), .B2(new_n17620_), .ZN(new_n17621_));
  OAI21_X1   g16601(.A1(new_n17621_), .A2(new_n17616_), .B(new_n17577_), .ZN(new_n17622_));
  OAI21_X1   g16602(.A1(new_n17561_), .A2(new_n17564_), .B(new_n17523_), .ZN(new_n17623_));
  AOI21_X1   g16603(.A1(new_n17623_), .A2(new_n17622_), .B(new_n17565_), .ZN(new_n17624_));
  INV_X1     g16604(.I(new_n13231_), .ZN(new_n17625_));
  AOI21_X1   g16605(.A1(new_n14724_), .A2(new_n14728_), .B(new_n14579_), .ZN(new_n17626_));
  INV_X1     g16606(.I(new_n14579_), .ZN(new_n17627_));
  OAI21_X1   g16607(.A1(new_n17490_), .A2(new_n17520_), .B(new_n14728_), .ZN(new_n17628_));
  NOR2_X1    g16608(.A1(new_n17628_), .A2(new_n17627_), .ZN(new_n17629_));
  OAI21_X1   g16609(.A1(new_n17629_), .A2(new_n17626_), .B(new_n17625_), .ZN(new_n17630_));
  NAND2_X1   g16610(.A1(new_n17628_), .A2(new_n17627_), .ZN(new_n17631_));
  NAND3_X1   g16611(.A1(new_n14724_), .A2(new_n14579_), .A3(new_n14728_), .ZN(new_n17632_));
  NAND3_X1   g16612(.A1(new_n17631_), .A2(new_n17632_), .A3(new_n13231_), .ZN(new_n17633_));
  NAND3_X1   g16613(.A1(new_n17562_), .A2(new_n17438_), .A3(new_n17454_), .ZN(new_n17634_));
  AOI21_X1   g16614(.A1(new_n17634_), .A2(new_n17483_), .B(new_n17313_), .ZN(new_n17635_));
  NOR2_X1    g16615(.A1(new_n17484_), .A2(new_n17312_), .ZN(new_n17636_));
  OAI21_X1   g16616(.A1(new_n17636_), .A2(new_n17635_), .B(new_n16018_), .ZN(new_n17637_));
  NAND2_X1   g16617(.A1(new_n17484_), .A2(new_n17312_), .ZN(new_n17638_));
  NAND3_X1   g16618(.A1(new_n17634_), .A2(new_n17313_), .A3(new_n17483_), .ZN(new_n17639_));
  NAND3_X1   g16619(.A1(new_n17638_), .A2(new_n17639_), .A3(new_n16019_), .ZN(new_n17640_));
  NAND4_X1   g16620(.A1(new_n17637_), .A2(new_n17640_), .A3(new_n17630_), .A4(new_n17633_), .ZN(new_n17641_));
  NAND2_X1   g16621(.A1(new_n17641_), .A2(new_n17624_), .ZN(new_n17642_));
  XOR2_X1    g16622(.A1(new_n14579_), .A2(new_n13231_), .Z(new_n17643_));
  XOR2_X1    g16623(.A1(new_n17312_), .A2(new_n16018_), .Z(new_n17644_));
  NOR4_X1    g16624(.A1(new_n17484_), .A2(new_n17644_), .A3(new_n17628_), .A4(new_n17643_), .ZN(new_n17645_));
  NOR4_X1    g16625(.A1(new_n17487_), .A2(new_n14580_), .A3(new_n14730_), .A4(new_n17314_), .ZN(new_n17648_));
  NOR2_X1    g16626(.A1(new_n7786_), .A2(new_n7790_), .ZN(new_n17649_));
  OAI21_X1   g16627(.A1(new_n11890_), .A2(new_n11875_), .B(new_n17649_), .ZN(new_n17650_));
  OAI22_X1   g16628(.A1(new_n11859_), .A2(new_n11830_), .B1(new_n11432_), .B2(new_n11873_), .ZN(new_n17651_));
  NAND2_X1   g16629(.A1(new_n11877_), .A2(new_n11878_), .ZN(new_n17652_));
  INV_X1     g16630(.I(new_n11883_), .ZN(new_n17653_));
  AOI21_X1   g16631(.A1(new_n17652_), .A2(new_n7782_), .B(new_n17653_), .ZN(new_n17654_));
  INV_X1     g16632(.I(new_n11889_), .ZN(new_n17655_));
  AOI21_X1   g16633(.A1(new_n17654_), .A2(new_n11879_), .B(new_n17655_), .ZN(new_n17656_));
  INV_X1     g16634(.I(new_n17649_), .ZN(new_n17657_));
  NAND3_X1   g16635(.A1(new_n17656_), .A2(new_n17657_), .A3(new_n17651_), .ZN(new_n17658_));
  AOI21_X1   g16636(.A1(new_n17650_), .A2(new_n17658_), .B(new_n17648_), .ZN(new_n17659_));
  NOR2_X1    g16637(.A1(new_n14730_), .A2(new_n14580_), .ZN(new_n17660_));
  INV_X1     g16638(.I(new_n17314_), .ZN(new_n17661_));
  NAND2_X1   g16639(.A1(new_n17486_), .A2(new_n17661_), .ZN(new_n17662_));
  AOI21_X1   g16640(.A1(new_n17642_), .A2(new_n17645_), .B(new_n17662_), .ZN(new_n17663_));
  NAND3_X1   g16641(.A1(new_n17642_), .A2(new_n17662_), .A3(new_n17645_), .ZN(new_n17664_));
  INV_X1     g16642(.I(new_n17664_), .ZN(new_n17665_));
  OAI21_X1   g16643(.A1(new_n17665_), .A2(new_n17663_), .B(new_n17660_), .ZN(new_n17666_));
  INV_X1     g16644(.I(new_n17660_), .ZN(new_n17667_));
  INV_X1     g16645(.I(new_n17663_), .ZN(new_n17668_));
  NAND3_X1   g16646(.A1(new_n17668_), .A2(new_n17667_), .A3(new_n17664_), .ZN(new_n17669_));
  NAND2_X1   g16647(.A1(new_n17669_), .A2(new_n17666_), .ZN(new_n17670_));
  NOR3_X1    g16648(.A1(new_n17653_), .A2(new_n7778_), .A3(new_n11888_), .ZN(new_n17671_));
  AOI21_X1   g16649(.A1(new_n7779_), .A2(new_n11887_), .B(new_n11883_), .ZN(new_n17672_));
  NOR2_X1    g16650(.A1(new_n17671_), .A2(new_n17672_), .ZN(new_n17673_));
  NOR2_X1    g16651(.A1(new_n17651_), .A2(new_n17673_), .ZN(new_n17674_));
  NAND2_X1   g16652(.A1(new_n17651_), .A2(new_n17673_), .ZN(new_n17675_));
  INV_X1     g16653(.I(new_n17675_), .ZN(new_n17676_));
  OAI21_X1   g16654(.A1(new_n17676_), .A2(new_n17674_), .B(new_n17670_), .ZN(new_n17677_));
  NOR2_X1    g16655(.A1(new_n11865_), .A2(new_n11864_), .ZN(new_n17678_));
  AOI21_X1   g16656(.A1(new_n7766_), .A2(new_n7770_), .B(new_n11860_), .ZN(new_n17679_));
  OAI21_X1   g16657(.A1(new_n17679_), .A2(new_n17678_), .B(new_n11868_), .ZN(new_n17680_));
  INV_X1     g16658(.I(new_n7771_), .ZN(new_n17681_));
  AOI22_X1   g16659(.A1(new_n7766_), .A2(new_n7770_), .B1(new_n7744_), .B2(new_n7748_), .ZN(new_n17682_));
  OAI21_X1   g16660(.A1(new_n17681_), .A2(new_n17682_), .B(new_n7727_), .ZN(new_n17683_));
  AOI21_X1   g16661(.A1(new_n17680_), .A2(new_n17683_), .B(new_n11831_), .ZN(new_n17684_));
  NOR3_X1    g16662(.A1(new_n11867_), .A2(new_n11432_), .A3(new_n11872_), .ZN(new_n17685_));
  NOR3_X1    g16663(.A1(new_n17684_), .A2(new_n11858_), .A3(new_n17685_), .ZN(new_n17686_));
  OAI21_X1   g16664(.A1(new_n11867_), .A2(new_n11872_), .B(new_n11432_), .ZN(new_n17687_));
  NAND3_X1   g16665(.A1(new_n17680_), .A2(new_n17683_), .A3(new_n11831_), .ZN(new_n17688_));
  AOI21_X1   g16666(.A1(new_n17688_), .A2(new_n17687_), .B(new_n11828_), .ZN(new_n17689_));
  NOR2_X1    g16667(.A1(new_n17686_), .A2(new_n17689_), .ZN(new_n17690_));
  NAND3_X1   g16668(.A1(new_n17688_), .A2(new_n17687_), .A3(new_n11828_), .ZN(new_n17691_));
  OAI21_X1   g16669(.A1(new_n17684_), .A2(new_n17685_), .B(new_n11858_), .ZN(new_n17692_));
  NAND2_X1   g16670(.A1(new_n17496_), .A2(new_n17499_), .ZN(new_n17693_));
  NAND2_X1   g16671(.A1(new_n17493_), .A2(new_n17494_), .ZN(new_n17694_));
  AOI21_X1   g16672(.A1(new_n17694_), .A2(new_n17693_), .B(new_n17519_), .ZN(new_n17695_));
  NAND2_X1   g16673(.A1(new_n17496_), .A2(new_n17494_), .ZN(new_n17696_));
  AOI21_X1   g16674(.A1(new_n17696_), .A2(new_n14723_), .B(new_n17490_), .ZN(new_n17697_));
  NOR2_X1    g16675(.A1(new_n17695_), .A2(new_n17697_), .ZN(new_n17698_));
  NOR2_X1    g16676(.A1(new_n17556_), .A2(new_n17559_), .ZN(new_n17699_));
  NOR2_X1    g16677(.A1(new_n17554_), .A2(new_n17553_), .ZN(new_n17700_));
  OAI21_X1   g16678(.A1(new_n17700_), .A2(new_n17699_), .B(new_n17455_), .ZN(new_n17701_));
  NOR2_X1    g16679(.A1(new_n17556_), .A2(new_n17554_), .ZN(new_n17702_));
  OAI21_X1   g16680(.A1(new_n17480_), .A2(new_n17702_), .B(new_n17550_), .ZN(new_n17703_));
  NAND3_X1   g16681(.A1(new_n17698_), .A2(new_n17703_), .A3(new_n17701_), .ZN(new_n17704_));
  AOI21_X1   g16682(.A1(new_n17438_), .A2(new_n17549_), .B(new_n17453_), .ZN(new_n17705_));
  NAND2_X1   g16683(.A1(new_n17437_), .A2(new_n17531_), .ZN(new_n17706_));
  OAI21_X1   g16684(.A1(new_n17582_), .A2(new_n17578_), .B(new_n17545_), .ZN(new_n17707_));
  NAND4_X1   g16685(.A1(new_n17707_), .A2(new_n17526_), .A3(new_n17530_), .A4(new_n17398_), .ZN(new_n17708_));
  AOI21_X1   g16686(.A1(new_n17706_), .A2(new_n17708_), .B(new_n17566_), .ZN(new_n17709_));
  NOR4_X1    g16687(.A1(new_n17705_), .A2(new_n17709_), .A3(new_n17574_), .A4(new_n17575_), .ZN(new_n17710_));
  NOR2_X1    g16688(.A1(new_n17582_), .A2(new_n17581_), .ZN(new_n17711_));
  NOR2_X1    g16689(.A1(new_n17579_), .A2(new_n17578_), .ZN(new_n17712_));
  OAI21_X1   g16690(.A1(new_n17712_), .A2(new_n17711_), .B(new_n17545_), .ZN(new_n17713_));
  INV_X1     g16691(.I(new_n17585_), .ZN(new_n17714_));
  INV_X1     g16692(.I(new_n17597_), .ZN(new_n17715_));
  NOR4_X1    g16693(.A1(new_n17715_), .A2(new_n17598_), .A3(new_n17605_), .A4(new_n17606_), .ZN(new_n17716_));
  NAND3_X1   g16694(.A1(new_n17714_), .A2(new_n17716_), .A3(new_n17713_), .ZN(new_n17717_));
  NAND2_X1   g16695(.A1(new_n17613_), .A2(new_n17610_), .ZN(new_n17718_));
  NAND2_X1   g16696(.A1(new_n17718_), .A2(new_n17611_), .ZN(new_n17719_));
  AOI21_X1   g16697(.A1(new_n17713_), .A2(new_n17714_), .B(new_n17716_), .ZN(new_n17720_));
  OAI21_X1   g16698(.A1(new_n17719_), .A2(new_n17720_), .B(new_n17717_), .ZN(new_n17721_));
  OAI22_X1   g16699(.A1(new_n17705_), .A2(new_n17709_), .B1(new_n17574_), .B2(new_n17575_), .ZN(new_n17722_));
  AOI21_X1   g16700(.A1(new_n17721_), .A2(new_n17722_), .B(new_n17710_), .ZN(new_n17723_));
  AOI21_X1   g16701(.A1(new_n17701_), .A2(new_n17703_), .B(new_n17698_), .ZN(new_n17724_));
  OAI21_X1   g16702(.A1(new_n17724_), .A2(new_n17723_), .B(new_n17704_), .ZN(new_n17725_));
  AOI21_X1   g16703(.A1(new_n17631_), .A2(new_n17632_), .B(new_n13231_), .ZN(new_n17726_));
  NOR3_X1    g16704(.A1(new_n17629_), .A2(new_n17626_), .A3(new_n17625_), .ZN(new_n17727_));
  NOR2_X1    g16705(.A1(new_n17727_), .A2(new_n17726_), .ZN(new_n17728_));
  AOI21_X1   g16706(.A1(new_n17638_), .A2(new_n17639_), .B(new_n16019_), .ZN(new_n17729_));
  NOR3_X1    g16707(.A1(new_n17636_), .A2(new_n17635_), .A3(new_n16018_), .ZN(new_n17730_));
  NOR3_X1    g16708(.A1(new_n17728_), .A2(new_n17729_), .A3(new_n17730_), .ZN(new_n17731_));
  NAND2_X1   g16709(.A1(new_n17630_), .A2(new_n17633_), .ZN(new_n17732_));
  AOI21_X1   g16710(.A1(new_n17637_), .A2(new_n17640_), .B(new_n17732_), .ZN(new_n17733_));
  OAI21_X1   g16711(.A1(new_n17733_), .A2(new_n17731_), .B(new_n17725_), .ZN(new_n17734_));
  NOR3_X1    g16712(.A1(new_n17732_), .A2(new_n17730_), .A3(new_n17729_), .ZN(new_n17735_));
  AOI22_X1   g16713(.A1(new_n17637_), .A2(new_n17640_), .B1(new_n17630_), .B2(new_n17633_), .ZN(new_n17736_));
  OAI21_X1   g16714(.A1(new_n17736_), .A2(new_n17735_), .B(new_n17624_), .ZN(new_n17737_));
  NAND2_X1   g16715(.A1(new_n17734_), .A2(new_n17737_), .ZN(new_n17738_));
  AOI21_X1   g16716(.A1(new_n17692_), .A2(new_n17691_), .B(new_n17738_), .ZN(new_n17739_));
  NAND3_X1   g16717(.A1(new_n17732_), .A2(new_n17637_), .A3(new_n17640_), .ZN(new_n17740_));
  OAI21_X1   g16718(.A1(new_n17729_), .A2(new_n17730_), .B(new_n17728_), .ZN(new_n17741_));
  AOI21_X1   g16719(.A1(new_n17741_), .A2(new_n17740_), .B(new_n17624_), .ZN(new_n17742_));
  OAI22_X1   g16720(.A1(new_n17730_), .A2(new_n17729_), .B1(new_n17726_), .B2(new_n17727_), .ZN(new_n17743_));
  AOI21_X1   g16721(.A1(new_n17743_), .A2(new_n17641_), .B(new_n17725_), .ZN(new_n17744_));
  NOR2_X1    g16722(.A1(new_n17742_), .A2(new_n17744_), .ZN(new_n17745_));
  NOR3_X1    g16723(.A1(new_n17686_), .A2(new_n17689_), .A3(new_n17745_), .ZN(new_n17746_));
  AOI21_X1   g16724(.A1(new_n11708_), .A2(new_n11736_), .B(new_n11740_), .ZN(new_n17747_));
  AOI21_X1   g16725(.A1(new_n11668_), .A2(new_n11684_), .B(new_n11698_), .ZN(new_n17748_));
  NOR3_X1    g16726(.A1(new_n11700_), .A2(new_n11699_), .A3(new_n11648_), .ZN(new_n17749_));
  NOR2_X1    g16727(.A1(new_n17749_), .A2(new_n17748_), .ZN(new_n17750_));
  NOR3_X1    g16728(.A1(new_n11743_), .A2(new_n11745_), .A3(new_n17750_), .ZN(new_n17751_));
  NOR3_X1    g16729(.A1(new_n17747_), .A2(new_n17751_), .A3(new_n11857_), .ZN(new_n17752_));
  OAI21_X1   g16730(.A1(new_n11743_), .A2(new_n11745_), .B(new_n11702_), .ZN(new_n17753_));
  OAI21_X1   g16731(.A1(new_n11700_), .A2(new_n11699_), .B(new_n11648_), .ZN(new_n17754_));
  NAND3_X1   g16732(.A1(new_n11668_), .A2(new_n11698_), .A3(new_n11684_), .ZN(new_n17755_));
  NAND2_X1   g16733(.A1(new_n17754_), .A2(new_n17755_), .ZN(new_n17756_));
  NAND3_X1   g16734(.A1(new_n11708_), .A2(new_n11736_), .A3(new_n17756_), .ZN(new_n17757_));
  AOI21_X1   g16735(.A1(new_n17753_), .A2(new_n17757_), .B(new_n11827_), .ZN(new_n17758_));
  NOR2_X1    g16736(.A1(new_n17752_), .A2(new_n17758_), .ZN(new_n17759_));
  NAND3_X1   g16737(.A1(new_n17753_), .A2(new_n17757_), .A3(new_n11827_), .ZN(new_n17760_));
  OAI21_X1   g16738(.A1(new_n17751_), .A2(new_n17747_), .B(new_n11857_), .ZN(new_n17761_));
  AOI21_X1   g16739(.A1(new_n17701_), .A2(new_n17703_), .B(new_n17523_), .ZN(new_n17762_));
  NOR3_X1    g16740(.A1(new_n17698_), .A2(new_n17561_), .A3(new_n17564_), .ZN(new_n17763_));
  OAI21_X1   g16741(.A1(new_n17762_), .A2(new_n17763_), .B(new_n17622_), .ZN(new_n17764_));
  OAI21_X1   g16742(.A1(new_n17724_), .A2(new_n17565_), .B(new_n17723_), .ZN(new_n17765_));
  NAND2_X1   g16743(.A1(new_n17764_), .A2(new_n17765_), .ZN(new_n17766_));
  AOI21_X1   g16744(.A1(new_n17761_), .A2(new_n17760_), .B(new_n17766_), .ZN(new_n17767_));
  OAI21_X1   g16745(.A1(new_n17561_), .A2(new_n17564_), .B(new_n17698_), .ZN(new_n17768_));
  NAND3_X1   g16746(.A1(new_n17523_), .A2(new_n17703_), .A3(new_n17701_), .ZN(new_n17769_));
  AOI21_X1   g16747(.A1(new_n17768_), .A2(new_n17769_), .B(new_n17723_), .ZN(new_n17770_));
  AOI21_X1   g16748(.A1(new_n17623_), .A2(new_n17704_), .B(new_n17622_), .ZN(new_n17771_));
  NOR2_X1    g16749(.A1(new_n17771_), .A2(new_n17770_), .ZN(new_n17772_));
  NOR3_X1    g16750(.A1(new_n17752_), .A2(new_n17758_), .A3(new_n17772_), .ZN(new_n17773_));
  NAND3_X1   g16751(.A1(new_n11856_), .A2(new_n11766_), .A3(new_n11855_), .ZN(new_n17774_));
  OAI21_X1   g16752(.A1(new_n11840_), .A2(new_n11826_), .B(new_n11825_), .ZN(new_n17775_));
  NOR3_X1    g16753(.A1(new_n17576_), .A2(new_n17705_), .A3(new_n17709_), .ZN(new_n17776_));
  NAND2_X1   g16754(.A1(new_n17619_), .A2(new_n17620_), .ZN(new_n17777_));
  AOI21_X1   g16755(.A1(new_n17568_), .A2(new_n17571_), .B(new_n17777_), .ZN(new_n17778_));
  OAI21_X1   g16756(.A1(new_n17778_), .A2(new_n17776_), .B(new_n17721_), .ZN(new_n17779_));
  OAI21_X1   g16757(.A1(new_n17621_), .A2(new_n17710_), .B(new_n17616_), .ZN(new_n17780_));
  NAND2_X1   g16758(.A1(new_n17779_), .A2(new_n17780_), .ZN(new_n17781_));
  AOI21_X1   g16759(.A1(new_n17775_), .A2(new_n17774_), .B(new_n17781_), .ZN(new_n17782_));
  NOR3_X1    g16760(.A1(new_n11840_), .A2(new_n11826_), .A3(new_n11825_), .ZN(new_n17783_));
  AOI21_X1   g16761(.A1(new_n11856_), .A2(new_n11766_), .B(new_n11855_), .ZN(new_n17784_));
  NAND3_X1   g16762(.A1(new_n17777_), .A2(new_n17568_), .A3(new_n17571_), .ZN(new_n17785_));
  OAI21_X1   g16763(.A1(new_n17705_), .A2(new_n17709_), .B(new_n17576_), .ZN(new_n17786_));
  AOI21_X1   g16764(.A1(new_n17786_), .A2(new_n17785_), .B(new_n17616_), .ZN(new_n17787_));
  AOI21_X1   g16765(.A1(new_n17577_), .A2(new_n17722_), .B(new_n17721_), .ZN(new_n17788_));
  NOR2_X1    g16766(.A1(new_n17787_), .A2(new_n17788_), .ZN(new_n17789_));
  NOR3_X1    g16767(.A1(new_n17783_), .A2(new_n17784_), .A3(new_n17789_), .ZN(new_n17790_));
  NOR3_X1    g16768(.A1(new_n17783_), .A2(new_n17784_), .A3(new_n17789_), .ZN(new_n17791_));
  NOR3_X1    g16769(.A1(new_n17790_), .A2(new_n17791_), .A3(new_n17782_), .ZN(new_n17792_));
  OAI22_X1   g16770(.A1(new_n17767_), .A2(new_n17773_), .B1(new_n17792_), .B2(new_n17759_), .ZN(new_n17793_));
  OAI22_X1   g16771(.A1(new_n17739_), .A2(new_n17746_), .B1(new_n17793_), .B2(new_n17690_), .ZN(new_n17794_));
  AOI21_X1   g16772(.A1(new_n17668_), .A2(new_n17664_), .B(new_n17667_), .ZN(new_n17795_));
  NOR3_X1    g16773(.A1(new_n17665_), .A2(new_n17660_), .A3(new_n17663_), .ZN(new_n17796_));
  NOR2_X1    g16774(.A1(new_n17795_), .A2(new_n17796_), .ZN(new_n17797_));
  INV_X1     g16775(.I(new_n17673_), .ZN(new_n17798_));
  NOR2_X1    g16776(.A1(new_n17798_), .A2(new_n17651_), .ZN(new_n17799_));
  NOR2_X1    g16777(.A1(new_n11875_), .A2(new_n17673_), .ZN(new_n17800_));
  OAI21_X1   g16778(.A1(new_n17800_), .A2(new_n17799_), .B(new_n17797_), .ZN(new_n17801_));
  NAND3_X1   g16779(.A1(new_n17801_), .A2(new_n17677_), .A3(new_n17794_), .ZN(new_n17802_));
  NOR3_X1    g16780(.A1(new_n17802_), .A2(new_n11892_), .A3(new_n17659_), .ZN(new_n17803_));
  INV_X1     g16781(.I(new_n11892_), .ZN(new_n17804_));
  INV_X1     g16782(.I(new_n17659_), .ZN(new_n17805_));
  INV_X1     g16783(.I(new_n17674_), .ZN(new_n17806_));
  AOI21_X1   g16784(.A1(new_n17806_), .A2(new_n17675_), .B(new_n17797_), .ZN(new_n17807_));
  NAND2_X1   g16785(.A1(new_n17692_), .A2(new_n17691_), .ZN(new_n17808_));
  OAI21_X1   g16786(.A1(new_n17686_), .A2(new_n17689_), .B(new_n17745_), .ZN(new_n17809_));
  NAND3_X1   g16787(.A1(new_n17692_), .A2(new_n17691_), .A3(new_n17738_), .ZN(new_n17810_));
  NAND2_X1   g16788(.A1(new_n17761_), .A2(new_n17760_), .ZN(new_n17811_));
  OAI21_X1   g16789(.A1(new_n17752_), .A2(new_n17758_), .B(new_n17772_), .ZN(new_n17812_));
  NAND3_X1   g16790(.A1(new_n17761_), .A2(new_n17760_), .A3(new_n17766_), .ZN(new_n17813_));
  OAI21_X1   g16791(.A1(new_n17783_), .A2(new_n17784_), .B(new_n17789_), .ZN(new_n17814_));
  NAND3_X1   g16792(.A1(new_n17775_), .A2(new_n17774_), .A3(new_n17781_), .ZN(new_n17815_));
  NAND3_X1   g16793(.A1(new_n17775_), .A2(new_n17774_), .A3(new_n17781_), .ZN(new_n17816_));
  NAND3_X1   g16794(.A1(new_n17814_), .A2(new_n17815_), .A3(new_n17816_), .ZN(new_n17817_));
  AOI22_X1   g16795(.A1(new_n17812_), .A2(new_n17813_), .B1(new_n17817_), .B2(new_n17811_), .ZN(new_n17818_));
  AOI22_X1   g16796(.A1(new_n17809_), .A2(new_n17810_), .B1(new_n17818_), .B2(new_n17808_), .ZN(new_n17819_));
  NAND2_X1   g16797(.A1(new_n11875_), .A2(new_n17673_), .ZN(new_n17820_));
  NAND2_X1   g16798(.A1(new_n17798_), .A2(new_n17651_), .ZN(new_n17821_));
  AOI21_X1   g16799(.A1(new_n17820_), .A2(new_n17821_), .B(new_n17670_), .ZN(new_n17822_));
  NOR3_X1    g16800(.A1(new_n17807_), .A2(new_n17822_), .A3(new_n17819_), .ZN(new_n17823_));
  AOI21_X1   g16801(.A1(new_n17823_), .A2(new_n17805_), .B(new_n17804_), .ZN(new_n17824_));
  NOR2_X1    g16802(.A1(new_n17824_), .A2(new_n17803_), .ZN(new_n17825_));
  NAND2_X1   g16803(.A1(new_n11850_), .A2(new_n11811_), .ZN(new_n17826_));
  XOR2_X1    g16804(.A1(new_n14681_), .A2(new_n14683_), .Z(new_n17827_));
  XOR2_X1    g16805(.A1(new_n17422_), .A2(new_n17424_), .Z(new_n17828_));
  NAND2_X1   g16806(.A1(new_n17828_), .A2(new_n17827_), .ZN(new_n17829_));
  INV_X1     g16807(.I(new_n17829_), .ZN(new_n17830_));
  NOR2_X1    g16808(.A1(new_n17828_), .A2(new_n17827_), .ZN(new_n17831_));
  XNOR2_X1   g16809(.A1(new_n11803_), .A2(new_n11806_), .ZN(new_n17832_));
  NOR3_X1    g16810(.A1(new_n17832_), .A2(new_n17830_), .A3(new_n17831_), .ZN(new_n17833_));
  XNOR2_X1   g16811(.A1(new_n17826_), .A2(new_n17833_), .ZN(new_n17834_));
  NOR2_X1    g16812(.A1(new_n14687_), .A2(new_n14685_), .ZN(new_n17835_));
  NAND2_X1   g16813(.A1(new_n17835_), .A2(new_n14688_), .ZN(new_n17836_));
  NAND2_X1   g16814(.A1(new_n17426_), .A2(new_n17427_), .ZN(new_n17837_));
  XOR2_X1    g16815(.A1(new_n17837_), .A2(new_n17430_), .Z(new_n17838_));
  XOR2_X1    g16816(.A1(new_n17838_), .A2(new_n17836_), .Z(new_n17839_));
  XOR2_X1    g16817(.A1(new_n17839_), .A2(new_n17830_), .Z(new_n17840_));
  INV_X1     g16818(.I(new_n17840_), .ZN(new_n17841_));
  AOI21_X1   g16819(.A1(new_n17841_), .A2(new_n17826_), .B(new_n17834_), .ZN(new_n17842_));
  INV_X1     g16820(.I(new_n17842_), .ZN(new_n17843_));
  NAND2_X1   g16821(.A1(new_n11797_), .A2(new_n11798_), .ZN(new_n17844_));
  NOR2_X1    g16822(.A1(new_n17715_), .A2(new_n17598_), .ZN(new_n17845_));
  NOR2_X1    g16823(.A1(new_n17845_), .A2(new_n17607_), .ZN(new_n17846_));
  NOR2_X1    g16824(.A1(new_n17846_), .A2(new_n17716_), .ZN(new_n17847_));
  NOR2_X1    g16825(.A1(new_n11851_), .A2(new_n11816_), .ZN(new_n17848_));
  NAND2_X1   g16826(.A1(new_n11793_), .A2(new_n11791_), .ZN(new_n17849_));
  NOR2_X1    g16827(.A1(new_n17849_), .A2(new_n11812_), .ZN(new_n17850_));
  OAI21_X1   g16828(.A1(new_n17850_), .A2(new_n17848_), .B(new_n17847_), .ZN(new_n17851_));
  NOR3_X1    g16829(.A1(new_n17850_), .A2(new_n17848_), .A3(new_n17847_), .ZN(new_n17852_));
  INV_X1     g16830(.I(new_n17852_), .ZN(new_n17853_));
  AOI21_X1   g16831(.A1(new_n17853_), .A2(new_n17851_), .B(new_n17844_), .ZN(new_n17854_));
  INV_X1     g16832(.I(new_n17851_), .ZN(new_n17855_));
  NOR3_X1    g16833(.A1(new_n17855_), .A2(new_n17852_), .A3(new_n11821_), .ZN(new_n17856_));
  OAI21_X1   g16834(.A1(new_n17856_), .A2(new_n17854_), .B(new_n17843_), .ZN(new_n17857_));
  OAI21_X1   g16835(.A1(new_n17855_), .A2(new_n17852_), .B(new_n11821_), .ZN(new_n17858_));
  NAND3_X1   g16836(.A1(new_n17853_), .A2(new_n17851_), .A3(new_n17844_), .ZN(new_n17859_));
  NAND3_X1   g16837(.A1(new_n17858_), .A2(new_n17859_), .A3(new_n17842_), .ZN(new_n17860_));
  NOR2_X1    g16838(.A1(new_n17830_), .A2(new_n17831_), .ZN(new_n17861_));
  XOR2_X1    g16839(.A1(new_n17861_), .A2(new_n11803_), .Z(new_n17862_));
  XOR2_X1    g16840(.A1(new_n17862_), .A2(new_n11806_), .Z(new_n17863_));
  NOR2_X1    g16841(.A1(new_n17863_), .A2(\A[1000] ), .ZN(new_n17864_));
  INV_X1     g16842(.I(new_n17864_), .ZN(new_n17865_));
  AOI21_X1   g16843(.A1(new_n17834_), .A2(new_n17840_), .B(new_n17865_), .ZN(new_n17866_));
  INV_X1     g16844(.I(new_n17866_), .ZN(new_n17867_));
  AOI21_X1   g16845(.A1(new_n17857_), .A2(new_n17860_), .B(new_n17867_), .ZN(new_n17868_));
  INV_X1     g16846(.I(new_n17868_), .ZN(new_n17869_));
  OAI21_X1   g16847(.A1(new_n17850_), .A2(new_n17848_), .B(new_n11821_), .ZN(new_n17870_));
  OR3_X2     g16848(.A1(new_n17850_), .A2(new_n17848_), .A3(new_n11821_), .Z(new_n17871_));
  NAND2_X1   g16849(.A1(new_n17871_), .A2(new_n17870_), .ZN(new_n17872_));
  NAND2_X1   g16850(.A1(new_n17872_), .A2(new_n17847_), .ZN(new_n17873_));
  OAI21_X1   g16851(.A1(new_n11822_), .A2(new_n11849_), .B(new_n11812_), .ZN(new_n17874_));
  NAND2_X1   g16852(.A1(new_n17844_), .A2(new_n11816_), .ZN(new_n17875_));
  NAND2_X1   g16853(.A1(new_n17849_), .A2(new_n11821_), .ZN(new_n17876_));
  NAND2_X1   g16854(.A1(new_n17876_), .A2(new_n17875_), .ZN(new_n17877_));
  NAND2_X1   g16855(.A1(new_n17877_), .A2(new_n11851_), .ZN(new_n17878_));
  NAND3_X1   g16856(.A1(new_n17878_), .A2(new_n17847_), .A3(new_n17874_), .ZN(new_n17879_));
  NAND2_X1   g16857(.A1(new_n17843_), .A2(new_n17879_), .ZN(new_n17880_));
  NAND2_X1   g16858(.A1(new_n17880_), .A2(new_n17873_), .ZN(new_n17881_));
  NAND3_X1   g16859(.A1(new_n11843_), .A2(new_n11781_), .A3(new_n11844_), .ZN(new_n17882_));
  OAI21_X1   g16860(.A1(new_n11773_), .A2(new_n11774_), .B(new_n11847_), .ZN(new_n17883_));
  AOI21_X1   g16861(.A1(new_n17883_), .A2(new_n17882_), .B(new_n11823_), .ZN(new_n17884_));
  INV_X1     g16862(.I(new_n17884_), .ZN(new_n17885_));
  AOI21_X1   g16863(.A1(new_n11848_), .A2(new_n11824_), .B(new_n11853_), .ZN(new_n17886_));
  INV_X1     g16864(.I(new_n17886_), .ZN(new_n17887_));
  NAND2_X1   g16865(.A1(new_n17615_), .A2(new_n17717_), .ZN(new_n17888_));
  NAND2_X1   g16866(.A1(new_n17888_), .A2(new_n17719_), .ZN(new_n17889_));
  NOR2_X1    g16867(.A1(new_n17584_), .A2(new_n17585_), .ZN(new_n17890_));
  XOR2_X1    g16868(.A1(new_n17890_), .A2(new_n17608_), .Z(new_n17891_));
  OAI21_X1   g16869(.A1(new_n17719_), .A2(new_n17891_), .B(new_n17889_), .ZN(new_n17892_));
  AOI21_X1   g16870(.A1(new_n17885_), .A2(new_n17887_), .B(new_n17892_), .ZN(new_n17893_));
  INV_X1     g16871(.I(new_n17893_), .ZN(new_n17894_));
  NAND3_X1   g16872(.A1(new_n17885_), .A2(new_n17887_), .A3(new_n17892_), .ZN(new_n17895_));
  NAND3_X1   g16873(.A1(new_n17881_), .A2(new_n17894_), .A3(new_n17895_), .ZN(new_n17896_));
  AOI22_X1   g16874(.A1(new_n17843_), .A2(new_n17879_), .B1(new_n17847_), .B2(new_n17872_), .ZN(new_n17897_));
  INV_X1     g16875(.I(new_n17895_), .ZN(new_n17898_));
  OAI21_X1   g16876(.A1(new_n17898_), .A2(new_n17893_), .B(new_n17897_), .ZN(new_n17899_));
  AOI21_X1   g16877(.A1(new_n17899_), .A2(new_n17896_), .B(new_n17869_), .ZN(new_n17900_));
  NAND2_X1   g16878(.A1(new_n11856_), .A2(new_n11766_), .ZN(new_n17901_));
  XOR2_X1    g16879(.A1(new_n17781_), .A2(new_n11855_), .Z(new_n17902_));
  NAND2_X1   g16880(.A1(new_n17902_), .A2(new_n17901_), .ZN(new_n17903_));
  XOR2_X1    g16881(.A1(new_n17781_), .A2(new_n11855_), .Z(new_n17904_));
  OAI21_X1   g16882(.A1(new_n17901_), .A2(new_n17904_), .B(new_n17903_), .ZN(new_n17905_));
  NAND2_X1   g16883(.A1(new_n17905_), .A2(new_n17900_), .ZN(new_n17906_));
  NOR2_X1    g16884(.A1(new_n17751_), .A2(new_n17747_), .ZN(new_n17907_));
  INV_X1     g16885(.I(new_n17907_), .ZN(new_n17908_));
  NAND2_X1   g16886(.A1(new_n17792_), .A2(new_n17908_), .ZN(new_n17909_));
  NAND2_X1   g16887(.A1(new_n17817_), .A2(new_n17907_), .ZN(new_n17910_));
  AOI21_X1   g16888(.A1(new_n17909_), .A2(new_n17910_), .B(new_n11827_), .ZN(new_n17911_));
  NOR2_X1    g16889(.A1(new_n17817_), .A2(new_n17907_), .ZN(new_n17912_));
  NOR2_X1    g16890(.A1(new_n17792_), .A2(new_n17908_), .ZN(new_n17913_));
  NOR3_X1    g16891(.A1(new_n17913_), .A2(new_n17912_), .A3(new_n11857_), .ZN(new_n17914_));
  OAI21_X1   g16892(.A1(new_n17911_), .A2(new_n17914_), .B(new_n17772_), .ZN(new_n17915_));
  OAI21_X1   g16893(.A1(new_n17913_), .A2(new_n17912_), .B(new_n11857_), .ZN(new_n17916_));
  NAND3_X1   g16894(.A1(new_n17909_), .A2(new_n17910_), .A3(new_n11827_), .ZN(new_n17917_));
  NAND3_X1   g16895(.A1(new_n17916_), .A2(new_n17917_), .A3(new_n17766_), .ZN(new_n17918_));
  AOI21_X1   g16896(.A1(new_n17915_), .A2(new_n17918_), .B(new_n17906_), .ZN(new_n17919_));
  NOR2_X1    g16897(.A1(new_n17684_), .A2(new_n17685_), .ZN(new_n17920_));
  INV_X1     g16898(.I(new_n17920_), .ZN(new_n17921_));
  NOR2_X1    g16899(.A1(new_n17738_), .A2(new_n11858_), .ZN(new_n17922_));
  NOR2_X1    g16900(.A1(new_n17745_), .A2(new_n11828_), .ZN(new_n17923_));
  OAI21_X1   g16901(.A1(new_n17922_), .A2(new_n17923_), .B(new_n17921_), .ZN(new_n17924_));
  NOR2_X1    g16902(.A1(new_n17745_), .A2(new_n11858_), .ZN(new_n17925_));
  NOR2_X1    g16903(.A1(new_n17738_), .A2(new_n11828_), .ZN(new_n17926_));
  OAI21_X1   g16904(.A1(new_n17926_), .A2(new_n17925_), .B(new_n17920_), .ZN(new_n17927_));
  NAND3_X1   g16905(.A1(new_n17924_), .A2(new_n17927_), .A3(new_n17818_), .ZN(new_n17928_));
  NAND2_X1   g16906(.A1(new_n17745_), .A2(new_n11828_), .ZN(new_n17929_));
  NAND2_X1   g16907(.A1(new_n17738_), .A2(new_n11858_), .ZN(new_n17930_));
  AOI21_X1   g16908(.A1(new_n17930_), .A2(new_n17929_), .B(new_n17920_), .ZN(new_n17931_));
  NAND2_X1   g16909(.A1(new_n17738_), .A2(new_n11828_), .ZN(new_n17932_));
  NAND2_X1   g16910(.A1(new_n17745_), .A2(new_n11858_), .ZN(new_n17933_));
  AOI21_X1   g16911(.A1(new_n17932_), .A2(new_n17933_), .B(new_n17921_), .ZN(new_n17934_));
  OAI21_X1   g16912(.A1(new_n17931_), .A2(new_n17934_), .B(new_n17793_), .ZN(new_n17935_));
  NAND2_X1   g16913(.A1(new_n17935_), .A2(new_n17928_), .ZN(new_n17936_));
  NAND2_X1   g16914(.A1(new_n17936_), .A2(new_n17919_), .ZN(new_n17937_));
  NAND2_X1   g16915(.A1(new_n17690_), .A2(new_n17738_), .ZN(new_n17938_));
  OAI21_X1   g16916(.A1(new_n17739_), .A2(new_n17746_), .B(new_n17793_), .ZN(new_n17939_));
  NAND3_X1   g16917(.A1(new_n17939_), .A2(new_n17798_), .A3(new_n17938_), .ZN(new_n17940_));
  NAND2_X1   g16918(.A1(new_n17819_), .A2(new_n17673_), .ZN(new_n17941_));
  AOI21_X1   g16919(.A1(new_n17941_), .A2(new_n17940_), .B(new_n11875_), .ZN(new_n17942_));
  NOR2_X1    g16920(.A1(new_n17819_), .A2(new_n17673_), .ZN(new_n17943_));
  NOR2_X1    g16921(.A1(new_n17794_), .A2(new_n17798_), .ZN(new_n17944_));
  NOR3_X1    g16922(.A1(new_n17944_), .A2(new_n17943_), .A3(new_n17651_), .ZN(new_n17945_));
  OAI21_X1   g16923(.A1(new_n17945_), .A2(new_n17942_), .B(new_n17797_), .ZN(new_n17946_));
  OAI21_X1   g16924(.A1(new_n17944_), .A2(new_n17943_), .B(new_n17651_), .ZN(new_n17947_));
  NAND3_X1   g16925(.A1(new_n17941_), .A2(new_n17940_), .A3(new_n11875_), .ZN(new_n17948_));
  NAND3_X1   g16926(.A1(new_n17947_), .A2(new_n17948_), .A3(new_n17670_), .ZN(new_n17949_));
  AOI21_X1   g16927(.A1(new_n17946_), .A2(new_n17949_), .B(new_n17937_), .ZN(new_n17950_));
  AOI21_X1   g16928(.A1(new_n17656_), .A2(new_n17651_), .B(new_n17657_), .ZN(new_n17951_));
  NOR3_X1    g16929(.A1(new_n11890_), .A2(new_n11875_), .A3(new_n17649_), .ZN(new_n17952_));
  NOR3_X1    g16930(.A1(new_n17952_), .A2(new_n17951_), .A3(new_n17648_), .ZN(new_n17953_));
  NAND2_X1   g16931(.A1(new_n17802_), .A2(new_n17953_), .ZN(new_n17954_));
  INV_X1     g16932(.I(new_n17648_), .ZN(new_n17955_));
  NAND3_X1   g16933(.A1(new_n17650_), .A2(new_n17658_), .A3(new_n17955_), .ZN(new_n17956_));
  NAND2_X1   g16934(.A1(new_n17823_), .A2(new_n17956_), .ZN(new_n17957_));
  NAND2_X1   g16935(.A1(new_n17957_), .A2(new_n17954_), .ZN(new_n17958_));
  NAND3_X1   g16936(.A1(new_n17950_), .A2(new_n17825_), .A3(new_n17958_), .ZN(new_n17959_));
  NAND3_X1   g16937(.A1(new_n17823_), .A2(new_n17805_), .A3(new_n17804_), .ZN(new_n17960_));
  OAI21_X1   g16938(.A1(new_n17802_), .A2(new_n17659_), .B(new_n11892_), .ZN(new_n17961_));
  NAND2_X1   g16939(.A1(new_n17960_), .A2(new_n17961_), .ZN(new_n17962_));
  NOR3_X1    g16940(.A1(new_n17898_), .A2(new_n17897_), .A3(new_n17893_), .ZN(new_n17963_));
  AOI21_X1   g16941(.A1(new_n17895_), .A2(new_n17894_), .B(new_n17881_), .ZN(new_n17964_));
  OAI21_X1   g16942(.A1(new_n17964_), .A2(new_n17963_), .B(new_n17868_), .ZN(new_n17965_));
  NOR2_X1    g16943(.A1(new_n17904_), .A2(new_n17901_), .ZN(new_n17966_));
  AOI21_X1   g16944(.A1(new_n17901_), .A2(new_n17902_), .B(new_n17966_), .ZN(new_n17967_));
  NOR2_X1    g16945(.A1(new_n17967_), .A2(new_n17965_), .ZN(new_n17968_));
  AOI21_X1   g16946(.A1(new_n17916_), .A2(new_n17917_), .B(new_n17766_), .ZN(new_n17969_));
  NOR3_X1    g16947(.A1(new_n17911_), .A2(new_n17914_), .A3(new_n17772_), .ZN(new_n17970_));
  OAI21_X1   g16948(.A1(new_n17970_), .A2(new_n17969_), .B(new_n17968_), .ZN(new_n17971_));
  NOR3_X1    g16949(.A1(new_n17931_), .A2(new_n17934_), .A3(new_n17793_), .ZN(new_n17972_));
  AOI21_X1   g16950(.A1(new_n17924_), .A2(new_n17927_), .B(new_n17818_), .ZN(new_n17973_));
  NOR2_X1    g16951(.A1(new_n17973_), .A2(new_n17972_), .ZN(new_n17974_));
  NOR2_X1    g16952(.A1(new_n17974_), .A2(new_n17971_), .ZN(new_n17975_));
  AOI21_X1   g16953(.A1(new_n17947_), .A2(new_n17948_), .B(new_n17670_), .ZN(new_n17976_));
  NOR3_X1    g16954(.A1(new_n17945_), .A2(new_n17942_), .A3(new_n17797_), .ZN(new_n17977_));
  OAI21_X1   g16955(.A1(new_n17977_), .A2(new_n17976_), .B(new_n17975_), .ZN(new_n17978_));
  NOR2_X1    g16956(.A1(new_n17823_), .A2(new_n17956_), .ZN(new_n17979_));
  NOR2_X1    g16957(.A1(new_n17802_), .A2(new_n17953_), .ZN(new_n17980_));
  NOR2_X1    g16958(.A1(new_n17979_), .A2(new_n17980_), .ZN(new_n17981_));
  OAI21_X1   g16959(.A1(new_n17978_), .A2(new_n17981_), .B(new_n17962_), .ZN(new_n17982_));
  NAND2_X1   g16960(.A1(new_n17982_), .A2(new_n17959_), .ZN(new_n17983_));
  AOI21_X1   g16961(.A1(new_n17915_), .A2(new_n17918_), .B(new_n17968_), .ZN(new_n17984_));
  NAND3_X1   g16962(.A1(new_n17915_), .A2(new_n17918_), .A3(new_n17968_), .ZN(new_n17985_));
  INV_X1     g16963(.I(new_n17985_), .ZN(new_n17986_));
  NAND2_X1   g16964(.A1(new_n17967_), .A2(new_n17900_), .ZN(new_n17987_));
  NAND2_X1   g16965(.A1(new_n17905_), .A2(new_n17965_), .ZN(new_n17988_));
  NAND2_X1   g16966(.A1(new_n17987_), .A2(new_n17988_), .ZN(new_n17989_));
  AOI21_X1   g16967(.A1(new_n17894_), .A2(new_n17895_), .B(new_n17897_), .ZN(new_n17990_));
  NOR3_X1    g16968(.A1(new_n17881_), .A2(new_n17898_), .A3(new_n17893_), .ZN(new_n17991_));
  OAI21_X1   g16969(.A1(new_n17991_), .A2(new_n17990_), .B(new_n17868_), .ZN(new_n17992_));
  OAI21_X1   g16970(.A1(new_n17963_), .A2(new_n17964_), .B(new_n17869_), .ZN(new_n17993_));
  NAND3_X1   g16971(.A1(new_n17834_), .A2(new_n17840_), .A3(new_n17865_), .ZN(new_n17994_));
  NAND2_X1   g16972(.A1(new_n17867_), .A2(new_n17994_), .ZN(new_n17995_));
  AOI21_X1   g16973(.A1(new_n17857_), .A2(new_n17860_), .B(new_n17866_), .ZN(new_n17996_));
  NAND2_X1   g16974(.A1(new_n17857_), .A2(new_n17860_), .ZN(new_n17997_));
  NOR2_X1    g16975(.A1(new_n17997_), .A2(new_n17867_), .ZN(new_n17998_));
  NOR2_X1    g16976(.A1(new_n17998_), .A2(new_n17996_), .ZN(new_n17999_));
  AOI22_X1   g16977(.A1(new_n17993_), .A2(new_n17992_), .B1(new_n17995_), .B2(new_n17999_), .ZN(new_n18000_));
  OAI22_X1   g16978(.A1(new_n17986_), .A2(new_n17984_), .B1(new_n17989_), .B2(new_n18000_), .ZN(new_n18001_));
  NOR2_X1    g16979(.A1(new_n17936_), .A2(new_n17971_), .ZN(new_n18002_));
  NOR2_X1    g16980(.A1(new_n17974_), .A2(new_n17919_), .ZN(new_n18003_));
  NOR2_X1    g16981(.A1(new_n18003_), .A2(new_n18002_), .ZN(new_n18004_));
  NOR2_X1    g16982(.A1(new_n18004_), .A2(new_n18001_), .ZN(new_n18005_));
  AOI21_X1   g16983(.A1(new_n17946_), .A2(new_n17949_), .B(new_n17975_), .ZN(new_n18006_));
  NOR3_X1    g16984(.A1(new_n17977_), .A2(new_n17976_), .A3(new_n17937_), .ZN(new_n18007_));
  OAI21_X1   g16985(.A1(new_n18006_), .A2(new_n18007_), .B(new_n18005_), .ZN(new_n18008_));
  NOR2_X1    g16986(.A1(new_n17950_), .A2(new_n17981_), .ZN(new_n18009_));
  NOR2_X1    g16987(.A1(new_n17978_), .A2(new_n17958_), .ZN(new_n18010_));
  NOR2_X1    g16988(.A1(new_n18010_), .A2(new_n18009_), .ZN(new_n18011_));
  NOR3_X1    g16989(.A1(new_n17983_), .A2(new_n18011_), .A3(new_n18008_), .ZN(new_n18012_));
  NOR2_X1    g16990(.A1(new_n17802_), .A2(new_n17659_), .ZN(new_n18013_));
  NOR2_X1    g16991(.A1(new_n18013_), .A2(new_n11892_), .ZN(new_n18014_));
  NAND4_X1   g16992(.A1(new_n17950_), .A2(new_n11892_), .A3(new_n17958_), .A4(new_n18013_), .ZN(new_n18015_));
  NAND2_X1   g16993(.A1(new_n17946_), .A2(new_n17949_), .ZN(new_n18016_));
  NAND2_X1   g16994(.A1(new_n17650_), .A2(new_n17658_), .ZN(new_n18017_));
  INV_X1     g16995(.I(new_n18017_), .ZN(new_n18018_));
  NAND4_X1   g16996(.A1(new_n17823_), .A2(new_n17804_), .A3(new_n18018_), .A4(new_n17955_), .ZN(new_n18019_));
  NOR2_X1    g16997(.A1(new_n17823_), .A2(new_n17953_), .ZN(new_n18020_));
  NOR4_X1    g16998(.A1(new_n18019_), .A2(new_n18013_), .A3(new_n18020_), .A4(new_n17937_), .ZN(new_n18021_));
  NAND3_X1   g16999(.A1(new_n18021_), .A2(new_n17825_), .A3(new_n18016_), .ZN(new_n18022_));
  NAND4_X1   g17000(.A1(new_n18022_), .A2(new_n18015_), .A3(new_n17982_), .A4(new_n18014_), .ZN(new_n18023_));
  NOR2_X1    g17001(.A1(new_n18012_), .A2(new_n18023_), .ZN(new_n18024_));
  NOR2_X1    g17002(.A1(new_n18011_), .A2(new_n18008_), .ZN(new_n18025_));
  NAND4_X1   g17003(.A1(new_n18025_), .A2(new_n18014_), .A3(new_n17959_), .A4(new_n17982_), .ZN(new_n18026_));
  OAI21_X1   g17004(.A1(new_n17970_), .A2(new_n17969_), .B(new_n17906_), .ZN(new_n18027_));
  NOR2_X1    g17005(.A1(new_n17989_), .A2(new_n18000_), .ZN(new_n18028_));
  AOI21_X1   g17006(.A1(new_n18027_), .A2(new_n17985_), .B(new_n18028_), .ZN(new_n18029_));
  OAI21_X1   g17007(.A1(new_n18002_), .A2(new_n18003_), .B(new_n18029_), .ZN(new_n18030_));
  NOR2_X1    g17008(.A1(new_n18007_), .A2(new_n18006_), .ZN(new_n18031_));
  NAND3_X1   g17009(.A1(new_n17993_), .A2(new_n17992_), .A3(new_n17999_), .ZN(new_n18032_));
  NAND3_X1   g17010(.A1(new_n17997_), .A2(new_n17867_), .A3(new_n17994_), .ZN(new_n18033_));
  XOR2_X1    g17011(.A1(new_n17862_), .A2(\A[1000] ), .Z(new_n18034_));
  XOR2_X1    g17012(.A1(new_n18034_), .A2(new_n11806_), .Z(new_n18035_));
  OAI21_X1   g17013(.A1(new_n17999_), .A2(new_n18035_), .B(new_n17995_), .ZN(new_n18036_));
  NAND2_X1   g17014(.A1(new_n18036_), .A2(new_n18033_), .ZN(new_n18037_));
  NAND2_X1   g17015(.A1(new_n18037_), .A2(new_n18032_), .ZN(new_n18038_));
  AOI22_X1   g17016(.A1(new_n18038_), .A2(new_n18000_), .B1(new_n17987_), .B2(new_n17988_), .ZN(new_n18039_));
  OAI21_X1   g17017(.A1(new_n17984_), .A2(new_n17986_), .B(new_n18039_), .ZN(new_n18040_));
  OAI21_X1   g17018(.A1(new_n18029_), .A2(new_n18004_), .B(new_n18040_), .ZN(new_n18041_));
  OAI21_X1   g17019(.A1(new_n18031_), .A2(new_n18030_), .B(new_n18041_), .ZN(new_n18042_));
  NAND2_X1   g17020(.A1(new_n17978_), .A2(new_n17958_), .ZN(new_n18043_));
  NAND2_X1   g17021(.A1(new_n17950_), .A2(new_n17981_), .ZN(new_n18044_));
  NAND3_X1   g17022(.A1(new_n18008_), .A2(new_n18043_), .A3(new_n18044_), .ZN(new_n18045_));
  OAI21_X1   g17023(.A1(new_n17977_), .A2(new_n17976_), .B(new_n17937_), .ZN(new_n18046_));
  NAND3_X1   g17024(.A1(new_n17946_), .A2(new_n17949_), .A3(new_n17975_), .ZN(new_n18047_));
  AOI21_X1   g17025(.A1(new_n18046_), .A2(new_n18047_), .B(new_n18030_), .ZN(new_n18048_));
  NAND3_X1   g17026(.A1(new_n18048_), .A2(new_n18043_), .A3(new_n18044_), .ZN(new_n18049_));
  AOI21_X1   g17027(.A1(new_n18045_), .A2(new_n18049_), .B(new_n18042_), .ZN(new_n18050_));
  NAND2_X1   g17028(.A1(new_n18050_), .A2(new_n18012_), .ZN(new_n18051_));
  AOI21_X1   g17029(.A1(new_n18051_), .A2(new_n18026_), .B(new_n18024_), .ZN(maj));
endmodule


