// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:30 2022

module ibm  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43,
    v44, v45, v46, v47,
    \v48.0 , \v48.1 , \v48.2 , \v48.3 , \v48.4 , \v48.5 , \v48.6 , \v48.7 ,
    \v48.8 , \v48.9 , \v48.10 , \v48.11 , \v48.12 , \v48.13 , \v48.14 ,
    \v48.15 , \v48.16   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42,
    v43, v44, v45, v46, v47;
  output \v48.0 , \v48.1 , \v48.2 , \v48.3 , \v48.4 , \v48.5 , \v48.6 ,
    \v48.7 , \v48.8 , \v48.9 , \v48.10 , \v48.11 , \v48.12 , \v48.13 ,
    \v48.14 , \v48.15 , \v48.16 ;
  wire new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_;
  assign new_n66_ = ~v3 & ~v9;
  assign new_n67_ = v0 & v1;
  assign new_n68_ = v2 & ~v5;
  assign new_n69_ = new_n67_ & new_n68_;
  assign new_n70_ = ~v2 & v5;
  assign new_n71_ = v12 & v13;
  assign new_n72_ = new_n70_ & new_n71_;
  assign new_n73_ = ~new_n69_ & ~new_n72_;
  assign new_n74_ = ~new_n66_ & ~new_n73_;
  assign new_n75_ = v9 & v11;
  assign new_n76_ = ~v9 & v12;
  assign new_n77_ = ~v3 & new_n76_;
  assign new_n78_ = ~new_n75_ & ~new_n77_;
  assign new_n79_ = v5 & ~new_n78_;
  assign new_n80_ = v2 & new_n79_;
  assign new_n81_ = ~new_n74_ & ~new_n80_;
  assign new_n82_ = v4 & ~new_n81_;
  assign new_n83_ = v2 & ~new_n66_;
  assign new_n84_ = ~v5 & ~new_n83_;
  assign new_n85_ = v4 & ~new_n84_;
  assign new_n86_ = v15 & ~new_n85_;
  assign new_n87_ = ~new_n82_ & ~new_n86_;
  assign new_n88_ = ~v8 & ~new_n87_;
  assign new_n89_ = v3 & v4;
  assign new_n90_ = v2 & new_n89_;
  assign new_n91_ = ~v10 & v11;
  assign new_n92_ = v5 & new_n91_;
  assign new_n93_ = new_n90_ & new_n92_;
  assign new_n94_ = ~v4 & ~v5;
  assign new_n95_ = v8 & ~v16;
  assign new_n96_ = new_n94_ & new_n95_;
  assign new_n97_ = ~new_n93_ & ~new_n96_;
  assign new_n98_ = ~new_n88_ & new_n97_;
  assign new_n99_ = v6 & ~new_n98_;
  assign new_n100_ = ~v4 & v5;
  assign new_n101_ = ~v8 & v15;
  assign new_n102_ = new_n100_ & new_n101_;
  assign new_n103_ = ~new_n99_ & ~new_n102_;
  assign new_n104_ = v7 & ~new_n103_;
  assign new_n105_ = v1 & new_n83_;
  assign new_n106_ = v0 & new_n105_;
  assign new_n107_ = v15 & ~new_n83_;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = v14 & ~new_n108_;
  assign new_n110_ = ~v7 & v15;
  assign new_n111_ = ~v6 & new_n110_;
  assign new_n112_ = new_n94_ & new_n111_;
  assign new_n113_ = ~new_n109_ & ~new_n112_;
  assign \v48.0  = new_n104_ | ~new_n113_;
  assign new_n115_ = ~v5 & v6;
  assign new_n116_ = ~v4 & new_n115_;
  assign new_n117_ = v7 & new_n95_;
  assign new_n118_ = new_n116_ & new_n117_;
  assign new_n119_ = ~v14 & ~new_n118_;
  assign new_n120_ = v2 & v11;
  assign new_n121_ = ~v2 & new_n71_;
  assign new_n122_ = ~new_n120_ & ~new_n121_;
  assign new_n123_ = ~new_n119_ & ~new_n122_;
  assign new_n124_ = v4 & ~v5;
  assign new_n125_ = v2 & new_n124_;
  assign new_n126_ = v6 & v7;
  assign new_n127_ = ~v8 & v11;
  assign new_n128_ = new_n126_ & new_n127_;
  assign new_n129_ = new_n125_ & new_n128_;
  assign new_n130_ = ~new_n123_ & ~new_n129_;
  assign new_n131_ = ~new_n66_ & ~new_n130_;
  assign new_n132_ = v12 & ~new_n119_;
  assign new_n133_ = v2 & new_n132_;
  assign new_n134_ = ~v8 & v17;
  assign new_n135_ = v7 & new_n134_;
  assign new_n136_ = new_n115_ & new_n135_;
  assign new_n137_ = ~new_n133_ & ~new_n136_;
  assign new_n138_ = ~v9 & ~new_n137_;
  assign new_n139_ = ~v3 & new_n138_;
  assign new_n140_ = v5 & ~v8;
  assign new_n141_ = ~new_n115_ & ~new_n140_;
  assign new_n142_ = ~v4 & ~new_n141_;
  assign new_n143_ = ~v2 & ~v5;
  assign new_n144_ = v6 & ~v8;
  assign new_n145_ = new_n143_ & new_n144_;
  assign new_n146_ = ~new_n142_ & ~new_n145_;
  assign new_n147_ = v17 & ~new_n146_;
  assign new_n148_ = v7 & new_n147_;
  assign new_n149_ = ~new_n139_ & ~new_n148_;
  assign \v48.1  = new_n131_ | ~new_n149_;
  assign new_n151_ = v4 & v6;
  assign new_n152_ = v7 & ~v8;
  assign new_n153_ = new_n151_ & new_n152_;
  assign new_n154_ = ~v14 & ~new_n153_;
  assign new_n155_ = ~v16 & ~new_n67_;
  assign new_n156_ = new_n83_ & ~new_n155_;
  assign new_n157_ = v18 & ~new_n156_;
  assign new_n158_ = v16 & v19;
  assign new_n159_ = ~new_n157_ & ~new_n158_;
  assign new_n160_ = ~new_n154_ & ~new_n159_;
  assign new_n161_ = ~v6 & ~v7;
  assign new_n162_ = ~new_n126_ & ~new_n161_;
  assign new_n163_ = ~v5 & ~new_n162_;
  assign new_n164_ = v5 & new_n152_;
  assign new_n165_ = ~new_n163_ & ~new_n164_;
  assign new_n166_ = v18 & ~new_n165_;
  assign new_n167_ = ~v4 & new_n166_;
  assign \v48.2  = new_n160_ | new_n167_;
  assign new_n169_ = v16 & v21;
  assign new_n170_ = ~v0 & ~v16;
  assign new_n171_ = ~new_n66_ & ~new_n170_;
  assign new_n172_ = v2 & new_n171_;
  assign new_n173_ = v20 & ~new_n172_;
  assign new_n174_ = ~new_n169_ & ~new_n173_;
  assign new_n175_ = ~new_n154_ & ~new_n174_;
  assign new_n176_ = ~v8 & v16;
  assign new_n177_ = v7 & new_n176_;
  assign new_n178_ = new_n151_ & new_n177_;
  assign new_n179_ = v14 & ~v16;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = ~v1 & ~new_n180_;
  assign new_n182_ = ~v4 & ~new_n165_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = v20 & ~new_n183_;
  assign \v48.3  = new_n175_ | new_n184_;
  assign new_n186_ = ~v0 & ~new_n180_;
  assign new_n187_ = ~v1 & ~v16;
  assign new_n188_ = ~new_n66_ & ~new_n187_;
  assign new_n189_ = v2 & new_n188_;
  assign new_n190_ = ~new_n154_ & ~new_n189_;
  assign new_n191_ = ~new_n182_ & ~new_n190_;
  assign new_n192_ = ~new_n186_ & new_n191_;
  assign new_n193_ = v22 & ~new_n192_;
  assign new_n194_ = v23 & ~new_n154_;
  assign new_n195_ = v16 & new_n194_;
  assign \v48.4  = new_n193_ | new_n195_;
  assign new_n197_ = v24 & ~new_n156_;
  assign new_n198_ = v16 & v25;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~new_n154_ & ~new_n199_;
  assign new_n201_ = v24 & ~new_n165_;
  assign new_n202_ = ~v4 & new_n201_;
  assign \v48.5  = new_n200_ | new_n202_;
  assign new_n204_ = v27 & ~new_n154_;
  assign new_n205_ = v16 & new_n204_;
  assign new_n206_ = v4 & v5;
  assign new_n207_ = new_n152_ & new_n206_;
  assign new_n208_ = ~v14 & ~new_n207_;
  assign new_n209_ = ~v0 & ~new_n208_;
  assign new_n210_ = ~v1 & ~new_n154_;
  assign new_n211_ = ~new_n209_ & ~new_n210_;
  assign new_n212_ = ~v16 & ~new_n211_;
  assign new_n213_ = ~new_n83_ & ~new_n154_;
  assign new_n214_ = ~v6 & v8;
  assign new_n215_ = v7 & ~new_n214_;
  assign new_n216_ = ~new_n161_ & ~new_n215_;
  assign new_n217_ = ~v5 & ~new_n216_;
  assign new_n218_ = ~v4 & new_n217_;
  assign new_n219_ = ~new_n213_ & ~new_n218_;
  assign new_n220_ = ~new_n212_ & new_n219_;
  assign new_n221_ = v26 & ~new_n220_;
  assign \v48.6  = new_n205_ | new_n221_;
  assign new_n223_ = v28 & ~new_n156_;
  assign new_n224_ = v16 & v29;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = ~new_n154_ & ~new_n225_;
  assign new_n227_ = v28 & ~new_n165_;
  assign new_n228_ = ~v4 & new_n227_;
  assign \v48.7  = new_n226_ | new_n228_;
  assign new_n230_ = ~v16 & v30;
  assign new_n231_ = v16 & v31;
  assign new_n232_ = ~new_n230_ & ~new_n231_;
  assign new_n233_ = ~new_n154_ & ~new_n232_;
  assign new_n234_ = ~v5 & ~v6;
  assign new_n235_ = ~new_n140_ & ~new_n234_;
  assign new_n236_ = v30 & ~new_n235_;
  assign new_n237_ = v7 & new_n236_;
  assign new_n238_ = ~v4 & new_n237_;
  assign \v48.8  = new_n233_ | new_n238_;
  assign new_n240_ = ~v16 & v32;
  assign new_n241_ = v16 & v33;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign new_n243_ = ~new_n154_ & ~new_n242_;
  assign new_n244_ = v32 & ~new_n165_;
  assign new_n245_ = ~v4 & new_n244_;
  assign \v48.9  = new_n243_ | new_n245_;
  assign new_n247_ = ~v16 & v34;
  assign new_n248_ = v16 & v35;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = ~new_n154_ & ~new_n249_;
  assign new_n251_ = v34 & ~new_n165_;
  assign new_n252_ = ~v4 & new_n251_;
  assign \v48.10  = new_n250_ | new_n252_;
  assign new_n254_ = ~v16 & v36;
  assign new_n255_ = v16 & v37;
  assign new_n256_ = ~new_n254_ & ~new_n255_;
  assign new_n257_ = ~new_n154_ & ~new_n256_;
  assign new_n258_ = v36 & ~new_n165_;
  assign new_n259_ = ~v4 & new_n258_;
  assign \v48.11  = new_n257_ | new_n259_;
  assign new_n261_ = ~v16 & v38;
  assign new_n262_ = v16 & v39;
  assign new_n263_ = ~new_n261_ & ~new_n262_;
  assign new_n264_ = ~new_n154_ & ~new_n263_;
  assign new_n265_ = v38 & ~new_n165_;
  assign new_n266_ = ~v4 & new_n265_;
  assign \v48.12  = new_n264_ | new_n266_;
  assign new_n268_ = ~v16 & v40;
  assign new_n269_ = v16 & v41;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = ~new_n154_ & ~new_n270_;
  assign new_n272_ = v40 & ~new_n165_;
  assign new_n273_ = ~v4 & new_n272_;
  assign \v48.13  = new_n271_ | new_n273_;
  assign new_n275_ = ~v16 & v42;
  assign new_n276_ = v16 & v43;
  assign new_n277_ = ~new_n275_ & ~new_n276_;
  assign new_n278_ = ~v8 & ~new_n277_;
  assign new_n279_ = v4 & new_n278_;
  assign new_n280_ = ~v5 & v42;
  assign new_n281_ = ~v4 & new_n280_;
  assign new_n282_ = ~new_n279_ & ~new_n281_;
  assign new_n283_ = v6 & ~new_n282_;
  assign new_n284_ = ~v8 & v42;
  assign new_n285_ = new_n100_ & new_n284_;
  assign new_n286_ = ~new_n283_ & ~new_n285_;
  assign new_n287_ = v7 & ~new_n286_;
  assign new_n288_ = v11 & ~v16;
  assign new_n289_ = ~new_n276_ & ~new_n288_;
  assign new_n290_ = v14 & ~new_n289_;
  assign new_n291_ = ~v7 & v42;
  assign new_n292_ = ~v6 & new_n291_;
  assign new_n293_ = new_n94_ & new_n292_;
  assign new_n294_ = ~new_n290_ & ~new_n293_;
  assign \v48.14  = new_n287_ | ~new_n294_;
  assign new_n296_ = ~v16 & v44;
  assign new_n297_ = v16 & v45;
  assign new_n298_ = ~new_n296_ & ~new_n297_;
  assign new_n299_ = ~new_n154_ & ~new_n298_;
  assign new_n300_ = v44 & ~new_n165_;
  assign new_n301_ = ~v4 & new_n300_;
  assign \v48.15  = new_n299_ | new_n301_;
  assign new_n303_ = ~v16 & v46;
  assign new_n304_ = v16 & v47;
  assign new_n305_ = ~new_n303_ & ~new_n304_;
  assign new_n306_ = ~new_n154_ & ~new_n305_;
  assign new_n307_ = v46 & ~new_n165_;
  assign new_n308_ = ~v4 & new_n307_;
  assign \v48.16  = new_n306_ | new_n308_;
endmodule


