// Benchmark "bar" written by ABC on Mon Sep  4 17:54:07 2023

module bar ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2564_, new_n2565_,
    new_n2567_, new_n2568_, new_n2570_, new_n2571_, new_n2573_, new_n2574_,
    new_n2576_, new_n2577_, new_n2579_, new_n2580_, new_n2582_, new_n2583_,
    new_n2585_, new_n2586_, new_n2588_, new_n2589_, new_n2591_, new_n2592_,
    new_n2594_, new_n2595_, new_n2597_, new_n2598_, new_n2600_, new_n2601_,
    new_n2603_, new_n2604_, new_n2606_, new_n2607_, new_n2609_, new_n2610_,
    new_n2612_, new_n2613_, new_n2615_, new_n2616_, new_n2618_, new_n2619_,
    new_n2621_, new_n2622_, new_n2624_, new_n2625_, new_n2627_, new_n2628_,
    new_n2630_, new_n2631_, new_n2633_, new_n2634_, new_n2636_, new_n2637_,
    new_n2639_, new_n2640_, new_n2642_, new_n2643_, new_n2645_, new_n2646_,
    new_n2648_, new_n2649_, new_n2651_, new_n2652_, new_n2654_, new_n2655_,
    new_n2657_, new_n2658_, new_n2660_, new_n2661_, new_n2663_, new_n2664_,
    new_n2666_, new_n2667_, new_n2669_, new_n2670_, new_n2672_, new_n2673_,
    new_n2675_, new_n2676_, new_n2678_, new_n2679_, new_n2681_, new_n2682_,
    new_n2684_, new_n2685_, new_n2687_, new_n2688_, new_n2690_, new_n2691_,
    new_n2693_, new_n2694_, new_n2696_, new_n2697_, new_n2699_, new_n2700_,
    new_n2702_, new_n2703_, new_n2705_, new_n2706_, new_n2708_, new_n2709_,
    new_n2711_, new_n2712_, new_n2714_, new_n2715_, new_n2717_, new_n2718_,
    new_n2720_, new_n2721_, new_n2723_, new_n2724_, new_n2726_, new_n2727_,
    new_n2729_, new_n2730_, new_n2732_, new_n2733_, new_n2735_, new_n2736_,
    new_n2738_, new_n2739_, new_n2741_, new_n2742_, new_n2744_, new_n2745_,
    new_n2747_, new_n2748_, new_n2750_, new_n2751_, new_n2753_, new_n2754_;
  INV_X1     g0000(.I(\shift[6] ), .ZN(new_n264_));
  NAND3_X1   g0001(.A1(\a[77] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n265_));
  INV_X1     g0002(.I(\shift[0] ), .ZN(new_n266_));
  NAND3_X1   g0003(.A1(new_n266_), .A2(\a[78] ), .A3(\shift[1] ), .ZN(new_n267_));
  NAND2_X1   g0004(.A1(new_n267_), .A2(new_n265_), .ZN(new_n268_));
  NAND2_X1   g0005(.A1(new_n266_), .A2(\a[80] ), .ZN(new_n269_));
  NAND2_X1   g0006(.A1(\a[79] ), .A2(\shift[0] ), .ZN(new_n270_));
  AOI21_X1   g0007(.A1(new_n269_), .A2(new_n270_), .B(\shift[1] ), .ZN(new_n271_));
  NOR2_X1    g0008(.A1(new_n271_), .A2(new_n268_), .ZN(new_n272_));
  NOR2_X1    g0009(.A1(\shift[2] ), .A2(\shift[3] ), .ZN(new_n273_));
  INV_X1     g0010(.I(new_n273_), .ZN(new_n274_));
  INV_X1     g0011(.I(\shift[1] ), .ZN(new_n275_));
  NAND2_X1   g0012(.A1(\a[73] ), .A2(\shift[0] ), .ZN(new_n276_));
  NAND2_X1   g0013(.A1(new_n266_), .A2(\a[74] ), .ZN(new_n277_));
  AOI21_X1   g0014(.A1(new_n277_), .A2(new_n276_), .B(new_n275_), .ZN(new_n278_));
  NAND2_X1   g0015(.A1(new_n266_), .A2(\a[76] ), .ZN(new_n279_));
  NAND2_X1   g0016(.A1(\a[75] ), .A2(\shift[0] ), .ZN(new_n280_));
  AOI21_X1   g0017(.A1(new_n279_), .A2(new_n280_), .B(\shift[1] ), .ZN(new_n281_));
  NOR2_X1    g0018(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1     g0019(.I(\shift[2] ), .ZN(new_n283_));
  NOR2_X1    g0020(.A1(new_n283_), .A2(\shift[3] ), .ZN(new_n284_));
  INV_X1     g0021(.I(new_n284_), .ZN(new_n285_));
  OAI22_X1   g0022(.A1(new_n282_), .A2(new_n285_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n286_));
  NAND2_X1   g0023(.A1(\a[65] ), .A2(\shift[0] ), .ZN(new_n287_));
  NAND2_X1   g0024(.A1(new_n266_), .A2(\a[66] ), .ZN(new_n288_));
  AOI21_X1   g0025(.A1(new_n288_), .A2(new_n287_), .B(new_n275_), .ZN(new_n289_));
  NAND2_X1   g0026(.A1(new_n266_), .A2(\a[68] ), .ZN(new_n290_));
  NAND2_X1   g0027(.A1(\a[67] ), .A2(\shift[0] ), .ZN(new_n291_));
  AOI21_X1   g0028(.A1(new_n290_), .A2(new_n291_), .B(\shift[1] ), .ZN(new_n292_));
  INV_X1     g0029(.I(\shift[3] ), .ZN(new_n293_));
  NOR2_X1    g0030(.A1(new_n283_), .A2(new_n293_), .ZN(new_n294_));
  OAI21_X1   g0031(.A1(new_n289_), .A2(new_n292_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1   g0032(.A1(\a[69] ), .A2(\shift[0] ), .ZN(new_n296_));
  NAND2_X1   g0033(.A1(new_n266_), .A2(\a[70] ), .ZN(new_n297_));
  AOI21_X1   g0034(.A1(new_n297_), .A2(new_n296_), .B(new_n275_), .ZN(new_n298_));
  NAND2_X1   g0035(.A1(new_n266_), .A2(\a[72] ), .ZN(new_n299_));
  NAND2_X1   g0036(.A1(\a[71] ), .A2(\shift[0] ), .ZN(new_n300_));
  AOI21_X1   g0037(.A1(new_n299_), .A2(new_n300_), .B(\shift[1] ), .ZN(new_n301_));
  NOR2_X1    g0038(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1    g0039(.A1(new_n293_), .A2(\shift[2] ), .ZN(new_n303_));
  INV_X1     g0040(.I(new_n303_), .ZN(new_n304_));
  OAI21_X1   g0041(.A1(new_n302_), .A2(new_n304_), .B(new_n295_), .ZN(new_n305_));
  INV_X1     g0042(.I(\shift[4] ), .ZN(new_n306_));
  INV_X1     g0043(.I(\shift[5] ), .ZN(new_n307_));
  NOR2_X1    g0044(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1   g0045(.A1(new_n286_), .A2(new_n305_), .B(new_n308_), .ZN(new_n309_));
  NAND3_X1   g0046(.A1(\a[93] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n310_));
  NAND3_X1   g0047(.A1(new_n266_), .A2(\a[94] ), .A3(\shift[1] ), .ZN(new_n311_));
  NAND2_X1   g0048(.A1(new_n311_), .A2(new_n310_), .ZN(new_n312_));
  NAND2_X1   g0049(.A1(new_n266_), .A2(\a[96] ), .ZN(new_n313_));
  NAND2_X1   g0050(.A1(\a[95] ), .A2(\shift[0] ), .ZN(new_n314_));
  AOI21_X1   g0051(.A1(new_n313_), .A2(new_n314_), .B(\shift[1] ), .ZN(new_n315_));
  NOR2_X1    g0052(.A1(new_n315_), .A2(new_n312_), .ZN(new_n316_));
  NAND2_X1   g0053(.A1(\a[89] ), .A2(\shift[0] ), .ZN(new_n317_));
  NAND2_X1   g0054(.A1(new_n266_), .A2(\a[90] ), .ZN(new_n318_));
  AOI21_X1   g0055(.A1(new_n318_), .A2(new_n317_), .B(new_n275_), .ZN(new_n319_));
  NAND2_X1   g0056(.A1(new_n266_), .A2(\a[92] ), .ZN(new_n320_));
  NAND2_X1   g0057(.A1(\a[91] ), .A2(\shift[0] ), .ZN(new_n321_));
  AOI21_X1   g0058(.A1(new_n320_), .A2(new_n321_), .B(\shift[1] ), .ZN(new_n322_));
  NOR2_X1    g0059(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  OAI22_X1   g0060(.A1(new_n285_), .A2(new_n323_), .B1(new_n316_), .B2(new_n274_), .ZN(new_n324_));
  NAND3_X1   g0061(.A1(\a[81] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n325_));
  NAND3_X1   g0062(.A1(new_n266_), .A2(\a[82] ), .A3(\shift[1] ), .ZN(new_n326_));
  NAND2_X1   g0063(.A1(new_n326_), .A2(new_n325_), .ZN(new_n327_));
  NAND2_X1   g0064(.A1(new_n266_), .A2(\a[84] ), .ZN(new_n328_));
  NAND2_X1   g0065(.A1(\a[83] ), .A2(\shift[0] ), .ZN(new_n329_));
  AOI21_X1   g0066(.A1(new_n328_), .A2(new_n329_), .B(\shift[1] ), .ZN(new_n330_));
  OAI21_X1   g0067(.A1(new_n330_), .A2(new_n327_), .B(new_n294_), .ZN(new_n331_));
  NAND2_X1   g0068(.A1(\a[85] ), .A2(\shift[0] ), .ZN(new_n332_));
  NAND2_X1   g0069(.A1(new_n266_), .A2(\a[86] ), .ZN(new_n333_));
  AOI21_X1   g0070(.A1(new_n333_), .A2(new_n332_), .B(new_n275_), .ZN(new_n334_));
  NAND2_X1   g0071(.A1(new_n266_), .A2(\a[88] ), .ZN(new_n335_));
  NAND2_X1   g0072(.A1(\a[87] ), .A2(\shift[0] ), .ZN(new_n336_));
  AOI21_X1   g0073(.A1(new_n335_), .A2(new_n336_), .B(\shift[1] ), .ZN(new_n337_));
  OAI21_X1   g0074(.A1(new_n334_), .A2(new_n337_), .B(new_n303_), .ZN(new_n338_));
  NAND2_X1   g0075(.A1(new_n338_), .A2(new_n331_), .ZN(new_n339_));
  NOR2_X1    g0076(.A1(new_n307_), .A2(\shift[4] ), .ZN(new_n340_));
  OAI21_X1   g0077(.A1(new_n324_), .A2(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1   g0078(.A1(new_n309_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1   g0079(.A1(\a[125] ), .A2(\shift[0] ), .ZN(new_n343_));
  NAND2_X1   g0080(.A1(new_n266_), .A2(\a[126] ), .ZN(new_n344_));
  AOI21_X1   g0081(.A1(new_n344_), .A2(new_n343_), .B(new_n275_), .ZN(new_n345_));
  NAND2_X1   g0082(.A1(new_n266_), .A2(\a[0] ), .ZN(new_n346_));
  NAND2_X1   g0083(.A1(\a[127] ), .A2(\shift[0] ), .ZN(new_n347_));
  AOI21_X1   g0084(.A1(new_n346_), .A2(new_n347_), .B(\shift[1] ), .ZN(new_n348_));
  OAI21_X1   g0085(.A1(new_n345_), .A2(new_n348_), .B(new_n273_), .ZN(new_n349_));
  NAND3_X1   g0086(.A1(\a[121] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n350_));
  NAND3_X1   g0087(.A1(new_n266_), .A2(\a[122] ), .A3(\shift[1] ), .ZN(new_n351_));
  NAND2_X1   g0088(.A1(new_n351_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1   g0089(.A1(new_n266_), .A2(\a[124] ), .ZN(new_n353_));
  NAND2_X1   g0090(.A1(\a[123] ), .A2(\shift[0] ), .ZN(new_n354_));
  AOI21_X1   g0091(.A1(new_n353_), .A2(new_n354_), .B(\shift[1] ), .ZN(new_n355_));
  OAI21_X1   g0092(.A1(new_n355_), .A2(new_n352_), .B(new_n284_), .ZN(new_n356_));
  NAND2_X1   g0093(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1   g0094(.A1(\a[113] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n358_));
  NAND3_X1   g0095(.A1(new_n266_), .A2(\a[114] ), .A3(\shift[1] ), .ZN(new_n359_));
  NAND2_X1   g0096(.A1(new_n359_), .A2(new_n358_), .ZN(new_n360_));
  NAND2_X1   g0097(.A1(new_n266_), .A2(\a[116] ), .ZN(new_n361_));
  NAND2_X1   g0098(.A1(\a[115] ), .A2(\shift[0] ), .ZN(new_n362_));
  AOI21_X1   g0099(.A1(new_n361_), .A2(new_n362_), .B(\shift[1] ), .ZN(new_n363_));
  OAI21_X1   g0100(.A1(new_n363_), .A2(new_n360_), .B(new_n294_), .ZN(new_n364_));
  NAND3_X1   g0101(.A1(\a[117] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n365_));
  NAND3_X1   g0102(.A1(new_n266_), .A2(\a[118] ), .A3(\shift[1] ), .ZN(new_n366_));
  NAND2_X1   g0103(.A1(new_n366_), .A2(new_n365_), .ZN(new_n367_));
  NAND2_X1   g0104(.A1(new_n266_), .A2(\a[120] ), .ZN(new_n368_));
  NAND2_X1   g0105(.A1(\a[119] ), .A2(\shift[0] ), .ZN(new_n369_));
  AOI21_X1   g0106(.A1(new_n368_), .A2(new_n369_), .B(\shift[1] ), .ZN(new_n370_));
  OAI21_X1   g0107(.A1(new_n370_), .A2(new_n367_), .B(new_n303_), .ZN(new_n371_));
  NAND2_X1   g0108(.A1(new_n364_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1    g0109(.A1(\shift[4] ), .A2(\shift[5] ), .ZN(new_n373_));
  OAI21_X1   g0110(.A1(new_n357_), .A2(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NAND3_X1   g0111(.A1(\a[109] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n375_));
  NAND3_X1   g0112(.A1(new_n266_), .A2(\a[110] ), .A3(\shift[1] ), .ZN(new_n376_));
  NAND2_X1   g0113(.A1(new_n376_), .A2(new_n375_), .ZN(new_n377_));
  NAND2_X1   g0114(.A1(new_n266_), .A2(\a[112] ), .ZN(new_n378_));
  NAND2_X1   g0115(.A1(\a[111] ), .A2(\shift[0] ), .ZN(new_n379_));
  AOI21_X1   g0116(.A1(new_n378_), .A2(new_n379_), .B(\shift[1] ), .ZN(new_n380_));
  OAI21_X1   g0117(.A1(new_n380_), .A2(new_n377_), .B(new_n273_), .ZN(new_n381_));
  NAND3_X1   g0118(.A1(\a[105] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n382_));
  NAND3_X1   g0119(.A1(new_n266_), .A2(\a[106] ), .A3(\shift[1] ), .ZN(new_n383_));
  NAND2_X1   g0120(.A1(new_n383_), .A2(new_n382_), .ZN(new_n384_));
  NAND2_X1   g0121(.A1(new_n266_), .A2(\a[108] ), .ZN(new_n385_));
  NAND2_X1   g0122(.A1(\a[107] ), .A2(\shift[0] ), .ZN(new_n386_));
  AOI21_X1   g0123(.A1(new_n385_), .A2(new_n386_), .B(\shift[1] ), .ZN(new_n387_));
  OAI21_X1   g0124(.A1(new_n387_), .A2(new_n384_), .B(new_n284_), .ZN(new_n388_));
  NAND2_X1   g0125(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1   g0126(.A1(\a[97] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n390_));
  NAND3_X1   g0127(.A1(new_n266_), .A2(\a[98] ), .A3(\shift[1] ), .ZN(new_n391_));
  NAND2_X1   g0128(.A1(new_n391_), .A2(new_n390_), .ZN(new_n392_));
  NAND2_X1   g0129(.A1(new_n266_), .A2(\a[100] ), .ZN(new_n393_));
  NAND2_X1   g0130(.A1(\a[99] ), .A2(\shift[0] ), .ZN(new_n394_));
  AOI21_X1   g0131(.A1(new_n393_), .A2(new_n394_), .B(\shift[1] ), .ZN(new_n395_));
  OAI21_X1   g0132(.A1(new_n395_), .A2(new_n392_), .B(new_n294_), .ZN(new_n396_));
  NAND3_X1   g0133(.A1(\a[101] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n397_));
  NAND3_X1   g0134(.A1(new_n266_), .A2(\a[102] ), .A3(\shift[1] ), .ZN(new_n398_));
  NAND2_X1   g0135(.A1(new_n398_), .A2(new_n397_), .ZN(new_n399_));
  NAND2_X1   g0136(.A1(new_n266_), .A2(\a[104] ), .ZN(new_n400_));
  NAND2_X1   g0137(.A1(\a[103] ), .A2(\shift[0] ), .ZN(new_n401_));
  AOI21_X1   g0138(.A1(new_n400_), .A2(new_n401_), .B(\shift[1] ), .ZN(new_n402_));
  OAI21_X1   g0139(.A1(new_n402_), .A2(new_n399_), .B(new_n303_), .ZN(new_n403_));
  NAND2_X1   g0140(.A1(new_n396_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1    g0141(.A1(new_n306_), .A2(\shift[5] ), .ZN(new_n405_));
  OAI21_X1   g0142(.A1(new_n389_), .A2(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1   g0143(.A1(new_n374_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1   g0144(.A1(new_n342_), .A2(new_n407_), .B(new_n264_), .ZN(new_n408_));
  NAND3_X1   g0145(.A1(\a[13] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n409_));
  NAND3_X1   g0146(.A1(new_n266_), .A2(\a[14] ), .A3(\shift[1] ), .ZN(new_n410_));
  NAND2_X1   g0147(.A1(new_n410_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1   g0148(.A1(new_n266_), .A2(\a[16] ), .ZN(new_n412_));
  NAND2_X1   g0149(.A1(\a[15] ), .A2(\shift[0] ), .ZN(new_n413_));
  AOI21_X1   g0150(.A1(new_n412_), .A2(new_n413_), .B(\shift[1] ), .ZN(new_n414_));
  OAI21_X1   g0151(.A1(new_n414_), .A2(new_n411_), .B(new_n273_), .ZN(new_n415_));
  NAND3_X1   g0152(.A1(\a[9] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n416_));
  NAND3_X1   g0153(.A1(new_n266_), .A2(\a[10] ), .A3(\shift[1] ), .ZN(new_n417_));
  NAND2_X1   g0154(.A1(new_n417_), .A2(new_n416_), .ZN(new_n418_));
  NAND2_X1   g0155(.A1(new_n266_), .A2(\a[12] ), .ZN(new_n419_));
  NAND2_X1   g0156(.A1(\a[11] ), .A2(\shift[0] ), .ZN(new_n420_));
  AOI21_X1   g0157(.A1(new_n419_), .A2(new_n420_), .B(\shift[1] ), .ZN(new_n421_));
  OAI21_X1   g0158(.A1(new_n421_), .A2(new_n418_), .B(new_n284_), .ZN(new_n422_));
  NAND2_X1   g0159(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1   g0160(.A1(\a[1] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n424_));
  NAND3_X1   g0161(.A1(new_n266_), .A2(\a[2] ), .A3(\shift[1] ), .ZN(new_n425_));
  NAND2_X1   g0162(.A1(new_n425_), .A2(new_n424_), .ZN(new_n426_));
  NAND2_X1   g0163(.A1(new_n266_), .A2(\a[4] ), .ZN(new_n427_));
  NAND2_X1   g0164(.A1(\a[3] ), .A2(\shift[0] ), .ZN(new_n428_));
  AOI21_X1   g0165(.A1(new_n427_), .A2(new_n428_), .B(\shift[1] ), .ZN(new_n429_));
  OAI21_X1   g0166(.A1(new_n429_), .A2(new_n426_), .B(new_n294_), .ZN(new_n430_));
  NAND3_X1   g0167(.A1(\a[5] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n431_));
  NAND3_X1   g0168(.A1(new_n266_), .A2(\a[6] ), .A3(\shift[1] ), .ZN(new_n432_));
  NAND2_X1   g0169(.A1(new_n432_), .A2(new_n431_), .ZN(new_n433_));
  NAND2_X1   g0170(.A1(new_n266_), .A2(\a[8] ), .ZN(new_n434_));
  NAND2_X1   g0171(.A1(\a[7] ), .A2(\shift[0] ), .ZN(new_n435_));
  AOI21_X1   g0172(.A1(new_n434_), .A2(new_n435_), .B(\shift[1] ), .ZN(new_n436_));
  OAI21_X1   g0173(.A1(new_n436_), .A2(new_n433_), .B(new_n303_), .ZN(new_n437_));
  NAND2_X1   g0174(.A1(new_n430_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1   g0175(.A1(new_n423_), .A2(new_n438_), .B(new_n308_), .ZN(new_n439_));
  NAND3_X1   g0176(.A1(\a[29] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n440_));
  NAND3_X1   g0177(.A1(new_n266_), .A2(\a[30] ), .A3(\shift[1] ), .ZN(new_n441_));
  NAND2_X1   g0178(.A1(new_n441_), .A2(new_n440_), .ZN(new_n442_));
  NAND2_X1   g0179(.A1(new_n266_), .A2(\a[32] ), .ZN(new_n443_));
  NAND2_X1   g0180(.A1(\a[31] ), .A2(\shift[0] ), .ZN(new_n444_));
  AOI21_X1   g0181(.A1(new_n443_), .A2(new_n444_), .B(\shift[1] ), .ZN(new_n445_));
  OAI21_X1   g0182(.A1(new_n445_), .A2(new_n442_), .B(new_n273_), .ZN(new_n446_));
  NAND2_X1   g0183(.A1(\a[25] ), .A2(\shift[0] ), .ZN(new_n447_));
  NAND2_X1   g0184(.A1(new_n266_), .A2(\a[26] ), .ZN(new_n448_));
  AOI21_X1   g0185(.A1(new_n448_), .A2(new_n447_), .B(new_n275_), .ZN(new_n449_));
  NAND2_X1   g0186(.A1(new_n266_), .A2(\a[28] ), .ZN(new_n450_));
  NAND2_X1   g0187(.A1(\a[27] ), .A2(\shift[0] ), .ZN(new_n451_));
  AOI21_X1   g0188(.A1(new_n450_), .A2(new_n451_), .B(\shift[1] ), .ZN(new_n452_));
  OAI21_X1   g0189(.A1(new_n449_), .A2(new_n452_), .B(new_n284_), .ZN(new_n453_));
  NAND2_X1   g0190(.A1(new_n453_), .A2(new_n446_), .ZN(new_n454_));
  NAND3_X1   g0191(.A1(\a[17] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n455_));
  NAND3_X1   g0192(.A1(new_n266_), .A2(\a[18] ), .A3(\shift[1] ), .ZN(new_n456_));
  NAND2_X1   g0193(.A1(new_n456_), .A2(new_n455_), .ZN(new_n457_));
  NAND2_X1   g0194(.A1(new_n266_), .A2(\a[20] ), .ZN(new_n458_));
  NAND2_X1   g0195(.A1(\a[19] ), .A2(\shift[0] ), .ZN(new_n459_));
  AOI21_X1   g0196(.A1(new_n458_), .A2(new_n459_), .B(\shift[1] ), .ZN(new_n460_));
  OAI21_X1   g0197(.A1(new_n460_), .A2(new_n457_), .B(new_n294_), .ZN(new_n461_));
  NAND3_X1   g0198(.A1(\a[21] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n462_));
  NAND3_X1   g0199(.A1(new_n266_), .A2(\a[22] ), .A3(\shift[1] ), .ZN(new_n463_));
  NAND2_X1   g0200(.A1(new_n463_), .A2(new_n462_), .ZN(new_n464_));
  NAND2_X1   g0201(.A1(new_n266_), .A2(\a[24] ), .ZN(new_n465_));
  NAND2_X1   g0202(.A1(\a[23] ), .A2(\shift[0] ), .ZN(new_n466_));
  AOI21_X1   g0203(.A1(new_n465_), .A2(new_n466_), .B(\shift[1] ), .ZN(new_n467_));
  OAI21_X1   g0204(.A1(new_n467_), .A2(new_n464_), .B(new_n303_), .ZN(new_n468_));
  NAND2_X1   g0205(.A1(new_n461_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1   g0206(.A1(new_n454_), .A2(new_n469_), .B(new_n340_), .ZN(new_n470_));
  NAND2_X1   g0207(.A1(new_n439_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1   g0208(.A1(\a[61] ), .A2(\shift[0] ), .ZN(new_n472_));
  NAND2_X1   g0209(.A1(new_n266_), .A2(\a[62] ), .ZN(new_n473_));
  AOI21_X1   g0210(.A1(new_n473_), .A2(new_n472_), .B(new_n275_), .ZN(new_n474_));
  NAND2_X1   g0211(.A1(new_n266_), .A2(\a[64] ), .ZN(new_n475_));
  NAND2_X1   g0212(.A1(\a[63] ), .A2(\shift[0] ), .ZN(new_n476_));
  AOI21_X1   g0213(.A1(new_n475_), .A2(new_n476_), .B(\shift[1] ), .ZN(new_n477_));
  NOR2_X1    g0214(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1   g0215(.A1(\a[57] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n479_));
  NAND3_X1   g0216(.A1(new_n266_), .A2(\a[58] ), .A3(\shift[1] ), .ZN(new_n480_));
  NAND2_X1   g0217(.A1(new_n480_), .A2(new_n479_), .ZN(new_n481_));
  NAND2_X1   g0218(.A1(new_n266_), .A2(\a[60] ), .ZN(new_n482_));
  NAND2_X1   g0219(.A1(\a[59] ), .A2(\shift[0] ), .ZN(new_n483_));
  AOI21_X1   g0220(.A1(new_n482_), .A2(new_n483_), .B(\shift[1] ), .ZN(new_n484_));
  NOR2_X1    g0221(.A1(new_n484_), .A2(new_n481_), .ZN(new_n485_));
  OAI22_X1   g0222(.A1(new_n274_), .A2(new_n478_), .B1(new_n485_), .B2(new_n285_), .ZN(new_n486_));
  NAND2_X1   g0223(.A1(\a[49] ), .A2(\shift[0] ), .ZN(new_n487_));
  NAND2_X1   g0224(.A1(new_n266_), .A2(\a[50] ), .ZN(new_n488_));
  AOI21_X1   g0225(.A1(new_n488_), .A2(new_n487_), .B(new_n275_), .ZN(new_n489_));
  NAND2_X1   g0226(.A1(new_n266_), .A2(\a[52] ), .ZN(new_n490_));
  NAND2_X1   g0227(.A1(\a[51] ), .A2(\shift[0] ), .ZN(new_n491_));
  AOI21_X1   g0228(.A1(new_n490_), .A2(new_n491_), .B(\shift[1] ), .ZN(new_n492_));
  OAI21_X1   g0229(.A1(new_n489_), .A2(new_n492_), .B(new_n294_), .ZN(new_n493_));
  NAND2_X1   g0230(.A1(\a[53] ), .A2(\shift[0] ), .ZN(new_n494_));
  NAND2_X1   g0231(.A1(new_n266_), .A2(\a[54] ), .ZN(new_n495_));
  AOI21_X1   g0232(.A1(new_n495_), .A2(new_n494_), .B(new_n275_), .ZN(new_n496_));
  NAND2_X1   g0233(.A1(new_n266_), .A2(\a[56] ), .ZN(new_n497_));
  NAND2_X1   g0234(.A1(\a[55] ), .A2(\shift[0] ), .ZN(new_n498_));
  AOI21_X1   g0235(.A1(new_n497_), .A2(new_n498_), .B(\shift[1] ), .ZN(new_n499_));
  OAI21_X1   g0236(.A1(new_n496_), .A2(new_n499_), .B(new_n303_), .ZN(new_n500_));
  NAND2_X1   g0237(.A1(new_n493_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1   g0238(.A1(new_n486_), .A2(new_n501_), .B(new_n373_), .ZN(new_n502_));
  NAND2_X1   g0239(.A1(\a[45] ), .A2(\shift[0] ), .ZN(new_n503_));
  NAND2_X1   g0240(.A1(new_n266_), .A2(\a[46] ), .ZN(new_n504_));
  AOI21_X1   g0241(.A1(new_n504_), .A2(new_n503_), .B(new_n275_), .ZN(new_n505_));
  NAND2_X1   g0242(.A1(new_n266_), .A2(\a[48] ), .ZN(new_n506_));
  NAND2_X1   g0243(.A1(\a[47] ), .A2(\shift[0] ), .ZN(new_n507_));
  AOI21_X1   g0244(.A1(new_n506_), .A2(new_n507_), .B(\shift[1] ), .ZN(new_n508_));
  OAI21_X1   g0245(.A1(new_n505_), .A2(new_n508_), .B(new_n273_), .ZN(new_n509_));
  NAND3_X1   g0246(.A1(\a[41] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n510_));
  NAND3_X1   g0247(.A1(new_n266_), .A2(\a[42] ), .A3(\shift[1] ), .ZN(new_n511_));
  NAND2_X1   g0248(.A1(new_n511_), .A2(new_n510_), .ZN(new_n512_));
  NAND2_X1   g0249(.A1(new_n266_), .A2(\a[44] ), .ZN(new_n513_));
  NAND2_X1   g0250(.A1(\a[43] ), .A2(\shift[0] ), .ZN(new_n514_));
  AOI21_X1   g0251(.A1(new_n513_), .A2(new_n514_), .B(\shift[1] ), .ZN(new_n515_));
  OAI21_X1   g0252(.A1(new_n515_), .A2(new_n512_), .B(new_n284_), .ZN(new_n516_));
  NAND2_X1   g0253(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1   g0254(.A1(\a[33] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n518_));
  NAND3_X1   g0255(.A1(new_n266_), .A2(\a[34] ), .A3(\shift[1] ), .ZN(new_n519_));
  NAND2_X1   g0256(.A1(new_n519_), .A2(new_n518_), .ZN(new_n520_));
  NAND2_X1   g0257(.A1(new_n266_), .A2(\a[36] ), .ZN(new_n521_));
  NAND2_X1   g0258(.A1(\a[35] ), .A2(\shift[0] ), .ZN(new_n522_));
  AOI21_X1   g0259(.A1(new_n521_), .A2(new_n522_), .B(\shift[1] ), .ZN(new_n523_));
  OAI21_X1   g0260(.A1(new_n523_), .A2(new_n520_), .B(new_n294_), .ZN(new_n524_));
  NAND2_X1   g0261(.A1(new_n266_), .A2(\a[40] ), .ZN(new_n525_));
  NAND3_X1   g0262(.A1(\a[37] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n526_));
  OAI21_X1   g0263(.A1(new_n525_), .A2(\shift[1] ), .B(new_n526_), .ZN(new_n527_));
  NAND3_X1   g0264(.A1(new_n275_), .A2(\a[39] ), .A3(\shift[0] ), .ZN(new_n528_));
  NAND3_X1   g0265(.A1(new_n266_), .A2(\a[38] ), .A3(\shift[1] ), .ZN(new_n529_));
  NAND2_X1   g0266(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1   g0267(.A1(new_n530_), .A2(new_n527_), .B(new_n303_), .ZN(new_n531_));
  NAND2_X1   g0268(.A1(new_n531_), .A2(new_n524_), .ZN(new_n532_));
  OAI21_X1   g0269(.A1(new_n517_), .A2(new_n532_), .B(new_n405_), .ZN(new_n533_));
  NAND2_X1   g0270(.A1(new_n502_), .A2(new_n533_), .ZN(new_n534_));
  OAI21_X1   g0271(.A1(new_n471_), .A2(new_n534_), .B(\shift[6] ), .ZN(new_n535_));
  NAND2_X1   g0272(.A1(new_n408_), .A2(new_n535_), .ZN(\result[0] ));
  INV_X1     g0273(.I(new_n308_), .ZN(new_n537_));
  INV_X1     g0274(.I(\a[81] ), .ZN(new_n538_));
  NOR3_X1    g0275(.A1(new_n538_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n539_));
  INV_X1     g0276(.I(\a[78] ), .ZN(new_n540_));
  NOR3_X1    g0277(.A1(new_n540_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n541_));
  NAND2_X1   g0278(.A1(\a[80] ), .A2(\shift[0] ), .ZN(new_n542_));
  NOR2_X1    g0279(.A1(new_n542_), .A2(\shift[1] ), .ZN(new_n543_));
  INV_X1     g0280(.I(\a[79] ), .ZN(new_n544_));
  NOR3_X1    g0281(.A1(new_n544_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n545_));
  NOR4_X1    g0282(.A1(new_n541_), .A2(new_n543_), .A3(new_n545_), .A4(new_n539_), .ZN(new_n546_));
  INV_X1     g0283(.I(\a[77] ), .ZN(new_n547_));
  NOR3_X1    g0284(.A1(new_n547_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n548_));
  INV_X1     g0285(.I(\a[74] ), .ZN(new_n549_));
  NOR3_X1    g0286(.A1(new_n549_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n550_));
  NAND2_X1   g0287(.A1(\a[76] ), .A2(\shift[0] ), .ZN(new_n551_));
  NOR2_X1    g0288(.A1(new_n551_), .A2(\shift[1] ), .ZN(new_n552_));
  INV_X1     g0289(.I(\a[75] ), .ZN(new_n553_));
  NOR3_X1    g0290(.A1(new_n553_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n554_));
  NOR4_X1    g0291(.A1(new_n550_), .A2(new_n552_), .A3(new_n554_), .A4(new_n548_), .ZN(new_n555_));
  OAI22_X1   g0292(.A1(new_n274_), .A2(new_n546_), .B1(new_n555_), .B2(new_n285_), .ZN(new_n556_));
  INV_X1     g0293(.I(new_n294_), .ZN(new_n557_));
  INV_X1     g0294(.I(\a[69] ), .ZN(new_n558_));
  NOR3_X1    g0295(.A1(new_n558_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n559_));
  INV_X1     g0296(.I(\a[66] ), .ZN(new_n560_));
  NOR3_X1    g0297(.A1(new_n560_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n561_));
  NAND2_X1   g0298(.A1(\a[68] ), .A2(\shift[0] ), .ZN(new_n562_));
  NOR2_X1    g0299(.A1(new_n562_), .A2(\shift[1] ), .ZN(new_n563_));
  INV_X1     g0300(.I(\a[67] ), .ZN(new_n564_));
  NOR3_X1    g0301(.A1(new_n564_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n565_));
  NOR4_X1    g0302(.A1(new_n561_), .A2(new_n563_), .A3(new_n565_), .A4(new_n559_), .ZN(new_n566_));
  INV_X1     g0303(.I(\a[73] ), .ZN(new_n567_));
  NOR3_X1    g0304(.A1(new_n567_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n568_));
  INV_X1     g0305(.I(\a[70] ), .ZN(new_n569_));
  NOR3_X1    g0306(.A1(new_n569_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n570_));
  NAND2_X1   g0307(.A1(\a[72] ), .A2(\shift[0] ), .ZN(new_n571_));
  NOR2_X1    g0308(.A1(new_n571_), .A2(\shift[1] ), .ZN(new_n572_));
  INV_X1     g0309(.I(\a[71] ), .ZN(new_n573_));
  NOR3_X1    g0310(.A1(new_n573_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n574_));
  NOR4_X1    g0311(.A1(new_n570_), .A2(new_n572_), .A3(new_n574_), .A4(new_n568_), .ZN(new_n575_));
  OAI22_X1   g0312(.A1(new_n557_), .A2(new_n566_), .B1(new_n575_), .B2(new_n304_), .ZN(new_n576_));
  NOR2_X1    g0313(.A1(new_n556_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1     g0314(.I(\a[97] ), .ZN(new_n578_));
  NOR3_X1    g0315(.A1(new_n578_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n579_));
  INV_X1     g0316(.I(\a[94] ), .ZN(new_n580_));
  NOR3_X1    g0317(.A1(new_n580_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n581_));
  INV_X1     g0318(.I(\a[96] ), .ZN(new_n582_));
  NOR3_X1    g0319(.A1(new_n582_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n583_));
  INV_X1     g0320(.I(\a[95] ), .ZN(new_n584_));
  NOR3_X1    g0321(.A1(new_n584_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n585_));
  NOR4_X1    g0322(.A1(new_n581_), .A2(new_n583_), .A3(new_n585_), .A4(new_n579_), .ZN(new_n586_));
  INV_X1     g0323(.I(\a[93] ), .ZN(new_n587_));
  NOR3_X1    g0324(.A1(new_n587_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n588_));
  INV_X1     g0325(.I(\a[90] ), .ZN(new_n589_));
  NOR3_X1    g0326(.A1(new_n589_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n590_));
  INV_X1     g0327(.I(\a[92] ), .ZN(new_n591_));
  NOR3_X1    g0328(.A1(new_n591_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n592_));
  INV_X1     g0329(.I(\a[91] ), .ZN(new_n593_));
  NOR3_X1    g0330(.A1(new_n593_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n594_));
  NOR4_X1    g0331(.A1(new_n590_), .A2(new_n592_), .A3(new_n594_), .A4(new_n588_), .ZN(new_n595_));
  OAI22_X1   g0332(.A1(new_n274_), .A2(new_n586_), .B1(new_n595_), .B2(new_n285_), .ZN(new_n596_));
  INV_X1     g0333(.I(\a[85] ), .ZN(new_n597_));
  NOR3_X1    g0334(.A1(new_n597_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n598_));
  INV_X1     g0335(.I(\a[82] ), .ZN(new_n599_));
  NOR3_X1    g0336(.A1(new_n599_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n600_));
  INV_X1     g0337(.I(\a[84] ), .ZN(new_n601_));
  NOR3_X1    g0338(.A1(new_n601_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n602_));
  INV_X1     g0339(.I(\a[83] ), .ZN(new_n603_));
  NOR3_X1    g0340(.A1(new_n603_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n604_));
  NOR4_X1    g0341(.A1(new_n600_), .A2(new_n602_), .A3(new_n604_), .A4(new_n598_), .ZN(new_n605_));
  INV_X1     g0342(.I(\a[89] ), .ZN(new_n606_));
  NOR3_X1    g0343(.A1(new_n606_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n607_));
  INV_X1     g0344(.I(\a[86] ), .ZN(new_n608_));
  NOR3_X1    g0345(.A1(new_n608_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n609_));
  NAND2_X1   g0346(.A1(\a[88] ), .A2(\shift[0] ), .ZN(new_n610_));
  NOR2_X1    g0347(.A1(new_n610_), .A2(\shift[1] ), .ZN(new_n611_));
  INV_X1     g0348(.I(\a[87] ), .ZN(new_n612_));
  NOR3_X1    g0349(.A1(new_n612_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n613_));
  NOR4_X1    g0350(.A1(new_n609_), .A2(new_n611_), .A3(new_n613_), .A4(new_n607_), .ZN(new_n614_));
  OAI22_X1   g0351(.A1(new_n557_), .A2(new_n605_), .B1(new_n614_), .B2(new_n304_), .ZN(new_n615_));
  OAI21_X1   g0352(.A1(new_n596_), .A2(new_n615_), .B(new_n340_), .ZN(new_n616_));
  OAI21_X1   g0353(.A1(new_n537_), .A2(new_n577_), .B(new_n616_), .ZN(new_n617_));
  INV_X1     g0354(.I(\a[1] ), .ZN(new_n618_));
  NOR3_X1    g0355(.A1(new_n618_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n619_));
  INV_X1     g0356(.I(\a[126] ), .ZN(new_n620_));
  NOR3_X1    g0357(.A1(new_n620_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n621_));
  INV_X1     g0358(.I(\a[0] ), .ZN(new_n622_));
  NOR3_X1    g0359(.A1(new_n622_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n623_));
  INV_X1     g0360(.I(\a[127] ), .ZN(new_n624_));
  NOR3_X1    g0361(.A1(new_n624_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n625_));
  NOR4_X1    g0362(.A1(new_n621_), .A2(new_n623_), .A3(new_n625_), .A4(new_n619_), .ZN(new_n626_));
  INV_X1     g0363(.I(\a[125] ), .ZN(new_n627_));
  NOR3_X1    g0364(.A1(new_n627_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n628_));
  INV_X1     g0365(.I(\a[122] ), .ZN(new_n629_));
  NOR3_X1    g0366(.A1(new_n629_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n630_));
  INV_X1     g0367(.I(\a[124] ), .ZN(new_n631_));
  NOR3_X1    g0368(.A1(new_n631_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n632_));
  INV_X1     g0369(.I(\a[123] ), .ZN(new_n633_));
  NOR3_X1    g0370(.A1(new_n633_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n634_));
  NOR4_X1    g0371(.A1(new_n630_), .A2(new_n632_), .A3(new_n634_), .A4(new_n628_), .ZN(new_n635_));
  OAI22_X1   g0372(.A1(new_n274_), .A2(new_n626_), .B1(new_n635_), .B2(new_n285_), .ZN(new_n636_));
  INV_X1     g0373(.I(\a[117] ), .ZN(new_n637_));
  NOR3_X1    g0374(.A1(new_n637_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n638_));
  INV_X1     g0375(.I(\a[114] ), .ZN(new_n639_));
  NOR3_X1    g0376(.A1(new_n639_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n640_));
  INV_X1     g0377(.I(\a[116] ), .ZN(new_n641_));
  NOR3_X1    g0378(.A1(new_n641_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n642_));
  INV_X1     g0379(.I(\a[115] ), .ZN(new_n643_));
  NOR3_X1    g0380(.A1(new_n643_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n644_));
  NOR4_X1    g0381(.A1(new_n640_), .A2(new_n642_), .A3(new_n644_), .A4(new_n638_), .ZN(new_n645_));
  INV_X1     g0382(.I(\a[121] ), .ZN(new_n646_));
  NOR3_X1    g0383(.A1(new_n646_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n647_));
  INV_X1     g0384(.I(\a[118] ), .ZN(new_n648_));
  NOR3_X1    g0385(.A1(new_n648_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n649_));
  INV_X1     g0386(.I(\a[120] ), .ZN(new_n650_));
  NOR3_X1    g0387(.A1(new_n650_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n651_));
  INV_X1     g0388(.I(\a[119] ), .ZN(new_n652_));
  NOR3_X1    g0389(.A1(new_n652_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n653_));
  NOR4_X1    g0390(.A1(new_n649_), .A2(new_n651_), .A3(new_n653_), .A4(new_n647_), .ZN(new_n654_));
  OAI22_X1   g0391(.A1(new_n557_), .A2(new_n645_), .B1(new_n654_), .B2(new_n304_), .ZN(new_n655_));
  OAI21_X1   g0392(.A1(new_n636_), .A2(new_n655_), .B(new_n373_), .ZN(new_n656_));
  INV_X1     g0393(.I(\a[113] ), .ZN(new_n657_));
  NOR3_X1    g0394(.A1(new_n657_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n658_));
  INV_X1     g0395(.I(\a[110] ), .ZN(new_n659_));
  NOR3_X1    g0396(.A1(new_n659_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n660_));
  INV_X1     g0397(.I(\a[112] ), .ZN(new_n661_));
  NOR3_X1    g0398(.A1(new_n661_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n662_));
  INV_X1     g0399(.I(\a[111] ), .ZN(new_n663_));
  NOR3_X1    g0400(.A1(new_n663_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n664_));
  NOR4_X1    g0401(.A1(new_n660_), .A2(new_n662_), .A3(new_n664_), .A4(new_n658_), .ZN(new_n665_));
  INV_X1     g0402(.I(\a[109] ), .ZN(new_n666_));
  NOR3_X1    g0403(.A1(new_n666_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n667_));
  INV_X1     g0404(.I(\a[106] ), .ZN(new_n668_));
  NOR3_X1    g0405(.A1(new_n668_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n669_));
  INV_X1     g0406(.I(\a[108] ), .ZN(new_n670_));
  NOR3_X1    g0407(.A1(new_n670_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n671_));
  INV_X1     g0408(.I(\a[107] ), .ZN(new_n672_));
  NOR3_X1    g0409(.A1(new_n672_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n673_));
  NOR4_X1    g0410(.A1(new_n669_), .A2(new_n671_), .A3(new_n673_), .A4(new_n667_), .ZN(new_n674_));
  OAI22_X1   g0411(.A1(new_n274_), .A2(new_n665_), .B1(new_n674_), .B2(new_n285_), .ZN(new_n675_));
  INV_X1     g0412(.I(\a[101] ), .ZN(new_n676_));
  NOR3_X1    g0413(.A1(new_n676_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n677_));
  INV_X1     g0414(.I(\a[98] ), .ZN(new_n678_));
  NOR3_X1    g0415(.A1(new_n678_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n679_));
  INV_X1     g0416(.I(\a[100] ), .ZN(new_n680_));
  NOR3_X1    g0417(.A1(new_n680_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n681_));
  INV_X1     g0418(.I(\a[99] ), .ZN(new_n682_));
  NOR3_X1    g0419(.A1(new_n682_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n683_));
  NOR4_X1    g0420(.A1(new_n679_), .A2(new_n681_), .A3(new_n683_), .A4(new_n677_), .ZN(new_n684_));
  INV_X1     g0421(.I(\a[105] ), .ZN(new_n685_));
  NOR3_X1    g0422(.A1(new_n685_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n686_));
  INV_X1     g0423(.I(\a[102] ), .ZN(new_n687_));
  NOR3_X1    g0424(.A1(new_n687_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n688_));
  INV_X1     g0425(.I(\a[104] ), .ZN(new_n689_));
  NOR3_X1    g0426(.A1(new_n689_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n690_));
  INV_X1     g0427(.I(\a[103] ), .ZN(new_n691_));
  NOR3_X1    g0428(.A1(new_n691_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n692_));
  NOR4_X1    g0429(.A1(new_n688_), .A2(new_n690_), .A3(new_n692_), .A4(new_n686_), .ZN(new_n693_));
  OAI22_X1   g0430(.A1(new_n557_), .A2(new_n684_), .B1(new_n693_), .B2(new_n304_), .ZN(new_n694_));
  OAI21_X1   g0431(.A1(new_n675_), .A2(new_n694_), .B(new_n405_), .ZN(new_n695_));
  NAND2_X1   g0432(.A1(new_n656_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1   g0433(.A1(new_n617_), .A2(new_n696_), .B(new_n264_), .ZN(new_n697_));
  INV_X1     g0434(.I(\a[65] ), .ZN(new_n698_));
  NOR3_X1    g0435(.A1(new_n698_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n699_));
  INV_X1     g0436(.I(\a[62] ), .ZN(new_n700_));
  NOR3_X1    g0437(.A1(new_n700_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n701_));
  INV_X1     g0438(.I(\a[64] ), .ZN(new_n702_));
  NOR3_X1    g0439(.A1(new_n702_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n703_));
  INV_X1     g0440(.I(\a[63] ), .ZN(new_n704_));
  NOR3_X1    g0441(.A1(new_n704_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n705_));
  NOR4_X1    g0442(.A1(new_n701_), .A2(new_n703_), .A3(new_n705_), .A4(new_n699_), .ZN(new_n706_));
  INV_X1     g0443(.I(\a[61] ), .ZN(new_n707_));
  NOR3_X1    g0444(.A1(new_n707_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n708_));
  INV_X1     g0445(.I(\a[58] ), .ZN(new_n709_));
  NOR3_X1    g0446(.A1(new_n709_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n710_));
  INV_X1     g0447(.I(\a[60] ), .ZN(new_n711_));
  NOR3_X1    g0448(.A1(new_n711_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n712_));
  INV_X1     g0449(.I(\a[59] ), .ZN(new_n713_));
  NOR3_X1    g0450(.A1(new_n713_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n714_));
  NOR4_X1    g0451(.A1(new_n710_), .A2(new_n712_), .A3(new_n714_), .A4(new_n708_), .ZN(new_n715_));
  OAI22_X1   g0452(.A1(new_n274_), .A2(new_n706_), .B1(new_n715_), .B2(new_n285_), .ZN(new_n716_));
  INV_X1     g0453(.I(\a[53] ), .ZN(new_n717_));
  NOR3_X1    g0454(.A1(new_n717_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n718_));
  INV_X1     g0455(.I(\a[50] ), .ZN(new_n719_));
  NOR3_X1    g0456(.A1(new_n719_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n720_));
  INV_X1     g0457(.I(\a[52] ), .ZN(new_n721_));
  NOR3_X1    g0458(.A1(new_n721_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n722_));
  INV_X1     g0459(.I(\a[51] ), .ZN(new_n723_));
  NOR3_X1    g0460(.A1(new_n723_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n724_));
  NOR4_X1    g0461(.A1(new_n720_), .A2(new_n722_), .A3(new_n724_), .A4(new_n718_), .ZN(new_n725_));
  INV_X1     g0462(.I(\a[57] ), .ZN(new_n726_));
  NOR3_X1    g0463(.A1(new_n726_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n727_));
  INV_X1     g0464(.I(\a[54] ), .ZN(new_n728_));
  NOR3_X1    g0465(.A1(new_n728_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n729_));
  INV_X1     g0466(.I(\a[56] ), .ZN(new_n730_));
  NOR3_X1    g0467(.A1(new_n730_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n731_));
  INV_X1     g0468(.I(\a[55] ), .ZN(new_n732_));
  NOR3_X1    g0469(.A1(new_n732_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n733_));
  NOR4_X1    g0470(.A1(new_n729_), .A2(new_n731_), .A3(new_n733_), .A4(new_n727_), .ZN(new_n734_));
  OAI22_X1   g0471(.A1(new_n557_), .A2(new_n725_), .B1(new_n734_), .B2(new_n304_), .ZN(new_n735_));
  OAI21_X1   g0472(.A1(new_n716_), .A2(new_n735_), .B(new_n373_), .ZN(new_n736_));
  INV_X1     g0473(.I(\a[17] ), .ZN(new_n737_));
  NOR3_X1    g0474(.A1(new_n737_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n738_));
  INV_X1     g0475(.I(\a[14] ), .ZN(new_n739_));
  NOR3_X1    g0476(.A1(new_n739_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n740_));
  NAND2_X1   g0477(.A1(\a[16] ), .A2(\shift[0] ), .ZN(new_n741_));
  NOR2_X1    g0478(.A1(new_n741_), .A2(\shift[1] ), .ZN(new_n742_));
  INV_X1     g0479(.I(\a[15] ), .ZN(new_n743_));
  NOR3_X1    g0480(.A1(new_n743_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n744_));
  NOR4_X1    g0481(.A1(new_n740_), .A2(new_n742_), .A3(new_n744_), .A4(new_n738_), .ZN(new_n745_));
  INV_X1     g0482(.I(\a[13] ), .ZN(new_n746_));
  NOR3_X1    g0483(.A1(new_n746_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n747_));
  INV_X1     g0484(.I(\a[10] ), .ZN(new_n748_));
  NOR3_X1    g0485(.A1(new_n748_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n749_));
  NAND2_X1   g0486(.A1(\a[12] ), .A2(\shift[0] ), .ZN(new_n750_));
  NOR2_X1    g0487(.A1(new_n750_), .A2(\shift[1] ), .ZN(new_n751_));
  INV_X1     g0488(.I(\a[11] ), .ZN(new_n752_));
  NOR3_X1    g0489(.A1(new_n752_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n753_));
  NOR4_X1    g0490(.A1(new_n749_), .A2(new_n751_), .A3(new_n753_), .A4(new_n747_), .ZN(new_n754_));
  OAI22_X1   g0491(.A1(new_n274_), .A2(new_n745_), .B1(new_n754_), .B2(new_n285_), .ZN(new_n755_));
  INV_X1     g0492(.I(\a[5] ), .ZN(new_n756_));
  NOR3_X1    g0493(.A1(new_n756_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n757_));
  INV_X1     g0494(.I(\a[2] ), .ZN(new_n758_));
  NOR3_X1    g0495(.A1(new_n758_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n759_));
  NAND2_X1   g0496(.A1(\a[4] ), .A2(\shift[0] ), .ZN(new_n760_));
  NOR2_X1    g0497(.A1(new_n760_), .A2(\shift[1] ), .ZN(new_n761_));
  INV_X1     g0498(.I(\a[3] ), .ZN(new_n762_));
  NOR3_X1    g0499(.A1(new_n762_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n763_));
  NOR4_X1    g0500(.A1(new_n759_), .A2(new_n761_), .A3(new_n763_), .A4(new_n757_), .ZN(new_n764_));
  INV_X1     g0501(.I(\a[9] ), .ZN(new_n765_));
  NOR3_X1    g0502(.A1(new_n765_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n766_));
  INV_X1     g0503(.I(\a[6] ), .ZN(new_n767_));
  NOR3_X1    g0504(.A1(new_n767_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n768_));
  NAND2_X1   g0505(.A1(\a[8] ), .A2(\shift[0] ), .ZN(new_n769_));
  NOR2_X1    g0506(.A1(new_n769_), .A2(\shift[1] ), .ZN(new_n770_));
  INV_X1     g0507(.I(\a[7] ), .ZN(new_n771_));
  NOR3_X1    g0508(.A1(new_n771_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n772_));
  NOR4_X1    g0509(.A1(new_n768_), .A2(new_n770_), .A3(new_n772_), .A4(new_n766_), .ZN(new_n773_));
  OAI22_X1   g0510(.A1(new_n557_), .A2(new_n764_), .B1(new_n773_), .B2(new_n304_), .ZN(new_n774_));
  OAI21_X1   g0511(.A1(new_n755_), .A2(new_n774_), .B(new_n308_), .ZN(new_n775_));
  NAND2_X1   g0512(.A1(new_n736_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1     g0513(.I(\a[49] ), .ZN(new_n777_));
  NOR3_X1    g0514(.A1(new_n777_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n778_));
  NAND3_X1   g0515(.A1(\a[46] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n779_));
  INV_X1     g0516(.I(new_n779_), .ZN(new_n780_));
  NAND2_X1   g0517(.A1(\a[48] ), .A2(\shift[0] ), .ZN(new_n781_));
  NOR2_X1    g0518(.A1(new_n781_), .A2(\shift[1] ), .ZN(new_n782_));
  INV_X1     g0519(.I(\a[47] ), .ZN(new_n783_));
  NOR3_X1    g0520(.A1(new_n783_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n784_));
  NOR4_X1    g0521(.A1(new_n780_), .A2(new_n782_), .A3(new_n784_), .A4(new_n778_), .ZN(new_n785_));
  NAND3_X1   g0522(.A1(\a[42] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n786_));
  NAND3_X1   g0523(.A1(new_n266_), .A2(\a[43] ), .A3(\shift[1] ), .ZN(new_n787_));
  NAND2_X1   g0524(.A1(new_n787_), .A2(new_n786_), .ZN(new_n788_));
  NAND2_X1   g0525(.A1(new_n266_), .A2(\a[45] ), .ZN(new_n789_));
  NAND2_X1   g0526(.A1(\a[44] ), .A2(\shift[0] ), .ZN(new_n790_));
  AOI21_X1   g0527(.A1(new_n789_), .A2(new_n790_), .B(\shift[1] ), .ZN(new_n791_));
  NOR2_X1    g0528(.A1(new_n791_), .A2(new_n788_), .ZN(new_n792_));
  OAI22_X1   g0529(.A1(new_n792_), .A2(new_n285_), .B1(new_n785_), .B2(new_n274_), .ZN(new_n793_));
  NAND2_X1   g0530(.A1(new_n266_), .A2(\a[37] ), .ZN(new_n794_));
  NAND3_X1   g0531(.A1(\a[34] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n795_));
  OAI21_X1   g0532(.A1(new_n794_), .A2(\shift[1] ), .B(new_n795_), .ZN(new_n796_));
  NAND3_X1   g0533(.A1(new_n275_), .A2(\a[36] ), .A3(\shift[0] ), .ZN(new_n797_));
  NAND3_X1   g0534(.A1(new_n266_), .A2(\a[35] ), .A3(\shift[1] ), .ZN(new_n798_));
  NAND2_X1   g0535(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1   g0536(.A1(new_n799_), .A2(new_n796_), .B(new_n294_), .ZN(new_n800_));
  NAND2_X1   g0537(.A1(new_n266_), .A2(\a[41] ), .ZN(new_n801_));
  NAND2_X1   g0538(.A1(\a[40] ), .A2(\shift[0] ), .ZN(new_n802_));
  AOI21_X1   g0539(.A1(new_n801_), .A2(new_n802_), .B(\shift[1] ), .ZN(new_n803_));
  NAND3_X1   g0540(.A1(new_n266_), .A2(\a[39] ), .A3(\shift[1] ), .ZN(new_n804_));
  NAND3_X1   g0541(.A1(\a[38] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n805_));
  NAND2_X1   g0542(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1   g0543(.A1(new_n803_), .A2(new_n806_), .B(new_n303_), .ZN(new_n807_));
  NAND2_X1   g0544(.A1(new_n800_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1   g0545(.A1(new_n793_), .A2(new_n808_), .B(new_n405_), .ZN(new_n809_));
  INV_X1     g0546(.I(\a[33] ), .ZN(new_n810_));
  NOR3_X1    g0547(.A1(new_n810_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n811_));
  INV_X1     g0548(.I(\a[30] ), .ZN(new_n812_));
  NOR3_X1    g0549(.A1(new_n812_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n813_));
  INV_X1     g0550(.I(\a[32] ), .ZN(new_n814_));
  NOR3_X1    g0551(.A1(new_n814_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n815_));
  INV_X1     g0552(.I(\a[31] ), .ZN(new_n816_));
  NOR3_X1    g0553(.A1(new_n816_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n817_));
  NOR4_X1    g0554(.A1(new_n813_), .A2(new_n815_), .A3(new_n817_), .A4(new_n811_), .ZN(new_n818_));
  INV_X1     g0555(.I(\a[29] ), .ZN(new_n819_));
  NOR3_X1    g0556(.A1(new_n819_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n820_));
  INV_X1     g0557(.I(\a[26] ), .ZN(new_n821_));
  NOR3_X1    g0558(.A1(new_n821_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n822_));
  NAND2_X1   g0559(.A1(\a[28] ), .A2(\shift[0] ), .ZN(new_n823_));
  NOR2_X1    g0560(.A1(new_n823_), .A2(\shift[1] ), .ZN(new_n824_));
  INV_X1     g0561(.I(\a[27] ), .ZN(new_n825_));
  NOR3_X1    g0562(.A1(new_n825_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n826_));
  NOR4_X1    g0563(.A1(new_n822_), .A2(new_n824_), .A3(new_n826_), .A4(new_n820_), .ZN(new_n827_));
  OAI22_X1   g0564(.A1(new_n274_), .A2(new_n818_), .B1(new_n827_), .B2(new_n285_), .ZN(new_n828_));
  INV_X1     g0565(.I(\a[21] ), .ZN(new_n829_));
  NOR3_X1    g0566(.A1(new_n829_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n830_));
  INV_X1     g0567(.I(\a[18] ), .ZN(new_n831_));
  NOR3_X1    g0568(.A1(new_n831_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n832_));
  INV_X1     g0569(.I(\a[20] ), .ZN(new_n833_));
  NOR3_X1    g0570(.A1(new_n833_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n834_));
  INV_X1     g0571(.I(\a[19] ), .ZN(new_n835_));
  NOR3_X1    g0572(.A1(new_n835_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n836_));
  NOR4_X1    g0573(.A1(new_n832_), .A2(new_n834_), .A3(new_n836_), .A4(new_n830_), .ZN(new_n837_));
  INV_X1     g0574(.I(\a[25] ), .ZN(new_n838_));
  NOR3_X1    g0575(.A1(new_n838_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n839_));
  INV_X1     g0576(.I(\a[22] ), .ZN(new_n840_));
  NOR3_X1    g0577(.A1(new_n840_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n841_));
  NAND2_X1   g0578(.A1(\a[24] ), .A2(\shift[0] ), .ZN(new_n842_));
  NOR2_X1    g0579(.A1(new_n842_), .A2(\shift[1] ), .ZN(new_n843_));
  INV_X1     g0580(.I(\a[23] ), .ZN(new_n844_));
  NOR3_X1    g0581(.A1(new_n844_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n845_));
  NOR4_X1    g0582(.A1(new_n841_), .A2(new_n843_), .A3(new_n845_), .A4(new_n839_), .ZN(new_n846_));
  OAI22_X1   g0583(.A1(new_n557_), .A2(new_n837_), .B1(new_n846_), .B2(new_n304_), .ZN(new_n847_));
  OAI21_X1   g0584(.A1(new_n828_), .A2(new_n847_), .B(new_n340_), .ZN(new_n848_));
  NAND2_X1   g0585(.A1(new_n848_), .A2(new_n809_), .ZN(new_n849_));
  OAI21_X1   g0586(.A1(new_n776_), .A2(new_n849_), .B(\shift[6] ), .ZN(new_n850_));
  NAND2_X1   g0587(.A1(new_n697_), .A2(new_n850_), .ZN(\result[1] ));
  NAND2_X1   g0588(.A1(\a[81] ), .A2(\shift[0] ), .ZN(new_n852_));
  NAND2_X1   g0589(.A1(new_n266_), .A2(\a[82] ), .ZN(new_n853_));
  AOI21_X1   g0590(.A1(new_n853_), .A2(new_n852_), .B(\shift[1] ), .ZN(new_n854_));
  NAND3_X1   g0591(.A1(new_n266_), .A2(\a[80] ), .A3(\shift[1] ), .ZN(new_n855_));
  NAND3_X1   g0592(.A1(\a[79] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n856_));
  NAND2_X1   g0593(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1    g0594(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1   g0595(.A1(\a[77] ), .A2(\shift[0] ), .ZN(new_n859_));
  NAND2_X1   g0596(.A1(new_n266_), .A2(\a[78] ), .ZN(new_n860_));
  AOI21_X1   g0597(.A1(new_n860_), .A2(new_n859_), .B(\shift[1] ), .ZN(new_n861_));
  AOI21_X1   g0598(.A1(new_n279_), .A2(new_n280_), .B(new_n275_), .ZN(new_n862_));
  NOR2_X1    g0599(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI22_X1   g0600(.A1(new_n285_), .A2(new_n863_), .B1(new_n858_), .B2(new_n274_), .ZN(new_n864_));
  AOI21_X1   g0601(.A1(new_n297_), .A2(new_n296_), .B(\shift[1] ), .ZN(new_n865_));
  AOI21_X1   g0602(.A1(new_n290_), .A2(new_n291_), .B(new_n275_), .ZN(new_n866_));
  OAI21_X1   g0603(.A1(new_n865_), .A2(new_n866_), .B(new_n294_), .ZN(new_n867_));
  AOI21_X1   g0604(.A1(new_n277_), .A2(new_n276_), .B(\shift[1] ), .ZN(new_n868_));
  AOI21_X1   g0605(.A1(new_n299_), .A2(new_n300_), .B(new_n275_), .ZN(new_n869_));
  OAI21_X1   g0606(.A1(new_n868_), .A2(new_n869_), .B(new_n303_), .ZN(new_n870_));
  NAND2_X1   g0607(.A1(new_n867_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1   g0608(.A1(new_n864_), .A2(new_n871_), .B(new_n308_), .ZN(new_n872_));
  NAND2_X1   g0609(.A1(\a[97] ), .A2(\shift[0] ), .ZN(new_n873_));
  NAND2_X1   g0610(.A1(new_n266_), .A2(\a[98] ), .ZN(new_n874_));
  AOI21_X1   g0611(.A1(new_n874_), .A2(new_n873_), .B(\shift[1] ), .ZN(new_n875_));
  NAND3_X1   g0612(.A1(new_n266_), .A2(\a[96] ), .A3(\shift[1] ), .ZN(new_n876_));
  NAND3_X1   g0613(.A1(\a[95] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n877_));
  NAND2_X1   g0614(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI21_X1   g0615(.A1(new_n875_), .A2(new_n878_), .B(new_n273_), .ZN(new_n879_));
  NAND2_X1   g0616(.A1(\a[93] ), .A2(\shift[0] ), .ZN(new_n880_));
  NAND2_X1   g0617(.A1(new_n266_), .A2(\a[94] ), .ZN(new_n881_));
  AOI21_X1   g0618(.A1(new_n881_), .A2(new_n880_), .B(\shift[1] ), .ZN(new_n882_));
  AOI21_X1   g0619(.A1(new_n320_), .A2(new_n321_), .B(new_n275_), .ZN(new_n883_));
  OAI21_X1   g0620(.A1(new_n882_), .A2(new_n883_), .B(new_n284_), .ZN(new_n884_));
  NAND2_X1   g0621(.A1(new_n884_), .A2(new_n879_), .ZN(new_n885_));
  AOI21_X1   g0622(.A1(new_n333_), .A2(new_n332_), .B(\shift[1] ), .ZN(new_n886_));
  NAND3_X1   g0623(.A1(new_n266_), .A2(\a[84] ), .A3(\shift[1] ), .ZN(new_n887_));
  NAND3_X1   g0624(.A1(\a[83] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n888_));
  NAND2_X1   g0625(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1   g0626(.A1(new_n886_), .A2(new_n889_), .B(new_n294_), .ZN(new_n890_));
  AOI21_X1   g0627(.A1(new_n318_), .A2(new_n317_), .B(\shift[1] ), .ZN(new_n891_));
  NAND3_X1   g0628(.A1(new_n266_), .A2(\a[88] ), .A3(\shift[1] ), .ZN(new_n892_));
  NAND3_X1   g0629(.A1(\a[87] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n893_));
  NAND2_X1   g0630(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1   g0631(.A1(new_n891_), .A2(new_n894_), .B(new_n303_), .ZN(new_n895_));
  NAND2_X1   g0632(.A1(new_n890_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1   g0633(.A1(new_n885_), .A2(new_n896_), .B(new_n340_), .ZN(new_n897_));
  NAND2_X1   g0634(.A1(new_n872_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1   g0635(.A1(\a[1] ), .A2(\shift[0] ), .ZN(new_n899_));
  NAND2_X1   g0636(.A1(new_n266_), .A2(\a[2] ), .ZN(new_n900_));
  AOI21_X1   g0637(.A1(new_n900_), .A2(new_n899_), .B(\shift[1] ), .ZN(new_n901_));
  NAND3_X1   g0638(.A1(new_n266_), .A2(\a[0] ), .A3(\shift[1] ), .ZN(new_n902_));
  NAND3_X1   g0639(.A1(\a[127] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n903_));
  NAND2_X1   g0640(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI21_X1   g0641(.A1(new_n901_), .A2(new_n904_), .B(new_n273_), .ZN(new_n905_));
  AOI21_X1   g0642(.A1(new_n344_), .A2(new_n343_), .B(\shift[1] ), .ZN(new_n906_));
  NAND3_X1   g0643(.A1(new_n266_), .A2(\a[124] ), .A3(\shift[1] ), .ZN(new_n907_));
  NAND3_X1   g0644(.A1(\a[123] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n908_));
  NAND2_X1   g0645(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI21_X1   g0646(.A1(new_n906_), .A2(new_n909_), .B(new_n284_), .ZN(new_n910_));
  NAND2_X1   g0647(.A1(new_n905_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1   g0648(.A1(\a[117] ), .A2(\shift[0] ), .ZN(new_n912_));
  NAND2_X1   g0649(.A1(new_n266_), .A2(\a[118] ), .ZN(new_n913_));
  AOI21_X1   g0650(.A1(new_n913_), .A2(new_n912_), .B(\shift[1] ), .ZN(new_n914_));
  NAND3_X1   g0651(.A1(new_n266_), .A2(\a[116] ), .A3(\shift[1] ), .ZN(new_n915_));
  NAND3_X1   g0652(.A1(\a[115] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n916_));
  NAND2_X1   g0653(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1   g0654(.A1(new_n914_), .A2(new_n917_), .B(new_n294_), .ZN(new_n918_));
  NAND2_X1   g0655(.A1(\a[121] ), .A2(\shift[0] ), .ZN(new_n919_));
  NAND2_X1   g0656(.A1(new_n266_), .A2(\a[122] ), .ZN(new_n920_));
  AOI21_X1   g0657(.A1(new_n920_), .A2(new_n919_), .B(\shift[1] ), .ZN(new_n921_));
  NAND3_X1   g0658(.A1(new_n266_), .A2(\a[120] ), .A3(\shift[1] ), .ZN(new_n922_));
  NAND3_X1   g0659(.A1(\a[119] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n923_));
  NAND2_X1   g0660(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OAI21_X1   g0661(.A1(new_n921_), .A2(new_n924_), .B(new_n303_), .ZN(new_n925_));
  NAND2_X1   g0662(.A1(new_n918_), .A2(new_n925_), .ZN(new_n926_));
  OAI21_X1   g0663(.A1(new_n911_), .A2(new_n926_), .B(new_n373_), .ZN(new_n927_));
  NAND2_X1   g0664(.A1(\a[113] ), .A2(\shift[0] ), .ZN(new_n928_));
  NAND2_X1   g0665(.A1(new_n266_), .A2(\a[114] ), .ZN(new_n929_));
  AOI21_X1   g0666(.A1(new_n929_), .A2(new_n928_), .B(\shift[1] ), .ZN(new_n930_));
  NAND3_X1   g0667(.A1(new_n266_), .A2(\a[112] ), .A3(\shift[1] ), .ZN(new_n931_));
  NAND3_X1   g0668(.A1(\a[111] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n932_));
  NAND2_X1   g0669(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1   g0670(.A1(new_n930_), .A2(new_n933_), .B(new_n273_), .ZN(new_n934_));
  NAND2_X1   g0671(.A1(\a[109] ), .A2(\shift[0] ), .ZN(new_n935_));
  NAND2_X1   g0672(.A1(new_n266_), .A2(\a[110] ), .ZN(new_n936_));
  AOI21_X1   g0673(.A1(new_n936_), .A2(new_n935_), .B(\shift[1] ), .ZN(new_n937_));
  NAND3_X1   g0674(.A1(new_n266_), .A2(\a[108] ), .A3(\shift[1] ), .ZN(new_n938_));
  NAND3_X1   g0675(.A1(\a[107] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n939_));
  NAND2_X1   g0676(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  OAI21_X1   g0677(.A1(new_n937_), .A2(new_n940_), .B(new_n284_), .ZN(new_n941_));
  NAND2_X1   g0678(.A1(new_n934_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1   g0679(.A1(\a[101] ), .A2(\shift[0] ), .ZN(new_n943_));
  NAND2_X1   g0680(.A1(new_n266_), .A2(\a[102] ), .ZN(new_n944_));
  AOI21_X1   g0681(.A1(new_n944_), .A2(new_n943_), .B(\shift[1] ), .ZN(new_n945_));
  NAND3_X1   g0682(.A1(new_n266_), .A2(\a[100] ), .A3(\shift[1] ), .ZN(new_n946_));
  NAND3_X1   g0683(.A1(\a[99] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n947_));
  NAND2_X1   g0684(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  OAI21_X1   g0685(.A1(new_n945_), .A2(new_n948_), .B(new_n294_), .ZN(new_n949_));
  NAND2_X1   g0686(.A1(\a[105] ), .A2(\shift[0] ), .ZN(new_n950_));
  NAND2_X1   g0687(.A1(new_n266_), .A2(\a[106] ), .ZN(new_n951_));
  AOI21_X1   g0688(.A1(new_n951_), .A2(new_n950_), .B(\shift[1] ), .ZN(new_n952_));
  NAND3_X1   g0689(.A1(new_n266_), .A2(\a[104] ), .A3(\shift[1] ), .ZN(new_n953_));
  NAND3_X1   g0690(.A1(\a[103] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n954_));
  NAND2_X1   g0691(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  OAI21_X1   g0692(.A1(new_n952_), .A2(new_n955_), .B(new_n303_), .ZN(new_n956_));
  NAND2_X1   g0693(.A1(new_n949_), .A2(new_n956_), .ZN(new_n957_));
  OAI21_X1   g0694(.A1(new_n942_), .A2(new_n957_), .B(new_n405_), .ZN(new_n958_));
  NAND2_X1   g0695(.A1(new_n927_), .A2(new_n958_), .ZN(new_n959_));
  OAI21_X1   g0696(.A1(new_n898_), .A2(new_n959_), .B(new_n264_), .ZN(new_n960_));
  AOI21_X1   g0697(.A1(new_n288_), .A2(new_n287_), .B(\shift[1] ), .ZN(new_n961_));
  AOI21_X1   g0698(.A1(new_n475_), .A2(new_n476_), .B(new_n275_), .ZN(new_n962_));
  NOR2_X1    g0699(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  AOI21_X1   g0700(.A1(new_n473_), .A2(new_n472_), .B(\shift[1] ), .ZN(new_n964_));
  NAND3_X1   g0701(.A1(new_n266_), .A2(\a[60] ), .A3(\shift[1] ), .ZN(new_n965_));
  NAND3_X1   g0702(.A1(\a[59] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n966_));
  NAND2_X1   g0703(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  NOR2_X1    g0704(.A1(new_n964_), .A2(new_n967_), .ZN(new_n968_));
  OAI22_X1   g0705(.A1(new_n274_), .A2(new_n963_), .B1(new_n968_), .B2(new_n285_), .ZN(new_n969_));
  AOI21_X1   g0706(.A1(new_n495_), .A2(new_n494_), .B(\shift[1] ), .ZN(new_n970_));
  AOI21_X1   g0707(.A1(new_n490_), .A2(new_n491_), .B(new_n275_), .ZN(new_n971_));
  OAI21_X1   g0708(.A1(new_n970_), .A2(new_n971_), .B(new_n294_), .ZN(new_n972_));
  NAND2_X1   g0709(.A1(\a[57] ), .A2(\shift[0] ), .ZN(new_n973_));
  NAND2_X1   g0710(.A1(new_n266_), .A2(\a[58] ), .ZN(new_n974_));
  AOI21_X1   g0711(.A1(new_n974_), .A2(new_n973_), .B(\shift[1] ), .ZN(new_n975_));
  AOI21_X1   g0712(.A1(new_n497_), .A2(new_n498_), .B(new_n275_), .ZN(new_n976_));
  NOR2_X1    g0713(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  OAI21_X1   g0714(.A1(new_n304_), .A2(new_n977_), .B(new_n972_), .ZN(new_n978_));
  OAI21_X1   g0715(.A1(new_n969_), .A2(new_n978_), .B(new_n373_), .ZN(new_n979_));
  NAND2_X1   g0716(.A1(\a[17] ), .A2(\shift[0] ), .ZN(new_n980_));
  NAND2_X1   g0717(.A1(new_n266_), .A2(\a[18] ), .ZN(new_n981_));
  AOI21_X1   g0718(.A1(new_n981_), .A2(new_n980_), .B(\shift[1] ), .ZN(new_n982_));
  NAND3_X1   g0719(.A1(new_n266_), .A2(\a[16] ), .A3(\shift[1] ), .ZN(new_n983_));
  NAND3_X1   g0720(.A1(\a[15] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n984_));
  NAND2_X1   g0721(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  OAI21_X1   g0722(.A1(new_n982_), .A2(new_n985_), .B(new_n273_), .ZN(new_n986_));
  NAND2_X1   g0723(.A1(\a[13] ), .A2(\shift[0] ), .ZN(new_n987_));
  NAND2_X1   g0724(.A1(new_n266_), .A2(\a[14] ), .ZN(new_n988_));
  AOI21_X1   g0725(.A1(new_n988_), .A2(new_n987_), .B(\shift[1] ), .ZN(new_n989_));
  NAND3_X1   g0726(.A1(new_n266_), .A2(\a[12] ), .A3(\shift[1] ), .ZN(new_n990_));
  NAND3_X1   g0727(.A1(\a[11] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n991_));
  NAND2_X1   g0728(.A1(new_n990_), .A2(new_n991_), .ZN(new_n992_));
  OAI21_X1   g0729(.A1(new_n989_), .A2(new_n992_), .B(new_n284_), .ZN(new_n993_));
  NAND2_X1   g0730(.A1(new_n986_), .A2(new_n993_), .ZN(new_n994_));
  NAND2_X1   g0731(.A1(\a[5] ), .A2(\shift[0] ), .ZN(new_n995_));
  NAND2_X1   g0732(.A1(new_n266_), .A2(\a[6] ), .ZN(new_n996_));
  AOI21_X1   g0733(.A1(new_n996_), .A2(new_n995_), .B(\shift[1] ), .ZN(new_n997_));
  NAND3_X1   g0734(.A1(new_n266_), .A2(\a[4] ), .A3(\shift[1] ), .ZN(new_n998_));
  NAND3_X1   g0735(.A1(\a[3] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n999_));
  NAND2_X1   g0736(.A1(new_n998_), .A2(new_n999_), .ZN(new_n1000_));
  OAI21_X1   g0737(.A1(new_n997_), .A2(new_n1000_), .B(new_n294_), .ZN(new_n1001_));
  NAND2_X1   g0738(.A1(\a[9] ), .A2(\shift[0] ), .ZN(new_n1002_));
  NAND2_X1   g0739(.A1(new_n266_), .A2(\a[10] ), .ZN(new_n1003_));
  AOI21_X1   g0740(.A1(new_n1003_), .A2(new_n1002_), .B(\shift[1] ), .ZN(new_n1004_));
  NAND3_X1   g0741(.A1(new_n266_), .A2(\a[8] ), .A3(\shift[1] ), .ZN(new_n1005_));
  NAND3_X1   g0742(.A1(\a[7] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1006_));
  NAND2_X1   g0743(.A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1007_));
  OAI21_X1   g0744(.A1(new_n1004_), .A2(new_n1007_), .B(new_n303_), .ZN(new_n1008_));
  NAND2_X1   g0745(.A1(new_n1001_), .A2(new_n1008_), .ZN(new_n1009_));
  OAI21_X1   g0746(.A1(new_n994_), .A2(new_n1009_), .B(new_n308_), .ZN(new_n1010_));
  NAND2_X1   g0747(.A1(new_n979_), .A2(new_n1010_), .ZN(new_n1011_));
  AOI21_X1   g0748(.A1(new_n488_), .A2(new_n487_), .B(\shift[1] ), .ZN(new_n1012_));
  AOI21_X1   g0749(.A1(new_n506_), .A2(new_n507_), .B(new_n275_), .ZN(new_n1013_));
  NOR2_X1    g0750(.A1(new_n1012_), .A2(new_n1013_), .ZN(new_n1014_));
  NAND3_X1   g0751(.A1(\a[43] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1015_));
  NAND3_X1   g0752(.A1(new_n266_), .A2(\a[44] ), .A3(\shift[1] ), .ZN(new_n1016_));
  NAND2_X1   g0753(.A1(new_n1016_), .A2(new_n1015_), .ZN(new_n1017_));
  AOI21_X1   g0754(.A1(new_n504_), .A2(new_n503_), .B(\shift[1] ), .ZN(new_n1018_));
  NOR2_X1    g0755(.A1(new_n1018_), .A2(new_n1017_), .ZN(new_n1019_));
  OAI22_X1   g0756(.A1(new_n274_), .A2(new_n1014_), .B1(new_n1019_), .B2(new_n285_), .ZN(new_n1020_));
  NAND2_X1   g0757(.A1(\a[37] ), .A2(\shift[0] ), .ZN(new_n1021_));
  NAND2_X1   g0758(.A1(new_n266_), .A2(\a[38] ), .ZN(new_n1022_));
  AOI21_X1   g0759(.A1(new_n1022_), .A2(new_n1021_), .B(\shift[1] ), .ZN(new_n1023_));
  AOI21_X1   g0760(.A1(new_n521_), .A2(new_n522_), .B(new_n275_), .ZN(new_n1024_));
  OAI21_X1   g0761(.A1(new_n1023_), .A2(new_n1024_), .B(new_n294_), .ZN(new_n1025_));
  NAND2_X1   g0762(.A1(\a[41] ), .A2(\shift[0] ), .ZN(new_n1026_));
  NAND2_X1   g0763(.A1(new_n266_), .A2(\a[42] ), .ZN(new_n1027_));
  AOI21_X1   g0764(.A1(new_n1027_), .A2(new_n1026_), .B(\shift[1] ), .ZN(new_n1028_));
  NAND2_X1   g0765(.A1(\a[39] ), .A2(\shift[0] ), .ZN(new_n1029_));
  AOI21_X1   g0766(.A1(new_n525_), .A2(new_n1029_), .B(new_n275_), .ZN(new_n1030_));
  OAI21_X1   g0767(.A1(new_n1028_), .A2(new_n1030_), .B(new_n303_), .ZN(new_n1031_));
  NAND2_X1   g0768(.A1(new_n1025_), .A2(new_n1031_), .ZN(new_n1032_));
  OAI21_X1   g0769(.A1(new_n1020_), .A2(new_n1032_), .B(new_n405_), .ZN(new_n1033_));
  NAND2_X1   g0770(.A1(\a[33] ), .A2(\shift[0] ), .ZN(new_n1034_));
  NAND2_X1   g0771(.A1(new_n266_), .A2(\a[34] ), .ZN(new_n1035_));
  AOI21_X1   g0772(.A1(new_n1035_), .A2(new_n1034_), .B(\shift[1] ), .ZN(new_n1036_));
  AOI21_X1   g0773(.A1(new_n443_), .A2(new_n444_), .B(new_n275_), .ZN(new_n1037_));
  OAI21_X1   g0774(.A1(new_n1036_), .A2(new_n1037_), .B(new_n273_), .ZN(new_n1038_));
  NAND2_X1   g0775(.A1(\a[29] ), .A2(\shift[0] ), .ZN(new_n1039_));
  NAND2_X1   g0776(.A1(new_n266_), .A2(\a[30] ), .ZN(new_n1040_));
  AOI21_X1   g0777(.A1(new_n1040_), .A2(new_n1039_), .B(\shift[1] ), .ZN(new_n1041_));
  AOI21_X1   g0778(.A1(new_n450_), .A2(new_n451_), .B(new_n275_), .ZN(new_n1042_));
  OAI21_X1   g0779(.A1(new_n1041_), .A2(new_n1042_), .B(new_n284_), .ZN(new_n1043_));
  NAND2_X1   g0780(.A1(new_n1038_), .A2(new_n1043_), .ZN(new_n1044_));
  NAND2_X1   g0781(.A1(\a[21] ), .A2(\shift[0] ), .ZN(new_n1045_));
  NAND2_X1   g0782(.A1(new_n266_), .A2(\a[22] ), .ZN(new_n1046_));
  AOI21_X1   g0783(.A1(new_n1046_), .A2(new_n1045_), .B(\shift[1] ), .ZN(new_n1047_));
  NAND3_X1   g0784(.A1(new_n266_), .A2(\a[20] ), .A3(\shift[1] ), .ZN(new_n1048_));
  NAND3_X1   g0785(.A1(\a[19] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1049_));
  NAND2_X1   g0786(.A1(new_n1048_), .A2(new_n1049_), .ZN(new_n1050_));
  OAI21_X1   g0787(.A1(new_n1047_), .A2(new_n1050_), .B(new_n294_), .ZN(new_n1051_));
  AOI21_X1   g0788(.A1(new_n448_), .A2(new_n447_), .B(\shift[1] ), .ZN(new_n1052_));
  NAND3_X1   g0789(.A1(new_n266_), .A2(\a[24] ), .A3(\shift[1] ), .ZN(new_n1053_));
  NAND3_X1   g0790(.A1(\a[23] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1054_));
  NAND2_X1   g0791(.A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_));
  OAI21_X1   g0792(.A1(new_n1052_), .A2(new_n1055_), .B(new_n303_), .ZN(new_n1056_));
  NAND2_X1   g0793(.A1(new_n1051_), .A2(new_n1056_), .ZN(new_n1057_));
  OAI21_X1   g0794(.A1(new_n1044_), .A2(new_n1057_), .B(new_n340_), .ZN(new_n1058_));
  NAND2_X1   g0795(.A1(new_n1033_), .A2(new_n1058_), .ZN(new_n1059_));
  OAI21_X1   g0796(.A1(new_n1011_), .A2(new_n1059_), .B(\shift[6] ), .ZN(new_n1060_));
  NAND2_X1   g0797(.A1(new_n960_), .A2(new_n1060_), .ZN(\result[2] ));
  INV_X1     g0798(.I(new_n340_), .ZN(new_n1062_));
  NOR3_X1    g0799(.A1(new_n657_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1063_));
  NOR3_X1    g0800(.A1(new_n639_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1064_));
  NOR3_X1    g0801(.A1(new_n661_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1065_));
  NOR3_X1    g0802(.A1(new_n643_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1066_));
  NOR4_X1    g0803(.A1(new_n1065_), .A2(new_n1063_), .A3(new_n1064_), .A4(new_n1066_), .ZN(new_n1067_));
  NOR3_X1    g0804(.A1(new_n666_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1068_));
  NOR3_X1    g0805(.A1(new_n659_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1069_));
  NOR3_X1    g0806(.A1(new_n670_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1070_));
  NOR3_X1    g0807(.A1(new_n663_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1071_));
  NOR4_X1    g0808(.A1(new_n1070_), .A2(new_n1068_), .A3(new_n1069_), .A4(new_n1071_), .ZN(new_n1072_));
  OAI22_X1   g0809(.A1(new_n274_), .A2(new_n1067_), .B1(new_n1072_), .B2(new_n285_), .ZN(new_n1073_));
  NOR3_X1    g0810(.A1(new_n676_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1074_));
  NOR3_X1    g0811(.A1(new_n687_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1075_));
  NOR3_X1    g0812(.A1(new_n680_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1076_));
  NOR3_X1    g0813(.A1(new_n691_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1077_));
  NOR4_X1    g0814(.A1(new_n1076_), .A2(new_n1074_), .A3(new_n1075_), .A4(new_n1077_), .ZN(new_n1078_));
  NOR3_X1    g0815(.A1(new_n685_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1079_));
  NOR3_X1    g0816(.A1(new_n668_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1080_));
  NOR3_X1    g0817(.A1(new_n689_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1081_));
  NOR3_X1    g0818(.A1(new_n672_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1082_));
  NOR4_X1    g0819(.A1(new_n1081_), .A2(new_n1079_), .A3(new_n1080_), .A4(new_n1082_), .ZN(new_n1083_));
  OAI22_X1   g0820(.A1(new_n557_), .A2(new_n1078_), .B1(new_n1083_), .B2(new_n304_), .ZN(new_n1084_));
  OAI21_X1   g0821(.A1(new_n1073_), .A2(new_n1084_), .B(new_n405_), .ZN(new_n1085_));
  NOR3_X1    g0822(.A1(new_n578_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1086_));
  NOR3_X1    g0823(.A1(new_n678_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1087_));
  NOR3_X1    g0824(.A1(new_n582_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1088_));
  NOR3_X1    g0825(.A1(new_n682_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1089_));
  NOR4_X1    g0826(.A1(new_n1088_), .A2(new_n1086_), .A3(new_n1087_), .A4(new_n1089_), .ZN(new_n1090_));
  NOR3_X1    g0827(.A1(new_n587_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1091_));
  NOR3_X1    g0828(.A1(new_n580_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1092_));
  NOR3_X1    g0829(.A1(new_n591_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1093_));
  NOR3_X1    g0830(.A1(new_n584_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1094_));
  NOR4_X1    g0831(.A1(new_n1093_), .A2(new_n1091_), .A3(new_n1092_), .A4(new_n1094_), .ZN(new_n1095_));
  OAI22_X1   g0832(.A1(new_n274_), .A2(new_n1090_), .B1(new_n1095_), .B2(new_n285_), .ZN(new_n1096_));
  NOR3_X1    g0833(.A1(new_n597_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1097_));
  NOR3_X1    g0834(.A1(new_n608_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1098_));
  NOR3_X1    g0835(.A1(new_n601_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1099_));
  NOR3_X1    g0836(.A1(new_n612_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1100_));
  NOR4_X1    g0837(.A1(new_n1099_), .A2(new_n1097_), .A3(new_n1098_), .A4(new_n1100_), .ZN(new_n1101_));
  NOR3_X1    g0838(.A1(new_n606_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1102_));
  NOR3_X1    g0839(.A1(new_n589_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1103_));
  NOR2_X1    g0840(.A1(new_n610_), .A2(new_n275_), .ZN(new_n1104_));
  NOR3_X1    g0841(.A1(new_n593_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1105_));
  NOR4_X1    g0842(.A1(new_n1102_), .A2(new_n1104_), .A3(new_n1103_), .A4(new_n1105_), .ZN(new_n1106_));
  OAI22_X1   g0843(.A1(new_n557_), .A2(new_n1101_), .B1(new_n1106_), .B2(new_n304_), .ZN(new_n1107_));
  NOR2_X1    g0844(.A1(new_n1096_), .A2(new_n1107_), .ZN(new_n1108_));
  OAI21_X1   g0845(.A1(new_n1062_), .A2(new_n1108_), .B(new_n1085_), .ZN(new_n1109_));
  NOR3_X1    g0846(.A1(new_n618_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1110_));
  NOR3_X1    g0847(.A1(new_n758_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1111_));
  NOR3_X1    g0848(.A1(new_n622_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1112_));
  NOR3_X1    g0849(.A1(new_n762_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1113_));
  NOR4_X1    g0850(.A1(new_n1112_), .A2(new_n1110_), .A3(new_n1111_), .A4(new_n1113_), .ZN(new_n1114_));
  NOR3_X1    g0851(.A1(new_n627_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1115_));
  NOR3_X1    g0852(.A1(new_n620_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1116_));
  NOR3_X1    g0853(.A1(new_n631_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1117_));
  NOR3_X1    g0854(.A1(new_n624_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1118_));
  NOR4_X1    g0855(.A1(new_n1117_), .A2(new_n1115_), .A3(new_n1116_), .A4(new_n1118_), .ZN(new_n1119_));
  OAI22_X1   g0856(.A1(new_n274_), .A2(new_n1114_), .B1(new_n1119_), .B2(new_n285_), .ZN(new_n1120_));
  NOR3_X1    g0857(.A1(new_n637_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1121_));
  NOR3_X1    g0858(.A1(new_n648_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1122_));
  NOR3_X1    g0859(.A1(new_n641_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1123_));
  NOR3_X1    g0860(.A1(new_n652_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1124_));
  NOR4_X1    g0861(.A1(new_n1123_), .A2(new_n1121_), .A3(new_n1122_), .A4(new_n1124_), .ZN(new_n1125_));
  NOR3_X1    g0862(.A1(new_n646_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1126_));
  NOR3_X1    g0863(.A1(new_n629_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1127_));
  NOR3_X1    g0864(.A1(new_n650_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1128_));
  NOR3_X1    g0865(.A1(new_n633_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1129_));
  NOR4_X1    g0866(.A1(new_n1128_), .A2(new_n1126_), .A3(new_n1127_), .A4(new_n1129_), .ZN(new_n1130_));
  OAI22_X1   g0867(.A1(new_n557_), .A2(new_n1125_), .B1(new_n1130_), .B2(new_n304_), .ZN(new_n1131_));
  OAI21_X1   g0868(.A1(new_n1120_), .A2(new_n1131_), .B(new_n373_), .ZN(new_n1132_));
  NOR3_X1    g0869(.A1(new_n538_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1133_));
  NOR3_X1    g0870(.A1(new_n599_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1134_));
  NOR2_X1    g0871(.A1(new_n542_), .A2(new_n275_), .ZN(new_n1135_));
  NOR3_X1    g0872(.A1(new_n603_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1136_));
  NOR4_X1    g0873(.A1(new_n1133_), .A2(new_n1135_), .A3(new_n1134_), .A4(new_n1136_), .ZN(new_n1137_));
  NOR3_X1    g0874(.A1(new_n547_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1138_));
  NOR3_X1    g0875(.A1(new_n540_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1139_));
  NOR2_X1    g0876(.A1(new_n551_), .A2(new_n275_), .ZN(new_n1140_));
  NOR3_X1    g0877(.A1(new_n544_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1141_));
  NOR4_X1    g0878(.A1(new_n1138_), .A2(new_n1140_), .A3(new_n1139_), .A4(new_n1141_), .ZN(new_n1142_));
  OAI22_X1   g0879(.A1(new_n274_), .A2(new_n1137_), .B1(new_n1142_), .B2(new_n285_), .ZN(new_n1143_));
  NOR3_X1    g0880(.A1(new_n558_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1144_));
  NOR3_X1    g0881(.A1(new_n569_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1145_));
  NOR2_X1    g0882(.A1(new_n562_), .A2(new_n275_), .ZN(new_n1146_));
  NOR3_X1    g0883(.A1(new_n573_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1147_));
  NOR4_X1    g0884(.A1(new_n1144_), .A2(new_n1146_), .A3(new_n1145_), .A4(new_n1147_), .ZN(new_n1148_));
  NOR3_X1    g0885(.A1(new_n567_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1149_));
  NOR3_X1    g0886(.A1(new_n549_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1150_));
  NOR2_X1    g0887(.A1(new_n571_), .A2(new_n275_), .ZN(new_n1151_));
  NOR3_X1    g0888(.A1(new_n553_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1152_));
  NOR4_X1    g0889(.A1(new_n1149_), .A2(new_n1151_), .A3(new_n1150_), .A4(new_n1152_), .ZN(new_n1153_));
  OAI22_X1   g0890(.A1(new_n557_), .A2(new_n1148_), .B1(new_n1153_), .B2(new_n304_), .ZN(new_n1154_));
  OAI21_X1   g0891(.A1(new_n1143_), .A2(new_n1154_), .B(new_n308_), .ZN(new_n1155_));
  NAND2_X1   g0892(.A1(new_n1132_), .A2(new_n1155_), .ZN(new_n1156_));
  OAI21_X1   g0893(.A1(new_n1109_), .A2(new_n1156_), .B(new_n264_), .ZN(new_n1157_));
  NOR3_X1    g0894(.A1(new_n698_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1158_));
  NOR3_X1    g0895(.A1(new_n560_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1159_));
  NOR3_X1    g0896(.A1(new_n702_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1160_));
  NOR3_X1    g0897(.A1(new_n564_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1161_));
  NOR4_X1    g0898(.A1(new_n1160_), .A2(new_n1158_), .A3(new_n1159_), .A4(new_n1161_), .ZN(new_n1162_));
  NOR3_X1    g0899(.A1(new_n707_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1163_));
  NOR3_X1    g0900(.A1(new_n700_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1164_));
  NOR3_X1    g0901(.A1(new_n711_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1165_));
  NOR3_X1    g0902(.A1(new_n704_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1166_));
  NOR4_X1    g0903(.A1(new_n1165_), .A2(new_n1163_), .A3(new_n1164_), .A4(new_n1166_), .ZN(new_n1167_));
  OAI22_X1   g0904(.A1(new_n274_), .A2(new_n1162_), .B1(new_n1167_), .B2(new_n285_), .ZN(new_n1168_));
  NOR3_X1    g0905(.A1(new_n717_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1169_));
  NOR3_X1    g0906(.A1(new_n728_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1170_));
  NAND3_X1   g0907(.A1(\a[52] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1171_));
  INV_X1     g0908(.I(new_n1171_), .ZN(new_n1172_));
  NOR3_X1    g0909(.A1(new_n732_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1173_));
  NOR4_X1    g0910(.A1(new_n1172_), .A2(new_n1169_), .A3(new_n1170_), .A4(new_n1173_), .ZN(new_n1174_));
  NOR3_X1    g0911(.A1(new_n726_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1175_));
  NOR3_X1    g0912(.A1(new_n709_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1176_));
  NOR3_X1    g0913(.A1(new_n730_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1177_));
  NOR3_X1    g0914(.A1(new_n713_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1178_));
  NOR4_X1    g0915(.A1(new_n1177_), .A2(new_n1175_), .A3(new_n1176_), .A4(new_n1178_), .ZN(new_n1179_));
  OAI22_X1   g0916(.A1(new_n557_), .A2(new_n1174_), .B1(new_n1179_), .B2(new_n304_), .ZN(new_n1180_));
  OAI21_X1   g0917(.A1(new_n1168_), .A2(new_n1180_), .B(new_n373_), .ZN(new_n1181_));
  NAND3_X1   g0918(.A1(new_n266_), .A2(\a[49] ), .A3(\shift[1] ), .ZN(new_n1182_));
  NAND3_X1   g0919(.A1(new_n275_), .A2(\a[50] ), .A3(\shift[0] ), .ZN(new_n1183_));
  NAND2_X1   g0920(.A1(new_n1182_), .A2(new_n1183_), .ZN(new_n1184_));
  NAND2_X1   g0921(.A1(new_n266_), .A2(\a[51] ), .ZN(new_n1185_));
  NAND3_X1   g0922(.A1(\a[48] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1186_));
  OAI21_X1   g0923(.A1(new_n1185_), .A2(\shift[1] ), .B(new_n1186_), .ZN(new_n1187_));
  OAI21_X1   g0924(.A1(new_n1184_), .A2(new_n1187_), .B(new_n273_), .ZN(new_n1188_));
  NAND3_X1   g0925(.A1(\a[44] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1189_));
  NAND3_X1   g0926(.A1(new_n266_), .A2(\a[45] ), .A3(\shift[1] ), .ZN(new_n1190_));
  NAND2_X1   g0927(.A1(new_n1190_), .A2(new_n1189_), .ZN(new_n1191_));
  NAND2_X1   g0928(.A1(\a[46] ), .A2(\shift[0] ), .ZN(new_n1192_));
  NAND2_X1   g0929(.A1(new_n266_), .A2(\a[47] ), .ZN(new_n1193_));
  AOI21_X1   g0930(.A1(new_n1193_), .A2(new_n1192_), .B(\shift[1] ), .ZN(new_n1194_));
  OAI21_X1   g0931(.A1(new_n1194_), .A2(new_n1191_), .B(new_n284_), .ZN(new_n1195_));
  NAND2_X1   g0932(.A1(new_n1188_), .A2(new_n1195_), .ZN(new_n1196_));
  INV_X1     g0933(.I(\a[37] ), .ZN(new_n1197_));
  NOR3_X1    g0934(.A1(new_n1197_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1198_));
  NAND2_X1   g0935(.A1(\a[38] ), .A2(\shift[0] ), .ZN(new_n1199_));
  NOR2_X1    g0936(.A1(new_n1199_), .A2(\shift[1] ), .ZN(new_n1200_));
  NAND2_X1   g0937(.A1(\a[36] ), .A2(\shift[0] ), .ZN(new_n1201_));
  NOR2_X1    g0938(.A1(new_n1201_), .A2(new_n275_), .ZN(new_n1202_));
  INV_X1     g0939(.I(\a[39] ), .ZN(new_n1203_));
  NOR3_X1    g0940(.A1(new_n1203_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1204_));
  NOR4_X1    g0941(.A1(new_n1200_), .A2(new_n1202_), .A3(new_n1198_), .A4(new_n1204_), .ZN(new_n1205_));
  INV_X1     g0942(.I(\a[41] ), .ZN(new_n1206_));
  NOR3_X1    g0943(.A1(new_n1206_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1207_));
  NAND2_X1   g0944(.A1(\a[42] ), .A2(\shift[0] ), .ZN(new_n1208_));
  NOR2_X1    g0945(.A1(new_n1208_), .A2(\shift[1] ), .ZN(new_n1209_));
  NAND3_X1   g0946(.A1(\a[40] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1210_));
  INV_X1     g0947(.I(new_n1210_), .ZN(new_n1211_));
  INV_X1     g0948(.I(\a[43] ), .ZN(new_n1212_));
  NOR3_X1    g0949(.A1(new_n1212_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1213_));
  NOR4_X1    g0950(.A1(new_n1209_), .A2(new_n1211_), .A3(new_n1207_), .A4(new_n1213_), .ZN(new_n1214_));
  OAI22_X1   g0951(.A1(new_n557_), .A2(new_n1205_), .B1(new_n1214_), .B2(new_n304_), .ZN(new_n1215_));
  OAI21_X1   g0952(.A1(new_n1215_), .A2(new_n1196_), .B(new_n405_), .ZN(new_n1216_));
  NAND2_X1   g0953(.A1(new_n1181_), .A2(new_n1216_), .ZN(new_n1217_));
  NOR3_X1    g0954(.A1(new_n737_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1218_));
  NOR3_X1    g0955(.A1(new_n831_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1219_));
  NOR2_X1    g0956(.A1(new_n741_), .A2(new_n275_), .ZN(new_n1220_));
  NOR3_X1    g0957(.A1(new_n835_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1221_));
  NOR4_X1    g0958(.A1(new_n1218_), .A2(new_n1220_), .A3(new_n1219_), .A4(new_n1221_), .ZN(new_n1222_));
  NOR3_X1    g0959(.A1(new_n746_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1223_));
  NOR3_X1    g0960(.A1(new_n739_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1224_));
  NOR2_X1    g0961(.A1(new_n750_), .A2(new_n275_), .ZN(new_n1225_));
  NOR3_X1    g0962(.A1(new_n743_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1226_));
  NOR4_X1    g0963(.A1(new_n1223_), .A2(new_n1225_), .A3(new_n1224_), .A4(new_n1226_), .ZN(new_n1227_));
  OAI22_X1   g0964(.A1(new_n274_), .A2(new_n1222_), .B1(new_n1227_), .B2(new_n285_), .ZN(new_n1228_));
  NOR3_X1    g0965(.A1(new_n756_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1229_));
  NOR3_X1    g0966(.A1(new_n767_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1230_));
  NOR2_X1    g0967(.A1(new_n760_), .A2(new_n275_), .ZN(new_n1231_));
  NOR3_X1    g0968(.A1(new_n771_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1232_));
  NOR4_X1    g0969(.A1(new_n1229_), .A2(new_n1231_), .A3(new_n1230_), .A4(new_n1232_), .ZN(new_n1233_));
  NOR3_X1    g0970(.A1(new_n765_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1234_));
  NOR3_X1    g0971(.A1(new_n748_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1235_));
  NOR2_X1    g0972(.A1(new_n769_), .A2(new_n275_), .ZN(new_n1236_));
  NOR3_X1    g0973(.A1(new_n752_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1237_));
  NOR4_X1    g0974(.A1(new_n1234_), .A2(new_n1236_), .A3(new_n1235_), .A4(new_n1237_), .ZN(new_n1238_));
  OAI22_X1   g0975(.A1(new_n557_), .A2(new_n1233_), .B1(new_n1238_), .B2(new_n304_), .ZN(new_n1239_));
  OAI21_X1   g0976(.A1(new_n1228_), .A2(new_n1239_), .B(new_n308_), .ZN(new_n1240_));
  NOR3_X1    g0977(.A1(new_n810_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1241_));
  NAND2_X1   g0978(.A1(\a[34] ), .A2(\shift[0] ), .ZN(new_n1242_));
  NOR2_X1    g0979(.A1(new_n1242_), .A2(\shift[1] ), .ZN(new_n1243_));
  NOR3_X1    g0980(.A1(new_n814_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1244_));
  INV_X1     g0981(.I(\a[35] ), .ZN(new_n1245_));
  NOR3_X1    g0982(.A1(new_n1245_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1246_));
  NOR4_X1    g0983(.A1(new_n1244_), .A2(new_n1243_), .A3(new_n1241_), .A4(new_n1246_), .ZN(new_n1247_));
  NOR3_X1    g0984(.A1(new_n819_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1248_));
  NOR3_X1    g0985(.A1(new_n812_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1249_));
  NOR2_X1    g0986(.A1(new_n823_), .A2(new_n275_), .ZN(new_n1250_));
  NOR3_X1    g0987(.A1(new_n816_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1251_));
  NOR4_X1    g0988(.A1(new_n1248_), .A2(new_n1250_), .A3(new_n1249_), .A4(new_n1251_), .ZN(new_n1252_));
  OAI22_X1   g0989(.A1(new_n274_), .A2(new_n1247_), .B1(new_n1252_), .B2(new_n285_), .ZN(new_n1253_));
  NOR3_X1    g0990(.A1(new_n829_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1254_));
  NOR3_X1    g0991(.A1(new_n840_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1255_));
  NOR3_X1    g0992(.A1(new_n833_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n1256_));
  NOR3_X1    g0993(.A1(new_n844_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1257_));
  NOR4_X1    g0994(.A1(new_n1256_), .A2(new_n1254_), .A3(new_n1255_), .A4(new_n1257_), .ZN(new_n1258_));
  NOR3_X1    g0995(.A1(new_n838_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1259_));
  NOR3_X1    g0996(.A1(new_n821_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1260_));
  NOR2_X1    g0997(.A1(new_n842_), .A2(new_n275_), .ZN(new_n1261_));
  NOR3_X1    g0998(.A1(new_n825_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1262_));
  NOR4_X1    g0999(.A1(new_n1259_), .A2(new_n1261_), .A3(new_n1260_), .A4(new_n1262_), .ZN(new_n1263_));
  OAI22_X1   g1000(.A1(new_n557_), .A2(new_n1258_), .B1(new_n1263_), .B2(new_n304_), .ZN(new_n1264_));
  OAI21_X1   g1001(.A1(new_n1253_), .A2(new_n1264_), .B(new_n340_), .ZN(new_n1265_));
  NAND2_X1   g1002(.A1(new_n1240_), .A2(new_n1265_), .ZN(new_n1266_));
  OAI21_X1   g1003(.A1(new_n1266_), .A2(new_n1217_), .B(\shift[6] ), .ZN(new_n1267_));
  NAND2_X1   g1004(.A1(new_n1157_), .A2(new_n1267_), .ZN(\result[3] ));
  NOR2_X1    g1005(.A1(new_n330_), .A2(new_n327_), .ZN(new_n1269_));
  OAI22_X1   g1006(.A1(new_n272_), .A2(new_n285_), .B1(new_n1269_), .B2(new_n274_), .ZN(new_n1270_));
  OAI21_X1   g1007(.A1(new_n298_), .A2(new_n301_), .B(new_n294_), .ZN(new_n1271_));
  OAI21_X1   g1008(.A1(new_n282_), .A2(new_n304_), .B(new_n1271_), .ZN(new_n1272_));
  OAI21_X1   g1009(.A1(new_n1270_), .A2(new_n1272_), .B(new_n308_), .ZN(new_n1273_));
  NOR2_X1    g1010(.A1(new_n395_), .A2(new_n392_), .ZN(new_n1274_));
  OAI22_X1   g1011(.A1(new_n274_), .A2(new_n1274_), .B1(new_n316_), .B2(new_n285_), .ZN(new_n1275_));
  OAI21_X1   g1012(.A1(new_n334_), .A2(new_n337_), .B(new_n294_), .ZN(new_n1276_));
  OAI21_X1   g1013(.A1(new_n319_), .A2(new_n322_), .B(new_n303_), .ZN(new_n1277_));
  NAND2_X1   g1014(.A1(new_n1276_), .A2(new_n1277_), .ZN(new_n1278_));
  OAI21_X1   g1015(.A1(new_n1275_), .A2(new_n1278_), .B(new_n340_), .ZN(new_n1279_));
  NAND2_X1   g1016(.A1(new_n1273_), .A2(new_n1279_), .ZN(new_n1280_));
  OAI21_X1   g1017(.A1(new_n429_), .A2(new_n426_), .B(new_n273_), .ZN(new_n1281_));
  OAI21_X1   g1018(.A1(new_n345_), .A2(new_n348_), .B(new_n284_), .ZN(new_n1282_));
  NAND2_X1   g1019(.A1(new_n1282_), .A2(new_n1281_), .ZN(new_n1283_));
  OAI21_X1   g1020(.A1(new_n370_), .A2(new_n367_), .B(new_n294_), .ZN(new_n1284_));
  OAI21_X1   g1021(.A1(new_n355_), .A2(new_n352_), .B(new_n303_), .ZN(new_n1285_));
  NAND2_X1   g1022(.A1(new_n1284_), .A2(new_n1285_), .ZN(new_n1286_));
  OAI21_X1   g1023(.A1(new_n1283_), .A2(new_n1286_), .B(new_n373_), .ZN(new_n1287_));
  OAI21_X1   g1024(.A1(new_n363_), .A2(new_n360_), .B(new_n273_), .ZN(new_n1288_));
  OAI21_X1   g1025(.A1(new_n380_), .A2(new_n377_), .B(new_n284_), .ZN(new_n1289_));
  NAND2_X1   g1026(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_));
  OAI21_X1   g1027(.A1(new_n402_), .A2(new_n399_), .B(new_n294_), .ZN(new_n1291_));
  OAI21_X1   g1028(.A1(new_n387_), .A2(new_n384_), .B(new_n303_), .ZN(new_n1292_));
  NAND2_X1   g1029(.A1(new_n1291_), .A2(new_n1292_), .ZN(new_n1293_));
  OAI21_X1   g1030(.A1(new_n1290_), .A2(new_n1293_), .B(new_n405_), .ZN(new_n1294_));
  NAND2_X1   g1031(.A1(new_n1287_), .A2(new_n1294_), .ZN(new_n1295_));
  OAI21_X1   g1032(.A1(new_n1280_), .A2(new_n1295_), .B(new_n264_), .ZN(new_n1296_));
  OAI21_X1   g1033(.A1(new_n489_), .A2(new_n492_), .B(new_n273_), .ZN(new_n1297_));
  OAI21_X1   g1034(.A1(new_n505_), .A2(new_n508_), .B(new_n284_), .ZN(new_n1298_));
  NAND2_X1   g1035(.A1(new_n1297_), .A2(new_n1298_), .ZN(new_n1299_));
  OAI21_X1   g1036(.A1(new_n530_), .A2(new_n527_), .B(new_n294_), .ZN(new_n1300_));
  OAI21_X1   g1037(.A1(new_n515_), .A2(new_n512_), .B(new_n303_), .ZN(new_n1301_));
  NAND2_X1   g1038(.A1(new_n1300_), .A2(new_n1301_), .ZN(new_n1302_));
  OAI21_X1   g1039(.A1(new_n1299_), .A2(new_n1302_), .B(new_n405_), .ZN(new_n1303_));
  OAI21_X1   g1040(.A1(new_n289_), .A2(new_n292_), .B(new_n273_), .ZN(new_n1304_));
  OAI21_X1   g1041(.A1(new_n474_), .A2(new_n477_), .B(new_n284_), .ZN(new_n1305_));
  NAND2_X1   g1042(.A1(new_n1304_), .A2(new_n1305_), .ZN(new_n1306_));
  OAI21_X1   g1043(.A1(new_n496_), .A2(new_n499_), .B(new_n294_), .ZN(new_n1307_));
  OAI21_X1   g1044(.A1(new_n484_), .A2(new_n481_), .B(new_n303_), .ZN(new_n1308_));
  NAND2_X1   g1045(.A1(new_n1307_), .A2(new_n1308_), .ZN(new_n1309_));
  OAI21_X1   g1046(.A1(new_n1306_), .A2(new_n1309_), .B(new_n373_), .ZN(new_n1310_));
  NAND2_X1   g1047(.A1(new_n1303_), .A2(new_n1310_), .ZN(new_n1311_));
  NOR2_X1    g1048(.A1(new_n445_), .A2(new_n442_), .ZN(new_n1312_));
  NOR2_X1    g1049(.A1(new_n523_), .A2(new_n520_), .ZN(new_n1313_));
  OAI22_X1   g1050(.A1(new_n274_), .A2(new_n1313_), .B1(new_n1312_), .B2(new_n285_), .ZN(new_n1314_));
  OAI21_X1   g1051(.A1(new_n467_), .A2(new_n464_), .B(new_n294_), .ZN(new_n1315_));
  OAI21_X1   g1052(.A1(new_n449_), .A2(new_n452_), .B(new_n303_), .ZN(new_n1316_));
  NAND2_X1   g1053(.A1(new_n1316_), .A2(new_n1315_), .ZN(new_n1317_));
  OAI21_X1   g1054(.A1(new_n1314_), .A2(new_n1317_), .B(new_n340_), .ZN(new_n1318_));
  OAI21_X1   g1055(.A1(new_n460_), .A2(new_n457_), .B(new_n273_), .ZN(new_n1319_));
  OAI21_X1   g1056(.A1(new_n414_), .A2(new_n411_), .B(new_n284_), .ZN(new_n1320_));
  NAND2_X1   g1057(.A1(new_n1319_), .A2(new_n1320_), .ZN(new_n1321_));
  OAI21_X1   g1058(.A1(new_n436_), .A2(new_n433_), .B(new_n294_), .ZN(new_n1322_));
  OAI21_X1   g1059(.A1(new_n421_), .A2(new_n418_), .B(new_n303_), .ZN(new_n1323_));
  NAND2_X1   g1060(.A1(new_n1322_), .A2(new_n1323_), .ZN(new_n1324_));
  OAI21_X1   g1061(.A1(new_n1321_), .A2(new_n1324_), .B(new_n308_), .ZN(new_n1325_));
  NAND2_X1   g1062(.A1(new_n1318_), .A2(new_n1325_), .ZN(new_n1326_));
  OAI21_X1   g1063(.A1(new_n1311_), .A2(new_n1326_), .B(\shift[6] ), .ZN(new_n1327_));
  NAND2_X1   g1064(.A1(new_n1296_), .A2(new_n1327_), .ZN(\result[4] ));
  OAI22_X1   g1065(.A1(new_n274_), .A2(new_n605_), .B1(new_n546_), .B2(new_n285_), .ZN(new_n1329_));
  OAI22_X1   g1066(.A1(new_n557_), .A2(new_n575_), .B1(new_n555_), .B2(new_n304_), .ZN(new_n1330_));
  NOR2_X1    g1067(.A1(new_n1329_), .A2(new_n1330_), .ZN(new_n1331_));
  OAI22_X1   g1068(.A1(new_n274_), .A2(new_n684_), .B1(new_n586_), .B2(new_n285_), .ZN(new_n1332_));
  OAI22_X1   g1069(.A1(new_n557_), .A2(new_n614_), .B1(new_n595_), .B2(new_n304_), .ZN(new_n1333_));
  OAI21_X1   g1070(.A1(new_n1332_), .A2(new_n1333_), .B(new_n340_), .ZN(new_n1334_));
  OAI21_X1   g1071(.A1(new_n537_), .A2(new_n1331_), .B(new_n1334_), .ZN(new_n1335_));
  OAI22_X1   g1072(.A1(new_n274_), .A2(new_n764_), .B1(new_n626_), .B2(new_n285_), .ZN(new_n1336_));
  OAI22_X1   g1073(.A1(new_n557_), .A2(new_n654_), .B1(new_n635_), .B2(new_n304_), .ZN(new_n1337_));
  OAI21_X1   g1074(.A1(new_n1336_), .A2(new_n1337_), .B(new_n373_), .ZN(new_n1338_));
  OAI22_X1   g1075(.A1(new_n274_), .A2(new_n645_), .B1(new_n665_), .B2(new_n285_), .ZN(new_n1339_));
  OAI22_X1   g1076(.A1(new_n557_), .A2(new_n693_), .B1(new_n674_), .B2(new_n304_), .ZN(new_n1340_));
  OAI21_X1   g1077(.A1(new_n1339_), .A2(new_n1340_), .B(new_n405_), .ZN(new_n1341_));
  NAND2_X1   g1078(.A1(new_n1338_), .A2(new_n1341_), .ZN(new_n1342_));
  OAI21_X1   g1079(.A1(new_n1335_), .A2(new_n1342_), .B(new_n264_), .ZN(new_n1343_));
  OAI22_X1   g1080(.A1(new_n274_), .A2(new_n725_), .B1(new_n785_), .B2(new_n285_), .ZN(new_n1344_));
  OAI21_X1   g1081(.A1(new_n803_), .A2(new_n806_), .B(new_n294_), .ZN(new_n1345_));
  OAI21_X1   g1082(.A1(new_n791_), .A2(new_n788_), .B(new_n303_), .ZN(new_n1346_));
  NAND2_X1   g1083(.A1(new_n1345_), .A2(new_n1346_), .ZN(new_n1347_));
  OAI21_X1   g1084(.A1(new_n1344_), .A2(new_n1347_), .B(new_n405_), .ZN(new_n1348_));
  OAI22_X1   g1085(.A1(new_n274_), .A2(new_n566_), .B1(new_n706_), .B2(new_n285_), .ZN(new_n1349_));
  OAI22_X1   g1086(.A1(new_n557_), .A2(new_n734_), .B1(new_n715_), .B2(new_n304_), .ZN(new_n1350_));
  OAI21_X1   g1087(.A1(new_n1349_), .A2(new_n1350_), .B(new_n373_), .ZN(new_n1351_));
  NAND2_X1   g1088(.A1(new_n1351_), .A2(new_n1348_), .ZN(new_n1352_));
  NOR3_X1    g1089(.A1(new_n1197_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1353_));
  INV_X1     g1090(.I(new_n795_), .ZN(new_n1354_));
  NOR2_X1    g1091(.A1(new_n1201_), .A2(\shift[1] ), .ZN(new_n1355_));
  NOR3_X1    g1092(.A1(new_n1245_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1356_));
  NOR4_X1    g1093(.A1(new_n1354_), .A2(new_n1355_), .A3(new_n1356_), .A4(new_n1353_), .ZN(new_n1357_));
  OAI22_X1   g1094(.A1(new_n274_), .A2(new_n1357_), .B1(new_n818_), .B2(new_n285_), .ZN(new_n1358_));
  OAI22_X1   g1095(.A1(new_n557_), .A2(new_n846_), .B1(new_n827_), .B2(new_n304_), .ZN(new_n1359_));
  OAI21_X1   g1096(.A1(new_n1358_), .A2(new_n1359_), .B(new_n340_), .ZN(new_n1360_));
  OAI22_X1   g1097(.A1(new_n274_), .A2(new_n837_), .B1(new_n745_), .B2(new_n285_), .ZN(new_n1361_));
  OAI22_X1   g1098(.A1(new_n557_), .A2(new_n773_), .B1(new_n754_), .B2(new_n304_), .ZN(new_n1362_));
  OAI21_X1   g1099(.A1(new_n1361_), .A2(new_n1362_), .B(new_n308_), .ZN(new_n1363_));
  NAND2_X1   g1100(.A1(new_n1360_), .A2(new_n1363_), .ZN(new_n1364_));
  OAI21_X1   g1101(.A1(new_n1364_), .A2(new_n1352_), .B(\shift[6] ), .ZN(new_n1365_));
  NAND2_X1   g1102(.A1(new_n1343_), .A2(new_n1365_), .ZN(\result[5] ));
  NOR2_X1    g1103(.A1(new_n886_), .A2(new_n889_), .ZN(new_n1367_));
  OAI22_X1   g1104(.A1(new_n274_), .A2(new_n1367_), .B1(new_n858_), .B2(new_n285_), .ZN(new_n1368_));
  OAI21_X1   g1105(.A1(new_n868_), .A2(new_n869_), .B(new_n294_), .ZN(new_n1369_));
  OAI21_X1   g1106(.A1(new_n304_), .A2(new_n863_), .B(new_n1369_), .ZN(new_n1370_));
  OAI21_X1   g1107(.A1(new_n1368_), .A2(new_n1370_), .B(new_n308_), .ZN(new_n1371_));
  NOR2_X1    g1108(.A1(new_n875_), .A2(new_n878_), .ZN(new_n1372_));
  NOR2_X1    g1109(.A1(new_n945_), .A2(new_n948_), .ZN(new_n1373_));
  OAI22_X1   g1110(.A1(new_n274_), .A2(new_n1373_), .B1(new_n1372_), .B2(new_n285_), .ZN(new_n1374_));
  OAI21_X1   g1111(.A1(new_n891_), .A2(new_n894_), .B(new_n294_), .ZN(new_n1375_));
  OAI21_X1   g1112(.A1(new_n882_), .A2(new_n883_), .B(new_n303_), .ZN(new_n1376_));
  NAND2_X1   g1113(.A1(new_n1376_), .A2(new_n1375_), .ZN(new_n1377_));
  OAI21_X1   g1114(.A1(new_n1374_), .A2(new_n1377_), .B(new_n340_), .ZN(new_n1378_));
  NAND2_X1   g1115(.A1(new_n1371_), .A2(new_n1378_), .ZN(new_n1379_));
  OAI21_X1   g1116(.A1(new_n997_), .A2(new_n1000_), .B(new_n273_), .ZN(new_n1380_));
  OAI21_X1   g1117(.A1(new_n901_), .A2(new_n904_), .B(new_n284_), .ZN(new_n1381_));
  NAND2_X1   g1118(.A1(new_n1380_), .A2(new_n1381_), .ZN(new_n1382_));
  OAI21_X1   g1119(.A1(new_n921_), .A2(new_n924_), .B(new_n294_), .ZN(new_n1383_));
  OAI21_X1   g1120(.A1(new_n906_), .A2(new_n909_), .B(new_n303_), .ZN(new_n1384_));
  NAND2_X1   g1121(.A1(new_n1383_), .A2(new_n1384_), .ZN(new_n1385_));
  OAI21_X1   g1122(.A1(new_n1382_), .A2(new_n1385_), .B(new_n373_), .ZN(new_n1386_));
  OAI21_X1   g1123(.A1(new_n914_), .A2(new_n917_), .B(new_n273_), .ZN(new_n1387_));
  OAI21_X1   g1124(.A1(new_n930_), .A2(new_n933_), .B(new_n284_), .ZN(new_n1388_));
  NAND2_X1   g1125(.A1(new_n1387_), .A2(new_n1388_), .ZN(new_n1389_));
  OAI21_X1   g1126(.A1(new_n952_), .A2(new_n955_), .B(new_n294_), .ZN(new_n1390_));
  OAI21_X1   g1127(.A1(new_n937_), .A2(new_n940_), .B(new_n303_), .ZN(new_n1391_));
  NAND2_X1   g1128(.A1(new_n1390_), .A2(new_n1391_), .ZN(new_n1392_));
  OAI21_X1   g1129(.A1(new_n1389_), .A2(new_n1392_), .B(new_n405_), .ZN(new_n1393_));
  NAND2_X1   g1130(.A1(new_n1386_), .A2(new_n1393_), .ZN(new_n1394_));
  OAI21_X1   g1131(.A1(new_n1379_), .A2(new_n1394_), .B(new_n264_), .ZN(new_n1395_));
  OAI21_X1   g1132(.A1(new_n970_), .A2(new_n971_), .B(new_n273_), .ZN(new_n1396_));
  OAI21_X1   g1133(.A1(new_n1012_), .A2(new_n1013_), .B(new_n284_), .ZN(new_n1397_));
  NAND2_X1   g1134(.A1(new_n1396_), .A2(new_n1397_), .ZN(new_n1398_));
  OAI21_X1   g1135(.A1(new_n1028_), .A2(new_n1030_), .B(new_n294_), .ZN(new_n1399_));
  OAI21_X1   g1136(.A1(new_n1018_), .A2(new_n1017_), .B(new_n303_), .ZN(new_n1400_));
  NAND2_X1   g1137(.A1(new_n1399_), .A2(new_n1400_), .ZN(new_n1401_));
  OAI21_X1   g1138(.A1(new_n1398_), .A2(new_n1401_), .B(new_n405_), .ZN(new_n1402_));
  OAI21_X1   g1139(.A1(new_n865_), .A2(new_n866_), .B(new_n273_), .ZN(new_n1403_));
  OAI21_X1   g1140(.A1(new_n961_), .A2(new_n962_), .B(new_n284_), .ZN(new_n1404_));
  NAND2_X1   g1141(.A1(new_n1403_), .A2(new_n1404_), .ZN(new_n1405_));
  OAI21_X1   g1142(.A1(new_n975_), .A2(new_n976_), .B(new_n294_), .ZN(new_n1406_));
  OAI21_X1   g1143(.A1(new_n964_), .A2(new_n967_), .B(new_n303_), .ZN(new_n1407_));
  NAND2_X1   g1144(.A1(new_n1406_), .A2(new_n1407_), .ZN(new_n1408_));
  OAI21_X1   g1145(.A1(new_n1405_), .A2(new_n1408_), .B(new_n373_), .ZN(new_n1409_));
  NAND2_X1   g1146(.A1(new_n1402_), .A2(new_n1409_), .ZN(new_n1410_));
  OAI21_X1   g1147(.A1(new_n1023_), .A2(new_n1024_), .B(new_n273_), .ZN(new_n1411_));
  OAI21_X1   g1148(.A1(new_n1036_), .A2(new_n1037_), .B(new_n284_), .ZN(new_n1412_));
  NAND2_X1   g1149(.A1(new_n1411_), .A2(new_n1412_), .ZN(new_n1413_));
  OAI21_X1   g1150(.A1(new_n1052_), .A2(new_n1055_), .B(new_n294_), .ZN(new_n1414_));
  OAI21_X1   g1151(.A1(new_n1041_), .A2(new_n1042_), .B(new_n303_), .ZN(new_n1415_));
  NAND2_X1   g1152(.A1(new_n1415_), .A2(new_n1414_), .ZN(new_n1416_));
  OAI21_X1   g1153(.A1(new_n1413_), .A2(new_n1416_), .B(new_n340_), .ZN(new_n1417_));
  OAI21_X1   g1154(.A1(new_n1047_), .A2(new_n1050_), .B(new_n273_), .ZN(new_n1418_));
  OAI21_X1   g1155(.A1(new_n982_), .A2(new_n985_), .B(new_n284_), .ZN(new_n1419_));
  NAND2_X1   g1156(.A1(new_n1418_), .A2(new_n1419_), .ZN(new_n1420_));
  OAI21_X1   g1157(.A1(new_n1004_), .A2(new_n1007_), .B(new_n294_), .ZN(new_n1421_));
  OAI21_X1   g1158(.A1(new_n989_), .A2(new_n992_), .B(new_n303_), .ZN(new_n1422_));
  NAND2_X1   g1159(.A1(new_n1421_), .A2(new_n1422_), .ZN(new_n1423_));
  OAI21_X1   g1160(.A1(new_n1420_), .A2(new_n1423_), .B(new_n308_), .ZN(new_n1424_));
  NAND2_X1   g1161(.A1(new_n1417_), .A2(new_n1424_), .ZN(new_n1425_));
  OAI21_X1   g1162(.A1(new_n1410_), .A2(new_n1425_), .B(\shift[6] ), .ZN(new_n1426_));
  NAND2_X1   g1163(.A1(new_n1395_), .A2(new_n1426_), .ZN(\result[6] ));
  OAI22_X1   g1164(.A1(new_n274_), .A2(new_n1101_), .B1(new_n1137_), .B2(new_n285_), .ZN(new_n1428_));
  OAI22_X1   g1165(.A1(new_n557_), .A2(new_n1153_), .B1(new_n1142_), .B2(new_n304_), .ZN(new_n1429_));
  NOR2_X1    g1166(.A1(new_n1428_), .A2(new_n1429_), .ZN(new_n1430_));
  OAI22_X1   g1167(.A1(new_n274_), .A2(new_n1078_), .B1(new_n1090_), .B2(new_n285_), .ZN(new_n1431_));
  OAI22_X1   g1168(.A1(new_n557_), .A2(new_n1106_), .B1(new_n1095_), .B2(new_n304_), .ZN(new_n1432_));
  OAI21_X1   g1169(.A1(new_n1431_), .A2(new_n1432_), .B(new_n340_), .ZN(new_n1433_));
  OAI21_X1   g1170(.A1(new_n537_), .A2(new_n1430_), .B(new_n1433_), .ZN(new_n1434_));
  OAI22_X1   g1171(.A1(new_n274_), .A2(new_n1233_), .B1(new_n1114_), .B2(new_n285_), .ZN(new_n1435_));
  OAI22_X1   g1172(.A1(new_n557_), .A2(new_n1130_), .B1(new_n1119_), .B2(new_n304_), .ZN(new_n1436_));
  OAI21_X1   g1173(.A1(new_n1435_), .A2(new_n1436_), .B(new_n373_), .ZN(new_n1437_));
  OAI22_X1   g1174(.A1(new_n274_), .A2(new_n1125_), .B1(new_n1067_), .B2(new_n285_), .ZN(new_n1438_));
  OAI22_X1   g1175(.A1(new_n557_), .A2(new_n1083_), .B1(new_n1072_), .B2(new_n304_), .ZN(new_n1439_));
  OAI21_X1   g1176(.A1(new_n1438_), .A2(new_n1439_), .B(new_n405_), .ZN(new_n1440_));
  NAND2_X1   g1177(.A1(new_n1437_), .A2(new_n1440_), .ZN(new_n1441_));
  OAI21_X1   g1178(.A1(new_n1434_), .A2(new_n1441_), .B(new_n264_), .ZN(new_n1442_));
  OAI21_X1   g1179(.A1(new_n1184_), .A2(new_n1187_), .B(new_n284_), .ZN(new_n1443_));
  OAI21_X1   g1180(.A1(new_n1194_), .A2(new_n1191_), .B(new_n303_), .ZN(new_n1444_));
  NAND2_X1   g1181(.A1(new_n1443_), .A2(new_n1444_), .ZN(new_n1445_));
  OAI22_X1   g1182(.A1(new_n274_), .A2(new_n1174_), .B1(new_n1214_), .B2(new_n557_), .ZN(new_n1446_));
  OAI21_X1   g1183(.A1(new_n1446_), .A2(new_n1445_), .B(new_n405_), .ZN(new_n1447_));
  OAI22_X1   g1184(.A1(new_n274_), .A2(new_n1148_), .B1(new_n1162_), .B2(new_n285_), .ZN(new_n1448_));
  OAI22_X1   g1185(.A1(new_n557_), .A2(new_n1179_), .B1(new_n1167_), .B2(new_n304_), .ZN(new_n1449_));
  OAI21_X1   g1186(.A1(new_n1448_), .A2(new_n1449_), .B(new_n373_), .ZN(new_n1450_));
  NAND2_X1   g1187(.A1(new_n1450_), .A2(new_n1447_), .ZN(new_n1451_));
  OAI22_X1   g1188(.A1(new_n274_), .A2(new_n1205_), .B1(new_n1247_), .B2(new_n285_), .ZN(new_n1452_));
  OAI22_X1   g1189(.A1(new_n557_), .A2(new_n1263_), .B1(new_n1252_), .B2(new_n304_), .ZN(new_n1453_));
  OAI21_X1   g1190(.A1(new_n1452_), .A2(new_n1453_), .B(new_n340_), .ZN(new_n1454_));
  OAI22_X1   g1191(.A1(new_n274_), .A2(new_n1258_), .B1(new_n1222_), .B2(new_n285_), .ZN(new_n1455_));
  OAI22_X1   g1192(.A1(new_n557_), .A2(new_n1238_), .B1(new_n1227_), .B2(new_n304_), .ZN(new_n1456_));
  OAI21_X1   g1193(.A1(new_n1455_), .A2(new_n1456_), .B(new_n308_), .ZN(new_n1457_));
  NAND2_X1   g1194(.A1(new_n1454_), .A2(new_n1457_), .ZN(new_n1458_));
  OAI21_X1   g1195(.A1(new_n1458_), .A2(new_n1451_), .B(\shift[6] ), .ZN(new_n1459_));
  NAND2_X1   g1196(.A1(new_n1442_), .A2(new_n1459_), .ZN(\result[7] ));
  OAI21_X1   g1197(.A1(new_n334_), .A2(new_n337_), .B(new_n273_), .ZN(new_n1461_));
  OAI21_X1   g1198(.A1(new_n330_), .A2(new_n327_), .B(new_n284_), .ZN(new_n1462_));
  NAND2_X1   g1199(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1463_));
  OAI21_X1   g1200(.A1(new_n278_), .A2(new_n281_), .B(new_n294_), .ZN(new_n1464_));
  OAI21_X1   g1201(.A1(new_n271_), .A2(new_n268_), .B(new_n303_), .ZN(new_n1465_));
  NAND2_X1   g1202(.A1(new_n1464_), .A2(new_n1465_), .ZN(new_n1466_));
  OAI21_X1   g1203(.A1(new_n1463_), .A2(new_n1466_), .B(new_n308_), .ZN(new_n1467_));
  OAI21_X1   g1204(.A1(new_n402_), .A2(new_n399_), .B(new_n273_), .ZN(new_n1468_));
  OAI21_X1   g1205(.A1(new_n395_), .A2(new_n392_), .B(new_n284_), .ZN(new_n1469_));
  NAND2_X1   g1206(.A1(new_n1468_), .A2(new_n1469_), .ZN(new_n1470_));
  OAI21_X1   g1207(.A1(new_n319_), .A2(new_n322_), .B(new_n294_), .ZN(new_n1471_));
  OAI21_X1   g1208(.A1(new_n315_), .A2(new_n312_), .B(new_n303_), .ZN(new_n1472_));
  NAND2_X1   g1209(.A1(new_n1471_), .A2(new_n1472_), .ZN(new_n1473_));
  OAI21_X1   g1210(.A1(new_n1470_), .A2(new_n1473_), .B(new_n340_), .ZN(new_n1474_));
  NAND2_X1   g1211(.A1(new_n1467_), .A2(new_n1474_), .ZN(new_n1475_));
  NOR2_X1    g1212(.A1(new_n429_), .A2(new_n426_), .ZN(new_n1476_));
  NOR2_X1    g1213(.A1(new_n436_), .A2(new_n433_), .ZN(new_n1477_));
  OAI22_X1   g1214(.A1(new_n274_), .A2(new_n1477_), .B1(new_n1476_), .B2(new_n285_), .ZN(new_n1478_));
  OAI21_X1   g1215(.A1(new_n355_), .A2(new_n352_), .B(new_n294_), .ZN(new_n1479_));
  OAI21_X1   g1216(.A1(new_n345_), .A2(new_n348_), .B(new_n303_), .ZN(new_n1480_));
  NAND2_X1   g1217(.A1(new_n1480_), .A2(new_n1479_), .ZN(new_n1481_));
  OAI21_X1   g1218(.A1(new_n1478_), .A2(new_n1481_), .B(new_n373_), .ZN(new_n1482_));
  OAI21_X1   g1219(.A1(new_n370_), .A2(new_n367_), .B(new_n273_), .ZN(new_n1483_));
  OAI21_X1   g1220(.A1(new_n363_), .A2(new_n360_), .B(new_n284_), .ZN(new_n1484_));
  NAND2_X1   g1221(.A1(new_n1483_), .A2(new_n1484_), .ZN(new_n1485_));
  OAI21_X1   g1222(.A1(new_n387_), .A2(new_n384_), .B(new_n294_), .ZN(new_n1486_));
  OAI21_X1   g1223(.A1(new_n380_), .A2(new_n377_), .B(new_n303_), .ZN(new_n1487_));
  NAND2_X1   g1224(.A1(new_n1486_), .A2(new_n1487_), .ZN(new_n1488_));
  OAI21_X1   g1225(.A1(new_n1485_), .A2(new_n1488_), .B(new_n405_), .ZN(new_n1489_));
  NAND2_X1   g1226(.A1(new_n1482_), .A2(new_n1489_), .ZN(new_n1490_));
  OAI21_X1   g1227(.A1(new_n1475_), .A2(new_n1490_), .B(new_n264_), .ZN(new_n1491_));
  NOR2_X1    g1228(.A1(new_n489_), .A2(new_n492_), .ZN(new_n1492_));
  NOR2_X1    g1229(.A1(new_n496_), .A2(new_n499_), .ZN(new_n1493_));
  OAI22_X1   g1230(.A1(new_n274_), .A2(new_n1493_), .B1(new_n1492_), .B2(new_n285_), .ZN(new_n1494_));
  NOR2_X1    g1231(.A1(new_n505_), .A2(new_n508_), .ZN(new_n1495_));
  NOR2_X1    g1232(.A1(new_n515_), .A2(new_n512_), .ZN(new_n1496_));
  OAI22_X1   g1233(.A1(new_n304_), .A2(new_n1495_), .B1(new_n1496_), .B2(new_n557_), .ZN(new_n1497_));
  OAI21_X1   g1234(.A1(new_n1494_), .A2(new_n1497_), .B(new_n405_), .ZN(new_n1498_));
  OAI21_X1   g1235(.A1(new_n289_), .A2(new_n292_), .B(new_n284_), .ZN(new_n1499_));
  OAI21_X1   g1236(.A1(new_n274_), .A2(new_n302_), .B(new_n1499_), .ZN(new_n1500_));
  OAI21_X1   g1237(.A1(new_n484_), .A2(new_n481_), .B(new_n294_), .ZN(new_n1501_));
  OAI21_X1   g1238(.A1(new_n474_), .A2(new_n477_), .B(new_n303_), .ZN(new_n1502_));
  NAND2_X1   g1239(.A1(new_n1502_), .A2(new_n1501_), .ZN(new_n1503_));
  OAI21_X1   g1240(.A1(new_n1500_), .A2(new_n1503_), .B(new_n373_), .ZN(new_n1504_));
  NAND2_X1   g1241(.A1(new_n1498_), .A2(new_n1504_), .ZN(new_n1505_));
  OAI21_X1   g1242(.A1(new_n530_), .A2(new_n527_), .B(new_n273_), .ZN(new_n1506_));
  OAI21_X1   g1243(.A1(new_n523_), .A2(new_n520_), .B(new_n284_), .ZN(new_n1507_));
  NAND2_X1   g1244(.A1(new_n1506_), .A2(new_n1507_), .ZN(new_n1508_));
  OAI21_X1   g1245(.A1(new_n449_), .A2(new_n452_), .B(new_n294_), .ZN(new_n1509_));
  OAI21_X1   g1246(.A1(new_n445_), .A2(new_n442_), .B(new_n303_), .ZN(new_n1510_));
  NAND2_X1   g1247(.A1(new_n1509_), .A2(new_n1510_), .ZN(new_n1511_));
  OAI21_X1   g1248(.A1(new_n1508_), .A2(new_n1511_), .B(new_n340_), .ZN(new_n1512_));
  OAI21_X1   g1249(.A1(new_n467_), .A2(new_n464_), .B(new_n273_), .ZN(new_n1513_));
  OAI21_X1   g1250(.A1(new_n460_), .A2(new_n457_), .B(new_n284_), .ZN(new_n1514_));
  NAND2_X1   g1251(.A1(new_n1513_), .A2(new_n1514_), .ZN(new_n1515_));
  OAI21_X1   g1252(.A1(new_n421_), .A2(new_n418_), .B(new_n294_), .ZN(new_n1516_));
  OAI21_X1   g1253(.A1(new_n414_), .A2(new_n411_), .B(new_n303_), .ZN(new_n1517_));
  NAND2_X1   g1254(.A1(new_n1516_), .A2(new_n1517_), .ZN(new_n1518_));
  OAI21_X1   g1255(.A1(new_n1515_), .A2(new_n1518_), .B(new_n308_), .ZN(new_n1519_));
  NAND2_X1   g1256(.A1(new_n1512_), .A2(new_n1519_), .ZN(new_n1520_));
  OAI21_X1   g1257(.A1(new_n1505_), .A2(new_n1520_), .B(\shift[6] ), .ZN(new_n1521_));
  NAND2_X1   g1258(.A1(new_n1491_), .A2(new_n1521_), .ZN(\result[8] ));
  OAI22_X1   g1259(.A1(new_n274_), .A2(new_n614_), .B1(new_n605_), .B2(new_n285_), .ZN(new_n1523_));
  OAI22_X1   g1260(.A1(new_n557_), .A2(new_n555_), .B1(new_n546_), .B2(new_n304_), .ZN(new_n1524_));
  OAI21_X1   g1261(.A1(new_n1523_), .A2(new_n1524_), .B(new_n308_), .ZN(new_n1525_));
  OAI22_X1   g1262(.A1(new_n274_), .A2(new_n693_), .B1(new_n684_), .B2(new_n285_), .ZN(new_n1526_));
  OAI22_X1   g1263(.A1(new_n557_), .A2(new_n595_), .B1(new_n586_), .B2(new_n304_), .ZN(new_n1527_));
  OAI21_X1   g1264(.A1(new_n1526_), .A2(new_n1527_), .B(new_n340_), .ZN(new_n1528_));
  NAND2_X1   g1265(.A1(new_n1525_), .A2(new_n1528_), .ZN(new_n1529_));
  OAI22_X1   g1266(.A1(new_n274_), .A2(new_n773_), .B1(new_n764_), .B2(new_n285_), .ZN(new_n1530_));
  OAI22_X1   g1267(.A1(new_n557_), .A2(new_n635_), .B1(new_n626_), .B2(new_n304_), .ZN(new_n1531_));
  OAI21_X1   g1268(.A1(new_n1530_), .A2(new_n1531_), .B(new_n373_), .ZN(new_n1532_));
  OAI22_X1   g1269(.A1(new_n274_), .A2(new_n654_), .B1(new_n645_), .B2(new_n285_), .ZN(new_n1533_));
  OAI22_X1   g1270(.A1(new_n557_), .A2(new_n674_), .B1(new_n665_), .B2(new_n304_), .ZN(new_n1534_));
  OAI21_X1   g1271(.A1(new_n1533_), .A2(new_n1534_), .B(new_n405_), .ZN(new_n1535_));
  NAND2_X1   g1272(.A1(new_n1532_), .A2(new_n1535_), .ZN(new_n1536_));
  OAI21_X1   g1273(.A1(new_n1529_), .A2(new_n1536_), .B(new_n264_), .ZN(new_n1537_));
  OAI22_X1   g1274(.A1(new_n274_), .A2(new_n734_), .B1(new_n725_), .B2(new_n285_), .ZN(new_n1538_));
  OAI21_X1   g1275(.A1(new_n791_), .A2(new_n788_), .B(new_n294_), .ZN(new_n1539_));
  NAND2_X1   g1276(.A1(new_n266_), .A2(\a[49] ), .ZN(new_n1540_));
  OAI21_X1   g1277(.A1(new_n1540_), .A2(\shift[1] ), .B(new_n779_), .ZN(new_n1541_));
  NAND3_X1   g1278(.A1(new_n275_), .A2(\a[48] ), .A3(\shift[0] ), .ZN(new_n1542_));
  NAND3_X1   g1279(.A1(new_n266_), .A2(\a[47] ), .A3(\shift[1] ), .ZN(new_n1543_));
  NAND2_X1   g1280(.A1(new_n1542_), .A2(new_n1543_), .ZN(new_n1544_));
  OAI21_X1   g1281(.A1(new_n1544_), .A2(new_n1541_), .B(new_n303_), .ZN(new_n1545_));
  NAND2_X1   g1282(.A1(new_n1545_), .A2(new_n1539_), .ZN(new_n1546_));
  OAI21_X1   g1283(.A1(new_n1538_), .A2(new_n1546_), .B(new_n405_), .ZN(new_n1547_));
  OAI22_X1   g1284(.A1(new_n274_), .A2(new_n575_), .B1(new_n566_), .B2(new_n285_), .ZN(new_n1548_));
  OAI22_X1   g1285(.A1(new_n557_), .A2(new_n715_), .B1(new_n706_), .B2(new_n304_), .ZN(new_n1549_));
  OAI21_X1   g1286(.A1(new_n1548_), .A2(new_n1549_), .B(new_n373_), .ZN(new_n1550_));
  NAND2_X1   g1287(.A1(new_n1550_), .A2(new_n1547_), .ZN(new_n1551_));
  OAI21_X1   g1288(.A1(new_n803_), .A2(new_n806_), .B(new_n273_), .ZN(new_n1552_));
  OAI21_X1   g1289(.A1(new_n799_), .A2(new_n796_), .B(new_n284_), .ZN(new_n1553_));
  NAND2_X1   g1290(.A1(new_n1553_), .A2(new_n1552_), .ZN(new_n1554_));
  OAI22_X1   g1291(.A1(new_n557_), .A2(new_n827_), .B1(new_n818_), .B2(new_n304_), .ZN(new_n1555_));
  OAI21_X1   g1292(.A1(new_n1555_), .A2(new_n1554_), .B(new_n340_), .ZN(new_n1556_));
  OAI22_X1   g1293(.A1(new_n274_), .A2(new_n846_), .B1(new_n837_), .B2(new_n285_), .ZN(new_n1557_));
  OAI22_X1   g1294(.A1(new_n557_), .A2(new_n754_), .B1(new_n745_), .B2(new_n304_), .ZN(new_n1558_));
  OAI21_X1   g1295(.A1(new_n1557_), .A2(new_n1558_), .B(new_n308_), .ZN(new_n1559_));
  NAND2_X1   g1296(.A1(new_n1559_), .A2(new_n1556_), .ZN(new_n1560_));
  OAI21_X1   g1297(.A1(new_n1551_), .A2(new_n1560_), .B(\shift[6] ), .ZN(new_n1561_));
  NAND2_X1   g1298(.A1(new_n1537_), .A2(new_n1561_), .ZN(\result[9] ));
  OAI21_X1   g1299(.A1(new_n891_), .A2(new_n894_), .B(new_n273_), .ZN(new_n1563_));
  OAI21_X1   g1300(.A1(new_n886_), .A2(new_n889_), .B(new_n284_), .ZN(new_n1564_));
  NAND2_X1   g1301(.A1(new_n1563_), .A2(new_n1564_), .ZN(new_n1565_));
  OAI21_X1   g1302(.A1(new_n861_), .A2(new_n862_), .B(new_n294_), .ZN(new_n1566_));
  OAI21_X1   g1303(.A1(new_n854_), .A2(new_n857_), .B(new_n303_), .ZN(new_n1567_));
  NAND2_X1   g1304(.A1(new_n1566_), .A2(new_n1567_), .ZN(new_n1568_));
  OAI21_X1   g1305(.A1(new_n1565_), .A2(new_n1568_), .B(new_n308_), .ZN(new_n1569_));
  OAI21_X1   g1306(.A1(new_n952_), .A2(new_n955_), .B(new_n273_), .ZN(new_n1570_));
  OAI21_X1   g1307(.A1(new_n945_), .A2(new_n948_), .B(new_n284_), .ZN(new_n1571_));
  NAND2_X1   g1308(.A1(new_n1570_), .A2(new_n1571_), .ZN(new_n1572_));
  OAI21_X1   g1309(.A1(new_n882_), .A2(new_n883_), .B(new_n294_), .ZN(new_n1573_));
  OAI21_X1   g1310(.A1(new_n875_), .A2(new_n878_), .B(new_n303_), .ZN(new_n1574_));
  NAND2_X1   g1311(.A1(new_n1573_), .A2(new_n1574_), .ZN(new_n1575_));
  OAI21_X1   g1312(.A1(new_n1572_), .A2(new_n1575_), .B(new_n340_), .ZN(new_n1576_));
  NAND2_X1   g1313(.A1(new_n1569_), .A2(new_n1576_), .ZN(new_n1577_));
  OAI21_X1   g1314(.A1(new_n1004_), .A2(new_n1007_), .B(new_n273_), .ZN(new_n1578_));
  OAI21_X1   g1315(.A1(new_n997_), .A2(new_n1000_), .B(new_n284_), .ZN(new_n1579_));
  NAND2_X1   g1316(.A1(new_n1578_), .A2(new_n1579_), .ZN(new_n1580_));
  OAI21_X1   g1317(.A1(new_n906_), .A2(new_n909_), .B(new_n294_), .ZN(new_n1581_));
  OAI21_X1   g1318(.A1(new_n901_), .A2(new_n904_), .B(new_n303_), .ZN(new_n1582_));
  NAND2_X1   g1319(.A1(new_n1581_), .A2(new_n1582_), .ZN(new_n1583_));
  OAI21_X1   g1320(.A1(new_n1580_), .A2(new_n1583_), .B(new_n373_), .ZN(new_n1584_));
  OAI21_X1   g1321(.A1(new_n921_), .A2(new_n924_), .B(new_n273_), .ZN(new_n1585_));
  OAI21_X1   g1322(.A1(new_n914_), .A2(new_n917_), .B(new_n284_), .ZN(new_n1586_));
  NAND2_X1   g1323(.A1(new_n1585_), .A2(new_n1586_), .ZN(new_n1587_));
  OAI21_X1   g1324(.A1(new_n937_), .A2(new_n940_), .B(new_n294_), .ZN(new_n1588_));
  OAI21_X1   g1325(.A1(new_n930_), .A2(new_n933_), .B(new_n303_), .ZN(new_n1589_));
  NAND2_X1   g1326(.A1(new_n1588_), .A2(new_n1589_), .ZN(new_n1590_));
  OAI21_X1   g1327(.A1(new_n1587_), .A2(new_n1590_), .B(new_n405_), .ZN(new_n1591_));
  NAND2_X1   g1328(.A1(new_n1584_), .A2(new_n1591_), .ZN(new_n1592_));
  OAI21_X1   g1329(.A1(new_n1577_), .A2(new_n1592_), .B(new_n264_), .ZN(new_n1593_));
  NOR2_X1    g1330(.A1(new_n970_), .A2(new_n971_), .ZN(new_n1594_));
  OAI22_X1   g1331(.A1(new_n274_), .A2(new_n977_), .B1(new_n1594_), .B2(new_n285_), .ZN(new_n1595_));
  OAI22_X1   g1332(.A1(new_n304_), .A2(new_n1014_), .B1(new_n1019_), .B2(new_n557_), .ZN(new_n1596_));
  OAI21_X1   g1333(.A1(new_n1595_), .A2(new_n1596_), .B(new_n405_), .ZN(new_n1597_));
  NOR2_X1    g1334(.A1(new_n868_), .A2(new_n869_), .ZN(new_n1598_));
  OAI21_X1   g1335(.A1(new_n865_), .A2(new_n866_), .B(new_n284_), .ZN(new_n1599_));
  OAI21_X1   g1336(.A1(new_n274_), .A2(new_n1598_), .B(new_n1599_), .ZN(new_n1600_));
  OAI21_X1   g1337(.A1(new_n964_), .A2(new_n967_), .B(new_n294_), .ZN(new_n1601_));
  OAI21_X1   g1338(.A1(new_n961_), .A2(new_n962_), .B(new_n303_), .ZN(new_n1602_));
  NAND2_X1   g1339(.A1(new_n1602_), .A2(new_n1601_), .ZN(new_n1603_));
  OAI21_X1   g1340(.A1(new_n1600_), .A2(new_n1603_), .B(new_n373_), .ZN(new_n1604_));
  NAND2_X1   g1341(.A1(new_n1597_), .A2(new_n1604_), .ZN(new_n1605_));
  NOR2_X1    g1342(.A1(new_n1028_), .A2(new_n1030_), .ZN(new_n1606_));
  OAI21_X1   g1343(.A1(new_n1023_), .A2(new_n1024_), .B(new_n284_), .ZN(new_n1607_));
  OAI21_X1   g1344(.A1(new_n274_), .A2(new_n1606_), .B(new_n1607_), .ZN(new_n1608_));
  OAI21_X1   g1345(.A1(new_n1041_), .A2(new_n1042_), .B(new_n294_), .ZN(new_n1609_));
  OAI21_X1   g1346(.A1(new_n1036_), .A2(new_n1037_), .B(new_n303_), .ZN(new_n1610_));
  NAND2_X1   g1347(.A1(new_n1609_), .A2(new_n1610_), .ZN(new_n1611_));
  OAI21_X1   g1348(.A1(new_n1608_), .A2(new_n1611_), .B(new_n340_), .ZN(new_n1612_));
  OAI21_X1   g1349(.A1(new_n1052_), .A2(new_n1055_), .B(new_n273_), .ZN(new_n1613_));
  OAI21_X1   g1350(.A1(new_n1047_), .A2(new_n1050_), .B(new_n284_), .ZN(new_n1614_));
  NAND2_X1   g1351(.A1(new_n1613_), .A2(new_n1614_), .ZN(new_n1615_));
  OAI21_X1   g1352(.A1(new_n989_), .A2(new_n992_), .B(new_n294_), .ZN(new_n1616_));
  OAI21_X1   g1353(.A1(new_n982_), .A2(new_n985_), .B(new_n303_), .ZN(new_n1617_));
  NAND2_X1   g1354(.A1(new_n1616_), .A2(new_n1617_), .ZN(new_n1618_));
  OAI21_X1   g1355(.A1(new_n1615_), .A2(new_n1618_), .B(new_n308_), .ZN(new_n1619_));
  NAND2_X1   g1356(.A1(new_n1612_), .A2(new_n1619_), .ZN(new_n1620_));
  OAI21_X1   g1357(.A1(new_n1605_), .A2(new_n1620_), .B(\shift[6] ), .ZN(new_n1621_));
  NAND2_X1   g1358(.A1(new_n1593_), .A2(new_n1621_), .ZN(\result[10] ));
  OAI22_X1   g1359(.A1(new_n274_), .A2(new_n1106_), .B1(new_n1101_), .B2(new_n285_), .ZN(new_n1623_));
  OAI22_X1   g1360(.A1(new_n557_), .A2(new_n1142_), .B1(new_n1137_), .B2(new_n304_), .ZN(new_n1624_));
  NOR2_X1    g1361(.A1(new_n1623_), .A2(new_n1624_), .ZN(new_n1625_));
  OAI22_X1   g1362(.A1(new_n274_), .A2(new_n1083_), .B1(new_n1078_), .B2(new_n285_), .ZN(new_n1626_));
  OAI22_X1   g1363(.A1(new_n557_), .A2(new_n1095_), .B1(new_n1090_), .B2(new_n304_), .ZN(new_n1627_));
  OAI21_X1   g1364(.A1(new_n1626_), .A2(new_n1627_), .B(new_n340_), .ZN(new_n1628_));
  OAI21_X1   g1365(.A1(new_n537_), .A2(new_n1625_), .B(new_n1628_), .ZN(new_n1629_));
  OAI22_X1   g1366(.A1(new_n274_), .A2(new_n1238_), .B1(new_n1233_), .B2(new_n285_), .ZN(new_n1630_));
  OAI22_X1   g1367(.A1(new_n557_), .A2(new_n1119_), .B1(new_n1114_), .B2(new_n304_), .ZN(new_n1631_));
  OAI21_X1   g1368(.A1(new_n1630_), .A2(new_n1631_), .B(new_n373_), .ZN(new_n1632_));
  OAI22_X1   g1369(.A1(new_n274_), .A2(new_n1130_), .B1(new_n1125_), .B2(new_n285_), .ZN(new_n1633_));
  OAI22_X1   g1370(.A1(new_n557_), .A2(new_n1072_), .B1(new_n1067_), .B2(new_n304_), .ZN(new_n1634_));
  OAI21_X1   g1371(.A1(new_n1633_), .A2(new_n1634_), .B(new_n405_), .ZN(new_n1635_));
  NAND2_X1   g1372(.A1(new_n1632_), .A2(new_n1635_), .ZN(new_n1636_));
  OAI21_X1   g1373(.A1(new_n1629_), .A2(new_n1636_), .B(new_n264_), .ZN(new_n1637_));
  NOR3_X1    g1374(.A1(new_n777_), .A2(new_n275_), .A3(\shift[0] ), .ZN(new_n1638_));
  NOR3_X1    g1375(.A1(new_n719_), .A2(new_n266_), .A3(\shift[1] ), .ZN(new_n1639_));
  INV_X1     g1376(.I(new_n1186_), .ZN(new_n1640_));
  NOR3_X1    g1377(.A1(new_n723_), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1641_));
  NOR4_X1    g1378(.A1(new_n1638_), .A2(new_n1640_), .A3(new_n1639_), .A4(new_n1641_), .ZN(new_n1642_));
  OAI22_X1   g1379(.A1(new_n274_), .A2(new_n1179_), .B1(new_n1642_), .B2(new_n304_), .ZN(new_n1643_));
  OAI21_X1   g1380(.A1(new_n1194_), .A2(new_n1191_), .B(new_n294_), .ZN(new_n1644_));
  NAND3_X1   g1381(.A1(new_n266_), .A2(\a[53] ), .A3(\shift[1] ), .ZN(new_n1645_));
  NAND3_X1   g1382(.A1(new_n275_), .A2(\a[54] ), .A3(\shift[0] ), .ZN(new_n1646_));
  NAND2_X1   g1383(.A1(new_n1645_), .A2(new_n1646_), .ZN(new_n1647_));
  NAND2_X1   g1384(.A1(new_n266_), .A2(\a[55] ), .ZN(new_n1648_));
  OAI21_X1   g1385(.A1(new_n1648_), .A2(\shift[1] ), .B(new_n1171_), .ZN(new_n1649_));
  OAI21_X1   g1386(.A1(new_n1647_), .A2(new_n1649_), .B(new_n284_), .ZN(new_n1650_));
  NAND2_X1   g1387(.A1(new_n1650_), .A2(new_n1644_), .ZN(new_n1651_));
  OAI21_X1   g1388(.A1(new_n1643_), .A2(new_n1651_), .B(new_n405_), .ZN(new_n1652_));
  OAI22_X1   g1389(.A1(new_n274_), .A2(new_n1153_), .B1(new_n1148_), .B2(new_n285_), .ZN(new_n1653_));
  OAI22_X1   g1390(.A1(new_n557_), .A2(new_n1167_), .B1(new_n1162_), .B2(new_n304_), .ZN(new_n1654_));
  OAI21_X1   g1391(.A1(new_n1653_), .A2(new_n1654_), .B(new_n373_), .ZN(new_n1655_));
  NAND2_X1   g1392(.A1(new_n1655_), .A2(new_n1652_), .ZN(new_n1656_));
  OAI22_X1   g1393(.A1(new_n274_), .A2(new_n1214_), .B1(new_n1205_), .B2(new_n285_), .ZN(new_n1657_));
  OAI22_X1   g1394(.A1(new_n557_), .A2(new_n1252_), .B1(new_n1247_), .B2(new_n304_), .ZN(new_n1658_));
  OAI21_X1   g1395(.A1(new_n1657_), .A2(new_n1658_), .B(new_n340_), .ZN(new_n1659_));
  OAI22_X1   g1396(.A1(new_n274_), .A2(new_n1263_), .B1(new_n1258_), .B2(new_n285_), .ZN(new_n1660_));
  OAI22_X1   g1397(.A1(new_n557_), .A2(new_n1227_), .B1(new_n1222_), .B2(new_n304_), .ZN(new_n1661_));
  OAI21_X1   g1398(.A1(new_n1660_), .A2(new_n1661_), .B(new_n308_), .ZN(new_n1662_));
  NAND2_X1   g1399(.A1(new_n1659_), .A2(new_n1662_), .ZN(new_n1663_));
  OAI21_X1   g1400(.A1(new_n1663_), .A2(new_n1656_), .B(\shift[6] ), .ZN(new_n1664_));
  NAND2_X1   g1401(.A1(new_n1637_), .A2(new_n1664_), .ZN(\result[11] ));
  OAI21_X1   g1402(.A1(new_n319_), .A2(new_n322_), .B(new_n273_), .ZN(new_n1666_));
  OAI21_X1   g1403(.A1(new_n334_), .A2(new_n337_), .B(new_n284_), .ZN(new_n1667_));
  NAND2_X1   g1404(.A1(new_n1666_), .A2(new_n1667_), .ZN(new_n1668_));
  OAI21_X1   g1405(.A1(new_n271_), .A2(new_n268_), .B(new_n294_), .ZN(new_n1669_));
  OAI21_X1   g1406(.A1(new_n330_), .A2(new_n327_), .B(new_n303_), .ZN(new_n1670_));
  NAND2_X1   g1407(.A1(new_n1669_), .A2(new_n1670_), .ZN(new_n1671_));
  OAI21_X1   g1408(.A1(new_n1668_), .A2(new_n1671_), .B(new_n308_), .ZN(new_n1672_));
  OAI21_X1   g1409(.A1(new_n387_), .A2(new_n384_), .B(new_n273_), .ZN(new_n1673_));
  OAI21_X1   g1410(.A1(new_n402_), .A2(new_n399_), .B(new_n284_), .ZN(new_n1674_));
  NAND2_X1   g1411(.A1(new_n1673_), .A2(new_n1674_), .ZN(new_n1675_));
  OAI21_X1   g1412(.A1(new_n315_), .A2(new_n312_), .B(new_n294_), .ZN(new_n1676_));
  OAI21_X1   g1413(.A1(new_n395_), .A2(new_n392_), .B(new_n303_), .ZN(new_n1677_));
  NAND2_X1   g1414(.A1(new_n1676_), .A2(new_n1677_), .ZN(new_n1678_));
  OAI21_X1   g1415(.A1(new_n1675_), .A2(new_n1678_), .B(new_n340_), .ZN(new_n1679_));
  NAND2_X1   g1416(.A1(new_n1672_), .A2(new_n1679_), .ZN(new_n1680_));
  OAI21_X1   g1417(.A1(new_n421_), .A2(new_n418_), .B(new_n273_), .ZN(new_n1681_));
  OAI21_X1   g1418(.A1(new_n436_), .A2(new_n433_), .B(new_n284_), .ZN(new_n1682_));
  NAND2_X1   g1419(.A1(new_n1681_), .A2(new_n1682_), .ZN(new_n1683_));
  OAI21_X1   g1420(.A1(new_n345_), .A2(new_n348_), .B(new_n294_), .ZN(new_n1684_));
  OAI21_X1   g1421(.A1(new_n429_), .A2(new_n426_), .B(new_n303_), .ZN(new_n1685_));
  NAND2_X1   g1422(.A1(new_n1684_), .A2(new_n1685_), .ZN(new_n1686_));
  OAI21_X1   g1423(.A1(new_n1683_), .A2(new_n1686_), .B(new_n373_), .ZN(new_n1687_));
  OAI21_X1   g1424(.A1(new_n355_), .A2(new_n352_), .B(new_n273_), .ZN(new_n1688_));
  OAI21_X1   g1425(.A1(new_n370_), .A2(new_n367_), .B(new_n284_), .ZN(new_n1689_));
  NAND2_X1   g1426(.A1(new_n1688_), .A2(new_n1689_), .ZN(new_n1690_));
  OAI21_X1   g1427(.A1(new_n380_), .A2(new_n377_), .B(new_n294_), .ZN(new_n1691_));
  OAI21_X1   g1428(.A1(new_n363_), .A2(new_n360_), .B(new_n303_), .ZN(new_n1692_));
  NAND2_X1   g1429(.A1(new_n1691_), .A2(new_n1692_), .ZN(new_n1693_));
  OAI21_X1   g1430(.A1(new_n1690_), .A2(new_n1693_), .B(new_n405_), .ZN(new_n1694_));
  NAND2_X1   g1431(.A1(new_n1687_), .A2(new_n1694_), .ZN(new_n1695_));
  OAI21_X1   g1432(.A1(new_n1680_), .A2(new_n1695_), .B(new_n264_), .ZN(new_n1696_));
  OAI22_X1   g1433(.A1(new_n285_), .A2(new_n1493_), .B1(new_n485_), .B2(new_n274_), .ZN(new_n1697_));
  OAI21_X1   g1434(.A1(new_n505_), .A2(new_n508_), .B(new_n294_), .ZN(new_n1698_));
  OAI21_X1   g1435(.A1(new_n304_), .A2(new_n1492_), .B(new_n1698_), .ZN(new_n1699_));
  OAI21_X1   g1436(.A1(new_n1697_), .A2(new_n1699_), .B(new_n405_), .ZN(new_n1700_));
  OAI21_X1   g1437(.A1(new_n278_), .A2(new_n281_), .B(new_n273_), .ZN(new_n1701_));
  OAI21_X1   g1438(.A1(new_n285_), .A2(new_n302_), .B(new_n1701_), .ZN(new_n1702_));
  OAI21_X1   g1439(.A1(new_n474_), .A2(new_n477_), .B(new_n294_), .ZN(new_n1703_));
  OAI21_X1   g1440(.A1(new_n289_), .A2(new_n292_), .B(new_n303_), .ZN(new_n1704_));
  NAND2_X1   g1441(.A1(new_n1703_), .A2(new_n1704_), .ZN(new_n1705_));
  OAI21_X1   g1442(.A1(new_n1702_), .A2(new_n1705_), .B(new_n373_), .ZN(new_n1706_));
  NAND2_X1   g1443(.A1(new_n1700_), .A2(new_n1706_), .ZN(new_n1707_));
  NOR2_X1    g1444(.A1(new_n530_), .A2(new_n527_), .ZN(new_n1708_));
  OAI22_X1   g1445(.A1(new_n285_), .A2(new_n1708_), .B1(new_n1496_), .B2(new_n274_), .ZN(new_n1709_));
  OAI21_X1   g1446(.A1(new_n445_), .A2(new_n442_), .B(new_n294_), .ZN(new_n1710_));
  OAI21_X1   g1447(.A1(new_n523_), .A2(new_n520_), .B(new_n303_), .ZN(new_n1711_));
  NAND2_X1   g1448(.A1(new_n1710_), .A2(new_n1711_), .ZN(new_n1712_));
  OAI21_X1   g1449(.A1(new_n1709_), .A2(new_n1712_), .B(new_n340_), .ZN(new_n1713_));
  OAI21_X1   g1450(.A1(new_n449_), .A2(new_n452_), .B(new_n273_), .ZN(new_n1714_));
  OAI21_X1   g1451(.A1(new_n467_), .A2(new_n464_), .B(new_n284_), .ZN(new_n1715_));
  NAND2_X1   g1452(.A1(new_n1714_), .A2(new_n1715_), .ZN(new_n1716_));
  OAI21_X1   g1453(.A1(new_n414_), .A2(new_n411_), .B(new_n294_), .ZN(new_n1717_));
  OAI21_X1   g1454(.A1(new_n460_), .A2(new_n457_), .B(new_n303_), .ZN(new_n1718_));
  NAND2_X1   g1455(.A1(new_n1717_), .A2(new_n1718_), .ZN(new_n1719_));
  OAI21_X1   g1456(.A1(new_n1716_), .A2(new_n1719_), .B(new_n308_), .ZN(new_n1720_));
  NAND2_X1   g1457(.A1(new_n1713_), .A2(new_n1720_), .ZN(new_n1721_));
  OAI21_X1   g1458(.A1(new_n1707_), .A2(new_n1721_), .B(\shift[6] ), .ZN(new_n1722_));
  NAND2_X1   g1459(.A1(new_n1696_), .A2(new_n1722_), .ZN(\result[12] ));
  OAI22_X1   g1460(.A1(new_n274_), .A2(new_n595_), .B1(new_n614_), .B2(new_n285_), .ZN(new_n1724_));
  OAI22_X1   g1461(.A1(new_n557_), .A2(new_n546_), .B1(new_n605_), .B2(new_n304_), .ZN(new_n1725_));
  NOR2_X1    g1462(.A1(new_n1724_), .A2(new_n1725_), .ZN(new_n1726_));
  OAI22_X1   g1463(.A1(new_n274_), .A2(new_n674_), .B1(new_n693_), .B2(new_n285_), .ZN(new_n1727_));
  OAI22_X1   g1464(.A1(new_n557_), .A2(new_n586_), .B1(new_n684_), .B2(new_n304_), .ZN(new_n1728_));
  OAI21_X1   g1465(.A1(new_n1727_), .A2(new_n1728_), .B(new_n340_), .ZN(new_n1729_));
  OAI21_X1   g1466(.A1(new_n537_), .A2(new_n1726_), .B(new_n1729_), .ZN(new_n1730_));
  OAI22_X1   g1467(.A1(new_n274_), .A2(new_n754_), .B1(new_n773_), .B2(new_n285_), .ZN(new_n1731_));
  OAI22_X1   g1468(.A1(new_n557_), .A2(new_n626_), .B1(new_n764_), .B2(new_n304_), .ZN(new_n1732_));
  OAI21_X1   g1469(.A1(new_n1731_), .A2(new_n1732_), .B(new_n373_), .ZN(new_n1733_));
  OAI22_X1   g1470(.A1(new_n274_), .A2(new_n635_), .B1(new_n654_), .B2(new_n285_), .ZN(new_n1734_));
  OAI22_X1   g1471(.A1(new_n557_), .A2(new_n665_), .B1(new_n645_), .B2(new_n304_), .ZN(new_n1735_));
  OAI21_X1   g1472(.A1(new_n1734_), .A2(new_n1735_), .B(new_n405_), .ZN(new_n1736_));
  NAND2_X1   g1473(.A1(new_n1733_), .A2(new_n1736_), .ZN(new_n1737_));
  OAI21_X1   g1474(.A1(new_n1730_), .A2(new_n1737_), .B(new_n264_), .ZN(new_n1738_));
  OAI22_X1   g1475(.A1(new_n274_), .A2(new_n715_), .B1(new_n734_), .B2(new_n285_), .ZN(new_n1739_));
  OAI22_X1   g1476(.A1(new_n557_), .A2(new_n785_), .B1(new_n725_), .B2(new_n304_), .ZN(new_n1740_));
  OAI21_X1   g1477(.A1(new_n1739_), .A2(new_n1740_), .B(new_n405_), .ZN(new_n1741_));
  OAI22_X1   g1478(.A1(new_n274_), .A2(new_n555_), .B1(new_n575_), .B2(new_n285_), .ZN(new_n1742_));
  OAI22_X1   g1479(.A1(new_n557_), .A2(new_n706_), .B1(new_n566_), .B2(new_n304_), .ZN(new_n1743_));
  OAI21_X1   g1480(.A1(new_n1742_), .A2(new_n1743_), .B(new_n373_), .ZN(new_n1744_));
  NAND2_X1   g1481(.A1(new_n1741_), .A2(new_n1744_), .ZN(new_n1745_));
  OAI21_X1   g1482(.A1(new_n791_), .A2(new_n788_), .B(new_n273_), .ZN(new_n1746_));
  OAI21_X1   g1483(.A1(new_n803_), .A2(new_n806_), .B(new_n284_), .ZN(new_n1747_));
  NAND2_X1   g1484(.A1(new_n1746_), .A2(new_n1747_), .ZN(new_n1748_));
  OAI22_X1   g1485(.A1(new_n557_), .A2(new_n818_), .B1(new_n1357_), .B2(new_n304_), .ZN(new_n1749_));
  OAI21_X1   g1486(.A1(new_n1749_), .A2(new_n1748_), .B(new_n340_), .ZN(new_n1750_));
  OAI22_X1   g1487(.A1(new_n274_), .A2(new_n827_), .B1(new_n846_), .B2(new_n285_), .ZN(new_n1751_));
  OAI22_X1   g1488(.A1(new_n557_), .A2(new_n745_), .B1(new_n837_), .B2(new_n304_), .ZN(new_n1752_));
  OAI21_X1   g1489(.A1(new_n1751_), .A2(new_n1752_), .B(new_n308_), .ZN(new_n1753_));
  NAND2_X1   g1490(.A1(new_n1753_), .A2(new_n1750_), .ZN(new_n1754_));
  OAI21_X1   g1491(.A1(new_n1745_), .A2(new_n1754_), .B(\shift[6] ), .ZN(new_n1755_));
  NAND2_X1   g1492(.A1(new_n1738_), .A2(new_n1755_), .ZN(\result[13] ));
  OAI21_X1   g1493(.A1(new_n882_), .A2(new_n883_), .B(new_n273_), .ZN(new_n1757_));
  OAI21_X1   g1494(.A1(new_n891_), .A2(new_n894_), .B(new_n284_), .ZN(new_n1758_));
  NAND2_X1   g1495(.A1(new_n1757_), .A2(new_n1758_), .ZN(new_n1759_));
  OAI21_X1   g1496(.A1(new_n854_), .A2(new_n857_), .B(new_n294_), .ZN(new_n1760_));
  OAI21_X1   g1497(.A1(new_n886_), .A2(new_n889_), .B(new_n303_), .ZN(new_n1761_));
  NAND2_X1   g1498(.A1(new_n1760_), .A2(new_n1761_), .ZN(new_n1762_));
  OAI21_X1   g1499(.A1(new_n1759_), .A2(new_n1762_), .B(new_n308_), .ZN(new_n1763_));
  OAI21_X1   g1500(.A1(new_n937_), .A2(new_n940_), .B(new_n273_), .ZN(new_n1764_));
  OAI21_X1   g1501(.A1(new_n952_), .A2(new_n955_), .B(new_n284_), .ZN(new_n1765_));
  NAND2_X1   g1502(.A1(new_n1764_), .A2(new_n1765_), .ZN(new_n1766_));
  OAI21_X1   g1503(.A1(new_n875_), .A2(new_n878_), .B(new_n294_), .ZN(new_n1767_));
  OAI21_X1   g1504(.A1(new_n945_), .A2(new_n948_), .B(new_n303_), .ZN(new_n1768_));
  NAND2_X1   g1505(.A1(new_n1767_), .A2(new_n1768_), .ZN(new_n1769_));
  OAI21_X1   g1506(.A1(new_n1766_), .A2(new_n1769_), .B(new_n340_), .ZN(new_n1770_));
  NAND2_X1   g1507(.A1(new_n1763_), .A2(new_n1770_), .ZN(new_n1771_));
  OAI21_X1   g1508(.A1(new_n989_), .A2(new_n992_), .B(new_n273_), .ZN(new_n1772_));
  OAI21_X1   g1509(.A1(new_n1004_), .A2(new_n1007_), .B(new_n284_), .ZN(new_n1773_));
  NAND2_X1   g1510(.A1(new_n1772_), .A2(new_n1773_), .ZN(new_n1774_));
  OAI21_X1   g1511(.A1(new_n901_), .A2(new_n904_), .B(new_n294_), .ZN(new_n1775_));
  OAI21_X1   g1512(.A1(new_n997_), .A2(new_n1000_), .B(new_n303_), .ZN(new_n1776_));
  NAND2_X1   g1513(.A1(new_n1775_), .A2(new_n1776_), .ZN(new_n1777_));
  OAI21_X1   g1514(.A1(new_n1774_), .A2(new_n1777_), .B(new_n373_), .ZN(new_n1778_));
  OAI21_X1   g1515(.A1(new_n906_), .A2(new_n909_), .B(new_n273_), .ZN(new_n1779_));
  OAI21_X1   g1516(.A1(new_n921_), .A2(new_n924_), .B(new_n284_), .ZN(new_n1780_));
  NAND2_X1   g1517(.A1(new_n1779_), .A2(new_n1780_), .ZN(new_n1781_));
  OAI21_X1   g1518(.A1(new_n930_), .A2(new_n933_), .B(new_n294_), .ZN(new_n1782_));
  OAI21_X1   g1519(.A1(new_n914_), .A2(new_n917_), .B(new_n303_), .ZN(new_n1783_));
  NAND2_X1   g1520(.A1(new_n1782_), .A2(new_n1783_), .ZN(new_n1784_));
  OAI21_X1   g1521(.A1(new_n1781_), .A2(new_n1784_), .B(new_n405_), .ZN(new_n1785_));
  NAND2_X1   g1522(.A1(new_n1778_), .A2(new_n1785_), .ZN(new_n1786_));
  OAI21_X1   g1523(.A1(new_n1771_), .A2(new_n1786_), .B(new_n264_), .ZN(new_n1787_));
  OAI22_X1   g1524(.A1(new_n285_), .A2(new_n977_), .B1(new_n968_), .B2(new_n274_), .ZN(new_n1788_));
  OAI21_X1   g1525(.A1(new_n1012_), .A2(new_n1013_), .B(new_n294_), .ZN(new_n1789_));
  OAI21_X1   g1526(.A1(new_n304_), .A2(new_n1594_), .B(new_n1789_), .ZN(new_n1790_));
  OAI21_X1   g1527(.A1(new_n1788_), .A2(new_n1790_), .B(new_n405_), .ZN(new_n1791_));
  OAI21_X1   g1528(.A1(new_n861_), .A2(new_n862_), .B(new_n273_), .ZN(new_n1792_));
  OAI21_X1   g1529(.A1(new_n285_), .A2(new_n1598_), .B(new_n1792_), .ZN(new_n1793_));
  OAI21_X1   g1530(.A1(new_n961_), .A2(new_n962_), .B(new_n294_), .ZN(new_n1794_));
  OAI21_X1   g1531(.A1(new_n865_), .A2(new_n866_), .B(new_n303_), .ZN(new_n1795_));
  NAND2_X1   g1532(.A1(new_n1794_), .A2(new_n1795_), .ZN(new_n1796_));
  OAI21_X1   g1533(.A1(new_n1793_), .A2(new_n1796_), .B(new_n373_), .ZN(new_n1797_));
  NAND2_X1   g1534(.A1(new_n1791_), .A2(new_n1797_), .ZN(new_n1798_));
  OAI22_X1   g1535(.A1(new_n285_), .A2(new_n1606_), .B1(new_n1019_), .B2(new_n274_), .ZN(new_n1799_));
  OAI21_X1   g1536(.A1(new_n1036_), .A2(new_n1037_), .B(new_n294_), .ZN(new_n1800_));
  OAI21_X1   g1537(.A1(new_n1023_), .A2(new_n1024_), .B(new_n303_), .ZN(new_n1801_));
  NAND2_X1   g1538(.A1(new_n1800_), .A2(new_n1801_), .ZN(new_n1802_));
  OAI21_X1   g1539(.A1(new_n1799_), .A2(new_n1802_), .B(new_n340_), .ZN(new_n1803_));
  OAI21_X1   g1540(.A1(new_n1041_), .A2(new_n1042_), .B(new_n273_), .ZN(new_n1804_));
  OAI21_X1   g1541(.A1(new_n1052_), .A2(new_n1055_), .B(new_n284_), .ZN(new_n1805_));
  NAND2_X1   g1542(.A1(new_n1804_), .A2(new_n1805_), .ZN(new_n1806_));
  OAI21_X1   g1543(.A1(new_n982_), .A2(new_n985_), .B(new_n294_), .ZN(new_n1807_));
  OAI21_X1   g1544(.A1(new_n1047_), .A2(new_n1050_), .B(new_n303_), .ZN(new_n1808_));
  NAND2_X1   g1545(.A1(new_n1807_), .A2(new_n1808_), .ZN(new_n1809_));
  OAI21_X1   g1546(.A1(new_n1806_), .A2(new_n1809_), .B(new_n308_), .ZN(new_n1810_));
  NAND2_X1   g1547(.A1(new_n1803_), .A2(new_n1810_), .ZN(new_n1811_));
  OAI21_X1   g1548(.A1(new_n1798_), .A2(new_n1811_), .B(\shift[6] ), .ZN(new_n1812_));
  NAND2_X1   g1549(.A1(new_n1787_), .A2(new_n1812_), .ZN(\result[14] ));
  OAI22_X1   g1550(.A1(new_n274_), .A2(new_n1095_), .B1(new_n1106_), .B2(new_n285_), .ZN(new_n1814_));
  OAI22_X1   g1551(.A1(new_n557_), .A2(new_n1137_), .B1(new_n1101_), .B2(new_n304_), .ZN(new_n1815_));
  OAI21_X1   g1552(.A1(new_n1814_), .A2(new_n1815_), .B(new_n308_), .ZN(new_n1816_));
  OAI22_X1   g1553(.A1(new_n274_), .A2(new_n1072_), .B1(new_n1083_), .B2(new_n285_), .ZN(new_n1817_));
  OAI22_X1   g1554(.A1(new_n557_), .A2(new_n1090_), .B1(new_n1078_), .B2(new_n304_), .ZN(new_n1818_));
  OAI21_X1   g1555(.A1(new_n1817_), .A2(new_n1818_), .B(new_n340_), .ZN(new_n1819_));
  NAND2_X1   g1556(.A1(new_n1816_), .A2(new_n1819_), .ZN(new_n1820_));
  OAI22_X1   g1557(.A1(new_n274_), .A2(new_n1227_), .B1(new_n1238_), .B2(new_n285_), .ZN(new_n1821_));
  OAI22_X1   g1558(.A1(new_n557_), .A2(new_n1114_), .B1(new_n1233_), .B2(new_n304_), .ZN(new_n1822_));
  OAI21_X1   g1559(.A1(new_n1821_), .A2(new_n1822_), .B(new_n373_), .ZN(new_n1823_));
  OAI22_X1   g1560(.A1(new_n274_), .A2(new_n1119_), .B1(new_n1130_), .B2(new_n285_), .ZN(new_n1824_));
  OAI22_X1   g1561(.A1(new_n557_), .A2(new_n1067_), .B1(new_n1125_), .B2(new_n304_), .ZN(new_n1825_));
  OAI21_X1   g1562(.A1(new_n1824_), .A2(new_n1825_), .B(new_n405_), .ZN(new_n1826_));
  NAND2_X1   g1563(.A1(new_n1823_), .A2(new_n1826_), .ZN(new_n1827_));
  OAI21_X1   g1564(.A1(new_n1820_), .A2(new_n1827_), .B(new_n264_), .ZN(new_n1828_));
  OAI22_X1   g1565(.A1(new_n274_), .A2(new_n1167_), .B1(new_n1179_), .B2(new_n285_), .ZN(new_n1829_));
  OAI22_X1   g1566(.A1(new_n557_), .A2(new_n1642_), .B1(new_n1174_), .B2(new_n304_), .ZN(new_n1830_));
  OAI21_X1   g1567(.A1(new_n1829_), .A2(new_n1830_), .B(new_n405_), .ZN(new_n1831_));
  OAI22_X1   g1568(.A1(new_n274_), .A2(new_n1142_), .B1(new_n1153_), .B2(new_n285_), .ZN(new_n1832_));
  OAI22_X1   g1569(.A1(new_n557_), .A2(new_n1162_), .B1(new_n1148_), .B2(new_n304_), .ZN(new_n1833_));
  OAI21_X1   g1570(.A1(new_n1832_), .A2(new_n1833_), .B(new_n373_), .ZN(new_n1834_));
  NAND2_X1   g1571(.A1(new_n1831_), .A2(new_n1834_), .ZN(new_n1835_));
  OAI21_X1   g1572(.A1(new_n1194_), .A2(new_n1191_), .B(new_n273_), .ZN(new_n1836_));
  NAND3_X1   g1573(.A1(new_n266_), .A2(\a[41] ), .A3(\shift[1] ), .ZN(new_n1837_));
  NAND3_X1   g1574(.A1(new_n275_), .A2(\a[42] ), .A3(\shift[0] ), .ZN(new_n1838_));
  NAND2_X1   g1575(.A1(new_n1837_), .A2(new_n1838_), .ZN(new_n1839_));
  NAND2_X1   g1576(.A1(new_n266_), .A2(\a[43] ), .ZN(new_n1840_));
  OAI21_X1   g1577(.A1(new_n1840_), .A2(\shift[1] ), .B(new_n1210_), .ZN(new_n1841_));
  OAI21_X1   g1578(.A1(new_n1839_), .A2(new_n1841_), .B(new_n284_), .ZN(new_n1842_));
  NAND2_X1   g1579(.A1(new_n1842_), .A2(new_n1836_), .ZN(new_n1843_));
  OAI22_X1   g1580(.A1(new_n557_), .A2(new_n1247_), .B1(new_n1205_), .B2(new_n304_), .ZN(new_n1844_));
  OAI21_X1   g1581(.A1(new_n1844_), .A2(new_n1843_), .B(new_n340_), .ZN(new_n1845_));
  OAI22_X1   g1582(.A1(new_n274_), .A2(new_n1252_), .B1(new_n1263_), .B2(new_n285_), .ZN(new_n1846_));
  OAI22_X1   g1583(.A1(new_n557_), .A2(new_n1222_), .B1(new_n1258_), .B2(new_n304_), .ZN(new_n1847_));
  OAI21_X1   g1584(.A1(new_n1846_), .A2(new_n1847_), .B(new_n308_), .ZN(new_n1848_));
  NAND2_X1   g1585(.A1(new_n1848_), .A2(new_n1845_), .ZN(new_n1849_));
  OAI21_X1   g1586(.A1(new_n1835_), .A2(new_n1849_), .B(\shift[6] ), .ZN(new_n1850_));
  NAND2_X1   g1587(.A1(new_n1828_), .A2(new_n1850_), .ZN(\result[15] ));
  OAI21_X1   g1588(.A1(new_n324_), .A2(new_n339_), .B(new_n308_), .ZN(new_n1852_));
  OAI21_X1   g1589(.A1(new_n389_), .A2(new_n404_), .B(new_n340_), .ZN(new_n1853_));
  NAND2_X1   g1590(.A1(new_n1852_), .A2(new_n1853_), .ZN(new_n1854_));
  OAI21_X1   g1591(.A1(new_n423_), .A2(new_n438_), .B(new_n373_), .ZN(new_n1855_));
  OAI21_X1   g1592(.A1(new_n357_), .A2(new_n372_), .B(new_n405_), .ZN(new_n1856_));
  NAND2_X1   g1593(.A1(new_n1855_), .A2(new_n1856_), .ZN(new_n1857_));
  OAI21_X1   g1594(.A1(new_n1854_), .A2(new_n1857_), .B(new_n264_), .ZN(new_n1858_));
  OAI21_X1   g1595(.A1(new_n286_), .A2(new_n305_), .B(new_n373_), .ZN(new_n1859_));
  OAI21_X1   g1596(.A1(new_n454_), .A2(new_n469_), .B(new_n308_), .ZN(new_n1860_));
  NAND2_X1   g1597(.A1(new_n1859_), .A2(new_n1860_), .ZN(new_n1861_));
  OAI21_X1   g1598(.A1(new_n486_), .A2(new_n501_), .B(new_n405_), .ZN(new_n1862_));
  OAI21_X1   g1599(.A1(new_n517_), .A2(new_n532_), .B(new_n340_), .ZN(new_n1863_));
  NAND2_X1   g1600(.A1(new_n1862_), .A2(new_n1863_), .ZN(new_n1864_));
  OAI21_X1   g1601(.A1(new_n1861_), .A2(new_n1864_), .B(\shift[6] ), .ZN(new_n1865_));
  NAND2_X1   g1602(.A1(new_n1858_), .A2(new_n1865_), .ZN(\result[16] ));
  NOR2_X1    g1603(.A1(new_n675_), .A2(new_n694_), .ZN(new_n1867_));
  OAI21_X1   g1604(.A1(new_n596_), .A2(new_n615_), .B(new_n308_), .ZN(new_n1868_));
  OAI21_X1   g1605(.A1(new_n1062_), .A2(new_n1867_), .B(new_n1868_), .ZN(new_n1869_));
  OAI21_X1   g1606(.A1(new_n755_), .A2(new_n774_), .B(new_n373_), .ZN(new_n1870_));
  OAI21_X1   g1607(.A1(new_n636_), .A2(new_n655_), .B(new_n405_), .ZN(new_n1871_));
  NAND2_X1   g1608(.A1(new_n1870_), .A2(new_n1871_), .ZN(new_n1872_));
  OAI21_X1   g1609(.A1(new_n1869_), .A2(new_n1872_), .B(new_n264_), .ZN(new_n1873_));
  OAI21_X1   g1610(.A1(new_n716_), .A2(new_n735_), .B(new_n405_), .ZN(new_n1874_));
  OAI21_X1   g1611(.A1(new_n556_), .A2(new_n576_), .B(new_n373_), .ZN(new_n1875_));
  NAND2_X1   g1612(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1876_));
  OAI21_X1   g1613(.A1(new_n793_), .A2(new_n808_), .B(new_n340_), .ZN(new_n1877_));
  OAI21_X1   g1614(.A1(new_n828_), .A2(new_n847_), .B(new_n308_), .ZN(new_n1878_));
  NAND2_X1   g1615(.A1(new_n1878_), .A2(new_n1877_), .ZN(new_n1879_));
  OAI21_X1   g1616(.A1(new_n1876_), .A2(new_n1879_), .B(\shift[6] ), .ZN(new_n1880_));
  NAND2_X1   g1617(.A1(new_n1873_), .A2(new_n1880_), .ZN(\result[17] ));
  OAI21_X1   g1618(.A1(new_n885_), .A2(new_n896_), .B(new_n308_), .ZN(new_n1882_));
  OAI21_X1   g1619(.A1(new_n942_), .A2(new_n957_), .B(new_n340_), .ZN(new_n1883_));
  NAND2_X1   g1620(.A1(new_n1882_), .A2(new_n1883_), .ZN(new_n1884_));
  OAI21_X1   g1621(.A1(new_n994_), .A2(new_n1009_), .B(new_n373_), .ZN(new_n1885_));
  OAI21_X1   g1622(.A1(new_n911_), .A2(new_n926_), .B(new_n405_), .ZN(new_n1886_));
  NAND2_X1   g1623(.A1(new_n1885_), .A2(new_n1886_), .ZN(new_n1887_));
  OAI21_X1   g1624(.A1(new_n1884_), .A2(new_n1887_), .B(new_n264_), .ZN(new_n1888_));
  OAI21_X1   g1625(.A1(new_n969_), .A2(new_n978_), .B(new_n405_), .ZN(new_n1889_));
  OAI21_X1   g1626(.A1(new_n864_), .A2(new_n871_), .B(new_n373_), .ZN(new_n1890_));
  NAND2_X1   g1627(.A1(new_n1889_), .A2(new_n1890_), .ZN(new_n1891_));
  OAI21_X1   g1628(.A1(new_n1020_), .A2(new_n1032_), .B(new_n340_), .ZN(new_n1892_));
  OAI21_X1   g1629(.A1(new_n1044_), .A2(new_n1057_), .B(new_n308_), .ZN(new_n1893_));
  NAND2_X1   g1630(.A1(new_n1892_), .A2(new_n1893_), .ZN(new_n1894_));
  OAI21_X1   g1631(.A1(new_n1891_), .A2(new_n1894_), .B(\shift[6] ), .ZN(new_n1895_));
  NAND2_X1   g1632(.A1(new_n1888_), .A2(new_n1895_), .ZN(\result[18] ));
  OAI21_X1   g1633(.A1(new_n1073_), .A2(new_n1084_), .B(new_n340_), .ZN(new_n1897_));
  OAI21_X1   g1634(.A1(new_n537_), .A2(new_n1108_), .B(new_n1897_), .ZN(new_n1898_));
  OAI21_X1   g1635(.A1(new_n1120_), .A2(new_n1131_), .B(new_n405_), .ZN(new_n1899_));
  OAI21_X1   g1636(.A1(new_n1228_), .A2(new_n1239_), .B(new_n373_), .ZN(new_n1900_));
  NAND2_X1   g1637(.A1(new_n1899_), .A2(new_n1900_), .ZN(new_n1901_));
  OAI21_X1   g1638(.A1(new_n1898_), .A2(new_n1901_), .B(new_n264_), .ZN(new_n1902_));
  OAI21_X1   g1639(.A1(new_n1168_), .A2(new_n1180_), .B(new_n405_), .ZN(new_n1903_));
  OAI21_X1   g1640(.A1(new_n1143_), .A2(new_n1154_), .B(new_n373_), .ZN(new_n1904_));
  NAND2_X1   g1641(.A1(new_n1903_), .A2(new_n1904_), .ZN(new_n1905_));
  OAI21_X1   g1642(.A1(new_n1253_), .A2(new_n1264_), .B(new_n308_), .ZN(new_n1906_));
  OAI21_X1   g1643(.A1(new_n1215_), .A2(new_n1196_), .B(new_n340_), .ZN(new_n1907_));
  NAND2_X1   g1644(.A1(new_n1906_), .A2(new_n1907_), .ZN(new_n1908_));
  OAI21_X1   g1645(.A1(new_n1905_), .A2(new_n1908_), .B(\shift[6] ), .ZN(new_n1909_));
  NAND2_X1   g1646(.A1(new_n1902_), .A2(new_n1909_), .ZN(\result[19] ));
  OAI21_X1   g1647(.A1(new_n1275_), .A2(new_n1278_), .B(new_n308_), .ZN(new_n1911_));
  OAI21_X1   g1648(.A1(new_n1290_), .A2(new_n1293_), .B(new_n340_), .ZN(new_n1912_));
  NAND2_X1   g1649(.A1(new_n1911_), .A2(new_n1912_), .ZN(new_n1913_));
  OAI21_X1   g1650(.A1(new_n1321_), .A2(new_n1324_), .B(new_n373_), .ZN(new_n1914_));
  OAI21_X1   g1651(.A1(new_n1283_), .A2(new_n1286_), .B(new_n405_), .ZN(new_n1915_));
  NAND2_X1   g1652(.A1(new_n1914_), .A2(new_n1915_), .ZN(new_n1916_));
  OAI21_X1   g1653(.A1(new_n1913_), .A2(new_n1916_), .B(new_n264_), .ZN(new_n1917_));
  OAI21_X1   g1654(.A1(new_n1270_), .A2(new_n1272_), .B(new_n373_), .ZN(new_n1918_));
  OAI21_X1   g1655(.A1(new_n1299_), .A2(new_n1302_), .B(new_n340_), .ZN(new_n1919_));
  NAND2_X1   g1656(.A1(new_n1918_), .A2(new_n1919_), .ZN(new_n1920_));
  OAI21_X1   g1657(.A1(new_n1314_), .A2(new_n1317_), .B(new_n308_), .ZN(new_n1921_));
  OAI21_X1   g1658(.A1(new_n1306_), .A2(new_n1309_), .B(new_n405_), .ZN(new_n1922_));
  NAND2_X1   g1659(.A1(new_n1921_), .A2(new_n1922_), .ZN(new_n1923_));
  OAI21_X1   g1660(.A1(new_n1920_), .A2(new_n1923_), .B(\shift[6] ), .ZN(new_n1924_));
  NAND2_X1   g1661(.A1(new_n1917_), .A2(new_n1924_), .ZN(\result[20] ));
  OAI21_X1   g1662(.A1(new_n1332_), .A2(new_n1333_), .B(new_n308_), .ZN(new_n1926_));
  OAI21_X1   g1663(.A1(new_n1339_), .A2(new_n1340_), .B(new_n340_), .ZN(new_n1927_));
  NAND2_X1   g1664(.A1(new_n1926_), .A2(new_n1927_), .ZN(new_n1928_));
  OAI21_X1   g1665(.A1(new_n1361_), .A2(new_n1362_), .B(new_n373_), .ZN(new_n1929_));
  OAI21_X1   g1666(.A1(new_n1336_), .A2(new_n1337_), .B(new_n405_), .ZN(new_n1930_));
  NAND2_X1   g1667(.A1(new_n1929_), .A2(new_n1930_), .ZN(new_n1931_));
  OAI21_X1   g1668(.A1(new_n1928_), .A2(new_n1931_), .B(new_n264_), .ZN(new_n1932_));
  OAI21_X1   g1669(.A1(new_n1329_), .A2(new_n1330_), .B(new_n373_), .ZN(new_n1933_));
  OAI21_X1   g1670(.A1(new_n1344_), .A2(new_n1347_), .B(new_n340_), .ZN(new_n1934_));
  NAND2_X1   g1671(.A1(new_n1933_), .A2(new_n1934_), .ZN(new_n1935_));
  OAI21_X1   g1672(.A1(new_n1358_), .A2(new_n1359_), .B(new_n308_), .ZN(new_n1936_));
  OAI21_X1   g1673(.A1(new_n1349_), .A2(new_n1350_), .B(new_n405_), .ZN(new_n1937_));
  NAND2_X1   g1674(.A1(new_n1936_), .A2(new_n1937_), .ZN(new_n1938_));
  OAI21_X1   g1675(.A1(new_n1938_), .A2(new_n1935_), .B(\shift[6] ), .ZN(new_n1939_));
  NAND2_X1   g1676(.A1(new_n1932_), .A2(new_n1939_), .ZN(\result[21] ));
  OAI21_X1   g1677(.A1(new_n1374_), .A2(new_n1377_), .B(new_n308_), .ZN(new_n1941_));
  OAI21_X1   g1678(.A1(new_n1389_), .A2(new_n1392_), .B(new_n340_), .ZN(new_n1942_));
  NAND2_X1   g1679(.A1(new_n1941_), .A2(new_n1942_), .ZN(new_n1943_));
  OAI21_X1   g1680(.A1(new_n1420_), .A2(new_n1423_), .B(new_n373_), .ZN(new_n1944_));
  OAI21_X1   g1681(.A1(new_n1382_), .A2(new_n1385_), .B(new_n405_), .ZN(new_n1945_));
  NAND2_X1   g1682(.A1(new_n1944_), .A2(new_n1945_), .ZN(new_n1946_));
  OAI21_X1   g1683(.A1(new_n1943_), .A2(new_n1946_), .B(new_n264_), .ZN(new_n1947_));
  OAI21_X1   g1684(.A1(new_n1368_), .A2(new_n1370_), .B(new_n373_), .ZN(new_n1948_));
  OAI21_X1   g1685(.A1(new_n1398_), .A2(new_n1401_), .B(new_n340_), .ZN(new_n1949_));
  NAND2_X1   g1686(.A1(new_n1948_), .A2(new_n1949_), .ZN(new_n1950_));
  OAI21_X1   g1687(.A1(new_n1413_), .A2(new_n1416_), .B(new_n308_), .ZN(new_n1951_));
  OAI21_X1   g1688(.A1(new_n1405_), .A2(new_n1408_), .B(new_n405_), .ZN(new_n1952_));
  NAND2_X1   g1689(.A1(new_n1951_), .A2(new_n1952_), .ZN(new_n1953_));
  OAI21_X1   g1690(.A1(new_n1950_), .A2(new_n1953_), .B(\shift[6] ), .ZN(new_n1954_));
  NAND2_X1   g1691(.A1(new_n1947_), .A2(new_n1954_), .ZN(\result[22] ));
  OAI21_X1   g1692(.A1(new_n1431_), .A2(new_n1432_), .B(new_n308_), .ZN(new_n1956_));
  OAI21_X1   g1693(.A1(new_n1455_), .A2(new_n1456_), .B(new_n373_), .ZN(new_n1957_));
  NAND2_X1   g1694(.A1(new_n1956_), .A2(new_n1957_), .ZN(new_n1958_));
  OAI21_X1   g1695(.A1(new_n1435_), .A2(new_n1436_), .B(new_n405_), .ZN(new_n1959_));
  OAI21_X1   g1696(.A1(new_n1438_), .A2(new_n1439_), .B(new_n340_), .ZN(new_n1960_));
  NAND2_X1   g1697(.A1(new_n1959_), .A2(new_n1960_), .ZN(new_n1961_));
  OAI21_X1   g1698(.A1(new_n1958_), .A2(new_n1961_), .B(new_n264_), .ZN(new_n1962_));
  OAI21_X1   g1699(.A1(new_n1446_), .A2(new_n1445_), .B(new_n340_), .ZN(new_n1963_));
  OAI21_X1   g1700(.A1(new_n1448_), .A2(new_n1449_), .B(new_n405_), .ZN(new_n1964_));
  NAND2_X1   g1701(.A1(new_n1964_), .A2(new_n1963_), .ZN(new_n1965_));
  OAI21_X1   g1702(.A1(new_n1452_), .A2(new_n1453_), .B(new_n308_), .ZN(new_n1966_));
  OAI21_X1   g1703(.A1(new_n1428_), .A2(new_n1429_), .B(new_n373_), .ZN(new_n1967_));
  NAND2_X1   g1704(.A1(new_n1966_), .A2(new_n1967_), .ZN(new_n1968_));
  OAI21_X1   g1705(.A1(new_n1968_), .A2(new_n1965_), .B(\shift[6] ), .ZN(new_n1969_));
  NAND2_X1   g1706(.A1(new_n1962_), .A2(new_n1969_), .ZN(\result[23] ));
  OAI21_X1   g1707(.A1(new_n1470_), .A2(new_n1473_), .B(new_n308_), .ZN(new_n1971_));
  OAI21_X1   g1708(.A1(new_n1515_), .A2(new_n1518_), .B(new_n373_), .ZN(new_n1972_));
  NAND2_X1   g1709(.A1(new_n1971_), .A2(new_n1972_), .ZN(new_n1973_));
  OAI21_X1   g1710(.A1(new_n1478_), .A2(new_n1481_), .B(new_n405_), .ZN(new_n1974_));
  OAI21_X1   g1711(.A1(new_n1485_), .A2(new_n1488_), .B(new_n340_), .ZN(new_n1975_));
  NAND2_X1   g1712(.A1(new_n1974_), .A2(new_n1975_), .ZN(new_n1976_));
  OAI21_X1   g1713(.A1(new_n1973_), .A2(new_n1976_), .B(new_n264_), .ZN(new_n1977_));
  OAI21_X1   g1714(.A1(new_n1494_), .A2(new_n1497_), .B(new_n340_), .ZN(new_n1978_));
  OAI21_X1   g1715(.A1(new_n1500_), .A2(new_n1503_), .B(new_n405_), .ZN(new_n1979_));
  NAND2_X1   g1716(.A1(new_n1978_), .A2(new_n1979_), .ZN(new_n1980_));
  OAI21_X1   g1717(.A1(new_n1508_), .A2(new_n1511_), .B(new_n308_), .ZN(new_n1981_));
  OAI21_X1   g1718(.A1(new_n1463_), .A2(new_n1466_), .B(new_n373_), .ZN(new_n1982_));
  NAND2_X1   g1719(.A1(new_n1981_), .A2(new_n1982_), .ZN(new_n1983_));
  OAI21_X1   g1720(.A1(new_n1980_), .A2(new_n1983_), .B(\shift[6] ), .ZN(new_n1984_));
  NAND2_X1   g1721(.A1(new_n1977_), .A2(new_n1984_), .ZN(\result[24] ));
  OAI21_X1   g1722(.A1(new_n1526_), .A2(new_n1527_), .B(new_n308_), .ZN(new_n1986_));
  OAI21_X1   g1723(.A1(new_n1557_), .A2(new_n1558_), .B(new_n373_), .ZN(new_n1987_));
  NAND2_X1   g1724(.A1(new_n1986_), .A2(new_n1987_), .ZN(new_n1988_));
  OAI21_X1   g1725(.A1(new_n1530_), .A2(new_n1531_), .B(new_n405_), .ZN(new_n1989_));
  OAI21_X1   g1726(.A1(new_n1533_), .A2(new_n1534_), .B(new_n340_), .ZN(new_n1990_));
  NAND2_X1   g1727(.A1(new_n1989_), .A2(new_n1990_), .ZN(new_n1991_));
  OAI21_X1   g1728(.A1(new_n1988_), .A2(new_n1991_), .B(new_n264_), .ZN(new_n1992_));
  OAI21_X1   g1729(.A1(new_n1538_), .A2(new_n1546_), .B(new_n340_), .ZN(new_n1993_));
  OAI21_X1   g1730(.A1(new_n1548_), .A2(new_n1549_), .B(new_n405_), .ZN(new_n1994_));
  NAND2_X1   g1731(.A1(new_n1994_), .A2(new_n1993_), .ZN(new_n1995_));
  OAI21_X1   g1732(.A1(new_n1555_), .A2(new_n1554_), .B(new_n308_), .ZN(new_n1996_));
  OAI21_X1   g1733(.A1(new_n1523_), .A2(new_n1524_), .B(new_n373_), .ZN(new_n1997_));
  NAND2_X1   g1734(.A1(new_n1997_), .A2(new_n1996_), .ZN(new_n1998_));
  OAI21_X1   g1735(.A1(new_n1995_), .A2(new_n1998_), .B(\shift[6] ), .ZN(new_n1999_));
  NAND2_X1   g1736(.A1(new_n1992_), .A2(new_n1999_), .ZN(\result[25] ));
  OAI21_X1   g1737(.A1(new_n1572_), .A2(new_n1575_), .B(new_n308_), .ZN(new_n2001_));
  OAI21_X1   g1738(.A1(new_n1587_), .A2(new_n1590_), .B(new_n340_), .ZN(new_n2002_));
  NAND2_X1   g1739(.A1(new_n2001_), .A2(new_n2002_), .ZN(new_n2003_));
  OAI21_X1   g1740(.A1(new_n1615_), .A2(new_n1618_), .B(new_n373_), .ZN(new_n2004_));
  OAI21_X1   g1741(.A1(new_n1580_), .A2(new_n1583_), .B(new_n405_), .ZN(new_n2005_));
  NAND2_X1   g1742(.A1(new_n2004_), .A2(new_n2005_), .ZN(new_n2006_));
  OAI21_X1   g1743(.A1(new_n2003_), .A2(new_n2006_), .B(new_n264_), .ZN(new_n2007_));
  OAI21_X1   g1744(.A1(new_n1595_), .A2(new_n1596_), .B(new_n340_), .ZN(new_n2008_));
  OAI21_X1   g1745(.A1(new_n1600_), .A2(new_n1603_), .B(new_n405_), .ZN(new_n2009_));
  NAND2_X1   g1746(.A1(new_n2008_), .A2(new_n2009_), .ZN(new_n2010_));
  OAI21_X1   g1747(.A1(new_n1608_), .A2(new_n1611_), .B(new_n308_), .ZN(new_n2011_));
  OAI21_X1   g1748(.A1(new_n1565_), .A2(new_n1568_), .B(new_n373_), .ZN(new_n2012_));
  NAND2_X1   g1749(.A1(new_n2011_), .A2(new_n2012_), .ZN(new_n2013_));
  OAI21_X1   g1750(.A1(new_n2010_), .A2(new_n2013_), .B(\shift[6] ), .ZN(new_n2014_));
  NAND2_X1   g1751(.A1(new_n2007_), .A2(new_n2014_), .ZN(\result[26] ));
  OAI21_X1   g1752(.A1(new_n1626_), .A2(new_n1627_), .B(new_n308_), .ZN(new_n2016_));
  OAI21_X1   g1753(.A1(new_n1633_), .A2(new_n1634_), .B(new_n340_), .ZN(new_n2017_));
  NAND2_X1   g1754(.A1(new_n2016_), .A2(new_n2017_), .ZN(new_n2018_));
  OAI21_X1   g1755(.A1(new_n1660_), .A2(new_n1661_), .B(new_n373_), .ZN(new_n2019_));
  OAI21_X1   g1756(.A1(new_n1630_), .A2(new_n1631_), .B(new_n405_), .ZN(new_n2020_));
  NAND2_X1   g1757(.A1(new_n2019_), .A2(new_n2020_), .ZN(new_n2021_));
  OAI21_X1   g1758(.A1(new_n2018_), .A2(new_n2021_), .B(new_n264_), .ZN(new_n2022_));
  OAI21_X1   g1759(.A1(new_n1643_), .A2(new_n1651_), .B(new_n340_), .ZN(new_n2023_));
  OAI21_X1   g1760(.A1(new_n1653_), .A2(new_n1654_), .B(new_n405_), .ZN(new_n2024_));
  NAND2_X1   g1761(.A1(new_n2024_), .A2(new_n2023_), .ZN(new_n2025_));
  OAI21_X1   g1762(.A1(new_n1657_), .A2(new_n1658_), .B(new_n308_), .ZN(new_n2026_));
  OAI21_X1   g1763(.A1(new_n1623_), .A2(new_n1624_), .B(new_n373_), .ZN(new_n2027_));
  NAND2_X1   g1764(.A1(new_n2026_), .A2(new_n2027_), .ZN(new_n2028_));
  OAI21_X1   g1765(.A1(new_n2028_), .A2(new_n2025_), .B(\shift[6] ), .ZN(new_n2029_));
  NAND2_X1   g1766(.A1(new_n2022_), .A2(new_n2029_), .ZN(\result[27] ));
  OAI21_X1   g1767(.A1(new_n1675_), .A2(new_n1678_), .B(new_n308_), .ZN(new_n2031_));
  OAI21_X1   g1768(.A1(new_n1690_), .A2(new_n1693_), .B(new_n340_), .ZN(new_n2032_));
  NAND2_X1   g1769(.A1(new_n2031_), .A2(new_n2032_), .ZN(new_n2033_));
  OAI21_X1   g1770(.A1(new_n1716_), .A2(new_n1719_), .B(new_n373_), .ZN(new_n2034_));
  OAI21_X1   g1771(.A1(new_n1683_), .A2(new_n1686_), .B(new_n405_), .ZN(new_n2035_));
  NAND2_X1   g1772(.A1(new_n2034_), .A2(new_n2035_), .ZN(new_n2036_));
  OAI21_X1   g1773(.A1(new_n2033_), .A2(new_n2036_), .B(new_n264_), .ZN(new_n2037_));
  OAI21_X1   g1774(.A1(new_n1697_), .A2(new_n1699_), .B(new_n340_), .ZN(new_n2038_));
  OAI21_X1   g1775(.A1(new_n1702_), .A2(new_n1705_), .B(new_n405_), .ZN(new_n2039_));
  NAND2_X1   g1776(.A1(new_n2038_), .A2(new_n2039_), .ZN(new_n2040_));
  OAI21_X1   g1777(.A1(new_n1709_), .A2(new_n1712_), .B(new_n308_), .ZN(new_n2041_));
  OAI21_X1   g1778(.A1(new_n1668_), .A2(new_n1671_), .B(new_n373_), .ZN(new_n2042_));
  NAND2_X1   g1779(.A1(new_n2041_), .A2(new_n2042_), .ZN(new_n2043_));
  OAI21_X1   g1780(.A1(new_n2040_), .A2(new_n2043_), .B(\shift[6] ), .ZN(new_n2044_));
  NAND2_X1   g1781(.A1(new_n2037_), .A2(new_n2044_), .ZN(\result[28] ));
  OAI21_X1   g1782(.A1(new_n1727_), .A2(new_n1728_), .B(new_n308_), .ZN(new_n2046_));
  OAI21_X1   g1783(.A1(new_n1734_), .A2(new_n1735_), .B(new_n340_), .ZN(new_n2047_));
  NAND2_X1   g1784(.A1(new_n2046_), .A2(new_n2047_), .ZN(new_n2048_));
  OAI21_X1   g1785(.A1(new_n1751_), .A2(new_n1752_), .B(new_n373_), .ZN(new_n2049_));
  OAI21_X1   g1786(.A1(new_n1731_), .A2(new_n1732_), .B(new_n405_), .ZN(new_n2050_));
  NAND2_X1   g1787(.A1(new_n2049_), .A2(new_n2050_), .ZN(new_n2051_));
  OAI21_X1   g1788(.A1(new_n2048_), .A2(new_n2051_), .B(new_n264_), .ZN(new_n2052_));
  OAI21_X1   g1789(.A1(new_n1739_), .A2(new_n1740_), .B(new_n340_), .ZN(new_n2053_));
  OAI21_X1   g1790(.A1(new_n1742_), .A2(new_n1743_), .B(new_n405_), .ZN(new_n2054_));
  NAND2_X1   g1791(.A1(new_n2053_), .A2(new_n2054_), .ZN(new_n2055_));
  OAI21_X1   g1792(.A1(new_n1749_), .A2(new_n1748_), .B(new_n308_), .ZN(new_n2056_));
  OAI21_X1   g1793(.A1(new_n1724_), .A2(new_n1725_), .B(new_n373_), .ZN(new_n2057_));
  NAND2_X1   g1794(.A1(new_n2057_), .A2(new_n2056_), .ZN(new_n2058_));
  OAI21_X1   g1795(.A1(new_n2055_), .A2(new_n2058_), .B(\shift[6] ), .ZN(new_n2059_));
  NAND2_X1   g1796(.A1(new_n2052_), .A2(new_n2059_), .ZN(\result[29] ));
  OAI21_X1   g1797(.A1(new_n1766_), .A2(new_n1769_), .B(new_n308_), .ZN(new_n2061_));
  OAI21_X1   g1798(.A1(new_n1781_), .A2(new_n1784_), .B(new_n340_), .ZN(new_n2062_));
  NAND2_X1   g1799(.A1(new_n2061_), .A2(new_n2062_), .ZN(new_n2063_));
  OAI21_X1   g1800(.A1(new_n1806_), .A2(new_n1809_), .B(new_n373_), .ZN(new_n2064_));
  OAI21_X1   g1801(.A1(new_n1774_), .A2(new_n1777_), .B(new_n405_), .ZN(new_n2065_));
  NAND2_X1   g1802(.A1(new_n2064_), .A2(new_n2065_), .ZN(new_n2066_));
  OAI21_X1   g1803(.A1(new_n2063_), .A2(new_n2066_), .B(new_n264_), .ZN(new_n2067_));
  OAI21_X1   g1804(.A1(new_n1788_), .A2(new_n1790_), .B(new_n340_), .ZN(new_n2068_));
  OAI21_X1   g1805(.A1(new_n1793_), .A2(new_n1796_), .B(new_n405_), .ZN(new_n2069_));
  NAND2_X1   g1806(.A1(new_n2068_), .A2(new_n2069_), .ZN(new_n2070_));
  OAI21_X1   g1807(.A1(new_n1799_), .A2(new_n1802_), .B(new_n308_), .ZN(new_n2071_));
  OAI21_X1   g1808(.A1(new_n1759_), .A2(new_n1762_), .B(new_n373_), .ZN(new_n2072_));
  NAND2_X1   g1809(.A1(new_n2071_), .A2(new_n2072_), .ZN(new_n2073_));
  OAI21_X1   g1810(.A1(new_n2070_), .A2(new_n2073_), .B(\shift[6] ), .ZN(new_n2074_));
  NAND2_X1   g1811(.A1(new_n2067_), .A2(new_n2074_), .ZN(\result[30] ));
  OAI21_X1   g1812(.A1(new_n1817_), .A2(new_n1818_), .B(new_n308_), .ZN(new_n2076_));
  OAI21_X1   g1813(.A1(new_n1824_), .A2(new_n1825_), .B(new_n340_), .ZN(new_n2077_));
  NAND2_X1   g1814(.A1(new_n2076_), .A2(new_n2077_), .ZN(new_n2078_));
  OAI21_X1   g1815(.A1(new_n1846_), .A2(new_n1847_), .B(new_n373_), .ZN(new_n2079_));
  OAI21_X1   g1816(.A1(new_n1821_), .A2(new_n1822_), .B(new_n405_), .ZN(new_n2080_));
  NAND2_X1   g1817(.A1(new_n2079_), .A2(new_n2080_), .ZN(new_n2081_));
  OAI21_X1   g1818(.A1(new_n2078_), .A2(new_n2081_), .B(new_n264_), .ZN(new_n2082_));
  OAI21_X1   g1819(.A1(new_n1829_), .A2(new_n1830_), .B(new_n340_), .ZN(new_n2083_));
  OAI21_X1   g1820(.A1(new_n1832_), .A2(new_n1833_), .B(new_n405_), .ZN(new_n2084_));
  NAND2_X1   g1821(.A1(new_n2083_), .A2(new_n2084_), .ZN(new_n2085_));
  OAI21_X1   g1822(.A1(new_n1844_), .A2(new_n1843_), .B(new_n308_), .ZN(new_n2086_));
  OAI21_X1   g1823(.A1(new_n1814_), .A2(new_n1815_), .B(new_n373_), .ZN(new_n2087_));
  NAND2_X1   g1824(.A1(new_n2087_), .A2(new_n2086_), .ZN(new_n2088_));
  OAI21_X1   g1825(.A1(new_n2085_), .A2(new_n2088_), .B(\shift[6] ), .ZN(new_n2089_));
  NAND2_X1   g1826(.A1(new_n2082_), .A2(new_n2089_), .ZN(\result[31] ));
  OAI21_X1   g1827(.A1(new_n389_), .A2(new_n404_), .B(new_n308_), .ZN(new_n2091_));
  OAI21_X1   g1828(.A1(new_n357_), .A2(new_n372_), .B(new_n340_), .ZN(new_n2092_));
  NAND2_X1   g1829(.A1(new_n2091_), .A2(new_n2092_), .ZN(new_n2093_));
  OAI21_X1   g1830(.A1(new_n454_), .A2(new_n469_), .B(new_n373_), .ZN(new_n2094_));
  OAI21_X1   g1831(.A1(new_n423_), .A2(new_n438_), .B(new_n405_), .ZN(new_n2095_));
  NAND2_X1   g1832(.A1(new_n2094_), .A2(new_n2095_), .ZN(new_n2096_));
  OAI21_X1   g1833(.A1(new_n2093_), .A2(new_n2096_), .B(new_n264_), .ZN(new_n2097_));
  OAI21_X1   g1834(.A1(new_n286_), .A2(new_n305_), .B(new_n405_), .ZN(new_n2098_));
  OAI21_X1   g1835(.A1(new_n324_), .A2(new_n339_), .B(new_n373_), .ZN(new_n2099_));
  NAND2_X1   g1836(.A1(new_n2098_), .A2(new_n2099_), .ZN(new_n2100_));
  OAI21_X1   g1837(.A1(new_n486_), .A2(new_n501_), .B(new_n340_), .ZN(new_n2101_));
  OAI21_X1   g1838(.A1(new_n517_), .A2(new_n532_), .B(new_n308_), .ZN(new_n2102_));
  NAND2_X1   g1839(.A1(new_n2101_), .A2(new_n2102_), .ZN(new_n2103_));
  OAI21_X1   g1840(.A1(new_n2100_), .A2(new_n2103_), .B(\shift[6] ), .ZN(new_n2104_));
  NAND2_X1   g1841(.A1(new_n2097_), .A2(new_n2104_), .ZN(\result[32] ));
  OAI21_X1   g1842(.A1(new_n636_), .A2(new_n655_), .B(new_n340_), .ZN(new_n2106_));
  OAI21_X1   g1843(.A1(new_n537_), .A2(new_n1867_), .B(new_n2106_), .ZN(new_n2107_));
  OAI21_X1   g1844(.A1(new_n828_), .A2(new_n847_), .B(new_n373_), .ZN(new_n2108_));
  OAI21_X1   g1845(.A1(new_n755_), .A2(new_n774_), .B(new_n405_), .ZN(new_n2109_));
  NAND2_X1   g1846(.A1(new_n2108_), .A2(new_n2109_), .ZN(new_n2110_));
  OAI21_X1   g1847(.A1(new_n2107_), .A2(new_n2110_), .B(new_n264_), .ZN(new_n2111_));
  OAI21_X1   g1848(.A1(new_n716_), .A2(new_n735_), .B(new_n340_), .ZN(new_n2112_));
  OAI21_X1   g1849(.A1(new_n556_), .A2(new_n576_), .B(new_n405_), .ZN(new_n2113_));
  NAND2_X1   g1850(.A1(new_n2112_), .A2(new_n2113_), .ZN(new_n2114_));
  OAI21_X1   g1851(.A1(new_n793_), .A2(new_n808_), .B(new_n308_), .ZN(new_n2115_));
  OAI21_X1   g1852(.A1(new_n596_), .A2(new_n615_), .B(new_n373_), .ZN(new_n2116_));
  NAND2_X1   g1853(.A1(new_n2116_), .A2(new_n2115_), .ZN(new_n2117_));
  OAI21_X1   g1854(.A1(new_n2114_), .A2(new_n2117_), .B(\shift[6] ), .ZN(new_n2118_));
  NAND2_X1   g1855(.A1(new_n2111_), .A2(new_n2118_), .ZN(\result[33] ));
  OAI21_X1   g1856(.A1(new_n942_), .A2(new_n957_), .B(new_n308_), .ZN(new_n2120_));
  OAI21_X1   g1857(.A1(new_n911_), .A2(new_n926_), .B(new_n340_), .ZN(new_n2121_));
  NAND2_X1   g1858(.A1(new_n2120_), .A2(new_n2121_), .ZN(new_n2122_));
  OAI21_X1   g1859(.A1(new_n1044_), .A2(new_n1057_), .B(new_n373_), .ZN(new_n2123_));
  OAI21_X1   g1860(.A1(new_n994_), .A2(new_n1009_), .B(new_n405_), .ZN(new_n2124_));
  NAND2_X1   g1861(.A1(new_n2123_), .A2(new_n2124_), .ZN(new_n2125_));
  OAI21_X1   g1862(.A1(new_n2122_), .A2(new_n2125_), .B(new_n264_), .ZN(new_n2126_));
  OAI21_X1   g1863(.A1(new_n969_), .A2(new_n978_), .B(new_n340_), .ZN(new_n2127_));
  OAI21_X1   g1864(.A1(new_n864_), .A2(new_n871_), .B(new_n405_), .ZN(new_n2128_));
  NAND2_X1   g1865(.A1(new_n2127_), .A2(new_n2128_), .ZN(new_n2129_));
  OAI21_X1   g1866(.A1(new_n1020_), .A2(new_n1032_), .B(new_n308_), .ZN(new_n2130_));
  OAI21_X1   g1867(.A1(new_n885_), .A2(new_n896_), .B(new_n373_), .ZN(new_n2131_));
  NAND2_X1   g1868(.A1(new_n2130_), .A2(new_n2131_), .ZN(new_n2132_));
  OAI21_X1   g1869(.A1(new_n2129_), .A2(new_n2132_), .B(\shift[6] ), .ZN(new_n2133_));
  NAND2_X1   g1870(.A1(new_n2126_), .A2(new_n2133_), .ZN(\result[34] ));
  OAI21_X1   g1871(.A1(new_n1073_), .A2(new_n1084_), .B(new_n308_), .ZN(new_n2135_));
  OAI21_X1   g1872(.A1(new_n1253_), .A2(new_n1264_), .B(new_n373_), .ZN(new_n2136_));
  NAND2_X1   g1873(.A1(new_n2135_), .A2(new_n2136_), .ZN(new_n2137_));
  OAI21_X1   g1874(.A1(new_n1120_), .A2(new_n1131_), .B(new_n340_), .ZN(new_n2138_));
  OAI21_X1   g1875(.A1(new_n1228_), .A2(new_n1239_), .B(new_n405_), .ZN(new_n2139_));
  NAND2_X1   g1876(.A1(new_n2138_), .A2(new_n2139_), .ZN(new_n2140_));
  OAI21_X1   g1877(.A1(new_n2137_), .A2(new_n2140_), .B(new_n264_), .ZN(new_n2141_));
  OAI21_X1   g1878(.A1(new_n1168_), .A2(new_n1180_), .B(new_n340_), .ZN(new_n2142_));
  OAI21_X1   g1879(.A1(new_n1096_), .A2(new_n1107_), .B(new_n373_), .ZN(new_n2143_));
  NAND2_X1   g1880(.A1(new_n2142_), .A2(new_n2143_), .ZN(new_n2144_));
  OAI21_X1   g1881(.A1(new_n1215_), .A2(new_n1196_), .B(new_n308_), .ZN(new_n2145_));
  OAI21_X1   g1882(.A1(new_n1143_), .A2(new_n1154_), .B(new_n405_), .ZN(new_n2146_));
  NAND2_X1   g1883(.A1(new_n2146_), .A2(new_n2145_), .ZN(new_n2147_));
  OAI21_X1   g1884(.A1(new_n2144_), .A2(new_n2147_), .B(\shift[6] ), .ZN(new_n2148_));
  NAND2_X1   g1885(.A1(new_n2141_), .A2(new_n2148_), .ZN(\result[35] ));
  OAI21_X1   g1886(.A1(new_n1290_), .A2(new_n1293_), .B(new_n308_), .ZN(new_n2150_));
  OAI21_X1   g1887(.A1(new_n1283_), .A2(new_n1286_), .B(new_n340_), .ZN(new_n2151_));
  NAND2_X1   g1888(.A1(new_n2150_), .A2(new_n2151_), .ZN(new_n2152_));
  OAI21_X1   g1889(.A1(new_n1314_), .A2(new_n1317_), .B(new_n373_), .ZN(new_n2153_));
  OAI21_X1   g1890(.A1(new_n1321_), .A2(new_n1324_), .B(new_n405_), .ZN(new_n2154_));
  NAND2_X1   g1891(.A1(new_n2153_), .A2(new_n2154_), .ZN(new_n2155_));
  OAI21_X1   g1892(.A1(new_n2152_), .A2(new_n2155_), .B(new_n264_), .ZN(new_n2156_));
  OAI21_X1   g1893(.A1(new_n1270_), .A2(new_n1272_), .B(new_n405_), .ZN(new_n2157_));
  OAI21_X1   g1894(.A1(new_n1275_), .A2(new_n1278_), .B(new_n373_), .ZN(new_n2158_));
  NAND2_X1   g1895(.A1(new_n2157_), .A2(new_n2158_), .ZN(new_n2159_));
  OAI21_X1   g1896(.A1(new_n1306_), .A2(new_n1309_), .B(new_n340_), .ZN(new_n2160_));
  OAI21_X1   g1897(.A1(new_n1299_), .A2(new_n1302_), .B(new_n308_), .ZN(new_n2161_));
  NAND2_X1   g1898(.A1(new_n2160_), .A2(new_n2161_), .ZN(new_n2162_));
  OAI21_X1   g1899(.A1(new_n2159_), .A2(new_n2162_), .B(\shift[6] ), .ZN(new_n2163_));
  NAND2_X1   g1900(.A1(new_n2156_), .A2(new_n2163_), .ZN(\result[36] ));
  OAI21_X1   g1901(.A1(new_n1339_), .A2(new_n1340_), .B(new_n308_), .ZN(new_n2165_));
  OAI21_X1   g1902(.A1(new_n1336_), .A2(new_n1337_), .B(new_n340_), .ZN(new_n2166_));
  NAND2_X1   g1903(.A1(new_n2165_), .A2(new_n2166_), .ZN(new_n2167_));
  OAI21_X1   g1904(.A1(new_n1358_), .A2(new_n1359_), .B(new_n373_), .ZN(new_n2168_));
  OAI21_X1   g1905(.A1(new_n1361_), .A2(new_n1362_), .B(new_n405_), .ZN(new_n2169_));
  NAND2_X1   g1906(.A1(new_n2168_), .A2(new_n2169_), .ZN(new_n2170_));
  OAI21_X1   g1907(.A1(new_n2167_), .A2(new_n2170_), .B(new_n264_), .ZN(new_n2171_));
  OAI21_X1   g1908(.A1(new_n1329_), .A2(new_n1330_), .B(new_n405_), .ZN(new_n2172_));
  OAI21_X1   g1909(.A1(new_n1332_), .A2(new_n1333_), .B(new_n373_), .ZN(new_n2173_));
  NAND2_X1   g1910(.A1(new_n2172_), .A2(new_n2173_), .ZN(new_n2174_));
  OAI21_X1   g1911(.A1(new_n1349_), .A2(new_n1350_), .B(new_n340_), .ZN(new_n2175_));
  OAI21_X1   g1912(.A1(new_n1344_), .A2(new_n1347_), .B(new_n308_), .ZN(new_n2176_));
  NAND2_X1   g1913(.A1(new_n2175_), .A2(new_n2176_), .ZN(new_n2177_));
  OAI21_X1   g1914(.A1(new_n2174_), .A2(new_n2177_), .B(\shift[6] ), .ZN(new_n2178_));
  NAND2_X1   g1915(.A1(new_n2171_), .A2(new_n2178_), .ZN(\result[37] ));
  OAI21_X1   g1916(.A1(new_n1389_), .A2(new_n1392_), .B(new_n308_), .ZN(new_n2180_));
  OAI21_X1   g1917(.A1(new_n1382_), .A2(new_n1385_), .B(new_n340_), .ZN(new_n2181_));
  NAND2_X1   g1918(.A1(new_n2180_), .A2(new_n2181_), .ZN(new_n2182_));
  OAI21_X1   g1919(.A1(new_n1413_), .A2(new_n1416_), .B(new_n373_), .ZN(new_n2183_));
  OAI21_X1   g1920(.A1(new_n1420_), .A2(new_n1423_), .B(new_n405_), .ZN(new_n2184_));
  NAND2_X1   g1921(.A1(new_n2183_), .A2(new_n2184_), .ZN(new_n2185_));
  OAI21_X1   g1922(.A1(new_n2182_), .A2(new_n2185_), .B(new_n264_), .ZN(new_n2186_));
  OAI21_X1   g1923(.A1(new_n1368_), .A2(new_n1370_), .B(new_n405_), .ZN(new_n2187_));
  OAI21_X1   g1924(.A1(new_n1374_), .A2(new_n1377_), .B(new_n373_), .ZN(new_n2188_));
  NAND2_X1   g1925(.A1(new_n2187_), .A2(new_n2188_), .ZN(new_n2189_));
  OAI21_X1   g1926(.A1(new_n1405_), .A2(new_n1408_), .B(new_n340_), .ZN(new_n2190_));
  OAI21_X1   g1927(.A1(new_n1398_), .A2(new_n1401_), .B(new_n308_), .ZN(new_n2191_));
  NAND2_X1   g1928(.A1(new_n2190_), .A2(new_n2191_), .ZN(new_n2192_));
  OAI21_X1   g1929(.A1(new_n2189_), .A2(new_n2192_), .B(\shift[6] ), .ZN(new_n2193_));
  NAND2_X1   g1930(.A1(new_n2186_), .A2(new_n2193_), .ZN(\result[38] ));
  OAI21_X1   g1931(.A1(new_n1455_), .A2(new_n1456_), .B(new_n405_), .ZN(new_n2195_));
  OAI21_X1   g1932(.A1(new_n1452_), .A2(new_n1453_), .B(new_n373_), .ZN(new_n2196_));
  NAND2_X1   g1933(.A1(new_n2195_), .A2(new_n2196_), .ZN(new_n2197_));
  OAI21_X1   g1934(.A1(new_n1435_), .A2(new_n1436_), .B(new_n340_), .ZN(new_n2198_));
  OAI21_X1   g1935(.A1(new_n1438_), .A2(new_n1439_), .B(new_n308_), .ZN(new_n2199_));
  NAND2_X1   g1936(.A1(new_n2198_), .A2(new_n2199_), .ZN(new_n2200_));
  OAI21_X1   g1937(.A1(new_n2197_), .A2(new_n2200_), .B(new_n264_), .ZN(new_n2201_));
  OAI21_X1   g1938(.A1(new_n1446_), .A2(new_n1445_), .B(new_n308_), .ZN(new_n2202_));
  OAI21_X1   g1939(.A1(new_n1448_), .A2(new_n1449_), .B(new_n340_), .ZN(new_n2203_));
  NAND2_X1   g1940(.A1(new_n2203_), .A2(new_n2202_), .ZN(new_n2204_));
  OAI21_X1   g1941(.A1(new_n1431_), .A2(new_n1432_), .B(new_n373_), .ZN(new_n2205_));
  OAI21_X1   g1942(.A1(new_n1428_), .A2(new_n1429_), .B(new_n405_), .ZN(new_n2206_));
  NAND2_X1   g1943(.A1(new_n2205_), .A2(new_n2206_), .ZN(new_n2207_));
  OAI21_X1   g1944(.A1(new_n2207_), .A2(new_n2204_), .B(\shift[6] ), .ZN(new_n2208_));
  NAND2_X1   g1945(.A1(new_n2201_), .A2(new_n2208_), .ZN(\result[39] ));
  OAI21_X1   g1946(.A1(new_n1515_), .A2(new_n1518_), .B(new_n405_), .ZN(new_n2210_));
  OAI21_X1   g1947(.A1(new_n1508_), .A2(new_n1511_), .B(new_n373_), .ZN(new_n2211_));
  NAND2_X1   g1948(.A1(new_n2210_), .A2(new_n2211_), .ZN(new_n2212_));
  OAI21_X1   g1949(.A1(new_n1478_), .A2(new_n1481_), .B(new_n340_), .ZN(new_n2213_));
  OAI21_X1   g1950(.A1(new_n1485_), .A2(new_n1488_), .B(new_n308_), .ZN(new_n2214_));
  NAND2_X1   g1951(.A1(new_n2213_), .A2(new_n2214_), .ZN(new_n2215_));
  OAI21_X1   g1952(.A1(new_n2212_), .A2(new_n2215_), .B(new_n264_), .ZN(new_n2216_));
  OAI21_X1   g1953(.A1(new_n1494_), .A2(new_n1497_), .B(new_n308_), .ZN(new_n2217_));
  OAI21_X1   g1954(.A1(new_n1500_), .A2(new_n1503_), .B(new_n340_), .ZN(new_n2218_));
  NAND2_X1   g1955(.A1(new_n2217_), .A2(new_n2218_), .ZN(new_n2219_));
  OAI21_X1   g1956(.A1(new_n1470_), .A2(new_n1473_), .B(new_n373_), .ZN(new_n2220_));
  OAI21_X1   g1957(.A1(new_n1463_), .A2(new_n1466_), .B(new_n405_), .ZN(new_n2221_));
  NAND2_X1   g1958(.A1(new_n2220_), .A2(new_n2221_), .ZN(new_n2222_));
  OAI21_X1   g1959(.A1(new_n2219_), .A2(new_n2222_), .B(\shift[6] ), .ZN(new_n2223_));
  NAND2_X1   g1960(.A1(new_n2216_), .A2(new_n2223_), .ZN(\result[40] ));
  OAI21_X1   g1961(.A1(new_n1557_), .A2(new_n1558_), .B(new_n405_), .ZN(new_n2225_));
  OAI21_X1   g1962(.A1(new_n1555_), .A2(new_n1554_), .B(new_n373_), .ZN(new_n2226_));
  NAND2_X1   g1963(.A1(new_n2225_), .A2(new_n2226_), .ZN(new_n2227_));
  OAI21_X1   g1964(.A1(new_n1530_), .A2(new_n1531_), .B(new_n340_), .ZN(new_n2228_));
  OAI21_X1   g1965(.A1(new_n1533_), .A2(new_n1534_), .B(new_n308_), .ZN(new_n2229_));
  NAND2_X1   g1966(.A1(new_n2228_), .A2(new_n2229_), .ZN(new_n2230_));
  OAI21_X1   g1967(.A1(new_n2230_), .A2(new_n2227_), .B(new_n264_), .ZN(new_n2231_));
  OAI21_X1   g1968(.A1(new_n1538_), .A2(new_n1546_), .B(new_n308_), .ZN(new_n2232_));
  OAI21_X1   g1969(.A1(new_n1548_), .A2(new_n1549_), .B(new_n340_), .ZN(new_n2233_));
  NAND2_X1   g1970(.A1(new_n2233_), .A2(new_n2232_), .ZN(new_n2234_));
  OAI21_X1   g1971(.A1(new_n1526_), .A2(new_n1527_), .B(new_n373_), .ZN(new_n2235_));
  OAI21_X1   g1972(.A1(new_n1523_), .A2(new_n1524_), .B(new_n405_), .ZN(new_n2236_));
  NAND2_X1   g1973(.A1(new_n2235_), .A2(new_n2236_), .ZN(new_n2237_));
  OAI21_X1   g1974(.A1(new_n2237_), .A2(new_n2234_), .B(\shift[6] ), .ZN(new_n2238_));
  NAND2_X1   g1975(.A1(new_n2231_), .A2(new_n2238_), .ZN(\result[41] ));
  OAI21_X1   g1976(.A1(new_n1587_), .A2(new_n1590_), .B(new_n308_), .ZN(new_n2240_));
  OAI21_X1   g1977(.A1(new_n1580_), .A2(new_n1583_), .B(new_n340_), .ZN(new_n2241_));
  NAND2_X1   g1978(.A1(new_n2240_), .A2(new_n2241_), .ZN(new_n2242_));
  OAI21_X1   g1979(.A1(new_n1608_), .A2(new_n1611_), .B(new_n373_), .ZN(new_n2243_));
  OAI21_X1   g1980(.A1(new_n1615_), .A2(new_n1618_), .B(new_n405_), .ZN(new_n2244_));
  NAND2_X1   g1981(.A1(new_n2243_), .A2(new_n2244_), .ZN(new_n2245_));
  OAI21_X1   g1982(.A1(new_n2242_), .A2(new_n2245_), .B(new_n264_), .ZN(new_n2246_));
  OAI21_X1   g1983(.A1(new_n1595_), .A2(new_n1596_), .B(new_n308_), .ZN(new_n2247_));
  OAI21_X1   g1984(.A1(new_n1600_), .A2(new_n1603_), .B(new_n340_), .ZN(new_n2248_));
  NAND2_X1   g1985(.A1(new_n2247_), .A2(new_n2248_), .ZN(new_n2249_));
  OAI21_X1   g1986(.A1(new_n1572_), .A2(new_n1575_), .B(new_n373_), .ZN(new_n2250_));
  OAI21_X1   g1987(.A1(new_n1565_), .A2(new_n1568_), .B(new_n405_), .ZN(new_n2251_));
  NAND2_X1   g1988(.A1(new_n2250_), .A2(new_n2251_), .ZN(new_n2252_));
  OAI21_X1   g1989(.A1(new_n2249_), .A2(new_n2252_), .B(\shift[6] ), .ZN(new_n2253_));
  NAND2_X1   g1990(.A1(new_n2246_), .A2(new_n2253_), .ZN(\result[42] ));
  OAI21_X1   g1991(.A1(new_n1633_), .A2(new_n1634_), .B(new_n308_), .ZN(new_n2255_));
  OAI21_X1   g1992(.A1(new_n1630_), .A2(new_n1631_), .B(new_n340_), .ZN(new_n2256_));
  NAND2_X1   g1993(.A1(new_n2255_), .A2(new_n2256_), .ZN(new_n2257_));
  OAI21_X1   g1994(.A1(new_n1657_), .A2(new_n1658_), .B(new_n373_), .ZN(new_n2258_));
  OAI21_X1   g1995(.A1(new_n1660_), .A2(new_n1661_), .B(new_n405_), .ZN(new_n2259_));
  NAND2_X1   g1996(.A1(new_n2258_), .A2(new_n2259_), .ZN(new_n2260_));
  OAI21_X1   g1997(.A1(new_n2257_), .A2(new_n2260_), .B(new_n264_), .ZN(new_n2261_));
  OAI21_X1   g1998(.A1(new_n1643_), .A2(new_n1651_), .B(new_n308_), .ZN(new_n2262_));
  OAI21_X1   g1999(.A1(new_n1653_), .A2(new_n1654_), .B(new_n340_), .ZN(new_n2263_));
  NAND2_X1   g2000(.A1(new_n2263_), .A2(new_n2262_), .ZN(new_n2264_));
  OAI21_X1   g2001(.A1(new_n1626_), .A2(new_n1627_), .B(new_n373_), .ZN(new_n2265_));
  OAI21_X1   g2002(.A1(new_n1623_), .A2(new_n1624_), .B(new_n405_), .ZN(new_n2266_));
  NAND2_X1   g2003(.A1(new_n2265_), .A2(new_n2266_), .ZN(new_n2267_));
  OAI21_X1   g2004(.A1(new_n2267_), .A2(new_n2264_), .B(\shift[6] ), .ZN(new_n2268_));
  NAND2_X1   g2005(.A1(new_n2261_), .A2(new_n2268_), .ZN(\result[43] ));
  OAI21_X1   g2006(.A1(new_n1690_), .A2(new_n1693_), .B(new_n308_), .ZN(new_n2270_));
  OAI21_X1   g2007(.A1(new_n1683_), .A2(new_n1686_), .B(new_n340_), .ZN(new_n2271_));
  NAND2_X1   g2008(.A1(new_n2270_), .A2(new_n2271_), .ZN(new_n2272_));
  OAI21_X1   g2009(.A1(new_n1709_), .A2(new_n1712_), .B(new_n373_), .ZN(new_n2273_));
  OAI21_X1   g2010(.A1(new_n1716_), .A2(new_n1719_), .B(new_n405_), .ZN(new_n2274_));
  NAND2_X1   g2011(.A1(new_n2273_), .A2(new_n2274_), .ZN(new_n2275_));
  OAI21_X1   g2012(.A1(new_n2272_), .A2(new_n2275_), .B(new_n264_), .ZN(new_n2276_));
  OAI21_X1   g2013(.A1(new_n1697_), .A2(new_n1699_), .B(new_n308_), .ZN(new_n2277_));
  OAI21_X1   g2014(.A1(new_n1702_), .A2(new_n1705_), .B(new_n340_), .ZN(new_n2278_));
  NAND2_X1   g2015(.A1(new_n2277_), .A2(new_n2278_), .ZN(new_n2279_));
  OAI21_X1   g2016(.A1(new_n1675_), .A2(new_n1678_), .B(new_n373_), .ZN(new_n2280_));
  OAI21_X1   g2017(.A1(new_n1668_), .A2(new_n1671_), .B(new_n405_), .ZN(new_n2281_));
  NAND2_X1   g2018(.A1(new_n2280_), .A2(new_n2281_), .ZN(new_n2282_));
  OAI21_X1   g2019(.A1(new_n2279_), .A2(new_n2282_), .B(\shift[6] ), .ZN(new_n2283_));
  NAND2_X1   g2020(.A1(new_n2276_), .A2(new_n2283_), .ZN(\result[44] ));
  OAI21_X1   g2021(.A1(new_n1734_), .A2(new_n1735_), .B(new_n308_), .ZN(new_n2285_));
  OAI21_X1   g2022(.A1(new_n1731_), .A2(new_n1732_), .B(new_n340_), .ZN(new_n2286_));
  NAND2_X1   g2023(.A1(new_n2285_), .A2(new_n2286_), .ZN(new_n2287_));
  OAI21_X1   g2024(.A1(new_n1749_), .A2(new_n1748_), .B(new_n373_), .ZN(new_n2288_));
  OAI21_X1   g2025(.A1(new_n1751_), .A2(new_n1752_), .B(new_n405_), .ZN(new_n2289_));
  NAND2_X1   g2026(.A1(new_n2289_), .A2(new_n2288_), .ZN(new_n2290_));
  OAI21_X1   g2027(.A1(new_n2287_), .A2(new_n2290_), .B(new_n264_), .ZN(new_n2291_));
  OAI21_X1   g2028(.A1(new_n1739_), .A2(new_n1740_), .B(new_n308_), .ZN(new_n2292_));
  OAI21_X1   g2029(.A1(new_n1742_), .A2(new_n1743_), .B(new_n340_), .ZN(new_n2293_));
  NAND2_X1   g2030(.A1(new_n2292_), .A2(new_n2293_), .ZN(new_n2294_));
  OAI21_X1   g2031(.A1(new_n1727_), .A2(new_n1728_), .B(new_n373_), .ZN(new_n2295_));
  OAI21_X1   g2032(.A1(new_n1724_), .A2(new_n1725_), .B(new_n405_), .ZN(new_n2296_));
  NAND2_X1   g2033(.A1(new_n2295_), .A2(new_n2296_), .ZN(new_n2297_));
  OAI21_X1   g2034(.A1(new_n2294_), .A2(new_n2297_), .B(\shift[6] ), .ZN(new_n2298_));
  NAND2_X1   g2035(.A1(new_n2298_), .A2(new_n2291_), .ZN(\result[45] ));
  OAI21_X1   g2036(.A1(new_n1781_), .A2(new_n1784_), .B(new_n308_), .ZN(new_n2300_));
  OAI21_X1   g2037(.A1(new_n1774_), .A2(new_n1777_), .B(new_n340_), .ZN(new_n2301_));
  NAND2_X1   g2038(.A1(new_n2300_), .A2(new_n2301_), .ZN(new_n2302_));
  OAI21_X1   g2039(.A1(new_n1799_), .A2(new_n1802_), .B(new_n373_), .ZN(new_n2303_));
  OAI21_X1   g2040(.A1(new_n1806_), .A2(new_n1809_), .B(new_n405_), .ZN(new_n2304_));
  NAND2_X1   g2041(.A1(new_n2303_), .A2(new_n2304_), .ZN(new_n2305_));
  OAI21_X1   g2042(.A1(new_n2302_), .A2(new_n2305_), .B(new_n264_), .ZN(new_n2306_));
  OAI21_X1   g2043(.A1(new_n1788_), .A2(new_n1790_), .B(new_n308_), .ZN(new_n2307_));
  OAI21_X1   g2044(.A1(new_n1793_), .A2(new_n1796_), .B(new_n340_), .ZN(new_n2308_));
  NAND2_X1   g2045(.A1(new_n2307_), .A2(new_n2308_), .ZN(new_n2309_));
  OAI21_X1   g2046(.A1(new_n1766_), .A2(new_n1769_), .B(new_n373_), .ZN(new_n2310_));
  OAI21_X1   g2047(.A1(new_n1759_), .A2(new_n1762_), .B(new_n405_), .ZN(new_n2311_));
  NAND2_X1   g2048(.A1(new_n2310_), .A2(new_n2311_), .ZN(new_n2312_));
  OAI21_X1   g2049(.A1(new_n2309_), .A2(new_n2312_), .B(\shift[6] ), .ZN(new_n2313_));
  NAND2_X1   g2050(.A1(new_n2306_), .A2(new_n2313_), .ZN(\result[46] ));
  OAI21_X1   g2051(.A1(new_n1824_), .A2(new_n1825_), .B(new_n308_), .ZN(new_n2315_));
  OAI21_X1   g2052(.A1(new_n1821_), .A2(new_n1822_), .B(new_n340_), .ZN(new_n2316_));
  NAND2_X1   g2053(.A1(new_n2315_), .A2(new_n2316_), .ZN(new_n2317_));
  OAI21_X1   g2054(.A1(new_n1844_), .A2(new_n1843_), .B(new_n373_), .ZN(new_n2318_));
  OAI21_X1   g2055(.A1(new_n1846_), .A2(new_n1847_), .B(new_n405_), .ZN(new_n2319_));
  NAND2_X1   g2056(.A1(new_n2319_), .A2(new_n2318_), .ZN(new_n2320_));
  OAI21_X1   g2057(.A1(new_n2317_), .A2(new_n2320_), .B(new_n264_), .ZN(new_n2321_));
  NOR2_X1    g2058(.A1(new_n1832_), .A2(new_n1833_), .ZN(new_n2322_));
  OAI21_X1   g2059(.A1(new_n1829_), .A2(new_n1830_), .B(new_n308_), .ZN(new_n2323_));
  OAI21_X1   g2060(.A1(new_n1062_), .A2(new_n2322_), .B(new_n2323_), .ZN(new_n2324_));
  OAI21_X1   g2061(.A1(new_n1817_), .A2(new_n1818_), .B(new_n373_), .ZN(new_n2325_));
  OAI21_X1   g2062(.A1(new_n1814_), .A2(new_n1815_), .B(new_n405_), .ZN(new_n2326_));
  NAND2_X1   g2063(.A1(new_n2325_), .A2(new_n2326_), .ZN(new_n2327_));
  OAI21_X1   g2064(.A1(new_n2324_), .A2(new_n2327_), .B(\shift[6] ), .ZN(new_n2328_));
  NAND2_X1   g2065(.A1(new_n2328_), .A2(new_n2321_), .ZN(\result[47] ));
  OAI21_X1   g2066(.A1(new_n357_), .A2(new_n372_), .B(new_n308_), .ZN(new_n2330_));
  OAI21_X1   g2067(.A1(new_n423_), .A2(new_n438_), .B(new_n340_), .ZN(new_n2331_));
  NAND2_X1   g2068(.A1(new_n2330_), .A2(new_n2331_), .ZN(new_n2332_));
  OAI21_X1   g2069(.A1(new_n517_), .A2(new_n532_), .B(new_n373_), .ZN(new_n2333_));
  OAI21_X1   g2070(.A1(new_n454_), .A2(new_n469_), .B(new_n405_), .ZN(new_n2334_));
  NAND2_X1   g2071(.A1(new_n2333_), .A2(new_n2334_), .ZN(new_n2335_));
  OAI21_X1   g2072(.A1(new_n2332_), .A2(new_n2335_), .B(new_n264_), .ZN(new_n2336_));
  OAI21_X1   g2073(.A1(new_n286_), .A2(new_n305_), .B(new_n340_), .ZN(new_n2337_));
  OAI21_X1   g2074(.A1(new_n324_), .A2(new_n339_), .B(new_n405_), .ZN(new_n2338_));
  NAND2_X1   g2075(.A1(new_n2337_), .A2(new_n2338_), .ZN(new_n2339_));
  OAI21_X1   g2076(.A1(new_n486_), .A2(new_n501_), .B(new_n308_), .ZN(new_n2340_));
  OAI21_X1   g2077(.A1(new_n389_), .A2(new_n404_), .B(new_n373_), .ZN(new_n2341_));
  NAND2_X1   g2078(.A1(new_n2340_), .A2(new_n2341_), .ZN(new_n2342_));
  OAI21_X1   g2079(.A1(new_n2339_), .A2(new_n2342_), .B(\shift[6] ), .ZN(new_n2343_));
  NAND2_X1   g2080(.A1(new_n2336_), .A2(new_n2343_), .ZN(\result[48] ));
  OAI21_X1   g2081(.A1(new_n636_), .A2(new_n655_), .B(new_n308_), .ZN(new_n2345_));
  OAI21_X1   g2082(.A1(new_n755_), .A2(new_n774_), .B(new_n340_), .ZN(new_n2346_));
  NAND2_X1   g2083(.A1(new_n2345_), .A2(new_n2346_), .ZN(new_n2347_));
  OAI21_X1   g2084(.A1(new_n793_), .A2(new_n808_), .B(new_n373_), .ZN(new_n2348_));
  OAI21_X1   g2085(.A1(new_n828_), .A2(new_n847_), .B(new_n405_), .ZN(new_n2349_));
  NAND2_X1   g2086(.A1(new_n2349_), .A2(new_n2348_), .ZN(new_n2350_));
  OAI21_X1   g2087(.A1(new_n2347_), .A2(new_n2350_), .B(new_n264_), .ZN(new_n2351_));
  OAI21_X1   g2088(.A1(new_n716_), .A2(new_n735_), .B(new_n308_), .ZN(new_n2352_));
  OAI21_X1   g2089(.A1(new_n1062_), .A2(new_n577_), .B(new_n2352_), .ZN(new_n2353_));
  OAI21_X1   g2090(.A1(new_n675_), .A2(new_n694_), .B(new_n373_), .ZN(new_n2354_));
  OAI21_X1   g2091(.A1(new_n596_), .A2(new_n615_), .B(new_n405_), .ZN(new_n2355_));
  NAND2_X1   g2092(.A1(new_n2354_), .A2(new_n2355_), .ZN(new_n2356_));
  OAI21_X1   g2093(.A1(new_n2353_), .A2(new_n2356_), .B(\shift[6] ), .ZN(new_n2357_));
  NAND2_X1   g2094(.A1(new_n2357_), .A2(new_n2351_), .ZN(\result[49] ));
  OAI21_X1   g2095(.A1(new_n911_), .A2(new_n926_), .B(new_n308_), .ZN(new_n2359_));
  OAI21_X1   g2096(.A1(new_n994_), .A2(new_n1009_), .B(new_n340_), .ZN(new_n2360_));
  NAND2_X1   g2097(.A1(new_n2359_), .A2(new_n2360_), .ZN(new_n2361_));
  OAI21_X1   g2098(.A1(new_n1020_), .A2(new_n1032_), .B(new_n373_), .ZN(new_n2362_));
  OAI21_X1   g2099(.A1(new_n1044_), .A2(new_n1057_), .B(new_n405_), .ZN(new_n2363_));
  NAND2_X1   g2100(.A1(new_n2362_), .A2(new_n2363_), .ZN(new_n2364_));
  OAI21_X1   g2101(.A1(new_n2361_), .A2(new_n2364_), .B(new_n264_), .ZN(new_n2365_));
  OAI21_X1   g2102(.A1(new_n969_), .A2(new_n978_), .B(new_n308_), .ZN(new_n2366_));
  OAI21_X1   g2103(.A1(new_n864_), .A2(new_n871_), .B(new_n340_), .ZN(new_n2367_));
  NAND2_X1   g2104(.A1(new_n2366_), .A2(new_n2367_), .ZN(new_n2368_));
  OAI21_X1   g2105(.A1(new_n942_), .A2(new_n957_), .B(new_n373_), .ZN(new_n2369_));
  OAI21_X1   g2106(.A1(new_n885_), .A2(new_n896_), .B(new_n405_), .ZN(new_n2370_));
  NAND2_X1   g2107(.A1(new_n2369_), .A2(new_n2370_), .ZN(new_n2371_));
  OAI21_X1   g2108(.A1(new_n2368_), .A2(new_n2371_), .B(\shift[6] ), .ZN(new_n2372_));
  NAND2_X1   g2109(.A1(new_n2365_), .A2(new_n2372_), .ZN(\result[50] ));
  OAI21_X1   g2110(.A1(new_n1215_), .A2(new_n1196_), .B(new_n373_), .ZN(new_n2374_));
  OAI21_X1   g2111(.A1(new_n1253_), .A2(new_n1264_), .B(new_n405_), .ZN(new_n2375_));
  NAND2_X1   g2112(.A1(new_n2375_), .A2(new_n2374_), .ZN(new_n2376_));
  OAI21_X1   g2113(.A1(new_n1120_), .A2(new_n1131_), .B(new_n308_), .ZN(new_n2377_));
  OAI21_X1   g2114(.A1(new_n1228_), .A2(new_n1239_), .B(new_n340_), .ZN(new_n2378_));
  NAND2_X1   g2115(.A1(new_n2377_), .A2(new_n2378_), .ZN(new_n2379_));
  OAI21_X1   g2116(.A1(new_n2379_), .A2(new_n2376_), .B(new_n264_), .ZN(new_n2380_));
  OAI21_X1   g2117(.A1(new_n1168_), .A2(new_n1180_), .B(new_n308_), .ZN(new_n2381_));
  OAI21_X1   g2118(.A1(new_n1073_), .A2(new_n1084_), .B(new_n373_), .ZN(new_n2382_));
  NAND2_X1   g2119(.A1(new_n2381_), .A2(new_n2382_), .ZN(new_n2383_));
  OAI21_X1   g2120(.A1(new_n1143_), .A2(new_n1154_), .B(new_n340_), .ZN(new_n2384_));
  OAI21_X1   g2121(.A1(new_n1096_), .A2(new_n1107_), .B(new_n405_), .ZN(new_n2385_));
  NAND2_X1   g2122(.A1(new_n2384_), .A2(new_n2385_), .ZN(new_n2386_));
  OAI21_X1   g2123(.A1(new_n2383_), .A2(new_n2386_), .B(\shift[6] ), .ZN(new_n2387_));
  NAND2_X1   g2124(.A1(new_n2387_), .A2(new_n2380_), .ZN(\result[51] ));
  OAI21_X1   g2125(.A1(new_n1299_), .A2(new_n1302_), .B(new_n373_), .ZN(new_n2389_));
  OAI21_X1   g2126(.A1(new_n1283_), .A2(new_n1286_), .B(new_n308_), .ZN(new_n2390_));
  NAND2_X1   g2127(.A1(new_n2389_), .A2(new_n2390_), .ZN(new_n2391_));
  OAI21_X1   g2128(.A1(new_n1314_), .A2(new_n1317_), .B(new_n405_), .ZN(new_n2392_));
  OAI21_X1   g2129(.A1(new_n1321_), .A2(new_n1324_), .B(new_n340_), .ZN(new_n2393_));
  NAND2_X1   g2130(.A1(new_n2392_), .A2(new_n2393_), .ZN(new_n2394_));
  OAI21_X1   g2131(.A1(new_n2391_), .A2(new_n2394_), .B(new_n264_), .ZN(new_n2395_));
  OAI21_X1   g2132(.A1(new_n1270_), .A2(new_n1272_), .B(new_n340_), .ZN(new_n2396_));
  OAI21_X1   g2133(.A1(new_n1275_), .A2(new_n1278_), .B(new_n405_), .ZN(new_n2397_));
  NAND2_X1   g2134(.A1(new_n2396_), .A2(new_n2397_), .ZN(new_n2398_));
  OAI21_X1   g2135(.A1(new_n1290_), .A2(new_n1293_), .B(new_n373_), .ZN(new_n2399_));
  OAI21_X1   g2136(.A1(new_n1306_), .A2(new_n1309_), .B(new_n308_), .ZN(new_n2400_));
  NAND2_X1   g2137(.A1(new_n2399_), .A2(new_n2400_), .ZN(new_n2401_));
  OAI21_X1   g2138(.A1(new_n2398_), .A2(new_n2401_), .B(\shift[6] ), .ZN(new_n2402_));
  NAND2_X1   g2139(.A1(new_n2395_), .A2(new_n2402_), .ZN(\result[52] ));
  OAI21_X1   g2140(.A1(new_n1344_), .A2(new_n1347_), .B(new_n373_), .ZN(new_n2404_));
  OAI21_X1   g2141(.A1(new_n1336_), .A2(new_n1337_), .B(new_n308_), .ZN(new_n2405_));
  NAND2_X1   g2142(.A1(new_n2405_), .A2(new_n2404_), .ZN(new_n2406_));
  OAI21_X1   g2143(.A1(new_n1358_), .A2(new_n1359_), .B(new_n405_), .ZN(new_n2407_));
  OAI21_X1   g2144(.A1(new_n1361_), .A2(new_n1362_), .B(new_n340_), .ZN(new_n2408_));
  NAND2_X1   g2145(.A1(new_n2407_), .A2(new_n2408_), .ZN(new_n2409_));
  OAI21_X1   g2146(.A1(new_n2409_), .A2(new_n2406_), .B(new_n264_), .ZN(new_n2410_));
  OAI21_X1   g2147(.A1(new_n1332_), .A2(new_n1333_), .B(new_n405_), .ZN(new_n2411_));
  OAI21_X1   g2148(.A1(new_n1062_), .A2(new_n1331_), .B(new_n2411_), .ZN(new_n2412_));
  OAI21_X1   g2149(.A1(new_n1339_), .A2(new_n1340_), .B(new_n373_), .ZN(new_n2413_));
  OAI21_X1   g2150(.A1(new_n1349_), .A2(new_n1350_), .B(new_n308_), .ZN(new_n2414_));
  NAND2_X1   g2151(.A1(new_n2413_), .A2(new_n2414_), .ZN(new_n2415_));
  OAI21_X1   g2152(.A1(new_n2412_), .A2(new_n2415_), .B(\shift[6] ), .ZN(new_n2416_));
  NAND2_X1   g2153(.A1(new_n2416_), .A2(new_n2410_), .ZN(\result[53] ));
  OAI21_X1   g2154(.A1(new_n1398_), .A2(new_n1401_), .B(new_n373_), .ZN(new_n2418_));
  OAI21_X1   g2155(.A1(new_n1382_), .A2(new_n1385_), .B(new_n308_), .ZN(new_n2419_));
  NAND2_X1   g2156(.A1(new_n2418_), .A2(new_n2419_), .ZN(new_n2420_));
  OAI21_X1   g2157(.A1(new_n1413_), .A2(new_n1416_), .B(new_n405_), .ZN(new_n2421_));
  OAI21_X1   g2158(.A1(new_n1420_), .A2(new_n1423_), .B(new_n340_), .ZN(new_n2422_));
  NAND2_X1   g2159(.A1(new_n2421_), .A2(new_n2422_), .ZN(new_n2423_));
  OAI21_X1   g2160(.A1(new_n2420_), .A2(new_n2423_), .B(new_n264_), .ZN(new_n2424_));
  OAI21_X1   g2161(.A1(new_n1368_), .A2(new_n1370_), .B(new_n340_), .ZN(new_n2425_));
  OAI21_X1   g2162(.A1(new_n1374_), .A2(new_n1377_), .B(new_n405_), .ZN(new_n2426_));
  NAND2_X1   g2163(.A1(new_n2425_), .A2(new_n2426_), .ZN(new_n2427_));
  OAI21_X1   g2164(.A1(new_n1389_), .A2(new_n1392_), .B(new_n373_), .ZN(new_n2428_));
  OAI21_X1   g2165(.A1(new_n1405_), .A2(new_n1408_), .B(new_n308_), .ZN(new_n2429_));
  NAND2_X1   g2166(.A1(new_n2428_), .A2(new_n2429_), .ZN(new_n2430_));
  OAI21_X1   g2167(.A1(new_n2427_), .A2(new_n2430_), .B(\shift[6] ), .ZN(new_n2431_));
  NAND2_X1   g2168(.A1(new_n2424_), .A2(new_n2431_), .ZN(\result[54] ));
  OAI21_X1   g2169(.A1(new_n1446_), .A2(new_n1445_), .B(new_n373_), .ZN(new_n2433_));
  OAI21_X1   g2170(.A1(new_n1455_), .A2(new_n1456_), .B(new_n340_), .ZN(new_n2434_));
  NAND2_X1   g2171(.A1(new_n2434_), .A2(new_n2433_), .ZN(new_n2435_));
  OAI21_X1   g2172(.A1(new_n1435_), .A2(new_n1436_), .B(new_n308_), .ZN(new_n2436_));
  OAI21_X1   g2173(.A1(new_n1452_), .A2(new_n1453_), .B(new_n405_), .ZN(new_n2437_));
  NAND2_X1   g2174(.A1(new_n2436_), .A2(new_n2437_), .ZN(new_n2438_));
  OAI21_X1   g2175(.A1(new_n2438_), .A2(new_n2435_), .B(new_n264_), .ZN(new_n2439_));
  OAI21_X1   g2176(.A1(new_n1448_), .A2(new_n1449_), .B(new_n308_), .ZN(new_n2440_));
  OAI21_X1   g2177(.A1(new_n1062_), .A2(new_n1430_), .B(new_n2440_), .ZN(new_n2441_));
  OAI21_X1   g2178(.A1(new_n1438_), .A2(new_n1439_), .B(new_n373_), .ZN(new_n2442_));
  OAI21_X1   g2179(.A1(new_n1431_), .A2(new_n1432_), .B(new_n405_), .ZN(new_n2443_));
  NAND2_X1   g2180(.A1(new_n2442_), .A2(new_n2443_), .ZN(new_n2444_));
  OAI21_X1   g2181(.A1(new_n2441_), .A2(new_n2444_), .B(\shift[6] ), .ZN(new_n2445_));
  NAND2_X1   g2182(.A1(new_n2445_), .A2(new_n2439_), .ZN(\result[55] ));
  OAI21_X1   g2183(.A1(new_n1494_), .A2(new_n1497_), .B(new_n373_), .ZN(new_n2447_));
  OAI21_X1   g2184(.A1(new_n1515_), .A2(new_n1518_), .B(new_n340_), .ZN(new_n2448_));
  NAND2_X1   g2185(.A1(new_n2447_), .A2(new_n2448_), .ZN(new_n2449_));
  OAI21_X1   g2186(.A1(new_n1478_), .A2(new_n1481_), .B(new_n308_), .ZN(new_n2450_));
  OAI21_X1   g2187(.A1(new_n1508_), .A2(new_n1511_), .B(new_n405_), .ZN(new_n2451_));
  NAND2_X1   g2188(.A1(new_n2450_), .A2(new_n2451_), .ZN(new_n2452_));
  OAI21_X1   g2189(.A1(new_n2449_), .A2(new_n2452_), .B(new_n264_), .ZN(new_n2453_));
  OAI21_X1   g2190(.A1(new_n1500_), .A2(new_n1503_), .B(new_n308_), .ZN(new_n2454_));
  OAI21_X1   g2191(.A1(new_n1463_), .A2(new_n1466_), .B(new_n340_), .ZN(new_n2455_));
  NAND2_X1   g2192(.A1(new_n2454_), .A2(new_n2455_), .ZN(new_n2456_));
  OAI21_X1   g2193(.A1(new_n1485_), .A2(new_n1488_), .B(new_n373_), .ZN(new_n2457_));
  OAI21_X1   g2194(.A1(new_n1470_), .A2(new_n1473_), .B(new_n405_), .ZN(new_n2458_));
  NAND2_X1   g2195(.A1(new_n2457_), .A2(new_n2458_), .ZN(new_n2459_));
  OAI21_X1   g2196(.A1(new_n2456_), .A2(new_n2459_), .B(\shift[6] ), .ZN(new_n2460_));
  NAND2_X1   g2197(.A1(new_n2453_), .A2(new_n2460_), .ZN(\result[56] ));
  OAI21_X1   g2198(.A1(new_n1538_), .A2(new_n1546_), .B(new_n373_), .ZN(new_n2462_));
  OAI21_X1   g2199(.A1(new_n1557_), .A2(new_n1558_), .B(new_n340_), .ZN(new_n2463_));
  NAND2_X1   g2200(.A1(new_n2463_), .A2(new_n2462_), .ZN(new_n2464_));
  OAI21_X1   g2201(.A1(new_n1530_), .A2(new_n1531_), .B(new_n308_), .ZN(new_n2465_));
  OAI21_X1   g2202(.A1(new_n1555_), .A2(new_n1554_), .B(new_n405_), .ZN(new_n2466_));
  NAND2_X1   g2203(.A1(new_n2465_), .A2(new_n2466_), .ZN(new_n2467_));
  OAI21_X1   g2204(.A1(new_n2464_), .A2(new_n2467_), .B(new_n264_), .ZN(new_n2468_));
  OAI21_X1   g2205(.A1(new_n1548_), .A2(new_n1549_), .B(new_n308_), .ZN(new_n2469_));
  OAI21_X1   g2206(.A1(new_n1523_), .A2(new_n1524_), .B(new_n340_), .ZN(new_n2470_));
  NAND2_X1   g2207(.A1(new_n2469_), .A2(new_n2470_), .ZN(new_n2471_));
  OAI21_X1   g2208(.A1(new_n1533_), .A2(new_n1534_), .B(new_n373_), .ZN(new_n2472_));
  OAI21_X1   g2209(.A1(new_n1526_), .A2(new_n1527_), .B(new_n405_), .ZN(new_n2473_));
  NAND2_X1   g2210(.A1(new_n2472_), .A2(new_n2473_), .ZN(new_n2474_));
  OAI21_X1   g2211(.A1(new_n2471_), .A2(new_n2474_), .B(\shift[6] ), .ZN(new_n2475_));
  NAND2_X1   g2212(.A1(new_n2475_), .A2(new_n2468_), .ZN(\result[57] ));
  OAI21_X1   g2213(.A1(new_n1595_), .A2(new_n1596_), .B(new_n373_), .ZN(new_n2477_));
  OAI21_X1   g2214(.A1(new_n1580_), .A2(new_n1583_), .B(new_n308_), .ZN(new_n2478_));
  NAND2_X1   g2215(.A1(new_n2477_), .A2(new_n2478_), .ZN(new_n2479_));
  OAI21_X1   g2216(.A1(new_n1608_), .A2(new_n1611_), .B(new_n405_), .ZN(new_n2480_));
  OAI21_X1   g2217(.A1(new_n1615_), .A2(new_n1618_), .B(new_n340_), .ZN(new_n2481_));
  NAND2_X1   g2218(.A1(new_n2480_), .A2(new_n2481_), .ZN(new_n2482_));
  OAI21_X1   g2219(.A1(new_n2479_), .A2(new_n2482_), .B(new_n264_), .ZN(new_n2483_));
  OAI21_X1   g2220(.A1(new_n1600_), .A2(new_n1603_), .B(new_n308_), .ZN(new_n2484_));
  OAI21_X1   g2221(.A1(new_n1565_), .A2(new_n1568_), .B(new_n340_), .ZN(new_n2485_));
  NAND2_X1   g2222(.A1(new_n2484_), .A2(new_n2485_), .ZN(new_n2486_));
  OAI21_X1   g2223(.A1(new_n1587_), .A2(new_n1590_), .B(new_n373_), .ZN(new_n2487_));
  OAI21_X1   g2224(.A1(new_n1572_), .A2(new_n1575_), .B(new_n405_), .ZN(new_n2488_));
  NAND2_X1   g2225(.A1(new_n2487_), .A2(new_n2488_), .ZN(new_n2489_));
  OAI21_X1   g2226(.A1(new_n2486_), .A2(new_n2489_), .B(\shift[6] ), .ZN(new_n2490_));
  NAND2_X1   g2227(.A1(new_n2483_), .A2(new_n2490_), .ZN(\result[58] ));
  OAI21_X1   g2228(.A1(new_n1643_), .A2(new_n1651_), .B(new_n373_), .ZN(new_n2492_));
  OAI21_X1   g2229(.A1(new_n1630_), .A2(new_n1631_), .B(new_n308_), .ZN(new_n2493_));
  NAND2_X1   g2230(.A1(new_n2493_), .A2(new_n2492_), .ZN(new_n2494_));
  OAI21_X1   g2231(.A1(new_n1657_), .A2(new_n1658_), .B(new_n405_), .ZN(new_n2495_));
  OAI21_X1   g2232(.A1(new_n1660_), .A2(new_n1661_), .B(new_n340_), .ZN(new_n2496_));
  NAND2_X1   g2233(.A1(new_n2495_), .A2(new_n2496_), .ZN(new_n2497_));
  OAI21_X1   g2234(.A1(new_n2497_), .A2(new_n2494_), .B(new_n264_), .ZN(new_n2498_));
  OAI21_X1   g2235(.A1(new_n1653_), .A2(new_n1654_), .B(new_n308_), .ZN(new_n2499_));
  OAI21_X1   g2236(.A1(new_n1062_), .A2(new_n1625_), .B(new_n2499_), .ZN(new_n2500_));
  OAI21_X1   g2237(.A1(new_n1633_), .A2(new_n1634_), .B(new_n373_), .ZN(new_n2501_));
  OAI21_X1   g2238(.A1(new_n1626_), .A2(new_n1627_), .B(new_n405_), .ZN(new_n2502_));
  NAND2_X1   g2239(.A1(new_n2501_), .A2(new_n2502_), .ZN(new_n2503_));
  OAI21_X1   g2240(.A1(new_n2500_), .A2(new_n2503_), .B(\shift[6] ), .ZN(new_n2504_));
  NAND2_X1   g2241(.A1(new_n2504_), .A2(new_n2498_), .ZN(\result[59] ));
  OAI21_X1   g2242(.A1(new_n1697_), .A2(new_n1699_), .B(new_n373_), .ZN(new_n2506_));
  OAI21_X1   g2243(.A1(new_n1683_), .A2(new_n1686_), .B(new_n308_), .ZN(new_n2507_));
  NAND2_X1   g2244(.A1(new_n2506_), .A2(new_n2507_), .ZN(new_n2508_));
  OAI21_X1   g2245(.A1(new_n1709_), .A2(new_n1712_), .B(new_n405_), .ZN(new_n2509_));
  OAI21_X1   g2246(.A1(new_n1716_), .A2(new_n1719_), .B(new_n340_), .ZN(new_n2510_));
  NAND2_X1   g2247(.A1(new_n2509_), .A2(new_n2510_), .ZN(new_n2511_));
  OAI21_X1   g2248(.A1(new_n2508_), .A2(new_n2511_), .B(new_n264_), .ZN(new_n2512_));
  OAI21_X1   g2249(.A1(new_n1702_), .A2(new_n1705_), .B(new_n308_), .ZN(new_n2513_));
  OAI21_X1   g2250(.A1(new_n1668_), .A2(new_n1671_), .B(new_n340_), .ZN(new_n2514_));
  NAND2_X1   g2251(.A1(new_n2513_), .A2(new_n2514_), .ZN(new_n2515_));
  OAI21_X1   g2252(.A1(new_n1690_), .A2(new_n1693_), .B(new_n373_), .ZN(new_n2516_));
  OAI21_X1   g2253(.A1(new_n1675_), .A2(new_n1678_), .B(new_n405_), .ZN(new_n2517_));
  NAND2_X1   g2254(.A1(new_n2516_), .A2(new_n2517_), .ZN(new_n2518_));
  OAI21_X1   g2255(.A1(new_n2515_), .A2(new_n2518_), .B(\shift[6] ), .ZN(new_n2519_));
  NAND2_X1   g2256(.A1(new_n2512_), .A2(new_n2519_), .ZN(\result[60] ));
  OAI21_X1   g2257(.A1(new_n1739_), .A2(new_n1740_), .B(new_n373_), .ZN(new_n2521_));
  OAI21_X1   g2258(.A1(new_n1731_), .A2(new_n1732_), .B(new_n308_), .ZN(new_n2522_));
  NAND2_X1   g2259(.A1(new_n2521_), .A2(new_n2522_), .ZN(new_n2523_));
  OAI21_X1   g2260(.A1(new_n1749_), .A2(new_n1748_), .B(new_n405_), .ZN(new_n2524_));
  OAI21_X1   g2261(.A1(new_n1751_), .A2(new_n1752_), .B(new_n340_), .ZN(new_n2525_));
  NAND2_X1   g2262(.A1(new_n2525_), .A2(new_n2524_), .ZN(new_n2526_));
  OAI21_X1   g2263(.A1(new_n2523_), .A2(new_n2526_), .B(new_n264_), .ZN(new_n2527_));
  OAI21_X1   g2264(.A1(new_n1742_), .A2(new_n1743_), .B(new_n308_), .ZN(new_n2528_));
  OAI21_X1   g2265(.A1(new_n1062_), .A2(new_n1726_), .B(new_n2528_), .ZN(new_n2529_));
  OAI21_X1   g2266(.A1(new_n1734_), .A2(new_n1735_), .B(new_n373_), .ZN(new_n2530_));
  OAI21_X1   g2267(.A1(new_n1727_), .A2(new_n1728_), .B(new_n405_), .ZN(new_n2531_));
  NAND2_X1   g2268(.A1(new_n2530_), .A2(new_n2531_), .ZN(new_n2532_));
  OAI21_X1   g2269(.A1(new_n2529_), .A2(new_n2532_), .B(\shift[6] ), .ZN(new_n2533_));
  NAND2_X1   g2270(.A1(new_n2533_), .A2(new_n2527_), .ZN(\result[61] ));
  OAI21_X1   g2271(.A1(new_n1788_), .A2(new_n1790_), .B(new_n373_), .ZN(new_n2535_));
  OAI21_X1   g2272(.A1(new_n1774_), .A2(new_n1777_), .B(new_n308_), .ZN(new_n2536_));
  NAND2_X1   g2273(.A1(new_n2535_), .A2(new_n2536_), .ZN(new_n2537_));
  OAI21_X1   g2274(.A1(new_n1799_), .A2(new_n1802_), .B(new_n405_), .ZN(new_n2538_));
  OAI21_X1   g2275(.A1(new_n1806_), .A2(new_n1809_), .B(new_n340_), .ZN(new_n2539_));
  NAND2_X1   g2276(.A1(new_n2538_), .A2(new_n2539_), .ZN(new_n2540_));
  OAI21_X1   g2277(.A1(new_n2537_), .A2(new_n2540_), .B(new_n264_), .ZN(new_n2541_));
  OAI21_X1   g2278(.A1(new_n1793_), .A2(new_n1796_), .B(new_n308_), .ZN(new_n2542_));
  OAI21_X1   g2279(.A1(new_n1759_), .A2(new_n1762_), .B(new_n340_), .ZN(new_n2543_));
  NAND2_X1   g2280(.A1(new_n2542_), .A2(new_n2543_), .ZN(new_n2544_));
  OAI21_X1   g2281(.A1(new_n1781_), .A2(new_n1784_), .B(new_n373_), .ZN(new_n2545_));
  OAI21_X1   g2282(.A1(new_n1766_), .A2(new_n1769_), .B(new_n405_), .ZN(new_n2546_));
  NAND2_X1   g2283(.A1(new_n2545_), .A2(new_n2546_), .ZN(new_n2547_));
  OAI21_X1   g2284(.A1(new_n2544_), .A2(new_n2547_), .B(\shift[6] ), .ZN(new_n2548_));
  NAND2_X1   g2285(.A1(new_n2541_), .A2(new_n2548_), .ZN(\result[62] ));
  OAI21_X1   g2286(.A1(new_n1829_), .A2(new_n1830_), .B(new_n373_), .ZN(new_n2550_));
  OAI21_X1   g2287(.A1(new_n1821_), .A2(new_n1822_), .B(new_n308_), .ZN(new_n2551_));
  NAND2_X1   g2288(.A1(new_n2550_), .A2(new_n2551_), .ZN(new_n2552_));
  OAI21_X1   g2289(.A1(new_n1844_), .A2(new_n1843_), .B(new_n405_), .ZN(new_n2553_));
  OAI21_X1   g2290(.A1(new_n1846_), .A2(new_n1847_), .B(new_n340_), .ZN(new_n2554_));
  NAND2_X1   g2291(.A1(new_n2554_), .A2(new_n2553_), .ZN(new_n2555_));
  OAI21_X1   g2292(.A1(new_n2552_), .A2(new_n2555_), .B(new_n264_), .ZN(new_n2556_));
  OAI21_X1   g2293(.A1(new_n1814_), .A2(new_n1815_), .B(new_n340_), .ZN(new_n2557_));
  OAI21_X1   g2294(.A1(new_n537_), .A2(new_n2322_), .B(new_n2557_), .ZN(new_n2558_));
  OAI21_X1   g2295(.A1(new_n1824_), .A2(new_n1825_), .B(new_n373_), .ZN(new_n2559_));
  OAI21_X1   g2296(.A1(new_n1817_), .A2(new_n1818_), .B(new_n405_), .ZN(new_n2560_));
  NAND2_X1   g2297(.A1(new_n2559_), .A2(new_n2560_), .ZN(new_n2561_));
  OAI21_X1   g2298(.A1(new_n2558_), .A2(new_n2561_), .B(\shift[6] ), .ZN(new_n2562_));
  NAND2_X1   g2299(.A1(new_n2562_), .A2(new_n2556_), .ZN(\result[63] ));
  OAI21_X1   g2300(.A1(new_n471_), .A2(new_n534_), .B(new_n264_), .ZN(new_n2564_));
  OAI21_X1   g2301(.A1(new_n342_), .A2(new_n407_), .B(\shift[6] ), .ZN(new_n2565_));
  NAND2_X1   g2302(.A1(new_n2564_), .A2(new_n2565_), .ZN(\result[64] ));
  OAI21_X1   g2303(.A1(new_n776_), .A2(new_n849_), .B(new_n264_), .ZN(new_n2567_));
  OAI21_X1   g2304(.A1(new_n617_), .A2(new_n696_), .B(\shift[6] ), .ZN(new_n2568_));
  NAND2_X1   g2305(.A1(new_n2568_), .A2(new_n2567_), .ZN(\result[65] ));
  OAI21_X1   g2306(.A1(new_n1011_), .A2(new_n1059_), .B(new_n264_), .ZN(new_n2570_));
  OAI21_X1   g2307(.A1(new_n898_), .A2(new_n959_), .B(\shift[6] ), .ZN(new_n2571_));
  NAND2_X1   g2308(.A1(new_n2570_), .A2(new_n2571_), .ZN(\result[66] ));
  OAI21_X1   g2309(.A1(new_n1266_), .A2(new_n1217_), .B(new_n264_), .ZN(new_n2573_));
  OAI21_X1   g2310(.A1(new_n1109_), .A2(new_n1156_), .B(\shift[6] ), .ZN(new_n2574_));
  NAND2_X1   g2311(.A1(new_n2574_), .A2(new_n2573_), .ZN(\result[67] ));
  OAI21_X1   g2312(.A1(new_n1311_), .A2(new_n1326_), .B(new_n264_), .ZN(new_n2576_));
  OAI21_X1   g2313(.A1(new_n1280_), .A2(new_n1295_), .B(\shift[6] ), .ZN(new_n2577_));
  NAND2_X1   g2314(.A1(new_n2576_), .A2(new_n2577_), .ZN(\result[68] ));
  OAI21_X1   g2315(.A1(new_n1364_), .A2(new_n1352_), .B(new_n264_), .ZN(new_n2579_));
  OAI21_X1   g2316(.A1(new_n1335_), .A2(new_n1342_), .B(\shift[6] ), .ZN(new_n2580_));
  NAND2_X1   g2317(.A1(new_n2580_), .A2(new_n2579_), .ZN(\result[69] ));
  OAI21_X1   g2318(.A1(new_n1410_), .A2(new_n1425_), .B(new_n264_), .ZN(new_n2582_));
  OAI21_X1   g2319(.A1(new_n1379_), .A2(new_n1394_), .B(\shift[6] ), .ZN(new_n2583_));
  NAND2_X1   g2320(.A1(new_n2582_), .A2(new_n2583_), .ZN(\result[70] ));
  OAI21_X1   g2321(.A1(new_n1458_), .A2(new_n1451_), .B(new_n264_), .ZN(new_n2585_));
  OAI21_X1   g2322(.A1(new_n1434_), .A2(new_n1441_), .B(\shift[6] ), .ZN(new_n2586_));
  NAND2_X1   g2323(.A1(new_n2586_), .A2(new_n2585_), .ZN(\result[71] ));
  OAI21_X1   g2324(.A1(new_n1505_), .A2(new_n1520_), .B(new_n264_), .ZN(new_n2588_));
  OAI21_X1   g2325(.A1(new_n1475_), .A2(new_n1490_), .B(\shift[6] ), .ZN(new_n2589_));
  NAND2_X1   g2326(.A1(new_n2588_), .A2(new_n2589_), .ZN(\result[72] ));
  OAI21_X1   g2327(.A1(new_n1551_), .A2(new_n1560_), .B(new_n264_), .ZN(new_n2591_));
  OAI21_X1   g2328(.A1(new_n1529_), .A2(new_n1536_), .B(\shift[6] ), .ZN(new_n2592_));
  NAND2_X1   g2329(.A1(new_n2592_), .A2(new_n2591_), .ZN(\result[73] ));
  OAI21_X1   g2330(.A1(new_n1605_), .A2(new_n1620_), .B(new_n264_), .ZN(new_n2594_));
  OAI21_X1   g2331(.A1(new_n1577_), .A2(new_n1592_), .B(\shift[6] ), .ZN(new_n2595_));
  NAND2_X1   g2332(.A1(new_n2594_), .A2(new_n2595_), .ZN(\result[74] ));
  OAI21_X1   g2333(.A1(new_n1663_), .A2(new_n1656_), .B(new_n264_), .ZN(new_n2597_));
  OAI21_X1   g2334(.A1(new_n1629_), .A2(new_n1636_), .B(\shift[6] ), .ZN(new_n2598_));
  NAND2_X1   g2335(.A1(new_n2598_), .A2(new_n2597_), .ZN(\result[75] ));
  OAI21_X1   g2336(.A1(new_n1707_), .A2(new_n1721_), .B(new_n264_), .ZN(new_n2600_));
  OAI21_X1   g2337(.A1(new_n1680_), .A2(new_n1695_), .B(\shift[6] ), .ZN(new_n2601_));
  NAND2_X1   g2338(.A1(new_n2600_), .A2(new_n2601_), .ZN(\result[76] ));
  OAI21_X1   g2339(.A1(new_n1745_), .A2(new_n1754_), .B(new_n264_), .ZN(new_n2603_));
  OAI21_X1   g2340(.A1(new_n1730_), .A2(new_n1737_), .B(\shift[6] ), .ZN(new_n2604_));
  NAND2_X1   g2341(.A1(new_n2604_), .A2(new_n2603_), .ZN(\result[77] ));
  OAI21_X1   g2342(.A1(new_n1798_), .A2(new_n1811_), .B(new_n264_), .ZN(new_n2606_));
  OAI21_X1   g2343(.A1(new_n1771_), .A2(new_n1786_), .B(\shift[6] ), .ZN(new_n2607_));
  NAND2_X1   g2344(.A1(new_n2606_), .A2(new_n2607_), .ZN(\result[78] ));
  OAI21_X1   g2345(.A1(new_n1835_), .A2(new_n1849_), .B(new_n264_), .ZN(new_n2609_));
  OAI21_X1   g2346(.A1(new_n1820_), .A2(new_n1827_), .B(\shift[6] ), .ZN(new_n2610_));
  NAND2_X1   g2347(.A1(new_n2610_), .A2(new_n2609_), .ZN(\result[79] ));
  OAI21_X1   g2348(.A1(new_n1861_), .A2(new_n1864_), .B(new_n264_), .ZN(new_n2612_));
  OAI21_X1   g2349(.A1(new_n1854_), .A2(new_n1857_), .B(\shift[6] ), .ZN(new_n2613_));
  NAND2_X1   g2350(.A1(new_n2612_), .A2(new_n2613_), .ZN(\result[80] ));
  OAI21_X1   g2351(.A1(new_n1876_), .A2(new_n1879_), .B(new_n264_), .ZN(new_n2615_));
  OAI21_X1   g2352(.A1(new_n1869_), .A2(new_n1872_), .B(\shift[6] ), .ZN(new_n2616_));
  NAND2_X1   g2353(.A1(new_n2616_), .A2(new_n2615_), .ZN(\result[81] ));
  OAI21_X1   g2354(.A1(new_n1891_), .A2(new_n1894_), .B(new_n264_), .ZN(new_n2618_));
  OAI21_X1   g2355(.A1(new_n1884_), .A2(new_n1887_), .B(\shift[6] ), .ZN(new_n2619_));
  NAND2_X1   g2356(.A1(new_n2618_), .A2(new_n2619_), .ZN(\result[82] ));
  OAI21_X1   g2357(.A1(new_n1905_), .A2(new_n1908_), .B(new_n264_), .ZN(new_n2621_));
  OAI21_X1   g2358(.A1(new_n1898_), .A2(new_n1901_), .B(\shift[6] ), .ZN(new_n2622_));
  NAND2_X1   g2359(.A1(new_n2622_), .A2(new_n2621_), .ZN(\result[83] ));
  OAI21_X1   g2360(.A1(new_n1920_), .A2(new_n1923_), .B(new_n264_), .ZN(new_n2624_));
  OAI21_X1   g2361(.A1(new_n1913_), .A2(new_n1916_), .B(\shift[6] ), .ZN(new_n2625_));
  NAND2_X1   g2362(.A1(new_n2624_), .A2(new_n2625_), .ZN(\result[84] ));
  OAI21_X1   g2363(.A1(new_n1938_), .A2(new_n1935_), .B(new_n264_), .ZN(new_n2627_));
  OAI21_X1   g2364(.A1(new_n1928_), .A2(new_n1931_), .B(\shift[6] ), .ZN(new_n2628_));
  NAND2_X1   g2365(.A1(new_n2628_), .A2(new_n2627_), .ZN(\result[85] ));
  OAI21_X1   g2366(.A1(new_n1950_), .A2(new_n1953_), .B(new_n264_), .ZN(new_n2630_));
  OAI21_X1   g2367(.A1(new_n1943_), .A2(new_n1946_), .B(\shift[6] ), .ZN(new_n2631_));
  NAND2_X1   g2368(.A1(new_n2630_), .A2(new_n2631_), .ZN(\result[86] ));
  OAI21_X1   g2369(.A1(new_n1968_), .A2(new_n1965_), .B(new_n264_), .ZN(new_n2633_));
  OAI21_X1   g2370(.A1(new_n1958_), .A2(new_n1961_), .B(\shift[6] ), .ZN(new_n2634_));
  NAND2_X1   g2371(.A1(new_n2634_), .A2(new_n2633_), .ZN(\result[87] ));
  OAI21_X1   g2372(.A1(new_n1980_), .A2(new_n1983_), .B(new_n264_), .ZN(new_n2636_));
  OAI21_X1   g2373(.A1(new_n1973_), .A2(new_n1976_), .B(\shift[6] ), .ZN(new_n2637_));
  NAND2_X1   g2374(.A1(new_n2636_), .A2(new_n2637_), .ZN(\result[88] ));
  OAI21_X1   g2375(.A1(new_n1995_), .A2(new_n1998_), .B(new_n264_), .ZN(new_n2639_));
  OAI21_X1   g2376(.A1(new_n1988_), .A2(new_n1991_), .B(\shift[6] ), .ZN(new_n2640_));
  NAND2_X1   g2377(.A1(new_n2640_), .A2(new_n2639_), .ZN(\result[89] ));
  OAI21_X1   g2378(.A1(new_n2010_), .A2(new_n2013_), .B(new_n264_), .ZN(new_n2642_));
  OAI21_X1   g2379(.A1(new_n2003_), .A2(new_n2006_), .B(\shift[6] ), .ZN(new_n2643_));
  NAND2_X1   g2380(.A1(new_n2642_), .A2(new_n2643_), .ZN(\result[90] ));
  OAI21_X1   g2381(.A1(new_n2028_), .A2(new_n2025_), .B(new_n264_), .ZN(new_n2645_));
  OAI21_X1   g2382(.A1(new_n2018_), .A2(new_n2021_), .B(\shift[6] ), .ZN(new_n2646_));
  NAND2_X1   g2383(.A1(new_n2646_), .A2(new_n2645_), .ZN(\result[91] ));
  OAI21_X1   g2384(.A1(new_n2040_), .A2(new_n2043_), .B(new_n264_), .ZN(new_n2648_));
  OAI21_X1   g2385(.A1(new_n2033_), .A2(new_n2036_), .B(\shift[6] ), .ZN(new_n2649_));
  NAND2_X1   g2386(.A1(new_n2648_), .A2(new_n2649_), .ZN(\result[92] ));
  OAI21_X1   g2387(.A1(new_n2055_), .A2(new_n2058_), .B(new_n264_), .ZN(new_n2651_));
  OAI21_X1   g2388(.A1(new_n2048_), .A2(new_n2051_), .B(\shift[6] ), .ZN(new_n2652_));
  NAND2_X1   g2389(.A1(new_n2652_), .A2(new_n2651_), .ZN(\result[93] ));
  OAI21_X1   g2390(.A1(new_n2070_), .A2(new_n2073_), .B(new_n264_), .ZN(new_n2654_));
  OAI21_X1   g2391(.A1(new_n2063_), .A2(new_n2066_), .B(\shift[6] ), .ZN(new_n2655_));
  NAND2_X1   g2392(.A1(new_n2654_), .A2(new_n2655_), .ZN(\result[94] ));
  OAI21_X1   g2393(.A1(new_n2085_), .A2(new_n2088_), .B(new_n264_), .ZN(new_n2657_));
  OAI21_X1   g2394(.A1(new_n2078_), .A2(new_n2081_), .B(\shift[6] ), .ZN(new_n2658_));
  NAND2_X1   g2395(.A1(new_n2658_), .A2(new_n2657_), .ZN(\result[95] ));
  OAI21_X1   g2396(.A1(new_n2100_), .A2(new_n2103_), .B(new_n264_), .ZN(new_n2660_));
  OAI21_X1   g2397(.A1(new_n2093_), .A2(new_n2096_), .B(\shift[6] ), .ZN(new_n2661_));
  NAND2_X1   g2398(.A1(new_n2660_), .A2(new_n2661_), .ZN(\result[96] ));
  OAI21_X1   g2399(.A1(new_n2114_), .A2(new_n2117_), .B(new_n264_), .ZN(new_n2663_));
  OAI21_X1   g2400(.A1(new_n2107_), .A2(new_n2110_), .B(\shift[6] ), .ZN(new_n2664_));
  NAND2_X1   g2401(.A1(new_n2664_), .A2(new_n2663_), .ZN(\result[97] ));
  OAI21_X1   g2402(.A1(new_n2129_), .A2(new_n2132_), .B(new_n264_), .ZN(new_n2666_));
  OAI21_X1   g2403(.A1(new_n2122_), .A2(new_n2125_), .B(\shift[6] ), .ZN(new_n2667_));
  NAND2_X1   g2404(.A1(new_n2666_), .A2(new_n2667_), .ZN(\result[98] ));
  OAI21_X1   g2405(.A1(new_n2144_), .A2(new_n2147_), .B(new_n264_), .ZN(new_n2669_));
  OAI21_X1   g2406(.A1(new_n2137_), .A2(new_n2140_), .B(\shift[6] ), .ZN(new_n2670_));
  NAND2_X1   g2407(.A1(new_n2670_), .A2(new_n2669_), .ZN(\result[99] ));
  OAI21_X1   g2408(.A1(new_n2159_), .A2(new_n2162_), .B(new_n264_), .ZN(new_n2672_));
  OAI21_X1   g2409(.A1(new_n2152_), .A2(new_n2155_), .B(\shift[6] ), .ZN(new_n2673_));
  NAND2_X1   g2410(.A1(new_n2672_), .A2(new_n2673_), .ZN(\result[100] ));
  OAI21_X1   g2411(.A1(new_n2174_), .A2(new_n2177_), .B(new_n264_), .ZN(new_n2675_));
  OAI21_X1   g2412(.A1(new_n2167_), .A2(new_n2170_), .B(\shift[6] ), .ZN(new_n2676_));
  NAND2_X1   g2413(.A1(new_n2676_), .A2(new_n2675_), .ZN(\result[101] ));
  OAI21_X1   g2414(.A1(new_n2189_), .A2(new_n2192_), .B(new_n264_), .ZN(new_n2678_));
  OAI21_X1   g2415(.A1(new_n2182_), .A2(new_n2185_), .B(\shift[6] ), .ZN(new_n2679_));
  NAND2_X1   g2416(.A1(new_n2678_), .A2(new_n2679_), .ZN(\result[102] ));
  OAI21_X1   g2417(.A1(new_n2207_), .A2(new_n2204_), .B(new_n264_), .ZN(new_n2681_));
  OAI21_X1   g2418(.A1(new_n2197_), .A2(new_n2200_), .B(\shift[6] ), .ZN(new_n2682_));
  NAND2_X1   g2419(.A1(new_n2682_), .A2(new_n2681_), .ZN(\result[103] ));
  OAI21_X1   g2420(.A1(new_n2219_), .A2(new_n2222_), .B(new_n264_), .ZN(new_n2684_));
  OAI21_X1   g2421(.A1(new_n2212_), .A2(new_n2215_), .B(\shift[6] ), .ZN(new_n2685_));
  NAND2_X1   g2422(.A1(new_n2684_), .A2(new_n2685_), .ZN(\result[104] ));
  OAI21_X1   g2423(.A1(new_n2237_), .A2(new_n2234_), .B(new_n264_), .ZN(new_n2687_));
  OAI21_X1   g2424(.A1(new_n2230_), .A2(new_n2227_), .B(\shift[6] ), .ZN(new_n2688_));
  NAND2_X1   g2425(.A1(new_n2687_), .A2(new_n2688_), .ZN(\result[105] ));
  OAI21_X1   g2426(.A1(new_n2249_), .A2(new_n2252_), .B(new_n264_), .ZN(new_n2690_));
  OAI21_X1   g2427(.A1(new_n2242_), .A2(new_n2245_), .B(\shift[6] ), .ZN(new_n2691_));
  NAND2_X1   g2428(.A1(new_n2690_), .A2(new_n2691_), .ZN(\result[106] ));
  OAI21_X1   g2429(.A1(new_n2267_), .A2(new_n2264_), .B(new_n264_), .ZN(new_n2693_));
  OAI21_X1   g2430(.A1(new_n2257_), .A2(new_n2260_), .B(\shift[6] ), .ZN(new_n2694_));
  NAND2_X1   g2431(.A1(new_n2694_), .A2(new_n2693_), .ZN(\result[107] ));
  OAI21_X1   g2432(.A1(new_n2279_), .A2(new_n2282_), .B(new_n264_), .ZN(new_n2696_));
  OAI21_X1   g2433(.A1(new_n2272_), .A2(new_n2275_), .B(\shift[6] ), .ZN(new_n2697_));
  NAND2_X1   g2434(.A1(new_n2696_), .A2(new_n2697_), .ZN(\result[108] ));
  OAI21_X1   g2435(.A1(new_n2294_), .A2(new_n2297_), .B(new_n264_), .ZN(new_n2699_));
  OAI21_X1   g2436(.A1(new_n2287_), .A2(new_n2290_), .B(\shift[6] ), .ZN(new_n2700_));
  NAND2_X1   g2437(.A1(new_n2699_), .A2(new_n2700_), .ZN(\result[109] ));
  OAI21_X1   g2438(.A1(new_n2309_), .A2(new_n2312_), .B(new_n264_), .ZN(new_n2702_));
  OAI21_X1   g2439(.A1(new_n2302_), .A2(new_n2305_), .B(\shift[6] ), .ZN(new_n2703_));
  NAND2_X1   g2440(.A1(new_n2702_), .A2(new_n2703_), .ZN(\result[110] ));
  OAI21_X1   g2441(.A1(new_n2324_), .A2(new_n2327_), .B(new_n264_), .ZN(new_n2705_));
  OAI21_X1   g2442(.A1(new_n2317_), .A2(new_n2320_), .B(\shift[6] ), .ZN(new_n2706_));
  NAND2_X1   g2443(.A1(new_n2705_), .A2(new_n2706_), .ZN(\result[111] ));
  OAI21_X1   g2444(.A1(new_n2339_), .A2(new_n2342_), .B(new_n264_), .ZN(new_n2708_));
  OAI21_X1   g2445(.A1(new_n2332_), .A2(new_n2335_), .B(\shift[6] ), .ZN(new_n2709_));
  NAND2_X1   g2446(.A1(new_n2708_), .A2(new_n2709_), .ZN(\result[112] ));
  OAI21_X1   g2447(.A1(new_n2353_), .A2(new_n2356_), .B(new_n264_), .ZN(new_n2711_));
  OAI21_X1   g2448(.A1(new_n2347_), .A2(new_n2350_), .B(\shift[6] ), .ZN(new_n2712_));
  NAND2_X1   g2449(.A1(new_n2711_), .A2(new_n2712_), .ZN(\result[113] ));
  OAI21_X1   g2450(.A1(new_n2368_), .A2(new_n2371_), .B(new_n264_), .ZN(new_n2714_));
  OAI21_X1   g2451(.A1(new_n2361_), .A2(new_n2364_), .B(\shift[6] ), .ZN(new_n2715_));
  NAND2_X1   g2452(.A1(new_n2714_), .A2(new_n2715_), .ZN(\result[114] ));
  OAI21_X1   g2453(.A1(new_n2383_), .A2(new_n2386_), .B(new_n264_), .ZN(new_n2717_));
  OAI21_X1   g2454(.A1(new_n2379_), .A2(new_n2376_), .B(\shift[6] ), .ZN(new_n2718_));
  NAND2_X1   g2455(.A1(new_n2717_), .A2(new_n2718_), .ZN(\result[115] ));
  OAI21_X1   g2456(.A1(new_n2398_), .A2(new_n2401_), .B(new_n264_), .ZN(new_n2720_));
  OAI21_X1   g2457(.A1(new_n2391_), .A2(new_n2394_), .B(\shift[6] ), .ZN(new_n2721_));
  NAND2_X1   g2458(.A1(new_n2720_), .A2(new_n2721_), .ZN(\result[116] ));
  OAI21_X1   g2459(.A1(new_n2412_), .A2(new_n2415_), .B(new_n264_), .ZN(new_n2723_));
  OAI21_X1   g2460(.A1(new_n2409_), .A2(new_n2406_), .B(\shift[6] ), .ZN(new_n2724_));
  NAND2_X1   g2461(.A1(new_n2723_), .A2(new_n2724_), .ZN(\result[117] ));
  OAI21_X1   g2462(.A1(new_n2427_), .A2(new_n2430_), .B(new_n264_), .ZN(new_n2726_));
  OAI21_X1   g2463(.A1(new_n2420_), .A2(new_n2423_), .B(\shift[6] ), .ZN(new_n2727_));
  NAND2_X1   g2464(.A1(new_n2726_), .A2(new_n2727_), .ZN(\result[118] ));
  OAI21_X1   g2465(.A1(new_n2441_), .A2(new_n2444_), .B(new_n264_), .ZN(new_n2729_));
  OAI21_X1   g2466(.A1(new_n2438_), .A2(new_n2435_), .B(\shift[6] ), .ZN(new_n2730_));
  NAND2_X1   g2467(.A1(new_n2729_), .A2(new_n2730_), .ZN(\result[119] ));
  OAI21_X1   g2468(.A1(new_n2456_), .A2(new_n2459_), .B(new_n264_), .ZN(new_n2732_));
  OAI21_X1   g2469(.A1(new_n2449_), .A2(new_n2452_), .B(\shift[6] ), .ZN(new_n2733_));
  NAND2_X1   g2470(.A1(new_n2732_), .A2(new_n2733_), .ZN(\result[120] ));
  OAI21_X1   g2471(.A1(new_n2471_), .A2(new_n2474_), .B(new_n264_), .ZN(new_n2735_));
  OAI21_X1   g2472(.A1(new_n2464_), .A2(new_n2467_), .B(\shift[6] ), .ZN(new_n2736_));
  NAND2_X1   g2473(.A1(new_n2735_), .A2(new_n2736_), .ZN(\result[121] ));
  OAI21_X1   g2474(.A1(new_n2486_), .A2(new_n2489_), .B(new_n264_), .ZN(new_n2738_));
  OAI21_X1   g2475(.A1(new_n2479_), .A2(new_n2482_), .B(\shift[6] ), .ZN(new_n2739_));
  NAND2_X1   g2476(.A1(new_n2738_), .A2(new_n2739_), .ZN(\result[122] ));
  OAI21_X1   g2477(.A1(new_n2500_), .A2(new_n2503_), .B(new_n264_), .ZN(new_n2741_));
  OAI21_X1   g2478(.A1(new_n2497_), .A2(new_n2494_), .B(\shift[6] ), .ZN(new_n2742_));
  NAND2_X1   g2479(.A1(new_n2741_), .A2(new_n2742_), .ZN(\result[123] ));
  OAI21_X1   g2480(.A1(new_n2515_), .A2(new_n2518_), .B(new_n264_), .ZN(new_n2744_));
  OAI21_X1   g2481(.A1(new_n2508_), .A2(new_n2511_), .B(\shift[6] ), .ZN(new_n2745_));
  NAND2_X1   g2482(.A1(new_n2744_), .A2(new_n2745_), .ZN(\result[124] ));
  OAI21_X1   g2483(.A1(new_n2529_), .A2(new_n2532_), .B(new_n264_), .ZN(new_n2747_));
  OAI21_X1   g2484(.A1(new_n2523_), .A2(new_n2526_), .B(\shift[6] ), .ZN(new_n2748_));
  NAND2_X1   g2485(.A1(new_n2747_), .A2(new_n2748_), .ZN(\result[125] ));
  OAI21_X1   g2486(.A1(new_n2544_), .A2(new_n2547_), .B(new_n264_), .ZN(new_n2750_));
  OAI21_X1   g2487(.A1(new_n2537_), .A2(new_n2540_), .B(\shift[6] ), .ZN(new_n2751_));
  NAND2_X1   g2488(.A1(new_n2750_), .A2(new_n2751_), .ZN(\result[126] ));
  OAI21_X1   g2489(.A1(new_n2558_), .A2(new_n2561_), .B(new_n264_), .ZN(new_n2753_));
  OAI21_X1   g2490(.A1(new_n2552_), .A2(new_n2555_), .B(\shift[6] ), .ZN(new_n2754_));
  NAND2_X1   g2491(.A1(new_n2753_), .A2(new_n2754_), .ZN(\result[127] ));
endmodule


