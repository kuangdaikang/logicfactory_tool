// Benchmark "example2.blif" written by ABC on Fri Feb 25 15:13:00 2022

module example2  ( 
    a, b, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1,
    j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2,
    b2, c2, d2, e2, f2, g2, h2,
    i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2,
    a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3,
    s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4,
    k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4  );
  input  a, b, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v,
    w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1,
    h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1,
    z1, a2, b2, c2, d2, e2, f2, g2, h2;
  output i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2,
    z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3,
    r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4,
    j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4;
  wire new_n152_, new_n153_, new_n154_, new_n156_, new_n157_, new_n158_,
    new_n160_, new_n161_, new_n162_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n170_, new_n171_, new_n173_, new_n174_,
    new_n176_, new_n177_, new_n179_, new_n180_, new_n182_, new_n183_,
    new_n185_, new_n186_, new_n188_, new_n189_, new_n191_, new_n192_,
    new_n194_, new_n195_, new_n197_, new_n198_, new_n200_, new_n201_,
    new_n203_, new_n204_, new_n206_, new_n207_, new_n209_, new_n210_,
    new_n212_, new_n213_, new_n215_, new_n216_, new_n218_, new_n219_,
    new_n221_, new_n222_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n242_, new_n243_, new_n244_, new_n246_, new_n247_,
    new_n248_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n279_, new_n280_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n336_, new_n337_, new_n338_, new_n339_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n351_, new_n352_, new_n354_, new_n355_, new_n356_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n373_, new_n374_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n412_, new_n413_, new_n416_, new_n417_, new_n418_, new_n419_;
  assign new_n152_ = a2 & b2;
  assign new_n153_ = ~b & c2;
  assign new_n154_ = ~b & ~new_n152_;
  assign m2 = new_n153_ | new_n154_;
  assign new_n156_ = ~b1 & ~m2;
  assign new_n157_ = p0 & ~new_n156_;
  assign new_n158_ = h & ~p0;
  assign i2 = new_n157_ | new_n158_;
  assign new_n160_ = ~a2 & ~b2;
  assign new_n161_ = c2 & ~new_n152_;
  assign new_n162_ = ~new_n160_ & new_n161_;
  assign j2 = ~b & ~new_n162_;
  assign new_n164_ = a2 & ~b2;
  assign new_n165_ = ~a2 & b2;
  assign new_n166_ = p1 & new_n164_;
  assign new_n167_ = y1 & new_n165_;
  assign new_n168_ = ~new_n166_ & ~new_n167_;
  assign k2 = new_n153_ & ~new_n168_;
  assign new_n170_ = b2 & ~c2;
  assign new_n171_ = ~b & b1;
  assign l2 = new_n170_ & new_n171_;
  assign new_n173_ = y & ~p0;
  assign new_n174_ = p0 & o1;
  assign n2 = new_n173_ | new_n174_;
  assign new_n176_ = z & ~p0;
  assign new_n177_ = p0 & n1;
  assign o2 = new_n176_ | new_n177_;
  assign new_n179_ = a0 & ~p0;
  assign new_n180_ = p0 & m1;
  assign p2 = new_n179_ | new_n180_;
  assign new_n182_ = b0 & ~p0;
  assign new_n183_ = p0 & l1;
  assign q2 = new_n182_ | new_n183_;
  assign new_n185_ = c0 & ~p0;
  assign new_n186_ = p0 & k1;
  assign r2 = new_n185_ | new_n186_;
  assign new_n188_ = d0 & ~p0;
  assign new_n189_ = p0 & j1;
  assign s2 = new_n188_ | new_n189_;
  assign new_n191_ = e0 & ~p0;
  assign new_n192_ = p0 & i1;
  assign t2 = new_n191_ | new_n192_;
  assign new_n194_ = f0 & ~p0;
  assign new_n195_ = p0 & h1;
  assign u2 = new_n194_ | new_n195_;
  assign new_n197_ = g0 & ~p0;
  assign new_n198_ = p0 & g1;
  assign v2 = new_n197_ | new_n198_;
  assign new_n200_ = h0 & ~p0;
  assign new_n201_ = p0 & a1;
  assign w2 = new_n200_ | new_n201_;
  assign new_n203_ = i0 & ~p0;
  assign new_n204_ = p0 & z0;
  assign x2 = new_n203_ | new_n204_;
  assign new_n206_ = j0 & ~p0;
  assign new_n207_ = p0 & y0;
  assign y2 = new_n206_ | new_n207_;
  assign new_n209_ = k0 & ~p0;
  assign new_n210_ = p0 & x0;
  assign z2 = new_n209_ | new_n210_;
  assign new_n212_ = l0 & ~p0;
  assign new_n213_ = p0 & w0;
  assign a3 = new_n212_ | new_n213_;
  assign new_n215_ = m0 & ~p0;
  assign new_n216_ = p0 & v0;
  assign b3 = new_n215_ | new_n216_;
  assign new_n218_ = n0 & ~p0;
  assign new_n219_ = p0 & u0;
  assign c3 = new_n218_ | new_n219_;
  assign new_n221_ = o0 & ~p0;
  assign new_n222_ = p0 & t0;
  assign d3 = new_n221_ | new_n222_;
  assign new_n224_ = f & b2;
  assign new_n225_ = f2 & ~g2;
  assign new_n226_ = h2 & new_n225_;
  assign new_n227_ = s0 & ~x1;
  assign new_n228_ = d2 & e2;
  assign new_n229_ = new_n227_ & new_n228_;
  assign new_n230_ = new_n226_ & new_n229_;
  assign new_n231_ = ~r0 & a2;
  assign new_n232_ = ~new_n230_ & new_n231_;
  assign new_n233_ = c2 & ~new_n232_;
  assign new_n234_ = ~b & ~new_n233_;
  assign new_n235_ = new_n224_ & new_n234_;
  assign new_n236_ = e2 & ~h2;
  assign new_n237_ = ~e2 & h2;
  assign new_n238_ = ~new_n236_ & ~new_n237_;
  assign new_n239_ = k2 & new_n238_;
  assign new_n240_ = ~q0 & new_n239_;
  assign e3 = new_n235_ | new_n240_;
  assign new_n242_ = ~f & ~c2;
  assign new_n243_ = g & new_n242_;
  assign new_n244_ = a & ~new_n243_;
  assign f3 = b | ~new_n244_;
  assign new_n246_ = ~s0 & ~new_n161_;
  assign new_n247_ = ~f & new_n246_;
  assign new_n248_ = g & new_n247_;
  assign g3 = ~b & new_n248_;
  assign new_n250_ = ~f & new_n153_;
  assign new_n251_ = new_n152_ & new_n250_;
  assign new_n252_ = ~e2 & ~f2;
  assign new_n253_ = e2 & f2;
  assign new_n254_ = ~new_n252_ & ~new_n253_;
  assign new_n255_ = ~h2 & new_n254_;
  assign new_n256_ = h2 & ~new_n254_;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = ~r0 & ~new_n257_;
  assign new_n259_ = new_n251_ & new_n258_;
  assign h3 = g & new_n259_;
  assign i3 = t0 & new_n259_;
  assign j3 = u0 & new_n259_;
  assign k3 = v0 & new_n259_;
  assign l3 = w0 & new_n259_;
  assign m3 = x0 & new_n259_;
  assign n3 = y0 & new_n259_;
  assign o3 = z0 & new_n259_;
  assign new_n268_ = g2 & ~new_n254_;
  assign new_n269_ = ~g2 & new_n254_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = h2 & new_n270_;
  assign new_n272_ = ~h2 & ~new_n270_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = a1 & new_n259_;
  assign new_n275_ = r0 & ~new_n273_;
  assign new_n276_ = g & new_n251_;
  assign new_n277_ = new_n275_ & new_n276_;
  assign p3 = new_n274_ | new_n277_;
  assign new_n279_ = new_n251_ & new_n275_;
  assign new_n280_ = ~new_n259_ & ~new_n279_;
  assign q3 = b1 & ~new_n280_;
  assign r3 = c1 & ~new_n280_;
  assign s3 = d1 & ~new_n280_;
  assign t3 = e1 & ~new_n280_;
  assign u3 = f1 & ~new_n280_;
  assign v3 = g1 & ~new_n280_;
  assign w3 = h1 & ~new_n280_;
  assign x3 = i1 & ~new_n280_;
  assign y3 = j1 & ~new_n280_;
  assign z3 = k1 & ~new_n280_;
  assign a4 = l1 & ~new_n280_;
  assign b4 = m1 & ~new_n280_;
  assign c4 = n1 & ~new_n280_;
  assign new_n294_ = f & l2;
  assign new_n295_ = ~a2 & new_n294_;
  assign new_n296_ = ~b & ~b1;
  assign new_n297_ = new_n170_ & new_n296_;
  assign new_n298_ = f & new_n297_;
  assign new_n299_ = ~a2 & new_n298_;
  assign new_n300_ = ~g2 & ~h2;
  assign new_n301_ = new_n252_ & new_n300_;
  assign new_n302_ = q0 & p1;
  assign new_n303_ = ~q0 & ~p1;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = d2 & ~new_n304_;
  assign new_n306_ = ~new_n238_ & new_n305_;
  assign new_n307_ = new_n301_ & new_n306_;
  assign new_n308_ = ~q1 & ~y1;
  assign new_n309_ = new_n238_ & ~new_n308_;
  assign new_n310_ = ~new_n307_ & ~new_n309_;
  assign new_n311_ = c2 & ~new_n310_;
  assign new_n312_ = ~b & new_n311_;
  assign new_n313_ = new_n164_ & new_n312_;
  assign new_n314_ = i & new_n299_;
  assign new_n315_ = q & new_n295_;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign d4 = new_n313_ | ~new_n316_;
  assign new_n318_ = ~b & new_n238_;
  assign new_n319_ = c2 & new_n318_;
  assign new_n320_ = new_n164_ & new_n319_;
  assign new_n321_ = r1 & new_n320_;
  assign new_n322_ = r & new_n295_;
  assign new_n323_ = j & new_n299_;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign e4 = new_n321_ | ~new_n324_;
  assign new_n326_ = s1 & new_n320_;
  assign new_n327_ = s & new_n295_;
  assign new_n328_ = k & new_n299_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign f4 = new_n326_ | ~new_n329_;
  assign new_n331_ = t1 & new_n320_;
  assign new_n332_ = t & new_n295_;
  assign new_n333_ = l & new_n299_;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign g4 = new_n331_ | ~new_n334_;
  assign new_n336_ = u1 & new_n320_;
  assign new_n337_ = u & new_n295_;
  assign new_n338_ = m & new_n299_;
  assign new_n339_ = ~new_n337_ & ~new_n338_;
  assign h4 = new_n336_ | ~new_n339_;
  assign new_n341_ = v1 & new_n320_;
  assign new_n342_ = v & new_n295_;
  assign new_n343_ = n & new_n299_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign i4 = new_n341_ | ~new_n344_;
  assign new_n346_ = w1 & new_n320_;
  assign new_n347_ = w & new_n295_;
  assign new_n348_ = o & new_n299_;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign j4 = new_n346_ | ~new_n349_;
  assign new_n351_ = x & new_n295_;
  assign new_n352_ = p & new_n299_;
  assign k4 = new_n351_ | new_n352_;
  assign new_n354_ = ~d2 & g2;
  assign new_n355_ = h2 & new_n354_;
  assign new_n356_ = new_n251_ & new_n355_;
  assign l4 = new_n252_ & new_n356_;
  assign new_n358_ = ~q0 & ~y1;
  assign new_n359_ = q0 & y1;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~a2 & ~new_n360_;
  assign new_n362_ = d2 & new_n301_;
  assign new_n363_ = ~new_n152_ & ~new_n362_;
  assign new_n364_ = ~new_n361_ & ~new_n363_;
  assign new_n365_ = ~new_n238_ & ~new_n364_;
  assign new_n366_ = z1 & new_n238_;
  assign new_n367_ = ~new_n152_ & new_n366_;
  assign new_n368_ = ~new_n365_ & ~new_n367_;
  assign new_n369_ = c2 & ~new_n368_;
  assign new_n370_ = a & ~new_n160_;
  assign new_n371_ = ~b & new_n370_;
  assign m4 = new_n369_ | ~new_n371_;
  assign new_n373_ = a & ~b;
  assign new_n374_ = ~d & new_n373_;
  assign n4 = e & new_n374_;
  assign new_n376_ = ~p0 & r0;
  assign new_n377_ = ~r0 & new_n230_;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = a2 & ~new_n378_;
  assign new_n380_ = new_n153_ & new_n379_;
  assign new_n381_ = new_n224_ & new_n380_;
  assign new_n382_ = ~r0 & new_n164_;
  assign new_n383_ = p0 & new_n382_;
  assign new_n384_ = ~new_n165_ & ~new_n383_;
  assign new_n385_ = f & new_n384_;
  assign new_n386_ = ~c2 & ~new_n385_;
  assign new_n387_ = ~b & new_n386_;
  assign o4 = new_n381_ | new_n387_;
  assign new_n389_ = new_n224_ & new_n232_;
  assign new_n390_ = ~new_n242_ & ~new_n389_;
  assign new_n391_ = c2 & ~new_n224_;
  assign new_n392_ = p0 & ~new_n391_;
  assign new_n393_ = ~new_n170_ & ~new_n392_;
  assign new_n394_ = a2 & ~new_n393_;
  assign new_n395_ = new_n390_ & ~new_n394_;
  assign p4 = ~b & ~new_n395_;
  assign new_n397_ = ~new_n170_ & new_n390_;
  assign new_n398_ = c2 & new_n164_;
  assign new_n399_ = ~new_n165_ & ~new_n398_;
  assign new_n400_ = ~new_n362_ & ~new_n399_;
  assign new_n401_ = ~new_n238_ & new_n400_;
  assign new_n402_ = new_n397_ & ~new_n401_;
  assign q4 = ~b & ~new_n402_;
  assign new_n404_ = ~new_n164_ & ~new_n165_;
  assign new_n405_ = new_n238_ & ~new_n404_;
  assign new_n406_ = ~f & new_n152_;
  assign new_n407_ = ~new_n405_ & ~new_n406_;
  assign new_n408_ = new_n301_ & ~new_n404_;
  assign new_n409_ = new_n407_ & ~new_n408_;
  assign new_n410_ = d2 & ~new_n409_;
  assign r4 = new_n153_ & new_n410_;
  assign new_n412_ = new_n153_ & ~new_n407_;
  assign new_n413_ = e2 & new_n412_;
  assign s4 = new_n235_ | new_n413_;
  assign t4 = f2 & new_n412_;
  assign new_n416_ = g2 & new_n412_;
  assign new_n417_ = ~b & new_n170_;
  assign new_n418_ = f & ~a2;
  assign new_n419_ = new_n417_ & new_n418_;
  assign u4 = new_n416_ | new_n419_;
  assign v4 = h2 & new_n412_;
endmodule


