// Benchmark "testing" written by ABC on Fri Feb 25 15:12:37 2022

module 25_16 ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A43  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A43;
  wire new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_,
    new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_;
  assign new_n27_ = A203 & ~A202;
  assign new_n28_ = A200 & new_n27_;
  assign new_n29_ = ~A203 & A202;
  assign new_n30_ = ~A200 & new_n29_;
  assign new_n31_ = ~new_n28_ & ~new_n30_;
  assign new_n32_ = ~A199 & ~new_n31_;
  assign new_n33_ = A199 & new_n29_;
  assign new_n34_ = ~A201 & ~new_n33_;
  assign new_n35_ = A200 & ~new_n34_;
  assign new_n36_ = ~A200 & new_n27_;
  assign new_n37_ = ~A201 & ~new_n36_;
  assign new_n38_ = A199 & ~new_n37_;
  assign new_n39_ = ~new_n35_ & ~new_n38_;
  assign new_n40_ = ~new_n32_ & new_n39_;
  assign new_n41_ = ~A169 & ~A170;
  assign new_n42_ = A168 & ~new_n41_;
  assign new_n43_ = ~A167 & new_n42_;
  assign new_n44_ = A166 & new_n43_;
  assign new_n45_ = ~A166 & A167;
  assign new_n46_ = ~new_n44_ & ~new_n45_;
  assign new_n47_ = ~new_n40_ & ~new_n46_;
  assign new_n48_ = A166 & new_n42_;
  assign new_n49_ = ~A167 & ~new_n48_;
  assign new_n50_ = A166 & A167;
  assign new_n51_ = ~new_n49_ & ~new_n50_;
  assign new_n52_ = A200 & ~A199;
  assign new_n53_ = ~A200 & A199;
  assign new_n54_ = ~new_n52_ & ~new_n53_;
  assign new_n55_ = ~new_n27_ & ~new_n54_;
  assign new_n56_ = A200 & ~new_n29_;
  assign new_n57_ = A199 & new_n56_;
  assign new_n58_ = ~new_n55_ & ~new_n57_;
  assign new_n59_ = ~new_n51_ & ~new_n58_;
  assign new_n60_ = ~A201 & new_n59_;
  assign new_n61_ = ~new_n29_ & ~new_n51_;
  assign new_n62_ = ~A200 & new_n61_;
  assign new_n63_ = ~A199 & new_n62_;
  assign new_n64_ = A269 & ~A268;
  assign new_n65_ = A266 & new_n64_;
  assign new_n66_ = ~A269 & A268;
  assign new_n67_ = ~A266 & new_n66_;
  assign new_n68_ = ~new_n65_ & ~new_n67_;
  assign new_n69_ = ~A265 & ~new_n68_;
  assign new_n70_ = A265 & new_n66_;
  assign new_n71_ = ~A267 & ~new_n70_;
  assign new_n72_ = A266 & ~new_n71_;
  assign new_n73_ = ~A266 & new_n64_;
  assign new_n74_ = ~A267 & ~new_n73_;
  assign new_n75_ = A265 & ~new_n74_;
  assign new_n76_ = A302 & ~A301;
  assign new_n77_ = A299 & new_n76_;
  assign new_n78_ = ~A302 & A301;
  assign new_n79_ = ~A299 & new_n78_;
  assign new_n80_ = ~new_n77_ & ~new_n79_;
  assign new_n81_ = ~A298 & ~new_n80_;
  assign new_n82_ = A298 & new_n78_;
  assign new_n83_ = ~A300 & ~new_n82_;
  assign new_n84_ = A299 & ~new_n83_;
  assign new_n85_ = ~A299 & new_n76_;
  assign new_n86_ = ~A300 & ~new_n85_;
  assign new_n87_ = A298 & ~new_n86_;
  assign new_n88_ = ~new_n84_ & ~new_n87_;
  assign new_n89_ = ~new_n81_ & new_n88_;
  assign new_n90_ = ~new_n75_ & new_n89_;
  assign new_n91_ = ~new_n72_ & new_n90_;
  assign new_n92_ = ~new_n69_ & new_n91_;
  assign new_n93_ = A236 & ~A235;
  assign new_n94_ = A233 & ~A232;
  assign new_n95_ = ~A233 & A232;
  assign new_n96_ = ~new_n94_ & ~new_n95_;
  assign new_n97_ = ~new_n93_ & ~new_n96_;
  assign new_n98_ = ~A236 & A235;
  assign new_n99_ = A233 & ~new_n98_;
  assign new_n100_ = A232 & new_n99_;
  assign new_n101_ = ~new_n97_ & ~new_n100_;
  assign new_n102_ = ~A234 & ~new_n101_;
  assign new_n103_ = ~A233 & ~new_n98_;
  assign new_n104_ = ~A232 & new_n103_;
  assign new_n105_ = ~new_n102_ & ~new_n104_;
  assign new_n106_ = ~new_n92_ & ~new_n105_;
  assign new_n107_ = A233 & new_n93_;
  assign new_n108_ = ~A233 & new_n98_;
  assign new_n109_ = ~new_n107_ & ~new_n108_;
  assign new_n110_ = ~A232 & ~new_n109_;
  assign new_n111_ = A232 & new_n98_;
  assign new_n112_ = ~A234 & ~new_n111_;
  assign new_n113_ = A233 & ~new_n112_;
  assign new_n114_ = ~A233 & new_n93_;
  assign new_n115_ = ~A234 & ~new_n114_;
  assign new_n116_ = A232 & ~new_n115_;
  assign new_n117_ = ~new_n113_ & ~new_n116_;
  assign new_n118_ = ~new_n110_ & new_n117_;
  assign new_n119_ = A299 & ~A298;
  assign new_n120_ = ~A299 & A298;
  assign new_n121_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = A266 & ~A265;
  assign new_n123_ = ~A266 & A265;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = ~new_n64_ & ~new_n124_;
  assign new_n126_ = A266 & ~new_n66_;
  assign new_n127_ = A265 & new_n126_;
  assign new_n128_ = ~new_n125_ & ~new_n127_;
  assign new_n129_ = ~new_n121_ & ~new_n128_;
  assign new_n130_ = ~new_n76_ & new_n129_;
  assign new_n131_ = ~new_n78_ & ~new_n128_;
  assign new_n132_ = A299 & new_n131_;
  assign new_n133_ = A298 & new_n132_;
  assign new_n134_ = ~new_n130_ & ~new_n133_;
  assign new_n135_ = ~new_n118_ & ~new_n134_;
  assign new_n136_ = ~A267 & new_n135_;
  assign new_n137_ = ~new_n76_ & ~new_n121_;
  assign new_n138_ = A299 & ~new_n78_;
  assign new_n139_ = A298 & new_n138_;
  assign new_n140_ = ~new_n137_ & ~new_n139_;
  assign new_n141_ = ~new_n118_ & ~new_n140_;
  assign new_n142_ = ~new_n66_ & new_n141_;
  assign new_n143_ = ~A266 & new_n142_;
  assign new_n144_ = ~A265 & new_n143_;
  assign new_n145_ = ~new_n136_ & ~new_n144_;
  assign new_n146_ = ~A300 & ~new_n145_;
  assign new_n147_ = ~new_n118_ & ~new_n128_;
  assign new_n148_ = ~A267 & new_n147_;
  assign new_n149_ = ~new_n66_ & ~new_n118_;
  assign new_n150_ = ~A266 & new_n149_;
  assign new_n151_ = ~A265 & new_n150_;
  assign new_n152_ = ~new_n148_ & ~new_n151_;
  assign new_n153_ = ~new_n78_ & ~new_n152_;
  assign new_n154_ = ~A299 & new_n153_;
  assign new_n155_ = ~A298 & new_n154_;
  assign new_n156_ = ~new_n146_ & ~new_n155_;
  assign new_n157_ = ~new_n106_ & new_n156_;
  assign new_n158_ = ~new_n63_ & new_n157_;
  assign new_n159_ = ~new_n60_ & new_n158_;
  assign A43 = ~new_n47_ & new_n159_;
endmodule


