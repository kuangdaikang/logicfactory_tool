// Benchmark "top" written by ABC on Fri Sep 15 19:21:45 2023

module top ( 
    n_1, n_2, n_3, n_4,
     );
  input  n_1, n_2, n_3, n_4;
  output;
endmodule


