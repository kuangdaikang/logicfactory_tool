// Benchmark "priority" written by ABC on Fri Sep 15 11:27:16 2023

module priority ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1037_,
    new_n1038_, new_n1039_;
  INV_X1     g000(.I(\A[4] ), .ZN(new_n137_));
  INV_X1     g001(.I(\A[12] ), .ZN(new_n138_));
  INV_X1     g002(.I(\A[16] ), .ZN(new_n139_));
  INV_X1     g003(.I(\A[20] ), .ZN(new_n140_));
  INV_X1     g004(.I(\A[24] ), .ZN(new_n141_));
  INV_X1     g005(.I(\A[28] ), .ZN(new_n142_));
  INV_X1     g006(.I(\A[32] ), .ZN(new_n143_));
  INV_X1     g007(.I(\A[36] ), .ZN(new_n144_));
  INV_X1     g008(.I(\A[40] ), .ZN(new_n145_));
  INV_X1     g009(.I(\A[44] ), .ZN(new_n146_));
  INV_X1     g010(.I(\A[48] ), .ZN(new_n147_));
  INV_X1     g011(.I(\A[52] ), .ZN(new_n148_));
  INV_X1     g012(.I(\A[56] ), .ZN(new_n149_));
  INV_X1     g013(.I(\A[60] ), .ZN(new_n150_));
  INV_X1     g014(.I(\A[64] ), .ZN(new_n151_));
  INV_X1     g015(.I(\A[68] ), .ZN(new_n152_));
  INV_X1     g016(.I(\A[72] ), .ZN(new_n153_));
  INV_X1     g017(.I(\A[76] ), .ZN(new_n154_));
  INV_X1     g018(.I(\A[80] ), .ZN(new_n155_));
  INV_X1     g019(.I(\A[84] ), .ZN(new_n156_));
  INV_X1     g020(.I(\A[88] ), .ZN(new_n157_));
  INV_X1     g021(.I(\A[92] ), .ZN(new_n158_));
  INV_X1     g022(.I(\A[96] ), .ZN(new_n159_));
  INV_X1     g023(.I(\A[100] ), .ZN(new_n160_));
  INV_X1     g024(.I(\A[104] ), .ZN(new_n161_));
  INV_X1     g025(.I(\A[108] ), .ZN(new_n162_));
  INV_X1     g026(.I(\A[112] ), .ZN(new_n163_));
  INV_X1     g027(.I(\A[116] ), .ZN(new_n164_));
  INV_X1     g028(.I(\A[125] ), .ZN(new_n165_));
  AOI21_X1   g029(.A1(new_n165_), .A2(\A[124] ), .B(\A[126] ), .ZN(new_n166_));
  INV_X1     g030(.I(\A[122] ), .ZN(new_n167_));
  NOR2_X1    g031(.A1(new_n167_), .A2(\A[123] ), .ZN(new_n168_));
  NOR3_X1    g032(.A1(new_n166_), .A2(new_n168_), .A3(\A[127] ), .ZN(new_n169_));
  NOR2_X1    g033(.A1(new_n165_), .A2(\A[126] ), .ZN(new_n170_));
  NOR4_X1    g034(.A1(new_n170_), .A2(new_n167_), .A3(\A[123] ), .A4(\A[127] ), .ZN(new_n171_));
  INV_X1     g035(.I(\A[120] ), .ZN(new_n172_));
  NOR2_X1    g036(.A1(new_n172_), .A2(\A[121] ), .ZN(new_n173_));
  INV_X1     g037(.I(new_n173_), .ZN(new_n174_));
  OAI21_X1   g038(.A1(new_n171_), .A2(new_n169_), .B(new_n174_), .ZN(new_n175_));
  NOR3_X1    g039(.A1(new_n170_), .A2(\A[123] ), .A3(\A[127] ), .ZN(new_n176_));
  INV_X1     g040(.I(\A[123] ), .ZN(new_n177_));
  NOR3_X1    g041(.A1(new_n166_), .A2(new_n177_), .A3(\A[127] ), .ZN(new_n178_));
  OAI21_X1   g042(.A1(new_n178_), .A2(new_n176_), .B(new_n173_), .ZN(new_n179_));
  INV_X1     g043(.I(\A[119] ), .ZN(new_n180_));
  NAND2_X1   g044(.A1(new_n180_), .A2(\A[118] ), .ZN(new_n181_));
  INV_X1     g045(.I(new_n181_), .ZN(new_n182_));
  AOI21_X1   g046(.A1(new_n175_), .A2(new_n179_), .B(new_n182_), .ZN(new_n183_));
  INV_X1     g047(.I(\A[121] ), .ZN(new_n184_));
  OAI21_X1   g048(.A1(new_n178_), .A2(new_n176_), .B(new_n184_), .ZN(new_n185_));
  OAI21_X1   g049(.A1(new_n171_), .A2(new_n169_), .B(\A[121] ), .ZN(new_n186_));
  AOI21_X1   g050(.A1(new_n186_), .A2(new_n185_), .B(new_n181_), .ZN(new_n187_));
  OAI22_X1   g051(.A1(new_n183_), .A2(new_n187_), .B1(new_n164_), .B2(\A[117] ), .ZN(new_n188_));
  NOR2_X1    g052(.A1(new_n164_), .A2(\A[117] ), .ZN(new_n189_));
  AOI21_X1   g053(.A1(new_n186_), .A2(new_n185_), .B(\A[119] ), .ZN(new_n190_));
  AOI21_X1   g054(.A1(new_n175_), .A2(new_n179_), .B(new_n180_), .ZN(new_n191_));
  OAI21_X1   g055(.A1(new_n190_), .A2(new_n191_), .B(new_n189_), .ZN(new_n192_));
  INV_X1     g056(.I(\A[114] ), .ZN(new_n193_));
  NOR2_X1    g057(.A1(new_n193_), .A2(\A[115] ), .ZN(new_n194_));
  AOI21_X1   g058(.A1(new_n188_), .A2(new_n192_), .B(new_n194_), .ZN(new_n195_));
  INV_X1     g059(.I(new_n194_), .ZN(new_n196_));
  INV_X1     g060(.I(\A[117] ), .ZN(new_n197_));
  OAI21_X1   g061(.A1(new_n190_), .A2(new_n191_), .B(new_n197_), .ZN(new_n198_));
  OAI21_X1   g062(.A1(new_n183_), .A2(new_n187_), .B(\A[117] ), .ZN(new_n199_));
  AOI21_X1   g063(.A1(new_n198_), .A2(new_n199_), .B(new_n196_), .ZN(new_n200_));
  OAI22_X1   g064(.A1(new_n195_), .A2(new_n200_), .B1(new_n163_), .B2(\A[113] ), .ZN(new_n201_));
  NOR2_X1    g065(.A1(new_n163_), .A2(\A[113] ), .ZN(new_n202_));
  AOI21_X1   g066(.A1(new_n198_), .A2(new_n199_), .B(\A[115] ), .ZN(new_n203_));
  INV_X1     g067(.I(\A[115] ), .ZN(new_n204_));
  AOI21_X1   g068(.A1(new_n188_), .A2(new_n192_), .B(new_n204_), .ZN(new_n205_));
  OAI21_X1   g069(.A1(new_n205_), .A2(new_n203_), .B(new_n202_), .ZN(new_n206_));
  INV_X1     g070(.I(\A[110] ), .ZN(new_n207_));
  NOR2_X1    g071(.A1(new_n207_), .A2(\A[111] ), .ZN(new_n208_));
  AOI21_X1   g072(.A1(new_n201_), .A2(new_n206_), .B(new_n208_), .ZN(new_n209_));
  INV_X1     g073(.I(new_n208_), .ZN(new_n210_));
  INV_X1     g074(.I(\A[113] ), .ZN(new_n211_));
  OAI21_X1   g075(.A1(new_n205_), .A2(new_n203_), .B(new_n211_), .ZN(new_n212_));
  OAI21_X1   g076(.A1(new_n195_), .A2(new_n200_), .B(\A[113] ), .ZN(new_n213_));
  AOI21_X1   g077(.A1(new_n212_), .A2(new_n213_), .B(new_n210_), .ZN(new_n214_));
  OAI22_X1   g078(.A1(new_n209_), .A2(new_n214_), .B1(new_n162_), .B2(\A[109] ), .ZN(new_n215_));
  NOR2_X1    g079(.A1(new_n162_), .A2(\A[109] ), .ZN(new_n216_));
  AOI21_X1   g080(.A1(new_n212_), .A2(new_n213_), .B(\A[111] ), .ZN(new_n217_));
  INV_X1     g081(.I(\A[111] ), .ZN(new_n218_));
  AOI21_X1   g082(.A1(new_n201_), .A2(new_n206_), .B(new_n218_), .ZN(new_n219_));
  OAI21_X1   g083(.A1(new_n219_), .A2(new_n217_), .B(new_n216_), .ZN(new_n220_));
  INV_X1     g084(.I(\A[106] ), .ZN(new_n221_));
  NOR2_X1    g085(.A1(new_n221_), .A2(\A[107] ), .ZN(new_n222_));
  AOI21_X1   g086(.A1(new_n215_), .A2(new_n220_), .B(new_n222_), .ZN(new_n223_));
  INV_X1     g087(.I(new_n222_), .ZN(new_n224_));
  INV_X1     g088(.I(\A[109] ), .ZN(new_n225_));
  OAI21_X1   g089(.A1(new_n219_), .A2(new_n217_), .B(new_n225_), .ZN(new_n226_));
  OAI21_X1   g090(.A1(new_n209_), .A2(new_n214_), .B(\A[109] ), .ZN(new_n227_));
  AOI21_X1   g091(.A1(new_n226_), .A2(new_n227_), .B(new_n224_), .ZN(new_n228_));
  OAI22_X1   g092(.A1(new_n223_), .A2(new_n228_), .B1(new_n161_), .B2(\A[105] ), .ZN(new_n229_));
  NOR2_X1    g093(.A1(new_n161_), .A2(\A[105] ), .ZN(new_n230_));
  AOI21_X1   g094(.A1(new_n226_), .A2(new_n227_), .B(\A[107] ), .ZN(new_n231_));
  INV_X1     g095(.I(\A[107] ), .ZN(new_n232_));
  AOI21_X1   g096(.A1(new_n215_), .A2(new_n220_), .B(new_n232_), .ZN(new_n233_));
  OAI21_X1   g097(.A1(new_n233_), .A2(new_n231_), .B(new_n230_), .ZN(new_n234_));
  INV_X1     g098(.I(\A[102] ), .ZN(new_n235_));
  NOR2_X1    g099(.A1(new_n235_), .A2(\A[103] ), .ZN(new_n236_));
  AOI21_X1   g100(.A1(new_n229_), .A2(new_n234_), .B(new_n236_), .ZN(new_n237_));
  INV_X1     g101(.I(new_n236_), .ZN(new_n238_));
  INV_X1     g102(.I(\A[105] ), .ZN(new_n239_));
  OAI21_X1   g103(.A1(new_n233_), .A2(new_n231_), .B(new_n239_), .ZN(new_n240_));
  OAI21_X1   g104(.A1(new_n223_), .A2(new_n228_), .B(\A[105] ), .ZN(new_n241_));
  AOI21_X1   g105(.A1(new_n240_), .A2(new_n241_), .B(new_n238_), .ZN(new_n242_));
  OAI22_X1   g106(.A1(new_n237_), .A2(new_n242_), .B1(new_n160_), .B2(\A[101] ), .ZN(new_n243_));
  NOR2_X1    g107(.A1(new_n160_), .A2(\A[101] ), .ZN(new_n244_));
  AOI21_X1   g108(.A1(new_n240_), .A2(new_n241_), .B(\A[103] ), .ZN(new_n245_));
  INV_X1     g109(.I(\A[103] ), .ZN(new_n246_));
  AOI21_X1   g110(.A1(new_n229_), .A2(new_n234_), .B(new_n246_), .ZN(new_n247_));
  OAI21_X1   g111(.A1(new_n247_), .A2(new_n245_), .B(new_n244_), .ZN(new_n248_));
  INV_X1     g112(.I(\A[98] ), .ZN(new_n249_));
  NOR2_X1    g113(.A1(new_n249_), .A2(\A[99] ), .ZN(new_n250_));
  AOI21_X1   g114(.A1(new_n243_), .A2(new_n248_), .B(new_n250_), .ZN(new_n251_));
  INV_X1     g115(.I(new_n250_), .ZN(new_n252_));
  INV_X1     g116(.I(\A[101] ), .ZN(new_n253_));
  OAI21_X1   g117(.A1(new_n247_), .A2(new_n245_), .B(new_n253_), .ZN(new_n254_));
  OAI21_X1   g118(.A1(new_n237_), .A2(new_n242_), .B(\A[101] ), .ZN(new_n255_));
  AOI21_X1   g119(.A1(new_n254_), .A2(new_n255_), .B(new_n252_), .ZN(new_n256_));
  OAI22_X1   g120(.A1(new_n251_), .A2(new_n256_), .B1(new_n159_), .B2(\A[97] ), .ZN(new_n257_));
  NOR2_X1    g121(.A1(new_n159_), .A2(\A[97] ), .ZN(new_n258_));
  AOI21_X1   g122(.A1(new_n254_), .A2(new_n255_), .B(\A[99] ), .ZN(new_n259_));
  INV_X1     g123(.I(\A[99] ), .ZN(new_n260_));
  AOI21_X1   g124(.A1(new_n243_), .A2(new_n248_), .B(new_n260_), .ZN(new_n261_));
  OAI21_X1   g125(.A1(new_n261_), .A2(new_n259_), .B(new_n258_), .ZN(new_n262_));
  INV_X1     g126(.I(\A[94] ), .ZN(new_n263_));
  NOR2_X1    g127(.A1(new_n263_), .A2(\A[95] ), .ZN(new_n264_));
  AOI21_X1   g128(.A1(new_n257_), .A2(new_n262_), .B(new_n264_), .ZN(new_n265_));
  INV_X1     g129(.I(new_n264_), .ZN(new_n266_));
  INV_X1     g130(.I(\A[97] ), .ZN(new_n267_));
  OAI21_X1   g131(.A1(new_n261_), .A2(new_n259_), .B(new_n267_), .ZN(new_n268_));
  OAI21_X1   g132(.A1(new_n251_), .A2(new_n256_), .B(\A[97] ), .ZN(new_n269_));
  AOI21_X1   g133(.A1(new_n268_), .A2(new_n269_), .B(new_n266_), .ZN(new_n270_));
  OAI22_X1   g134(.A1(new_n265_), .A2(new_n270_), .B1(new_n158_), .B2(\A[93] ), .ZN(new_n271_));
  NOR2_X1    g135(.A1(new_n158_), .A2(\A[93] ), .ZN(new_n272_));
  AOI21_X1   g136(.A1(new_n268_), .A2(new_n269_), .B(\A[95] ), .ZN(new_n273_));
  INV_X1     g137(.I(\A[95] ), .ZN(new_n274_));
  AOI21_X1   g138(.A1(new_n257_), .A2(new_n262_), .B(new_n274_), .ZN(new_n275_));
  OAI21_X1   g139(.A1(new_n275_), .A2(new_n273_), .B(new_n272_), .ZN(new_n276_));
  INV_X1     g140(.I(\A[90] ), .ZN(new_n277_));
  NOR2_X1    g141(.A1(new_n277_), .A2(\A[91] ), .ZN(new_n278_));
  AOI21_X1   g142(.A1(new_n271_), .A2(new_n276_), .B(new_n278_), .ZN(new_n279_));
  INV_X1     g143(.I(new_n278_), .ZN(new_n280_));
  INV_X1     g144(.I(\A[93] ), .ZN(new_n281_));
  OAI21_X1   g145(.A1(new_n275_), .A2(new_n273_), .B(new_n281_), .ZN(new_n282_));
  OAI21_X1   g146(.A1(new_n265_), .A2(new_n270_), .B(\A[93] ), .ZN(new_n283_));
  AOI21_X1   g147(.A1(new_n282_), .A2(new_n283_), .B(new_n280_), .ZN(new_n284_));
  OAI22_X1   g148(.A1(new_n279_), .A2(new_n284_), .B1(new_n157_), .B2(\A[89] ), .ZN(new_n285_));
  NOR2_X1    g149(.A1(new_n157_), .A2(\A[89] ), .ZN(new_n286_));
  AOI21_X1   g150(.A1(new_n282_), .A2(new_n283_), .B(\A[91] ), .ZN(new_n287_));
  INV_X1     g151(.I(\A[91] ), .ZN(new_n288_));
  AOI21_X1   g152(.A1(new_n271_), .A2(new_n276_), .B(new_n288_), .ZN(new_n289_));
  OAI21_X1   g153(.A1(new_n289_), .A2(new_n287_), .B(new_n286_), .ZN(new_n290_));
  INV_X1     g154(.I(\A[86] ), .ZN(new_n291_));
  NOR2_X1    g155(.A1(new_n291_), .A2(\A[87] ), .ZN(new_n292_));
  AOI21_X1   g156(.A1(new_n285_), .A2(new_n290_), .B(new_n292_), .ZN(new_n293_));
  INV_X1     g157(.I(new_n292_), .ZN(new_n294_));
  INV_X1     g158(.I(\A[89] ), .ZN(new_n295_));
  OAI21_X1   g159(.A1(new_n289_), .A2(new_n287_), .B(new_n295_), .ZN(new_n296_));
  OAI21_X1   g160(.A1(new_n279_), .A2(new_n284_), .B(\A[89] ), .ZN(new_n297_));
  AOI21_X1   g161(.A1(new_n296_), .A2(new_n297_), .B(new_n294_), .ZN(new_n298_));
  OAI22_X1   g162(.A1(new_n293_), .A2(new_n298_), .B1(new_n156_), .B2(\A[85] ), .ZN(new_n299_));
  NOR2_X1    g163(.A1(new_n156_), .A2(\A[85] ), .ZN(new_n300_));
  AOI21_X1   g164(.A1(new_n296_), .A2(new_n297_), .B(\A[87] ), .ZN(new_n301_));
  INV_X1     g165(.I(\A[87] ), .ZN(new_n302_));
  AOI21_X1   g166(.A1(new_n285_), .A2(new_n290_), .B(new_n302_), .ZN(new_n303_));
  OAI21_X1   g167(.A1(new_n303_), .A2(new_n301_), .B(new_n300_), .ZN(new_n304_));
  INV_X1     g168(.I(\A[82] ), .ZN(new_n305_));
  NOR2_X1    g169(.A1(new_n305_), .A2(\A[83] ), .ZN(new_n306_));
  AOI21_X1   g170(.A1(new_n299_), .A2(new_n304_), .B(new_n306_), .ZN(new_n307_));
  INV_X1     g171(.I(new_n306_), .ZN(new_n308_));
  INV_X1     g172(.I(\A[85] ), .ZN(new_n309_));
  OAI21_X1   g173(.A1(new_n303_), .A2(new_n301_), .B(new_n309_), .ZN(new_n310_));
  OAI21_X1   g174(.A1(new_n293_), .A2(new_n298_), .B(\A[85] ), .ZN(new_n311_));
  AOI21_X1   g175(.A1(new_n310_), .A2(new_n311_), .B(new_n308_), .ZN(new_n312_));
  OAI22_X1   g176(.A1(new_n307_), .A2(new_n312_), .B1(new_n155_), .B2(\A[81] ), .ZN(new_n313_));
  NOR2_X1    g177(.A1(new_n155_), .A2(\A[81] ), .ZN(new_n314_));
  AOI21_X1   g178(.A1(new_n310_), .A2(new_n311_), .B(\A[83] ), .ZN(new_n315_));
  INV_X1     g179(.I(\A[83] ), .ZN(new_n316_));
  AOI21_X1   g180(.A1(new_n299_), .A2(new_n304_), .B(new_n316_), .ZN(new_n317_));
  OAI21_X1   g181(.A1(new_n317_), .A2(new_n315_), .B(new_n314_), .ZN(new_n318_));
  INV_X1     g182(.I(\A[78] ), .ZN(new_n319_));
  NOR2_X1    g183(.A1(new_n319_), .A2(\A[79] ), .ZN(new_n320_));
  AOI21_X1   g184(.A1(new_n313_), .A2(new_n318_), .B(new_n320_), .ZN(new_n321_));
  INV_X1     g185(.I(new_n320_), .ZN(new_n322_));
  INV_X1     g186(.I(\A[81] ), .ZN(new_n323_));
  OAI21_X1   g187(.A1(new_n317_), .A2(new_n315_), .B(new_n323_), .ZN(new_n324_));
  OAI21_X1   g188(.A1(new_n307_), .A2(new_n312_), .B(\A[81] ), .ZN(new_n325_));
  AOI21_X1   g189(.A1(new_n324_), .A2(new_n325_), .B(new_n322_), .ZN(new_n326_));
  OAI22_X1   g190(.A1(new_n321_), .A2(new_n326_), .B1(new_n154_), .B2(\A[77] ), .ZN(new_n327_));
  NOR2_X1    g191(.A1(new_n154_), .A2(\A[77] ), .ZN(new_n328_));
  AOI21_X1   g192(.A1(new_n324_), .A2(new_n325_), .B(\A[79] ), .ZN(new_n329_));
  INV_X1     g193(.I(\A[79] ), .ZN(new_n330_));
  AOI21_X1   g194(.A1(new_n313_), .A2(new_n318_), .B(new_n330_), .ZN(new_n331_));
  OAI21_X1   g195(.A1(new_n331_), .A2(new_n329_), .B(new_n328_), .ZN(new_n332_));
  INV_X1     g196(.I(\A[74] ), .ZN(new_n333_));
  NOR2_X1    g197(.A1(new_n333_), .A2(\A[75] ), .ZN(new_n334_));
  AOI21_X1   g198(.A1(new_n327_), .A2(new_n332_), .B(new_n334_), .ZN(new_n335_));
  INV_X1     g199(.I(new_n334_), .ZN(new_n336_));
  INV_X1     g200(.I(\A[77] ), .ZN(new_n337_));
  OAI21_X1   g201(.A1(new_n331_), .A2(new_n329_), .B(new_n337_), .ZN(new_n338_));
  OAI21_X1   g202(.A1(new_n321_), .A2(new_n326_), .B(\A[77] ), .ZN(new_n339_));
  AOI21_X1   g203(.A1(new_n338_), .A2(new_n339_), .B(new_n336_), .ZN(new_n340_));
  OAI22_X1   g204(.A1(new_n335_), .A2(new_n340_), .B1(new_n153_), .B2(\A[73] ), .ZN(new_n341_));
  NOR2_X1    g205(.A1(new_n153_), .A2(\A[73] ), .ZN(new_n342_));
  AOI21_X1   g206(.A1(new_n338_), .A2(new_n339_), .B(\A[75] ), .ZN(new_n343_));
  INV_X1     g207(.I(\A[75] ), .ZN(new_n344_));
  AOI21_X1   g208(.A1(new_n327_), .A2(new_n332_), .B(new_n344_), .ZN(new_n345_));
  OAI21_X1   g209(.A1(new_n345_), .A2(new_n343_), .B(new_n342_), .ZN(new_n346_));
  INV_X1     g210(.I(\A[70] ), .ZN(new_n347_));
  NOR2_X1    g211(.A1(new_n347_), .A2(\A[71] ), .ZN(new_n348_));
  AOI21_X1   g212(.A1(new_n341_), .A2(new_n346_), .B(new_n348_), .ZN(new_n349_));
  INV_X1     g213(.I(new_n348_), .ZN(new_n350_));
  INV_X1     g214(.I(\A[73] ), .ZN(new_n351_));
  OAI21_X1   g215(.A1(new_n345_), .A2(new_n343_), .B(new_n351_), .ZN(new_n352_));
  OAI21_X1   g216(.A1(new_n335_), .A2(new_n340_), .B(\A[73] ), .ZN(new_n353_));
  AOI21_X1   g217(.A1(new_n352_), .A2(new_n353_), .B(new_n350_), .ZN(new_n354_));
  OAI22_X1   g218(.A1(new_n349_), .A2(new_n354_), .B1(new_n152_), .B2(\A[69] ), .ZN(new_n355_));
  NOR2_X1    g219(.A1(new_n152_), .A2(\A[69] ), .ZN(new_n356_));
  AOI21_X1   g220(.A1(new_n352_), .A2(new_n353_), .B(\A[71] ), .ZN(new_n357_));
  INV_X1     g221(.I(\A[71] ), .ZN(new_n358_));
  AOI21_X1   g222(.A1(new_n341_), .A2(new_n346_), .B(new_n358_), .ZN(new_n359_));
  OAI21_X1   g223(.A1(new_n359_), .A2(new_n357_), .B(new_n356_), .ZN(new_n360_));
  INV_X1     g224(.I(\A[66] ), .ZN(new_n361_));
  NOR2_X1    g225(.A1(new_n361_), .A2(\A[67] ), .ZN(new_n362_));
  AOI21_X1   g226(.A1(new_n355_), .A2(new_n360_), .B(new_n362_), .ZN(new_n363_));
  INV_X1     g227(.I(new_n362_), .ZN(new_n364_));
  INV_X1     g228(.I(\A[69] ), .ZN(new_n365_));
  OAI21_X1   g229(.A1(new_n359_), .A2(new_n357_), .B(new_n365_), .ZN(new_n366_));
  OAI21_X1   g230(.A1(new_n349_), .A2(new_n354_), .B(\A[69] ), .ZN(new_n367_));
  AOI21_X1   g231(.A1(new_n366_), .A2(new_n367_), .B(new_n364_), .ZN(new_n368_));
  OAI22_X1   g232(.A1(new_n363_), .A2(new_n368_), .B1(new_n151_), .B2(\A[65] ), .ZN(new_n369_));
  NOR2_X1    g233(.A1(new_n151_), .A2(\A[65] ), .ZN(new_n370_));
  AOI21_X1   g234(.A1(new_n366_), .A2(new_n367_), .B(\A[67] ), .ZN(new_n371_));
  INV_X1     g235(.I(\A[67] ), .ZN(new_n372_));
  AOI21_X1   g236(.A1(new_n355_), .A2(new_n360_), .B(new_n372_), .ZN(new_n373_));
  OAI21_X1   g237(.A1(new_n373_), .A2(new_n371_), .B(new_n370_), .ZN(new_n374_));
  INV_X1     g238(.I(\A[62] ), .ZN(new_n375_));
  NOR2_X1    g239(.A1(new_n375_), .A2(\A[63] ), .ZN(new_n376_));
  AOI21_X1   g240(.A1(new_n369_), .A2(new_n374_), .B(new_n376_), .ZN(new_n377_));
  INV_X1     g241(.I(new_n376_), .ZN(new_n378_));
  INV_X1     g242(.I(\A[65] ), .ZN(new_n379_));
  OAI21_X1   g243(.A1(new_n373_), .A2(new_n371_), .B(new_n379_), .ZN(new_n380_));
  OAI21_X1   g244(.A1(new_n363_), .A2(new_n368_), .B(\A[65] ), .ZN(new_n381_));
  AOI21_X1   g245(.A1(new_n380_), .A2(new_n381_), .B(new_n378_), .ZN(new_n382_));
  OAI22_X1   g246(.A1(new_n377_), .A2(new_n382_), .B1(new_n150_), .B2(\A[61] ), .ZN(new_n383_));
  NOR2_X1    g247(.A1(new_n150_), .A2(\A[61] ), .ZN(new_n384_));
  AOI21_X1   g248(.A1(new_n380_), .A2(new_n381_), .B(\A[63] ), .ZN(new_n385_));
  INV_X1     g249(.I(\A[63] ), .ZN(new_n386_));
  AOI21_X1   g250(.A1(new_n369_), .A2(new_n374_), .B(new_n386_), .ZN(new_n387_));
  OAI21_X1   g251(.A1(new_n387_), .A2(new_n385_), .B(new_n384_), .ZN(new_n388_));
  INV_X1     g252(.I(\A[58] ), .ZN(new_n389_));
  NOR2_X1    g253(.A1(new_n389_), .A2(\A[59] ), .ZN(new_n390_));
  AOI21_X1   g254(.A1(new_n383_), .A2(new_n388_), .B(new_n390_), .ZN(new_n391_));
  INV_X1     g255(.I(new_n390_), .ZN(new_n392_));
  INV_X1     g256(.I(\A[61] ), .ZN(new_n393_));
  OAI21_X1   g257(.A1(new_n387_), .A2(new_n385_), .B(new_n393_), .ZN(new_n394_));
  OAI21_X1   g258(.A1(new_n377_), .A2(new_n382_), .B(\A[61] ), .ZN(new_n395_));
  AOI21_X1   g259(.A1(new_n394_), .A2(new_n395_), .B(new_n392_), .ZN(new_n396_));
  OAI22_X1   g260(.A1(new_n391_), .A2(new_n396_), .B1(new_n149_), .B2(\A[57] ), .ZN(new_n397_));
  NOR2_X1    g261(.A1(new_n149_), .A2(\A[57] ), .ZN(new_n398_));
  AOI21_X1   g262(.A1(new_n394_), .A2(new_n395_), .B(\A[59] ), .ZN(new_n399_));
  INV_X1     g263(.I(\A[59] ), .ZN(new_n400_));
  AOI21_X1   g264(.A1(new_n383_), .A2(new_n388_), .B(new_n400_), .ZN(new_n401_));
  OAI21_X1   g265(.A1(new_n401_), .A2(new_n399_), .B(new_n398_), .ZN(new_n402_));
  INV_X1     g266(.I(\A[54] ), .ZN(new_n403_));
  NOR2_X1    g267(.A1(new_n403_), .A2(\A[55] ), .ZN(new_n404_));
  AOI21_X1   g268(.A1(new_n397_), .A2(new_n402_), .B(new_n404_), .ZN(new_n405_));
  INV_X1     g269(.I(new_n404_), .ZN(new_n406_));
  INV_X1     g270(.I(\A[57] ), .ZN(new_n407_));
  OAI21_X1   g271(.A1(new_n401_), .A2(new_n399_), .B(new_n407_), .ZN(new_n408_));
  OAI21_X1   g272(.A1(new_n391_), .A2(new_n396_), .B(\A[57] ), .ZN(new_n409_));
  AOI21_X1   g273(.A1(new_n408_), .A2(new_n409_), .B(new_n406_), .ZN(new_n410_));
  OAI22_X1   g274(.A1(new_n405_), .A2(new_n410_), .B1(new_n148_), .B2(\A[53] ), .ZN(new_n411_));
  NOR2_X1    g275(.A1(new_n148_), .A2(\A[53] ), .ZN(new_n412_));
  AOI21_X1   g276(.A1(new_n408_), .A2(new_n409_), .B(\A[55] ), .ZN(new_n413_));
  INV_X1     g277(.I(\A[55] ), .ZN(new_n414_));
  AOI21_X1   g278(.A1(new_n397_), .A2(new_n402_), .B(new_n414_), .ZN(new_n415_));
  OAI21_X1   g279(.A1(new_n415_), .A2(new_n413_), .B(new_n412_), .ZN(new_n416_));
  INV_X1     g280(.I(\A[50] ), .ZN(new_n417_));
  NOR2_X1    g281(.A1(new_n417_), .A2(\A[51] ), .ZN(new_n418_));
  AOI21_X1   g282(.A1(new_n411_), .A2(new_n416_), .B(new_n418_), .ZN(new_n419_));
  INV_X1     g283(.I(new_n418_), .ZN(new_n420_));
  INV_X1     g284(.I(\A[53] ), .ZN(new_n421_));
  OAI21_X1   g285(.A1(new_n415_), .A2(new_n413_), .B(new_n421_), .ZN(new_n422_));
  OAI21_X1   g286(.A1(new_n405_), .A2(new_n410_), .B(\A[53] ), .ZN(new_n423_));
  AOI21_X1   g287(.A1(new_n422_), .A2(new_n423_), .B(new_n420_), .ZN(new_n424_));
  OAI22_X1   g288(.A1(new_n419_), .A2(new_n424_), .B1(new_n147_), .B2(\A[49] ), .ZN(new_n425_));
  NOR2_X1    g289(.A1(new_n147_), .A2(\A[49] ), .ZN(new_n426_));
  AOI21_X1   g290(.A1(new_n422_), .A2(new_n423_), .B(\A[51] ), .ZN(new_n427_));
  INV_X1     g291(.I(\A[51] ), .ZN(new_n428_));
  AOI21_X1   g292(.A1(new_n411_), .A2(new_n416_), .B(new_n428_), .ZN(new_n429_));
  OAI21_X1   g293(.A1(new_n429_), .A2(new_n427_), .B(new_n426_), .ZN(new_n430_));
  INV_X1     g294(.I(\A[46] ), .ZN(new_n431_));
  NOR2_X1    g295(.A1(new_n431_), .A2(\A[47] ), .ZN(new_n432_));
  AOI21_X1   g296(.A1(new_n425_), .A2(new_n430_), .B(new_n432_), .ZN(new_n433_));
  INV_X1     g297(.I(new_n432_), .ZN(new_n434_));
  INV_X1     g298(.I(\A[49] ), .ZN(new_n435_));
  OAI21_X1   g299(.A1(new_n429_), .A2(new_n427_), .B(new_n435_), .ZN(new_n436_));
  OAI21_X1   g300(.A1(new_n419_), .A2(new_n424_), .B(\A[49] ), .ZN(new_n437_));
  AOI21_X1   g301(.A1(new_n436_), .A2(new_n437_), .B(new_n434_), .ZN(new_n438_));
  OAI22_X1   g302(.A1(new_n433_), .A2(new_n438_), .B1(new_n146_), .B2(\A[45] ), .ZN(new_n439_));
  NOR2_X1    g303(.A1(new_n146_), .A2(\A[45] ), .ZN(new_n440_));
  AOI21_X1   g304(.A1(new_n436_), .A2(new_n437_), .B(\A[47] ), .ZN(new_n441_));
  INV_X1     g305(.I(\A[47] ), .ZN(new_n442_));
  AOI21_X1   g306(.A1(new_n425_), .A2(new_n430_), .B(new_n442_), .ZN(new_n443_));
  OAI21_X1   g307(.A1(new_n443_), .A2(new_n441_), .B(new_n440_), .ZN(new_n444_));
  INV_X1     g308(.I(\A[42] ), .ZN(new_n445_));
  NOR2_X1    g309(.A1(new_n445_), .A2(\A[43] ), .ZN(new_n446_));
  AOI21_X1   g310(.A1(new_n439_), .A2(new_n444_), .B(new_n446_), .ZN(new_n447_));
  INV_X1     g311(.I(new_n446_), .ZN(new_n448_));
  INV_X1     g312(.I(\A[45] ), .ZN(new_n449_));
  OAI21_X1   g313(.A1(new_n443_), .A2(new_n441_), .B(new_n449_), .ZN(new_n450_));
  OAI21_X1   g314(.A1(new_n433_), .A2(new_n438_), .B(\A[45] ), .ZN(new_n451_));
  AOI21_X1   g315(.A1(new_n450_), .A2(new_n451_), .B(new_n448_), .ZN(new_n452_));
  OAI22_X1   g316(.A1(new_n447_), .A2(new_n452_), .B1(new_n145_), .B2(\A[41] ), .ZN(new_n453_));
  NOR2_X1    g317(.A1(new_n145_), .A2(\A[41] ), .ZN(new_n454_));
  AOI21_X1   g318(.A1(new_n450_), .A2(new_n451_), .B(\A[43] ), .ZN(new_n455_));
  INV_X1     g319(.I(\A[43] ), .ZN(new_n456_));
  AOI21_X1   g320(.A1(new_n439_), .A2(new_n444_), .B(new_n456_), .ZN(new_n457_));
  OAI21_X1   g321(.A1(new_n457_), .A2(new_n455_), .B(new_n454_), .ZN(new_n458_));
  INV_X1     g322(.I(\A[38] ), .ZN(new_n459_));
  NOR2_X1    g323(.A1(new_n459_), .A2(\A[39] ), .ZN(new_n460_));
  AOI21_X1   g324(.A1(new_n453_), .A2(new_n458_), .B(new_n460_), .ZN(new_n461_));
  INV_X1     g325(.I(new_n460_), .ZN(new_n462_));
  INV_X1     g326(.I(\A[41] ), .ZN(new_n463_));
  OAI21_X1   g327(.A1(new_n457_), .A2(new_n455_), .B(new_n463_), .ZN(new_n464_));
  OAI21_X1   g328(.A1(new_n447_), .A2(new_n452_), .B(\A[41] ), .ZN(new_n465_));
  AOI21_X1   g329(.A1(new_n464_), .A2(new_n465_), .B(new_n462_), .ZN(new_n466_));
  OAI22_X1   g330(.A1(new_n461_), .A2(new_n466_), .B1(new_n144_), .B2(\A[37] ), .ZN(new_n467_));
  NOR2_X1    g331(.A1(new_n144_), .A2(\A[37] ), .ZN(new_n468_));
  AOI21_X1   g332(.A1(new_n464_), .A2(new_n465_), .B(\A[39] ), .ZN(new_n469_));
  INV_X1     g333(.I(\A[39] ), .ZN(new_n470_));
  AOI21_X1   g334(.A1(new_n453_), .A2(new_n458_), .B(new_n470_), .ZN(new_n471_));
  OAI21_X1   g335(.A1(new_n471_), .A2(new_n469_), .B(new_n468_), .ZN(new_n472_));
  INV_X1     g336(.I(\A[34] ), .ZN(new_n473_));
  NOR2_X1    g337(.A1(new_n473_), .A2(\A[35] ), .ZN(new_n474_));
  AOI21_X1   g338(.A1(new_n467_), .A2(new_n472_), .B(new_n474_), .ZN(new_n475_));
  INV_X1     g339(.I(new_n474_), .ZN(new_n476_));
  INV_X1     g340(.I(\A[37] ), .ZN(new_n477_));
  OAI21_X1   g341(.A1(new_n471_), .A2(new_n469_), .B(new_n477_), .ZN(new_n478_));
  OAI21_X1   g342(.A1(new_n461_), .A2(new_n466_), .B(\A[37] ), .ZN(new_n479_));
  AOI21_X1   g343(.A1(new_n478_), .A2(new_n479_), .B(new_n476_), .ZN(new_n480_));
  OAI22_X1   g344(.A1(new_n475_), .A2(new_n480_), .B1(new_n143_), .B2(\A[33] ), .ZN(new_n481_));
  NOR2_X1    g345(.A1(new_n143_), .A2(\A[33] ), .ZN(new_n482_));
  AOI21_X1   g346(.A1(new_n478_), .A2(new_n479_), .B(\A[35] ), .ZN(new_n483_));
  INV_X1     g347(.I(\A[35] ), .ZN(new_n484_));
  AOI21_X1   g348(.A1(new_n467_), .A2(new_n472_), .B(new_n484_), .ZN(new_n485_));
  OAI21_X1   g349(.A1(new_n485_), .A2(new_n483_), .B(new_n482_), .ZN(new_n486_));
  INV_X1     g350(.I(\A[30] ), .ZN(new_n487_));
  NOR2_X1    g351(.A1(new_n487_), .A2(\A[31] ), .ZN(new_n488_));
  AOI21_X1   g352(.A1(new_n481_), .A2(new_n486_), .B(new_n488_), .ZN(new_n489_));
  INV_X1     g353(.I(new_n488_), .ZN(new_n490_));
  INV_X1     g354(.I(\A[33] ), .ZN(new_n491_));
  OAI21_X1   g355(.A1(new_n485_), .A2(new_n483_), .B(new_n491_), .ZN(new_n492_));
  OAI21_X1   g356(.A1(new_n475_), .A2(new_n480_), .B(\A[33] ), .ZN(new_n493_));
  AOI21_X1   g357(.A1(new_n492_), .A2(new_n493_), .B(new_n490_), .ZN(new_n494_));
  OAI22_X1   g358(.A1(new_n489_), .A2(new_n494_), .B1(new_n142_), .B2(\A[29] ), .ZN(new_n495_));
  NOR2_X1    g359(.A1(new_n142_), .A2(\A[29] ), .ZN(new_n496_));
  AOI21_X1   g360(.A1(new_n492_), .A2(new_n493_), .B(\A[31] ), .ZN(new_n497_));
  INV_X1     g361(.I(\A[31] ), .ZN(new_n498_));
  AOI21_X1   g362(.A1(new_n481_), .A2(new_n486_), .B(new_n498_), .ZN(new_n499_));
  OAI21_X1   g363(.A1(new_n499_), .A2(new_n497_), .B(new_n496_), .ZN(new_n500_));
  INV_X1     g364(.I(\A[26] ), .ZN(new_n501_));
  NOR2_X1    g365(.A1(new_n501_), .A2(\A[27] ), .ZN(new_n502_));
  AOI21_X1   g366(.A1(new_n495_), .A2(new_n500_), .B(new_n502_), .ZN(new_n503_));
  INV_X1     g367(.I(new_n502_), .ZN(new_n504_));
  INV_X1     g368(.I(\A[29] ), .ZN(new_n505_));
  OAI21_X1   g369(.A1(new_n499_), .A2(new_n497_), .B(new_n505_), .ZN(new_n506_));
  OAI21_X1   g370(.A1(new_n489_), .A2(new_n494_), .B(\A[29] ), .ZN(new_n507_));
  AOI21_X1   g371(.A1(new_n506_), .A2(new_n507_), .B(new_n504_), .ZN(new_n508_));
  OAI22_X1   g372(.A1(new_n503_), .A2(new_n508_), .B1(new_n141_), .B2(\A[25] ), .ZN(new_n509_));
  NOR2_X1    g373(.A1(new_n141_), .A2(\A[25] ), .ZN(new_n510_));
  AOI21_X1   g374(.A1(new_n506_), .A2(new_n507_), .B(\A[27] ), .ZN(new_n511_));
  INV_X1     g375(.I(\A[27] ), .ZN(new_n512_));
  AOI21_X1   g376(.A1(new_n495_), .A2(new_n500_), .B(new_n512_), .ZN(new_n513_));
  OAI21_X1   g377(.A1(new_n513_), .A2(new_n511_), .B(new_n510_), .ZN(new_n514_));
  INV_X1     g378(.I(\A[22] ), .ZN(new_n515_));
  NOR2_X1    g379(.A1(new_n515_), .A2(\A[23] ), .ZN(new_n516_));
  AOI21_X1   g380(.A1(new_n509_), .A2(new_n514_), .B(new_n516_), .ZN(new_n517_));
  INV_X1     g381(.I(new_n516_), .ZN(new_n518_));
  INV_X1     g382(.I(\A[25] ), .ZN(new_n519_));
  OAI21_X1   g383(.A1(new_n513_), .A2(new_n511_), .B(new_n519_), .ZN(new_n520_));
  OAI21_X1   g384(.A1(new_n503_), .A2(new_n508_), .B(\A[25] ), .ZN(new_n521_));
  AOI21_X1   g385(.A1(new_n520_), .A2(new_n521_), .B(new_n518_), .ZN(new_n522_));
  OAI22_X1   g386(.A1(new_n517_), .A2(new_n522_), .B1(new_n140_), .B2(\A[21] ), .ZN(new_n523_));
  NOR2_X1    g387(.A1(new_n140_), .A2(\A[21] ), .ZN(new_n524_));
  AOI21_X1   g388(.A1(new_n520_), .A2(new_n521_), .B(\A[23] ), .ZN(new_n525_));
  INV_X1     g389(.I(\A[23] ), .ZN(new_n526_));
  AOI21_X1   g390(.A1(new_n509_), .A2(new_n514_), .B(new_n526_), .ZN(new_n527_));
  OAI21_X1   g391(.A1(new_n527_), .A2(new_n525_), .B(new_n524_), .ZN(new_n528_));
  INV_X1     g392(.I(\A[18] ), .ZN(new_n529_));
  NOR2_X1    g393(.A1(new_n529_), .A2(\A[19] ), .ZN(new_n530_));
  AOI21_X1   g394(.A1(new_n523_), .A2(new_n528_), .B(new_n530_), .ZN(new_n531_));
  INV_X1     g395(.I(new_n530_), .ZN(new_n532_));
  INV_X1     g396(.I(\A[21] ), .ZN(new_n533_));
  OAI21_X1   g397(.A1(new_n527_), .A2(new_n525_), .B(new_n533_), .ZN(new_n534_));
  OAI21_X1   g398(.A1(new_n517_), .A2(new_n522_), .B(\A[21] ), .ZN(new_n535_));
  AOI21_X1   g399(.A1(new_n534_), .A2(new_n535_), .B(new_n532_), .ZN(new_n536_));
  OAI22_X1   g400(.A1(new_n531_), .A2(new_n536_), .B1(new_n139_), .B2(\A[17] ), .ZN(new_n537_));
  NOR2_X1    g401(.A1(new_n139_), .A2(\A[17] ), .ZN(new_n538_));
  AOI21_X1   g402(.A1(new_n534_), .A2(new_n535_), .B(\A[19] ), .ZN(new_n539_));
  INV_X1     g403(.I(\A[19] ), .ZN(new_n540_));
  AOI21_X1   g404(.A1(new_n523_), .A2(new_n528_), .B(new_n540_), .ZN(new_n541_));
  OAI21_X1   g405(.A1(new_n541_), .A2(new_n539_), .B(new_n538_), .ZN(new_n542_));
  INV_X1     g406(.I(\A[14] ), .ZN(new_n543_));
  NOR2_X1    g407(.A1(new_n543_), .A2(\A[15] ), .ZN(new_n544_));
  AOI21_X1   g408(.A1(new_n537_), .A2(new_n542_), .B(new_n544_), .ZN(new_n545_));
  INV_X1     g409(.I(new_n544_), .ZN(new_n546_));
  INV_X1     g410(.I(\A[17] ), .ZN(new_n547_));
  OAI21_X1   g411(.A1(new_n541_), .A2(new_n539_), .B(new_n547_), .ZN(new_n548_));
  OAI21_X1   g412(.A1(new_n531_), .A2(new_n536_), .B(\A[17] ), .ZN(new_n549_));
  AOI21_X1   g413(.A1(new_n548_), .A2(new_n549_), .B(new_n546_), .ZN(new_n550_));
  OAI22_X1   g414(.A1(new_n545_), .A2(new_n550_), .B1(new_n138_), .B2(\A[13] ), .ZN(new_n551_));
  NOR2_X1    g415(.A1(new_n138_), .A2(\A[13] ), .ZN(new_n552_));
  AOI21_X1   g416(.A1(new_n548_), .A2(new_n549_), .B(\A[15] ), .ZN(new_n553_));
  INV_X1     g417(.I(\A[15] ), .ZN(new_n554_));
  AOI21_X1   g418(.A1(new_n537_), .A2(new_n542_), .B(new_n554_), .ZN(new_n555_));
  OAI21_X1   g419(.A1(new_n555_), .A2(new_n553_), .B(new_n552_), .ZN(new_n556_));
  INV_X1     g420(.I(\A[10] ), .ZN(new_n557_));
  NOR2_X1    g421(.A1(new_n557_), .A2(\A[11] ), .ZN(new_n558_));
  AOI21_X1   g422(.A1(new_n551_), .A2(new_n556_), .B(new_n558_), .ZN(new_n559_));
  INV_X1     g423(.I(new_n558_), .ZN(new_n560_));
  INV_X1     g424(.I(\A[13] ), .ZN(new_n561_));
  OAI21_X1   g425(.A1(new_n555_), .A2(new_n553_), .B(new_n561_), .ZN(new_n562_));
  OAI21_X1   g426(.A1(new_n545_), .A2(new_n550_), .B(\A[13] ), .ZN(new_n563_));
  AOI21_X1   g427(.A1(new_n562_), .A2(new_n563_), .B(new_n560_), .ZN(new_n564_));
  INV_X1     g428(.I(\A[9] ), .ZN(new_n565_));
  NAND2_X1   g429(.A1(new_n565_), .A2(\A[8] ), .ZN(new_n566_));
  OAI21_X1   g430(.A1(new_n559_), .A2(new_n564_), .B(new_n566_), .ZN(new_n567_));
  INV_X1     g431(.I(new_n566_), .ZN(new_n568_));
  AOI21_X1   g432(.A1(new_n562_), .A2(new_n563_), .B(\A[11] ), .ZN(new_n569_));
  INV_X1     g433(.I(\A[11] ), .ZN(new_n570_));
  AOI21_X1   g434(.A1(new_n551_), .A2(new_n556_), .B(new_n570_), .ZN(new_n571_));
  OAI21_X1   g435(.A1(new_n571_), .A2(new_n569_), .B(new_n568_), .ZN(new_n572_));
  INV_X1     g436(.I(\A[6] ), .ZN(new_n573_));
  NOR2_X1    g437(.A1(new_n573_), .A2(\A[7] ), .ZN(new_n574_));
  AOI21_X1   g438(.A1(new_n567_), .A2(new_n572_), .B(new_n574_), .ZN(new_n575_));
  INV_X1     g439(.I(new_n574_), .ZN(new_n576_));
  OAI21_X1   g440(.A1(new_n571_), .A2(new_n569_), .B(new_n565_), .ZN(new_n577_));
  OAI21_X1   g441(.A1(new_n559_), .A2(new_n564_), .B(\A[9] ), .ZN(new_n578_));
  AOI21_X1   g442(.A1(new_n577_), .A2(new_n578_), .B(new_n576_), .ZN(new_n579_));
  OAI22_X1   g443(.A1(new_n575_), .A2(new_n579_), .B1(new_n137_), .B2(\A[5] ), .ZN(new_n580_));
  NOR2_X1    g444(.A1(new_n137_), .A2(\A[5] ), .ZN(new_n581_));
  AOI21_X1   g445(.A1(new_n577_), .A2(new_n578_), .B(\A[7] ), .ZN(new_n582_));
  INV_X1     g446(.I(\A[7] ), .ZN(new_n583_));
  AOI21_X1   g447(.A1(new_n567_), .A2(new_n572_), .B(new_n583_), .ZN(new_n584_));
  OAI21_X1   g448(.A1(new_n582_), .A2(new_n584_), .B(new_n581_), .ZN(new_n585_));
  INV_X1     g449(.I(\A[2] ), .ZN(new_n586_));
  AOI21_X1   g450(.A1(new_n586_), .A2(\A[1] ), .B(\A[3] ), .ZN(new_n587_));
  INV_X1     g451(.I(new_n587_), .ZN(new_n588_));
  NAND3_X1   g452(.A1(new_n580_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1     g453(.I(\A[5] ), .ZN(new_n590_));
  OAI21_X1   g454(.A1(new_n582_), .A2(new_n584_), .B(new_n590_), .ZN(new_n591_));
  OAI21_X1   g455(.A1(new_n575_), .A2(new_n579_), .B(\A[5] ), .ZN(new_n592_));
  NAND3_X1   g456(.A1(new_n591_), .A2(new_n592_), .A3(new_n587_), .ZN(new_n593_));
  NAND2_X1   g457(.A1(new_n589_), .A2(new_n593_), .ZN(\P[0] ));
  NOR2_X1    g458(.A1(\A[10] ), .A2(\A[11] ), .ZN(new_n595_));
  NOR2_X1    g459(.A1(\A[102] ), .A2(\A[103] ), .ZN(new_n596_));
  NOR2_X1    g460(.A1(\A[126] ), .A2(\A[127] ), .ZN(new_n597_));
  NOR2_X1    g461(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n598_));
  OR2_X2     g462(.A1(\A[124] ), .A2(\A[125] ), .Z(new_n599_));
  OAI21_X1   g463(.A1(new_n599_), .A2(new_n598_), .B(new_n597_), .ZN(new_n600_));
  NOR2_X1    g464(.A1(new_n600_), .A2(new_n172_), .ZN(new_n601_));
  INV_X1     g465(.I(new_n599_), .ZN(new_n602_));
  NAND2_X1   g466(.A1(new_n597_), .A2(new_n172_), .ZN(new_n603_));
  NAND2_X1   g467(.A1(new_n598_), .A2(\A[121] ), .ZN(new_n604_));
  AOI21_X1   g468(.A1(new_n602_), .A2(new_n604_), .B(new_n603_), .ZN(new_n605_));
  OR2_X2     g469(.A1(new_n601_), .A2(new_n605_), .Z(new_n606_));
  NOR2_X1    g470(.A1(\A[118] ), .A2(\A[119] ), .ZN(new_n607_));
  NAND2_X1   g471(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1   g472(.A1(new_n606_), .A2(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1    g473(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n610_));
  NOR2_X1    g474(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X2    g475(.A1(new_n606_), .A2(new_n610_), .Z(new_n612_));
  OR2_X2     g476(.A1(new_n611_), .A2(new_n612_), .Z(new_n613_));
  NOR2_X1    g477(.A1(\A[114] ), .A2(\A[115] ), .ZN(new_n614_));
  NAND2_X1   g478(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1   g479(.A1(new_n613_), .A2(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1    g480(.A1(\A[112] ), .A2(\A[113] ), .ZN(new_n617_));
  NOR2_X1    g481(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X2    g482(.A1(new_n613_), .A2(new_n617_), .Z(new_n619_));
  OR2_X2     g483(.A1(new_n618_), .A2(new_n619_), .Z(new_n620_));
  NOR2_X1    g484(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n621_));
  NAND2_X1   g485(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1   g486(.A1(new_n620_), .A2(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NOR2_X1    g487(.A1(\A[108] ), .A2(\A[109] ), .ZN(new_n624_));
  NOR2_X1    g488(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X2    g489(.A1(new_n620_), .A2(new_n624_), .Z(new_n626_));
  NOR2_X1    g490(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1    g491(.A1(\A[106] ), .A2(\A[107] ), .ZN(new_n628_));
  INV_X1     g492(.I(new_n628_), .ZN(new_n629_));
  NAND2_X1   g493(.A1(new_n623_), .A2(new_n628_), .ZN(new_n630_));
  INV_X1     g494(.I(new_n630_), .ZN(new_n631_));
  AOI21_X1   g495(.A1(new_n627_), .A2(new_n629_), .B(new_n631_), .ZN(new_n632_));
  NOR3_X1    g496(.A1(new_n632_), .A2(\A[102] ), .A3(\A[103] ), .ZN(new_n633_));
  INV_X1     g497(.I(new_n633_), .ZN(new_n634_));
  NOR2_X1    g498(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n635_));
  INV_X1     g499(.I(new_n635_), .ZN(new_n636_));
  NAND2_X1   g500(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1   g501(.A1(new_n627_), .A2(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OAI21_X1   g502(.A1(new_n638_), .A2(new_n596_), .B(new_n634_), .ZN(new_n639_));
  NOR2_X1    g503(.A1(\A[100] ), .A2(\A[101] ), .ZN(new_n640_));
  NOR2_X1    g504(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X2    g505(.A1(new_n638_), .A2(new_n640_), .Z(new_n642_));
  NOR2_X1    g506(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1     g507(.I(new_n643_), .ZN(new_n644_));
  NOR2_X1    g508(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n645_));
  NAND2_X1   g509(.A1(new_n639_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1   g510(.A1(new_n644_), .A2(new_n645_), .B(new_n646_), .ZN(new_n647_));
  NOR2_X1    g511(.A1(\A[96] ), .A2(\A[97] ), .ZN(new_n648_));
  NOR2_X1    g512(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1    g513(.A1(new_n643_), .A2(\A[96] ), .A3(\A[97] ), .ZN(new_n650_));
  NOR2_X1    g514(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1     g515(.I(new_n651_), .ZN(new_n652_));
  NOR2_X1    g516(.A1(\A[94] ), .A2(\A[95] ), .ZN(new_n653_));
  NAND2_X1   g517(.A1(new_n647_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1   g518(.A1(new_n652_), .A2(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NOR2_X1    g519(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n656_));
  NAND2_X1   g520(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1   g521(.A1(new_n655_), .A2(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NOR2_X1    g522(.A1(\A[90] ), .A2(\A[91] ), .ZN(new_n659_));
  NAND2_X1   g523(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1   g524(.A1(new_n658_), .A2(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NOR2_X1    g525(.A1(\A[88] ), .A2(\A[89] ), .ZN(new_n662_));
  NOR2_X1    g526(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND2_X2    g527(.A1(new_n658_), .A2(new_n662_), .Z(new_n664_));
  NOR2_X1    g528(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n665_));
  OR3_X2     g529(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .Z(new_n666_));
  NAND2_X1   g530(.A1(new_n661_), .A2(new_n665_), .ZN(new_n667_));
  NAND2_X1   g531(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1    g532(.A1(\A[84] ), .A2(\A[85] ), .ZN(new_n669_));
  OR2_X2     g533(.A1(new_n668_), .A2(new_n669_), .Z(new_n670_));
  OAI21_X1   g534(.A1(new_n663_), .A2(new_n664_), .B(new_n669_), .ZN(new_n671_));
  NOR2_X1    g535(.A1(\A[82] ), .A2(\A[83] ), .ZN(new_n672_));
  INV_X1     g536(.I(new_n672_), .ZN(new_n673_));
  NAND3_X1   g537(.A1(new_n670_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1   g538(.A1(new_n668_), .A2(new_n672_), .ZN(new_n675_));
  NOR2_X1    g539(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n676_));
  INV_X1     g540(.I(new_n676_), .ZN(new_n677_));
  NAND3_X1   g541(.A1(new_n674_), .A2(new_n675_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1   g542(.A1(new_n670_), .A2(new_n671_), .ZN(new_n679_));
  NAND2_X1   g543(.A1(new_n679_), .A2(new_n676_), .ZN(new_n680_));
  NAND2_X1   g544(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1    g545(.A1(\A[76] ), .A2(\A[77] ), .ZN(new_n682_));
  NAND2_X1   g546(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1     g547(.I(new_n682_), .ZN(new_n684_));
  NAND2_X1   g548(.A1(new_n674_), .A2(new_n675_), .ZN(new_n685_));
  NOR2_X1    g549(.A1(\A[78] ), .A2(\A[79] ), .ZN(new_n686_));
  NAND2_X1   g550(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1     g551(.I(new_n686_), .ZN(new_n688_));
  NAND3_X1   g552(.A1(new_n678_), .A2(new_n680_), .A3(new_n688_), .ZN(new_n689_));
  NAND3_X1   g553(.A1(new_n689_), .A2(new_n684_), .A3(new_n687_), .ZN(new_n690_));
  NOR2_X1    g554(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n691_));
  INV_X1     g555(.I(new_n691_), .ZN(new_n692_));
  NAND3_X1   g556(.A1(new_n690_), .A2(new_n683_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1   g557(.A1(new_n689_), .A2(new_n687_), .ZN(new_n694_));
  NAND2_X1   g558(.A1(new_n694_), .A2(new_n691_), .ZN(new_n695_));
  NOR2_X1    g559(.A1(\A[72] ), .A2(\A[73] ), .ZN(new_n696_));
  INV_X1     g560(.I(new_n696_), .ZN(new_n697_));
  NAND3_X1   g561(.A1(new_n693_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1   g562(.A1(new_n690_), .A2(new_n683_), .ZN(new_n699_));
  NAND2_X1   g563(.A1(new_n699_), .A2(new_n696_), .ZN(new_n700_));
  NOR2_X1    g564(.A1(\A[70] ), .A2(\A[71] ), .ZN(new_n701_));
  INV_X1     g565(.I(new_n701_), .ZN(new_n702_));
  NAND3_X1   g566(.A1(new_n698_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1   g567(.A1(new_n693_), .A2(new_n695_), .ZN(new_n704_));
  NAND2_X1   g568(.A1(new_n704_), .A2(new_n701_), .ZN(new_n705_));
  NOR2_X1    g569(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n706_));
  INV_X1     g570(.I(new_n706_), .ZN(new_n707_));
  NAND3_X1   g571(.A1(new_n703_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1   g572(.A1(new_n698_), .A2(new_n700_), .ZN(new_n709_));
  NAND2_X1   g573(.A1(new_n709_), .A2(new_n706_), .ZN(new_n710_));
  NOR2_X1    g574(.A1(\A[66] ), .A2(\A[67] ), .ZN(new_n711_));
  INV_X1     g575(.I(new_n711_), .ZN(new_n712_));
  NAND3_X1   g576(.A1(new_n708_), .A2(new_n710_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1   g577(.A1(new_n703_), .A2(new_n705_), .ZN(new_n714_));
  NAND2_X1   g578(.A1(new_n714_), .A2(new_n711_), .ZN(new_n715_));
  NOR2_X1    g579(.A1(\A[64] ), .A2(\A[65] ), .ZN(new_n716_));
  INV_X1     g580(.I(new_n716_), .ZN(new_n717_));
  NAND3_X1   g581(.A1(new_n713_), .A2(new_n715_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1   g582(.A1(new_n708_), .A2(new_n710_), .ZN(new_n719_));
  NAND2_X1   g583(.A1(new_n719_), .A2(new_n716_), .ZN(new_n720_));
  NOR2_X1    g584(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n721_));
  INV_X1     g585(.I(new_n721_), .ZN(new_n722_));
  NAND3_X1   g586(.A1(new_n718_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1   g587(.A1(new_n713_), .A2(new_n715_), .ZN(new_n724_));
  NAND2_X1   g588(.A1(new_n724_), .A2(new_n721_), .ZN(new_n725_));
  NOR2_X1    g589(.A1(\A[60] ), .A2(\A[61] ), .ZN(new_n726_));
  INV_X1     g590(.I(new_n726_), .ZN(new_n727_));
  NAND3_X1   g591(.A1(new_n723_), .A2(new_n725_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1   g592(.A1(new_n718_), .A2(new_n720_), .ZN(new_n729_));
  NAND2_X1   g593(.A1(new_n729_), .A2(new_n726_), .ZN(new_n730_));
  NOR2_X1    g594(.A1(\A[58] ), .A2(\A[59] ), .ZN(new_n731_));
  INV_X1     g595(.I(new_n731_), .ZN(new_n732_));
  NAND3_X1   g596(.A1(new_n728_), .A2(new_n730_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1   g597(.A1(new_n723_), .A2(new_n725_), .ZN(new_n734_));
  NAND2_X1   g598(.A1(new_n734_), .A2(new_n731_), .ZN(new_n735_));
  NOR2_X1    g599(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n736_));
  INV_X1     g600(.I(new_n736_), .ZN(new_n737_));
  NAND3_X1   g601(.A1(new_n733_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1   g602(.A1(new_n728_), .A2(new_n730_), .ZN(new_n739_));
  NAND2_X1   g603(.A1(new_n739_), .A2(new_n736_), .ZN(new_n740_));
  NOR2_X1    g604(.A1(\A[54] ), .A2(\A[55] ), .ZN(new_n741_));
  INV_X1     g605(.I(new_n741_), .ZN(new_n742_));
  NAND3_X1   g606(.A1(new_n738_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1   g607(.A1(new_n733_), .A2(new_n735_), .ZN(new_n744_));
  NAND2_X1   g608(.A1(new_n744_), .A2(new_n741_), .ZN(new_n745_));
  NOR2_X1    g609(.A1(\A[52] ), .A2(\A[53] ), .ZN(new_n746_));
  INV_X1     g610(.I(new_n746_), .ZN(new_n747_));
  NAND3_X1   g611(.A1(new_n743_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1   g612(.A1(new_n738_), .A2(new_n740_), .ZN(new_n749_));
  NAND2_X1   g613(.A1(new_n749_), .A2(new_n746_), .ZN(new_n750_));
  NOR2_X1    g614(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n751_));
  INV_X1     g615(.I(new_n751_), .ZN(new_n752_));
  NAND3_X1   g616(.A1(new_n748_), .A2(new_n750_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1   g617(.A1(new_n743_), .A2(new_n745_), .ZN(new_n754_));
  NAND2_X1   g618(.A1(new_n754_), .A2(new_n751_), .ZN(new_n755_));
  NOR2_X1    g619(.A1(\A[48] ), .A2(\A[49] ), .ZN(new_n756_));
  INV_X1     g620(.I(new_n756_), .ZN(new_n757_));
  NAND3_X1   g621(.A1(new_n753_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1   g622(.A1(new_n748_), .A2(new_n750_), .ZN(new_n759_));
  NAND2_X1   g623(.A1(new_n759_), .A2(new_n756_), .ZN(new_n760_));
  NOR2_X1    g624(.A1(\A[46] ), .A2(\A[47] ), .ZN(new_n761_));
  INV_X1     g625(.I(new_n761_), .ZN(new_n762_));
  NAND3_X1   g626(.A1(new_n758_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1   g627(.A1(new_n753_), .A2(new_n755_), .ZN(new_n764_));
  NAND2_X1   g628(.A1(new_n764_), .A2(new_n761_), .ZN(new_n765_));
  NOR2_X1    g629(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n766_));
  INV_X1     g630(.I(new_n766_), .ZN(new_n767_));
  NAND3_X1   g631(.A1(new_n763_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1   g632(.A1(new_n758_), .A2(new_n760_), .ZN(new_n769_));
  NAND2_X1   g633(.A1(new_n769_), .A2(new_n766_), .ZN(new_n770_));
  NOR2_X1    g634(.A1(\A[42] ), .A2(\A[43] ), .ZN(new_n771_));
  INV_X1     g635(.I(new_n771_), .ZN(new_n772_));
  NAND3_X1   g636(.A1(new_n768_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1   g637(.A1(new_n763_), .A2(new_n765_), .ZN(new_n774_));
  NAND2_X1   g638(.A1(new_n774_), .A2(new_n771_), .ZN(new_n775_));
  NOR2_X1    g639(.A1(\A[40] ), .A2(\A[41] ), .ZN(new_n776_));
  INV_X1     g640(.I(new_n776_), .ZN(new_n777_));
  NAND3_X1   g641(.A1(new_n773_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1   g642(.A1(new_n768_), .A2(new_n770_), .ZN(new_n779_));
  NAND2_X1   g643(.A1(new_n779_), .A2(new_n776_), .ZN(new_n780_));
  NOR2_X1    g644(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n781_));
  INV_X1     g645(.I(new_n781_), .ZN(new_n782_));
  NAND3_X1   g646(.A1(new_n778_), .A2(new_n780_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1   g647(.A1(new_n773_), .A2(new_n775_), .ZN(new_n784_));
  NAND2_X1   g648(.A1(new_n784_), .A2(new_n781_), .ZN(new_n785_));
  NOR2_X1    g649(.A1(\A[36] ), .A2(\A[37] ), .ZN(new_n786_));
  INV_X1     g650(.I(new_n786_), .ZN(new_n787_));
  NAND3_X1   g651(.A1(new_n783_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1   g652(.A1(new_n778_), .A2(new_n780_), .ZN(new_n789_));
  NAND2_X1   g653(.A1(new_n789_), .A2(new_n786_), .ZN(new_n790_));
  NOR2_X1    g654(.A1(\A[34] ), .A2(\A[35] ), .ZN(new_n791_));
  INV_X1     g655(.I(new_n791_), .ZN(new_n792_));
  NAND3_X1   g656(.A1(new_n788_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1   g657(.A1(new_n783_), .A2(new_n785_), .ZN(new_n794_));
  NAND2_X1   g658(.A1(new_n794_), .A2(new_n791_), .ZN(new_n795_));
  NOR2_X1    g659(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n796_));
  INV_X1     g660(.I(new_n796_), .ZN(new_n797_));
  NAND3_X1   g661(.A1(new_n793_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1   g662(.A1(new_n788_), .A2(new_n790_), .ZN(new_n799_));
  NAND2_X1   g663(.A1(new_n799_), .A2(new_n796_), .ZN(new_n800_));
  NAND2_X1   g664(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1    g665(.A1(\A[30] ), .A2(\A[31] ), .ZN(new_n802_));
  OR2_X2     g666(.A1(new_n801_), .A2(new_n802_), .Z(new_n803_));
  NAND2_X1   g667(.A1(new_n793_), .A2(new_n795_), .ZN(new_n804_));
  NAND2_X1   g668(.A1(new_n804_), .A2(new_n802_), .ZN(new_n805_));
  NOR2_X1    g669(.A1(\A[28] ), .A2(\A[29] ), .ZN(new_n806_));
  INV_X1     g670(.I(new_n806_), .ZN(new_n807_));
  NAND3_X1   g671(.A1(new_n803_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1   g672(.A1(new_n801_), .A2(new_n806_), .ZN(new_n809_));
  NOR2_X1    g673(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n810_));
  INV_X1     g674(.I(new_n810_), .ZN(new_n811_));
  NAND3_X1   g675(.A1(new_n808_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1   g676(.A1(new_n803_), .A2(new_n805_), .ZN(new_n813_));
  NAND2_X1   g677(.A1(new_n813_), .A2(new_n810_), .ZN(new_n814_));
  NOR2_X1    g678(.A1(\A[24] ), .A2(\A[25] ), .ZN(new_n815_));
  INV_X1     g679(.I(new_n815_), .ZN(new_n816_));
  NAND3_X1   g680(.A1(new_n812_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1   g681(.A1(new_n808_), .A2(new_n809_), .ZN(new_n818_));
  NAND2_X1   g682(.A1(new_n818_), .A2(new_n815_), .ZN(new_n819_));
  NOR2_X1    g683(.A1(\A[22] ), .A2(\A[23] ), .ZN(new_n820_));
  INV_X1     g684(.I(new_n820_), .ZN(new_n821_));
  NAND3_X1   g685(.A1(new_n817_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1   g686(.A1(new_n812_), .A2(new_n814_), .ZN(new_n823_));
  NAND2_X1   g687(.A1(new_n823_), .A2(new_n820_), .ZN(new_n824_));
  NOR2_X1    g688(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n825_));
  INV_X1     g689(.I(new_n825_), .ZN(new_n826_));
  NAND3_X1   g690(.A1(new_n822_), .A2(new_n824_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1   g691(.A1(new_n817_), .A2(new_n819_), .ZN(new_n828_));
  NAND2_X1   g692(.A1(new_n828_), .A2(new_n825_), .ZN(new_n829_));
  NOR2_X1    g693(.A1(\A[18] ), .A2(\A[19] ), .ZN(new_n830_));
  INV_X1     g694(.I(new_n830_), .ZN(new_n831_));
  NAND3_X1   g695(.A1(new_n827_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1   g696(.A1(new_n822_), .A2(new_n824_), .ZN(new_n833_));
  NAND2_X1   g697(.A1(new_n833_), .A2(new_n830_), .ZN(new_n834_));
  NAND2_X1   g698(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1    g699(.A1(\A[16] ), .A2(\A[17] ), .ZN(new_n836_));
  NAND2_X1   g700(.A1(new_n827_), .A2(new_n829_), .ZN(new_n837_));
  NAND2_X1   g701(.A1(new_n837_), .A2(new_n836_), .ZN(new_n838_));
  OAI21_X1   g702(.A1(new_n835_), .A2(new_n836_), .B(new_n838_), .ZN(new_n839_));
  NOR2_X1    g703(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n840_));
  NAND2_X1   g704(.A1(new_n835_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1   g705(.A1(new_n839_), .A2(new_n840_), .B(new_n841_), .ZN(new_n842_));
  NAND2_X1   g706(.A1(new_n842_), .A2(new_n595_), .ZN(new_n843_));
  NOR2_X1    g707(.A1(\A[12] ), .A2(\A[13] ), .ZN(new_n844_));
  NAND2_X1   g708(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1   g709(.A1(new_n842_), .A2(new_n844_), .B(new_n845_), .ZN(new_n846_));
  OAI21_X1   g710(.A1(new_n846_), .A2(new_n595_), .B(new_n843_), .ZN(new_n847_));
  NOR2_X1    g711(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n848_));
  NAND2_X1   g712(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1   g713(.A1(new_n847_), .A2(new_n848_), .B(new_n849_), .ZN(new_n850_));
  NAND2_X1   g714(.A1(new_n573_), .A2(new_n583_), .ZN(new_n851_));
  OR2_X2     g715(.A1(\A[2] ), .A2(\A[3] ), .Z(new_n852_));
  NOR2_X1    g716(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n853_));
  AOI21_X1   g717(.A1(new_n852_), .A2(new_n853_), .B(new_n851_), .ZN(new_n854_));
  NAND2_X1   g718(.A1(new_n847_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1   g719(.A1(new_n850_), .A2(new_n854_), .B(new_n855_), .ZN(\P[1] ));
  NOR3_X1    g720(.A1(new_n831_), .A2(\A[16] ), .A3(\A[17] ), .ZN(new_n857_));
  INV_X1     g721(.I(new_n857_), .ZN(new_n858_));
  NAND2_X1   g722(.A1(new_n810_), .A2(new_n815_), .ZN(new_n859_));
  NOR2_X1    g723(.A1(new_n792_), .A2(new_n797_), .ZN(new_n860_));
  INV_X1     g724(.I(new_n860_), .ZN(new_n861_));
  NOR2_X1    g725(.A1(new_n772_), .A2(new_n777_), .ZN(new_n862_));
  INV_X1     g726(.I(new_n862_), .ZN(new_n863_));
  NOR2_X1    g727(.A1(new_n752_), .A2(new_n757_), .ZN(new_n864_));
  INV_X1     g728(.I(new_n864_), .ZN(new_n865_));
  NOR2_X1    g729(.A1(new_n732_), .A2(new_n737_), .ZN(new_n866_));
  INV_X1     g730(.I(new_n866_), .ZN(new_n867_));
  NOR2_X1    g731(.A1(new_n712_), .A2(new_n717_), .ZN(new_n868_));
  INV_X1     g732(.I(new_n868_), .ZN(new_n869_));
  NOR2_X1    g733(.A1(new_n692_), .A2(new_n697_), .ZN(new_n870_));
  INV_X1     g734(.I(new_n870_), .ZN(new_n871_));
  NOR2_X1    g735(.A1(new_n673_), .A2(new_n677_), .ZN(new_n872_));
  INV_X1     g736(.I(new_n872_), .ZN(new_n873_));
  NAND2_X1   g737(.A1(new_n659_), .A2(new_n662_), .ZN(new_n874_));
  NAND2_X1   g738(.A1(new_n645_), .A2(new_n648_), .ZN(new_n875_));
  NOR2_X1    g739(.A1(new_n629_), .A2(new_n636_), .ZN(new_n876_));
  INV_X1     g740(.I(new_n876_), .ZN(new_n877_));
  NAND2_X1   g741(.A1(new_n602_), .A2(new_n597_), .ZN(new_n878_));
  INV_X1     g742(.I(new_n878_), .ZN(new_n879_));
  NAND3_X1   g743(.A1(new_n598_), .A2(new_n172_), .A3(new_n184_), .ZN(new_n880_));
  NAND2_X1   g744(.A1(new_n607_), .A2(new_n610_), .ZN(new_n881_));
  INV_X1     g745(.I(new_n881_), .ZN(new_n882_));
  OAI21_X1   g746(.A1(new_n880_), .A2(new_n882_), .B(new_n879_), .ZN(new_n883_));
  NAND2_X1   g747(.A1(new_n617_), .A2(new_n193_), .ZN(new_n884_));
  INV_X1     g748(.I(new_n884_), .ZN(new_n885_));
  NOR2_X1    g749(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1   g750(.A1(new_n882_), .A2(\A[115] ), .B(new_n880_), .ZN(new_n887_));
  NOR3_X1    g751(.A1(new_n887_), .A2(new_n878_), .A3(new_n884_), .ZN(new_n888_));
  NOR3_X1    g752(.A1(new_n886_), .A2(new_n888_), .A3(new_n877_), .ZN(new_n889_));
  NOR2_X1    g753(.A1(new_n886_), .A2(new_n888_), .ZN(new_n890_));
  INV_X1     g754(.I(new_n890_), .ZN(new_n891_));
  NAND2_X1   g755(.A1(new_n621_), .A2(new_n624_), .ZN(new_n892_));
  NOR2_X1    g756(.A1(new_n883_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1   g757(.A1(new_n891_), .A2(new_n892_), .B(new_n893_), .ZN(new_n894_));
  AOI21_X1   g758(.A1(new_n894_), .A2(new_n877_), .B(new_n889_), .ZN(new_n895_));
  NOR2_X1    g759(.A1(new_n895_), .A2(new_n875_), .ZN(new_n896_));
  NAND2_X1   g760(.A1(new_n596_), .A2(new_n640_), .ZN(new_n897_));
  NOR2_X1    g761(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1   g762(.A1(new_n895_), .A2(new_n897_), .B(new_n898_), .ZN(new_n899_));
  AOI21_X1   g763(.A1(new_n899_), .A2(new_n875_), .B(new_n896_), .ZN(new_n900_));
  NOR2_X1    g764(.A1(new_n900_), .A2(new_n874_), .ZN(new_n901_));
  NAND2_X1   g765(.A1(new_n653_), .A2(new_n656_), .ZN(new_n902_));
  NOR2_X1    g766(.A1(new_n899_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1   g767(.A1(new_n900_), .A2(new_n902_), .B(new_n903_), .ZN(new_n904_));
  AOI21_X1   g768(.A1(new_n904_), .A2(new_n874_), .B(new_n901_), .ZN(new_n905_));
  NOR2_X1    g769(.A1(new_n905_), .A2(new_n873_), .ZN(new_n906_));
  NAND2_X1   g770(.A1(new_n665_), .A2(new_n669_), .ZN(new_n907_));
  NOR2_X1    g771(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1   g772(.A1(new_n905_), .A2(new_n907_), .B(new_n908_), .ZN(new_n909_));
  AOI21_X1   g773(.A1(new_n909_), .A2(new_n873_), .B(new_n906_), .ZN(new_n910_));
  NOR2_X1    g774(.A1(new_n910_), .A2(new_n871_), .ZN(new_n911_));
  NOR2_X1    g775(.A1(new_n684_), .A2(new_n688_), .ZN(new_n912_));
  INV_X1     g776(.I(new_n912_), .ZN(new_n913_));
  NOR2_X1    g777(.A1(new_n909_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1   g778(.A1(new_n910_), .A2(new_n913_), .B(new_n914_), .ZN(new_n915_));
  AOI21_X1   g779(.A1(new_n915_), .A2(new_n871_), .B(new_n911_), .ZN(new_n916_));
  NOR2_X1    g780(.A1(new_n916_), .A2(new_n869_), .ZN(new_n917_));
  NOR2_X1    g781(.A1(new_n702_), .A2(new_n707_), .ZN(new_n918_));
  INV_X1     g782(.I(new_n918_), .ZN(new_n919_));
  NOR2_X1    g783(.A1(new_n915_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1   g784(.A1(new_n916_), .A2(new_n919_), .B(new_n920_), .ZN(new_n921_));
  AOI21_X1   g785(.A1(new_n921_), .A2(new_n869_), .B(new_n917_), .ZN(new_n922_));
  NOR2_X1    g786(.A1(new_n922_), .A2(new_n867_), .ZN(new_n923_));
  NOR2_X1    g787(.A1(new_n722_), .A2(new_n727_), .ZN(new_n924_));
  INV_X1     g788(.I(new_n924_), .ZN(new_n925_));
  NOR2_X1    g789(.A1(new_n921_), .A2(new_n925_), .ZN(new_n926_));
  AOI21_X1   g790(.A1(new_n922_), .A2(new_n925_), .B(new_n926_), .ZN(new_n927_));
  AOI21_X1   g791(.A1(new_n927_), .A2(new_n867_), .B(new_n923_), .ZN(new_n928_));
  NOR2_X1    g792(.A1(new_n928_), .A2(new_n865_), .ZN(new_n929_));
  NOR2_X1    g793(.A1(new_n742_), .A2(new_n747_), .ZN(new_n930_));
  INV_X1     g794(.I(new_n930_), .ZN(new_n931_));
  NOR2_X1    g795(.A1(new_n927_), .A2(new_n931_), .ZN(new_n932_));
  AOI21_X1   g796(.A1(new_n928_), .A2(new_n931_), .B(new_n932_), .ZN(new_n933_));
  AOI21_X1   g797(.A1(new_n933_), .A2(new_n865_), .B(new_n929_), .ZN(new_n934_));
  NOR2_X1    g798(.A1(new_n934_), .A2(new_n863_), .ZN(new_n935_));
  NOR2_X1    g799(.A1(new_n762_), .A2(new_n767_), .ZN(new_n936_));
  INV_X1     g800(.I(new_n936_), .ZN(new_n937_));
  NOR2_X1    g801(.A1(new_n933_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1   g802(.A1(new_n934_), .A2(new_n937_), .B(new_n938_), .ZN(new_n939_));
  AOI21_X1   g803(.A1(new_n939_), .A2(new_n863_), .B(new_n935_), .ZN(new_n940_));
  NOR2_X1    g804(.A1(new_n940_), .A2(new_n861_), .ZN(new_n941_));
  NOR2_X1    g805(.A1(new_n782_), .A2(new_n787_), .ZN(new_n942_));
  INV_X1     g806(.I(new_n942_), .ZN(new_n943_));
  NOR2_X1    g807(.A1(new_n939_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1   g808(.A1(new_n940_), .A2(new_n943_), .B(new_n944_), .ZN(new_n945_));
  AOI21_X1   g809(.A1(new_n945_), .A2(new_n861_), .B(new_n941_), .ZN(new_n946_));
  NOR2_X1    g810(.A1(new_n946_), .A2(new_n859_), .ZN(new_n947_));
  NAND2_X1   g811(.A1(new_n802_), .A2(new_n806_), .ZN(new_n948_));
  NOR2_X1    g812(.A1(new_n945_), .A2(new_n948_), .ZN(new_n949_));
  AOI21_X1   g813(.A1(new_n946_), .A2(new_n948_), .B(new_n949_), .ZN(new_n950_));
  AOI21_X1   g814(.A1(new_n950_), .A2(new_n859_), .B(new_n947_), .ZN(new_n951_));
  NOR2_X1    g815(.A1(new_n951_), .A2(new_n858_), .ZN(new_n952_));
  NOR2_X1    g816(.A1(new_n821_), .A2(new_n826_), .ZN(new_n953_));
  INV_X1     g817(.I(new_n953_), .ZN(new_n954_));
  NOR2_X1    g818(.A1(new_n950_), .A2(new_n954_), .ZN(new_n955_));
  AOI21_X1   g819(.A1(new_n951_), .A2(new_n954_), .B(new_n955_), .ZN(new_n956_));
  AOI21_X1   g820(.A1(new_n956_), .A2(new_n858_), .B(new_n952_), .ZN(new_n957_));
  NOR3_X1    g821(.A1(new_n851_), .A2(\A[4] ), .A3(\A[5] ), .ZN(new_n958_));
  NAND2_X1   g822(.A1(new_n595_), .A2(new_n848_), .ZN(new_n959_));
  NOR4_X1    g823(.A1(\A[12] ), .A2(\A[13] ), .A3(\A[14] ), .A4(\A[15] ), .ZN(new_n960_));
  OAI21_X1   g824(.A1(new_n958_), .A2(new_n959_), .B(new_n960_), .ZN(new_n961_));
  NOR2_X1    g825(.A1(new_n956_), .A2(new_n961_), .ZN(new_n962_));
  AOI21_X1   g826(.A1(new_n957_), .A2(new_n961_), .B(new_n962_), .ZN(\P[2] ));
  NOR2_X1    g827(.A1(new_n861_), .A2(new_n943_), .ZN(new_n964_));
  INV_X1     g828(.I(new_n964_), .ZN(new_n965_));
  NOR2_X1    g829(.A1(new_n865_), .A2(new_n931_), .ZN(new_n966_));
  INV_X1     g830(.I(new_n966_), .ZN(new_n967_));
  NOR2_X1    g831(.A1(new_n869_), .A2(new_n919_), .ZN(new_n968_));
  INV_X1     g832(.I(new_n968_), .ZN(new_n969_));
  NOR2_X1    g833(.A1(new_n873_), .A2(new_n907_), .ZN(new_n970_));
  INV_X1     g834(.I(new_n970_), .ZN(new_n971_));
  NOR2_X1    g835(.A1(new_n878_), .A2(new_n880_), .ZN(new_n972_));
  INV_X1     g836(.I(new_n972_), .ZN(new_n973_));
  NOR2_X1    g837(.A1(new_n877_), .A2(new_n892_), .ZN(new_n974_));
  INV_X1     g838(.I(new_n974_), .ZN(new_n975_));
  NOR3_X1    g839(.A1(new_n881_), .A2(new_n884_), .A3(\A[115] ), .ZN(new_n976_));
  AOI21_X1   g840(.A1(new_n975_), .A2(new_n976_), .B(new_n973_), .ZN(new_n977_));
  INV_X1     g841(.I(new_n875_), .ZN(new_n978_));
  NAND3_X1   g842(.A1(new_n978_), .A2(new_n235_), .A3(new_n640_), .ZN(new_n979_));
  AND2_X2    g843(.A1(new_n977_), .A2(new_n979_), .Z(new_n980_));
  INV_X1     g844(.I(new_n976_), .ZN(new_n981_));
  AOI21_X1   g845(.A1(new_n974_), .A2(\A[103] ), .B(new_n981_), .ZN(new_n982_));
  NOR3_X1    g846(.A1(new_n982_), .A2(new_n973_), .A3(new_n979_), .ZN(new_n983_));
  NOR3_X1    g847(.A1(new_n980_), .A2(new_n983_), .A3(new_n971_), .ZN(new_n984_));
  NOR2_X1    g848(.A1(new_n874_), .A2(new_n902_), .ZN(new_n985_));
  NOR2_X1    g849(.A1(new_n980_), .A2(new_n983_), .ZN(new_n986_));
  NOR2_X1    g850(.A1(new_n986_), .A2(new_n985_), .ZN(new_n987_));
  AOI21_X1   g851(.A1(new_n977_), .A2(new_n985_), .B(new_n987_), .ZN(new_n988_));
  AOI21_X1   g852(.A1(new_n988_), .A2(new_n971_), .B(new_n984_), .ZN(new_n989_));
  NOR2_X1    g853(.A1(new_n989_), .A2(new_n969_), .ZN(new_n990_));
  NOR2_X1    g854(.A1(new_n871_), .A2(new_n913_), .ZN(new_n991_));
  INV_X1     g855(.I(new_n991_), .ZN(new_n992_));
  NOR2_X1    g856(.A1(new_n988_), .A2(new_n992_), .ZN(new_n993_));
  AOI21_X1   g857(.A1(new_n989_), .A2(new_n992_), .B(new_n993_), .ZN(new_n994_));
  AOI21_X1   g858(.A1(new_n994_), .A2(new_n969_), .B(new_n990_), .ZN(new_n995_));
  NOR2_X1    g859(.A1(new_n995_), .A2(new_n967_), .ZN(new_n996_));
  NOR2_X1    g860(.A1(new_n867_), .A2(new_n925_), .ZN(new_n997_));
  INV_X1     g861(.I(new_n997_), .ZN(new_n998_));
  NOR2_X1    g862(.A1(new_n994_), .A2(new_n998_), .ZN(new_n999_));
  AOI21_X1   g863(.A1(new_n995_), .A2(new_n998_), .B(new_n999_), .ZN(new_n1000_));
  AOI21_X1   g864(.A1(new_n1000_), .A2(new_n967_), .B(new_n996_), .ZN(new_n1001_));
  NOR2_X1    g865(.A1(new_n1001_), .A2(new_n965_), .ZN(new_n1002_));
  NOR2_X1    g866(.A1(new_n863_), .A2(new_n937_), .ZN(new_n1003_));
  INV_X1     g867(.I(new_n1003_), .ZN(new_n1004_));
  NOR2_X1    g868(.A1(new_n1000_), .A2(new_n1004_), .ZN(new_n1005_));
  AOI21_X1   g869(.A1(new_n1001_), .A2(new_n1004_), .B(new_n1005_), .ZN(new_n1006_));
  AOI21_X1   g870(.A1(new_n1006_), .A2(new_n965_), .B(new_n1002_), .ZN(new_n1007_));
  NOR2_X1    g871(.A1(new_n859_), .A2(new_n948_), .ZN(new_n1008_));
  NAND3_X1   g872(.A1(new_n960_), .A2(new_n595_), .A3(new_n848_), .ZN(new_n1009_));
  NOR2_X1    g873(.A1(new_n858_), .A2(new_n954_), .ZN(new_n1010_));
  NAND2_X1   g874(.A1(new_n1010_), .A2(new_n1009_), .ZN(new_n1011_));
  NAND2_X1   g875(.A1(new_n1011_), .A2(new_n1008_), .ZN(new_n1012_));
  NOR2_X1    g876(.A1(new_n1006_), .A2(new_n1012_), .ZN(new_n1013_));
  AOI21_X1   g877(.A1(new_n1007_), .A2(new_n1012_), .B(new_n1013_), .ZN(\P[3] ));
  NAND2_X1   g878(.A1(new_n972_), .A2(new_n976_), .ZN(new_n1015_));
  INV_X1     g879(.I(new_n1015_), .ZN(new_n1016_));
  NAND2_X1   g880(.A1(new_n970_), .A2(new_n985_), .ZN(new_n1017_));
  INV_X1     g881(.I(new_n1017_), .ZN(new_n1018_));
  NAND4_X1   g882(.A1(new_n974_), .A2(new_n596_), .A3(new_n640_), .A4(new_n978_), .ZN(new_n1019_));
  OAI21_X1   g883(.A1(new_n1018_), .A2(new_n1019_), .B(new_n1016_), .ZN(new_n1020_));
  NOR4_X1    g884(.A1(new_n969_), .A2(\A[78] ), .A3(new_n684_), .A4(new_n871_), .ZN(new_n1021_));
  AOI21_X1   g885(.A1(new_n1018_), .A2(\A[79] ), .B(new_n1019_), .ZN(new_n1022_));
  NAND2_X1   g886(.A1(new_n1021_), .A2(new_n1016_), .ZN(new_n1023_));
  OAI22_X1   g887(.A1(new_n1023_), .A2(new_n1022_), .B1(new_n1020_), .B2(new_n1021_), .ZN(new_n1024_));
  NAND2_X1   g888(.A1(new_n966_), .A2(new_n997_), .ZN(new_n1025_));
  NAND2_X1   g889(.A1(new_n1010_), .A2(new_n1008_), .ZN(new_n1026_));
  NOR2_X1    g890(.A1(new_n965_), .A2(new_n1004_), .ZN(new_n1027_));
  AOI21_X1   g891(.A1(new_n1027_), .A2(new_n1026_), .B(new_n1025_), .ZN(new_n1028_));
  NAND2_X1   g892(.A1(new_n1028_), .A2(new_n1020_), .ZN(new_n1029_));
  OAI21_X1   g893(.A1(new_n1024_), .A2(new_n1028_), .B(new_n1029_), .ZN(\P[4] ));
  NOR2_X1    g894(.A1(new_n1019_), .A2(new_n1015_), .ZN(new_n1031_));
  NOR3_X1    g895(.A1(new_n1025_), .A2(new_n965_), .A3(new_n1004_), .ZN(new_n1032_));
  NOR3_X1    g896(.A1(new_n1017_), .A2(new_n969_), .A3(new_n992_), .ZN(new_n1033_));
  INV_X1     g897(.I(new_n1033_), .ZN(new_n1034_));
  OAI21_X1   g898(.A1(new_n1034_), .A2(new_n1032_), .B(new_n1031_), .ZN(\P[5] ));
  NAND2_X1   g899(.A1(new_n1033_), .A2(new_n1031_), .ZN(\P[6] ));
  NOR3_X1    g900(.A1(new_n852_), .A2(\A[0] ), .A3(\A[1] ), .ZN(new_n1037_));
  NOR2_X1    g901(.A1(new_n1026_), .A2(new_n1009_), .ZN(new_n1038_));
  NOR4_X1    g902(.A1(\P[6] ), .A2(new_n965_), .A3(new_n1004_), .A4(new_n1025_), .ZN(new_n1039_));
  NAND4_X1   g903(.A1(new_n1039_), .A2(new_n958_), .A3(new_n1037_), .A4(new_n1038_), .ZN(F));
endmodule


