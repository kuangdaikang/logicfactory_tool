// Benchmark "testing" written by ABC on Fri Feb 25 15:13:07 2022

module g36 ( 
    A743, A742, A741, A740, A739, A738, A676, A675, A674, A673, A672, A671,
    A609, A608, A607, A606, A605, A604, A542, A541, A540, A539, A538, A537,
    A475, A474, A473, A472, A471, A470, A403, A404, A405, A406, A407, A408,
    A347, A346, A345, A344, A343, A342, A280, A279, A278, A277, A276, A275,
    A213, A212, A211, A210, A209, A208, A146, A145, A144, A143, A142, A141,
    A79, A78, A77, A76, A75, A74, A7, A8, A9, A10, A11, A12  );
  input  A743, A742, A741, A740, A739, A738, A676, A675, A674, A673,
    A672, A671, A609, A608, A607, A606, A605, A604, A542, A541, A540, A539,
    A538, A537, A475, A474, A473, A472, A471, A470, A403, A404, A405, A406,
    A407, A408;
  output A347, A346, A345, A344, A343, A342, A280, A279, A278, A277, A276,
    A275, A213, A212, A211, A210, A209, A208, A146, A145, A144, A143, A142,
    A141, A79, A78, A77, A76, A75, A74, A7, A8, A9, A10, A11, A12;
  wire new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n261_, new_n262_, new_n263_,
    new_n265_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n287_, new_n288_, new_n289_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n345_, new_n346_, new_n347_,
    new_n349_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n371_, new_n372_, new_n373_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n423_, new_n424_, new_n425_,
    new_n427_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n449_, new_n450_, new_n451_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n518_, new_n519_, new_n520_, new_n522_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_;
  assign new_n73_ = ~A471 & A470;
  assign new_n74_ = ~A471 & ~new_n73_;
  assign new_n75_ = A471 & ~A470;
  assign new_n76_ = ~new_n73_ & ~new_n75_;
  assign new_n77_ = ~A472 & new_n76_;
  assign new_n78_ = ~A473 & ~A472;
  assign new_n79_ = ~new_n77_ & new_n78_;
  assign new_n80_ = new_n77_ & ~new_n78_;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign new_n82_ = A475 & ~new_n76_;
  assign new_n83_ = A475 & new_n76_;
  assign new_n84_ = ~A475 & ~new_n76_;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = ~new_n82_ & new_n85_;
  assign new_n87_ = ~A474 & ~new_n86_;
  assign new_n88_ = ~A475 & new_n76_;
  assign new_n89_ = ~new_n83_ & ~new_n88_;
  assign new_n90_ = ~new_n84_ & new_n89_;
  assign new_n91_ = A474 & ~new_n90_;
  assign new_n92_ = ~new_n87_ & ~new_n91_;
  assign new_n93_ = ~new_n81_ & new_n92_;
  assign new_n94_ = new_n78_ & new_n93_;
  assign new_n95_ = ~new_n78_ & ~new_n93_;
  assign new_n96_ = ~new_n94_ & ~new_n95_;
  assign new_n97_ = ~A474 & new_n96_;
  assign new_n98_ = new_n74_ & ~new_n97_;
  assign new_n99_ = new_n74_ & ~new_n98_;
  assign new_n100_ = A403 & ~A404;
  assign new_n101_ = ~A404 & ~new_n100_;
  assign new_n102_ = ~A405 & ~new_n101_;
  assign new_n103_ = A405 & new_n101_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = A405 & ~A406;
  assign new_n106_ = ~A405 & A406;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = ~new_n104_ & ~new_n107_;
  assign new_n109_ = ~A403 & A404;
  assign new_n110_ = ~new_n100_ & ~new_n109_;
  assign new_n111_ = A408 & ~new_n110_;
  assign new_n112_ = A408 & new_n110_;
  assign new_n113_ = ~A408 & ~new_n110_;
  assign new_n114_ = ~new_n112_ & ~new_n113_;
  assign new_n115_ = ~new_n111_ & new_n114_;
  assign new_n116_ = ~A407 & ~new_n115_;
  assign new_n117_ = ~A408 & new_n110_;
  assign new_n118_ = ~new_n112_ & ~new_n117_;
  assign new_n119_ = ~new_n113_ & new_n118_;
  assign new_n120_ = A407 & ~new_n119_;
  assign new_n121_ = ~new_n116_ & ~new_n120_;
  assign new_n122_ = new_n108_ & new_n121_;
  assign new_n123_ = ~new_n108_ & ~new_n121_;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = ~new_n101_ & ~new_n124_;
  assign new_n126_ = new_n99_ & new_n125_;
  assign new_n127_ = new_n99_ & ~new_n126_;
  assign new_n128_ = ~A672 & A671;
  assign new_n129_ = ~A672 & ~new_n128_;
  assign new_n130_ = A672 & ~A671;
  assign new_n131_ = ~new_n128_ & ~new_n130_;
  assign new_n132_ = ~A673 & new_n131_;
  assign new_n133_ = ~A674 & ~A673;
  assign new_n134_ = ~new_n132_ & new_n133_;
  assign new_n135_ = new_n132_ & ~new_n133_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = A676 & ~new_n131_;
  assign new_n138_ = A676 & new_n131_;
  assign new_n139_ = ~A676 & ~new_n131_;
  assign new_n140_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = ~new_n137_ & new_n140_;
  assign new_n142_ = ~A675 & ~new_n141_;
  assign new_n143_ = ~A676 & new_n131_;
  assign new_n144_ = ~new_n138_ & ~new_n143_;
  assign new_n145_ = ~new_n139_ & new_n144_;
  assign new_n146_ = A675 & ~new_n145_;
  assign new_n147_ = ~new_n142_ & ~new_n146_;
  assign new_n148_ = ~new_n136_ & new_n147_;
  assign new_n149_ = new_n133_ & new_n148_;
  assign new_n150_ = ~new_n133_ & ~new_n148_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = ~A675 & new_n151_;
  assign new_n153_ = new_n129_ & ~new_n152_;
  assign new_n154_ = new_n129_ & ~new_n153_;
  assign new_n155_ = ~A538 & A537;
  assign new_n156_ = ~A538 & ~new_n155_;
  assign new_n157_ = A538 & ~A537;
  assign new_n158_ = ~new_n155_ & ~new_n157_;
  assign new_n159_ = ~A539 & new_n158_;
  assign new_n160_ = ~A540 & ~A539;
  assign new_n161_ = ~new_n159_ & new_n160_;
  assign new_n162_ = new_n159_ & ~new_n160_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = A542 & ~new_n158_;
  assign new_n165_ = A542 & new_n158_;
  assign new_n166_ = ~A542 & ~new_n158_;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = ~new_n164_ & new_n167_;
  assign new_n169_ = ~A541 & ~new_n168_;
  assign new_n170_ = ~A542 & new_n158_;
  assign new_n171_ = ~new_n165_ & ~new_n170_;
  assign new_n172_ = ~new_n166_ & new_n171_;
  assign new_n173_ = A541 & ~new_n172_;
  assign new_n174_ = ~new_n169_ & ~new_n173_;
  assign new_n175_ = ~new_n163_ & new_n174_;
  assign new_n176_ = new_n160_ & new_n175_;
  assign new_n177_ = ~new_n160_ & ~new_n175_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~A541 & new_n178_;
  assign new_n180_ = new_n156_ & ~new_n179_;
  assign new_n181_ = new_n156_ & ~new_n180_;
  assign new_n182_ = ~new_n99_ & ~new_n125_;
  assign new_n183_ = ~new_n126_ & ~new_n182_;
  assign new_n184_ = new_n181_ & new_n183_;
  assign new_n185_ = ~A605 & A604;
  assign new_n186_ = ~A605 & ~new_n185_;
  assign new_n187_ = A605 & ~A604;
  assign new_n188_ = ~new_n185_ & ~new_n187_;
  assign new_n189_ = ~A606 & new_n188_;
  assign new_n190_ = ~A607 & ~A606;
  assign new_n191_ = ~new_n189_ & new_n190_;
  assign new_n192_ = new_n189_ & ~new_n190_;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = A609 & ~new_n188_;
  assign new_n195_ = A609 & new_n188_;
  assign new_n196_ = ~A609 & ~new_n188_;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = ~new_n194_ & new_n197_;
  assign new_n199_ = ~A608 & ~new_n198_;
  assign new_n200_ = ~A609 & new_n188_;
  assign new_n201_ = ~new_n195_ & ~new_n200_;
  assign new_n202_ = ~new_n196_ & new_n201_;
  assign new_n203_ = A608 & ~new_n202_;
  assign new_n204_ = ~new_n199_ & ~new_n203_;
  assign new_n205_ = ~new_n193_ & new_n204_;
  assign new_n206_ = new_n190_ & new_n205_;
  assign new_n207_ = ~new_n190_ & ~new_n205_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = ~A608 & new_n208_;
  assign new_n210_ = new_n186_ & ~new_n209_;
  assign new_n211_ = new_n186_ & ~new_n210_;
  assign new_n212_ = new_n181_ & new_n211_;
  assign new_n213_ = ~new_n184_ & new_n212_;
  assign new_n214_ = new_n184_ & ~new_n212_;
  assign new_n215_ = ~new_n213_ & ~new_n214_;
  assign new_n216_ = ~A739 & A738;
  assign new_n217_ = ~A739 & ~new_n216_;
  assign new_n218_ = A739 & ~A738;
  assign new_n219_ = ~new_n216_ & ~new_n218_;
  assign new_n220_ = ~A740 & new_n219_;
  assign new_n221_ = ~A741 & ~A740;
  assign new_n222_ = ~new_n220_ & new_n221_;
  assign new_n223_ = new_n220_ & ~new_n221_;
  assign new_n224_ = ~new_n222_ & ~new_n223_;
  assign new_n225_ = A743 & ~new_n219_;
  assign new_n226_ = A743 & new_n219_;
  assign new_n227_ = ~A743 & ~new_n219_;
  assign new_n228_ = ~new_n226_ & ~new_n227_;
  assign new_n229_ = ~new_n225_ & new_n228_;
  assign new_n230_ = ~A742 & ~new_n229_;
  assign new_n231_ = ~A743 & new_n219_;
  assign new_n232_ = ~new_n226_ & ~new_n231_;
  assign new_n233_ = ~new_n227_ & new_n232_;
  assign new_n234_ = A742 & ~new_n233_;
  assign new_n235_ = ~new_n230_ & ~new_n234_;
  assign new_n236_ = ~new_n224_ & new_n235_;
  assign new_n237_ = new_n221_ & new_n236_;
  assign new_n238_ = ~new_n221_ & ~new_n236_;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign new_n240_ = ~A742 & new_n239_;
  assign new_n241_ = new_n217_ & ~new_n240_;
  assign new_n242_ = new_n217_ & ~new_n241_;
  assign new_n243_ = ~new_n183_ & ~new_n242_;
  assign new_n244_ = new_n183_ & ~new_n242_;
  assign new_n245_ = ~new_n183_ & new_n242_;
  assign new_n246_ = ~new_n244_ & ~new_n245_;
  assign new_n247_ = ~new_n243_ & new_n246_;
  assign new_n248_ = new_n154_ & ~new_n247_;
  assign new_n249_ = new_n183_ & new_n242_;
  assign new_n250_ = ~new_n244_ & ~new_n249_;
  assign new_n251_ = ~new_n245_ & new_n250_;
  assign new_n252_ = ~new_n154_ & ~new_n251_;
  assign new_n253_ = ~new_n248_ & ~new_n252_;
  assign new_n254_ = ~new_n215_ & new_n253_;
  assign new_n255_ = new_n212_ & new_n254_;
  assign new_n256_ = ~new_n212_ & ~new_n254_;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = new_n154_ & new_n257_;
  assign new_n259_ = new_n127_ & ~new_n258_;
  assign A347 = ~new_n127_ | new_n259_;
  assign new_n261_ = new_n215_ & new_n253_;
  assign new_n262_ = ~new_n215_ & ~new_n253_;
  assign new_n263_ = ~new_n261_ & ~new_n262_;
  assign A346 = ~new_n183_ & ~new_n263_;
  assign new_n265_ = new_n99_ & new_n254_;
  assign A345 = ~new_n183_ & ~new_n265_;
  assign new_n267_ = ~new_n99_ & ~new_n253_;
  assign new_n268_ = ~new_n183_ & ~new_n267_;
  assign new_n269_ = new_n183_ & ~new_n268_;
  assign new_n270_ = new_n183_ & new_n267_;
  assign new_n271_ = new_n269_ & ~new_n270_;
  assign new_n272_ = ~new_n253_ & ~new_n271_;
  assign A344 = ~new_n215_ | new_n272_;
  assign new_n274_ = ~new_n127_ & ~new_n267_;
  assign new_n275_ = new_n127_ & ~new_n274_;
  assign new_n276_ = new_n127_ & new_n267_;
  assign new_n277_ = new_n275_ & ~new_n276_;
  assign new_n278_ = ~new_n253_ & ~new_n277_;
  assign new_n279_ = ~new_n127_ & new_n181_;
  assign new_n280_ = new_n127_ & ~new_n181_;
  assign new_n281_ = ~new_n279_ & ~new_n280_;
  assign new_n282_ = ~new_n181_ & new_n211_;
  assign new_n283_ = new_n181_ & ~new_n211_;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = ~new_n281_ & ~new_n284_;
  assign A343 = new_n278_ | new_n285_;
  assign new_n287_ = new_n253_ & new_n285_;
  assign new_n288_ = ~new_n253_ & ~new_n285_;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign A342 = ~new_n127_ & ~new_n289_;
  assign new_n291_ = new_n81_ & new_n92_;
  assign new_n292_ = ~new_n81_ & ~new_n92_;
  assign new_n293_ = ~new_n291_ & ~new_n292_;
  assign new_n294_ = ~new_n76_ & ~new_n293_;
  assign new_n295_ = A404 & ~new_n121_;
  assign new_n296_ = ~new_n101_ & ~new_n295_;
  assign new_n297_ = new_n101_ & ~new_n296_;
  assign new_n298_ = new_n101_ & new_n295_;
  assign new_n299_ = new_n297_ & ~new_n298_;
  assign new_n300_ = ~new_n121_ & ~new_n299_;
  assign new_n301_ = ~new_n108_ & ~new_n300_;
  assign new_n302_ = ~new_n294_ & ~new_n301_;
  assign new_n303_ = ~new_n294_ & ~new_n302_;
  assign new_n304_ = new_n136_ & new_n147_;
  assign new_n305_ = ~new_n136_ & ~new_n147_;
  assign new_n306_ = ~new_n304_ & ~new_n305_;
  assign new_n307_ = ~new_n131_ & ~new_n306_;
  assign new_n308_ = new_n163_ & new_n174_;
  assign new_n309_ = ~new_n163_ & ~new_n174_;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = ~new_n158_ & ~new_n310_;
  assign new_n312_ = new_n294_ & new_n301_;
  assign new_n313_ = ~new_n302_ & ~new_n312_;
  assign new_n314_ = ~new_n311_ & new_n313_;
  assign new_n315_ = new_n193_ & new_n204_;
  assign new_n316_ = ~new_n193_ & ~new_n204_;
  assign new_n317_ = ~new_n315_ & ~new_n316_;
  assign new_n318_ = ~new_n188_ & ~new_n317_;
  assign new_n319_ = ~new_n311_ & ~new_n318_;
  assign new_n320_ = ~new_n314_ & new_n319_;
  assign new_n321_ = new_n314_ & ~new_n319_;
  assign new_n322_ = ~new_n320_ & ~new_n321_;
  assign new_n323_ = new_n224_ & new_n235_;
  assign new_n324_ = ~new_n224_ & ~new_n235_;
  assign new_n325_ = ~new_n323_ & ~new_n324_;
  assign new_n326_ = ~new_n219_ & ~new_n325_;
  assign new_n327_ = ~new_n313_ & new_n326_;
  assign new_n328_ = new_n313_ & new_n326_;
  assign new_n329_ = ~new_n313_ & ~new_n326_;
  assign new_n330_ = ~new_n328_ & ~new_n329_;
  assign new_n331_ = ~new_n327_ & new_n330_;
  assign new_n332_ = ~new_n307_ & ~new_n331_;
  assign new_n333_ = new_n313_ & ~new_n326_;
  assign new_n334_ = ~new_n328_ & ~new_n333_;
  assign new_n335_ = ~new_n329_ & new_n334_;
  assign new_n336_ = new_n307_ & ~new_n335_;
  assign new_n337_ = ~new_n332_ & ~new_n336_;
  assign new_n338_ = ~new_n322_ & new_n337_;
  assign new_n339_ = new_n319_ & new_n338_;
  assign new_n340_ = ~new_n319_ & ~new_n338_;
  assign new_n341_ = ~new_n339_ & ~new_n340_;
  assign new_n342_ = ~new_n307_ & new_n341_;
  assign new_n343_ = new_n303_ & ~new_n342_;
  assign A280 = ~new_n303_ | new_n343_;
  assign new_n345_ = new_n322_ & new_n337_;
  assign new_n346_ = ~new_n322_ & ~new_n337_;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign A279 = ~new_n313_ & ~new_n347_;
  assign new_n349_ = ~new_n294_ & new_n338_;
  assign A278 = ~new_n313_ & ~new_n349_;
  assign new_n351_ = new_n294_ & ~new_n337_;
  assign new_n352_ = ~new_n313_ & ~new_n351_;
  assign new_n353_ = new_n313_ & ~new_n352_;
  assign new_n354_ = new_n313_ & new_n351_;
  assign new_n355_ = new_n353_ & ~new_n354_;
  assign new_n356_ = ~new_n337_ & ~new_n355_;
  assign A277 = ~new_n322_ | new_n356_;
  assign new_n358_ = ~new_n303_ & ~new_n351_;
  assign new_n359_ = new_n303_ & ~new_n358_;
  assign new_n360_ = new_n303_ & new_n351_;
  assign new_n361_ = new_n359_ & ~new_n360_;
  assign new_n362_ = ~new_n337_ & ~new_n361_;
  assign new_n363_ = ~new_n303_ & ~new_n311_;
  assign new_n364_ = new_n303_ & new_n311_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = new_n311_ & ~new_n318_;
  assign new_n367_ = ~new_n311_ & new_n318_;
  assign new_n368_ = ~new_n366_ & ~new_n367_;
  assign new_n369_ = ~new_n365_ & ~new_n368_;
  assign A276 = new_n362_ | new_n369_;
  assign new_n371_ = new_n337_ & new_n369_;
  assign new_n372_ = ~new_n337_ & ~new_n369_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign A275 = ~new_n303_ & ~new_n373_;
  assign new_n375_ = ~A471 & new_n93_;
  assign new_n376_ = ~new_n76_ & ~new_n375_;
  assign new_n377_ = ~new_n110_ & ~new_n295_;
  assign new_n378_ = new_n110_ & ~new_n377_;
  assign new_n379_ = new_n110_ & new_n295_;
  assign new_n380_ = new_n378_ & ~new_n379_;
  assign new_n381_ = ~new_n121_ & ~new_n380_;
  assign new_n382_ = ~A405 & new_n110_;
  assign new_n383_ = ~A405 & ~A406;
  assign new_n384_ = ~new_n382_ & new_n383_;
  assign new_n385_ = new_n382_ & ~new_n383_;
  assign new_n386_ = ~new_n384_ & ~new_n385_;
  assign new_n387_ = ~new_n381_ & new_n386_;
  assign new_n388_ = ~new_n376_ & ~new_n387_;
  assign new_n389_ = ~new_n376_ & ~new_n388_;
  assign new_n390_ = ~A672 & new_n148_;
  assign new_n391_ = ~new_n131_ & ~new_n390_;
  assign new_n392_ = ~A538 & new_n175_;
  assign new_n393_ = ~new_n158_ & ~new_n392_;
  assign new_n394_ = new_n376_ & new_n387_;
  assign new_n395_ = ~new_n388_ & ~new_n394_;
  assign new_n396_ = ~new_n393_ & new_n395_;
  assign new_n397_ = ~A605 & new_n205_;
  assign new_n398_ = ~new_n188_ & ~new_n397_;
  assign new_n399_ = ~new_n393_ & ~new_n398_;
  assign new_n400_ = ~new_n396_ & new_n399_;
  assign new_n401_ = new_n396_ & ~new_n399_;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign new_n403_ = ~A739 & new_n236_;
  assign new_n404_ = ~new_n219_ & ~new_n403_;
  assign new_n405_ = ~new_n395_ & new_n404_;
  assign new_n406_ = new_n395_ & new_n404_;
  assign new_n407_ = ~new_n395_ & ~new_n404_;
  assign new_n408_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = ~new_n405_ & new_n408_;
  assign new_n410_ = ~new_n391_ & ~new_n409_;
  assign new_n411_ = new_n395_ & ~new_n404_;
  assign new_n412_ = ~new_n406_ & ~new_n411_;
  assign new_n413_ = ~new_n407_ & new_n412_;
  assign new_n414_ = new_n391_ & ~new_n413_;
  assign new_n415_ = ~new_n410_ & ~new_n414_;
  assign new_n416_ = ~new_n402_ & new_n415_;
  assign new_n417_ = new_n399_ & new_n416_;
  assign new_n418_ = ~new_n399_ & ~new_n416_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = ~new_n391_ & new_n419_;
  assign new_n421_ = new_n389_ & ~new_n420_;
  assign A213 = ~new_n389_ | new_n421_;
  assign new_n423_ = new_n402_ & new_n415_;
  assign new_n424_ = ~new_n402_ & ~new_n415_;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign A212 = ~new_n395_ & ~new_n425_;
  assign new_n427_ = ~new_n376_ & new_n416_;
  assign A211 = ~new_n395_ & ~new_n427_;
  assign new_n429_ = new_n376_ & ~new_n415_;
  assign new_n430_ = ~new_n395_ & ~new_n429_;
  assign new_n431_ = new_n395_ & ~new_n430_;
  assign new_n432_ = new_n395_ & new_n429_;
  assign new_n433_ = new_n431_ & ~new_n432_;
  assign new_n434_ = ~new_n415_ & ~new_n433_;
  assign A210 = ~new_n402_ | new_n434_;
  assign new_n436_ = ~new_n389_ & ~new_n429_;
  assign new_n437_ = new_n389_ & ~new_n436_;
  assign new_n438_ = new_n389_ & new_n429_;
  assign new_n439_ = new_n437_ & ~new_n438_;
  assign new_n440_ = ~new_n415_ & ~new_n439_;
  assign new_n441_ = ~new_n389_ & ~new_n393_;
  assign new_n442_ = new_n389_ & new_n393_;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign new_n444_ = new_n393_ & ~new_n398_;
  assign new_n445_ = ~new_n393_ & new_n398_;
  assign new_n446_ = ~new_n444_ & ~new_n445_;
  assign new_n447_ = ~new_n443_ & ~new_n446_;
  assign A209 = new_n440_ | new_n447_;
  assign new_n449_ = new_n415_ & new_n447_;
  assign new_n450_ = ~new_n415_ & ~new_n447_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign A208 = ~new_n389_ & ~new_n451_;
  assign new_n453_ = A471 & ~new_n92_;
  assign new_n454_ = ~new_n76_ & ~new_n453_;
  assign new_n455_ = new_n76_ & ~new_n454_;
  assign new_n456_ = new_n76_ & new_n453_;
  assign new_n457_ = new_n455_ & ~new_n456_;
  assign new_n458_ = ~new_n92_ & ~new_n457_;
  assign new_n459_ = new_n81_ & ~new_n458_;
  assign new_n460_ = new_n121_ & ~new_n386_;
  assign new_n461_ = ~A404 & new_n460_;
  assign new_n462_ = ~new_n110_ & ~new_n461_;
  assign new_n463_ = new_n459_ & new_n462_;
  assign new_n464_ = new_n459_ & ~new_n463_;
  assign new_n465_ = A672 & ~new_n147_;
  assign new_n466_ = ~new_n131_ & ~new_n465_;
  assign new_n467_ = new_n131_ & ~new_n466_;
  assign new_n468_ = new_n131_ & new_n465_;
  assign new_n469_ = new_n467_ & ~new_n468_;
  assign new_n470_ = ~new_n147_ & ~new_n469_;
  assign new_n471_ = new_n136_ & ~new_n470_;
  assign new_n472_ = A538 & ~new_n174_;
  assign new_n473_ = ~new_n158_ & ~new_n472_;
  assign new_n474_ = new_n158_ & ~new_n473_;
  assign new_n475_ = new_n158_ & new_n472_;
  assign new_n476_ = new_n474_ & ~new_n475_;
  assign new_n477_ = ~new_n174_ & ~new_n476_;
  assign new_n478_ = new_n163_ & ~new_n477_;
  assign new_n479_ = ~new_n459_ & ~new_n462_;
  assign new_n480_ = ~new_n463_ & ~new_n479_;
  assign new_n481_ = new_n478_ & new_n480_;
  assign new_n482_ = A605 & ~new_n204_;
  assign new_n483_ = ~new_n188_ & ~new_n482_;
  assign new_n484_ = new_n188_ & ~new_n483_;
  assign new_n485_ = new_n188_ & new_n482_;
  assign new_n486_ = new_n484_ & ~new_n485_;
  assign new_n487_ = ~new_n204_ & ~new_n486_;
  assign new_n488_ = new_n193_ & ~new_n487_;
  assign new_n489_ = new_n478_ & new_n488_;
  assign new_n490_ = ~new_n481_ & new_n489_;
  assign new_n491_ = new_n481_ & ~new_n489_;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = A739 & ~new_n235_;
  assign new_n494_ = ~new_n219_ & ~new_n493_;
  assign new_n495_ = new_n219_ & ~new_n494_;
  assign new_n496_ = new_n219_ & new_n493_;
  assign new_n497_ = new_n495_ & ~new_n496_;
  assign new_n498_ = ~new_n235_ & ~new_n497_;
  assign new_n499_ = new_n224_ & ~new_n498_;
  assign new_n500_ = ~new_n480_ & ~new_n499_;
  assign new_n501_ = new_n480_ & ~new_n499_;
  assign new_n502_ = ~new_n480_ & new_n499_;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign new_n504_ = ~new_n500_ & new_n503_;
  assign new_n505_ = new_n471_ & ~new_n504_;
  assign new_n506_ = new_n480_ & new_n499_;
  assign new_n507_ = ~new_n501_ & ~new_n506_;
  assign new_n508_ = ~new_n502_ & new_n507_;
  assign new_n509_ = ~new_n471_ & ~new_n508_;
  assign new_n510_ = ~new_n505_ & ~new_n509_;
  assign new_n511_ = ~new_n492_ & new_n510_;
  assign new_n512_ = new_n489_ & new_n511_;
  assign new_n513_ = ~new_n489_ & ~new_n511_;
  assign new_n514_ = ~new_n512_ & ~new_n513_;
  assign new_n515_ = new_n471_ & new_n514_;
  assign new_n516_ = new_n464_ & ~new_n515_;
  assign A146 = ~new_n464_ | new_n516_;
  assign new_n518_ = new_n492_ & new_n510_;
  assign new_n519_ = ~new_n492_ & ~new_n510_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign A145 = ~new_n480_ & ~new_n520_;
  assign new_n522_ = new_n459_ & new_n511_;
  assign A144 = ~new_n480_ & ~new_n522_;
  assign new_n524_ = ~new_n459_ & ~new_n510_;
  assign new_n525_ = ~new_n480_ & ~new_n524_;
  assign new_n526_ = new_n480_ & ~new_n525_;
  assign new_n527_ = new_n480_ & new_n524_;
  assign new_n528_ = new_n526_ & ~new_n527_;
  assign new_n529_ = ~new_n510_ & ~new_n528_;
  assign A143 = ~new_n492_ | new_n529_;
  assign new_n531_ = ~new_n464_ & ~new_n524_;
  assign new_n532_ = new_n464_ & ~new_n531_;
  assign new_n533_ = new_n464_ & new_n524_;
  assign new_n534_ = new_n532_ & ~new_n533_;
  assign new_n535_ = ~new_n510_ & ~new_n534_;
  assign new_n536_ = ~new_n464_ & new_n478_;
  assign new_n537_ = new_n464_ & ~new_n478_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~new_n478_ & new_n488_;
  assign new_n540_ = new_n478_ & ~new_n488_;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = ~new_n538_ & ~new_n541_;
  assign A142 = new_n535_ | new_n542_;
  assign new_n544_ = new_n510_ & new_n542_;
  assign new_n545_ = ~new_n510_ & ~new_n542_;
  assign new_n546_ = ~new_n544_ & ~new_n545_;
  assign A141 = ~new_n464_ & ~new_n546_;
  assign new_n548_ = ~new_n74_ & ~new_n453_;
  assign new_n549_ = new_n74_ & ~new_n548_;
  assign new_n550_ = new_n74_ & new_n453_;
  assign new_n551_ = new_n549_ & ~new_n550_;
  assign new_n552_ = ~new_n92_ & ~new_n551_;
  assign new_n553_ = ~A472 & ~new_n74_;
  assign new_n554_ = A472 & new_n74_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = ~A473 & A472;
  assign new_n557_ = A473 & ~A472;
  assign new_n558_ = ~new_n556_ & ~new_n557_;
  assign new_n559_ = ~new_n555_ & ~new_n558_;
  assign new_n560_ = ~new_n552_ & ~new_n559_;
  assign new_n561_ = new_n121_ & new_n386_;
  assign new_n562_ = ~new_n121_ & ~new_n386_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = ~new_n110_ & ~new_n563_;
  assign new_n565_ = new_n560_ & new_n564_;
  assign new_n566_ = new_n560_ & ~new_n565_;
  assign new_n567_ = ~new_n129_ & ~new_n465_;
  assign new_n568_ = new_n129_ & ~new_n567_;
  assign new_n569_ = new_n129_ & new_n465_;
  assign new_n570_ = new_n568_ & ~new_n569_;
  assign new_n571_ = ~new_n147_ & ~new_n570_;
  assign new_n572_ = ~A673 & ~new_n129_;
  assign new_n573_ = A673 & new_n129_;
  assign new_n574_ = ~new_n572_ & ~new_n573_;
  assign new_n575_ = ~A674 & A673;
  assign new_n576_ = A674 & ~A673;
  assign new_n577_ = ~new_n575_ & ~new_n576_;
  assign new_n578_ = ~new_n574_ & ~new_n577_;
  assign new_n579_ = ~new_n571_ & ~new_n578_;
  assign new_n580_ = ~new_n156_ & ~new_n472_;
  assign new_n581_ = new_n156_ & ~new_n580_;
  assign new_n582_ = new_n156_ & new_n472_;
  assign new_n583_ = new_n581_ & ~new_n582_;
  assign new_n584_ = ~new_n174_ & ~new_n583_;
  assign new_n585_ = ~A539 & ~new_n156_;
  assign new_n586_ = A539 & new_n156_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~A540 & A539;
  assign new_n589_ = A540 & ~A539;
  assign new_n590_ = ~new_n588_ & ~new_n589_;
  assign new_n591_ = ~new_n587_ & ~new_n590_;
  assign new_n592_ = ~new_n584_ & ~new_n591_;
  assign new_n593_ = ~new_n560_ & ~new_n564_;
  assign new_n594_ = ~new_n565_ & ~new_n593_;
  assign new_n595_ = new_n592_ & new_n594_;
  assign new_n596_ = ~new_n186_ & ~new_n482_;
  assign new_n597_ = new_n186_ & ~new_n596_;
  assign new_n598_ = new_n186_ & new_n482_;
  assign new_n599_ = new_n597_ & ~new_n598_;
  assign new_n600_ = ~new_n204_ & ~new_n599_;
  assign new_n601_ = ~A606 & ~new_n186_;
  assign new_n602_ = A606 & new_n186_;
  assign new_n603_ = ~new_n601_ & ~new_n602_;
  assign new_n604_ = ~A607 & A606;
  assign new_n605_ = A607 & ~A606;
  assign new_n606_ = ~new_n604_ & ~new_n605_;
  assign new_n607_ = ~new_n603_ & ~new_n606_;
  assign new_n608_ = ~new_n600_ & ~new_n607_;
  assign new_n609_ = new_n592_ & new_n608_;
  assign new_n610_ = ~new_n595_ & new_n609_;
  assign new_n611_ = new_n595_ & ~new_n609_;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = ~new_n217_ & ~new_n493_;
  assign new_n614_ = new_n217_ & ~new_n613_;
  assign new_n615_ = new_n217_ & new_n493_;
  assign new_n616_ = new_n614_ & ~new_n615_;
  assign new_n617_ = ~new_n235_ & ~new_n616_;
  assign new_n618_ = ~A740 & ~new_n217_;
  assign new_n619_ = A740 & new_n217_;
  assign new_n620_ = ~new_n618_ & ~new_n619_;
  assign new_n621_ = ~A741 & A740;
  assign new_n622_ = A741 & ~A740;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_ = ~new_n620_ & ~new_n623_;
  assign new_n625_ = ~new_n617_ & ~new_n624_;
  assign new_n626_ = ~new_n594_ & ~new_n625_;
  assign new_n627_ = new_n594_ & ~new_n625_;
  assign new_n628_ = ~new_n594_ & new_n625_;
  assign new_n629_ = ~new_n627_ & ~new_n628_;
  assign new_n630_ = ~new_n626_ & new_n629_;
  assign new_n631_ = new_n579_ & ~new_n630_;
  assign new_n632_ = new_n594_ & new_n625_;
  assign new_n633_ = ~new_n627_ & ~new_n632_;
  assign new_n634_ = ~new_n628_ & new_n633_;
  assign new_n635_ = ~new_n579_ & ~new_n634_;
  assign new_n636_ = ~new_n631_ & ~new_n635_;
  assign new_n637_ = ~new_n612_ & new_n636_;
  assign new_n638_ = new_n609_ & new_n637_;
  assign new_n639_ = ~new_n609_ & ~new_n637_;
  assign new_n640_ = ~new_n638_ & ~new_n639_;
  assign new_n641_ = new_n579_ & new_n640_;
  assign new_n642_ = new_n566_ & ~new_n641_;
  assign A79 = ~new_n566_ | new_n642_;
  assign new_n644_ = new_n612_ & new_n636_;
  assign new_n645_ = ~new_n612_ & ~new_n636_;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign A78 = ~new_n594_ & ~new_n646_;
  assign new_n648_ = new_n560_ & new_n637_;
  assign A77 = ~new_n594_ & ~new_n648_;
  assign new_n650_ = ~new_n560_ & ~new_n636_;
  assign new_n651_ = ~new_n594_ & ~new_n650_;
  assign new_n652_ = new_n594_ & ~new_n651_;
  assign new_n653_ = new_n594_ & new_n650_;
  assign new_n654_ = new_n652_ & ~new_n653_;
  assign new_n655_ = ~new_n636_ & ~new_n654_;
  assign A76 = ~new_n612_ | new_n655_;
  assign new_n657_ = ~new_n566_ & ~new_n650_;
  assign new_n658_ = new_n566_ & ~new_n657_;
  assign new_n659_ = new_n566_ & new_n650_;
  assign new_n660_ = new_n658_ & ~new_n659_;
  assign new_n661_ = ~new_n636_ & ~new_n660_;
  assign new_n662_ = ~new_n566_ & new_n592_;
  assign new_n663_ = new_n566_ & ~new_n592_;
  assign new_n664_ = ~new_n662_ & ~new_n663_;
  assign new_n665_ = ~new_n592_ & new_n608_;
  assign new_n666_ = new_n592_ & ~new_n608_;
  assign new_n667_ = ~new_n665_ & ~new_n666_;
  assign new_n668_ = ~new_n664_ & ~new_n667_;
  assign A75 = new_n661_ | new_n668_;
  assign new_n670_ = new_n636_ & new_n668_;
  assign new_n671_ = ~new_n636_ & ~new_n668_;
  assign new_n672_ = ~new_n670_ & ~new_n671_;
  assign A74 = ~new_n566_ & ~new_n672_;
  assign new_n674_ = new_n204_ & new_n607_;
  assign new_n675_ = ~new_n204_ & ~new_n607_;
  assign new_n676_ = ~new_n674_ & ~new_n675_;
  assign new_n677_ = ~new_n186_ & ~new_n676_;
  assign new_n678_ = new_n147_ & new_n578_;
  assign new_n679_ = ~new_n147_ & ~new_n578_;
  assign new_n680_ = ~new_n678_ & ~new_n679_;
  assign new_n681_ = ~new_n129_ & ~new_n680_;
  assign new_n682_ = new_n235_ & new_n624_;
  assign new_n683_ = ~new_n235_ & ~new_n624_;
  assign new_n684_ = ~new_n682_ & ~new_n683_;
  assign new_n685_ = ~new_n217_ & ~new_n684_;
  assign new_n686_ = ~new_n681_ & new_n685_;
  assign new_n687_ = ~new_n681_ & ~new_n686_;
  assign new_n688_ = ~new_n677_ & ~new_n687_;
  assign new_n689_ = new_n677_ & new_n687_;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = new_n174_ & new_n591_;
  assign new_n692_ = ~new_n174_ & ~new_n591_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = ~new_n156_ & ~new_n693_;
  assign new_n695_ = new_n677_ & ~new_n694_;
  assign new_n696_ = ~new_n677_ & new_n694_;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~new_n690_ & ~new_n697_;
  assign new_n699_ = new_n92_ & new_n559_;
  assign new_n700_ = ~new_n92_ & ~new_n559_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = ~new_n74_ & ~new_n701_;
  assign new_n703_ = new_n383_ & new_n460_;
  assign new_n704_ = ~new_n383_ & ~new_n460_;
  assign new_n705_ = ~new_n703_ & ~new_n704_;
  assign new_n706_ = ~A407 & new_n705_;
  assign new_n707_ = new_n101_ & ~new_n706_;
  assign new_n708_ = new_n101_ & ~new_n707_;
  assign new_n709_ = new_n681_ & ~new_n685_;
  assign new_n710_ = ~new_n686_ & ~new_n709_;
  assign new_n711_ = ~new_n708_ & ~new_n710_;
  assign new_n712_ = ~new_n708_ & new_n710_;
  assign new_n713_ = new_n708_ & ~new_n710_;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = ~new_n711_ & new_n714_;
  assign new_n716_ = ~new_n702_ & ~new_n715_;
  assign new_n717_ = new_n708_ & new_n710_;
  assign new_n718_ = ~new_n712_ & ~new_n717_;
  assign new_n719_ = ~new_n713_ & new_n718_;
  assign new_n720_ = new_n702_ & ~new_n719_;
  assign new_n721_ = ~new_n716_ & ~new_n720_;
  assign new_n722_ = new_n698_ & new_n721_;
  assign new_n723_ = ~new_n698_ & ~new_n721_;
  assign new_n724_ = ~new_n722_ & ~new_n723_;
  assign A7 = ~new_n687_ & ~new_n724_;
  assign new_n726_ = new_n681_ & ~new_n721_;
  assign new_n727_ = ~new_n687_ & ~new_n726_;
  assign new_n728_ = new_n687_ & ~new_n727_;
  assign new_n729_ = new_n687_ & new_n726_;
  assign new_n730_ = new_n728_ & ~new_n729_;
  assign new_n731_ = ~new_n721_ & ~new_n730_;
  assign A8 = new_n698_ | new_n731_;
  assign new_n733_ = ~new_n710_ & ~new_n726_;
  assign new_n734_ = new_n710_ & ~new_n733_;
  assign new_n735_ = new_n710_ & new_n726_;
  assign new_n736_ = new_n734_ & ~new_n735_;
  assign new_n737_ = ~new_n721_ & ~new_n736_;
  assign new_n738_ = ~new_n677_ & new_n710_;
  assign new_n739_ = ~new_n677_ & ~new_n694_;
  assign new_n740_ = ~new_n738_ & new_n739_;
  assign new_n741_ = new_n738_ & ~new_n739_;
  assign new_n742_ = ~new_n740_ & ~new_n741_;
  assign A9 = new_n737_ | ~new_n742_;
  assign new_n744_ = new_n721_ & ~new_n742_;
  assign new_n745_ = ~new_n681_ & new_n744_;
  assign A10 = ~new_n710_ & ~new_n745_;
  assign new_n747_ = new_n721_ & new_n742_;
  assign new_n748_ = ~new_n721_ & ~new_n742_;
  assign new_n749_ = ~new_n747_ & ~new_n748_;
  assign A11 = ~new_n710_ & ~new_n749_;
  assign new_n751_ = new_n739_ & new_n744_;
  assign new_n752_ = ~new_n739_ & ~new_n744_;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = ~new_n702_ & new_n753_;
  assign new_n755_ = new_n687_ & ~new_n754_;
  assign A12 = ~new_n687_ | new_n755_;
endmodule


