// Benchmark "adder" written by ABC on Mon Sep  4 17:55:01 2023

module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n431_, new_n432_, new_n433_, new_n434_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n467_, new_n468_, new_n469_, new_n470_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n503_, new_n504_, new_n505_, new_n506_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n539_, new_n540_, new_n541_, new_n542_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n575_, new_n576_, new_n577_, new_n578_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_;
  XOR2_X1    g000(.A1(\a[0] ), .A2(\b[0] ), .Z(\f[0] ));
  NAND2_X1   g001(.A1(\a[0] ), .A2(\b[0] ), .ZN(new_n387_));
  NOR2_X1    g002(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n388_));
  INV_X1     g003(.I(new_n388_), .ZN(new_n389_));
  NAND2_X1   g004(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n390_));
  NAND2_X1   g005(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1    g006(.A1(new_n391_), .A2(new_n387_), .Z(\f[1] ));
  OAI21_X1   g007(.A1(new_n387_), .A2(new_n388_), .B(new_n390_), .ZN(new_n393_));
  INV_X1     g008(.I(\a[2] ), .ZN(new_n394_));
  INV_X1     g009(.I(\b[2] ), .ZN(new_n395_));
  NAND2_X1   g010(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1     g011(.I(new_n396_), .ZN(new_n397_));
  NOR2_X1    g012(.A1(new_n394_), .A2(new_n395_), .ZN(new_n398_));
  NOR2_X1    g013(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XOR2_X1    g014(.A1(new_n399_), .A2(new_n393_), .Z(\f[2] ));
  AOI21_X1   g015(.A1(new_n393_), .A2(new_n396_), .B(new_n398_), .ZN(new_n401_));
  NOR2_X1    g016(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n402_));
  INV_X1     g017(.I(new_n402_), .ZN(new_n403_));
  NAND2_X1   g018(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n404_));
  NAND2_X1   g019(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1    g020(.A1(new_n401_), .A2(new_n405_), .Z(\f[3] ));
  OAI21_X1   g021(.A1(new_n401_), .A2(new_n402_), .B(new_n404_), .ZN(new_n407_));
  NOR2_X1    g022(.A1(\a[4] ), .A2(\b[4] ), .ZN(new_n408_));
  AND2_X2    g023(.A1(\a[4] ), .A2(\b[4] ), .Z(new_n409_));
  NOR2_X1    g024(.A1(new_n409_), .A2(new_n408_), .ZN(new_n410_));
  XOR2_X1    g025(.A1(new_n407_), .A2(new_n410_), .Z(\f[4] ));
  INV_X1     g026(.I(new_n408_), .ZN(new_n412_));
  AOI21_X1   g027(.A1(new_n407_), .A2(new_n412_), .B(new_n409_), .ZN(new_n413_));
  NOR2_X1    g028(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n414_));
  INV_X1     g029(.I(new_n414_), .ZN(new_n415_));
  NAND2_X1   g030(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n416_));
  NAND2_X1   g031(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XOR2_X1    g032(.A1(new_n413_), .A2(new_n417_), .Z(\f[5] ));
  OAI21_X1   g033(.A1(new_n413_), .A2(new_n414_), .B(new_n416_), .ZN(new_n419_));
  NOR2_X1    g034(.A1(\a[6] ), .A2(\b[6] ), .ZN(new_n420_));
  AND2_X2    g035(.A1(\a[6] ), .A2(\b[6] ), .Z(new_n421_));
  NOR2_X1    g036(.A1(new_n421_), .A2(new_n420_), .ZN(new_n422_));
  XOR2_X1    g037(.A1(new_n419_), .A2(new_n422_), .Z(\f[6] ));
  INV_X1     g038(.I(new_n420_), .ZN(new_n424_));
  AOI21_X1   g039(.A1(new_n419_), .A2(new_n424_), .B(new_n421_), .ZN(new_n425_));
  NOR2_X1    g040(.A1(\a[7] ), .A2(\b[7] ), .ZN(new_n426_));
  INV_X1     g041(.I(new_n426_), .ZN(new_n427_));
  NAND2_X1   g042(.A1(\a[7] ), .A2(\b[7] ), .ZN(new_n428_));
  NAND2_X1   g043(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XOR2_X1    g044(.A1(new_n425_), .A2(new_n429_), .Z(\f[7] ));
  OAI21_X1   g045(.A1(new_n425_), .A2(new_n426_), .B(new_n428_), .ZN(new_n431_));
  NOR2_X1    g046(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n432_));
  AND2_X2    g047(.A1(\a[8] ), .A2(\b[8] ), .Z(new_n433_));
  NOR2_X1    g048(.A1(new_n433_), .A2(new_n432_), .ZN(new_n434_));
  XOR2_X1    g049(.A1(new_n431_), .A2(new_n434_), .Z(\f[8] ));
  INV_X1     g050(.I(new_n432_), .ZN(new_n436_));
  AOI21_X1   g051(.A1(new_n431_), .A2(new_n436_), .B(new_n433_), .ZN(new_n437_));
  NOR2_X1    g052(.A1(\a[9] ), .A2(\b[9] ), .ZN(new_n438_));
  INV_X1     g053(.I(new_n438_), .ZN(new_n439_));
  NAND2_X1   g054(.A1(\a[9] ), .A2(\b[9] ), .ZN(new_n440_));
  NAND2_X1   g055(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1    g056(.A1(new_n437_), .A2(new_n441_), .Z(\f[9] ));
  OAI21_X1   g057(.A1(new_n437_), .A2(new_n438_), .B(new_n440_), .ZN(new_n443_));
  NOR2_X1    g058(.A1(\a[10] ), .A2(\b[10] ), .ZN(new_n444_));
  AND2_X2    g059(.A1(\a[10] ), .A2(\b[10] ), .Z(new_n445_));
  NOR2_X1    g060(.A1(new_n445_), .A2(new_n444_), .ZN(new_n446_));
  XOR2_X1    g061(.A1(new_n443_), .A2(new_n446_), .Z(\f[10] ));
  INV_X1     g062(.I(new_n444_), .ZN(new_n448_));
  AOI21_X1   g063(.A1(new_n443_), .A2(new_n448_), .B(new_n445_), .ZN(new_n449_));
  NOR2_X1    g064(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n450_));
  INV_X1     g065(.I(new_n450_), .ZN(new_n451_));
  NAND2_X1   g066(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n452_));
  NAND2_X1   g067(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1    g068(.A1(new_n449_), .A2(new_n453_), .Z(\f[11] ));
  OAI21_X1   g069(.A1(new_n449_), .A2(new_n450_), .B(new_n452_), .ZN(new_n455_));
  NOR2_X1    g070(.A1(\a[12] ), .A2(\b[12] ), .ZN(new_n456_));
  AND2_X2    g071(.A1(\a[12] ), .A2(\b[12] ), .Z(new_n457_));
  NOR2_X1    g072(.A1(new_n457_), .A2(new_n456_), .ZN(new_n458_));
  XOR2_X1    g073(.A1(new_n455_), .A2(new_n458_), .Z(\f[12] ));
  INV_X1     g074(.I(new_n456_), .ZN(new_n460_));
  AOI21_X1   g075(.A1(new_n455_), .A2(new_n460_), .B(new_n457_), .ZN(new_n461_));
  NOR2_X1    g076(.A1(\a[13] ), .A2(\b[13] ), .ZN(new_n462_));
  INV_X1     g077(.I(new_n462_), .ZN(new_n463_));
  NAND2_X1   g078(.A1(\a[13] ), .A2(\b[13] ), .ZN(new_n464_));
  NAND2_X1   g079(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1    g080(.A1(new_n461_), .A2(new_n465_), .Z(\f[13] ));
  OAI21_X1   g081(.A1(new_n461_), .A2(new_n462_), .B(new_n464_), .ZN(new_n467_));
  NOR2_X1    g082(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n468_));
  AND2_X2    g083(.A1(\a[14] ), .A2(\b[14] ), .Z(new_n469_));
  NOR2_X1    g084(.A1(new_n469_), .A2(new_n468_), .ZN(new_n470_));
  XOR2_X1    g085(.A1(new_n467_), .A2(new_n470_), .Z(\f[14] ));
  INV_X1     g086(.I(new_n468_), .ZN(new_n472_));
  AOI21_X1   g087(.A1(new_n467_), .A2(new_n472_), .B(new_n469_), .ZN(new_n473_));
  NOR2_X1    g088(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n474_));
  INV_X1     g089(.I(new_n474_), .ZN(new_n475_));
  NAND2_X1   g090(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n476_));
  NAND2_X1   g091(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1    g092(.A1(new_n473_), .A2(new_n477_), .Z(\f[15] ));
  OAI21_X1   g093(.A1(new_n473_), .A2(new_n474_), .B(new_n476_), .ZN(new_n479_));
  NOR2_X1    g094(.A1(\a[16] ), .A2(\b[16] ), .ZN(new_n480_));
  AND2_X2    g095(.A1(\a[16] ), .A2(\b[16] ), .Z(new_n481_));
  NOR2_X1    g096(.A1(new_n481_), .A2(new_n480_), .ZN(new_n482_));
  XOR2_X1    g097(.A1(new_n479_), .A2(new_n482_), .Z(\f[16] ));
  INV_X1     g098(.I(new_n480_), .ZN(new_n484_));
  AOI21_X1   g099(.A1(new_n479_), .A2(new_n484_), .B(new_n481_), .ZN(new_n485_));
  NOR2_X1    g100(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n486_));
  INV_X1     g101(.I(new_n486_), .ZN(new_n487_));
  NAND2_X1   g102(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n488_));
  NAND2_X1   g103(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1    g104(.A1(new_n485_), .A2(new_n489_), .Z(\f[17] ));
  OAI21_X1   g105(.A1(new_n485_), .A2(new_n486_), .B(new_n488_), .ZN(new_n491_));
  NOR2_X1    g106(.A1(\a[18] ), .A2(\b[18] ), .ZN(new_n492_));
  AND2_X2    g107(.A1(\a[18] ), .A2(\b[18] ), .Z(new_n493_));
  NOR2_X1    g108(.A1(new_n493_), .A2(new_n492_), .ZN(new_n494_));
  XOR2_X1    g109(.A1(new_n491_), .A2(new_n494_), .Z(\f[18] ));
  INV_X1     g110(.I(new_n492_), .ZN(new_n496_));
  AOI21_X1   g111(.A1(new_n491_), .A2(new_n496_), .B(new_n493_), .ZN(new_n497_));
  NOR2_X1    g112(.A1(\a[19] ), .A2(\b[19] ), .ZN(new_n498_));
  INV_X1     g113(.I(new_n498_), .ZN(new_n499_));
  NAND2_X1   g114(.A1(\a[19] ), .A2(\b[19] ), .ZN(new_n500_));
  NAND2_X1   g115(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1    g116(.A1(new_n497_), .A2(new_n501_), .Z(\f[19] ));
  OAI21_X1   g117(.A1(new_n497_), .A2(new_n498_), .B(new_n500_), .ZN(new_n503_));
  NOR2_X1    g118(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n504_));
  AND2_X2    g119(.A1(\a[20] ), .A2(\b[20] ), .Z(new_n505_));
  NOR2_X1    g120(.A1(new_n505_), .A2(new_n504_), .ZN(new_n506_));
  XOR2_X1    g121(.A1(new_n503_), .A2(new_n506_), .Z(\f[20] ));
  INV_X1     g122(.I(new_n504_), .ZN(new_n508_));
  AOI21_X1   g123(.A1(new_n503_), .A2(new_n508_), .B(new_n505_), .ZN(new_n509_));
  NOR2_X1    g124(.A1(\a[21] ), .A2(\b[21] ), .ZN(new_n510_));
  INV_X1     g125(.I(new_n510_), .ZN(new_n511_));
  NAND2_X1   g126(.A1(\a[21] ), .A2(\b[21] ), .ZN(new_n512_));
  NAND2_X1   g127(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1    g128(.A1(new_n509_), .A2(new_n513_), .Z(\f[21] ));
  OAI21_X1   g129(.A1(new_n509_), .A2(new_n510_), .B(new_n512_), .ZN(new_n515_));
  NOR2_X1    g130(.A1(\a[22] ), .A2(\b[22] ), .ZN(new_n516_));
  AND2_X2    g131(.A1(\a[22] ), .A2(\b[22] ), .Z(new_n517_));
  NOR2_X1    g132(.A1(new_n517_), .A2(new_n516_), .ZN(new_n518_));
  XOR2_X1    g133(.A1(new_n515_), .A2(new_n518_), .Z(\f[22] ));
  INV_X1     g134(.I(new_n516_), .ZN(new_n520_));
  AOI21_X1   g135(.A1(new_n515_), .A2(new_n520_), .B(new_n517_), .ZN(new_n521_));
  NOR2_X1    g136(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n522_));
  INV_X1     g137(.I(new_n522_), .ZN(new_n523_));
  NAND2_X1   g138(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n524_));
  NAND2_X1   g139(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1    g140(.A1(new_n521_), .A2(new_n525_), .Z(\f[23] ));
  OAI21_X1   g141(.A1(new_n521_), .A2(new_n522_), .B(new_n524_), .ZN(new_n527_));
  NOR2_X1    g142(.A1(\a[24] ), .A2(\b[24] ), .ZN(new_n528_));
  AND2_X2    g143(.A1(\a[24] ), .A2(\b[24] ), .Z(new_n529_));
  NOR2_X1    g144(.A1(new_n529_), .A2(new_n528_), .ZN(new_n530_));
  XOR2_X1    g145(.A1(new_n527_), .A2(new_n530_), .Z(\f[24] ));
  INV_X1     g146(.I(new_n528_), .ZN(new_n532_));
  AOI21_X1   g147(.A1(new_n527_), .A2(new_n532_), .B(new_n529_), .ZN(new_n533_));
  NOR2_X1    g148(.A1(\a[25] ), .A2(\b[25] ), .ZN(new_n534_));
  INV_X1     g149(.I(new_n534_), .ZN(new_n535_));
  NAND2_X1   g150(.A1(\a[25] ), .A2(\b[25] ), .ZN(new_n536_));
  NAND2_X1   g151(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1    g152(.A1(new_n533_), .A2(new_n537_), .Z(\f[25] ));
  OAI21_X1   g153(.A1(new_n533_), .A2(new_n534_), .B(new_n536_), .ZN(new_n539_));
  NOR2_X1    g154(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n540_));
  AND2_X2    g155(.A1(\a[26] ), .A2(\b[26] ), .Z(new_n541_));
  NOR2_X1    g156(.A1(new_n541_), .A2(new_n540_), .ZN(new_n542_));
  XOR2_X1    g157(.A1(new_n539_), .A2(new_n542_), .Z(\f[26] ));
  INV_X1     g158(.I(new_n540_), .ZN(new_n544_));
  AOI21_X1   g159(.A1(new_n539_), .A2(new_n544_), .B(new_n541_), .ZN(new_n545_));
  NOR2_X1    g160(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n546_));
  INV_X1     g161(.I(new_n546_), .ZN(new_n547_));
  NAND2_X1   g162(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n548_));
  NAND2_X1   g163(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1    g164(.A1(new_n545_), .A2(new_n549_), .Z(\f[27] ));
  OAI21_X1   g165(.A1(new_n545_), .A2(new_n546_), .B(new_n548_), .ZN(new_n551_));
  NOR2_X1    g166(.A1(\a[28] ), .A2(\b[28] ), .ZN(new_n552_));
  AND2_X2    g167(.A1(\a[28] ), .A2(\b[28] ), .Z(new_n553_));
  NOR2_X1    g168(.A1(new_n553_), .A2(new_n552_), .ZN(new_n554_));
  XOR2_X1    g169(.A1(new_n551_), .A2(new_n554_), .Z(\f[28] ));
  INV_X1     g170(.I(new_n552_), .ZN(new_n556_));
  AOI21_X1   g171(.A1(new_n551_), .A2(new_n556_), .B(new_n553_), .ZN(new_n557_));
  NOR2_X1    g172(.A1(\a[29] ), .A2(\b[29] ), .ZN(new_n558_));
  INV_X1     g173(.I(new_n558_), .ZN(new_n559_));
  NAND2_X1   g174(.A1(\a[29] ), .A2(\b[29] ), .ZN(new_n560_));
  NAND2_X1   g175(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1    g176(.A1(new_n557_), .A2(new_n561_), .Z(\f[29] ));
  OAI21_X1   g177(.A1(new_n557_), .A2(new_n558_), .B(new_n560_), .ZN(new_n563_));
  NOR2_X1    g178(.A1(\a[30] ), .A2(\b[30] ), .ZN(new_n564_));
  AND2_X2    g179(.A1(\a[30] ), .A2(\b[30] ), .Z(new_n565_));
  NOR2_X1    g180(.A1(new_n565_), .A2(new_n564_), .ZN(new_n566_));
  XOR2_X1    g181(.A1(new_n563_), .A2(new_n566_), .Z(\f[30] ));
  INV_X1     g182(.I(new_n564_), .ZN(new_n568_));
  AOI21_X1   g183(.A1(new_n563_), .A2(new_n568_), .B(new_n565_), .ZN(new_n569_));
  NOR2_X1    g184(.A1(\a[31] ), .A2(\b[31] ), .ZN(new_n570_));
  INV_X1     g185(.I(new_n570_), .ZN(new_n571_));
  NAND2_X1   g186(.A1(\a[31] ), .A2(\b[31] ), .ZN(new_n572_));
  NAND2_X1   g187(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1    g188(.A1(new_n569_), .A2(new_n573_), .Z(\f[31] ));
  OAI21_X1   g189(.A1(new_n569_), .A2(new_n570_), .B(new_n572_), .ZN(new_n575_));
  NOR2_X1    g190(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n576_));
  AND2_X2    g191(.A1(\a[32] ), .A2(\b[32] ), .Z(new_n577_));
  NOR2_X1    g192(.A1(new_n577_), .A2(new_n576_), .ZN(new_n578_));
  XOR2_X1    g193(.A1(new_n575_), .A2(new_n578_), .Z(\f[32] ));
  INV_X1     g194(.I(new_n576_), .ZN(new_n580_));
  AOI21_X1   g195(.A1(new_n575_), .A2(new_n580_), .B(new_n577_), .ZN(new_n581_));
  NOR2_X1    g196(.A1(\a[33] ), .A2(\b[33] ), .ZN(new_n582_));
  INV_X1     g197(.I(new_n582_), .ZN(new_n583_));
  NAND2_X1   g198(.A1(\a[33] ), .A2(\b[33] ), .ZN(new_n584_));
  NAND2_X1   g199(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1    g200(.A1(new_n581_), .A2(new_n585_), .Z(\f[33] ));
  OAI21_X1   g201(.A1(new_n581_), .A2(new_n582_), .B(new_n584_), .ZN(new_n587_));
  NOR2_X1    g202(.A1(\a[34] ), .A2(\b[34] ), .ZN(new_n588_));
  AND2_X2    g203(.A1(\a[34] ), .A2(\b[34] ), .Z(new_n589_));
  NOR2_X1    g204(.A1(new_n589_), .A2(new_n588_), .ZN(new_n590_));
  XOR2_X1    g205(.A1(new_n587_), .A2(new_n590_), .Z(\f[34] ));
  INV_X1     g206(.I(new_n588_), .ZN(new_n592_));
  AOI21_X1   g207(.A1(new_n587_), .A2(new_n592_), .B(new_n589_), .ZN(new_n593_));
  NOR2_X1    g208(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n594_));
  INV_X1     g209(.I(new_n594_), .ZN(new_n595_));
  NAND2_X1   g210(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n596_));
  NAND2_X1   g211(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1    g212(.A1(new_n593_), .A2(new_n597_), .Z(\f[35] ));
  OAI21_X1   g213(.A1(new_n593_), .A2(new_n594_), .B(new_n596_), .ZN(new_n599_));
  NOR2_X1    g214(.A1(\a[36] ), .A2(\b[36] ), .ZN(new_n600_));
  AND2_X2    g215(.A1(\a[36] ), .A2(\b[36] ), .Z(new_n601_));
  NOR2_X1    g216(.A1(new_n601_), .A2(new_n600_), .ZN(new_n602_));
  XOR2_X1    g217(.A1(new_n599_), .A2(new_n602_), .Z(\f[36] ));
  INV_X1     g218(.I(new_n600_), .ZN(new_n604_));
  AOI21_X1   g219(.A1(new_n599_), .A2(new_n604_), .B(new_n601_), .ZN(new_n605_));
  NOR2_X1    g220(.A1(\a[37] ), .A2(\b[37] ), .ZN(new_n606_));
  INV_X1     g221(.I(new_n606_), .ZN(new_n607_));
  NAND2_X1   g222(.A1(\a[37] ), .A2(\b[37] ), .ZN(new_n608_));
  NAND2_X1   g223(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1    g224(.A1(new_n605_), .A2(new_n609_), .Z(\f[37] ));
  OAI21_X1   g225(.A1(new_n605_), .A2(new_n606_), .B(new_n608_), .ZN(new_n611_));
  NOR2_X1    g226(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n612_));
  AND2_X2    g227(.A1(\a[38] ), .A2(\b[38] ), .Z(new_n613_));
  NOR2_X1    g228(.A1(new_n613_), .A2(new_n612_), .ZN(new_n614_));
  XOR2_X1    g229(.A1(new_n611_), .A2(new_n614_), .Z(\f[38] ));
  INV_X1     g230(.I(new_n612_), .ZN(new_n616_));
  AOI21_X1   g231(.A1(new_n611_), .A2(new_n616_), .B(new_n613_), .ZN(new_n617_));
  NOR2_X1    g232(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n618_));
  INV_X1     g233(.I(new_n618_), .ZN(new_n619_));
  NAND2_X1   g234(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n620_));
  NAND2_X1   g235(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1    g236(.A1(new_n617_), .A2(new_n621_), .Z(\f[39] ));
  OAI21_X1   g237(.A1(new_n617_), .A2(new_n618_), .B(new_n620_), .ZN(new_n623_));
  NOR2_X1    g238(.A1(\a[40] ), .A2(\b[40] ), .ZN(new_n624_));
  AND2_X2    g239(.A1(\a[40] ), .A2(\b[40] ), .Z(new_n625_));
  NOR2_X1    g240(.A1(new_n625_), .A2(new_n624_), .ZN(new_n626_));
  XOR2_X1    g241(.A1(new_n623_), .A2(new_n626_), .Z(\f[40] ));
  INV_X1     g242(.I(new_n624_), .ZN(new_n628_));
  AOI21_X1   g243(.A1(new_n623_), .A2(new_n628_), .B(new_n625_), .ZN(new_n629_));
  NOR2_X1    g244(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n630_));
  INV_X1     g245(.I(new_n630_), .ZN(new_n631_));
  NAND2_X1   g246(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n632_));
  NAND2_X1   g247(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1    g248(.A1(new_n629_), .A2(new_n633_), .Z(\f[41] ));
  OAI21_X1   g249(.A1(new_n629_), .A2(new_n630_), .B(new_n632_), .ZN(new_n635_));
  NOR2_X1    g250(.A1(\a[42] ), .A2(\b[42] ), .ZN(new_n636_));
  AND2_X2    g251(.A1(\a[42] ), .A2(\b[42] ), .Z(new_n637_));
  NOR2_X1    g252(.A1(new_n637_), .A2(new_n636_), .ZN(new_n638_));
  XOR2_X1    g253(.A1(new_n635_), .A2(new_n638_), .Z(\f[42] ));
  INV_X1     g254(.I(new_n636_), .ZN(new_n640_));
  AOI21_X1   g255(.A1(new_n635_), .A2(new_n640_), .B(new_n637_), .ZN(new_n641_));
  NOR2_X1    g256(.A1(\a[43] ), .A2(\b[43] ), .ZN(new_n642_));
  INV_X1     g257(.I(new_n642_), .ZN(new_n643_));
  NAND2_X1   g258(.A1(\a[43] ), .A2(\b[43] ), .ZN(new_n644_));
  NAND2_X1   g259(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1    g260(.A1(new_n641_), .A2(new_n645_), .Z(\f[43] ));
  OAI21_X1   g261(.A1(new_n641_), .A2(new_n642_), .B(new_n644_), .ZN(new_n647_));
  NOR2_X1    g262(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n648_));
  AND2_X2    g263(.A1(\a[44] ), .A2(\b[44] ), .Z(new_n649_));
  NOR2_X1    g264(.A1(new_n649_), .A2(new_n648_), .ZN(new_n650_));
  XOR2_X1    g265(.A1(new_n647_), .A2(new_n650_), .Z(\f[44] ));
  INV_X1     g266(.I(new_n648_), .ZN(new_n652_));
  AOI21_X1   g267(.A1(new_n647_), .A2(new_n652_), .B(new_n649_), .ZN(new_n653_));
  NOR2_X1    g268(.A1(\a[45] ), .A2(\b[45] ), .ZN(new_n654_));
  INV_X1     g269(.I(new_n654_), .ZN(new_n655_));
  NAND2_X1   g270(.A1(\a[45] ), .A2(\b[45] ), .ZN(new_n656_));
  NAND2_X1   g271(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  XOR2_X1    g272(.A1(new_n653_), .A2(new_n657_), .Z(\f[45] ));
  OAI21_X1   g273(.A1(new_n653_), .A2(new_n654_), .B(new_n656_), .ZN(new_n659_));
  NOR2_X1    g274(.A1(\a[46] ), .A2(\b[46] ), .ZN(new_n660_));
  AND2_X2    g275(.A1(\a[46] ), .A2(\b[46] ), .Z(new_n661_));
  NOR2_X1    g276(.A1(new_n661_), .A2(new_n660_), .ZN(new_n662_));
  XOR2_X1    g277(.A1(new_n659_), .A2(new_n662_), .Z(\f[46] ));
  INV_X1     g278(.I(new_n660_), .ZN(new_n664_));
  AOI21_X1   g279(.A1(new_n659_), .A2(new_n664_), .B(new_n661_), .ZN(new_n665_));
  NOR2_X1    g280(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n666_));
  INV_X1     g281(.I(new_n666_), .ZN(new_n667_));
  NAND2_X1   g282(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n668_));
  NAND2_X1   g283(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  XOR2_X1    g284(.A1(new_n665_), .A2(new_n669_), .Z(\f[47] ));
  OAI21_X1   g285(.A1(new_n665_), .A2(new_n666_), .B(new_n668_), .ZN(new_n671_));
  NOR2_X1    g286(.A1(\a[48] ), .A2(\b[48] ), .ZN(new_n672_));
  AND2_X2    g287(.A1(\a[48] ), .A2(\b[48] ), .Z(new_n673_));
  NOR2_X1    g288(.A1(new_n673_), .A2(new_n672_), .ZN(new_n674_));
  XOR2_X1    g289(.A1(new_n671_), .A2(new_n674_), .Z(\f[48] ));
  INV_X1     g290(.I(new_n672_), .ZN(new_n676_));
  AOI21_X1   g291(.A1(new_n671_), .A2(new_n676_), .B(new_n673_), .ZN(new_n677_));
  NOR2_X1    g292(.A1(\a[49] ), .A2(\b[49] ), .ZN(new_n678_));
  INV_X1     g293(.I(new_n678_), .ZN(new_n679_));
  NAND2_X1   g294(.A1(\a[49] ), .A2(\b[49] ), .ZN(new_n680_));
  NAND2_X1   g295(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  XOR2_X1    g296(.A1(new_n677_), .A2(new_n681_), .Z(\f[49] ));
  OAI21_X1   g297(.A1(new_n677_), .A2(new_n678_), .B(new_n680_), .ZN(new_n683_));
  NOR2_X1    g298(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n684_));
  AND2_X2    g299(.A1(\a[50] ), .A2(\b[50] ), .Z(new_n685_));
  NOR2_X1    g300(.A1(new_n685_), .A2(new_n684_), .ZN(new_n686_));
  XOR2_X1    g301(.A1(new_n683_), .A2(new_n686_), .Z(\f[50] ));
  INV_X1     g302(.I(new_n684_), .ZN(new_n688_));
  AOI21_X1   g303(.A1(new_n683_), .A2(new_n688_), .B(new_n685_), .ZN(new_n689_));
  NOR2_X1    g304(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n690_));
  INV_X1     g305(.I(new_n690_), .ZN(new_n691_));
  NAND2_X1   g306(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n692_));
  NAND2_X1   g307(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XOR2_X1    g308(.A1(new_n689_), .A2(new_n693_), .Z(\f[51] ));
  OAI21_X1   g309(.A1(new_n689_), .A2(new_n690_), .B(new_n692_), .ZN(new_n695_));
  NOR2_X1    g310(.A1(\a[52] ), .A2(\b[52] ), .ZN(new_n696_));
  AND2_X2    g311(.A1(\a[52] ), .A2(\b[52] ), .Z(new_n697_));
  NOR2_X1    g312(.A1(new_n697_), .A2(new_n696_), .ZN(new_n698_));
  XOR2_X1    g313(.A1(new_n695_), .A2(new_n698_), .Z(\f[52] ));
  INV_X1     g314(.I(new_n696_), .ZN(new_n700_));
  AOI21_X1   g315(.A1(new_n695_), .A2(new_n700_), .B(new_n697_), .ZN(new_n701_));
  NOR2_X1    g316(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n702_));
  INV_X1     g317(.I(new_n702_), .ZN(new_n703_));
  NAND2_X1   g318(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n704_));
  NAND2_X1   g319(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  XOR2_X1    g320(.A1(new_n701_), .A2(new_n705_), .Z(\f[53] ));
  OAI21_X1   g321(.A1(new_n701_), .A2(new_n702_), .B(new_n704_), .ZN(new_n707_));
  NOR2_X1    g322(.A1(\a[54] ), .A2(\b[54] ), .ZN(new_n708_));
  AND2_X2    g323(.A1(\a[54] ), .A2(\b[54] ), .Z(new_n709_));
  NOR2_X1    g324(.A1(new_n709_), .A2(new_n708_), .ZN(new_n710_));
  XOR2_X1    g325(.A1(new_n707_), .A2(new_n710_), .Z(\f[54] ));
  INV_X1     g326(.I(new_n708_), .ZN(new_n712_));
  AOI21_X1   g327(.A1(new_n707_), .A2(new_n712_), .B(new_n709_), .ZN(new_n713_));
  NOR2_X1    g328(.A1(\a[55] ), .A2(\b[55] ), .ZN(new_n714_));
  INV_X1     g329(.I(new_n714_), .ZN(new_n715_));
  NAND2_X1   g330(.A1(\a[55] ), .A2(\b[55] ), .ZN(new_n716_));
  NAND2_X1   g331(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  XOR2_X1    g332(.A1(new_n713_), .A2(new_n717_), .Z(\f[55] ));
  OAI21_X1   g333(.A1(new_n713_), .A2(new_n714_), .B(new_n716_), .ZN(new_n719_));
  NOR2_X1    g334(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n720_));
  AND2_X2    g335(.A1(\a[56] ), .A2(\b[56] ), .Z(new_n721_));
  NOR2_X1    g336(.A1(new_n721_), .A2(new_n720_), .ZN(new_n722_));
  XOR2_X1    g337(.A1(new_n719_), .A2(new_n722_), .Z(\f[56] ));
  INV_X1     g338(.I(new_n720_), .ZN(new_n724_));
  AOI21_X1   g339(.A1(new_n719_), .A2(new_n724_), .B(new_n721_), .ZN(new_n725_));
  NOR2_X1    g340(.A1(\a[57] ), .A2(\b[57] ), .ZN(new_n726_));
  INV_X1     g341(.I(new_n726_), .ZN(new_n727_));
  NAND2_X1   g342(.A1(\a[57] ), .A2(\b[57] ), .ZN(new_n728_));
  NAND2_X1   g343(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  XOR2_X1    g344(.A1(new_n725_), .A2(new_n729_), .Z(\f[57] ));
  OAI21_X1   g345(.A1(new_n725_), .A2(new_n726_), .B(new_n728_), .ZN(new_n731_));
  NOR2_X1    g346(.A1(\a[58] ), .A2(\b[58] ), .ZN(new_n732_));
  AND2_X2    g347(.A1(\a[58] ), .A2(\b[58] ), .Z(new_n733_));
  NOR2_X1    g348(.A1(new_n733_), .A2(new_n732_), .ZN(new_n734_));
  XOR2_X1    g349(.A1(new_n731_), .A2(new_n734_), .Z(\f[58] ));
  INV_X1     g350(.I(new_n732_), .ZN(new_n736_));
  AOI21_X1   g351(.A1(new_n731_), .A2(new_n736_), .B(new_n733_), .ZN(new_n737_));
  NOR2_X1    g352(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n738_));
  INV_X1     g353(.I(new_n738_), .ZN(new_n739_));
  NAND2_X1   g354(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n740_));
  NAND2_X1   g355(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XOR2_X1    g356(.A1(new_n737_), .A2(new_n741_), .Z(\f[59] ));
  OAI21_X1   g357(.A1(new_n737_), .A2(new_n738_), .B(new_n740_), .ZN(new_n743_));
  NOR2_X1    g358(.A1(\a[60] ), .A2(\b[60] ), .ZN(new_n744_));
  AND2_X2    g359(.A1(\a[60] ), .A2(\b[60] ), .Z(new_n745_));
  NOR2_X1    g360(.A1(new_n745_), .A2(new_n744_), .ZN(new_n746_));
  XOR2_X1    g361(.A1(new_n743_), .A2(new_n746_), .Z(\f[60] ));
  INV_X1     g362(.I(new_n744_), .ZN(new_n748_));
  AOI21_X1   g363(.A1(new_n743_), .A2(new_n748_), .B(new_n745_), .ZN(new_n749_));
  NOR2_X1    g364(.A1(\a[61] ), .A2(\b[61] ), .ZN(new_n750_));
  INV_X1     g365(.I(new_n750_), .ZN(new_n751_));
  NAND2_X1   g366(.A1(\a[61] ), .A2(\b[61] ), .ZN(new_n752_));
  NAND2_X1   g367(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  XOR2_X1    g368(.A1(new_n749_), .A2(new_n753_), .Z(\f[61] ));
  OAI21_X1   g369(.A1(new_n749_), .A2(new_n750_), .B(new_n752_), .ZN(new_n755_));
  NOR2_X1    g370(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n756_));
  AND2_X2    g371(.A1(\a[62] ), .A2(\b[62] ), .Z(new_n757_));
  NOR2_X1    g372(.A1(new_n757_), .A2(new_n756_), .ZN(new_n758_));
  XOR2_X1    g373(.A1(new_n755_), .A2(new_n758_), .Z(\f[62] ));
  INV_X1     g374(.I(new_n756_), .ZN(new_n760_));
  AOI21_X1   g375(.A1(new_n755_), .A2(new_n760_), .B(new_n757_), .ZN(new_n761_));
  NOR2_X1    g376(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n762_));
  INV_X1     g377(.I(new_n762_), .ZN(new_n763_));
  NAND2_X1   g378(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n764_));
  NAND2_X1   g379(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  XOR2_X1    g380(.A1(new_n761_), .A2(new_n765_), .Z(\f[63] ));
  OAI21_X1   g381(.A1(new_n761_), .A2(new_n762_), .B(new_n764_), .ZN(new_n767_));
  NOR2_X1    g382(.A1(\a[64] ), .A2(\b[64] ), .ZN(new_n768_));
  AND2_X2    g383(.A1(\a[64] ), .A2(\b[64] ), .Z(new_n769_));
  NOR2_X1    g384(.A1(new_n769_), .A2(new_n768_), .ZN(new_n770_));
  XOR2_X1    g385(.A1(new_n767_), .A2(new_n770_), .Z(\f[64] ));
  INV_X1     g386(.I(new_n768_), .ZN(new_n772_));
  AOI21_X1   g387(.A1(new_n767_), .A2(new_n772_), .B(new_n769_), .ZN(new_n773_));
  NOR2_X1    g388(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n774_));
  INV_X1     g389(.I(new_n774_), .ZN(new_n775_));
  NAND2_X1   g390(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n776_));
  NAND2_X1   g391(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  XOR2_X1    g392(.A1(new_n773_), .A2(new_n777_), .Z(\f[65] ));
  OAI21_X1   g393(.A1(new_n773_), .A2(new_n774_), .B(new_n776_), .ZN(new_n779_));
  NOR2_X1    g394(.A1(\a[66] ), .A2(\b[66] ), .ZN(new_n780_));
  AND2_X2    g395(.A1(\a[66] ), .A2(\b[66] ), .Z(new_n781_));
  NOR2_X1    g396(.A1(new_n781_), .A2(new_n780_), .ZN(new_n782_));
  XOR2_X1    g397(.A1(new_n779_), .A2(new_n782_), .Z(\f[66] ));
  INV_X1     g398(.I(new_n780_), .ZN(new_n784_));
  AOI21_X1   g399(.A1(new_n779_), .A2(new_n784_), .B(new_n781_), .ZN(new_n785_));
  NOR2_X1    g400(.A1(\a[67] ), .A2(\b[67] ), .ZN(new_n786_));
  INV_X1     g401(.I(new_n786_), .ZN(new_n787_));
  NAND2_X1   g402(.A1(\a[67] ), .A2(\b[67] ), .ZN(new_n788_));
  NAND2_X1   g403(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  XOR2_X1    g404(.A1(new_n785_), .A2(new_n789_), .Z(\f[67] ));
  OAI21_X1   g405(.A1(new_n785_), .A2(new_n786_), .B(new_n788_), .ZN(new_n791_));
  NOR2_X1    g406(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n792_));
  AND2_X2    g407(.A1(\a[68] ), .A2(\b[68] ), .Z(new_n793_));
  NOR2_X1    g408(.A1(new_n793_), .A2(new_n792_), .ZN(new_n794_));
  XOR2_X1    g409(.A1(new_n791_), .A2(new_n794_), .Z(\f[68] ));
  INV_X1     g410(.I(new_n792_), .ZN(new_n796_));
  AOI21_X1   g411(.A1(new_n791_), .A2(new_n796_), .B(new_n793_), .ZN(new_n797_));
  NOR2_X1    g412(.A1(\a[69] ), .A2(\b[69] ), .ZN(new_n798_));
  INV_X1     g413(.I(new_n798_), .ZN(new_n799_));
  NAND2_X1   g414(.A1(\a[69] ), .A2(\b[69] ), .ZN(new_n800_));
  NAND2_X1   g415(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  XOR2_X1    g416(.A1(new_n797_), .A2(new_n801_), .Z(\f[69] ));
  OAI21_X1   g417(.A1(new_n797_), .A2(new_n798_), .B(new_n800_), .ZN(new_n803_));
  NOR2_X1    g418(.A1(\a[70] ), .A2(\b[70] ), .ZN(new_n804_));
  AND2_X2    g419(.A1(\a[70] ), .A2(\b[70] ), .Z(new_n805_));
  NOR2_X1    g420(.A1(new_n805_), .A2(new_n804_), .ZN(new_n806_));
  XOR2_X1    g421(.A1(new_n803_), .A2(new_n806_), .Z(\f[70] ));
  INV_X1     g422(.I(new_n804_), .ZN(new_n808_));
  AOI21_X1   g423(.A1(new_n803_), .A2(new_n808_), .B(new_n805_), .ZN(new_n809_));
  NOR2_X1    g424(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n810_));
  INV_X1     g425(.I(new_n810_), .ZN(new_n811_));
  NAND2_X1   g426(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n812_));
  NAND2_X1   g427(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  XOR2_X1    g428(.A1(new_n809_), .A2(new_n813_), .Z(\f[71] ));
  OAI21_X1   g429(.A1(new_n809_), .A2(new_n810_), .B(new_n812_), .ZN(new_n815_));
  NOR2_X1    g430(.A1(\a[72] ), .A2(\b[72] ), .ZN(new_n816_));
  AND2_X2    g431(.A1(\a[72] ), .A2(\b[72] ), .Z(new_n817_));
  NOR2_X1    g432(.A1(new_n817_), .A2(new_n816_), .ZN(new_n818_));
  XOR2_X1    g433(.A1(new_n815_), .A2(new_n818_), .Z(\f[72] ));
  INV_X1     g434(.I(new_n816_), .ZN(new_n820_));
  AOI21_X1   g435(.A1(new_n815_), .A2(new_n820_), .B(new_n817_), .ZN(new_n821_));
  NOR2_X1    g436(.A1(\a[73] ), .A2(\b[73] ), .ZN(new_n822_));
  INV_X1     g437(.I(new_n822_), .ZN(new_n823_));
  NAND2_X1   g438(.A1(\a[73] ), .A2(\b[73] ), .ZN(new_n824_));
  NAND2_X1   g439(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  XOR2_X1    g440(.A1(new_n821_), .A2(new_n825_), .Z(\f[73] ));
  OAI21_X1   g441(.A1(new_n821_), .A2(new_n822_), .B(new_n824_), .ZN(new_n827_));
  NOR2_X1    g442(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n828_));
  AND2_X2    g443(.A1(\a[74] ), .A2(\b[74] ), .Z(new_n829_));
  NOR2_X1    g444(.A1(new_n829_), .A2(new_n828_), .ZN(new_n830_));
  XOR2_X1    g445(.A1(new_n827_), .A2(new_n830_), .Z(\f[74] ));
  INV_X1     g446(.I(new_n828_), .ZN(new_n832_));
  AOI21_X1   g447(.A1(new_n827_), .A2(new_n832_), .B(new_n829_), .ZN(new_n833_));
  NOR2_X1    g448(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n834_));
  INV_X1     g449(.I(new_n834_), .ZN(new_n835_));
  NAND2_X1   g450(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n836_));
  NAND2_X1   g451(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  XOR2_X1    g452(.A1(new_n833_), .A2(new_n837_), .Z(\f[75] ));
  OAI21_X1   g453(.A1(new_n833_), .A2(new_n834_), .B(new_n836_), .ZN(new_n839_));
  NOR2_X1    g454(.A1(\a[76] ), .A2(\b[76] ), .ZN(new_n840_));
  AND2_X2    g455(.A1(\a[76] ), .A2(\b[76] ), .Z(new_n841_));
  NOR2_X1    g456(.A1(new_n841_), .A2(new_n840_), .ZN(new_n842_));
  XOR2_X1    g457(.A1(new_n839_), .A2(new_n842_), .Z(\f[76] ));
  INV_X1     g458(.I(new_n840_), .ZN(new_n844_));
  AOI21_X1   g459(.A1(new_n839_), .A2(new_n844_), .B(new_n841_), .ZN(new_n845_));
  NOR2_X1    g460(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n846_));
  INV_X1     g461(.I(new_n846_), .ZN(new_n847_));
  NAND2_X1   g462(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n848_));
  NAND2_X1   g463(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  XOR2_X1    g464(.A1(new_n845_), .A2(new_n849_), .Z(\f[77] ));
  OAI21_X1   g465(.A1(new_n845_), .A2(new_n846_), .B(new_n848_), .ZN(new_n851_));
  NOR2_X1    g466(.A1(\a[78] ), .A2(\b[78] ), .ZN(new_n852_));
  AND2_X2    g467(.A1(\a[78] ), .A2(\b[78] ), .Z(new_n853_));
  NOR2_X1    g468(.A1(new_n853_), .A2(new_n852_), .ZN(new_n854_));
  XOR2_X1    g469(.A1(new_n851_), .A2(new_n854_), .Z(\f[78] ));
  INV_X1     g470(.I(new_n852_), .ZN(new_n856_));
  AOI21_X1   g471(.A1(new_n851_), .A2(new_n856_), .B(new_n853_), .ZN(new_n857_));
  NOR2_X1    g472(.A1(\a[79] ), .A2(\b[79] ), .ZN(new_n858_));
  INV_X1     g473(.I(new_n858_), .ZN(new_n859_));
  NAND2_X1   g474(.A1(\a[79] ), .A2(\b[79] ), .ZN(new_n860_));
  NAND2_X1   g475(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  XOR2_X1    g476(.A1(new_n857_), .A2(new_n861_), .Z(\f[79] ));
  OAI21_X1   g477(.A1(new_n857_), .A2(new_n858_), .B(new_n860_), .ZN(new_n863_));
  NOR2_X1    g478(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n864_));
  AND2_X2    g479(.A1(\a[80] ), .A2(\b[80] ), .Z(new_n865_));
  NOR2_X1    g480(.A1(new_n865_), .A2(new_n864_), .ZN(new_n866_));
  XOR2_X1    g481(.A1(new_n863_), .A2(new_n866_), .Z(\f[80] ));
  INV_X1     g482(.I(new_n864_), .ZN(new_n868_));
  AOI21_X1   g483(.A1(new_n863_), .A2(new_n868_), .B(new_n865_), .ZN(new_n869_));
  NOR2_X1    g484(.A1(\a[81] ), .A2(\b[81] ), .ZN(new_n870_));
  INV_X1     g485(.I(new_n870_), .ZN(new_n871_));
  NAND2_X1   g486(.A1(\a[81] ), .A2(\b[81] ), .ZN(new_n872_));
  NAND2_X1   g487(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  XOR2_X1    g488(.A1(new_n869_), .A2(new_n873_), .Z(\f[81] ));
  OAI21_X1   g489(.A1(new_n869_), .A2(new_n870_), .B(new_n872_), .ZN(new_n875_));
  NOR2_X1    g490(.A1(\a[82] ), .A2(\b[82] ), .ZN(new_n876_));
  AND2_X2    g491(.A1(\a[82] ), .A2(\b[82] ), .Z(new_n877_));
  NOR2_X1    g492(.A1(new_n877_), .A2(new_n876_), .ZN(new_n878_));
  XOR2_X1    g493(.A1(new_n875_), .A2(new_n878_), .Z(\f[82] ));
  INV_X1     g494(.I(new_n876_), .ZN(new_n880_));
  AOI21_X1   g495(.A1(new_n875_), .A2(new_n880_), .B(new_n877_), .ZN(new_n881_));
  NOR2_X1    g496(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n882_));
  INV_X1     g497(.I(new_n882_), .ZN(new_n883_));
  NAND2_X1   g498(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n884_));
  NAND2_X1   g499(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  XOR2_X1    g500(.A1(new_n881_), .A2(new_n885_), .Z(\f[83] ));
  OAI21_X1   g501(.A1(new_n881_), .A2(new_n882_), .B(new_n884_), .ZN(new_n887_));
  NOR2_X1    g502(.A1(\a[84] ), .A2(\b[84] ), .ZN(new_n888_));
  AND2_X2    g503(.A1(\a[84] ), .A2(\b[84] ), .Z(new_n889_));
  NOR2_X1    g504(.A1(new_n889_), .A2(new_n888_), .ZN(new_n890_));
  XOR2_X1    g505(.A1(new_n887_), .A2(new_n890_), .Z(\f[84] ));
  INV_X1     g506(.I(new_n888_), .ZN(new_n892_));
  AOI21_X1   g507(.A1(new_n887_), .A2(new_n892_), .B(new_n889_), .ZN(new_n893_));
  NOR2_X1    g508(.A1(\a[85] ), .A2(\b[85] ), .ZN(new_n894_));
  INV_X1     g509(.I(new_n894_), .ZN(new_n895_));
  NAND2_X1   g510(.A1(\a[85] ), .A2(\b[85] ), .ZN(new_n896_));
  NAND2_X1   g511(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  XOR2_X1    g512(.A1(new_n893_), .A2(new_n897_), .Z(\f[85] ));
  OAI21_X1   g513(.A1(new_n893_), .A2(new_n894_), .B(new_n896_), .ZN(new_n899_));
  NOR2_X1    g514(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n900_));
  AND2_X2    g515(.A1(\a[86] ), .A2(\b[86] ), .Z(new_n901_));
  NOR2_X1    g516(.A1(new_n901_), .A2(new_n900_), .ZN(new_n902_));
  XOR2_X1    g517(.A1(new_n899_), .A2(new_n902_), .Z(\f[86] ));
  INV_X1     g518(.I(new_n900_), .ZN(new_n904_));
  AOI21_X1   g519(.A1(new_n899_), .A2(new_n904_), .B(new_n901_), .ZN(new_n905_));
  NOR2_X1    g520(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n906_));
  INV_X1     g521(.I(new_n906_), .ZN(new_n907_));
  NAND2_X1   g522(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n908_));
  NAND2_X1   g523(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  XOR2_X1    g524(.A1(new_n905_), .A2(new_n909_), .Z(\f[87] ));
  OAI21_X1   g525(.A1(new_n905_), .A2(new_n906_), .B(new_n908_), .ZN(new_n911_));
  NOR2_X1    g526(.A1(\a[88] ), .A2(\b[88] ), .ZN(new_n912_));
  AND2_X2    g527(.A1(\a[88] ), .A2(\b[88] ), .Z(new_n913_));
  NOR2_X1    g528(.A1(new_n913_), .A2(new_n912_), .ZN(new_n914_));
  XOR2_X1    g529(.A1(new_n911_), .A2(new_n914_), .Z(\f[88] ));
  INV_X1     g530(.I(new_n912_), .ZN(new_n916_));
  AOI21_X1   g531(.A1(new_n911_), .A2(new_n916_), .B(new_n913_), .ZN(new_n917_));
  NOR2_X1    g532(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n918_));
  INV_X1     g533(.I(new_n918_), .ZN(new_n919_));
  NAND2_X1   g534(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n920_));
  NAND2_X1   g535(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  XOR2_X1    g536(.A1(new_n917_), .A2(new_n921_), .Z(\f[89] ));
  OAI21_X1   g537(.A1(new_n917_), .A2(new_n918_), .B(new_n920_), .ZN(new_n923_));
  NOR2_X1    g538(.A1(\a[90] ), .A2(\b[90] ), .ZN(new_n924_));
  AND2_X2    g539(.A1(\a[90] ), .A2(\b[90] ), .Z(new_n925_));
  NOR2_X1    g540(.A1(new_n925_), .A2(new_n924_), .ZN(new_n926_));
  XOR2_X1    g541(.A1(new_n923_), .A2(new_n926_), .Z(\f[90] ));
  INV_X1     g542(.I(new_n924_), .ZN(new_n928_));
  AOI21_X1   g543(.A1(new_n923_), .A2(new_n928_), .B(new_n925_), .ZN(new_n929_));
  NOR2_X1    g544(.A1(\a[91] ), .A2(\b[91] ), .ZN(new_n930_));
  INV_X1     g545(.I(new_n930_), .ZN(new_n931_));
  NAND2_X1   g546(.A1(\a[91] ), .A2(\b[91] ), .ZN(new_n932_));
  NAND2_X1   g547(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  XOR2_X1    g548(.A1(new_n929_), .A2(new_n933_), .Z(\f[91] ));
  OAI21_X1   g549(.A1(new_n929_), .A2(new_n930_), .B(new_n932_), .ZN(new_n935_));
  NOR2_X1    g550(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n936_));
  AND2_X2    g551(.A1(\a[92] ), .A2(\b[92] ), .Z(new_n937_));
  NOR2_X1    g552(.A1(new_n937_), .A2(new_n936_), .ZN(new_n938_));
  XOR2_X1    g553(.A1(new_n935_), .A2(new_n938_), .Z(\f[92] ));
  INV_X1     g554(.I(new_n936_), .ZN(new_n940_));
  AOI21_X1   g555(.A1(new_n935_), .A2(new_n940_), .B(new_n937_), .ZN(new_n941_));
  NOR2_X1    g556(.A1(\a[93] ), .A2(\b[93] ), .ZN(new_n942_));
  INV_X1     g557(.I(new_n942_), .ZN(new_n943_));
  NAND2_X1   g558(.A1(\a[93] ), .A2(\b[93] ), .ZN(new_n944_));
  NAND2_X1   g559(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  XOR2_X1    g560(.A1(new_n941_), .A2(new_n945_), .Z(\f[93] ));
  OAI21_X1   g561(.A1(new_n941_), .A2(new_n942_), .B(new_n944_), .ZN(new_n947_));
  NOR2_X1    g562(.A1(\a[94] ), .A2(\b[94] ), .ZN(new_n948_));
  AND2_X2    g563(.A1(\a[94] ), .A2(\b[94] ), .Z(new_n949_));
  NOR2_X1    g564(.A1(new_n949_), .A2(new_n948_), .ZN(new_n950_));
  XOR2_X1    g565(.A1(new_n947_), .A2(new_n950_), .Z(\f[94] ));
  INV_X1     g566(.I(new_n948_), .ZN(new_n952_));
  AOI21_X1   g567(.A1(new_n947_), .A2(new_n952_), .B(new_n949_), .ZN(new_n953_));
  NOR2_X1    g568(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n954_));
  INV_X1     g569(.I(new_n954_), .ZN(new_n955_));
  NAND2_X1   g570(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n956_));
  NAND2_X1   g571(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  XOR2_X1    g572(.A1(new_n953_), .A2(new_n957_), .Z(\f[95] ));
  OAI21_X1   g573(.A1(new_n953_), .A2(new_n954_), .B(new_n956_), .ZN(new_n959_));
  NOR2_X1    g574(.A1(\a[96] ), .A2(\b[96] ), .ZN(new_n960_));
  AND2_X2    g575(.A1(\a[96] ), .A2(\b[96] ), .Z(new_n961_));
  NOR2_X1    g576(.A1(new_n961_), .A2(new_n960_), .ZN(new_n962_));
  XOR2_X1    g577(.A1(new_n959_), .A2(new_n962_), .Z(\f[96] ));
  INV_X1     g578(.I(new_n960_), .ZN(new_n964_));
  AOI21_X1   g579(.A1(new_n959_), .A2(new_n964_), .B(new_n961_), .ZN(new_n965_));
  NOR2_X1    g580(.A1(\a[97] ), .A2(\b[97] ), .ZN(new_n966_));
  INV_X1     g581(.I(new_n966_), .ZN(new_n967_));
  NAND2_X1   g582(.A1(\a[97] ), .A2(\b[97] ), .ZN(new_n968_));
  NAND2_X1   g583(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  XOR2_X1    g584(.A1(new_n965_), .A2(new_n969_), .Z(\f[97] ));
  OAI21_X1   g585(.A1(new_n965_), .A2(new_n966_), .B(new_n968_), .ZN(new_n971_));
  NOR2_X1    g586(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n972_));
  AND2_X2    g587(.A1(\a[98] ), .A2(\b[98] ), .Z(new_n973_));
  NOR2_X1    g588(.A1(new_n973_), .A2(new_n972_), .ZN(new_n974_));
  XOR2_X1    g589(.A1(new_n971_), .A2(new_n974_), .Z(\f[98] ));
  INV_X1     g590(.I(new_n972_), .ZN(new_n976_));
  AOI21_X1   g591(.A1(new_n971_), .A2(new_n976_), .B(new_n973_), .ZN(new_n977_));
  NOR2_X1    g592(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n978_));
  INV_X1     g593(.I(new_n978_), .ZN(new_n979_));
  NAND2_X1   g594(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n980_));
  NAND2_X1   g595(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  XOR2_X1    g596(.A1(new_n977_), .A2(new_n981_), .Z(\f[99] ));
  OAI21_X1   g597(.A1(new_n977_), .A2(new_n978_), .B(new_n980_), .ZN(new_n983_));
  NOR2_X1    g598(.A1(\a[100] ), .A2(\b[100] ), .ZN(new_n984_));
  AND2_X2    g599(.A1(\a[100] ), .A2(\b[100] ), .Z(new_n985_));
  NOR2_X1    g600(.A1(new_n985_), .A2(new_n984_), .ZN(new_n986_));
  XOR2_X1    g601(.A1(new_n983_), .A2(new_n986_), .Z(\f[100] ));
  INV_X1     g602(.I(new_n984_), .ZN(new_n988_));
  AOI21_X1   g603(.A1(new_n983_), .A2(new_n988_), .B(new_n985_), .ZN(new_n989_));
  NOR2_X1    g604(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n990_));
  INV_X1     g605(.I(new_n990_), .ZN(new_n991_));
  NAND2_X1   g606(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n992_));
  NAND2_X1   g607(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  XOR2_X1    g608(.A1(new_n989_), .A2(new_n993_), .Z(\f[101] ));
  OAI21_X1   g609(.A1(new_n989_), .A2(new_n990_), .B(new_n992_), .ZN(new_n995_));
  NOR2_X1    g610(.A1(\a[102] ), .A2(\b[102] ), .ZN(new_n996_));
  AND2_X2    g611(.A1(\a[102] ), .A2(\b[102] ), .Z(new_n997_));
  NOR2_X1    g612(.A1(new_n997_), .A2(new_n996_), .ZN(new_n998_));
  XOR2_X1    g613(.A1(new_n995_), .A2(new_n998_), .Z(\f[102] ));
  INV_X1     g614(.I(new_n996_), .ZN(new_n1000_));
  AOI21_X1   g615(.A1(new_n995_), .A2(new_n1000_), .B(new_n997_), .ZN(new_n1001_));
  NOR2_X1    g616(.A1(\a[103] ), .A2(\b[103] ), .ZN(new_n1002_));
  INV_X1     g617(.I(new_n1002_), .ZN(new_n1003_));
  NAND2_X1   g618(.A1(\a[103] ), .A2(\b[103] ), .ZN(new_n1004_));
  NAND2_X1   g619(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1005_));
  XOR2_X1    g620(.A1(new_n1001_), .A2(new_n1005_), .Z(\f[103] ));
  OAI21_X1   g621(.A1(new_n1001_), .A2(new_n1002_), .B(new_n1004_), .ZN(new_n1007_));
  NOR2_X1    g622(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1008_));
  AND2_X2    g623(.A1(\a[104] ), .A2(\b[104] ), .Z(new_n1009_));
  NOR2_X1    g624(.A1(new_n1009_), .A2(new_n1008_), .ZN(new_n1010_));
  XOR2_X1    g625(.A1(new_n1007_), .A2(new_n1010_), .Z(\f[104] ));
  INV_X1     g626(.I(new_n1008_), .ZN(new_n1012_));
  AOI21_X1   g627(.A1(new_n1007_), .A2(new_n1012_), .B(new_n1009_), .ZN(new_n1013_));
  NOR2_X1    g628(.A1(\a[105] ), .A2(\b[105] ), .ZN(new_n1014_));
  INV_X1     g629(.I(new_n1014_), .ZN(new_n1015_));
  NAND2_X1   g630(.A1(\a[105] ), .A2(\b[105] ), .ZN(new_n1016_));
  NAND2_X1   g631(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  XOR2_X1    g632(.A1(new_n1013_), .A2(new_n1017_), .Z(\f[105] ));
  OAI21_X1   g633(.A1(new_n1013_), .A2(new_n1014_), .B(new_n1016_), .ZN(new_n1019_));
  NOR2_X1    g634(.A1(\a[106] ), .A2(\b[106] ), .ZN(new_n1020_));
  AND2_X2    g635(.A1(\a[106] ), .A2(\b[106] ), .Z(new_n1021_));
  NOR2_X1    g636(.A1(new_n1021_), .A2(new_n1020_), .ZN(new_n1022_));
  XOR2_X1    g637(.A1(new_n1019_), .A2(new_n1022_), .Z(\f[106] ));
  INV_X1     g638(.I(new_n1020_), .ZN(new_n1024_));
  AOI21_X1   g639(.A1(new_n1019_), .A2(new_n1024_), .B(new_n1021_), .ZN(new_n1025_));
  NOR2_X1    g640(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1026_));
  INV_X1     g641(.I(new_n1026_), .ZN(new_n1027_));
  NAND2_X1   g642(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1028_));
  NAND2_X1   g643(.A1(new_n1027_), .A2(new_n1028_), .ZN(new_n1029_));
  XOR2_X1    g644(.A1(new_n1025_), .A2(new_n1029_), .Z(\f[107] ));
  OAI21_X1   g645(.A1(new_n1025_), .A2(new_n1026_), .B(new_n1028_), .ZN(new_n1031_));
  NOR2_X1    g646(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1032_));
  AND2_X2    g647(.A1(\a[108] ), .A2(\b[108] ), .Z(new_n1033_));
  NOR2_X1    g648(.A1(new_n1033_), .A2(new_n1032_), .ZN(new_n1034_));
  XOR2_X1    g649(.A1(new_n1031_), .A2(new_n1034_), .Z(\f[108] ));
  INV_X1     g650(.I(new_n1032_), .ZN(new_n1036_));
  AOI21_X1   g651(.A1(new_n1031_), .A2(new_n1036_), .B(new_n1033_), .ZN(new_n1037_));
  NOR2_X1    g652(.A1(\a[109] ), .A2(\b[109] ), .ZN(new_n1038_));
  INV_X1     g653(.I(new_n1038_), .ZN(new_n1039_));
  NAND2_X1   g654(.A1(\a[109] ), .A2(\b[109] ), .ZN(new_n1040_));
  NAND2_X1   g655(.A1(new_n1039_), .A2(new_n1040_), .ZN(new_n1041_));
  XOR2_X1    g656(.A1(new_n1037_), .A2(new_n1041_), .Z(\f[109] ));
  OAI21_X1   g657(.A1(new_n1037_), .A2(new_n1038_), .B(new_n1040_), .ZN(new_n1043_));
  NOR2_X1    g658(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1044_));
  AND2_X2    g659(.A1(\a[110] ), .A2(\b[110] ), .Z(new_n1045_));
  NOR2_X1    g660(.A1(new_n1045_), .A2(new_n1044_), .ZN(new_n1046_));
  XOR2_X1    g661(.A1(new_n1043_), .A2(new_n1046_), .Z(\f[110] ));
  INV_X1     g662(.I(new_n1044_), .ZN(new_n1048_));
  AOI21_X1   g663(.A1(new_n1043_), .A2(new_n1048_), .B(new_n1045_), .ZN(new_n1049_));
  NOR2_X1    g664(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1050_));
  INV_X1     g665(.I(new_n1050_), .ZN(new_n1051_));
  NAND2_X1   g666(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1052_));
  NAND2_X1   g667(.A1(new_n1051_), .A2(new_n1052_), .ZN(new_n1053_));
  XOR2_X1    g668(.A1(new_n1049_), .A2(new_n1053_), .Z(\f[111] ));
  OAI21_X1   g669(.A1(new_n1049_), .A2(new_n1050_), .B(new_n1052_), .ZN(new_n1055_));
  NOR2_X1    g670(.A1(\a[112] ), .A2(\b[112] ), .ZN(new_n1056_));
  AND2_X2    g671(.A1(\a[112] ), .A2(\b[112] ), .Z(new_n1057_));
  NOR2_X1    g672(.A1(new_n1057_), .A2(new_n1056_), .ZN(new_n1058_));
  XOR2_X1    g673(.A1(new_n1055_), .A2(new_n1058_), .Z(\f[112] ));
  INV_X1     g674(.I(new_n1056_), .ZN(new_n1060_));
  AOI21_X1   g675(.A1(new_n1055_), .A2(new_n1060_), .B(new_n1057_), .ZN(new_n1061_));
  NOR2_X1    g676(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1062_));
  INV_X1     g677(.I(new_n1062_), .ZN(new_n1063_));
  NAND2_X1   g678(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1064_));
  NAND2_X1   g679(.A1(new_n1063_), .A2(new_n1064_), .ZN(new_n1065_));
  XOR2_X1    g680(.A1(new_n1061_), .A2(new_n1065_), .Z(\f[113] ));
  OAI21_X1   g681(.A1(new_n1061_), .A2(new_n1062_), .B(new_n1064_), .ZN(new_n1067_));
  NOR2_X1    g682(.A1(\a[114] ), .A2(\b[114] ), .ZN(new_n1068_));
  AND2_X2    g683(.A1(\a[114] ), .A2(\b[114] ), .Z(new_n1069_));
  NOR2_X1    g684(.A1(new_n1069_), .A2(new_n1068_), .ZN(new_n1070_));
  XOR2_X1    g685(.A1(new_n1067_), .A2(new_n1070_), .Z(\f[114] ));
  INV_X1     g686(.I(new_n1068_), .ZN(new_n1072_));
  AOI21_X1   g687(.A1(new_n1067_), .A2(new_n1072_), .B(new_n1069_), .ZN(new_n1073_));
  NOR2_X1    g688(.A1(\a[115] ), .A2(\b[115] ), .ZN(new_n1074_));
  INV_X1     g689(.I(new_n1074_), .ZN(new_n1075_));
  NAND2_X1   g690(.A1(\a[115] ), .A2(\b[115] ), .ZN(new_n1076_));
  NAND2_X1   g691(.A1(new_n1075_), .A2(new_n1076_), .ZN(new_n1077_));
  XOR2_X1    g692(.A1(new_n1073_), .A2(new_n1077_), .Z(\f[115] ));
  OAI21_X1   g693(.A1(new_n1073_), .A2(new_n1074_), .B(new_n1076_), .ZN(new_n1079_));
  NOR2_X1    g694(.A1(\a[116] ), .A2(\b[116] ), .ZN(new_n1080_));
  AND2_X2    g695(.A1(\a[116] ), .A2(\b[116] ), .Z(new_n1081_));
  NOR2_X1    g696(.A1(new_n1081_), .A2(new_n1080_), .ZN(new_n1082_));
  XOR2_X1    g697(.A1(new_n1079_), .A2(new_n1082_), .Z(\f[116] ));
  INV_X1     g698(.I(new_n1080_), .ZN(new_n1084_));
  AOI21_X1   g699(.A1(new_n1079_), .A2(new_n1084_), .B(new_n1081_), .ZN(new_n1085_));
  NOR2_X1    g700(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1086_));
  INV_X1     g701(.I(new_n1086_), .ZN(new_n1087_));
  NAND2_X1   g702(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1088_));
  NAND2_X1   g703(.A1(new_n1087_), .A2(new_n1088_), .ZN(new_n1089_));
  XOR2_X1    g704(.A1(new_n1085_), .A2(new_n1089_), .Z(\f[117] ));
  OAI21_X1   g705(.A1(new_n1085_), .A2(new_n1086_), .B(new_n1088_), .ZN(new_n1091_));
  NOR2_X1    g706(.A1(\a[118] ), .A2(\b[118] ), .ZN(new_n1092_));
  AND2_X2    g707(.A1(\a[118] ), .A2(\b[118] ), .Z(new_n1093_));
  NOR2_X1    g708(.A1(new_n1093_), .A2(new_n1092_), .ZN(new_n1094_));
  XOR2_X1    g709(.A1(new_n1091_), .A2(new_n1094_), .Z(\f[118] ));
  INV_X1     g710(.I(new_n1092_), .ZN(new_n1096_));
  AOI21_X1   g711(.A1(new_n1091_), .A2(new_n1096_), .B(new_n1093_), .ZN(new_n1097_));
  NOR2_X1    g712(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1098_));
  INV_X1     g713(.I(new_n1098_), .ZN(new_n1099_));
  NAND2_X1   g714(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1100_));
  NAND2_X1   g715(.A1(new_n1099_), .A2(new_n1100_), .ZN(new_n1101_));
  XOR2_X1    g716(.A1(new_n1097_), .A2(new_n1101_), .Z(\f[119] ));
  OAI21_X1   g717(.A1(new_n1097_), .A2(new_n1098_), .B(new_n1100_), .ZN(new_n1103_));
  NOR2_X1    g718(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1104_));
  AND2_X2    g719(.A1(\a[120] ), .A2(\b[120] ), .Z(new_n1105_));
  NOR2_X1    g720(.A1(new_n1105_), .A2(new_n1104_), .ZN(new_n1106_));
  XOR2_X1    g721(.A1(new_n1103_), .A2(new_n1106_), .Z(\f[120] ));
  INV_X1     g722(.I(new_n1104_), .ZN(new_n1108_));
  AOI21_X1   g723(.A1(new_n1103_), .A2(new_n1108_), .B(new_n1105_), .ZN(new_n1109_));
  NOR2_X1    g724(.A1(\a[121] ), .A2(\b[121] ), .ZN(new_n1110_));
  INV_X1     g725(.I(new_n1110_), .ZN(new_n1111_));
  NAND2_X1   g726(.A1(\a[121] ), .A2(\b[121] ), .ZN(new_n1112_));
  NAND2_X1   g727(.A1(new_n1111_), .A2(new_n1112_), .ZN(new_n1113_));
  XOR2_X1    g728(.A1(new_n1109_), .A2(new_n1113_), .Z(\f[121] ));
  OAI21_X1   g729(.A1(new_n1109_), .A2(new_n1110_), .B(new_n1112_), .ZN(new_n1115_));
  NOR2_X1    g730(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1116_));
  AND2_X2    g731(.A1(\a[122] ), .A2(\b[122] ), .Z(new_n1117_));
  NOR2_X1    g732(.A1(new_n1117_), .A2(new_n1116_), .ZN(new_n1118_));
  XOR2_X1    g733(.A1(new_n1115_), .A2(new_n1118_), .Z(\f[122] ));
  INV_X1     g734(.I(new_n1116_), .ZN(new_n1120_));
  AOI21_X1   g735(.A1(new_n1115_), .A2(new_n1120_), .B(new_n1117_), .ZN(new_n1121_));
  NOR2_X1    g736(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1122_));
  INV_X1     g737(.I(new_n1122_), .ZN(new_n1123_));
  NAND2_X1   g738(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1124_));
  NAND2_X1   g739(.A1(new_n1123_), .A2(new_n1124_), .ZN(new_n1125_));
  XOR2_X1    g740(.A1(new_n1121_), .A2(new_n1125_), .Z(\f[123] ));
  OAI21_X1   g741(.A1(new_n1121_), .A2(new_n1122_), .B(new_n1124_), .ZN(new_n1127_));
  NOR2_X1    g742(.A1(\a[124] ), .A2(\b[124] ), .ZN(new_n1128_));
  AND2_X2    g743(.A1(\a[124] ), .A2(\b[124] ), .Z(new_n1129_));
  NOR2_X1    g744(.A1(new_n1129_), .A2(new_n1128_), .ZN(new_n1130_));
  XOR2_X1    g745(.A1(new_n1127_), .A2(new_n1130_), .Z(\f[124] ));
  INV_X1     g746(.I(new_n1128_), .ZN(new_n1132_));
  AOI21_X1   g747(.A1(new_n1127_), .A2(new_n1132_), .B(new_n1129_), .ZN(new_n1133_));
  NOR2_X1    g748(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1134_));
  INV_X1     g749(.I(new_n1134_), .ZN(new_n1135_));
  NAND2_X1   g750(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1136_));
  NAND2_X1   g751(.A1(new_n1135_), .A2(new_n1136_), .ZN(new_n1137_));
  XOR2_X1    g752(.A1(new_n1133_), .A2(new_n1137_), .Z(\f[125] ));
  OAI21_X1   g753(.A1(new_n1133_), .A2(new_n1134_), .B(new_n1136_), .ZN(new_n1139_));
  NOR2_X1    g754(.A1(\a[126] ), .A2(\b[126] ), .ZN(new_n1140_));
  AND2_X2    g755(.A1(\a[126] ), .A2(\b[126] ), .Z(new_n1141_));
  NOR2_X1    g756(.A1(new_n1141_), .A2(new_n1140_), .ZN(new_n1142_));
  XOR2_X1    g757(.A1(new_n1139_), .A2(new_n1142_), .Z(\f[126] ));
  INV_X1     g758(.I(new_n1140_), .ZN(new_n1144_));
  AOI21_X1   g759(.A1(new_n1139_), .A2(new_n1144_), .B(new_n1141_), .ZN(new_n1145_));
  NOR2_X1    g760(.A1(\a[127] ), .A2(\b[127] ), .ZN(new_n1146_));
  INV_X1     g761(.I(new_n1146_), .ZN(new_n1147_));
  NAND2_X1   g762(.A1(\a[127] ), .A2(\b[127] ), .ZN(new_n1148_));
  NAND2_X1   g763(.A1(new_n1147_), .A2(new_n1148_), .ZN(new_n1149_));
  XOR2_X1    g764(.A1(new_n1145_), .A2(new_n1149_), .Z(\f[127] ));
  OAI21_X1   g765(.A1(new_n1145_), .A2(new_n1146_), .B(new_n1148_), .ZN(cOut));
endmodule


