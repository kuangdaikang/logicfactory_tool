// Benchmark "multiplier" written by ABC on Thu Sep 14 20:20:10 2023

module multiplier ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257_, new_n258_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_,
    new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_,
    new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_,
    new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3735_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_,
    new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_,
    new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_,
    new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_,
    new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_,
    new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_,
    new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_,
    new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_,
    new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_,
    new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_,
    new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_,
    new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_,
    new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_,
    new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_,
    new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_,
    new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_,
    new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4265_, new_n4266_, new_n4267_, new_n4268_,
    new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_,
    new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_,
    new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_,
    new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_,
    new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_,
    new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_,
    new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_,
    new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_,
    new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_,
    new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_,
    new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_,
    new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_,
    new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_,
    new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_,
    new_n4353_, new_n4354_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_,
    new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_,
    new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_,
    new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_,
    new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_,
    new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_,
    new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_,
    new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_,
    new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_,
    new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_,
    new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_,
    new_n4505_, new_n4506_, new_n4507_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4792_, new_n4793_, new_n4794_,
    new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_,
    new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_,
    new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_,
    new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_,
    new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_,
    new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_,
    new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_,
    new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_,
    new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_,
    new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_,
    new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_,
    new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_,
    new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_,
    new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_,
    new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_,
    new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_,
    new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_,
    new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_,
    new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_,
    new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_,
    new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5216_,
    new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_,
    new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_,
    new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_,
    new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_,
    new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_,
    new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_,
    new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_,
    new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_,
    new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_,
    new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_,
    new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_,
    new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_,
    new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_,
    new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_,
    new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_,
    new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_,
    new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_,
    new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_,
    new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_,
    new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_,
    new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_,
    new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_,
    new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_,
    new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_,
    new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_,
    new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_,
    new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_,
    new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_,
    new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_,
    new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_,
    new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_,
    new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_,
    new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_,
    new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_,
    new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_,
    new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_,
    new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_,
    new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_,
    new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_,
    new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_,
    new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_,
    new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_,
    new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_,
    new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_,
    new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_,
    new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_,
    new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_,
    new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_,
    new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_,
    new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_,
    new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_,
    new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_,
    new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_,
    new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_,
    new_n7127_, new_n7128_, new_n7129_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_,
    new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_,
    new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_,
    new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_,
    new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_,
    new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_,
    new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_,
    new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_,
    new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_,
    new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_,
    new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_,
    new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_,
    new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_,
    new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_,
    new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_,
    new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_,
    new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_,
    new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_,
    new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_,
    new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_,
    new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_,
    new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_,
    new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_,
    new_n7983_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_,
    new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_,
    new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_,
    new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_,
    new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_,
    new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_,
    new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_,
    new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_,
    new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_,
    new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_,
    new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_,
    new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_,
    new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_,
    new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_,
    new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_,
    new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_,
    new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_,
    new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_,
    new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_,
    new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_,
    new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_,
    new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_,
    new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_,
    new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_,
    new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_,
    new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_,
    new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_,
    new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_,
    new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_,
    new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_,
    new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_,
    new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_,
    new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_,
    new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_,
    new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_,
    new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_,
    new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_,
    new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_,
    new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_,
    new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_,
    new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_,
    new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_,
    new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_,
    new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_,
    new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_,
    new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_,
    new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_,
    new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_,
    new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_,
    new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_,
    new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_,
    new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_,
    new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_,
    new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_,
    new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_,
    new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_,
    new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_,
    new_n9997_, new_n9998_, new_n9999_, new_n10000_, new_n10001_,
    new_n10002_, new_n10003_, new_n10004_, new_n10005_, new_n10006_,
    new_n10007_, new_n10008_, new_n10009_, new_n10010_, new_n10011_,
    new_n10012_, new_n10013_, new_n10014_, new_n10015_, new_n10016_,
    new_n10017_, new_n10018_, new_n10019_, new_n10020_, new_n10021_,
    new_n10022_, new_n10023_, new_n10024_, new_n10025_, new_n10026_,
    new_n10027_, new_n10028_, new_n10029_, new_n10030_, new_n10031_,
    new_n10032_, new_n10033_, new_n10034_, new_n10035_, new_n10036_,
    new_n10037_, new_n10038_, new_n10039_, new_n10040_, new_n10041_,
    new_n10042_, new_n10043_, new_n10044_, new_n10045_, new_n10046_,
    new_n10047_, new_n10048_, new_n10049_, new_n10050_, new_n10051_,
    new_n10052_, new_n10053_, new_n10054_, new_n10055_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10114_, new_n10115_, new_n10116_, new_n10117_,
    new_n10118_, new_n10119_, new_n10120_, new_n10121_, new_n10122_,
    new_n10123_, new_n10124_, new_n10125_, new_n10126_, new_n10127_,
    new_n10128_, new_n10129_, new_n10130_, new_n10131_, new_n10132_,
    new_n10133_, new_n10134_, new_n10135_, new_n10136_, new_n10137_,
    new_n10138_, new_n10139_, new_n10140_, new_n10141_, new_n10142_,
    new_n10143_, new_n10144_, new_n10145_, new_n10146_, new_n10147_,
    new_n10148_, new_n10149_, new_n10150_, new_n10151_, new_n10152_,
    new_n10153_, new_n10154_, new_n10155_, new_n10156_, new_n10157_,
    new_n10158_, new_n10159_, new_n10160_, new_n10161_, new_n10162_,
    new_n10163_, new_n10164_, new_n10165_, new_n10166_, new_n10167_,
    new_n10168_, new_n10169_, new_n10170_, new_n10171_, new_n10172_,
    new_n10173_, new_n10174_, new_n10175_, new_n10176_, new_n10177_,
    new_n10178_, new_n10179_, new_n10180_, new_n10181_, new_n10182_,
    new_n10183_, new_n10184_, new_n10185_, new_n10186_, new_n10187_,
    new_n10188_, new_n10189_, new_n10190_, new_n10191_, new_n10192_,
    new_n10193_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10200_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10205_, new_n10206_, new_n10207_,
    new_n10208_, new_n10209_, new_n10210_, new_n10211_, new_n10212_,
    new_n10213_, new_n10214_, new_n10215_, new_n10216_, new_n10217_,
    new_n10218_, new_n10219_, new_n10220_, new_n10221_, new_n10222_,
    new_n10223_, new_n10224_, new_n10225_, new_n10226_, new_n10227_,
    new_n10228_, new_n10229_, new_n10230_, new_n10231_, new_n10232_,
    new_n10233_, new_n10234_, new_n10235_, new_n10236_, new_n10237_,
    new_n10238_, new_n10239_, new_n10240_, new_n10241_, new_n10242_,
    new_n10243_, new_n10244_, new_n10245_, new_n10246_, new_n10247_,
    new_n10248_, new_n10249_, new_n10250_, new_n10251_, new_n10252_,
    new_n10253_, new_n10254_, new_n10255_, new_n10256_, new_n10257_,
    new_n10258_, new_n10259_, new_n10260_, new_n10261_, new_n10262_,
    new_n10263_, new_n10264_, new_n10265_, new_n10266_, new_n10267_,
    new_n10268_, new_n10269_, new_n10270_, new_n10271_, new_n10272_,
    new_n10273_, new_n10274_, new_n10275_, new_n10276_, new_n10277_,
    new_n10278_, new_n10279_, new_n10280_, new_n10281_, new_n10282_,
    new_n10283_, new_n10284_, new_n10285_, new_n10286_, new_n10287_,
    new_n10288_, new_n10289_, new_n10290_, new_n10291_, new_n10292_,
    new_n10293_, new_n10294_, new_n10295_, new_n10296_, new_n10297_,
    new_n10298_, new_n10299_, new_n10300_, new_n10301_, new_n10302_,
    new_n10303_, new_n10304_, new_n10305_, new_n10306_, new_n10307_,
    new_n10308_, new_n10309_, new_n10310_, new_n10311_, new_n10312_,
    new_n10313_, new_n10314_, new_n10315_, new_n10316_, new_n10317_,
    new_n10318_, new_n10319_, new_n10320_, new_n10321_, new_n10322_,
    new_n10323_, new_n10324_, new_n10325_, new_n10326_, new_n10327_,
    new_n10328_, new_n10329_, new_n10330_, new_n10331_, new_n10332_,
    new_n10333_, new_n10334_, new_n10335_, new_n10336_, new_n10337_,
    new_n10338_, new_n10339_, new_n10340_, new_n10341_, new_n10342_,
    new_n10343_, new_n10344_, new_n10345_, new_n10346_, new_n10347_,
    new_n10348_, new_n10349_, new_n10350_, new_n10352_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10359_, new_n10360_, new_n10361_, new_n10362_, new_n10363_,
    new_n10364_, new_n10365_, new_n10366_, new_n10367_, new_n10368_,
    new_n10369_, new_n10370_, new_n10371_, new_n10372_, new_n10373_,
    new_n10374_, new_n10375_, new_n10376_, new_n10377_, new_n10378_,
    new_n10379_, new_n10380_, new_n10381_, new_n10382_, new_n10383_,
    new_n10384_, new_n10385_, new_n10386_, new_n10387_, new_n10388_,
    new_n10389_, new_n10390_, new_n10391_, new_n10392_, new_n10393_,
    new_n10394_, new_n10395_, new_n10396_, new_n10397_, new_n10398_,
    new_n10399_, new_n10400_, new_n10401_, new_n10402_, new_n10403_,
    new_n10404_, new_n10405_, new_n10406_, new_n10407_, new_n10408_,
    new_n10409_, new_n10410_, new_n10411_, new_n10412_, new_n10413_,
    new_n10414_, new_n10415_, new_n10416_, new_n10417_, new_n10418_,
    new_n10419_, new_n10420_, new_n10421_, new_n10422_, new_n10423_,
    new_n10424_, new_n10425_, new_n10426_, new_n10427_, new_n10428_,
    new_n10429_, new_n10430_, new_n10431_, new_n10432_, new_n10433_,
    new_n10434_, new_n10435_, new_n10436_, new_n10437_, new_n10438_,
    new_n10439_, new_n10440_, new_n10441_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10448_,
    new_n10449_, new_n10450_, new_n10451_, new_n10452_, new_n10453_,
    new_n10454_, new_n10455_, new_n10456_, new_n10457_, new_n10458_,
    new_n10459_, new_n10460_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10890_, new_n10891_,
    new_n10892_, new_n10893_, new_n10894_, new_n10895_, new_n10896_,
    new_n10897_, new_n10898_, new_n10899_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11221_,
    new_n11222_, new_n11223_, new_n11224_, new_n11225_, new_n11226_,
    new_n11227_, new_n11228_, new_n11229_, new_n11230_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11452_, new_n11453_,
    new_n11454_, new_n11455_, new_n11456_, new_n11457_, new_n11458_,
    new_n11459_, new_n11460_, new_n11461_, new_n11462_, new_n11463_,
    new_n11464_, new_n11465_, new_n11466_, new_n11467_, new_n11468_,
    new_n11469_, new_n11470_, new_n11471_, new_n11472_, new_n11473_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11761_, new_n11762_, new_n11763_,
    new_n11764_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11771_, new_n11772_, new_n11773_,
    new_n11774_, new_n11775_, new_n11776_, new_n11777_, new_n11778_,
    new_n11779_, new_n11780_, new_n11781_, new_n11782_, new_n11783_,
    new_n11784_, new_n11785_, new_n11786_, new_n11787_, new_n11788_,
    new_n11789_, new_n11790_, new_n11791_, new_n11792_, new_n11793_,
    new_n11794_, new_n11795_, new_n11796_, new_n11797_, new_n11798_,
    new_n11799_, new_n11800_, new_n11801_, new_n11802_, new_n11803_,
    new_n11804_, new_n11805_, new_n11806_, new_n11807_, new_n11808_,
    new_n11809_, new_n11810_, new_n11811_, new_n11812_, new_n11813_,
    new_n11814_, new_n11815_, new_n11816_, new_n11817_, new_n11818_,
    new_n11819_, new_n11820_, new_n11821_, new_n11822_, new_n11823_,
    new_n11824_, new_n11825_, new_n11826_, new_n11827_, new_n11828_,
    new_n11829_, new_n11830_, new_n11831_, new_n11832_, new_n11833_,
    new_n11834_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11855_, new_n11856_, new_n11857_, new_n11858_,
    new_n11859_, new_n11860_, new_n11861_, new_n11862_, new_n11863_,
    new_n11864_, new_n11865_, new_n11866_, new_n11867_, new_n11868_,
    new_n11869_, new_n11870_, new_n11871_, new_n11872_, new_n11873_,
    new_n11874_, new_n11875_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11906_, new_n11907_, new_n11908_,
    new_n11909_, new_n11910_, new_n11911_, new_n11912_, new_n11913_,
    new_n11914_, new_n11915_, new_n11916_, new_n11917_, new_n11918_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12130_, new_n12131_, new_n12132_, new_n12133_,
    new_n12134_, new_n12135_, new_n12136_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12278_, new_n12279_,
    new_n12280_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12286_, new_n12287_, new_n12288_, new_n12289_,
    new_n12290_, new_n12291_, new_n12292_, new_n12293_, new_n12294_,
    new_n12295_, new_n12296_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12961_,
    new_n12962_, new_n12963_, new_n12964_, new_n12965_, new_n12966_,
    new_n12967_, new_n12968_, new_n12969_, new_n12970_, new_n12971_,
    new_n12972_, new_n12973_, new_n12974_, new_n12975_, new_n12976_,
    new_n12977_, new_n12978_, new_n12979_, new_n12980_, new_n12981_,
    new_n12982_, new_n12983_, new_n12984_, new_n12985_, new_n12986_,
    new_n12987_, new_n12988_, new_n12989_, new_n12990_, new_n12991_,
    new_n12992_, new_n12993_, new_n12994_, new_n12995_, new_n12996_,
    new_n12997_, new_n12998_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13010_, new_n13011_, new_n13012_, new_n13013_,
    new_n13014_, new_n13015_, new_n13016_, new_n13017_, new_n13018_,
    new_n13019_, new_n13020_, new_n13021_, new_n13022_, new_n13023_,
    new_n13024_, new_n13025_, new_n13026_, new_n13027_, new_n13028_,
    new_n13029_, new_n13030_, new_n13031_, new_n13032_, new_n13033_,
    new_n13034_, new_n13035_, new_n13036_, new_n13037_, new_n13038_,
    new_n13039_, new_n13040_, new_n13041_, new_n13042_, new_n13043_,
    new_n13044_, new_n13045_, new_n13046_, new_n13047_, new_n13048_,
    new_n13049_, new_n13050_, new_n13051_, new_n13052_, new_n13053_,
    new_n13054_, new_n13055_, new_n13056_, new_n13057_, new_n13058_,
    new_n13059_, new_n13060_, new_n13061_, new_n13062_, new_n13063_,
    new_n13064_, new_n13065_, new_n13066_, new_n13067_, new_n13068_,
    new_n13069_, new_n13070_, new_n13071_, new_n13072_, new_n13073_,
    new_n13074_, new_n13075_, new_n13076_, new_n13077_, new_n13078_,
    new_n13079_, new_n13080_, new_n13081_, new_n13082_, new_n13083_,
    new_n13084_, new_n13085_, new_n13086_, new_n13087_, new_n13088_,
    new_n13089_, new_n13090_, new_n13091_, new_n13092_, new_n13093_,
    new_n13094_, new_n13095_, new_n13096_, new_n13097_, new_n13098_,
    new_n13099_, new_n13100_, new_n13101_, new_n13102_, new_n13103_,
    new_n13104_, new_n13105_, new_n13106_, new_n13107_, new_n13108_,
    new_n13109_, new_n13110_, new_n13111_, new_n13112_, new_n13113_,
    new_n13114_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13120_, new_n13121_, new_n13122_, new_n13123_,
    new_n13124_, new_n13125_, new_n13126_, new_n13127_, new_n13128_,
    new_n13129_, new_n13130_, new_n13131_, new_n13132_, new_n13133_,
    new_n13134_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13139_, new_n13140_, new_n13141_, new_n13142_, new_n13143_,
    new_n13144_, new_n13145_, new_n13146_, new_n13147_, new_n13148_,
    new_n13149_, new_n13150_, new_n13151_, new_n13152_, new_n13153_,
    new_n13154_, new_n13155_, new_n13156_, new_n13157_, new_n13158_,
    new_n13159_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13167_, new_n13168_,
    new_n13169_, new_n13170_, new_n13171_, new_n13172_, new_n13173_,
    new_n13174_, new_n13175_, new_n13176_, new_n13177_, new_n13178_,
    new_n13179_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13185_, new_n13186_, new_n13187_, new_n13188_,
    new_n13189_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13195_, new_n13196_, new_n13197_, new_n13198_,
    new_n13199_, new_n13200_, new_n13201_, new_n13202_, new_n13203_,
    new_n13204_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13218_,
    new_n13219_, new_n13220_, new_n13221_, new_n13222_, new_n13223_,
    new_n13224_, new_n13225_, new_n13226_, new_n13227_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13233_,
    new_n13234_, new_n13235_, new_n13236_, new_n13237_, new_n13238_,
    new_n13239_, new_n13240_, new_n13241_, new_n13242_, new_n13243_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13250_, new_n13251_, new_n13252_, new_n13253_,
    new_n13254_, new_n13255_, new_n13256_, new_n13257_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13263_,
    new_n13264_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13269_, new_n13270_, new_n13271_, new_n13272_, new_n13273_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_,
    new_n13359_, new_n13360_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13367_, new_n13368_,
    new_n13369_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13376_, new_n13377_, new_n13378_,
    new_n13379_, new_n13380_, new_n13381_, new_n13382_, new_n13383_,
    new_n13384_, new_n13385_, new_n13386_, new_n13387_, new_n13388_,
    new_n13389_, new_n13390_, new_n13391_, new_n13392_, new_n13393_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13562_, new_n13563_, new_n13564_,
    new_n13565_, new_n13566_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13695_, new_n13696_, new_n13697_, new_n13698_, new_n13699_,
    new_n13700_, new_n13701_, new_n13702_, new_n13703_, new_n13704_,
    new_n13705_, new_n13706_, new_n13707_, new_n13708_, new_n13709_,
    new_n13710_, new_n13711_, new_n13712_, new_n13713_, new_n13714_,
    new_n13715_, new_n13716_, new_n13717_, new_n13718_, new_n13719_,
    new_n13720_, new_n13721_, new_n13722_, new_n13723_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13730_, new_n13731_, new_n13732_, new_n13733_, new_n13734_,
    new_n13735_, new_n13736_, new_n13737_, new_n13738_, new_n13739_,
    new_n13740_, new_n13741_, new_n13742_, new_n13743_, new_n13744_,
    new_n13745_, new_n13746_, new_n13747_, new_n13748_, new_n13749_,
    new_n13750_, new_n13751_, new_n13752_, new_n13753_, new_n13754_,
    new_n13755_, new_n13756_, new_n13757_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13766_, new_n13767_, new_n13768_, new_n13769_,
    new_n13770_, new_n13771_, new_n13772_, new_n13773_, new_n13774_,
    new_n13775_, new_n13776_, new_n13777_, new_n13778_, new_n13779_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14238_,
    new_n14239_, new_n14240_, new_n14241_, new_n14242_, new_n14243_,
    new_n14244_, new_n14245_, new_n14246_, new_n14247_, new_n14248_,
    new_n14249_, new_n14250_, new_n14251_, new_n14252_, new_n14253_,
    new_n14254_, new_n14255_, new_n14256_, new_n14257_, new_n14258_,
    new_n14259_, new_n14260_, new_n14261_, new_n14262_, new_n14263_,
    new_n14264_, new_n14265_, new_n14266_, new_n14267_, new_n14268_,
    new_n14269_, new_n14270_, new_n14271_, new_n14272_, new_n14273_,
    new_n14274_, new_n14275_, new_n14276_, new_n14277_, new_n14278_,
    new_n14279_, new_n14280_, new_n14281_, new_n14282_, new_n14283_,
    new_n14284_, new_n14285_, new_n14286_, new_n14287_, new_n14288_,
    new_n14289_, new_n14290_, new_n14291_, new_n14292_, new_n14293_,
    new_n14294_, new_n14295_, new_n14296_, new_n14297_, new_n14298_,
    new_n14299_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14351_, new_n14352_, new_n14353_,
    new_n14354_, new_n14355_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14362_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14370_, new_n14371_, new_n14372_, new_n14373_,
    new_n14374_, new_n14375_, new_n14376_, new_n14377_, new_n14378_,
    new_n14379_, new_n14380_, new_n14381_, new_n14382_, new_n14383_,
    new_n14384_, new_n14385_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14398_,
    new_n14399_, new_n14400_, new_n14401_, new_n14402_, new_n14403_,
    new_n14404_, new_n14405_, new_n14406_, new_n14407_, new_n14408_,
    new_n14409_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14416_, new_n14417_, new_n14418_,
    new_n14419_, new_n14420_, new_n14421_, new_n14422_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14435_, new_n14436_, new_n14437_, new_n14438_,
    new_n14439_, new_n14440_, new_n14441_, new_n14442_, new_n14443_,
    new_n14444_, new_n14445_, new_n14446_, new_n14447_, new_n14448_,
    new_n14449_, new_n14450_, new_n14451_, new_n14452_, new_n14453_,
    new_n14454_, new_n14455_, new_n14456_, new_n14457_, new_n14458_,
    new_n14459_, new_n14460_, new_n14461_, new_n14462_, new_n14463_,
    new_n14464_, new_n14465_, new_n14466_, new_n14467_, new_n14468_,
    new_n14469_, new_n14470_, new_n14471_, new_n14472_, new_n14473_,
    new_n14474_, new_n14475_, new_n14476_, new_n14477_, new_n14478_,
    new_n14479_, new_n14480_, new_n14481_, new_n14482_, new_n14483_,
    new_n14484_, new_n14485_, new_n14486_, new_n14487_, new_n14488_,
    new_n14489_, new_n14490_, new_n14491_, new_n14492_, new_n14493_,
    new_n14494_, new_n14495_, new_n14496_, new_n14497_, new_n14498_,
    new_n14499_, new_n14500_, new_n14501_, new_n14502_, new_n14503_,
    new_n14504_, new_n14505_, new_n14506_, new_n14507_, new_n14508_,
    new_n14509_, new_n14510_, new_n14511_, new_n14512_, new_n14513_,
    new_n14514_, new_n14515_, new_n14516_, new_n14517_, new_n14518_,
    new_n14519_, new_n14520_, new_n14521_, new_n14522_, new_n14523_,
    new_n14524_, new_n14525_, new_n14526_, new_n14527_, new_n14528_,
    new_n14529_, new_n14530_, new_n14531_, new_n14532_, new_n14533_,
    new_n14534_, new_n14535_, new_n14536_, new_n14537_, new_n14538_,
    new_n14539_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14608_,
    new_n14609_, new_n14610_, new_n14611_, new_n14612_, new_n14613_,
    new_n14614_, new_n14615_, new_n14616_, new_n14617_, new_n14618_,
    new_n14619_, new_n14620_, new_n14621_, new_n14622_, new_n14623_,
    new_n14624_, new_n14625_, new_n14626_, new_n14627_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14633_,
    new_n14634_, new_n14636_, new_n14637_, new_n14638_, new_n14639_,
    new_n14640_, new_n14641_, new_n14642_, new_n14643_, new_n14644_,
    new_n14645_, new_n14646_, new_n14647_, new_n14648_, new_n14649_,
    new_n14650_, new_n14651_, new_n14652_, new_n14653_, new_n14654_,
    new_n14655_, new_n14656_, new_n14657_, new_n14658_, new_n14659_,
    new_n14660_, new_n14661_, new_n14662_, new_n14663_, new_n14664_,
    new_n14665_, new_n14666_, new_n14667_, new_n14668_, new_n14669_,
    new_n14670_, new_n14671_, new_n14672_, new_n14673_, new_n14674_,
    new_n14675_, new_n14676_, new_n14677_, new_n14678_, new_n14679_,
    new_n14680_, new_n14681_, new_n14682_, new_n14683_, new_n14684_,
    new_n14685_, new_n14686_, new_n14687_, new_n14688_, new_n14689_,
    new_n14690_, new_n14691_, new_n14692_, new_n14693_, new_n14694_,
    new_n14695_, new_n14696_, new_n14697_, new_n14698_, new_n14699_,
    new_n14700_, new_n14701_, new_n14702_, new_n14703_, new_n14704_,
    new_n14705_, new_n14706_, new_n14707_, new_n14708_, new_n14709_,
    new_n14710_, new_n14711_, new_n14712_, new_n14713_, new_n14714_,
    new_n14715_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14733_, new_n14734_,
    new_n14735_, new_n14736_, new_n14737_, new_n14738_, new_n14739_,
    new_n14740_, new_n14741_, new_n14742_, new_n14743_, new_n14744_,
    new_n14745_, new_n14746_, new_n14747_, new_n14748_, new_n14749_,
    new_n14750_, new_n14751_, new_n14752_, new_n14753_, new_n14754_,
    new_n14755_, new_n14756_, new_n14757_, new_n14758_, new_n14759_,
    new_n14760_, new_n14761_, new_n14762_, new_n14763_, new_n14764_,
    new_n14765_, new_n14766_, new_n14767_, new_n14768_, new_n14769_,
    new_n14770_, new_n14771_, new_n14772_, new_n14773_, new_n14774_,
    new_n14775_, new_n14776_, new_n14777_, new_n14778_, new_n14779_,
    new_n14780_, new_n14781_, new_n14782_, new_n14783_, new_n14784_,
    new_n14785_, new_n14786_, new_n14787_, new_n14788_, new_n14789_,
    new_n14790_, new_n14791_, new_n14792_, new_n14793_, new_n14794_,
    new_n14795_, new_n14796_, new_n14797_, new_n14798_, new_n14799_,
    new_n14800_, new_n14801_, new_n14802_, new_n14803_, new_n14804_,
    new_n14805_, new_n14806_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14823_, new_n14824_,
    new_n14825_, new_n14826_, new_n14827_, new_n14828_, new_n14829_,
    new_n14830_, new_n14831_, new_n14832_, new_n14833_, new_n14834_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14908_, new_n14909_,
    new_n14910_, new_n14911_, new_n14912_, new_n14913_, new_n14914_,
    new_n14915_, new_n14916_, new_n14917_, new_n14918_, new_n14919_,
    new_n14920_, new_n14921_, new_n14922_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14930_, new_n14931_, new_n14932_, new_n14933_, new_n14934_,
    new_n14935_, new_n14936_, new_n14937_, new_n14938_, new_n14939_,
    new_n14940_, new_n14941_, new_n14942_, new_n14943_, new_n14944_,
    new_n14945_, new_n14946_, new_n14947_, new_n14948_, new_n14949_,
    new_n14950_, new_n14951_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14964_,
    new_n14965_, new_n14966_, new_n14967_, new_n14968_, new_n14969_,
    new_n14970_, new_n14971_, new_n14972_, new_n14973_, new_n14974_,
    new_n14975_, new_n14976_, new_n14977_, new_n14978_, new_n14979_,
    new_n14980_, new_n14981_, new_n14982_, new_n14983_, new_n14984_,
    new_n14985_, new_n14986_, new_n14987_, new_n14988_, new_n14989_,
    new_n14990_, new_n14991_, new_n14992_, new_n14993_, new_n14994_,
    new_n14995_, new_n14996_, new_n14997_, new_n14998_, new_n14999_,
    new_n15000_, new_n15001_, new_n15002_, new_n15003_, new_n15004_,
    new_n15005_, new_n15006_, new_n15007_, new_n15008_, new_n15009_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15307_, new_n15308_, new_n15309_, new_n15310_, new_n15311_,
    new_n15312_, new_n15313_, new_n15314_, new_n15315_, new_n15316_,
    new_n15317_, new_n15318_, new_n15319_, new_n15320_, new_n15321_,
    new_n15322_, new_n15323_, new_n15324_, new_n15325_, new_n15326_,
    new_n15327_, new_n15328_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15367_,
    new_n15368_, new_n15369_, new_n15370_, new_n15371_, new_n15372_,
    new_n15373_, new_n15374_, new_n15375_, new_n15376_, new_n15377_,
    new_n15378_, new_n15379_, new_n15380_, new_n15381_, new_n15382_,
    new_n15383_, new_n15384_, new_n15385_, new_n15386_, new_n15387_,
    new_n15388_, new_n15389_, new_n15390_, new_n15391_, new_n15392_,
    new_n15393_, new_n15394_, new_n15395_, new_n15396_, new_n15397_,
    new_n15398_, new_n15399_, new_n15400_, new_n15401_, new_n15402_,
    new_n15403_, new_n15404_, new_n15405_, new_n15406_, new_n15407_,
    new_n15408_, new_n15409_, new_n15410_, new_n15411_, new_n15412_,
    new_n15413_, new_n15414_, new_n15415_, new_n15416_, new_n15417_,
    new_n15418_, new_n15419_, new_n15420_, new_n15421_, new_n15422_,
    new_n15423_, new_n15424_, new_n15426_, new_n15427_, new_n15428_,
    new_n15429_, new_n15430_, new_n15431_, new_n15432_, new_n15433_,
    new_n15434_, new_n15435_, new_n15436_, new_n15437_, new_n15438_,
    new_n15439_, new_n15440_, new_n15441_, new_n15442_, new_n15443_,
    new_n15444_, new_n15445_, new_n15446_, new_n15447_, new_n15448_,
    new_n15449_, new_n15450_, new_n15451_, new_n15452_, new_n15453_,
    new_n15454_, new_n15455_, new_n15456_, new_n15457_, new_n15458_,
    new_n15459_, new_n15460_, new_n15461_, new_n15462_, new_n15463_,
    new_n15464_, new_n15465_, new_n15466_, new_n15467_, new_n15468_,
    new_n15469_, new_n15470_, new_n15471_, new_n15472_, new_n15473_,
    new_n15474_, new_n15475_, new_n15476_, new_n15477_, new_n15478_,
    new_n15479_, new_n15480_, new_n15481_, new_n15482_, new_n15483_,
    new_n15484_, new_n15485_, new_n15486_, new_n15487_, new_n15488_,
    new_n15489_, new_n15490_, new_n15491_, new_n15492_, new_n15493_,
    new_n15494_, new_n15495_, new_n15496_, new_n15497_, new_n15498_,
    new_n15499_, new_n15500_, new_n15501_, new_n15502_, new_n15503_,
    new_n15504_, new_n15505_, new_n15506_, new_n15507_, new_n15508_,
    new_n15509_, new_n15510_, new_n15511_, new_n15512_, new_n15513_,
    new_n15514_, new_n15515_, new_n15516_, new_n15517_, new_n15518_,
    new_n15519_, new_n15520_, new_n15521_, new_n15522_, new_n15523_,
    new_n15524_, new_n15525_, new_n15526_, new_n15527_, new_n15528_,
    new_n15529_, new_n15530_, new_n15531_, new_n15532_, new_n15533_,
    new_n15534_, new_n15535_, new_n15536_, new_n15537_, new_n15538_,
    new_n15539_, new_n15540_, new_n15541_, new_n15542_, new_n15543_,
    new_n15544_, new_n15545_, new_n15546_, new_n15547_, new_n15548_,
    new_n15549_, new_n15550_, new_n15551_, new_n15552_, new_n15553_,
    new_n15554_, new_n15555_, new_n15556_, new_n15557_, new_n15558_,
    new_n15559_, new_n15560_, new_n15561_, new_n15562_, new_n15563_,
    new_n15564_, new_n15565_, new_n15566_, new_n15567_, new_n15568_,
    new_n15569_, new_n15570_, new_n15571_, new_n15572_, new_n15573_,
    new_n15574_, new_n15575_, new_n15576_, new_n15577_, new_n15578_,
    new_n15579_, new_n15580_, new_n15581_, new_n15582_, new_n15583_,
    new_n15584_, new_n15585_, new_n15586_, new_n15587_, new_n15588_,
    new_n15589_, new_n15590_, new_n15591_, new_n15592_, new_n15593_,
    new_n15594_, new_n15595_, new_n15596_, new_n15597_, new_n15598_,
    new_n15599_, new_n15600_, new_n15601_, new_n15602_, new_n15603_,
    new_n15604_, new_n15605_, new_n15606_, new_n15607_, new_n15608_,
    new_n15609_, new_n15610_, new_n15611_, new_n15612_, new_n15613_,
    new_n15614_, new_n15615_, new_n15616_, new_n15617_, new_n15618_,
    new_n15619_, new_n15620_, new_n15621_, new_n15622_, new_n15623_,
    new_n15624_, new_n15625_, new_n15626_, new_n15627_, new_n15628_,
    new_n15629_, new_n15630_, new_n15631_, new_n15632_, new_n15633_,
    new_n15634_, new_n15635_, new_n15636_, new_n15637_, new_n15638_,
    new_n15639_, new_n15640_, new_n15641_, new_n15642_, new_n15643_,
    new_n15644_, new_n15645_, new_n15646_, new_n15647_, new_n15648_,
    new_n15649_, new_n15650_, new_n15651_, new_n15652_, new_n15653_,
    new_n15654_, new_n15655_, new_n15656_, new_n15657_, new_n15658_,
    new_n15659_, new_n15660_, new_n15661_, new_n15662_, new_n15663_,
    new_n15664_, new_n15665_, new_n15666_, new_n15667_, new_n15668_,
    new_n15669_, new_n15670_, new_n15671_, new_n15672_, new_n15673_,
    new_n15674_, new_n15675_, new_n15676_, new_n15677_, new_n15678_,
    new_n15679_, new_n15680_, new_n15681_, new_n15682_, new_n15683_,
    new_n15684_, new_n15685_, new_n15686_, new_n15687_, new_n15688_,
    new_n15689_, new_n15690_, new_n15691_, new_n15692_, new_n15693_,
    new_n15694_, new_n15695_, new_n15696_, new_n15697_, new_n15698_,
    new_n15699_, new_n15700_, new_n15701_, new_n15702_, new_n15703_,
    new_n15704_, new_n15705_, new_n15706_, new_n15707_, new_n15708_,
    new_n15709_, new_n15710_, new_n15711_, new_n15712_, new_n15713_,
    new_n15714_, new_n15715_, new_n15716_, new_n15717_, new_n15718_,
    new_n15719_, new_n15720_, new_n15721_, new_n15722_, new_n15723_,
    new_n15724_, new_n15725_, new_n15726_, new_n15727_, new_n15728_,
    new_n15729_, new_n15730_, new_n15731_, new_n15732_, new_n15733_,
    new_n15734_, new_n15735_, new_n15736_, new_n15737_, new_n15738_,
    new_n15739_, new_n15740_, new_n15741_, new_n15742_, new_n15743_,
    new_n15744_, new_n15745_, new_n15746_, new_n15747_, new_n15748_,
    new_n15749_, new_n15750_, new_n15751_, new_n15752_, new_n15753_,
    new_n15754_, new_n15755_, new_n15756_, new_n15757_, new_n15758_,
    new_n15759_, new_n15760_, new_n15761_, new_n15762_, new_n15763_,
    new_n15764_, new_n15765_, new_n15766_, new_n15767_, new_n15768_,
    new_n15769_, new_n15770_, new_n15771_, new_n15772_, new_n15773_,
    new_n15774_, new_n15775_, new_n15776_, new_n15777_, new_n15778_,
    new_n15779_, new_n15780_, new_n15781_, new_n15782_, new_n15783_,
    new_n15784_, new_n15785_, new_n15786_, new_n15787_, new_n15788_,
    new_n15789_, new_n15790_, new_n15791_, new_n15792_, new_n15793_,
    new_n15794_, new_n15795_, new_n15796_, new_n15797_, new_n15798_,
    new_n15799_, new_n15800_, new_n15801_, new_n15802_, new_n15803_,
    new_n15804_, new_n15805_, new_n15806_, new_n15807_, new_n15808_,
    new_n15809_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16074_,
    new_n16075_, new_n16076_, new_n16077_, new_n16078_, new_n16079_,
    new_n16080_, new_n16081_, new_n16082_, new_n16083_, new_n16084_,
    new_n16085_, new_n16086_, new_n16087_, new_n16088_, new_n16089_,
    new_n16090_, new_n16091_, new_n16092_, new_n16093_, new_n16094_,
    new_n16095_, new_n16096_, new_n16097_, new_n16098_, new_n16099_,
    new_n16100_, new_n16101_, new_n16102_, new_n16103_, new_n16104_,
    new_n16105_, new_n16106_, new_n16107_, new_n16108_, new_n16109_,
    new_n16110_, new_n16111_, new_n16112_, new_n16113_, new_n16114_,
    new_n16115_, new_n16116_, new_n16117_, new_n16118_, new_n16119_,
    new_n16120_, new_n16121_, new_n16122_, new_n16123_, new_n16124_,
    new_n16125_, new_n16126_, new_n16127_, new_n16128_, new_n16129_,
    new_n16130_, new_n16131_, new_n16132_, new_n16133_, new_n16134_,
    new_n16135_, new_n16136_, new_n16137_, new_n16138_, new_n16139_,
    new_n16140_, new_n16141_, new_n16142_, new_n16143_, new_n16144_,
    new_n16145_, new_n16146_, new_n16147_, new_n16148_, new_n16149_,
    new_n16150_, new_n16151_, new_n16152_, new_n16153_, new_n16154_,
    new_n16155_, new_n16156_, new_n16157_, new_n16158_, new_n16159_,
    new_n16160_, new_n16161_, new_n16162_, new_n16163_, new_n16164_,
    new_n16165_, new_n16166_, new_n16167_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16830_, new_n16831_, new_n16832_,
    new_n16833_, new_n16834_, new_n16835_, new_n16836_, new_n16837_,
    new_n16838_, new_n16839_, new_n16840_, new_n16841_, new_n16842_,
    new_n16843_, new_n16844_, new_n16845_, new_n16846_, new_n16847_,
    new_n16848_, new_n16849_, new_n16850_, new_n16851_, new_n16852_,
    new_n16853_, new_n16854_, new_n16855_, new_n16856_, new_n16857_,
    new_n16858_, new_n16859_, new_n16860_, new_n16861_, new_n16862_,
    new_n16863_, new_n16864_, new_n16865_, new_n16866_, new_n16867_,
    new_n16868_, new_n16869_, new_n16870_, new_n16871_, new_n16872_,
    new_n16873_, new_n16874_, new_n16875_, new_n16876_, new_n16877_,
    new_n16878_, new_n16879_, new_n16880_, new_n16881_, new_n16882_,
    new_n16883_, new_n16884_, new_n16885_, new_n16886_, new_n16887_,
    new_n16888_, new_n16889_, new_n16890_, new_n16891_, new_n16892_,
    new_n16893_, new_n16894_, new_n16895_, new_n16896_, new_n16897_,
    new_n16898_, new_n16899_, new_n16900_, new_n16901_, new_n16902_,
    new_n16903_, new_n16904_, new_n16905_, new_n16906_, new_n16907_,
    new_n16908_, new_n16909_, new_n16910_, new_n16911_, new_n16912_,
    new_n16913_, new_n16914_, new_n16915_, new_n16916_, new_n16917_,
    new_n16918_, new_n16919_, new_n16920_, new_n16921_, new_n16922_,
    new_n16923_, new_n16924_, new_n16925_, new_n16926_, new_n16927_,
    new_n16928_, new_n16929_, new_n16930_, new_n16931_, new_n16932_,
    new_n16933_, new_n16934_, new_n16935_, new_n16936_, new_n16937_,
    new_n16938_, new_n16939_, new_n16940_, new_n16941_, new_n16942_,
    new_n16943_, new_n16944_, new_n16945_, new_n16946_, new_n16947_,
    new_n16948_, new_n16949_, new_n16950_, new_n16951_, new_n16952_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16966_, new_n16967_,
    new_n16968_, new_n16969_, new_n16970_, new_n16971_, new_n16972_,
    new_n16973_, new_n16974_, new_n16975_, new_n16976_, new_n16977_,
    new_n16978_, new_n16979_, new_n16980_, new_n16981_, new_n16982_,
    new_n16983_, new_n16984_, new_n16985_, new_n16986_, new_n16987_,
    new_n16988_, new_n16989_, new_n16990_, new_n16991_, new_n16992_,
    new_n16993_, new_n16994_, new_n16995_, new_n16996_, new_n16997_,
    new_n16998_, new_n16999_, new_n17000_, new_n17001_, new_n17002_,
    new_n17003_, new_n17004_, new_n17005_, new_n17006_, new_n17007_,
    new_n17008_, new_n17009_, new_n17010_, new_n17011_, new_n17012_,
    new_n17013_, new_n17014_, new_n17015_, new_n17016_, new_n17017_,
    new_n17018_, new_n17019_, new_n17020_, new_n17021_, new_n17022_,
    new_n17023_, new_n17024_, new_n17025_, new_n17026_, new_n17027_,
    new_n17028_, new_n17029_, new_n17030_, new_n17031_, new_n17032_,
    new_n17033_, new_n17034_, new_n17035_, new_n17036_, new_n17037_,
    new_n17038_, new_n17039_, new_n17040_, new_n17041_, new_n17042_,
    new_n17043_, new_n17044_, new_n17045_, new_n17046_, new_n17047_,
    new_n17048_, new_n17049_, new_n17050_, new_n17051_, new_n17052_,
    new_n17053_, new_n17054_, new_n17055_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17070_, new_n17071_, new_n17072_,
    new_n17073_, new_n17074_, new_n17075_, new_n17076_, new_n17077_,
    new_n17078_, new_n17079_, new_n17080_, new_n17081_, new_n17082_,
    new_n17083_, new_n17084_, new_n17085_, new_n17086_, new_n17087_,
    new_n17088_, new_n17089_, new_n17090_, new_n17091_, new_n17092_,
    new_n17093_, new_n17094_, new_n17095_, new_n17096_, new_n17097_,
    new_n17098_, new_n17099_, new_n17100_, new_n17101_, new_n17102_,
    new_n17103_, new_n17104_, new_n17105_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17120_, new_n17121_, new_n17122_, new_n17123_,
    new_n17124_, new_n17125_, new_n17126_, new_n17127_, new_n17128_,
    new_n17129_, new_n17130_, new_n17131_, new_n17132_, new_n17133_,
    new_n17134_, new_n17135_, new_n17136_, new_n17137_, new_n17138_,
    new_n17139_, new_n17140_, new_n17141_, new_n17142_, new_n17143_,
    new_n17144_, new_n17145_, new_n17146_, new_n17147_, new_n17148_,
    new_n17149_, new_n17150_, new_n17151_, new_n17152_, new_n17153_,
    new_n17154_, new_n17155_, new_n17156_, new_n17157_, new_n17158_,
    new_n17159_, new_n17160_, new_n17161_, new_n17162_, new_n17163_,
    new_n17164_, new_n17165_, new_n17166_, new_n17167_, new_n17168_,
    new_n17169_, new_n17170_, new_n17171_, new_n17172_, new_n17173_,
    new_n17174_, new_n17175_, new_n17176_, new_n17177_, new_n17178_,
    new_n17179_, new_n17180_, new_n17181_, new_n17182_, new_n17183_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17229_, new_n17230_, new_n17231_, new_n17232_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17311_, new_n17312_, new_n17313_,
    new_n17314_, new_n17315_, new_n17316_, new_n17317_, new_n17318_,
    new_n17319_, new_n17320_, new_n17321_, new_n17322_, new_n17323_,
    new_n17324_, new_n17325_, new_n17326_, new_n17327_, new_n17328_,
    new_n17329_, new_n17330_, new_n17331_, new_n17332_, new_n17333_,
    new_n17334_, new_n17335_, new_n17336_, new_n17337_, new_n17338_,
    new_n17339_, new_n17340_, new_n17341_, new_n17342_, new_n17343_,
    new_n17344_, new_n17345_, new_n17346_, new_n17347_, new_n17348_,
    new_n17349_, new_n17350_, new_n17351_, new_n17352_, new_n17353_,
    new_n17354_, new_n17355_, new_n17356_, new_n17357_, new_n17358_,
    new_n17359_, new_n17360_, new_n17361_, new_n17362_, new_n17363_,
    new_n17364_, new_n17365_, new_n17366_, new_n17367_, new_n17368_,
    new_n17369_, new_n17370_, new_n17371_, new_n17372_, new_n17373_,
    new_n17374_, new_n17375_, new_n17376_, new_n17377_, new_n17378_,
    new_n17379_, new_n17380_, new_n17381_, new_n17382_, new_n17383_,
    new_n17384_, new_n17385_, new_n17386_, new_n17387_, new_n17388_,
    new_n17389_, new_n17390_, new_n17391_, new_n17392_, new_n17393_,
    new_n17394_, new_n17395_, new_n17396_, new_n17397_, new_n17398_,
    new_n17399_, new_n17400_, new_n17401_, new_n17402_, new_n17403_,
    new_n17404_, new_n17405_, new_n17406_, new_n17407_, new_n17408_,
    new_n17409_, new_n17410_, new_n17411_, new_n17412_, new_n17414_,
    new_n17415_, new_n17416_, new_n17417_, new_n17418_, new_n17419_,
    new_n17420_, new_n17421_, new_n17422_, new_n17423_, new_n17424_,
    new_n17425_, new_n17426_, new_n17427_, new_n17428_, new_n17429_,
    new_n17430_, new_n17431_, new_n17432_, new_n17433_, new_n17434_,
    new_n17435_, new_n17436_, new_n17437_, new_n17438_, new_n17439_,
    new_n17440_, new_n17441_, new_n17442_, new_n17443_, new_n17444_,
    new_n17445_, new_n17446_, new_n17447_, new_n17448_, new_n17449_,
    new_n17450_, new_n17451_, new_n17452_, new_n17453_, new_n17454_,
    new_n17455_, new_n17456_, new_n17457_, new_n17458_, new_n17459_,
    new_n17460_, new_n17461_, new_n17462_, new_n17463_, new_n17464_,
    new_n17465_, new_n17466_, new_n17467_, new_n17468_, new_n17469_,
    new_n17470_, new_n17471_, new_n17472_, new_n17473_, new_n17474_,
    new_n17475_, new_n17476_, new_n17477_, new_n17478_, new_n17479_,
    new_n17480_, new_n17481_, new_n17482_, new_n17483_, new_n17484_,
    new_n17485_, new_n17486_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17492_, new_n17493_, new_n17494_,
    new_n17495_, new_n17496_, new_n17497_, new_n17498_, new_n17499_,
    new_n17500_, new_n17501_, new_n17502_, new_n17503_, new_n17504_,
    new_n17505_, new_n17506_, new_n17507_, new_n17508_, new_n17509_,
    new_n17510_, new_n17511_, new_n17512_, new_n17513_, new_n17514_,
    new_n17515_, new_n17516_, new_n17517_, new_n17518_, new_n17519_,
    new_n17520_, new_n17521_, new_n17522_, new_n17523_, new_n17524_,
    new_n17525_, new_n17526_, new_n17527_, new_n17528_, new_n17529_,
    new_n17530_, new_n17531_, new_n17532_, new_n17533_, new_n17534_,
    new_n17535_, new_n17536_, new_n17537_, new_n17538_, new_n17539_,
    new_n17540_, new_n17541_, new_n17542_, new_n17543_, new_n17544_,
    new_n17545_, new_n17546_, new_n17547_, new_n17548_, new_n17549_,
    new_n17550_, new_n17551_, new_n17552_, new_n17553_, new_n17554_,
    new_n17555_, new_n17556_, new_n17557_, new_n17558_, new_n17559_,
    new_n17560_, new_n17561_, new_n17562_, new_n17563_, new_n17564_,
    new_n17565_, new_n17566_, new_n17567_, new_n17568_, new_n17569_,
    new_n17570_, new_n17571_, new_n17572_, new_n17573_, new_n17574_,
    new_n17575_, new_n17576_, new_n17577_, new_n17578_, new_n17579_,
    new_n17580_, new_n17581_, new_n17582_, new_n17583_, new_n17584_,
    new_n17585_, new_n17586_, new_n17587_, new_n17588_, new_n17589_,
    new_n17590_, new_n17591_, new_n17592_, new_n17593_, new_n17594_,
    new_n17595_, new_n17596_, new_n17597_, new_n17598_, new_n17599_,
    new_n17600_, new_n17601_, new_n17602_, new_n17603_, new_n17604_,
    new_n17605_, new_n17606_, new_n17607_, new_n17608_, new_n17609_,
    new_n17610_, new_n17611_, new_n17612_, new_n17613_, new_n17614_,
    new_n17615_, new_n17616_, new_n17617_, new_n17618_, new_n17619_,
    new_n17620_, new_n17621_, new_n17622_, new_n17623_, new_n17624_,
    new_n17625_, new_n17626_, new_n17627_, new_n17628_, new_n17629_,
    new_n17630_, new_n17631_, new_n17632_, new_n17633_, new_n17634_,
    new_n17635_, new_n17636_, new_n17637_, new_n17638_, new_n17639_,
    new_n17640_, new_n17641_, new_n17642_, new_n17643_, new_n17644_,
    new_n17645_, new_n17646_, new_n17647_, new_n17648_, new_n17649_,
    new_n17650_, new_n17651_, new_n17652_, new_n17653_, new_n17654_,
    new_n17655_, new_n17656_, new_n17657_, new_n17658_, new_n17659_,
    new_n17660_, new_n17661_, new_n17662_, new_n17663_, new_n17664_,
    new_n17665_, new_n17666_, new_n17667_, new_n17668_, new_n17669_,
    new_n17670_, new_n17671_, new_n17672_, new_n17673_, new_n17674_,
    new_n17675_, new_n17676_, new_n17677_, new_n17678_, new_n17679_,
    new_n17680_, new_n17681_, new_n17682_, new_n17683_, new_n17684_,
    new_n17685_, new_n17686_, new_n17687_, new_n17688_, new_n17689_,
    new_n17690_, new_n17691_, new_n17692_, new_n17693_, new_n17694_,
    new_n17695_, new_n17696_, new_n17697_, new_n17698_, new_n17699_,
    new_n17700_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17747_, new_n17748_, new_n17749_, new_n17750_,
    new_n17751_, new_n17752_, new_n17753_, new_n17754_, new_n17755_,
    new_n17756_, new_n17757_, new_n17758_, new_n17759_, new_n17760_,
    new_n17761_, new_n17762_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17791_, new_n17792_, new_n17793_, new_n17794_, new_n17795_,
    new_n17796_, new_n17797_, new_n17798_, new_n17799_, new_n17800_,
    new_n17801_, new_n17802_, new_n17803_, new_n17804_, new_n17805_,
    new_n17806_, new_n17807_, new_n17808_, new_n17809_, new_n17810_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17832_, new_n17833_, new_n17834_, new_n17835_,
    new_n17836_, new_n17837_, new_n17838_, new_n17839_, new_n17840_,
    new_n17841_, new_n17842_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17887_, new_n17888_, new_n17889_, new_n17890_,
    new_n17891_, new_n17892_, new_n17893_, new_n17894_, new_n17895_,
    new_n17896_, new_n17897_, new_n17898_, new_n17899_, new_n17900_,
    new_n17901_, new_n17902_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17974_, new_n17975_, new_n17976_,
    new_n17977_, new_n17978_, new_n17979_, new_n17980_, new_n17981_,
    new_n17982_, new_n17983_, new_n17984_, new_n17985_, new_n17986_,
    new_n17987_, new_n17988_, new_n17989_, new_n17990_, new_n17991_,
    new_n17992_, new_n17993_, new_n17994_, new_n17995_, new_n17996_,
    new_n17997_, new_n17998_, new_n17999_, new_n18000_, new_n18001_,
    new_n18002_, new_n18003_, new_n18004_, new_n18005_, new_n18006_,
    new_n18007_, new_n18008_, new_n18009_, new_n18010_, new_n18011_,
    new_n18012_, new_n18013_, new_n18014_, new_n18015_, new_n18016_,
    new_n18017_, new_n18018_, new_n18019_, new_n18020_, new_n18021_,
    new_n18022_, new_n18023_, new_n18024_, new_n18025_, new_n18026_,
    new_n18027_, new_n18028_, new_n18029_, new_n18030_, new_n18031_,
    new_n18032_, new_n18033_, new_n18034_, new_n18035_, new_n18036_,
    new_n18037_, new_n18038_, new_n18039_, new_n18040_, new_n18041_,
    new_n18042_, new_n18043_, new_n18044_, new_n18045_, new_n18046_,
    new_n18047_, new_n18048_, new_n18049_, new_n18050_, new_n18051_,
    new_n18052_, new_n18053_, new_n18054_, new_n18055_, new_n18056_,
    new_n18057_, new_n18058_, new_n18059_, new_n18060_, new_n18061_,
    new_n18062_, new_n18063_, new_n18064_, new_n18065_, new_n18066_,
    new_n18067_, new_n18068_, new_n18069_, new_n18070_, new_n18071_,
    new_n18072_, new_n18073_, new_n18074_, new_n18075_, new_n18076_,
    new_n18077_, new_n18078_, new_n18079_, new_n18080_, new_n18081_,
    new_n18082_, new_n18083_, new_n18084_, new_n18085_, new_n18086_,
    new_n18087_, new_n18088_, new_n18089_, new_n18090_, new_n18091_,
    new_n18092_, new_n18093_, new_n18094_, new_n18095_, new_n18096_,
    new_n18097_, new_n18098_, new_n18099_, new_n18100_, new_n18101_,
    new_n18102_, new_n18103_, new_n18104_, new_n18105_, new_n18106_,
    new_n18107_, new_n18108_, new_n18109_, new_n18110_, new_n18111_,
    new_n18112_, new_n18113_, new_n18114_, new_n18115_, new_n18116_,
    new_n18117_, new_n18118_, new_n18119_, new_n18120_, new_n18121_,
    new_n18122_, new_n18123_, new_n18124_, new_n18125_, new_n18126_,
    new_n18127_, new_n18128_, new_n18129_, new_n18130_, new_n18131_,
    new_n18132_, new_n18133_, new_n18134_, new_n18135_, new_n18136_,
    new_n18137_, new_n18138_, new_n18139_, new_n18140_, new_n18141_,
    new_n18142_, new_n18143_, new_n18144_, new_n18145_, new_n18146_,
    new_n18147_, new_n18148_, new_n18149_, new_n18150_, new_n18151_,
    new_n18152_, new_n18153_, new_n18154_, new_n18155_, new_n18156_,
    new_n18157_, new_n18158_, new_n18159_, new_n18160_, new_n18161_,
    new_n18162_, new_n18163_, new_n18164_, new_n18165_, new_n18166_,
    new_n18167_, new_n18168_, new_n18169_, new_n18170_, new_n18171_,
    new_n18172_, new_n18173_, new_n18174_, new_n18175_, new_n18176_,
    new_n18177_, new_n18178_, new_n18179_, new_n18180_, new_n18181_,
    new_n18182_, new_n18183_, new_n18184_, new_n18185_, new_n18186_,
    new_n18187_, new_n18188_, new_n18189_, new_n18190_, new_n18191_,
    new_n18192_, new_n18193_, new_n18194_, new_n18195_, new_n18196_,
    new_n18197_, new_n18198_, new_n18199_, new_n18200_, new_n18201_,
    new_n18202_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18210_, new_n18211_,
    new_n18212_, new_n18213_, new_n18214_, new_n18215_, new_n18216_,
    new_n18217_, new_n18219_, new_n18220_, new_n18221_, new_n18222_,
    new_n18223_, new_n18224_, new_n18225_, new_n18226_, new_n18227_,
    new_n18228_, new_n18229_, new_n18230_, new_n18231_, new_n18232_,
    new_n18233_, new_n18234_, new_n18235_, new_n18236_, new_n18237_,
    new_n18238_, new_n18239_, new_n18240_, new_n18241_, new_n18242_,
    new_n18243_, new_n18244_, new_n18245_, new_n18246_, new_n18247_,
    new_n18248_, new_n18249_, new_n18250_, new_n18251_, new_n18252_,
    new_n18253_, new_n18254_, new_n18255_, new_n18256_, new_n18257_,
    new_n18258_, new_n18259_, new_n18260_, new_n18261_, new_n18262_,
    new_n18263_, new_n18264_, new_n18265_, new_n18266_, new_n18267_,
    new_n18268_, new_n18269_, new_n18270_, new_n18271_, new_n18272_,
    new_n18273_, new_n18274_, new_n18275_, new_n18276_, new_n18277_,
    new_n18278_, new_n18279_, new_n18280_, new_n18281_, new_n18282_,
    new_n18283_, new_n18284_, new_n18285_, new_n18286_, new_n18287_,
    new_n18288_, new_n18289_, new_n18290_, new_n18291_, new_n18292_,
    new_n18293_, new_n18294_, new_n18295_, new_n18296_, new_n18297_,
    new_n18298_, new_n18299_, new_n18300_, new_n18301_, new_n18302_,
    new_n18303_, new_n18304_, new_n18305_, new_n18306_, new_n18307_,
    new_n18308_, new_n18309_, new_n18310_, new_n18311_, new_n18312_,
    new_n18313_, new_n18314_, new_n18315_, new_n18316_, new_n18317_,
    new_n18318_, new_n18319_, new_n18320_, new_n18321_, new_n18322_,
    new_n18323_, new_n18324_, new_n18325_, new_n18326_, new_n18327_,
    new_n18328_, new_n18329_, new_n18330_, new_n18331_, new_n18332_,
    new_n18333_, new_n18334_, new_n18335_, new_n18336_, new_n18337_,
    new_n18338_, new_n18339_, new_n18340_, new_n18341_, new_n18342_,
    new_n18343_, new_n18344_, new_n18345_, new_n18346_, new_n18347_,
    new_n18348_, new_n18349_, new_n18350_, new_n18351_, new_n18352_,
    new_n18353_, new_n18354_, new_n18355_, new_n18356_, new_n18357_,
    new_n18358_, new_n18359_, new_n18360_, new_n18361_, new_n18362_,
    new_n18363_, new_n18364_, new_n18365_, new_n18366_, new_n18367_,
    new_n18368_, new_n18369_, new_n18370_, new_n18371_, new_n18372_,
    new_n18373_, new_n18374_, new_n18375_, new_n18376_, new_n18377_,
    new_n18378_, new_n18379_, new_n18380_, new_n18381_, new_n18382_,
    new_n18383_, new_n18384_, new_n18385_, new_n18386_, new_n18387_,
    new_n18388_, new_n18389_, new_n18390_, new_n18391_, new_n18392_,
    new_n18393_, new_n18394_, new_n18395_, new_n18396_, new_n18397_,
    new_n18398_, new_n18399_, new_n18400_, new_n18401_, new_n18402_,
    new_n18403_, new_n18404_, new_n18405_, new_n18406_, new_n18407_,
    new_n18408_, new_n18409_, new_n18410_, new_n18411_, new_n18412_,
    new_n18413_, new_n18414_, new_n18415_, new_n18416_, new_n18417_,
    new_n18418_, new_n18419_, new_n18420_, new_n18421_, new_n18422_,
    new_n18423_, new_n18424_, new_n18425_, new_n18426_, new_n18427_,
    new_n18428_, new_n18429_, new_n18430_, new_n18431_, new_n18432_,
    new_n18433_, new_n18434_, new_n18435_, new_n18436_, new_n18437_,
    new_n18438_, new_n18439_, new_n18440_, new_n18441_, new_n18442_,
    new_n18443_, new_n18444_, new_n18445_, new_n18446_, new_n18447_,
    new_n18448_, new_n18449_, new_n18450_, new_n18451_, new_n18452_,
    new_n18453_, new_n18454_, new_n18455_, new_n18456_, new_n18457_,
    new_n18458_, new_n18459_, new_n18460_, new_n18461_, new_n18462_,
    new_n18463_, new_n18464_, new_n18465_, new_n18466_, new_n18467_,
    new_n18468_, new_n18469_, new_n18470_, new_n18471_, new_n18472_,
    new_n18473_, new_n18474_, new_n18475_, new_n18476_, new_n18477_,
    new_n18478_, new_n18479_, new_n18480_, new_n18481_, new_n18482_,
    new_n18483_, new_n18485_, new_n18486_, new_n18487_, new_n18488_,
    new_n18489_, new_n18490_, new_n18491_, new_n18492_, new_n18493_,
    new_n18494_, new_n18495_, new_n18496_, new_n18497_, new_n18498_,
    new_n18499_, new_n18500_, new_n18501_, new_n18502_, new_n18503_,
    new_n18504_, new_n18505_, new_n18506_, new_n18507_, new_n18508_,
    new_n18509_, new_n18510_, new_n18511_, new_n18512_, new_n18513_,
    new_n18514_, new_n18515_, new_n18516_, new_n18517_, new_n18518_,
    new_n18519_, new_n18520_, new_n18521_, new_n18522_, new_n18523_,
    new_n18524_, new_n18525_, new_n18526_, new_n18527_, new_n18528_,
    new_n18529_, new_n18530_, new_n18531_, new_n18532_, new_n18533_,
    new_n18534_, new_n18535_, new_n18536_, new_n18537_, new_n18538_,
    new_n18539_, new_n18540_, new_n18541_, new_n18542_, new_n18543_,
    new_n18544_, new_n18545_, new_n18546_, new_n18547_, new_n18548_,
    new_n18549_, new_n18550_, new_n18551_, new_n18552_, new_n18553_,
    new_n18554_, new_n18555_, new_n18556_, new_n18557_, new_n18558_,
    new_n18559_, new_n18560_, new_n18561_, new_n18562_, new_n18563_,
    new_n18564_, new_n18565_, new_n18566_, new_n18567_, new_n18568_,
    new_n18569_, new_n18570_, new_n18571_, new_n18572_, new_n18573_,
    new_n18574_, new_n18575_, new_n18576_, new_n18577_, new_n18578_,
    new_n18579_, new_n18580_, new_n18581_, new_n18582_, new_n18583_,
    new_n18584_, new_n18585_, new_n18586_, new_n18587_, new_n18588_,
    new_n18589_, new_n18590_, new_n18591_, new_n18592_, new_n18593_,
    new_n18594_, new_n18595_, new_n18596_, new_n18597_, new_n18598_,
    new_n18599_, new_n18600_, new_n18601_, new_n18602_, new_n18603_,
    new_n18604_, new_n18605_, new_n18606_, new_n18607_, new_n18608_,
    new_n18609_, new_n18610_, new_n18611_, new_n18612_, new_n18613_,
    new_n18614_, new_n18615_, new_n18616_, new_n18617_, new_n18618_,
    new_n18619_, new_n18620_, new_n18621_, new_n18622_, new_n18623_,
    new_n18624_, new_n18625_, new_n18626_, new_n18627_, new_n18628_,
    new_n18629_, new_n18630_, new_n18631_, new_n18632_, new_n18633_,
    new_n18634_, new_n18635_, new_n18636_, new_n18637_, new_n18638_,
    new_n18639_, new_n18640_, new_n18641_, new_n18642_, new_n18643_,
    new_n18644_, new_n18645_, new_n18646_, new_n18647_, new_n18648_,
    new_n18649_, new_n18650_, new_n18651_, new_n18652_, new_n18653_,
    new_n18654_, new_n18655_, new_n18656_, new_n18657_, new_n18658_,
    new_n18659_, new_n18660_, new_n18661_, new_n18662_, new_n18663_,
    new_n18664_, new_n18665_, new_n18666_, new_n18667_, new_n18668_,
    new_n18669_, new_n18670_, new_n18671_, new_n18672_, new_n18673_,
    new_n18674_, new_n18675_, new_n18676_, new_n18677_, new_n18678_,
    new_n18679_, new_n18680_, new_n18681_, new_n18682_, new_n18683_,
    new_n18684_, new_n18685_, new_n18686_, new_n18687_, new_n18688_,
    new_n18689_, new_n18690_, new_n18691_, new_n18692_, new_n18693_,
    new_n18694_, new_n18695_, new_n18696_, new_n18697_, new_n18698_,
    new_n18699_, new_n18700_, new_n18701_, new_n18702_, new_n18703_,
    new_n18704_, new_n18705_, new_n18706_, new_n18707_, new_n18708_,
    new_n18709_, new_n18710_, new_n18711_, new_n18712_, new_n18713_,
    new_n18714_, new_n18715_, new_n18716_, new_n18717_, new_n18718_,
    new_n18719_, new_n18720_, new_n18721_, new_n18722_, new_n18723_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19112_, new_n19113_, new_n19114_, new_n19115_,
    new_n19116_, new_n19117_, new_n19118_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19124_, new_n19125_,
    new_n19126_, new_n19127_, new_n19128_, new_n19129_, new_n19130_,
    new_n19131_, new_n19132_, new_n19133_, new_n19134_, new_n19135_,
    new_n19136_, new_n19137_, new_n19138_, new_n19139_, new_n19140_,
    new_n19141_, new_n19142_, new_n19143_, new_n19144_, new_n19145_,
    new_n19146_, new_n19147_, new_n19148_, new_n19149_, new_n19150_,
    new_n19151_, new_n19152_, new_n19153_, new_n19154_, new_n19155_,
    new_n19156_, new_n19157_, new_n19158_, new_n19159_, new_n19160_,
    new_n19161_, new_n19162_, new_n19163_, new_n19164_, new_n19165_,
    new_n19166_, new_n19167_, new_n19168_, new_n19169_, new_n19170_,
    new_n19171_, new_n19172_, new_n19173_, new_n19174_, new_n19175_,
    new_n19176_, new_n19177_, new_n19178_, new_n19179_, new_n19180_,
    new_n19181_, new_n19182_, new_n19183_, new_n19184_, new_n19185_,
    new_n19186_, new_n19187_, new_n19188_, new_n19189_, new_n19190_,
    new_n19191_, new_n19192_, new_n19193_, new_n19194_, new_n19195_,
    new_n19196_, new_n19197_, new_n19198_, new_n19199_, new_n19200_,
    new_n19201_, new_n19202_, new_n19203_, new_n19204_, new_n19205_,
    new_n19206_, new_n19207_, new_n19208_, new_n19209_, new_n19210_,
    new_n19211_, new_n19212_, new_n19213_, new_n19214_, new_n19215_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19227_, new_n19228_, new_n19229_, new_n19230_, new_n19231_,
    new_n19232_, new_n19233_, new_n19234_, new_n19235_, new_n19236_,
    new_n19237_, new_n19238_, new_n19239_, new_n19240_, new_n19241_,
    new_n19242_, new_n19243_, new_n19244_, new_n19245_, new_n19246_,
    new_n19247_, new_n19248_, new_n19249_, new_n19250_, new_n19251_,
    new_n19252_, new_n19253_, new_n19254_, new_n19255_, new_n19256_,
    new_n19257_, new_n19258_, new_n19259_, new_n19260_, new_n19261_,
    new_n19262_, new_n19263_, new_n19264_, new_n19265_, new_n19266_,
    new_n19267_, new_n19268_, new_n19269_, new_n19270_, new_n19271_,
    new_n19272_, new_n19273_, new_n19274_, new_n19275_, new_n19276_,
    new_n19277_, new_n19278_, new_n19279_, new_n19280_, new_n19281_,
    new_n19282_, new_n19283_, new_n19284_, new_n19285_, new_n19286_,
    new_n19287_, new_n19288_, new_n19289_, new_n19290_, new_n19291_,
    new_n19292_, new_n19293_, new_n19294_, new_n19295_, new_n19296_,
    new_n19297_, new_n19298_, new_n19299_, new_n19300_, new_n19301_,
    new_n19302_, new_n19303_, new_n19304_, new_n19305_, new_n19306_,
    new_n19307_, new_n19308_, new_n19309_, new_n19310_, new_n19311_,
    new_n19312_, new_n19313_, new_n19314_, new_n19315_, new_n19316_,
    new_n19317_, new_n19318_, new_n19319_, new_n19320_, new_n19321_,
    new_n19322_, new_n19323_, new_n19324_, new_n19325_, new_n19326_,
    new_n19327_, new_n19328_, new_n19329_, new_n19330_, new_n19331_,
    new_n19332_, new_n19333_, new_n19334_, new_n19335_, new_n19336_,
    new_n19337_, new_n19338_, new_n19339_, new_n19340_, new_n19341_,
    new_n19342_, new_n19343_, new_n19344_, new_n19345_, new_n19346_,
    new_n19347_, new_n19348_, new_n19349_, new_n19350_, new_n19351_,
    new_n19352_, new_n19353_, new_n19354_, new_n19355_, new_n19356_,
    new_n19357_, new_n19358_, new_n19359_, new_n19360_, new_n19361_,
    new_n19362_, new_n19363_, new_n19364_, new_n19365_, new_n19366_,
    new_n19367_, new_n19368_, new_n19369_, new_n19370_, new_n19371_,
    new_n19372_, new_n19373_, new_n19374_, new_n19375_, new_n19376_,
    new_n19377_, new_n19378_, new_n19379_, new_n19380_, new_n19381_,
    new_n19382_, new_n19383_, new_n19384_, new_n19385_, new_n19386_,
    new_n19387_, new_n19388_, new_n19389_, new_n19390_, new_n19391_,
    new_n19392_, new_n19393_, new_n19394_, new_n19395_, new_n19396_,
    new_n19397_, new_n19398_, new_n19399_, new_n19400_, new_n19401_,
    new_n19402_, new_n19403_, new_n19404_, new_n19405_, new_n19406_,
    new_n19407_, new_n19408_, new_n19409_, new_n19410_, new_n19411_,
    new_n19412_, new_n19413_, new_n19414_, new_n19415_, new_n19416_,
    new_n19417_, new_n19418_, new_n19419_, new_n19420_, new_n19421_,
    new_n19422_, new_n19423_, new_n19424_, new_n19425_, new_n19426_,
    new_n19427_, new_n19428_, new_n19429_, new_n19430_, new_n19431_,
    new_n19432_, new_n19433_, new_n19434_, new_n19435_, new_n19436_,
    new_n19437_, new_n19438_, new_n19439_, new_n19441_, new_n19442_,
    new_n19443_, new_n19444_, new_n19445_, new_n19446_, new_n19447_,
    new_n19448_, new_n19449_, new_n19450_, new_n19451_, new_n19452_,
    new_n19453_, new_n19454_, new_n19455_, new_n19456_, new_n19457_,
    new_n19458_, new_n19459_, new_n19460_, new_n19461_, new_n19462_,
    new_n19463_, new_n19464_, new_n19465_, new_n19466_, new_n19467_,
    new_n19468_, new_n19469_, new_n19470_, new_n19471_, new_n19472_,
    new_n19473_, new_n19474_, new_n19475_, new_n19476_, new_n19477_,
    new_n19478_, new_n19479_, new_n19480_, new_n19481_, new_n19482_,
    new_n19483_, new_n19484_, new_n19485_, new_n19486_, new_n19487_,
    new_n19488_, new_n19489_, new_n19490_, new_n19491_, new_n19492_,
    new_n19493_, new_n19494_, new_n19495_, new_n19496_, new_n19497_,
    new_n19498_, new_n19499_, new_n19500_, new_n19501_, new_n19502_,
    new_n19503_, new_n19504_, new_n19505_, new_n19506_, new_n19507_,
    new_n19508_, new_n19509_, new_n19510_, new_n19511_, new_n19512_,
    new_n19513_, new_n19514_, new_n19515_, new_n19516_, new_n19517_,
    new_n19518_, new_n19519_, new_n19520_, new_n19521_, new_n19522_,
    new_n19523_, new_n19524_, new_n19525_, new_n19526_, new_n19527_,
    new_n19528_, new_n19529_, new_n19530_, new_n19531_, new_n19532_,
    new_n19533_, new_n19534_, new_n19535_, new_n19536_, new_n19537_,
    new_n19538_, new_n19539_, new_n19540_, new_n19541_, new_n19542_,
    new_n19543_, new_n19544_, new_n19545_, new_n19546_, new_n19547_,
    new_n19548_, new_n19549_, new_n19550_, new_n19551_, new_n19552_,
    new_n19553_, new_n19554_, new_n19555_, new_n19556_, new_n19557_,
    new_n19558_, new_n19559_, new_n19560_, new_n19561_, new_n19562_,
    new_n19563_, new_n19564_, new_n19565_, new_n19566_, new_n19567_,
    new_n19568_, new_n19569_, new_n19570_, new_n19571_, new_n19572_,
    new_n19573_, new_n19574_, new_n19575_, new_n19576_, new_n19577_,
    new_n19578_, new_n19579_, new_n19580_, new_n19581_, new_n19582_,
    new_n19583_, new_n19584_, new_n19585_, new_n19586_, new_n19587_,
    new_n19588_, new_n19589_, new_n19590_, new_n19591_, new_n19592_,
    new_n19593_, new_n19594_, new_n19595_, new_n19596_, new_n19597_,
    new_n19598_, new_n19599_, new_n19600_, new_n19601_, new_n19602_,
    new_n19603_, new_n19604_, new_n19605_, new_n19606_, new_n19607_,
    new_n19608_, new_n19609_, new_n19610_, new_n19611_, new_n19612_,
    new_n19613_, new_n19614_, new_n19615_, new_n19616_, new_n19617_,
    new_n19618_, new_n19619_, new_n19620_, new_n19621_, new_n19622_,
    new_n19623_, new_n19624_, new_n19625_, new_n19626_, new_n19627_,
    new_n19628_, new_n19629_, new_n19630_, new_n19631_, new_n19632_,
    new_n19633_, new_n19634_, new_n19635_, new_n19636_, new_n19637_,
    new_n19638_, new_n19639_, new_n19640_, new_n19641_, new_n19642_,
    new_n19643_, new_n19644_, new_n19645_, new_n19646_, new_n19647_,
    new_n19648_, new_n19649_, new_n19650_, new_n19651_, new_n19652_,
    new_n19653_, new_n19654_, new_n19656_, new_n19657_, new_n19658_,
    new_n19659_, new_n19660_, new_n19661_, new_n19662_, new_n19663_,
    new_n19664_, new_n19665_, new_n19666_, new_n19667_, new_n19668_,
    new_n19669_, new_n19670_, new_n19671_, new_n19672_, new_n19673_,
    new_n19674_, new_n19675_, new_n19676_, new_n19677_, new_n19678_,
    new_n19679_, new_n19680_, new_n19681_, new_n19682_, new_n19683_,
    new_n19684_, new_n19685_, new_n19686_, new_n19687_, new_n19688_,
    new_n19689_, new_n19690_, new_n19691_, new_n19692_, new_n19693_,
    new_n19694_, new_n19695_, new_n19696_, new_n19697_, new_n19698_,
    new_n19699_, new_n19700_, new_n19701_, new_n19702_, new_n19703_,
    new_n19704_, new_n19705_, new_n19706_, new_n19707_, new_n19708_,
    new_n19709_, new_n19710_, new_n19711_, new_n19712_, new_n19713_,
    new_n19714_, new_n19715_, new_n19716_, new_n19717_, new_n19718_,
    new_n19719_, new_n19720_, new_n19721_, new_n19722_, new_n19723_,
    new_n19724_, new_n19725_, new_n19726_, new_n19727_, new_n19728_,
    new_n19729_, new_n19730_, new_n19731_, new_n19732_, new_n19733_,
    new_n19734_, new_n19735_, new_n19736_, new_n19737_, new_n19738_,
    new_n19739_, new_n19740_, new_n19741_, new_n19742_, new_n19743_,
    new_n19744_, new_n19745_, new_n19746_, new_n19747_, new_n19748_,
    new_n19749_, new_n19750_, new_n19751_, new_n19752_, new_n19753_,
    new_n19754_, new_n19755_, new_n19756_, new_n19757_, new_n19758_,
    new_n19759_, new_n19760_, new_n19761_, new_n19762_, new_n19763_,
    new_n19764_, new_n19765_, new_n19766_, new_n19767_, new_n19768_,
    new_n19769_, new_n19770_, new_n19771_, new_n19772_, new_n19773_,
    new_n19774_, new_n19775_, new_n19776_, new_n19777_, new_n19778_,
    new_n19779_, new_n19780_, new_n19781_, new_n19782_, new_n19783_,
    new_n19784_, new_n19785_, new_n19786_, new_n19787_, new_n19788_,
    new_n19789_, new_n19790_, new_n19791_, new_n19792_, new_n19793_,
    new_n19794_, new_n19795_, new_n19796_, new_n19797_, new_n19798_,
    new_n19799_, new_n19800_, new_n19801_, new_n19802_, new_n19803_,
    new_n19804_, new_n19805_, new_n19806_, new_n19807_, new_n19808_,
    new_n19809_, new_n19810_, new_n19811_, new_n19812_, new_n19813_,
    new_n19814_, new_n19815_, new_n19816_, new_n19817_, new_n19818_,
    new_n19819_, new_n19820_, new_n19821_, new_n19822_, new_n19823_,
    new_n19824_, new_n19825_, new_n19826_, new_n19827_, new_n19828_,
    new_n19829_, new_n19830_, new_n19831_, new_n19832_, new_n19833_,
    new_n19834_, new_n19835_, new_n19836_, new_n19837_, new_n19838_,
    new_n19839_, new_n19840_, new_n19841_, new_n19842_, new_n19843_,
    new_n19844_, new_n19845_, new_n19846_, new_n19847_, new_n19848_,
    new_n19849_, new_n19850_, new_n19851_, new_n19852_, new_n19853_,
    new_n19854_, new_n19855_, new_n19856_, new_n19857_, new_n19858_,
    new_n19859_, new_n19860_, new_n19861_, new_n19862_, new_n19863_,
    new_n19864_, new_n19865_, new_n19866_, new_n19867_, new_n19868_,
    new_n19869_, new_n19870_, new_n19871_, new_n19872_, new_n19873_,
    new_n19874_, new_n19875_, new_n19876_, new_n19877_, new_n19878_,
    new_n19879_, new_n19880_, new_n19881_, new_n19882_, new_n19883_,
    new_n19884_, new_n19885_, new_n19886_, new_n19888_, new_n19889_,
    new_n19890_, new_n19891_, new_n19892_, new_n19893_, new_n19894_,
    new_n19895_, new_n19896_, new_n19897_, new_n19898_, new_n19899_,
    new_n19900_, new_n19901_, new_n19902_, new_n19903_, new_n19904_,
    new_n19905_, new_n19906_, new_n19907_, new_n19908_, new_n19909_,
    new_n19910_, new_n19911_, new_n19912_, new_n19913_, new_n19914_,
    new_n19915_, new_n19916_, new_n19917_, new_n19918_, new_n19919_,
    new_n19920_, new_n19921_, new_n19922_, new_n19923_, new_n19924_,
    new_n19925_, new_n19926_, new_n19927_, new_n19928_, new_n19929_,
    new_n19930_, new_n19931_, new_n19932_, new_n19933_, new_n19934_,
    new_n19935_, new_n19936_, new_n19937_, new_n19938_, new_n19939_,
    new_n19940_, new_n19941_, new_n19942_, new_n19943_, new_n19944_,
    new_n19945_, new_n19946_, new_n19947_, new_n19948_, new_n19949_,
    new_n19950_, new_n19951_, new_n19952_, new_n19953_, new_n19954_,
    new_n19955_, new_n19956_, new_n19957_, new_n19958_, new_n19959_,
    new_n19960_, new_n19961_, new_n19962_, new_n19963_, new_n19964_,
    new_n19965_, new_n19966_, new_n19967_, new_n19968_, new_n19969_,
    new_n19970_, new_n19971_, new_n19972_, new_n19973_, new_n19974_,
    new_n19975_, new_n19976_, new_n19977_, new_n19978_, new_n19979_,
    new_n19980_, new_n19981_, new_n19982_, new_n19983_, new_n19984_,
    new_n19985_, new_n19986_, new_n19987_, new_n19988_, new_n19989_,
    new_n19990_, new_n19991_, new_n19992_, new_n19993_, new_n19994_,
    new_n19995_, new_n19996_, new_n19997_, new_n19998_, new_n19999_,
    new_n20000_, new_n20001_, new_n20002_, new_n20003_, new_n20004_,
    new_n20005_, new_n20006_, new_n20007_, new_n20008_, new_n20009_,
    new_n20010_, new_n20011_, new_n20012_, new_n20013_, new_n20014_,
    new_n20015_, new_n20016_, new_n20017_, new_n20018_, new_n20019_,
    new_n20020_, new_n20021_, new_n20022_, new_n20023_, new_n20024_,
    new_n20025_, new_n20026_, new_n20027_, new_n20028_, new_n20029_,
    new_n20030_, new_n20031_, new_n20032_, new_n20033_, new_n20034_,
    new_n20035_, new_n20036_, new_n20037_, new_n20038_, new_n20039_,
    new_n20040_, new_n20041_, new_n20042_, new_n20043_, new_n20044_,
    new_n20045_, new_n20046_, new_n20047_, new_n20048_, new_n20049_,
    new_n20050_, new_n20051_, new_n20052_, new_n20053_, new_n20054_,
    new_n20055_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20104_, new_n20105_,
    new_n20106_, new_n20107_, new_n20108_, new_n20109_, new_n20110_,
    new_n20111_, new_n20112_, new_n20113_, new_n20114_, new_n20115_,
    new_n20116_, new_n20117_, new_n20118_, new_n20119_, new_n20120_,
    new_n20121_, new_n20122_, new_n20123_, new_n20124_, new_n20125_,
    new_n20126_, new_n20127_, new_n20128_, new_n20129_, new_n20130_,
    new_n20131_, new_n20132_, new_n20133_, new_n20134_, new_n20135_,
    new_n20136_, new_n20137_, new_n20138_, new_n20139_, new_n20140_,
    new_n20141_, new_n20142_, new_n20143_, new_n20144_, new_n20145_,
    new_n20146_, new_n20147_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20199_, new_n20200_,
    new_n20201_, new_n20202_, new_n20203_, new_n20204_, new_n20205_,
    new_n20206_, new_n20207_, new_n20208_, new_n20209_, new_n20210_,
    new_n20211_, new_n20212_, new_n20213_, new_n20214_, new_n20215_,
    new_n20216_, new_n20217_, new_n20218_, new_n20219_, new_n20220_,
    new_n20221_, new_n20222_, new_n20223_, new_n20224_, new_n20225_,
    new_n20226_, new_n20227_, new_n20228_, new_n20229_, new_n20230_,
    new_n20231_, new_n20232_, new_n20233_, new_n20234_, new_n20235_,
    new_n20236_, new_n20237_, new_n20238_, new_n20239_, new_n20240_,
    new_n20241_, new_n20242_, new_n20243_, new_n20244_, new_n20245_,
    new_n20246_, new_n20247_, new_n20248_, new_n20249_, new_n20250_,
    new_n20251_, new_n20252_, new_n20253_, new_n20254_, new_n20255_,
    new_n20256_, new_n20257_, new_n20258_, new_n20259_, new_n20260_,
    new_n20261_, new_n20262_, new_n20263_, new_n20264_, new_n20265_,
    new_n20266_, new_n20267_, new_n20268_, new_n20269_, new_n20270_,
    new_n20271_, new_n20272_, new_n20273_, new_n20274_, new_n20275_,
    new_n20276_, new_n20277_, new_n20278_, new_n20279_, new_n20280_,
    new_n20281_, new_n20282_, new_n20283_, new_n20284_, new_n20285_,
    new_n20286_, new_n20287_, new_n20288_, new_n20289_, new_n20290_,
    new_n20291_, new_n20292_, new_n20293_, new_n20294_, new_n20295_,
    new_n20296_, new_n20297_, new_n20298_, new_n20299_, new_n20300_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20321_,
    new_n20322_, new_n20323_, new_n20324_, new_n20325_, new_n20326_,
    new_n20327_, new_n20328_, new_n20329_, new_n20330_, new_n20331_,
    new_n20332_, new_n20333_, new_n20334_, new_n20335_, new_n20336_,
    new_n20337_, new_n20338_, new_n20339_, new_n20340_, new_n20341_,
    new_n20342_, new_n20343_, new_n20344_, new_n20345_, new_n20346_,
    new_n20347_, new_n20348_, new_n20349_, new_n20350_, new_n20351_,
    new_n20352_, new_n20353_, new_n20354_, new_n20355_, new_n20356_,
    new_n20357_, new_n20358_, new_n20359_, new_n20360_, new_n20361_,
    new_n20362_, new_n20363_, new_n20364_, new_n20365_, new_n20366_,
    new_n20367_, new_n20368_, new_n20369_, new_n20370_, new_n20371_,
    new_n20372_, new_n20373_, new_n20374_, new_n20375_, new_n20376_,
    new_n20377_, new_n20378_, new_n20379_, new_n20380_, new_n20381_,
    new_n20382_, new_n20383_, new_n20384_, new_n20385_, new_n20386_,
    new_n20387_, new_n20388_, new_n20389_, new_n20390_, new_n20391_,
    new_n20392_, new_n20393_, new_n20394_, new_n20395_, new_n20396_,
    new_n20397_, new_n20398_, new_n20399_, new_n20400_, new_n20401_,
    new_n20402_, new_n20403_, new_n20404_, new_n20405_, new_n20406_,
    new_n20407_, new_n20408_, new_n20409_, new_n20410_, new_n20411_,
    new_n20412_, new_n20413_, new_n20414_, new_n20415_, new_n20416_,
    new_n20417_, new_n20418_, new_n20419_, new_n20420_, new_n20421_,
    new_n20422_, new_n20423_, new_n20424_, new_n20425_, new_n20426_,
    new_n20427_, new_n20428_, new_n20429_, new_n20430_, new_n20431_,
    new_n20432_, new_n20433_, new_n20434_, new_n20435_, new_n20436_,
    new_n20437_, new_n20438_, new_n20439_, new_n20440_, new_n20441_,
    new_n20442_, new_n20443_, new_n20444_, new_n20445_, new_n20446_,
    new_n20447_, new_n20448_, new_n20449_, new_n20450_, new_n20451_,
    new_n20452_, new_n20453_, new_n20454_, new_n20455_, new_n20456_,
    new_n20457_, new_n20458_, new_n20459_, new_n20460_, new_n20461_,
    new_n20462_, new_n20463_, new_n20464_, new_n20465_, new_n20466_,
    new_n20467_, new_n20468_, new_n20469_, new_n20470_, new_n20471_,
    new_n20472_, new_n20473_, new_n20474_, new_n20475_, new_n20476_,
    new_n20477_, new_n20478_, new_n20479_, new_n20480_, new_n20481_,
    new_n20482_, new_n20483_, new_n20484_, new_n20485_, new_n20486_,
    new_n20487_, new_n20488_, new_n20489_, new_n20490_, new_n20491_,
    new_n20492_, new_n20493_, new_n20494_, new_n20495_, new_n20496_,
    new_n20497_, new_n20498_, new_n20499_, new_n20500_, new_n20501_,
    new_n20502_, new_n20503_, new_n20504_, new_n20505_, new_n20506_,
    new_n20507_, new_n20508_, new_n20509_, new_n20511_, new_n20512_,
    new_n20513_, new_n20514_, new_n20515_, new_n20516_, new_n20517_,
    new_n20518_, new_n20519_, new_n20520_, new_n20521_, new_n20522_,
    new_n20523_, new_n20524_, new_n20525_, new_n20526_, new_n20527_,
    new_n20528_, new_n20529_, new_n20530_, new_n20531_, new_n20532_,
    new_n20533_, new_n20534_, new_n20535_, new_n20536_, new_n20537_,
    new_n20538_, new_n20539_, new_n20540_, new_n20541_, new_n20542_,
    new_n20543_, new_n20544_, new_n20545_, new_n20546_, new_n20547_,
    new_n20548_, new_n20549_, new_n20550_, new_n20551_, new_n20552_,
    new_n20553_, new_n20554_, new_n20555_, new_n20556_, new_n20557_,
    new_n20558_, new_n20559_, new_n20560_, new_n20561_, new_n20562_,
    new_n20563_, new_n20564_, new_n20565_, new_n20566_, new_n20567_,
    new_n20568_, new_n20569_, new_n20570_, new_n20571_, new_n20572_,
    new_n20573_, new_n20574_, new_n20575_, new_n20576_, new_n20577_,
    new_n20578_, new_n20579_, new_n20580_, new_n20581_, new_n20582_,
    new_n20583_, new_n20584_, new_n20585_, new_n20586_, new_n20587_,
    new_n20588_, new_n20589_, new_n20590_, new_n20591_, new_n20592_,
    new_n20593_, new_n20594_, new_n20595_, new_n20596_, new_n20597_,
    new_n20598_, new_n20599_, new_n20600_, new_n20601_, new_n20602_,
    new_n20603_, new_n20604_, new_n20605_, new_n20606_, new_n20607_,
    new_n20608_, new_n20609_, new_n20610_, new_n20611_, new_n20612_,
    new_n20613_, new_n20614_, new_n20615_, new_n20616_, new_n20617_,
    new_n20618_, new_n20619_, new_n20620_, new_n20621_, new_n20622_,
    new_n20623_, new_n20624_, new_n20625_, new_n20626_, new_n20627_,
    new_n20628_, new_n20629_, new_n20630_, new_n20631_, new_n20632_,
    new_n20633_, new_n20634_, new_n20635_, new_n20636_, new_n20637_,
    new_n20638_, new_n20639_, new_n20640_, new_n20641_, new_n20642_,
    new_n20643_, new_n20644_, new_n20645_, new_n20646_, new_n20647_,
    new_n20648_, new_n20649_, new_n20650_, new_n20651_, new_n20652_,
    new_n20653_, new_n20654_, new_n20655_, new_n20656_, new_n20657_,
    new_n20658_, new_n20659_, new_n20660_, new_n20661_, new_n20662_,
    new_n20663_, new_n20664_, new_n20665_, new_n20666_, new_n20667_,
    new_n20668_, new_n20669_, new_n20670_, new_n20671_, new_n20672_,
    new_n20673_, new_n20674_, new_n20675_, new_n20676_, new_n20677_,
    new_n20678_, new_n20679_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20714_, new_n20715_, new_n20716_, new_n20717_, new_n20718_,
    new_n20719_, new_n20720_, new_n20721_, new_n20722_, new_n20723_,
    new_n20724_, new_n20725_, new_n20726_, new_n20727_, new_n20728_,
    new_n20729_, new_n20730_, new_n20731_, new_n20732_, new_n20733_,
    new_n20734_, new_n20735_, new_n20736_, new_n20737_, new_n20738_,
    new_n20739_, new_n20740_, new_n20741_, new_n20742_, new_n20743_,
    new_n20744_, new_n20745_, new_n20746_, new_n20747_, new_n20748_,
    new_n20749_, new_n20750_, new_n20751_, new_n20752_, new_n20753_,
    new_n20754_, new_n20755_, new_n20756_, new_n20757_, new_n20758_,
    new_n20759_, new_n20760_, new_n20761_, new_n20762_, new_n20763_,
    new_n20764_, new_n20765_, new_n20766_, new_n20767_, new_n20768_,
    new_n20769_, new_n20770_, new_n20771_, new_n20772_, new_n20773_,
    new_n20774_, new_n20775_, new_n20776_, new_n20777_, new_n20778_,
    new_n20779_, new_n20780_, new_n20781_, new_n20782_, new_n20783_,
    new_n20784_, new_n20785_, new_n20786_, new_n20787_, new_n20788_,
    new_n20789_, new_n20790_, new_n20791_, new_n20792_, new_n20793_,
    new_n20794_, new_n20795_, new_n20796_, new_n20797_, new_n20798_,
    new_n20799_, new_n20800_, new_n20801_, new_n20802_, new_n20803_,
    new_n20804_, new_n20805_, new_n20806_, new_n20807_, new_n20808_,
    new_n20809_, new_n20810_, new_n20811_, new_n20812_, new_n20813_,
    new_n20814_, new_n20815_, new_n20816_, new_n20817_, new_n20818_,
    new_n20819_, new_n20820_, new_n20821_, new_n20822_, new_n20823_,
    new_n20824_, new_n20825_, new_n20826_, new_n20827_, new_n20828_,
    new_n20829_, new_n20830_, new_n20831_, new_n20832_, new_n20833_,
    new_n20834_, new_n20835_, new_n20836_, new_n20837_, new_n20838_,
    new_n20839_, new_n20840_, new_n20841_, new_n20842_, new_n20843_,
    new_n20844_, new_n20845_, new_n20846_, new_n20847_, new_n20848_,
    new_n20849_, new_n20850_, new_n20851_, new_n20852_, new_n20853_,
    new_n20854_, new_n20855_, new_n20856_, new_n20857_, new_n20858_,
    new_n20859_, new_n20860_, new_n20861_, new_n20862_, new_n20863_,
    new_n20864_, new_n20865_, new_n20866_, new_n20867_, new_n20868_,
    new_n20869_, new_n20870_, new_n20871_, new_n20872_, new_n20873_,
    new_n20874_, new_n20875_, new_n20876_, new_n20877_, new_n20878_,
    new_n20879_, new_n20880_, new_n20881_, new_n20882_, new_n20883_,
    new_n20884_, new_n20885_, new_n20886_, new_n20887_, new_n20888_,
    new_n20889_, new_n20890_, new_n20891_, new_n20892_, new_n20893_,
    new_n20894_, new_n20895_, new_n20896_, new_n20897_, new_n20898_,
    new_n20899_, new_n20901_, new_n20902_, new_n20903_, new_n20904_,
    new_n20905_, new_n20906_, new_n20907_, new_n20908_, new_n20909_,
    new_n20910_, new_n20911_, new_n20912_, new_n20913_, new_n20914_,
    new_n20915_, new_n20916_, new_n20917_, new_n20918_, new_n20919_,
    new_n20920_, new_n20921_, new_n20922_, new_n20923_, new_n20924_,
    new_n20925_, new_n20926_, new_n20927_, new_n20928_, new_n20929_,
    new_n20930_, new_n20931_, new_n20932_, new_n20933_, new_n20934_,
    new_n20935_, new_n20936_, new_n20937_, new_n20938_, new_n20939_,
    new_n20940_, new_n20941_, new_n20942_, new_n20943_, new_n20944_,
    new_n20945_, new_n20946_, new_n20947_, new_n20948_, new_n20949_,
    new_n20950_, new_n20951_, new_n20952_, new_n20953_, new_n20954_,
    new_n20955_, new_n20956_, new_n20957_, new_n20958_, new_n20959_,
    new_n20960_, new_n20961_, new_n20962_, new_n20963_, new_n20964_,
    new_n20965_, new_n20966_, new_n20967_, new_n20968_, new_n20969_,
    new_n20970_, new_n20971_, new_n20972_, new_n20973_, new_n20974_,
    new_n20975_, new_n20976_, new_n20977_, new_n20978_, new_n20979_,
    new_n20980_, new_n20981_, new_n20982_, new_n20983_, new_n20984_,
    new_n20985_, new_n20986_, new_n20987_, new_n20988_, new_n20989_,
    new_n20990_, new_n20991_, new_n20992_, new_n20993_, new_n20994_,
    new_n20995_, new_n20996_, new_n20997_, new_n20998_, new_n20999_,
    new_n21000_, new_n21001_, new_n21002_, new_n21003_, new_n21004_,
    new_n21005_, new_n21006_, new_n21007_, new_n21008_, new_n21009_,
    new_n21010_, new_n21011_, new_n21012_, new_n21013_, new_n21014_,
    new_n21015_, new_n21016_, new_n21017_, new_n21018_, new_n21019_,
    new_n21020_, new_n21021_, new_n21022_, new_n21023_, new_n21024_,
    new_n21025_, new_n21026_, new_n21027_, new_n21028_, new_n21029_,
    new_n21030_, new_n21031_, new_n21032_, new_n21033_, new_n21034_,
    new_n21035_, new_n21036_, new_n21037_, new_n21038_, new_n21039_,
    new_n21040_, new_n21041_, new_n21042_, new_n21043_, new_n21044_,
    new_n21045_, new_n21046_, new_n21047_, new_n21048_, new_n21049_,
    new_n21050_, new_n21051_, new_n21052_, new_n21053_, new_n21054_,
    new_n21055_, new_n21056_, new_n21057_, new_n21058_, new_n21059_,
    new_n21060_, new_n21061_, new_n21062_, new_n21063_, new_n21064_,
    new_n21065_, new_n21066_, new_n21067_, new_n21068_, new_n21069_,
    new_n21070_, new_n21071_, new_n21072_, new_n21073_, new_n21074_,
    new_n21075_, new_n21076_, new_n21077_, new_n21078_, new_n21079_,
    new_n21080_, new_n21081_, new_n21082_, new_n21083_, new_n21084_,
    new_n21085_, new_n21086_, new_n21087_, new_n21088_, new_n21089_,
    new_n21090_, new_n21091_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21100_,
    new_n21101_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21385_, new_n21386_,
    new_n21387_, new_n21388_, new_n21389_, new_n21390_, new_n21391_,
    new_n21392_, new_n21393_, new_n21394_, new_n21395_, new_n21396_,
    new_n21397_, new_n21398_, new_n21399_, new_n21400_, new_n21401_,
    new_n21402_, new_n21403_, new_n21404_, new_n21405_, new_n21406_,
    new_n21407_, new_n21408_, new_n21409_, new_n21410_, new_n21411_,
    new_n21412_, new_n21413_, new_n21414_, new_n21415_, new_n21416_,
    new_n21417_, new_n21418_, new_n21419_, new_n21420_, new_n21421_,
    new_n21422_, new_n21423_, new_n21424_, new_n21425_, new_n21426_,
    new_n21427_, new_n21428_, new_n21429_, new_n21430_, new_n21431_,
    new_n21432_, new_n21433_, new_n21434_, new_n21435_, new_n21436_,
    new_n21437_, new_n21438_, new_n21439_, new_n21440_, new_n21441_,
    new_n21442_, new_n21443_, new_n21444_, new_n21445_, new_n21446_,
    new_n21447_, new_n21448_, new_n21449_, new_n21450_, new_n21451_,
    new_n21452_, new_n21453_, new_n21454_, new_n21455_, new_n21456_,
    new_n21457_, new_n21458_, new_n21459_, new_n21461_, new_n21462_,
    new_n21463_, new_n21464_, new_n21465_, new_n21466_, new_n21467_,
    new_n21468_, new_n21469_, new_n21470_, new_n21471_, new_n21472_,
    new_n21473_, new_n21474_, new_n21475_, new_n21476_, new_n21477_,
    new_n21478_, new_n21479_, new_n21480_, new_n21481_, new_n21482_,
    new_n21483_, new_n21484_, new_n21485_, new_n21486_, new_n21487_,
    new_n21488_, new_n21489_, new_n21490_, new_n21491_, new_n21492_,
    new_n21493_, new_n21494_, new_n21495_, new_n21496_, new_n21497_,
    new_n21498_, new_n21499_, new_n21500_, new_n21501_, new_n21502_,
    new_n21503_, new_n21504_, new_n21505_, new_n21506_, new_n21507_,
    new_n21508_, new_n21509_, new_n21510_, new_n21511_, new_n21512_,
    new_n21513_, new_n21514_, new_n21515_, new_n21516_, new_n21517_,
    new_n21518_, new_n21519_, new_n21520_, new_n21521_, new_n21522_,
    new_n21523_, new_n21524_, new_n21525_, new_n21526_, new_n21527_,
    new_n21528_, new_n21529_, new_n21530_, new_n21531_, new_n21532_,
    new_n21533_, new_n21534_, new_n21535_, new_n21536_, new_n21537_,
    new_n21538_, new_n21539_, new_n21540_, new_n21541_, new_n21542_,
    new_n21543_, new_n21544_, new_n21545_, new_n21546_, new_n21547_,
    new_n21548_, new_n21549_, new_n21550_, new_n21551_, new_n21552_,
    new_n21553_, new_n21554_, new_n21555_, new_n21556_, new_n21557_,
    new_n21558_, new_n21559_, new_n21560_, new_n21561_, new_n21562_,
    new_n21563_, new_n21564_, new_n21565_, new_n21566_, new_n21567_,
    new_n21568_, new_n21569_, new_n21570_, new_n21571_, new_n21572_,
    new_n21573_, new_n21574_, new_n21575_, new_n21576_, new_n21577_,
    new_n21578_, new_n21579_, new_n21580_, new_n21581_, new_n21582_,
    new_n21583_, new_n21584_, new_n21585_, new_n21586_, new_n21587_,
    new_n21588_, new_n21589_, new_n21590_, new_n21591_, new_n21592_,
    new_n21593_, new_n21594_, new_n21595_, new_n21596_, new_n21597_,
    new_n21598_, new_n21599_, new_n21600_, new_n21601_, new_n21602_,
    new_n21603_, new_n21604_, new_n21605_, new_n21606_, new_n21607_,
    new_n21608_, new_n21609_, new_n21610_, new_n21611_, new_n21612_,
    new_n21613_, new_n21614_, new_n21615_, new_n21616_, new_n21617_,
    new_n21618_, new_n21619_, new_n21620_, new_n21621_, new_n21622_,
    new_n21623_, new_n21624_, new_n21625_, new_n21626_, new_n21627_,
    new_n21628_, new_n21629_, new_n21630_, new_n21631_, new_n21632_,
    new_n21633_, new_n21634_, new_n21635_, new_n21636_, new_n21637_,
    new_n21638_, new_n21639_, new_n21641_, new_n21642_, new_n21643_,
    new_n21644_, new_n21645_, new_n21646_, new_n21647_, new_n21648_,
    new_n21649_, new_n21650_, new_n21651_, new_n21652_, new_n21653_,
    new_n21654_, new_n21655_, new_n21656_, new_n21657_, new_n21658_,
    new_n21659_, new_n21660_, new_n21661_, new_n21662_, new_n21663_,
    new_n21664_, new_n21665_, new_n21666_, new_n21667_, new_n21668_,
    new_n21669_, new_n21670_, new_n21671_, new_n21672_, new_n21673_,
    new_n21674_, new_n21675_, new_n21676_, new_n21677_, new_n21678_,
    new_n21679_, new_n21680_, new_n21681_, new_n21682_, new_n21683_,
    new_n21684_, new_n21685_, new_n21686_, new_n21687_, new_n21688_,
    new_n21689_, new_n21690_, new_n21691_, new_n21692_, new_n21693_,
    new_n21694_, new_n21695_, new_n21696_, new_n21697_, new_n21698_,
    new_n21699_, new_n21700_, new_n21701_, new_n21702_, new_n21703_,
    new_n21704_, new_n21705_, new_n21706_, new_n21707_, new_n21708_,
    new_n21709_, new_n21710_, new_n21711_, new_n21712_, new_n21713_,
    new_n21714_, new_n21715_, new_n21716_, new_n21717_, new_n21718_,
    new_n21719_, new_n21720_, new_n21721_, new_n21722_, new_n21723_,
    new_n21724_, new_n21725_, new_n21726_, new_n21727_, new_n21728_,
    new_n21729_, new_n21730_, new_n21731_, new_n21732_, new_n21733_,
    new_n21734_, new_n21735_, new_n21736_, new_n21737_, new_n21738_,
    new_n21739_, new_n21740_, new_n21741_, new_n21742_, new_n21743_,
    new_n21744_, new_n21745_, new_n21746_, new_n21747_, new_n21748_,
    new_n21749_, new_n21750_, new_n21751_, new_n21752_, new_n21753_,
    new_n21754_, new_n21755_, new_n21756_, new_n21757_, new_n21758_,
    new_n21759_, new_n21760_, new_n21761_, new_n21762_, new_n21763_,
    new_n21764_, new_n21765_, new_n21766_, new_n21767_, new_n21768_,
    new_n21769_, new_n21770_, new_n21771_, new_n21772_, new_n21773_,
    new_n21774_, new_n21775_, new_n21776_, new_n21777_, new_n21778_,
    new_n21779_, new_n21780_, new_n21781_, new_n21782_, new_n21783_,
    new_n21784_, new_n21785_, new_n21786_, new_n21787_, new_n21788_,
    new_n21789_, new_n21790_, new_n21791_, new_n21792_, new_n21793_,
    new_n21794_, new_n21795_, new_n21796_, new_n21797_, new_n21798_,
    new_n21799_, new_n21800_, new_n21801_, new_n21802_, new_n21803_,
    new_n21804_, new_n21805_, new_n21806_, new_n21807_, new_n21808_,
    new_n21809_, new_n21810_, new_n21811_, new_n21812_, new_n21813_,
    new_n21814_, new_n21815_, new_n21816_, new_n21817_, new_n21818_,
    new_n21819_, new_n21821_, new_n21822_, new_n21823_, new_n21824_,
    new_n21825_, new_n21826_, new_n21827_, new_n21828_, new_n21829_,
    new_n21830_, new_n21831_, new_n21832_, new_n21833_, new_n21834_,
    new_n21835_, new_n21836_, new_n21837_, new_n21838_, new_n21839_,
    new_n21840_, new_n21841_, new_n21842_, new_n21843_, new_n21844_,
    new_n21845_, new_n21846_, new_n21847_, new_n21848_, new_n21849_,
    new_n21850_, new_n21851_, new_n21852_, new_n21853_, new_n21854_,
    new_n21855_, new_n21856_, new_n21857_, new_n21858_, new_n21859_,
    new_n21860_, new_n21861_, new_n21862_, new_n21863_, new_n21864_,
    new_n21865_, new_n21866_, new_n21867_, new_n21868_, new_n21869_,
    new_n21870_, new_n21871_, new_n21872_, new_n21873_, new_n21874_,
    new_n21875_, new_n21876_, new_n21877_, new_n21878_, new_n21879_,
    new_n21880_, new_n21881_, new_n21882_, new_n21883_, new_n21884_,
    new_n21885_, new_n21886_, new_n21887_, new_n21888_, new_n21889_,
    new_n21890_, new_n21891_, new_n21892_, new_n21893_, new_n21894_,
    new_n21895_, new_n21896_, new_n21897_, new_n21898_, new_n21899_,
    new_n21900_, new_n21901_, new_n21902_, new_n21903_, new_n21904_,
    new_n21905_, new_n21906_, new_n21907_, new_n21908_, new_n21909_,
    new_n21910_, new_n21911_, new_n21912_, new_n21913_, new_n21914_,
    new_n21915_, new_n21916_, new_n21917_, new_n21918_, new_n21919_,
    new_n21920_, new_n21921_, new_n21922_, new_n21923_, new_n21924_,
    new_n21925_, new_n21926_, new_n21927_, new_n21928_, new_n21929_,
    new_n21930_, new_n21931_, new_n21932_, new_n21933_, new_n21934_,
    new_n21935_, new_n21936_, new_n21937_, new_n21938_, new_n21939_,
    new_n21940_, new_n21941_, new_n21942_, new_n21943_, new_n21944_,
    new_n21945_, new_n21946_, new_n21947_, new_n21948_, new_n21949_,
    new_n21950_, new_n21951_, new_n21952_, new_n21953_, new_n21954_,
    new_n21955_, new_n21956_, new_n21957_, new_n21958_, new_n21959_,
    new_n21960_, new_n21961_, new_n21962_, new_n21963_, new_n21964_,
    new_n21965_, new_n21966_, new_n21967_, new_n21968_, new_n21969_,
    new_n21970_, new_n21971_, new_n21972_, new_n21973_, new_n21974_,
    new_n21975_, new_n21976_, new_n21977_, new_n21978_, new_n21979_,
    new_n21980_, new_n21981_, new_n21982_, new_n21983_, new_n21985_,
    new_n21986_, new_n21987_, new_n21988_, new_n21989_, new_n21990_,
    new_n21991_, new_n21992_, new_n21993_, new_n21994_, new_n21995_,
    new_n21996_, new_n21997_, new_n21998_, new_n21999_, new_n22000_,
    new_n22001_, new_n22002_, new_n22003_, new_n22004_, new_n22005_,
    new_n22006_, new_n22007_, new_n22008_, new_n22009_, new_n22010_,
    new_n22011_, new_n22012_, new_n22013_, new_n22014_, new_n22015_,
    new_n22016_, new_n22017_, new_n22018_, new_n22019_, new_n22020_,
    new_n22021_, new_n22022_, new_n22023_, new_n22024_, new_n22025_,
    new_n22026_, new_n22027_, new_n22028_, new_n22029_, new_n22030_,
    new_n22031_, new_n22032_, new_n22033_, new_n22034_, new_n22035_,
    new_n22036_, new_n22037_, new_n22038_, new_n22039_, new_n22040_,
    new_n22041_, new_n22042_, new_n22043_, new_n22044_, new_n22045_,
    new_n22046_, new_n22047_, new_n22048_, new_n22049_, new_n22050_,
    new_n22051_, new_n22052_, new_n22053_, new_n22054_, new_n22055_,
    new_n22056_, new_n22057_, new_n22058_, new_n22059_, new_n22060_,
    new_n22061_, new_n22062_, new_n22063_, new_n22064_, new_n22065_,
    new_n22066_, new_n22067_, new_n22068_, new_n22069_, new_n22070_,
    new_n22071_, new_n22072_, new_n22073_, new_n22074_, new_n22075_,
    new_n22076_, new_n22077_, new_n22078_, new_n22079_, new_n22080_,
    new_n22081_, new_n22082_, new_n22083_, new_n22084_, new_n22085_,
    new_n22086_, new_n22087_, new_n22088_, new_n22089_, new_n22090_,
    new_n22091_, new_n22092_, new_n22093_, new_n22094_, new_n22095_,
    new_n22096_, new_n22097_, new_n22098_, new_n22099_, new_n22100_,
    new_n22101_, new_n22102_, new_n22103_, new_n22104_, new_n22105_,
    new_n22106_, new_n22107_, new_n22108_, new_n22109_, new_n22110_,
    new_n22111_, new_n22112_, new_n22113_, new_n22114_, new_n22115_,
    new_n22116_, new_n22117_, new_n22118_, new_n22119_, new_n22120_,
    new_n22121_, new_n22122_, new_n22123_, new_n22124_, new_n22125_,
    new_n22126_, new_n22127_, new_n22128_, new_n22129_, new_n22130_,
    new_n22131_, new_n22132_, new_n22133_, new_n22134_, new_n22135_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22304_, new_n22305_, new_n22306_, new_n22307_,
    new_n22308_, new_n22309_, new_n22310_, new_n22311_, new_n22312_,
    new_n22313_, new_n22314_, new_n22315_, new_n22316_, new_n22317_,
    new_n22318_, new_n22319_, new_n22320_, new_n22321_, new_n22322_,
    new_n22323_, new_n22324_, new_n22325_, new_n22326_, new_n22327_,
    new_n22328_, new_n22329_, new_n22330_, new_n22331_, new_n22332_,
    new_n22333_, new_n22334_, new_n22335_, new_n22336_, new_n22337_,
    new_n22338_, new_n22339_, new_n22340_, new_n22341_, new_n22342_,
    new_n22343_, new_n22344_, new_n22345_, new_n22346_, new_n22347_,
    new_n22348_, new_n22349_, new_n22350_, new_n22351_, new_n22352_,
    new_n22353_, new_n22354_, new_n22355_, new_n22356_, new_n22357_,
    new_n22358_, new_n22359_, new_n22360_, new_n22361_, new_n22362_,
    new_n22363_, new_n22364_, new_n22365_, new_n22366_, new_n22367_,
    new_n22368_, new_n22369_, new_n22370_, new_n22371_, new_n22372_,
    new_n22373_, new_n22374_, new_n22375_, new_n22376_, new_n22377_,
    new_n22378_, new_n22379_, new_n22380_, new_n22381_, new_n22382_,
    new_n22383_, new_n22384_, new_n22385_, new_n22386_, new_n22387_,
    new_n22388_, new_n22389_, new_n22390_, new_n22391_, new_n22392_,
    new_n22393_, new_n22394_, new_n22395_, new_n22396_, new_n22397_,
    new_n22398_, new_n22399_, new_n22400_, new_n22401_, new_n22402_,
    new_n22403_, new_n22404_, new_n22405_, new_n22406_, new_n22407_,
    new_n22408_, new_n22409_, new_n22410_, new_n22411_, new_n22412_,
    new_n22413_, new_n22414_, new_n22415_, new_n22416_, new_n22417_,
    new_n22418_, new_n22419_, new_n22420_, new_n22421_, new_n22422_,
    new_n22423_, new_n22424_, new_n22425_, new_n22426_, new_n22427_,
    new_n22428_, new_n22429_, new_n22430_, new_n22431_, new_n22432_,
    new_n22433_, new_n22434_, new_n22435_, new_n22436_, new_n22437_,
    new_n22438_, new_n22439_, new_n22440_, new_n22441_, new_n22442_,
    new_n22443_, new_n22444_, new_n22445_, new_n22446_, new_n22447_,
    new_n22448_, new_n22449_, new_n22450_, new_n22451_, new_n22453_,
    new_n22454_, new_n22455_, new_n22456_, new_n22457_, new_n22458_,
    new_n22459_, new_n22460_, new_n22461_, new_n22462_, new_n22463_,
    new_n22464_, new_n22465_, new_n22466_, new_n22467_, new_n22468_,
    new_n22469_, new_n22470_, new_n22471_, new_n22472_, new_n22473_,
    new_n22474_, new_n22475_, new_n22476_, new_n22477_, new_n22478_,
    new_n22479_, new_n22480_, new_n22481_, new_n22482_, new_n22483_,
    new_n22484_, new_n22485_, new_n22486_, new_n22487_, new_n22488_,
    new_n22489_, new_n22490_, new_n22491_, new_n22492_, new_n22493_,
    new_n22494_, new_n22495_, new_n22496_, new_n22497_, new_n22498_,
    new_n22499_, new_n22500_, new_n22501_, new_n22502_, new_n22503_,
    new_n22504_, new_n22505_, new_n22506_, new_n22507_, new_n22508_,
    new_n22509_, new_n22510_, new_n22511_, new_n22512_, new_n22513_,
    new_n22514_, new_n22515_, new_n22516_, new_n22517_, new_n22518_,
    new_n22519_, new_n22520_, new_n22521_, new_n22522_, new_n22523_,
    new_n22524_, new_n22525_, new_n22526_, new_n22527_, new_n22528_,
    new_n22529_, new_n22530_, new_n22531_, new_n22532_, new_n22533_,
    new_n22534_, new_n22535_, new_n22536_, new_n22537_, new_n22538_,
    new_n22539_, new_n22540_, new_n22541_, new_n22542_, new_n22543_,
    new_n22544_, new_n22545_, new_n22546_, new_n22547_, new_n22548_,
    new_n22549_, new_n22550_, new_n22551_, new_n22552_, new_n22553_,
    new_n22554_, new_n22555_, new_n22556_, new_n22557_, new_n22558_,
    new_n22559_, new_n22560_, new_n22561_, new_n22562_, new_n22563_,
    new_n22564_, new_n22565_, new_n22566_, new_n22567_, new_n22568_,
    new_n22569_, new_n22570_, new_n22571_, new_n22572_, new_n22573_,
    new_n22574_, new_n22575_, new_n22576_, new_n22577_, new_n22578_,
    new_n22579_, new_n22580_, new_n22581_, new_n22582_, new_n22583_,
    new_n22584_, new_n22585_, new_n22586_, new_n22587_, new_n22588_,
    new_n22589_, new_n22590_, new_n22591_, new_n22592_, new_n22593_,
    new_n22594_, new_n22596_, new_n22597_, new_n22598_, new_n22599_,
    new_n22600_, new_n22601_, new_n22602_, new_n22603_, new_n22604_,
    new_n22605_, new_n22606_, new_n22607_, new_n22608_, new_n22609_,
    new_n22610_, new_n22611_, new_n22612_, new_n22613_, new_n22614_,
    new_n22615_, new_n22616_, new_n22617_, new_n22618_, new_n22619_,
    new_n22620_, new_n22621_, new_n22622_, new_n22623_, new_n22624_,
    new_n22625_, new_n22626_, new_n22627_, new_n22628_, new_n22629_,
    new_n22630_, new_n22631_, new_n22632_, new_n22633_, new_n22634_,
    new_n22635_, new_n22636_, new_n22637_, new_n22638_, new_n22639_,
    new_n22640_, new_n22641_, new_n22642_, new_n22643_, new_n22644_,
    new_n22645_, new_n22646_, new_n22647_, new_n22648_, new_n22649_,
    new_n22650_, new_n22651_, new_n22652_, new_n22653_, new_n22654_,
    new_n22655_, new_n22656_, new_n22657_, new_n22658_, new_n22659_,
    new_n22660_, new_n22661_, new_n22662_, new_n22663_, new_n22664_,
    new_n22665_, new_n22666_, new_n22667_, new_n22668_, new_n22669_,
    new_n22670_, new_n22671_, new_n22672_, new_n22673_, new_n22674_,
    new_n22675_, new_n22676_, new_n22677_, new_n22678_, new_n22679_,
    new_n22680_, new_n22681_, new_n22682_, new_n22683_, new_n22684_,
    new_n22685_, new_n22686_, new_n22687_, new_n22688_, new_n22689_,
    new_n22690_, new_n22691_, new_n22692_, new_n22693_, new_n22694_,
    new_n22695_, new_n22696_, new_n22697_, new_n22698_, new_n22699_,
    new_n22700_, new_n22701_, new_n22702_, new_n22703_, new_n22704_,
    new_n22705_, new_n22706_, new_n22707_, new_n22708_, new_n22709_,
    new_n22710_, new_n22711_, new_n22712_, new_n22713_, new_n22714_,
    new_n22715_, new_n22716_, new_n22717_, new_n22718_, new_n22719_,
    new_n22720_, new_n22721_, new_n22722_, new_n22723_, new_n22724_,
    new_n22725_, new_n22726_, new_n22727_, new_n22728_, new_n22729_,
    new_n22730_, new_n22731_, new_n22732_, new_n22733_, new_n22734_,
    new_n22735_, new_n22736_, new_n22737_, new_n22738_, new_n22739_,
    new_n22740_, new_n22741_, new_n22742_, new_n22743_, new_n22744_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22892_, new_n22893_, new_n22894_, new_n22895_, new_n22896_,
    new_n22897_, new_n22898_, new_n22899_, new_n22900_, new_n22901_,
    new_n22902_, new_n22903_, new_n22904_, new_n22905_, new_n22906_,
    new_n22907_, new_n22908_, new_n22909_, new_n22910_, new_n22911_,
    new_n22912_, new_n22913_, new_n22914_, new_n22915_, new_n22916_,
    new_n22917_, new_n22918_, new_n22919_, new_n22920_, new_n22921_,
    new_n22922_, new_n22923_, new_n22924_, new_n22925_, new_n22926_,
    new_n22927_, new_n22928_, new_n22929_, new_n22930_, new_n22931_,
    new_n22932_, new_n22933_, new_n22934_, new_n22935_, new_n22936_,
    new_n22937_, new_n22938_, new_n22939_, new_n22940_, new_n22941_,
    new_n22942_, new_n22943_, new_n22944_, new_n22945_, new_n22946_,
    new_n22947_, new_n22948_, new_n22949_, new_n22950_, new_n22951_,
    new_n22952_, new_n22953_, new_n22954_, new_n22955_, new_n22956_,
    new_n22957_, new_n22958_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23023_, new_n23024_, new_n23025_, new_n23026_,
    new_n23027_, new_n23028_, new_n23029_, new_n23031_, new_n23032_,
    new_n23033_, new_n23034_, new_n23035_, new_n23036_, new_n23037_,
    new_n23038_, new_n23039_, new_n23040_, new_n23041_, new_n23042_,
    new_n23043_, new_n23044_, new_n23045_, new_n23046_, new_n23047_,
    new_n23048_, new_n23049_, new_n23050_, new_n23051_, new_n23052_,
    new_n23053_, new_n23054_, new_n23055_, new_n23056_, new_n23057_,
    new_n23058_, new_n23059_, new_n23060_, new_n23061_, new_n23062_,
    new_n23063_, new_n23064_, new_n23065_, new_n23066_, new_n23067_,
    new_n23068_, new_n23069_, new_n23070_, new_n23071_, new_n23072_,
    new_n23073_, new_n23074_, new_n23075_, new_n23076_, new_n23077_,
    new_n23078_, new_n23079_, new_n23080_, new_n23081_, new_n23082_,
    new_n23083_, new_n23084_, new_n23085_, new_n23086_, new_n23087_,
    new_n23088_, new_n23089_, new_n23090_, new_n23091_, new_n23092_,
    new_n23093_, new_n23094_, new_n23095_, new_n23096_, new_n23097_,
    new_n23098_, new_n23099_, new_n23100_, new_n23101_, new_n23102_,
    new_n23103_, new_n23104_, new_n23105_, new_n23106_, new_n23107_,
    new_n23108_, new_n23109_, new_n23110_, new_n23111_, new_n23112_,
    new_n23113_, new_n23114_, new_n23115_, new_n23116_, new_n23117_,
    new_n23118_, new_n23119_, new_n23120_, new_n23121_, new_n23122_,
    new_n23123_, new_n23124_, new_n23125_, new_n23126_, new_n23127_,
    new_n23128_, new_n23129_, new_n23130_, new_n23131_, new_n23132_,
    new_n23133_, new_n23134_, new_n23135_, new_n23136_, new_n23137_,
    new_n23138_, new_n23139_, new_n23140_, new_n23141_, new_n23142_,
    new_n23143_, new_n23144_, new_n23145_, new_n23146_, new_n23147_,
    new_n23148_, new_n23149_, new_n23150_, new_n23151_, new_n23152_,
    new_n23153_, new_n23154_, new_n23155_, new_n23156_, new_n23157_,
    new_n23158_, new_n23159_, new_n23160_, new_n23161_, new_n23162_,
    new_n23163_, new_n23164_, new_n23165_, new_n23166_, new_n23167_,
    new_n23168_, new_n23170_, new_n23171_, new_n23172_, new_n23173_,
    new_n23174_, new_n23175_, new_n23176_, new_n23177_, new_n23178_,
    new_n23179_, new_n23180_, new_n23181_, new_n23182_, new_n23183_,
    new_n23184_, new_n23185_, new_n23186_, new_n23187_, new_n23188_,
    new_n23189_, new_n23190_, new_n23191_, new_n23192_, new_n23193_,
    new_n23194_, new_n23195_, new_n23196_, new_n23197_, new_n23198_,
    new_n23199_, new_n23200_, new_n23201_, new_n23202_, new_n23203_,
    new_n23204_, new_n23205_, new_n23206_, new_n23207_, new_n23208_,
    new_n23209_, new_n23210_, new_n23211_, new_n23212_, new_n23213_,
    new_n23214_, new_n23215_, new_n23216_, new_n23217_, new_n23218_,
    new_n23219_, new_n23220_, new_n23221_, new_n23222_, new_n23223_,
    new_n23224_, new_n23225_, new_n23226_, new_n23227_, new_n23228_,
    new_n23229_, new_n23230_, new_n23231_, new_n23232_, new_n23233_,
    new_n23234_, new_n23235_, new_n23236_, new_n23237_, new_n23238_,
    new_n23239_, new_n23240_, new_n23241_, new_n23242_, new_n23243_,
    new_n23244_, new_n23245_, new_n23246_, new_n23247_, new_n23248_,
    new_n23249_, new_n23250_, new_n23251_, new_n23252_, new_n23253_,
    new_n23254_, new_n23255_, new_n23256_, new_n23257_, new_n23258_,
    new_n23259_, new_n23260_, new_n23261_, new_n23262_, new_n23263_,
    new_n23264_, new_n23265_, new_n23266_, new_n23267_, new_n23268_,
    new_n23269_, new_n23270_, new_n23271_, new_n23272_, new_n23273_,
    new_n23274_, new_n23275_, new_n23276_, new_n23277_, new_n23278_,
    new_n23279_, new_n23280_, new_n23281_, new_n23282_, new_n23283_,
    new_n23284_, new_n23285_, new_n23286_, new_n23287_, new_n23288_,
    new_n23289_, new_n23290_, new_n23291_, new_n23292_, new_n23293_,
    new_n23294_, new_n23295_, new_n23296_, new_n23298_, new_n23299_,
    new_n23300_, new_n23301_, new_n23302_, new_n23303_, new_n23304_,
    new_n23305_, new_n23306_, new_n23307_, new_n23308_, new_n23309_,
    new_n23310_, new_n23311_, new_n23312_, new_n23313_, new_n23314_,
    new_n23315_, new_n23316_, new_n23317_, new_n23318_, new_n23319_,
    new_n23320_, new_n23321_, new_n23322_, new_n23323_, new_n23324_,
    new_n23325_, new_n23326_, new_n23327_, new_n23328_, new_n23329_,
    new_n23330_, new_n23331_, new_n23332_, new_n23333_, new_n23334_,
    new_n23335_, new_n23336_, new_n23337_, new_n23338_, new_n23339_,
    new_n23340_, new_n23341_, new_n23342_, new_n23343_, new_n23344_,
    new_n23345_, new_n23346_, new_n23347_, new_n23348_, new_n23349_,
    new_n23350_, new_n23351_, new_n23352_, new_n23353_, new_n23354_,
    new_n23355_, new_n23356_, new_n23357_, new_n23358_, new_n23359_,
    new_n23360_, new_n23361_, new_n23362_, new_n23363_, new_n23364_,
    new_n23365_, new_n23366_, new_n23367_, new_n23368_, new_n23369_,
    new_n23370_, new_n23371_, new_n23372_, new_n23373_, new_n23374_,
    new_n23375_, new_n23376_, new_n23377_, new_n23378_, new_n23379_,
    new_n23380_, new_n23381_, new_n23382_, new_n23383_, new_n23384_,
    new_n23385_, new_n23386_, new_n23387_, new_n23388_, new_n23389_,
    new_n23390_, new_n23391_, new_n23392_, new_n23393_, new_n23394_,
    new_n23395_, new_n23396_, new_n23397_, new_n23398_, new_n23399_,
    new_n23400_, new_n23401_, new_n23402_, new_n23403_, new_n23404_,
    new_n23405_, new_n23406_, new_n23407_, new_n23408_, new_n23409_,
    new_n23410_, new_n23411_, new_n23412_, new_n23413_, new_n23414_,
    new_n23415_, new_n23416_, new_n23417_, new_n23418_, new_n23419_,
    new_n23420_, new_n23421_, new_n23423_, new_n23424_, new_n23425_,
    new_n23426_, new_n23427_, new_n23428_, new_n23429_, new_n23430_,
    new_n23431_, new_n23432_, new_n23433_, new_n23434_, new_n23435_,
    new_n23436_, new_n23437_, new_n23438_, new_n23439_, new_n23440_,
    new_n23441_, new_n23442_, new_n23443_, new_n23444_, new_n23445_,
    new_n23446_, new_n23447_, new_n23448_, new_n23449_, new_n23450_,
    new_n23451_, new_n23452_, new_n23453_, new_n23454_, new_n23455_,
    new_n23456_, new_n23457_, new_n23458_, new_n23459_, new_n23460_,
    new_n23461_, new_n23462_, new_n23463_, new_n23464_, new_n23465_,
    new_n23466_, new_n23467_, new_n23468_, new_n23469_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23501_, new_n23502_, new_n23503_, new_n23504_, new_n23505_,
    new_n23506_, new_n23507_, new_n23508_, new_n23509_, new_n23510_,
    new_n23511_, new_n23512_, new_n23513_, new_n23514_, new_n23515_,
    new_n23516_, new_n23517_, new_n23518_, new_n23519_, new_n23520_,
    new_n23521_, new_n23522_, new_n23523_, new_n23524_, new_n23525_,
    new_n23526_, new_n23527_, new_n23528_, new_n23529_, new_n23530_,
    new_n23531_, new_n23532_, new_n23533_, new_n23534_, new_n23535_,
    new_n23536_, new_n23537_, new_n23538_, new_n23539_, new_n23540_,
    new_n23541_, new_n23542_, new_n23543_, new_n23544_, new_n23545_,
    new_n23547_, new_n23548_, new_n23549_, new_n23550_, new_n23551_,
    new_n23552_, new_n23553_, new_n23554_, new_n23555_, new_n23556_,
    new_n23557_, new_n23558_, new_n23559_, new_n23560_, new_n23561_,
    new_n23562_, new_n23563_, new_n23564_, new_n23565_, new_n23566_,
    new_n23567_, new_n23568_, new_n23569_, new_n23570_, new_n23571_,
    new_n23572_, new_n23573_, new_n23574_, new_n23575_, new_n23576_,
    new_n23577_, new_n23578_, new_n23579_, new_n23580_, new_n23581_,
    new_n23582_, new_n23583_, new_n23584_, new_n23585_, new_n23586_,
    new_n23587_, new_n23588_, new_n23589_, new_n23590_, new_n23591_,
    new_n23592_, new_n23593_, new_n23594_, new_n23595_, new_n23596_,
    new_n23597_, new_n23598_, new_n23599_, new_n23600_, new_n23601_,
    new_n23602_, new_n23603_, new_n23604_, new_n23605_, new_n23606_,
    new_n23607_, new_n23608_, new_n23609_, new_n23610_, new_n23611_,
    new_n23612_, new_n23613_, new_n23614_, new_n23615_, new_n23616_,
    new_n23617_, new_n23618_, new_n23619_, new_n23620_, new_n23621_,
    new_n23622_, new_n23623_, new_n23624_, new_n23625_, new_n23626_,
    new_n23627_, new_n23628_, new_n23629_, new_n23630_, new_n23631_,
    new_n23632_, new_n23633_, new_n23634_, new_n23635_, new_n23636_,
    new_n23637_, new_n23638_, new_n23639_, new_n23640_, new_n23641_,
    new_n23642_, new_n23643_, new_n23644_, new_n23645_, new_n23646_,
    new_n23647_, new_n23648_, new_n23649_, new_n23650_, new_n23651_,
    new_n23652_, new_n23653_, new_n23654_, new_n23655_, new_n23656_,
    new_n23657_, new_n23658_, new_n23659_, new_n23660_, new_n23661_,
    new_n23662_, new_n23663_, new_n23664_, new_n23665_, new_n23666_,
    new_n23667_, new_n23669_, new_n23670_, new_n23671_, new_n23672_,
    new_n23673_, new_n23674_, new_n23675_, new_n23676_, new_n23677_,
    new_n23678_, new_n23679_, new_n23680_, new_n23681_, new_n23682_,
    new_n23683_, new_n23684_, new_n23685_, new_n23686_, new_n23687_,
    new_n23688_, new_n23689_, new_n23690_, new_n23691_, new_n23692_,
    new_n23693_, new_n23694_, new_n23695_, new_n23696_, new_n23697_,
    new_n23698_, new_n23699_, new_n23700_, new_n23701_, new_n23702_,
    new_n23703_, new_n23704_, new_n23705_, new_n23706_, new_n23707_,
    new_n23708_, new_n23709_, new_n23710_, new_n23711_, new_n23712_,
    new_n23713_, new_n23714_, new_n23715_, new_n23716_, new_n23717_,
    new_n23718_, new_n23719_, new_n23720_, new_n23721_, new_n23722_,
    new_n23723_, new_n23724_, new_n23725_, new_n23726_, new_n23727_,
    new_n23728_, new_n23729_, new_n23730_, new_n23731_, new_n23732_,
    new_n23733_, new_n23734_, new_n23735_, new_n23736_, new_n23737_,
    new_n23738_, new_n23739_, new_n23740_, new_n23741_, new_n23742_,
    new_n23743_, new_n23744_, new_n23745_, new_n23746_, new_n23747_,
    new_n23748_, new_n23749_, new_n23750_, new_n23751_, new_n23752_,
    new_n23753_, new_n23754_, new_n23755_, new_n23756_, new_n23757_,
    new_n23758_, new_n23759_, new_n23760_, new_n23761_, new_n23762_,
    new_n23763_, new_n23764_, new_n23765_, new_n23766_, new_n23767_,
    new_n23768_, new_n23769_, new_n23770_, new_n23771_, new_n23772_,
    new_n23773_, new_n23774_, new_n23775_, new_n23776_, new_n23777_,
    new_n23778_, new_n23779_, new_n23780_, new_n23782_, new_n23783_,
    new_n23784_, new_n23785_, new_n23786_, new_n23787_, new_n23788_,
    new_n23789_, new_n23790_, new_n23791_, new_n23792_, new_n23793_,
    new_n23794_, new_n23795_, new_n23796_, new_n23797_, new_n23798_,
    new_n23799_, new_n23800_, new_n23801_, new_n23802_, new_n23803_,
    new_n23804_, new_n23805_, new_n23806_, new_n23807_, new_n23808_,
    new_n23809_, new_n23810_, new_n23811_, new_n23812_, new_n23813_,
    new_n23814_, new_n23815_, new_n23816_, new_n23817_, new_n23818_,
    new_n23819_, new_n23820_, new_n23821_, new_n23822_, new_n23823_,
    new_n23824_, new_n23825_, new_n23826_, new_n23827_, new_n23828_,
    new_n23829_, new_n23830_, new_n23831_, new_n23832_, new_n23833_,
    new_n23834_, new_n23835_, new_n23836_, new_n23837_, new_n23838_,
    new_n23839_, new_n23840_, new_n23841_, new_n23842_, new_n23843_,
    new_n23844_, new_n23845_, new_n23846_, new_n23847_, new_n23848_,
    new_n23849_, new_n23850_, new_n23851_, new_n23852_, new_n23853_,
    new_n23854_, new_n23855_, new_n23856_, new_n23857_, new_n23858_,
    new_n23859_, new_n23860_, new_n23861_, new_n23862_, new_n23863_,
    new_n23864_, new_n23865_, new_n23866_, new_n23867_, new_n23868_,
    new_n23869_, new_n23870_, new_n23871_, new_n23872_, new_n23873_,
    new_n23874_, new_n23875_, new_n23876_, new_n23877_, new_n23878_,
    new_n23879_, new_n23880_, new_n23881_, new_n23882_, new_n23883_,
    new_n23884_, new_n23885_, new_n23886_, new_n23887_, new_n23888_,
    new_n23889_, new_n23890_, new_n23891_, new_n23892_, new_n23893_,
    new_n23894_, new_n23896_, new_n23897_, new_n23898_, new_n23899_,
    new_n23900_, new_n23901_, new_n23902_, new_n23903_, new_n23904_,
    new_n23905_, new_n23906_, new_n23907_, new_n23908_, new_n23909_,
    new_n23910_, new_n23911_, new_n23912_, new_n23913_, new_n23914_,
    new_n23915_, new_n23916_, new_n23917_, new_n23918_, new_n23919_,
    new_n23920_, new_n23921_, new_n23922_, new_n23923_, new_n23924_,
    new_n23925_, new_n23926_, new_n23927_, new_n23928_, new_n23929_,
    new_n23930_, new_n23931_, new_n23932_, new_n23933_, new_n23934_,
    new_n23935_, new_n23936_, new_n23937_, new_n23938_, new_n23939_,
    new_n23940_, new_n23941_, new_n23942_, new_n23943_, new_n23944_,
    new_n23945_, new_n23946_, new_n23947_, new_n23948_, new_n23949_,
    new_n23950_, new_n23951_, new_n23952_, new_n23953_, new_n23954_,
    new_n23955_, new_n23956_, new_n23957_, new_n23958_, new_n23959_,
    new_n23960_, new_n23961_, new_n23962_, new_n23963_, new_n23964_,
    new_n23965_, new_n23966_, new_n23967_, new_n23968_, new_n23969_,
    new_n23970_, new_n23971_, new_n23972_, new_n23973_, new_n23974_,
    new_n23975_, new_n23976_, new_n23977_, new_n23978_, new_n23979_,
    new_n23980_, new_n23981_, new_n23982_, new_n23983_, new_n23984_,
    new_n23985_, new_n23986_, new_n23987_, new_n23988_, new_n23989_,
    new_n23990_, new_n23991_, new_n23992_, new_n23993_, new_n23995_,
    new_n23996_, new_n23997_, new_n23998_, new_n23999_, new_n24000_,
    new_n24001_, new_n24002_, new_n24003_, new_n24004_, new_n24005_,
    new_n24006_, new_n24007_, new_n24008_, new_n24009_, new_n24010_,
    new_n24011_, new_n24012_, new_n24013_, new_n24014_, new_n24015_,
    new_n24016_, new_n24017_, new_n24018_, new_n24019_, new_n24020_,
    new_n24021_, new_n24022_, new_n24023_, new_n24024_, new_n24025_,
    new_n24026_, new_n24027_, new_n24028_, new_n24029_, new_n24030_,
    new_n24031_, new_n24032_, new_n24033_, new_n24034_, new_n24035_,
    new_n24036_, new_n24037_, new_n24038_, new_n24039_, new_n24040_,
    new_n24041_, new_n24042_, new_n24043_, new_n24044_, new_n24045_,
    new_n24046_, new_n24047_, new_n24048_, new_n24049_, new_n24050_,
    new_n24051_, new_n24052_, new_n24053_, new_n24054_, new_n24055_,
    new_n24056_, new_n24057_, new_n24058_, new_n24059_, new_n24060_,
    new_n24061_, new_n24062_, new_n24063_, new_n24064_, new_n24065_,
    new_n24066_, new_n24067_, new_n24068_, new_n24069_, new_n24070_,
    new_n24071_, new_n24072_, new_n24073_, new_n24074_, new_n24075_,
    new_n24076_, new_n24077_, new_n24078_, new_n24079_, new_n24080_,
    new_n24081_, new_n24082_, new_n24083_, new_n24084_, new_n24085_,
    new_n24086_, new_n24087_, new_n24088_, new_n24089_, new_n24090_,
    new_n24091_, new_n24092_, new_n24093_, new_n24094_, new_n24095_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24193_, new_n24194_, new_n24195_, new_n24196_, new_n24197_,
    new_n24198_, new_n24199_, new_n24200_, new_n24201_, new_n24202_,
    new_n24203_, new_n24204_, new_n24205_, new_n24206_, new_n24207_,
    new_n24208_, new_n24209_, new_n24210_, new_n24211_, new_n24212_,
    new_n24213_, new_n24214_, new_n24215_, new_n24216_, new_n24217_,
    new_n24218_, new_n24219_, new_n24220_, new_n24221_, new_n24222_,
    new_n24223_, new_n24224_, new_n24225_, new_n24226_, new_n24227_,
    new_n24228_, new_n24229_, new_n24230_, new_n24231_, new_n24232_,
    new_n24233_, new_n24234_, new_n24235_, new_n24236_, new_n24237_,
    new_n24238_, new_n24239_, new_n24240_, new_n24241_, new_n24242_,
    new_n24243_, new_n24244_, new_n24245_, new_n24246_, new_n24247_,
    new_n24248_, new_n24249_, new_n24250_, new_n24251_, new_n24252_,
    new_n24253_, new_n24254_, new_n24255_, new_n24256_, new_n24257_,
    new_n24258_, new_n24259_, new_n24260_, new_n24261_, new_n24262_,
    new_n24263_, new_n24264_, new_n24265_, new_n24266_, new_n24267_,
    new_n24268_, new_n24269_, new_n24270_, new_n24271_, new_n24272_,
    new_n24273_, new_n24274_, new_n24275_, new_n24276_, new_n24277_,
    new_n24278_, new_n24279_, new_n24280_, new_n24281_, new_n24282_,
    new_n24283_, new_n24285_, new_n24286_, new_n24287_, new_n24288_,
    new_n24289_, new_n24290_, new_n24291_, new_n24292_, new_n24293_,
    new_n24294_, new_n24295_, new_n24296_, new_n24297_, new_n24298_,
    new_n24299_, new_n24300_, new_n24301_, new_n24302_, new_n24303_,
    new_n24304_, new_n24305_, new_n24306_, new_n24307_, new_n24308_,
    new_n24309_, new_n24310_, new_n24311_, new_n24312_, new_n24313_,
    new_n24314_, new_n24315_, new_n24316_, new_n24317_, new_n24318_,
    new_n24319_, new_n24320_, new_n24321_, new_n24322_, new_n24323_,
    new_n24324_, new_n24325_, new_n24326_, new_n24327_, new_n24328_,
    new_n24329_, new_n24330_, new_n24331_, new_n24332_, new_n24333_,
    new_n24334_, new_n24335_, new_n24336_, new_n24337_, new_n24338_,
    new_n24339_, new_n24340_, new_n24341_, new_n24342_, new_n24343_,
    new_n24344_, new_n24345_, new_n24346_, new_n24347_, new_n24348_,
    new_n24349_, new_n24350_, new_n24351_, new_n24352_, new_n24353_,
    new_n24354_, new_n24355_, new_n24356_, new_n24357_, new_n24358_,
    new_n24359_, new_n24360_, new_n24361_, new_n24362_, new_n24363_,
    new_n24364_, new_n24365_, new_n24366_, new_n24367_, new_n24369_,
    new_n24370_, new_n24371_, new_n24372_, new_n24373_, new_n24374_,
    new_n24375_, new_n24376_, new_n24377_, new_n24378_, new_n24379_,
    new_n24380_, new_n24381_, new_n24382_, new_n24383_, new_n24384_,
    new_n24385_, new_n24386_, new_n24387_, new_n24388_, new_n24389_,
    new_n24390_, new_n24391_, new_n24392_, new_n24393_, new_n24394_,
    new_n24395_, new_n24396_, new_n24397_, new_n24398_, new_n24399_,
    new_n24400_, new_n24401_, new_n24402_, new_n24403_, new_n24404_,
    new_n24405_, new_n24406_, new_n24407_, new_n24408_, new_n24409_,
    new_n24410_, new_n24411_, new_n24412_, new_n24413_, new_n24414_,
    new_n24415_, new_n24416_, new_n24417_, new_n24418_, new_n24419_,
    new_n24420_, new_n24421_, new_n24422_, new_n24423_, new_n24424_,
    new_n24425_, new_n24426_, new_n24427_, new_n24428_, new_n24429_,
    new_n24430_, new_n24431_, new_n24432_, new_n24433_, new_n24434_,
    new_n24435_, new_n24436_, new_n24437_, new_n24438_, new_n24439_,
    new_n24440_, new_n24441_, new_n24442_, new_n24443_, new_n24444_,
    new_n24446_, new_n24447_, new_n24448_, new_n24449_, new_n24450_,
    new_n24451_, new_n24452_, new_n24453_, new_n24454_, new_n24455_,
    new_n24456_, new_n24457_, new_n24458_, new_n24459_, new_n24460_,
    new_n24461_, new_n24462_, new_n24463_, new_n24464_, new_n24465_,
    new_n24466_, new_n24467_, new_n24468_, new_n24469_, new_n24470_,
    new_n24471_, new_n24472_, new_n24473_, new_n24474_, new_n24475_,
    new_n24476_, new_n24477_, new_n24478_, new_n24479_, new_n24480_,
    new_n24481_, new_n24482_, new_n24483_, new_n24484_, new_n24485_,
    new_n24486_, new_n24487_, new_n24488_, new_n24489_, new_n24490_,
    new_n24491_, new_n24492_, new_n24493_, new_n24494_, new_n24495_,
    new_n24496_, new_n24497_, new_n24498_, new_n24499_, new_n24500_,
    new_n24501_, new_n24502_, new_n24503_, new_n24504_, new_n24505_,
    new_n24506_, new_n24507_, new_n24508_, new_n24509_, new_n24510_,
    new_n24511_, new_n24512_, new_n24513_, new_n24514_, new_n24515_,
    new_n24516_, new_n24517_, new_n24518_, new_n24519_, new_n24521_,
    new_n24522_, new_n24523_, new_n24524_, new_n24525_, new_n24526_,
    new_n24527_, new_n24528_, new_n24529_, new_n24530_, new_n24531_,
    new_n24532_, new_n24533_, new_n24534_, new_n24535_, new_n24536_,
    new_n24537_, new_n24538_, new_n24539_, new_n24540_, new_n24541_,
    new_n24542_, new_n24543_, new_n24544_, new_n24545_, new_n24546_,
    new_n24547_, new_n24548_, new_n24549_, new_n24550_, new_n24551_,
    new_n24552_, new_n24553_, new_n24554_, new_n24555_, new_n24556_,
    new_n24557_, new_n24558_, new_n24559_, new_n24560_, new_n24561_,
    new_n24562_, new_n24563_, new_n24564_, new_n24565_, new_n24566_,
    new_n24567_, new_n24568_, new_n24569_, new_n24570_, new_n24571_,
    new_n24572_, new_n24573_, new_n24574_, new_n24575_, new_n24576_,
    new_n24577_, new_n24578_, new_n24579_, new_n24580_, new_n24581_,
    new_n24582_, new_n24583_, new_n24584_, new_n24585_, new_n24586_,
    new_n24587_, new_n24588_, new_n24589_, new_n24590_, new_n24591_,
    new_n24592_, new_n24594_, new_n24595_, new_n24596_, new_n24597_,
    new_n24598_, new_n24599_, new_n24600_, new_n24601_, new_n24602_,
    new_n24603_, new_n24604_, new_n24605_, new_n24606_, new_n24607_,
    new_n24608_, new_n24609_, new_n24610_, new_n24611_, new_n24612_,
    new_n24613_, new_n24614_, new_n24615_, new_n24616_, new_n24617_,
    new_n24618_, new_n24619_, new_n24620_, new_n24621_, new_n24622_,
    new_n24623_, new_n24624_, new_n24625_, new_n24626_, new_n24627_,
    new_n24628_, new_n24629_, new_n24630_, new_n24631_, new_n24632_,
    new_n24633_, new_n24634_, new_n24635_, new_n24636_, new_n24637_,
    new_n24638_, new_n24639_, new_n24640_, new_n24641_, new_n24642_,
    new_n24643_, new_n24644_, new_n24645_, new_n24646_, new_n24647_,
    new_n24648_, new_n24649_, new_n24650_, new_n24651_, new_n24652_,
    new_n24653_, new_n24654_, new_n24655_, new_n24656_, new_n24657_,
    new_n24658_, new_n24659_, new_n24660_, new_n24661_, new_n24662_,
    new_n24663_, new_n24665_, new_n24666_, new_n24667_, new_n24668_,
    new_n24669_, new_n24670_, new_n24671_, new_n24672_, new_n24673_,
    new_n24674_, new_n24675_, new_n24676_, new_n24677_, new_n24678_,
    new_n24679_, new_n24680_, new_n24681_, new_n24682_, new_n24683_,
    new_n24684_, new_n24685_, new_n24686_, new_n24687_, new_n24688_,
    new_n24689_, new_n24690_, new_n24691_, new_n24692_, new_n24693_,
    new_n24694_, new_n24695_, new_n24696_, new_n24697_, new_n24698_,
    new_n24699_, new_n24700_, new_n24701_, new_n24702_, new_n24703_,
    new_n24704_, new_n24705_, new_n24706_, new_n24707_, new_n24708_,
    new_n24709_, new_n24710_, new_n24711_, new_n24712_, new_n24713_,
    new_n24714_, new_n24715_, new_n24716_, new_n24717_, new_n24718_,
    new_n24719_, new_n24720_, new_n24721_, new_n24722_, new_n24723_,
    new_n24724_, new_n24725_, new_n24726_, new_n24727_, new_n24728_,
    new_n24729_, new_n24730_, new_n24731_, new_n24732_, new_n24734_,
    new_n24735_, new_n24736_, new_n24737_, new_n24738_, new_n24739_,
    new_n24740_, new_n24741_, new_n24742_, new_n24743_, new_n24744_,
    new_n24745_, new_n24746_, new_n24747_, new_n24748_, new_n24749_,
    new_n24750_, new_n24751_, new_n24752_, new_n24753_, new_n24754_,
    new_n24755_, new_n24756_, new_n24757_, new_n24758_, new_n24759_,
    new_n24760_, new_n24761_, new_n24762_, new_n24763_, new_n24764_,
    new_n24765_, new_n24766_, new_n24767_, new_n24768_, new_n24769_,
    new_n24770_, new_n24771_, new_n24772_, new_n24773_, new_n24774_,
    new_n24775_, new_n24776_, new_n24777_, new_n24778_, new_n24779_,
    new_n24780_, new_n24781_, new_n24782_, new_n24783_, new_n24784_,
    new_n24785_, new_n24786_, new_n24787_, new_n24788_, new_n24789_,
    new_n24790_, new_n24791_, new_n24792_, new_n24794_, new_n24795_,
    new_n24796_, new_n24797_, new_n24798_, new_n24799_, new_n24800_,
    new_n24801_, new_n24802_, new_n24803_, new_n24804_, new_n24805_,
    new_n24806_, new_n24807_, new_n24808_, new_n24809_, new_n24810_,
    new_n24811_, new_n24812_, new_n24813_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24820_,
    new_n24821_, new_n24822_, new_n24823_, new_n24824_, new_n24825_,
    new_n24826_, new_n24827_, new_n24828_, new_n24829_, new_n24830_,
    new_n24831_, new_n24832_, new_n24833_, new_n24834_, new_n24835_,
    new_n24836_, new_n24837_, new_n24838_, new_n24839_, new_n24840_,
    new_n24841_, new_n24842_, new_n24844_, new_n24845_, new_n24846_,
    new_n24847_, new_n24848_, new_n24849_, new_n24850_, new_n24851_,
    new_n24852_, new_n24853_, new_n24854_, new_n24855_, new_n24856_,
    new_n24857_, new_n24858_, new_n24859_, new_n24860_, new_n24861_,
    new_n24862_, new_n24863_, new_n24864_, new_n24865_, new_n24866_,
    new_n24867_, new_n24868_, new_n24869_, new_n24870_, new_n24871_,
    new_n24872_, new_n24873_, new_n24874_, new_n24875_, new_n24876_,
    new_n24877_, new_n24878_, new_n24879_, new_n24880_, new_n24881_,
    new_n24882_, new_n24883_, new_n24884_, new_n24885_, new_n24886_,
    new_n24887_, new_n24888_, new_n24889_, new_n24890_, new_n24891_,
    new_n24893_, new_n24894_, new_n24895_, new_n24896_, new_n24897_,
    new_n24898_, new_n24899_, new_n24900_, new_n24901_, new_n24902_,
    new_n24903_, new_n24904_, new_n24905_, new_n24906_, new_n24907_,
    new_n24908_, new_n24909_, new_n24910_, new_n24911_, new_n24912_,
    new_n24913_, new_n24914_, new_n24915_, new_n24916_, new_n24917_,
    new_n24918_, new_n24919_, new_n24920_, new_n24921_, new_n24922_,
    new_n24923_, new_n24924_, new_n24925_, new_n24926_, new_n24927_,
    new_n24928_, new_n24929_, new_n24930_, new_n24931_, new_n24932_,
    new_n24933_, new_n24934_, new_n24935_, new_n24936_, new_n24937_,
    new_n24938_, new_n24939_, new_n24940_, new_n24942_, new_n24943_,
    new_n24944_, new_n24945_, new_n24946_, new_n24947_, new_n24948_,
    new_n24949_, new_n24950_, new_n24951_, new_n24952_, new_n24953_,
    new_n24954_, new_n24955_, new_n24956_, new_n24957_, new_n24958_,
    new_n24959_, new_n24960_, new_n24961_, new_n24962_, new_n24963_,
    new_n24964_, new_n24965_, new_n24966_, new_n24967_, new_n24968_,
    new_n24969_, new_n24970_, new_n24971_, new_n24972_, new_n24973_,
    new_n24974_, new_n24975_, new_n24976_, new_n24977_, new_n24978_,
    new_n24979_, new_n24980_, new_n24981_, new_n24982_, new_n24984_,
    new_n24985_, new_n24986_, new_n24987_, new_n24988_, new_n24989_,
    new_n24990_, new_n24991_, new_n24992_, new_n24993_, new_n24994_,
    new_n24995_, new_n24996_, new_n24997_, new_n24998_, new_n24999_,
    new_n25000_, new_n25001_, new_n25002_, new_n25003_, new_n25004_,
    new_n25005_, new_n25006_, new_n25007_, new_n25008_, new_n25009_,
    new_n25010_, new_n25011_, new_n25012_, new_n25013_, new_n25014_,
    new_n25016_, new_n25017_, new_n25018_, new_n25019_, new_n25020_,
    new_n25021_, new_n25022_, new_n25023_, new_n25024_, new_n25025_,
    new_n25026_, new_n25027_, new_n25028_, new_n25029_, new_n25030_,
    new_n25031_, new_n25032_, new_n25033_, new_n25034_, new_n25035_,
    new_n25036_, new_n25037_, new_n25038_, new_n25039_, new_n25040_,
    new_n25041_, new_n25042_, new_n25043_, new_n25044_, new_n25045_,
    new_n25046_, new_n25047_, new_n25049_, new_n25050_, new_n25051_,
    new_n25052_, new_n25053_, new_n25054_, new_n25055_, new_n25056_,
    new_n25057_, new_n25058_, new_n25059_, new_n25060_, new_n25061_,
    new_n25062_, new_n25063_, new_n25064_, new_n25065_, new_n25066_,
    new_n25067_, new_n25068_, new_n25069_, new_n25070_, new_n25071_,
    new_n25072_, new_n25073_, new_n25074_, new_n25075_, new_n25076_,
    new_n25077_, new_n25078_, new_n25079_, new_n25081_, new_n25082_,
    new_n25083_, new_n25084_, new_n25085_, new_n25086_, new_n25087_,
    new_n25088_, new_n25089_, new_n25090_, new_n25091_, new_n25092_,
    new_n25093_, new_n25094_, new_n25095_, new_n25096_, new_n25097_,
    new_n25098_, new_n25099_, new_n25100_, new_n25101_, new_n25103_,
    new_n25104_, new_n25105_, new_n25106_, new_n25107_, new_n25108_,
    new_n25109_, new_n25110_, new_n25111_, new_n25112_, new_n25113_,
    new_n25114_, new_n25115_, new_n25116_, new_n25117_, new_n25118_,
    new_n25119_, new_n25120_, new_n25121_, new_n25122_, new_n25123_,
    new_n25124_, new_n25126_, new_n25127_, new_n25128_, new_n25129_,
    new_n25130_, new_n25131_, new_n25132_, new_n25133_, new_n25134_;
  INV_X1     g00000(.I(\a[0] ), .ZN(new_n257_));
  INV_X1     g00001(.I(\b[0] ), .ZN(new_n258_));
  NOR2_X1    g00002(.A1(new_n257_), .A2(new_n258_), .ZN(\f[0] ));
  INV_X1     g00003(.I(\a[2] ), .ZN(new_n260_));
  INV_X1     g00004(.I(\a[1] ), .ZN(new_n261_));
  NOR2_X1    g00005(.A1(new_n261_), .A2(\a[0] ), .ZN(new_n262_));
  INV_X1     g00006(.I(new_n262_), .ZN(new_n263_));
  XNOR2_X1   g00007(.A1(\a[0] ), .A2(\b[1] ), .ZN(new_n264_));
  NOR2_X1    g00008(.A1(new_n261_), .A2(new_n260_), .ZN(new_n265_));
  INV_X1     g00009(.I(new_n265_), .ZN(new_n266_));
  OAI22_X1   g00010(.A1(new_n264_), .A2(new_n266_), .B1(new_n263_), .B2(new_n258_), .ZN(new_n267_));
  NAND2_X1   g00011(.A1(\b[0] ), .A2(\b[1] ), .ZN(new_n268_));
  INV_X1     g00012(.I(\b[1] ), .ZN(new_n269_));
  NAND2_X1   g00013(.A1(new_n258_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1   g00014(.A1(new_n270_), .A2(new_n268_), .ZN(new_n271_));
  XNOR2_X1   g00015(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n272_));
  NOR2_X1    g00016(.A1(new_n272_), .A2(new_n257_), .ZN(new_n273_));
  NAND3_X1   g00017(.A1(new_n267_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  NOR3_X1    g00018(.A1(new_n274_), .A2(new_n260_), .A3(new_n258_), .ZN(new_n275_));
  XOR2_X1    g00019(.A1(new_n275_), .A2(\a[0] ), .Z(\f[1] ));
  NAND2_X1   g00020(.A1(new_n274_), .A2(new_n260_), .ZN(new_n277_));
  AND2_X2    g00021(.A1(new_n277_), .A2(\f[0] ), .Z(new_n278_));
  OAI21_X1   g00022(.A1(new_n269_), .A2(\b[0] ), .B(\b[2] ), .ZN(new_n279_));
  INV_X1     g00023(.I(\b[2] ), .ZN(new_n280_));
  NAND3_X1   g00024(.A1(new_n258_), .A2(new_n280_), .A3(\b[1] ), .ZN(new_n281_));
  NAND2_X1   g00025(.A1(new_n281_), .A2(new_n279_), .ZN(new_n282_));
  NAND2_X1   g00026(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1    g00027(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n284_));
  NOR2_X1    g00028(.A1(new_n265_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1    g00029(.A1(new_n285_), .A2(new_n257_), .ZN(new_n286_));
  AOI22_X1   g00030(.A1(new_n286_), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n262_), .ZN(new_n287_));
  NOR2_X1    g00031(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n288_));
  NAND2_X1   g00032(.A1(new_n288_), .A2(\a[2] ), .ZN(new_n289_));
  NOR4_X1    g00033(.A1(new_n287_), .A2(new_n260_), .A3(new_n258_), .A4(new_n289_), .ZN(new_n290_));
  XOR2_X1    g00034(.A1(new_n290_), .A2(new_n283_), .Z(new_n291_));
  XOR2_X1    g00035(.A1(new_n291_), .A2(new_n278_), .Z(\f[2] ));
  INV_X1     g00036(.I(new_n278_), .ZN(new_n293_));
  XNOR2_X1   g00037(.A1(\b[0] ), .A2(\b[2] ), .ZN(new_n294_));
  AOI21_X1   g00038(.A1(new_n269_), .A2(new_n280_), .B(\b[3] ), .ZN(new_n295_));
  NAND2_X1   g00039(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1    g00040(.A1(\b[0] ), .A2(\b[2] ), .Z(new_n297_));
  INV_X1     g00041(.I(\b[3] ), .ZN(new_n298_));
  OAI21_X1   g00042(.A1(\b[1] ), .A2(\b[2] ), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1   g00043(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1   g00044(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1    g00045(.A1(\a[0] ), .A2(\b[3] ), .Z(new_n302_));
  AOI22_X1   g00046(.A1(new_n302_), .A2(new_n265_), .B1(\b[2] ), .B2(new_n262_), .ZN(new_n303_));
  INV_X1     g00047(.I(new_n289_), .ZN(new_n304_));
  NAND2_X1   g00048(.A1(new_n304_), .A2(\b[1] ), .ZN(new_n305_));
  OAI21_X1   g00049(.A1(new_n303_), .A2(new_n305_), .B(new_n260_), .ZN(new_n306_));
  NAND2_X1   g00050(.A1(new_n306_), .A2(new_n301_), .ZN(new_n307_));
  XOR2_X1    g00051(.A1(new_n307_), .A2(new_n273_), .Z(new_n308_));
  XNOR2_X1   g00052(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n309_));
  NOR2_X1    g00053(.A1(new_n309_), .A2(new_n258_), .ZN(new_n310_));
  INV_X1     g00054(.I(new_n310_), .ZN(new_n311_));
  NOR2_X1    g00055(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1    g00056(.A1(new_n312_), .A2(new_n291_), .Z(new_n313_));
  XOR2_X1    g00057(.A1(new_n313_), .A2(new_n293_), .Z(\f[3] ));
  NOR3_X1    g00058(.A1(new_n269_), .A2(new_n298_), .A3(\b[0] ), .ZN(new_n315_));
  AOI21_X1   g00059(.A1(\b[1] ), .A2(\b[3] ), .B(new_n258_), .ZN(new_n316_));
  OAI21_X1   g00060(.A1(new_n316_), .A2(new_n315_), .B(\b[2] ), .ZN(new_n317_));
  NAND2_X1   g00061(.A1(new_n317_), .A2(new_n268_), .ZN(new_n318_));
  INV_X1     g00062(.I(new_n268_), .ZN(new_n319_));
  NAND3_X1   g00063(.A1(new_n258_), .A2(\b[1] ), .A3(\b[3] ), .ZN(new_n320_));
  OAI21_X1   g00064(.A1(new_n269_), .A2(new_n298_), .B(\b[0] ), .ZN(new_n321_));
  AOI21_X1   g00065(.A1(new_n321_), .A2(new_n320_), .B(new_n280_), .ZN(new_n322_));
  XOR2_X1    g00066(.A1(\b[3] ), .A2(\b[4] ), .Z(new_n323_));
  OAI21_X1   g00067(.A1(new_n322_), .A2(new_n319_), .B(new_n323_), .ZN(new_n324_));
  INV_X1     g00068(.I(\b[4] ), .ZN(new_n325_));
  NOR2_X1    g00069(.A1(new_n298_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1    g00070(.A1(\b[3] ), .A2(\b[4] ), .ZN(new_n327_));
  NOR2_X1    g00071(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1   g00072(.A1(new_n318_), .A2(new_n328_), .B(new_n324_), .ZN(new_n329_));
  INV_X1     g00073(.I(new_n286_), .ZN(new_n330_));
  AOI22_X1   g00074(.A1(new_n304_), .A2(\b[2] ), .B1(new_n262_), .B2(\b[4] ), .ZN(new_n331_));
  OAI21_X1   g00075(.A1(new_n330_), .A2(new_n298_), .B(new_n331_), .ZN(new_n332_));
  NAND3_X1   g00076(.A1(new_n329_), .A2(new_n332_), .A3(new_n273_), .ZN(new_n333_));
  INV_X1     g00077(.I(\a[5] ), .ZN(new_n334_));
  XNOR2_X1   g00078(.A1(\a[3] ), .A2(\a[5] ), .ZN(new_n335_));
  INV_X1     g00079(.I(\a[4] ), .ZN(new_n336_));
  NOR2_X1    g00080(.A1(new_n336_), .A2(\a[2] ), .ZN(new_n337_));
  NOR2_X1    g00081(.A1(new_n260_), .A2(\a[4] ), .ZN(new_n338_));
  NOR2_X1    g00082(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1    g00083(.A1(new_n339_), .A2(new_n335_), .ZN(new_n340_));
  INV_X1     g00084(.I(new_n340_), .ZN(new_n341_));
  NOR2_X1    g00085(.A1(new_n341_), .A2(new_n271_), .ZN(new_n342_));
  INV_X1     g00086(.I(\a[3] ), .ZN(new_n343_));
  NAND2_X1   g00087(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1   g00088(.A1(new_n338_), .A2(\a[3] ), .ZN(new_n345_));
  NAND2_X1   g00089(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI22_X1   g00090(.A1(\b[0] ), .A2(new_n340_), .B1(new_n346_), .B2(\b[1] ), .ZN(new_n347_));
  NOR2_X1    g00091(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1    g00092(.A1(new_n348_), .A2(new_n334_), .ZN(new_n349_));
  NOR3_X1    g00093(.A1(new_n342_), .A2(new_n347_), .A3(\a[5] ), .ZN(new_n350_));
  NOR2_X1    g00094(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1    g00095(.A1(new_n310_), .A2(new_n334_), .ZN(new_n352_));
  XOR2_X1    g00096(.A1(new_n351_), .A2(new_n352_), .Z(new_n353_));
  XOR2_X1    g00097(.A1(new_n353_), .A2(new_n333_), .Z(new_n354_));
  XOR2_X1    g00098(.A1(new_n354_), .A2(\a[2] ), .Z(new_n355_));
  NOR2_X1    g00099(.A1(new_n291_), .A2(new_n308_), .ZN(new_n356_));
  NAND2_X1   g00100(.A1(new_n291_), .A2(new_n308_), .ZN(new_n357_));
  NOR2_X1    g00101(.A1(new_n293_), .A2(new_n311_), .ZN(new_n358_));
  AOI21_X1   g00102(.A1(new_n357_), .A2(new_n358_), .B(new_n356_), .ZN(new_n359_));
  INV_X1     g00103(.I(new_n359_), .ZN(new_n360_));
  XOR2_X1    g00104(.A1(new_n355_), .A2(new_n360_), .Z(\f[4] ));
  XOR2_X1    g00105(.A1(new_n333_), .A2(\a[2] ), .Z(new_n362_));
  NOR2_X1    g00106(.A1(new_n353_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1   g00107(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n364_));
  NOR3_X1    g00108(.A1(new_n339_), .A2(new_n309_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1     g00109(.I(new_n365_), .ZN(new_n366_));
  AOI22_X1   g00110(.A1(\b[1] ), .A2(new_n340_), .B1(new_n346_), .B2(\b[2] ), .ZN(new_n367_));
  OAI21_X1   g00111(.A1(new_n258_), .A2(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND3_X1   g00112(.A1(new_n368_), .A2(new_n282_), .A3(new_n340_), .ZN(new_n369_));
  INV_X1     g00113(.I(new_n369_), .ZN(new_n370_));
  INV_X1     g00114(.I(new_n342_), .ZN(new_n371_));
  NOR4_X1    g00115(.A1(new_n371_), .A2(new_n334_), .A3(new_n311_), .A4(new_n347_), .ZN(new_n372_));
  XOR2_X1    g00116(.A1(\b[3] ), .A2(\b[5] ), .Z(new_n373_));
  NAND4_X1   g00117(.A1(new_n317_), .A2(new_n268_), .A3(new_n323_), .A4(new_n373_), .ZN(new_n374_));
  XNOR2_X1   g00118(.A1(\b[3] ), .A2(\b[4] ), .ZN(new_n375_));
  XNOR2_X1   g00119(.A1(\b[3] ), .A2(\b[5] ), .ZN(new_n376_));
  OAI22_X1   g00120(.A1(new_n322_), .A2(new_n319_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1   g00121(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NOR3_X1    g00122(.A1(new_n257_), .A2(new_n260_), .A3(\a[1] ), .ZN(new_n381_));
  XOR2_X1    g00123(.A1(new_n378_), .A2(new_n381_), .Z(new_n382_));
  XOR2_X1    g00124(.A1(new_n382_), .A2(new_n372_), .Z(new_n383_));
  XOR2_X1    g00125(.A1(new_n383_), .A2(new_n370_), .Z(new_n384_));
  XOR2_X1    g00126(.A1(new_n384_), .A2(\a[5] ), .Z(new_n385_));
  OAI21_X1   g00127(.A1(new_n385_), .A2(new_n363_), .B(new_n360_), .ZN(new_n386_));
  XNOR2_X1   g00128(.A1(new_n386_), .A2(new_n355_), .ZN(\f[5] ));
  XOR2_X1    g00129(.A1(new_n369_), .A2(new_n372_), .Z(new_n388_));
  XOR2_X1    g00130(.A1(new_n388_), .A2(new_n334_), .Z(new_n389_));
  NAND2_X1   g00131(.A1(new_n389_), .A2(new_n382_), .ZN(new_n390_));
  NAND2_X1   g00132(.A1(new_n385_), .A2(new_n363_), .ZN(new_n391_));
  NAND2_X1   g00133(.A1(new_n391_), .A2(new_n359_), .ZN(new_n392_));
  NAND2_X1   g00134(.A1(new_n392_), .A2(new_n355_), .ZN(new_n393_));
  INV_X1     g00135(.I(\a[6] ), .ZN(new_n394_));
  NOR2_X1    g00136(.A1(new_n334_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1    g00137(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n396_));
  NOR2_X1    g00138(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1     g00139(.I(new_n397_), .ZN(new_n398_));
  NOR2_X1    g00140(.A1(new_n398_), .A2(new_n258_), .ZN(new_n399_));
  XOR2_X1    g00141(.A1(new_n399_), .A2(new_n334_), .Z(new_n400_));
  NOR2_X1    g00142(.A1(new_n369_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1   g00143(.A1(new_n401_), .A2(new_n372_), .ZN(new_n402_));
  INV_X1     g00144(.I(new_n301_), .ZN(new_n403_));
  INV_X1     g00145(.I(new_n346_), .ZN(new_n404_));
  OAI22_X1   g00146(.A1(new_n280_), .A2(new_n341_), .B1(new_n404_), .B2(new_n298_), .ZN(new_n405_));
  OAI21_X1   g00147(.A1(new_n269_), .A2(new_n366_), .B(new_n405_), .ZN(new_n406_));
  AOI21_X1   g00148(.A1(new_n406_), .A2(new_n334_), .B(new_n341_), .ZN(new_n407_));
  XOR2_X1    g00149(.A1(new_n407_), .A2(new_n403_), .Z(new_n408_));
  XOR2_X1    g00150(.A1(new_n402_), .A2(new_n408_), .Z(new_n409_));
  NOR2_X1    g00151(.A1(new_n322_), .A2(new_n319_), .ZN(new_n410_));
  NOR2_X1    g00152(.A1(\b[4] ), .A2(\b[5] ), .ZN(new_n411_));
  AOI21_X1   g00153(.A1(new_n410_), .A2(new_n411_), .B(new_n298_), .ZN(new_n412_));
  NAND2_X1   g00154(.A1(\b[4] ), .A2(\b[5] ), .ZN(new_n413_));
  NOR2_X1    g00155(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1    g00156(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1   g00157(.A1(\b[5] ), .A2(\b[6] ), .ZN(new_n416_));
  NOR2_X1    g00158(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1     g00159(.I(new_n415_), .ZN(new_n418_));
  INV_X1     g00160(.I(\b[5] ), .ZN(new_n419_));
  INV_X1     g00161(.I(\b[6] ), .ZN(new_n420_));
  NOR2_X1    g00162(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1    g00163(.A1(\b[5] ), .A2(\b[6] ), .ZN(new_n422_));
  NOR2_X1    g00164(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1    g00165(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1    g00166(.A1(new_n424_), .A2(new_n417_), .ZN(new_n425_));
  INV_X1     g00167(.I(new_n273_), .ZN(new_n426_));
  OAI22_X1   g00168(.A1(new_n330_), .A2(new_n419_), .B1(new_n420_), .B2(new_n263_), .ZN(new_n427_));
  OAI21_X1   g00169(.A1(new_n325_), .A2(new_n289_), .B(new_n427_), .ZN(new_n428_));
  AOI21_X1   g00170(.A1(new_n428_), .A2(new_n260_), .B(new_n426_), .ZN(new_n429_));
  XOR2_X1    g00171(.A1(new_n425_), .A2(new_n429_), .Z(new_n430_));
  NOR2_X1    g00172(.A1(new_n409_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1    g00173(.A1(new_n393_), .A2(new_n431_), .Z(new_n432_));
  XOR2_X1    g00174(.A1(new_n432_), .A2(new_n390_), .Z(\f[6] ));
  NAND2_X1   g00175(.A1(new_n393_), .A2(new_n409_), .ZN(new_n434_));
  NOR2_X1    g00176(.A1(new_n390_), .A2(new_n430_), .ZN(new_n435_));
  NAND2_X1   g00177(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1   g00178(.A1(new_n393_), .A2(new_n409_), .B(new_n436_), .ZN(new_n437_));
  NOR2_X1    g00179(.A1(new_n370_), .A2(new_n334_), .ZN(new_n438_));
  NOR2_X1    g00180(.A1(new_n369_), .A2(\a[5] ), .ZN(new_n439_));
  OAI21_X1   g00181(.A1(new_n438_), .A2(new_n439_), .B(new_n372_), .ZN(new_n440_));
  NAND2_X1   g00182(.A1(new_n408_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1   g00183(.A1(new_n441_), .A2(\b[0] ), .A3(new_n398_), .ZN(new_n442_));
  OAI21_X1   g00184(.A1(new_n408_), .A2(new_n440_), .B(new_n442_), .ZN(new_n443_));
  INV_X1     g00185(.I(new_n271_), .ZN(new_n444_));
  XNOR2_X1   g00186(.A1(\a[6] ), .A2(\a[8] ), .ZN(new_n445_));
  XNOR2_X1   g00187(.A1(\a[5] ), .A2(\a[7] ), .ZN(new_n446_));
  NOR2_X1    g00188(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1     g00189(.I(new_n447_), .ZN(new_n448_));
  NOR3_X1    g00190(.A1(new_n334_), .A2(new_n394_), .A3(\a[7] ), .ZN(new_n449_));
  AOI21_X1   g00191(.A1(\a[7] ), .A2(new_n396_), .B(new_n449_), .ZN(new_n450_));
  INV_X1     g00192(.I(new_n450_), .ZN(new_n451_));
  INV_X1     g00193(.I(\a[8] ), .ZN(new_n452_));
  OAI21_X1   g00194(.A1(new_n448_), .A2(new_n258_), .B(new_n452_), .ZN(new_n453_));
  AOI21_X1   g00195(.A1(\b[1] ), .A2(new_n451_), .B(new_n453_), .ZN(new_n454_));
  NOR2_X1    g00196(.A1(new_n454_), .A2(new_n448_), .ZN(new_n455_));
  XOR2_X1    g00197(.A1(new_n455_), .A2(new_n444_), .Z(new_n456_));
  NOR2_X1    g00198(.A1(new_n399_), .A2(new_n452_), .ZN(new_n457_));
  NAND2_X1   g00199(.A1(new_n365_), .A2(\b[2] ), .ZN(new_n458_));
  AOI22_X1   g00200(.A1(\b[3] ), .A2(new_n340_), .B1(new_n346_), .B2(\b[4] ), .ZN(new_n459_));
  NAND2_X1   g00201(.A1(new_n459_), .A2(new_n458_), .ZN(new_n460_));
  NAND3_X1   g00202(.A1(new_n460_), .A2(new_n329_), .A3(new_n340_), .ZN(new_n461_));
  XOR2_X1    g00203(.A1(new_n461_), .A2(new_n457_), .Z(new_n462_));
  XOR2_X1    g00204(.A1(new_n456_), .A2(new_n462_), .Z(new_n463_));
  XOR2_X1    g00205(.A1(new_n463_), .A2(new_n334_), .Z(new_n464_));
  NOR2_X1    g00206(.A1(new_n464_), .A2(new_n443_), .ZN(new_n465_));
  AND2_X2    g00207(.A1(new_n464_), .A2(new_n443_), .Z(new_n466_));
  NOR2_X1    g00208(.A1(new_n466_), .A2(new_n465_), .ZN(new_n467_));
  INV_X1     g00209(.I(new_n467_), .ZN(new_n468_));
  XNOR2_X1   g00210(.A1(\b[5] ), .A2(\b[7] ), .ZN(new_n469_));
  NOR2_X1    g00211(.A1(new_n469_), .A2(new_n416_), .ZN(new_n470_));
  XOR2_X1    g00212(.A1(new_n415_), .A2(new_n470_), .Z(new_n471_));
  INV_X1     g00213(.I(\b[7] ), .ZN(new_n472_));
  OAI22_X1   g00214(.A1(new_n330_), .A2(new_n420_), .B1(new_n472_), .B2(new_n263_), .ZN(new_n473_));
  OAI21_X1   g00215(.A1(new_n419_), .A2(new_n289_), .B(new_n473_), .ZN(new_n474_));
  AOI21_X1   g00216(.A1(new_n474_), .A2(new_n260_), .B(new_n426_), .ZN(new_n475_));
  XOR2_X1    g00217(.A1(new_n471_), .A2(new_n475_), .Z(new_n476_));
  INV_X1     g00218(.I(new_n476_), .ZN(new_n477_));
  NAND2_X1   g00219(.A1(new_n468_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1   g00220(.A1(new_n467_), .A2(new_n476_), .ZN(new_n479_));
  NAND2_X1   g00221(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1    g00222(.A1(new_n467_), .A2(new_n476_), .Z(new_n481_));
  MUX2_X1    g00223(.I0(new_n481_), .I1(new_n480_), .S(new_n437_), .Z(\f[7] ));
  XOR2_X1    g00224(.A1(new_n461_), .A2(\a[5] ), .Z(new_n483_));
  XOR2_X1    g00225(.A1(new_n456_), .A2(new_n457_), .Z(new_n484_));
  NOR2_X1    g00226(.A1(new_n484_), .A2(new_n483_), .ZN(new_n485_));
  INV_X1     g00227(.I(new_n399_), .ZN(new_n486_));
  OAI21_X1   g00228(.A1(new_n464_), .A2(new_n486_), .B(new_n408_), .ZN(new_n487_));
  AOI21_X1   g00229(.A1(new_n464_), .A2(new_n486_), .B(new_n440_), .ZN(new_n488_));
  NAND2_X1   g00230(.A1(new_n488_), .A2(new_n487_), .ZN(new_n489_));
  AND2_X2    g00231(.A1(new_n281_), .A2(new_n279_), .Z(new_n490_));
  AOI21_X1   g00232(.A1(new_n269_), .A2(new_n490_), .B(new_n448_), .ZN(new_n491_));
  AOI21_X1   g00233(.A1(\b[2] ), .A2(new_n451_), .B(new_n491_), .ZN(new_n492_));
  INV_X1     g00234(.I(new_n446_), .ZN(new_n493_));
  XOR2_X1    g00235(.A1(\a[5] ), .A2(\a[6] ), .Z(new_n494_));
  XOR2_X1    g00236(.A1(\a[5] ), .A2(\a[8] ), .Z(new_n495_));
  NAND3_X1   g00237(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  NOR3_X1    g00238(.A1(new_n492_), .A2(new_n258_), .A3(new_n496_), .ZN(new_n497_));
  XOR2_X1    g00239(.A1(new_n497_), .A2(new_n452_), .Z(new_n498_));
  INV_X1     g00240(.I(new_n498_), .ZN(new_n499_));
  NAND2_X1   g00241(.A1(new_n456_), .A2(new_n457_), .ZN(new_n500_));
  OAI22_X1   g00242(.A1(new_n325_), .A2(new_n341_), .B1(new_n404_), .B2(new_n419_), .ZN(new_n501_));
  OAI21_X1   g00243(.A1(new_n298_), .A2(new_n366_), .B(new_n501_), .ZN(new_n502_));
  AOI21_X1   g00244(.A1(new_n340_), .A2(new_n378_), .B(new_n502_), .ZN(new_n503_));
  XOR2_X1    g00245(.A1(new_n500_), .A2(new_n503_), .Z(new_n504_));
  XOR2_X1    g00246(.A1(new_n504_), .A2(new_n499_), .Z(new_n505_));
  XOR2_X1    g00247(.A1(new_n505_), .A2(new_n334_), .Z(new_n506_));
  NOR2_X1    g00248(.A1(\b[6] ), .A2(\b[7] ), .ZN(new_n507_));
  AOI21_X1   g00249(.A1(new_n415_), .A2(new_n507_), .B(new_n419_), .ZN(new_n508_));
  NOR2_X1    g00250(.A1(new_n420_), .A2(new_n472_), .ZN(new_n509_));
  INV_X1     g00251(.I(new_n509_), .ZN(new_n510_));
  NOR2_X1    g00252(.A1(new_n415_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1   g00253(.A1(\b[7] ), .A2(\b[8] ), .ZN(new_n512_));
  INV_X1     g00254(.I(new_n512_), .ZN(new_n513_));
  OAI21_X1   g00255(.A1(new_n508_), .A2(new_n511_), .B(new_n513_), .ZN(new_n514_));
  INV_X1     g00256(.I(\b[8] ), .ZN(new_n515_));
  NOR2_X1    g00257(.A1(new_n472_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1     g00258(.I(new_n516_), .ZN(new_n517_));
  NAND2_X1   g00259(.A1(new_n472_), .A2(new_n515_), .ZN(new_n518_));
  AND2_X2    g00260(.A1(new_n517_), .A2(new_n518_), .Z(new_n519_));
  NOR3_X1    g00261(.A1(new_n508_), .A2(new_n511_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1     g00262(.I(new_n520_), .ZN(new_n521_));
  NAND2_X1   g00263(.A1(new_n521_), .A2(new_n514_), .ZN(new_n522_));
  OAI22_X1   g00264(.A1(new_n330_), .A2(new_n472_), .B1(new_n515_), .B2(new_n263_), .ZN(new_n523_));
  OAI21_X1   g00265(.A1(new_n420_), .A2(new_n289_), .B(new_n523_), .ZN(new_n524_));
  AOI21_X1   g00266(.A1(new_n524_), .A2(new_n260_), .B(new_n426_), .ZN(new_n525_));
  XOR2_X1    g00267(.A1(new_n522_), .A2(new_n525_), .Z(new_n526_));
  NAND2_X1   g00268(.A1(new_n506_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1   g00269(.A1(new_n527_), .A2(new_n489_), .ZN(new_n528_));
  XOR2_X1    g00270(.A1(new_n528_), .A2(new_n485_), .Z(new_n529_));
  INV_X1     g00271(.I(new_n529_), .ZN(new_n530_));
  NAND2_X1   g00272(.A1(new_n530_), .A2(new_n481_), .ZN(new_n531_));
  XOR2_X1    g00273(.A1(new_n531_), .A2(new_n478_), .Z(new_n532_));
  XOR2_X1    g00274(.A1(new_n532_), .A2(new_n437_), .Z(\f[8] ));
  XOR2_X1    g00275(.A1(new_n500_), .A2(new_n498_), .Z(new_n534_));
  NOR2_X1    g00276(.A1(new_n489_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X2    g00277(.A1(new_n489_), .A2(new_n534_), .Z(new_n536_));
  XOR2_X1    g00278(.A1(new_n503_), .A2(new_n334_), .Z(new_n537_));
  NOR4_X1    g00279(.A1(new_n536_), .A2(new_n483_), .A3(new_n484_), .A4(new_n537_), .ZN(new_n538_));
  NOR2_X1    g00280(.A1(new_n538_), .A2(new_n535_), .ZN(new_n539_));
  INV_X1     g00281(.I(new_n539_), .ZN(new_n540_));
  XOR2_X1    g00282(.A1(\a[8] ), .A2(\a[9] ), .Z(new_n541_));
  NAND2_X1   g00283(.A1(new_n541_), .A2(\b[0] ), .ZN(new_n542_));
  INV_X1     g00284(.I(new_n542_), .ZN(new_n543_));
  AOI22_X1   g00285(.A1(new_n451_), .A2(\b[3] ), .B1(\b[2] ), .B2(new_n447_), .ZN(new_n544_));
  NOR2_X1    g00286(.A1(new_n496_), .A2(new_n269_), .ZN(new_n545_));
  OAI21_X1   g00287(.A1(new_n544_), .A2(new_n545_), .B(new_n452_), .ZN(new_n546_));
  NAND2_X1   g00288(.A1(new_n546_), .A2(new_n447_), .ZN(new_n547_));
  NOR2_X1    g00289(.A1(new_n547_), .A2(new_n301_), .ZN(new_n548_));
  NAND2_X1   g00290(.A1(new_n547_), .A2(new_n301_), .ZN(new_n549_));
  INV_X1     g00291(.I(new_n549_), .ZN(new_n550_));
  NOR2_X1    g00292(.A1(new_n550_), .A2(new_n548_), .ZN(new_n551_));
  INV_X1     g00293(.I(new_n551_), .ZN(new_n552_));
  NOR2_X1    g00294(.A1(new_n499_), .A2(new_n500_), .ZN(new_n553_));
  INV_X1     g00295(.I(new_n417_), .ZN(new_n554_));
  OAI21_X1   g00296(.A1(new_n421_), .A2(new_n422_), .B(new_n415_), .ZN(new_n555_));
  NAND2_X1   g00297(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AOI22_X1   g00298(.A1(\b[5] ), .A2(new_n340_), .B1(new_n346_), .B2(\b[6] ), .ZN(new_n557_));
  AOI21_X1   g00299(.A1(\b[4] ), .A2(new_n365_), .B(new_n557_), .ZN(new_n558_));
  OAI21_X1   g00300(.A1(new_n558_), .A2(\a[5] ), .B(new_n340_), .ZN(new_n559_));
  XOR2_X1    g00301(.A1(new_n556_), .A2(new_n559_), .Z(new_n560_));
  XOR2_X1    g00302(.A1(new_n553_), .A2(new_n560_), .Z(new_n561_));
  XOR2_X1    g00303(.A1(new_n561_), .A2(new_n552_), .Z(new_n562_));
  XOR2_X1    g00304(.A1(new_n562_), .A2(new_n543_), .Z(new_n563_));
  NOR2_X1    g00305(.A1(new_n508_), .A2(new_n511_), .ZN(new_n564_));
  INV_X1     g00306(.I(\b[9] ), .ZN(new_n565_));
  NOR2_X1    g00307(.A1(new_n565_), .A2(\b[7] ), .ZN(new_n566_));
  NOR2_X1    g00308(.A1(new_n472_), .A2(\b[9] ), .ZN(new_n567_));
  OAI21_X1   g00309(.A1(new_n566_), .A2(new_n567_), .B(new_n513_), .ZN(new_n568_));
  XOR2_X1    g00310(.A1(new_n564_), .A2(new_n568_), .Z(new_n569_));
  NAND2_X1   g00311(.A1(new_n286_), .A2(\b[8] ), .ZN(new_n570_));
  AOI22_X1   g00312(.A1(new_n304_), .A2(\b[7] ), .B1(new_n262_), .B2(\b[9] ), .ZN(new_n571_));
  AOI21_X1   g00313(.A1(new_n570_), .A2(new_n571_), .B(new_n426_), .ZN(new_n572_));
  NAND2_X1   g00314(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1   g00315(.A1(new_n563_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1    g00316(.A1(new_n574_), .A2(new_n540_), .Z(new_n575_));
  XOR2_X1    g00317(.A1(new_n575_), .A2(\a[2] ), .Z(new_n576_));
  AOI21_X1   g00318(.A1(new_n530_), .A2(new_n468_), .B(new_n477_), .ZN(new_n577_));
  OAI21_X1   g00319(.A1(new_n530_), .A2(new_n468_), .B(new_n437_), .ZN(new_n578_));
  NOR2_X1    g00320(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1    g00321(.A1(new_n527_), .A2(new_n485_), .Z(new_n580_));
  NOR2_X1    g00322(.A1(new_n580_), .A2(new_n489_), .ZN(new_n581_));
  NOR2_X1    g00323(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1   g00324(.A1(new_n582_), .A2(new_n576_), .ZN(\f[9] ));
  XOR2_X1    g00325(.A1(new_n539_), .A2(\a[2] ), .Z(new_n584_));
  NOR3_X1    g00326(.A1(new_n576_), .A2(new_n574_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1   g00327(.A1(new_n585_), .A2(new_n581_), .B(new_n579_), .ZN(new_n586_));
  XOR2_X1    g00328(.A1(new_n551_), .A2(new_n542_), .Z(new_n587_));
  XOR2_X1    g00329(.A1(new_n551_), .A2(new_n542_), .Z(new_n588_));
  NOR2_X1    g00330(.A1(new_n588_), .A2(new_n553_), .ZN(new_n589_));
  AOI21_X1   g00331(.A1(new_n553_), .A2(new_n587_), .B(new_n589_), .ZN(new_n590_));
  INV_X1     g00332(.I(new_n590_), .ZN(new_n591_));
  NOR2_X1    g00333(.A1(new_n539_), .A2(new_n560_), .ZN(new_n592_));
  NOR2_X1    g00334(.A1(new_n498_), .A2(new_n551_), .ZN(new_n593_));
  NOR2_X1    g00335(.A1(new_n499_), .A2(new_n552_), .ZN(new_n594_));
  INV_X1     g00336(.I(new_n594_), .ZN(new_n595_));
  NOR2_X1    g00337(.A1(new_n500_), .A2(new_n542_), .ZN(new_n596_));
  AOI21_X1   g00338(.A1(new_n595_), .A2(new_n596_), .B(new_n593_), .ZN(new_n597_));
  OAI22_X1   g00339(.A1(new_n448_), .A2(new_n298_), .B1(new_n325_), .B2(new_n450_), .ZN(new_n598_));
  OAI21_X1   g00340(.A1(new_n280_), .A2(new_n496_), .B(new_n598_), .ZN(new_n599_));
  AOI21_X1   g00341(.A1(new_n329_), .A2(new_n447_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1   g00342(.A1(\a[9] ), .A2(\a[11] ), .ZN(new_n601_));
  INV_X1     g00343(.I(\a[10] ), .ZN(new_n602_));
  NOR2_X1    g00344(.A1(new_n602_), .A2(\a[8] ), .ZN(new_n603_));
  NOR2_X1    g00345(.A1(new_n452_), .A2(\a[10] ), .ZN(new_n604_));
  NOR2_X1    g00346(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1    g00347(.A1(new_n605_), .A2(new_n601_), .ZN(new_n606_));
  INV_X1     g00348(.I(new_n606_), .ZN(new_n607_));
  NOR3_X1    g00349(.A1(new_n602_), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n608_));
  AND2_X2    g00350(.A1(new_n604_), .A2(\a[9] ), .Z(new_n609_));
  NOR2_X1    g00351(.A1(new_n609_), .A2(new_n608_), .ZN(new_n610_));
  INV_X1     g00352(.I(new_n610_), .ZN(new_n611_));
  INV_X1     g00353(.I(\a[11] ), .ZN(new_n612_));
  OAI21_X1   g00354(.A1(new_n607_), .A2(new_n258_), .B(new_n612_), .ZN(new_n613_));
  AOI21_X1   g00355(.A1(\b[1] ), .A2(new_n611_), .B(new_n613_), .ZN(new_n614_));
  NOR3_X1    g00356(.A1(new_n614_), .A2(new_n271_), .A3(new_n607_), .ZN(new_n615_));
  NOR2_X1    g00357(.A1(new_n614_), .A2(new_n607_), .ZN(new_n616_));
  NOR2_X1    g00358(.A1(new_n616_), .A2(new_n444_), .ZN(new_n617_));
  NOR2_X1    g00359(.A1(new_n617_), .A2(new_n615_), .ZN(new_n618_));
  INV_X1     g00360(.I(new_n618_), .ZN(new_n619_));
  NOR2_X1    g00361(.A1(new_n543_), .A2(new_n612_), .ZN(new_n620_));
  NOR2_X1    g00362(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1     g00363(.I(new_n620_), .ZN(new_n622_));
  NOR2_X1    g00364(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1    g00365(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1     g00366(.I(new_n624_), .ZN(new_n625_));
  NOR2_X1    g00367(.A1(new_n625_), .A2(new_n452_), .ZN(new_n626_));
  NOR2_X1    g00368(.A1(new_n624_), .A2(\a[8] ), .ZN(new_n627_));
  OAI21_X1   g00369(.A1(new_n626_), .A2(new_n627_), .B(new_n600_), .ZN(new_n628_));
  NOR2_X1    g00370(.A1(new_n624_), .A2(new_n452_), .ZN(new_n629_));
  NOR2_X1    g00371(.A1(new_n625_), .A2(\a[8] ), .ZN(new_n630_));
  NOR2_X1    g00372(.A1(new_n630_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1   g00373(.A1(new_n600_), .A2(new_n631_), .B(new_n628_), .ZN(new_n632_));
  AOI22_X1   g00374(.A1(\b[6] ), .A2(new_n340_), .B1(new_n346_), .B2(\b[7] ), .ZN(new_n633_));
  AOI21_X1   g00375(.A1(\b[5] ), .A2(new_n365_), .B(new_n633_), .ZN(new_n634_));
  OAI21_X1   g00376(.A1(new_n634_), .A2(\a[5] ), .B(new_n340_), .ZN(new_n635_));
  XNOR2_X1   g00377(.A1(new_n471_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1    g00378(.A1(new_n632_), .A2(new_n636_), .Z(new_n637_));
  NOR2_X1    g00379(.A1(new_n637_), .A2(new_n597_), .ZN(new_n638_));
  INV_X1     g00380(.I(new_n597_), .ZN(new_n639_));
  INV_X1     g00381(.I(new_n636_), .ZN(new_n640_));
  XOR2_X1    g00382(.A1(new_n632_), .A2(new_n640_), .Z(new_n641_));
  NOR2_X1    g00383(.A1(new_n641_), .A2(new_n639_), .ZN(new_n642_));
  XOR2_X1    g00384(.A1(new_n539_), .A2(new_n560_), .Z(new_n643_));
  OAI21_X1   g00385(.A1(new_n638_), .A2(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XOR2_X1    g00386(.A1(new_n644_), .A2(new_n592_), .Z(new_n645_));
  XOR2_X1    g00387(.A1(new_n645_), .A2(new_n591_), .Z(new_n646_));
  NOR2_X1    g00388(.A1(\b[8] ), .A2(\b[9] ), .ZN(new_n647_));
  AOI21_X1   g00389(.A1(new_n564_), .A2(new_n647_), .B(new_n472_), .ZN(new_n648_));
  NOR2_X1    g00390(.A1(new_n515_), .A2(new_n565_), .ZN(new_n649_));
  INV_X1     g00391(.I(new_n649_), .ZN(new_n650_));
  NOR2_X1    g00392(.A1(new_n564_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1   g00393(.A1(\b[9] ), .A2(\b[10] ), .ZN(new_n652_));
  INV_X1     g00394(.I(new_n652_), .ZN(new_n653_));
  OAI21_X1   g00395(.A1(new_n648_), .A2(new_n651_), .B(new_n653_), .ZN(new_n654_));
  NOR2_X1    g00396(.A1(new_n648_), .A2(new_n651_), .ZN(new_n655_));
  INV_X1     g00397(.I(\b[10] ), .ZN(new_n656_));
  NOR2_X1    g00398(.A1(new_n565_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1    g00399(.A1(\b[9] ), .A2(\b[10] ), .ZN(new_n658_));
  OAI21_X1   g00400(.A1(new_n657_), .A2(new_n658_), .B(new_n655_), .ZN(new_n659_));
  NAND2_X1   g00401(.A1(new_n659_), .A2(new_n654_), .ZN(new_n660_));
  OAI22_X1   g00402(.A1(new_n330_), .A2(new_n565_), .B1(new_n656_), .B2(new_n263_), .ZN(new_n661_));
  OAI21_X1   g00403(.A1(new_n515_), .A2(new_n289_), .B(new_n661_), .ZN(new_n662_));
  AOI21_X1   g00404(.A1(new_n662_), .A2(new_n260_), .B(new_n426_), .ZN(new_n663_));
  XNOR2_X1   g00405(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  XOR2_X1    g00406(.A1(new_n646_), .A2(new_n664_), .Z(new_n665_));
  XOR2_X1    g00407(.A1(new_n646_), .A2(new_n664_), .Z(new_n666_));
  NAND2_X1   g00408(.A1(new_n666_), .A2(new_n586_), .ZN(new_n667_));
  OAI21_X1   g00409(.A1(new_n586_), .A2(new_n665_), .B(new_n667_), .ZN(\f[10] ));
  NOR2_X1    g00410(.A1(new_n646_), .A2(new_n664_), .ZN(new_n669_));
  XOR2_X1    g00411(.A1(new_n632_), .A2(new_n639_), .Z(new_n670_));
  NOR2_X1    g00412(.A1(new_n670_), .A2(new_n640_), .ZN(new_n671_));
  NOR2_X1    g00413(.A1(new_n638_), .A2(new_n642_), .ZN(new_n672_));
  OAI21_X1   g00414(.A1(new_n672_), .A2(new_n560_), .B(new_n539_), .ZN(new_n673_));
  AOI21_X1   g00415(.A1(new_n672_), .A2(new_n560_), .B(new_n590_), .ZN(new_n674_));
  NAND2_X1   g00416(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1     g00417(.I(new_n675_), .ZN(new_n676_));
  XOR2_X1    g00418(.A1(new_n600_), .A2(new_n452_), .Z(new_n677_));
  INV_X1     g00419(.I(new_n677_), .ZN(new_n678_));
  NAND2_X1   g00420(.A1(new_n625_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1   g00421(.A1(new_n269_), .A2(new_n490_), .B(new_n607_), .ZN(new_n680_));
  AOI21_X1   g00422(.A1(\b[2] ), .A2(new_n611_), .B(new_n680_), .ZN(new_n681_));
  INV_X1     g00423(.I(new_n605_), .ZN(new_n682_));
  XOR2_X1    g00424(.A1(\a[8] ), .A2(\a[11] ), .Z(new_n683_));
  NAND3_X1   g00425(.A1(new_n682_), .A2(new_n541_), .A3(new_n683_), .ZN(new_n684_));
  NOR3_X1    g00426(.A1(new_n681_), .A2(new_n258_), .A3(new_n684_), .ZN(new_n685_));
  XOR2_X1    g00427(.A1(new_n685_), .A2(new_n612_), .Z(new_n686_));
  INV_X1     g00428(.I(new_n686_), .ZN(new_n687_));
  NAND2_X1   g00429(.A1(new_n618_), .A2(new_n620_), .ZN(new_n688_));
  OAI22_X1   g00430(.A1(new_n448_), .A2(new_n325_), .B1(new_n419_), .B2(new_n450_), .ZN(new_n689_));
  OAI21_X1   g00431(.A1(new_n298_), .A2(new_n496_), .B(new_n689_), .ZN(new_n690_));
  AOI21_X1   g00432(.A1(new_n378_), .A2(new_n447_), .B(new_n690_), .ZN(new_n691_));
  XOR2_X1    g00433(.A1(new_n688_), .A2(new_n691_), .Z(new_n692_));
  XOR2_X1    g00434(.A1(new_n692_), .A2(new_n687_), .Z(new_n693_));
  XOR2_X1    g00435(.A1(new_n693_), .A2(new_n452_), .Z(new_n694_));
  XOR2_X1    g00436(.A1(new_n624_), .A2(new_n677_), .Z(new_n695_));
  NAND2_X1   g00437(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  XOR2_X1    g00438(.A1(new_n696_), .A2(new_n679_), .Z(new_n697_));
  XOR2_X1    g00439(.A1(new_n697_), .A2(new_n597_), .Z(new_n698_));
  INV_X1     g00440(.I(new_n514_), .ZN(new_n699_));
  NOR2_X1    g00441(.A1(new_n699_), .A2(new_n520_), .ZN(new_n700_));
  OAI22_X1   g00442(.A1(new_n472_), .A2(new_n341_), .B1(new_n404_), .B2(new_n515_), .ZN(new_n701_));
  OAI21_X1   g00443(.A1(new_n420_), .A2(new_n366_), .B(new_n701_), .ZN(new_n702_));
  AOI21_X1   g00444(.A1(new_n702_), .A2(new_n334_), .B(new_n341_), .ZN(new_n703_));
  XOR2_X1    g00445(.A1(new_n700_), .A2(new_n703_), .Z(new_n704_));
  XOR2_X1    g00446(.A1(new_n698_), .A2(new_n704_), .Z(new_n705_));
  INV_X1     g00447(.I(\b[11] ), .ZN(new_n706_));
  NOR2_X1    g00448(.A1(new_n706_), .A2(\b[9] ), .ZN(new_n707_));
  NOR2_X1    g00449(.A1(new_n565_), .A2(\b[11] ), .ZN(new_n708_));
  OAI21_X1   g00450(.A1(new_n707_), .A2(new_n708_), .B(new_n653_), .ZN(new_n709_));
  XOR2_X1    g00451(.A1(new_n655_), .A2(new_n709_), .Z(new_n710_));
  OAI22_X1   g00452(.A1(new_n330_), .A2(new_n656_), .B1(new_n706_), .B2(new_n263_), .ZN(new_n711_));
  OAI21_X1   g00453(.A1(new_n565_), .A2(new_n289_), .B(new_n711_), .ZN(new_n712_));
  AOI21_X1   g00454(.A1(new_n712_), .A2(new_n260_), .B(new_n426_), .ZN(new_n713_));
  XOR2_X1    g00455(.A1(new_n710_), .A2(new_n713_), .Z(new_n714_));
  NAND2_X1   g00456(.A1(new_n705_), .A2(new_n714_), .ZN(new_n715_));
  XOR2_X1    g00457(.A1(new_n715_), .A2(new_n676_), .Z(new_n716_));
  XOR2_X1    g00458(.A1(new_n716_), .A2(new_n671_), .Z(new_n717_));
  INV_X1     g00459(.I(new_n717_), .ZN(new_n718_));
  NAND2_X1   g00460(.A1(new_n718_), .A2(new_n666_), .ZN(new_n719_));
  XOR2_X1    g00461(.A1(new_n719_), .A2(new_n669_), .Z(new_n720_));
  XOR2_X1    g00462(.A1(new_n720_), .A2(new_n586_), .Z(\f[11] ));
  INV_X1     g00463(.I(new_n671_), .ZN(new_n722_));
  XOR2_X1    g00464(.A1(new_n715_), .A2(new_n722_), .Z(new_n723_));
  NAND2_X1   g00465(.A1(new_n723_), .A2(new_n676_), .ZN(new_n724_));
  OAI21_X1   g00466(.A1(new_n717_), .A2(new_n646_), .B(new_n664_), .ZN(new_n725_));
  AOI21_X1   g00467(.A1(new_n717_), .A2(new_n646_), .B(new_n586_), .ZN(new_n726_));
  NAND2_X1   g00468(.A1(new_n726_), .A2(new_n725_), .ZN(new_n727_));
  AND2_X2    g00469(.A1(new_n698_), .A2(new_n722_), .Z(new_n728_));
  OR3_X2     g00470(.A1(new_n728_), .A2(new_n675_), .A3(new_n704_), .Z(new_n729_));
  OAI21_X1   g00471(.A1(new_n722_), .A2(new_n698_), .B(new_n729_), .ZN(new_n730_));
  XOR2_X1    g00472(.A1(new_n691_), .A2(new_n452_), .Z(new_n731_));
  XNOR2_X1   g00473(.A1(new_n686_), .A2(new_n688_), .ZN(new_n732_));
  NOR2_X1    g00474(.A1(new_n732_), .A2(new_n731_), .ZN(new_n733_));
  INV_X1     g00475(.I(new_n733_), .ZN(new_n734_));
  AOI21_X1   g00476(.A1(new_n694_), .A2(new_n625_), .B(new_n678_), .ZN(new_n735_));
  OAI21_X1   g00477(.A1(new_n694_), .A2(new_n625_), .B(new_n639_), .ZN(new_n736_));
  NOR2_X1    g00478(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1     g00479(.I(new_n688_), .ZN(new_n738_));
  INV_X1     g00480(.I(new_n684_), .ZN(new_n739_));
  OAI22_X1   g00481(.A1(new_n607_), .A2(new_n280_), .B1(new_n610_), .B2(new_n298_), .ZN(new_n740_));
  AOI21_X1   g00482(.A1(\b[1] ), .A2(new_n739_), .B(new_n740_), .ZN(new_n741_));
  NOR3_X1    g00483(.A1(new_n741_), .A2(new_n403_), .A3(new_n607_), .ZN(new_n742_));
  XOR2_X1    g00484(.A1(new_n742_), .A2(new_n612_), .Z(new_n743_));
  XOR2_X1    g00485(.A1(\a[11] ), .A2(\a[12] ), .Z(new_n744_));
  NAND2_X1   g00486(.A1(new_n744_), .A2(\b[0] ), .ZN(new_n745_));
  NOR2_X1    g00487(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  XOR2_X1    g00488(.A1(new_n746_), .A2(new_n686_), .Z(new_n747_));
  XOR2_X1    g00489(.A1(new_n747_), .A2(new_n738_), .Z(new_n748_));
  INV_X1     g00490(.I(new_n496_), .ZN(new_n749_));
  AOI22_X1   g00491(.A1(new_n451_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n447_), .ZN(new_n750_));
  AOI21_X1   g00492(.A1(\b[4] ), .A2(new_n749_), .B(new_n750_), .ZN(new_n751_));
  OAI21_X1   g00493(.A1(new_n751_), .A2(\a[8] ), .B(new_n447_), .ZN(new_n752_));
  XOR2_X1    g00494(.A1(new_n556_), .A2(new_n752_), .Z(new_n753_));
  NOR2_X1    g00495(.A1(new_n748_), .A2(new_n753_), .ZN(new_n754_));
  XOR2_X1    g00496(.A1(new_n737_), .A2(new_n754_), .Z(new_n755_));
  NAND2_X1   g00497(.A1(new_n755_), .A2(new_n734_), .ZN(new_n756_));
  OR2_X2     g00498(.A1(new_n755_), .A2(new_n734_), .Z(new_n757_));
  NAND2_X1   g00499(.A1(new_n757_), .A2(new_n756_), .ZN(new_n758_));
  XNOR2_X1   g00500(.A1(new_n564_), .A2(new_n568_), .ZN(new_n759_));
  OAI22_X1   g00501(.A1(new_n515_), .A2(new_n341_), .B1(new_n404_), .B2(new_n565_), .ZN(new_n760_));
  OAI21_X1   g00502(.A1(new_n472_), .A2(new_n366_), .B(new_n760_), .ZN(new_n761_));
  AOI21_X1   g00503(.A1(new_n761_), .A2(new_n334_), .B(new_n341_), .ZN(new_n762_));
  XOR2_X1    g00504(.A1(new_n759_), .A2(new_n762_), .Z(new_n763_));
  XOR2_X1    g00505(.A1(new_n758_), .A2(new_n763_), .Z(new_n764_));
  NOR2_X1    g00506(.A1(new_n758_), .A2(new_n763_), .ZN(new_n765_));
  INV_X1     g00507(.I(new_n765_), .ZN(new_n766_));
  NAND2_X1   g00508(.A1(new_n758_), .A2(new_n763_), .ZN(new_n767_));
  AOI21_X1   g00509(.A1(new_n766_), .A2(new_n767_), .B(new_n730_), .ZN(new_n768_));
  AOI21_X1   g00510(.A1(new_n730_), .A2(new_n764_), .B(new_n768_), .ZN(new_n769_));
  NOR2_X1    g00511(.A1(\b[10] ), .A2(\b[11] ), .ZN(new_n770_));
  AOI21_X1   g00512(.A1(new_n655_), .A2(new_n770_), .B(new_n565_), .ZN(new_n771_));
  NOR2_X1    g00513(.A1(new_n656_), .A2(new_n706_), .ZN(new_n772_));
  INV_X1     g00514(.I(new_n772_), .ZN(new_n773_));
  NOR2_X1    g00515(.A1(new_n655_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1    g00516(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  XNOR2_X1   g00517(.A1(\b[11] ), .A2(\b[12] ), .ZN(new_n776_));
  NOR2_X1    g00518(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NOR4_X1    g00519(.A1(new_n648_), .A2(new_n651_), .A3(\b[10] ), .A4(\b[11] ), .ZN(new_n778_));
  OAI22_X1   g00520(.A1(new_n778_), .A2(new_n565_), .B1(new_n655_), .B2(new_n773_), .ZN(new_n779_));
  INV_X1     g00521(.I(\b[12] ), .ZN(new_n780_));
  NOR2_X1    g00522(.A1(new_n706_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1    g00523(.A1(\b[11] ), .A2(\b[12] ), .ZN(new_n782_));
  NOR2_X1    g00524(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1    g00525(.A1(new_n779_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1    g00526(.A1(new_n777_), .A2(new_n784_), .ZN(new_n785_));
  OAI22_X1   g00527(.A1(new_n330_), .A2(new_n706_), .B1(new_n780_), .B2(new_n263_), .ZN(new_n786_));
  OAI21_X1   g00528(.A1(new_n656_), .A2(new_n289_), .B(new_n786_), .ZN(new_n787_));
  AOI21_X1   g00529(.A1(new_n787_), .A2(new_n260_), .B(new_n426_), .ZN(new_n788_));
  XOR2_X1    g00530(.A1(new_n785_), .A2(new_n788_), .Z(new_n789_));
  NOR2_X1    g00531(.A1(new_n769_), .A2(new_n789_), .ZN(new_n790_));
  XOR2_X1    g00532(.A1(new_n727_), .A2(new_n790_), .Z(new_n791_));
  XOR2_X1    g00533(.A1(new_n791_), .A2(new_n724_), .Z(\f[12] ));
  NOR2_X1    g00534(.A1(new_n727_), .A2(new_n769_), .ZN(new_n793_));
  OR2_X2     g00535(.A1(new_n724_), .A2(new_n789_), .Z(new_n794_));
  AOI21_X1   g00536(.A1(new_n727_), .A2(new_n769_), .B(new_n794_), .ZN(new_n795_));
  NOR2_X1    g00537(.A1(new_n795_), .A2(new_n793_), .ZN(new_n796_));
  INV_X1     g00538(.I(new_n796_), .ZN(new_n797_));
  NAND2_X1   g00539(.A1(new_n730_), .A2(new_n767_), .ZN(new_n798_));
  INV_X1     g00540(.I(new_n798_), .ZN(new_n799_));
  OR2_X2     g00541(.A1(new_n686_), .A2(new_n743_), .Z(new_n800_));
  INV_X1     g00542(.I(new_n745_), .ZN(new_n801_));
  NAND2_X1   g00543(.A1(new_n686_), .A2(new_n743_), .ZN(new_n802_));
  NAND3_X1   g00544(.A1(new_n802_), .A2(new_n738_), .A3(new_n801_), .ZN(new_n803_));
  NAND2_X1   g00545(.A1(new_n803_), .A2(new_n800_), .ZN(new_n804_));
  INV_X1     g00546(.I(new_n804_), .ZN(new_n805_));
  NOR3_X1    g00547(.A1(new_n322_), .A2(new_n319_), .A3(new_n328_), .ZN(new_n806_));
  AOI21_X1   g00548(.A1(new_n318_), .A2(new_n323_), .B(new_n806_), .ZN(new_n807_));
  OAI22_X1   g00549(.A1(new_n607_), .A2(new_n298_), .B1(new_n610_), .B2(new_n325_), .ZN(new_n808_));
  OAI21_X1   g00550(.A1(new_n280_), .A2(new_n684_), .B(new_n808_), .ZN(new_n809_));
  AOI21_X1   g00551(.A1(new_n809_), .A2(new_n612_), .B(new_n607_), .ZN(new_n810_));
  XOR2_X1    g00552(.A1(new_n810_), .A2(new_n807_), .Z(new_n811_));
  XNOR2_X1   g00553(.A1(\a[12] ), .A2(\a[14] ), .ZN(new_n812_));
  INV_X1     g00554(.I(\a[13] ), .ZN(new_n813_));
  NOR2_X1    g00555(.A1(new_n813_), .A2(\a[11] ), .ZN(new_n814_));
  NOR2_X1    g00556(.A1(new_n612_), .A2(\a[13] ), .ZN(new_n815_));
  NOR2_X1    g00557(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1    g00558(.A1(new_n816_), .A2(new_n812_), .ZN(new_n817_));
  NOR3_X1    g00559(.A1(new_n813_), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n818_));
  AND3_X2    g00560(.A1(new_n813_), .A2(\a[11] ), .A3(\a[12] ), .Z(new_n819_));
  NOR2_X1    g00561(.A1(new_n819_), .A2(new_n818_), .ZN(new_n820_));
  AOI21_X1   g00562(.A1(new_n817_), .A2(\b[0] ), .B(\a[14] ), .ZN(new_n821_));
  OAI21_X1   g00563(.A1(new_n269_), .A2(new_n820_), .B(new_n821_), .ZN(new_n822_));
  NAND2_X1   g00564(.A1(new_n822_), .A2(new_n817_), .ZN(new_n823_));
  NOR2_X1    g00565(.A1(new_n823_), .A2(new_n271_), .ZN(new_n824_));
  AOI21_X1   g00566(.A1(new_n822_), .A2(new_n817_), .B(new_n444_), .ZN(new_n825_));
  NOR2_X1    g00567(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1     g00568(.I(\a[14] ), .ZN(new_n827_));
  NOR2_X1    g00569(.A1(new_n801_), .A2(new_n827_), .ZN(new_n828_));
  XOR2_X1    g00570(.A1(new_n826_), .A2(new_n828_), .Z(new_n829_));
  XNOR2_X1   g00571(.A1(new_n829_), .A2(new_n811_), .ZN(new_n830_));
  NAND2_X1   g00572(.A1(new_n829_), .A2(new_n811_), .ZN(new_n831_));
  NOR2_X1    g00573(.A1(new_n829_), .A2(new_n811_), .ZN(new_n832_));
  INV_X1     g00574(.I(new_n832_), .ZN(new_n833_));
  NAND2_X1   g00575(.A1(new_n833_), .A2(new_n831_), .ZN(new_n834_));
  NAND2_X1   g00576(.A1(new_n805_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1   g00577(.A1(new_n805_), .A2(new_n830_), .B(new_n835_), .ZN(new_n836_));
  AOI22_X1   g00578(.A1(new_n451_), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n447_), .ZN(new_n837_));
  AOI21_X1   g00579(.A1(\b[5] ), .A2(new_n749_), .B(new_n837_), .ZN(new_n838_));
  OAI21_X1   g00580(.A1(new_n838_), .A2(\a[8] ), .B(new_n447_), .ZN(new_n839_));
  XNOR2_X1   g00581(.A1(new_n471_), .A2(new_n839_), .ZN(new_n840_));
  XOR2_X1    g00582(.A1(new_n836_), .A2(new_n840_), .Z(new_n841_));
  AOI21_X1   g00583(.A1(new_n748_), .A2(new_n734_), .B(new_n753_), .ZN(new_n842_));
  NAND2_X1   g00584(.A1(new_n737_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1   g00585(.A1(new_n734_), .A2(new_n748_), .B(new_n843_), .ZN(new_n844_));
  XOR2_X1    g00586(.A1(new_n844_), .A2(new_n841_), .Z(new_n845_));
  INV_X1     g00587(.I(new_n845_), .ZN(new_n846_));
  OAI22_X1   g00588(.A1(new_n565_), .A2(new_n341_), .B1(new_n404_), .B2(new_n656_), .ZN(new_n847_));
  OAI21_X1   g00589(.A1(new_n515_), .A2(new_n366_), .B(new_n847_), .ZN(new_n848_));
  AOI21_X1   g00590(.A1(new_n848_), .A2(new_n334_), .B(new_n341_), .ZN(new_n849_));
  XNOR2_X1   g00591(.A1(new_n660_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1    g00592(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1   g00593(.A1(new_n846_), .A2(new_n850_), .ZN(new_n852_));
  INV_X1     g00594(.I(new_n852_), .ZN(new_n853_));
  OAI22_X1   g00595(.A1(new_n799_), .A2(new_n765_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  XNOR2_X1   g00596(.A1(new_n845_), .A2(new_n850_), .ZN(new_n855_));
  NAND3_X1   g00597(.A1(new_n798_), .A2(new_n766_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1   g00598(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  XNOR2_X1   g00599(.A1(\b[11] ), .A2(\b[13] ), .ZN(new_n858_));
  NOR2_X1    g00600(.A1(new_n858_), .A2(new_n776_), .ZN(new_n859_));
  XOR2_X1    g00601(.A1(new_n779_), .A2(new_n859_), .Z(new_n860_));
  INV_X1     g00602(.I(\b[13] ), .ZN(new_n861_));
  OAI22_X1   g00603(.A1(new_n330_), .A2(new_n780_), .B1(new_n861_), .B2(new_n263_), .ZN(new_n862_));
  OAI21_X1   g00604(.A1(new_n706_), .A2(new_n289_), .B(new_n862_), .ZN(new_n863_));
  AOI21_X1   g00605(.A1(new_n863_), .A2(new_n260_), .B(new_n426_), .ZN(new_n864_));
  XNOR2_X1   g00606(.A1(new_n860_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1     g00607(.I(new_n865_), .ZN(new_n866_));
  XOR2_X1    g00608(.A1(new_n857_), .A2(new_n866_), .Z(new_n867_));
  NAND2_X1   g00609(.A1(new_n797_), .A2(new_n867_), .ZN(new_n868_));
  XOR2_X1    g00610(.A1(new_n857_), .A2(new_n866_), .Z(new_n869_));
  OAI21_X1   g00611(.A1(new_n797_), .A2(new_n869_), .B(new_n868_), .ZN(\f[13] ));
  NAND2_X1   g00612(.A1(new_n857_), .A2(new_n866_), .ZN(new_n871_));
  INV_X1     g00613(.I(new_n841_), .ZN(new_n872_));
  XNOR2_X1   g00614(.A1(new_n844_), .A2(new_n850_), .ZN(new_n873_));
  NAND2_X1   g00615(.A1(new_n873_), .A2(new_n872_), .ZN(new_n874_));
  XOR2_X1    g00616(.A1(new_n844_), .A2(new_n850_), .Z(new_n875_));
  NAND2_X1   g00617(.A1(new_n875_), .A2(new_n841_), .ZN(new_n876_));
  NAND2_X1   g00618(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1   g00619(.A1(new_n877_), .A2(new_n758_), .ZN(new_n878_));
  NAND2_X1   g00620(.A1(new_n878_), .A2(new_n763_), .ZN(new_n879_));
  NAND4_X1   g00621(.A1(new_n874_), .A2(new_n876_), .A3(new_n756_), .A4(new_n757_), .ZN(new_n880_));
  NAND3_X1   g00622(.A1(new_n879_), .A2(new_n730_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1     g00623(.I(new_n881_), .ZN(new_n882_));
  INV_X1     g00624(.I(new_n840_), .ZN(new_n883_));
  NAND2_X1   g00625(.A1(new_n836_), .A2(new_n883_), .ZN(new_n884_));
  OAI22_X1   g00626(.A1(new_n448_), .A2(new_n472_), .B1(new_n515_), .B2(new_n450_), .ZN(new_n885_));
  OAI21_X1   g00627(.A1(new_n420_), .A2(new_n496_), .B(new_n885_), .ZN(new_n886_));
  AOI21_X1   g00628(.A1(new_n886_), .A2(new_n452_), .B(new_n448_), .ZN(new_n887_));
  XOR2_X1    g00629(.A1(new_n700_), .A2(new_n887_), .Z(new_n888_));
  NOR4_X1    g00630(.A1(new_n824_), .A2(new_n827_), .A3(new_n801_), .A4(new_n825_), .ZN(new_n889_));
  OAI21_X1   g00631(.A1(\b[1] ), .A2(new_n282_), .B(new_n817_), .ZN(new_n890_));
  OAI21_X1   g00632(.A1(new_n280_), .A2(new_n820_), .B(new_n890_), .ZN(new_n891_));
  INV_X1     g00633(.I(new_n816_), .ZN(new_n892_));
  XOR2_X1    g00634(.A1(\a[11] ), .A2(\a[14] ), .Z(new_n893_));
  NAND3_X1   g00635(.A1(new_n892_), .A2(new_n744_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1     g00636(.I(new_n894_), .ZN(new_n895_));
  NAND3_X1   g00637(.A1(new_n891_), .A2(\b[0] ), .A3(new_n895_), .ZN(new_n896_));
  XOR2_X1    g00638(.A1(new_n896_), .A2(\a[14] ), .Z(new_n897_));
  XNOR2_X1   g00639(.A1(new_n897_), .A2(new_n889_), .ZN(new_n898_));
  INV_X1     g00640(.I(new_n898_), .ZN(new_n899_));
  NAND2_X1   g00641(.A1(new_n804_), .A2(new_n831_), .ZN(new_n900_));
  NAND2_X1   g00642(.A1(new_n900_), .A2(new_n833_), .ZN(new_n901_));
  OAI22_X1   g00643(.A1(new_n607_), .A2(new_n325_), .B1(new_n610_), .B2(new_n419_), .ZN(new_n902_));
  OAI21_X1   g00644(.A1(new_n298_), .A2(new_n684_), .B(new_n902_), .ZN(new_n903_));
  AOI21_X1   g00645(.A1(new_n378_), .A2(new_n606_), .B(new_n903_), .ZN(new_n904_));
  XOR2_X1    g00646(.A1(new_n904_), .A2(new_n612_), .Z(new_n905_));
  XOR2_X1    g00647(.A1(new_n901_), .A2(new_n905_), .Z(new_n906_));
  XOR2_X1    g00648(.A1(new_n906_), .A2(new_n899_), .Z(new_n907_));
  XOR2_X1    g00649(.A1(new_n907_), .A2(new_n888_), .Z(new_n908_));
  NAND2_X1   g00650(.A1(new_n908_), .A2(new_n872_), .ZN(new_n909_));
  XNOR2_X1   g00651(.A1(new_n909_), .A2(new_n884_), .ZN(new_n910_));
  XOR2_X1    g00652(.A1(new_n910_), .A2(new_n844_), .Z(new_n911_));
  OAI22_X1   g00653(.A1(new_n656_), .A2(new_n341_), .B1(new_n404_), .B2(new_n706_), .ZN(new_n912_));
  OAI21_X1   g00654(.A1(new_n565_), .A2(new_n366_), .B(new_n912_), .ZN(new_n913_));
  AOI21_X1   g00655(.A1(new_n913_), .A2(new_n334_), .B(new_n341_), .ZN(new_n914_));
  XNOR2_X1   g00656(.A1(new_n710_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1     g00657(.I(new_n915_), .ZN(new_n916_));
  XOR2_X1    g00658(.A1(new_n911_), .A2(new_n916_), .Z(new_n917_));
  NOR2_X1    g00659(.A1(\b[12] ), .A2(\b[13] ), .ZN(new_n918_));
  INV_X1     g00660(.I(new_n918_), .ZN(new_n919_));
  OAI21_X1   g00661(.A1(new_n779_), .A2(new_n919_), .B(\b[11] ), .ZN(new_n920_));
  NOR2_X1    g00662(.A1(new_n780_), .A2(new_n861_), .ZN(new_n921_));
  NAND2_X1   g00663(.A1(new_n779_), .A2(new_n921_), .ZN(new_n922_));
  XNOR2_X1   g00664(.A1(\b[13] ), .A2(\b[14] ), .ZN(new_n923_));
  AOI21_X1   g00665(.A1(new_n920_), .A2(new_n922_), .B(new_n923_), .ZN(new_n924_));
  INV_X1     g00666(.I(new_n924_), .ZN(new_n925_));
  AOI21_X1   g00667(.A1(new_n775_), .A2(new_n918_), .B(new_n706_), .ZN(new_n926_));
  INV_X1     g00668(.I(new_n921_), .ZN(new_n927_));
  NOR2_X1    g00669(.A1(new_n775_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1    g00670(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1     g00671(.I(\b[14] ), .ZN(new_n930_));
  NOR2_X1    g00672(.A1(new_n861_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1     g00673(.I(new_n931_), .ZN(new_n932_));
  NAND2_X1   g00674(.A1(new_n861_), .A2(new_n930_), .ZN(new_n933_));
  AND2_X2    g00675(.A1(new_n932_), .A2(new_n933_), .Z(new_n934_));
  INV_X1     g00676(.I(new_n934_), .ZN(new_n935_));
  NAND2_X1   g00677(.A1(new_n929_), .A2(new_n935_), .ZN(new_n936_));
  NAND2_X1   g00678(.A1(new_n936_), .A2(new_n925_), .ZN(new_n937_));
  OAI22_X1   g00679(.A1(new_n330_), .A2(new_n861_), .B1(new_n930_), .B2(new_n263_), .ZN(new_n938_));
  OAI21_X1   g00680(.A1(new_n780_), .A2(new_n289_), .B(new_n938_), .ZN(new_n939_));
  AOI21_X1   g00681(.A1(new_n939_), .A2(new_n260_), .B(new_n426_), .ZN(new_n940_));
  XOR2_X1    g00682(.A1(new_n937_), .A2(new_n940_), .Z(new_n941_));
  NAND2_X1   g00683(.A1(new_n917_), .A2(new_n941_), .ZN(new_n942_));
  XOR2_X1    g00684(.A1(new_n942_), .A2(new_n853_), .Z(new_n943_));
  XOR2_X1    g00685(.A1(new_n943_), .A2(new_n882_), .Z(new_n944_));
  INV_X1     g00686(.I(new_n944_), .ZN(new_n945_));
  NAND2_X1   g00687(.A1(new_n945_), .A2(new_n867_), .ZN(new_n946_));
  XOR2_X1    g00688(.A1(new_n946_), .A2(new_n871_), .Z(new_n947_));
  XOR2_X1    g00689(.A1(new_n947_), .A2(new_n797_), .Z(\f[14] ));
  XOR2_X1    g00690(.A1(new_n942_), .A2(new_n881_), .Z(new_n949_));
  NAND2_X1   g00691(.A1(new_n949_), .A2(new_n853_), .ZN(new_n950_));
  AOI21_X1   g00692(.A1(new_n945_), .A2(new_n866_), .B(new_n857_), .ZN(new_n951_));
  OAI21_X1   g00693(.A1(new_n945_), .A2(new_n866_), .B(new_n797_), .ZN(new_n952_));
  NOR2_X1    g00694(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  OR2_X2     g00695(.A1(new_n881_), .A2(new_n911_), .Z(new_n954_));
  NAND2_X1   g00696(.A1(new_n881_), .A2(new_n911_), .ZN(new_n955_));
  NAND3_X1   g00697(.A1(new_n955_), .A2(new_n853_), .A3(new_n916_), .ZN(new_n956_));
  NAND2_X1   g00698(.A1(new_n956_), .A2(new_n954_), .ZN(new_n957_));
  INV_X1     g00699(.I(new_n957_), .ZN(new_n958_));
  INV_X1     g00700(.I(new_n897_), .ZN(new_n959_));
  XOR2_X1    g00701(.A1(new_n889_), .A2(new_n904_), .Z(new_n960_));
  XOR2_X1    g00702(.A1(new_n960_), .A2(new_n959_), .Z(new_n961_));
  XOR2_X1    g00703(.A1(new_n961_), .A2(\a[11] ), .Z(new_n962_));
  NAND2_X1   g00704(.A1(new_n962_), .A2(new_n829_), .ZN(new_n963_));
  NAND2_X1   g00705(.A1(new_n963_), .A2(new_n811_), .ZN(new_n964_));
  NOR2_X1    g00706(.A1(new_n962_), .A2(new_n829_), .ZN(new_n965_));
  NOR2_X1    g00707(.A1(new_n965_), .A2(new_n805_), .ZN(new_n966_));
  NAND2_X1   g00708(.A1(new_n966_), .A2(new_n964_), .ZN(new_n967_));
  NAND2_X1   g00709(.A1(new_n899_), .A2(new_n905_), .ZN(new_n968_));
  INV_X1     g00710(.I(new_n968_), .ZN(new_n969_));
  INV_X1     g00711(.I(new_n817_), .ZN(new_n970_));
  OAI22_X1   g00712(.A1(new_n970_), .A2(new_n280_), .B1(new_n298_), .B2(new_n820_), .ZN(new_n971_));
  AOI21_X1   g00713(.A1(\b[1] ), .A2(new_n895_), .B(new_n971_), .ZN(new_n972_));
  NOR3_X1    g00714(.A1(new_n972_), .A2(new_n403_), .A3(new_n970_), .ZN(new_n973_));
  XOR2_X1    g00715(.A1(new_n973_), .A2(new_n827_), .Z(new_n974_));
  XOR2_X1    g00716(.A1(\a[14] ), .A2(\a[15] ), .Z(new_n975_));
  NAND2_X1   g00717(.A1(new_n975_), .A2(\b[0] ), .ZN(new_n976_));
  NOR2_X1    g00718(.A1(new_n974_), .A2(new_n976_), .ZN(new_n977_));
  XOR2_X1    g00719(.A1(new_n977_), .A2(new_n897_), .Z(new_n978_));
  XOR2_X1    g00720(.A1(new_n978_), .A2(new_n889_), .Z(new_n979_));
  INV_X1     g00721(.I(new_n979_), .ZN(new_n980_));
  OAI22_X1   g00722(.A1(new_n607_), .A2(new_n419_), .B1(new_n610_), .B2(new_n420_), .ZN(new_n981_));
  OAI21_X1   g00723(.A1(new_n325_), .A2(new_n684_), .B(new_n981_), .ZN(new_n982_));
  AOI21_X1   g00724(.A1(new_n982_), .A2(new_n612_), .B(new_n607_), .ZN(new_n983_));
  XOR2_X1    g00725(.A1(new_n556_), .A2(new_n983_), .Z(new_n984_));
  NAND2_X1   g00726(.A1(new_n980_), .A2(new_n984_), .ZN(new_n985_));
  XOR2_X1    g00727(.A1(new_n985_), .A2(new_n969_), .Z(new_n986_));
  XNOR2_X1   g00728(.A1(new_n986_), .A2(new_n967_), .ZN(new_n987_));
  OAI22_X1   g00729(.A1(new_n448_), .A2(new_n515_), .B1(new_n565_), .B2(new_n450_), .ZN(new_n988_));
  OAI21_X1   g00730(.A1(new_n472_), .A2(new_n496_), .B(new_n988_), .ZN(new_n989_));
  AOI21_X1   g00731(.A1(new_n989_), .A2(new_n452_), .B(new_n448_), .ZN(new_n990_));
  XOR2_X1    g00732(.A1(new_n759_), .A2(new_n990_), .Z(new_n991_));
  INV_X1     g00733(.I(new_n991_), .ZN(new_n992_));
  XOR2_X1    g00734(.A1(new_n987_), .A2(new_n992_), .Z(new_n993_));
  INV_X1     g00735(.I(new_n993_), .ZN(new_n994_));
  AOI21_X1   g00736(.A1(new_n908_), .A2(new_n836_), .B(new_n883_), .ZN(new_n995_));
  OAI21_X1   g00737(.A1(new_n908_), .A2(new_n836_), .B(new_n844_), .ZN(new_n996_));
  XOR2_X1    g00738(.A1(new_n901_), .A2(new_n898_), .Z(new_n997_));
  XNOR2_X1   g00739(.A1(new_n997_), .A2(new_n905_), .ZN(new_n998_));
  NOR2_X1    g00740(.A1(new_n998_), .A2(new_n888_), .ZN(new_n999_));
  INV_X1     g00741(.I(new_n999_), .ZN(new_n1000_));
  OAI21_X1   g00742(.A1(new_n995_), .A2(new_n996_), .B(new_n1000_), .ZN(new_n1001_));
  NOR2_X1    g00743(.A1(new_n995_), .A2(new_n996_), .ZN(new_n1002_));
  NOR3_X1    g00744(.A1(new_n994_), .A2(new_n1002_), .A3(new_n999_), .ZN(new_n1003_));
  AOI21_X1   g00745(.A1(new_n994_), .A2(new_n1001_), .B(new_n1003_), .ZN(new_n1004_));
  OAI22_X1   g00746(.A1(new_n706_), .A2(new_n341_), .B1(new_n404_), .B2(new_n780_), .ZN(new_n1005_));
  OAI21_X1   g00747(.A1(new_n656_), .A2(new_n366_), .B(new_n1005_), .ZN(new_n1006_));
  AOI21_X1   g00748(.A1(new_n1006_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1007_));
  XOR2_X1    g00749(.A1(new_n785_), .A2(new_n1007_), .Z(new_n1008_));
  OR2_X2     g00750(.A1(new_n1004_), .A2(new_n1008_), .Z(new_n1009_));
  NAND2_X1   g00751(.A1(new_n1004_), .A2(new_n1008_), .ZN(new_n1010_));
  AOI21_X1   g00752(.A1(new_n1009_), .A2(new_n1010_), .B(new_n958_), .ZN(new_n1011_));
  XNOR2_X1   g00753(.A1(new_n1004_), .A2(new_n1008_), .ZN(new_n1012_));
  NOR2_X1    g00754(.A1(new_n957_), .A2(new_n1012_), .ZN(new_n1013_));
  NOR2_X1    g00755(.A1(new_n1011_), .A2(new_n1013_), .ZN(new_n1014_));
  NAND2_X1   g00756(.A1(new_n920_), .A2(new_n922_), .ZN(new_n1015_));
  INV_X1     g00757(.I(new_n923_), .ZN(new_n1016_));
  INV_X1     g00758(.I(\b[15] ), .ZN(new_n1017_));
  NOR2_X1    g00759(.A1(new_n1017_), .A2(\b[13] ), .ZN(new_n1018_));
  NOR2_X1    g00760(.A1(new_n861_), .A2(\b[15] ), .ZN(new_n1019_));
  OAI21_X1   g00761(.A1(new_n1018_), .A2(new_n1019_), .B(new_n1016_), .ZN(new_n1020_));
  NOR2_X1    g00762(.A1(new_n1015_), .A2(new_n1020_), .ZN(new_n1021_));
  NAND2_X1   g00763(.A1(new_n1015_), .A2(new_n1020_), .ZN(new_n1022_));
  INV_X1     g00764(.I(new_n1022_), .ZN(new_n1023_));
  NOR2_X1    g00765(.A1(new_n1023_), .A2(new_n1021_), .ZN(new_n1024_));
  OAI22_X1   g00766(.A1(new_n330_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n263_), .ZN(new_n1025_));
  OAI21_X1   g00767(.A1(new_n861_), .A2(new_n289_), .B(new_n1025_), .ZN(new_n1026_));
  AOI21_X1   g00768(.A1(new_n1026_), .A2(new_n260_), .B(new_n426_), .ZN(new_n1027_));
  XOR2_X1    g00769(.A1(new_n1024_), .A2(new_n1027_), .Z(new_n1028_));
  NOR2_X1    g00770(.A1(new_n1014_), .A2(new_n1028_), .ZN(new_n1029_));
  XNOR2_X1   g00771(.A1(new_n953_), .A2(new_n1029_), .ZN(new_n1030_));
  XOR2_X1    g00772(.A1(new_n1030_), .A2(new_n950_), .Z(\f[15] ));
  OAI21_X1   g00773(.A1(new_n1011_), .A2(new_n1013_), .B(new_n953_), .ZN(new_n1032_));
  INV_X1     g00774(.I(new_n1014_), .ZN(new_n1033_));
  NOR2_X1    g00775(.A1(new_n950_), .A2(new_n1028_), .ZN(new_n1034_));
  OAI21_X1   g00776(.A1(new_n953_), .A2(new_n1033_), .B(new_n1034_), .ZN(new_n1035_));
  NAND2_X1   g00777(.A1(new_n1032_), .A2(new_n1035_), .ZN(new_n1036_));
  NOR2_X1    g00778(.A1(new_n987_), .A2(new_n1000_), .ZN(new_n1037_));
  NAND2_X1   g00779(.A1(new_n987_), .A2(new_n1000_), .ZN(new_n1038_));
  AND3_X2    g00780(.A1(new_n1002_), .A2(new_n992_), .A3(new_n1038_), .Z(new_n1039_));
  NOR2_X1    g00781(.A1(new_n1039_), .A2(new_n1037_), .ZN(new_n1040_));
  NOR2_X1    g00782(.A1(new_n967_), .A2(new_n979_), .ZN(new_n1041_));
  NAND2_X1   g00783(.A1(new_n969_), .A2(new_n984_), .ZN(new_n1042_));
  AOI21_X1   g00784(.A1(new_n967_), .A2(new_n979_), .B(new_n1042_), .ZN(new_n1043_));
  NOR2_X1    g00785(.A1(new_n1043_), .A2(new_n1041_), .ZN(new_n1044_));
  INV_X1     g00786(.I(new_n976_), .ZN(new_n1045_));
  NAND2_X1   g00787(.A1(new_n974_), .A2(new_n897_), .ZN(new_n1046_));
  NAND3_X1   g00788(.A1(new_n1046_), .A2(new_n889_), .A3(new_n1045_), .ZN(new_n1047_));
  OAI21_X1   g00789(.A1(new_n897_), .A2(new_n974_), .B(new_n1047_), .ZN(new_n1048_));
  OAI22_X1   g00790(.A1(new_n970_), .A2(new_n298_), .B1(new_n325_), .B2(new_n820_), .ZN(new_n1049_));
  OAI21_X1   g00791(.A1(new_n280_), .A2(new_n894_), .B(new_n1049_), .ZN(new_n1050_));
  AOI21_X1   g00792(.A1(new_n1050_), .A2(new_n827_), .B(new_n970_), .ZN(new_n1051_));
  XOR2_X1    g00793(.A1(new_n1051_), .A2(new_n807_), .Z(new_n1052_));
  XOR2_X1    g00794(.A1(\a[15] ), .A2(\a[17] ), .Z(new_n1053_));
  XOR2_X1    g00795(.A1(\a[14] ), .A2(\a[16] ), .Z(new_n1054_));
  NAND2_X1   g00796(.A1(new_n1054_), .A2(new_n1053_), .ZN(new_n1055_));
  INV_X1     g00797(.I(new_n1055_), .ZN(new_n1056_));
  INV_X1     g00798(.I(\a[17] ), .ZN(new_n1057_));
  INV_X1     g00799(.I(\a[15] ), .ZN(new_n1058_));
  AND3_X2    g00800(.A1(new_n827_), .A2(new_n1058_), .A3(\a[16] ), .Z(new_n1059_));
  NOR3_X1    g00801(.A1(new_n827_), .A2(new_n1058_), .A3(\a[16] ), .ZN(new_n1060_));
  NOR2_X1    g00802(.A1(new_n1059_), .A2(new_n1060_), .ZN(new_n1061_));
  NOR2_X1    g00803(.A1(new_n1061_), .A2(new_n269_), .ZN(new_n1062_));
  INV_X1     g00804(.I(new_n1062_), .ZN(new_n1063_));
  NAND2_X1   g00805(.A1(new_n1056_), .A2(\b[0] ), .ZN(new_n1064_));
  NAND3_X1   g00806(.A1(new_n1064_), .A2(new_n1063_), .A3(new_n1057_), .ZN(new_n1065_));
  NAND2_X1   g00807(.A1(new_n1065_), .A2(new_n1056_), .ZN(new_n1066_));
  NOR2_X1    g00808(.A1(new_n1066_), .A2(new_n271_), .ZN(new_n1067_));
  AOI21_X1   g00809(.A1(new_n1065_), .A2(new_n1056_), .B(new_n444_), .ZN(new_n1068_));
  NOR2_X1    g00810(.A1(new_n1067_), .A2(new_n1068_), .ZN(new_n1069_));
  NOR2_X1    g00811(.A1(new_n1045_), .A2(new_n1057_), .ZN(new_n1070_));
  XOR2_X1    g00812(.A1(new_n1069_), .A2(new_n1070_), .Z(new_n1071_));
  XOR2_X1    g00813(.A1(new_n1071_), .A2(new_n1052_), .Z(new_n1072_));
  NAND2_X1   g00814(.A1(new_n1071_), .A2(new_n1052_), .ZN(new_n1073_));
  OR2_X2     g00815(.A1(new_n1071_), .A2(new_n1052_), .Z(new_n1074_));
  NAND2_X1   g00816(.A1(new_n1074_), .A2(new_n1073_), .ZN(new_n1075_));
  MUX2_X1    g00817(.I0(new_n1075_), .I1(new_n1072_), .S(new_n1048_), .Z(new_n1076_));
  AOI22_X1   g00818(.A1(new_n611_), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n606_), .ZN(new_n1077_));
  AOI21_X1   g00819(.A1(\b[5] ), .A2(new_n739_), .B(new_n1077_), .ZN(new_n1078_));
  OAI21_X1   g00820(.A1(new_n1078_), .A2(\a[11] ), .B(new_n606_), .ZN(new_n1079_));
  XNOR2_X1   g00821(.A1(new_n1079_), .A2(new_n471_), .ZN(new_n1080_));
  INV_X1     g00822(.I(new_n1080_), .ZN(new_n1081_));
  XOR2_X1    g00823(.A1(new_n1076_), .A2(new_n1081_), .Z(new_n1082_));
  NOR2_X1    g00824(.A1(new_n1044_), .A2(new_n1082_), .ZN(new_n1083_));
  XOR2_X1    g00825(.A1(new_n1076_), .A2(new_n1081_), .Z(new_n1084_));
  AND2_X2    g00826(.A1(new_n1044_), .A2(new_n1084_), .Z(new_n1085_));
  NOR2_X1    g00827(.A1(new_n1085_), .A2(new_n1083_), .ZN(new_n1086_));
  OAI22_X1   g00828(.A1(new_n448_), .A2(new_n565_), .B1(new_n656_), .B2(new_n450_), .ZN(new_n1087_));
  OAI21_X1   g00829(.A1(new_n515_), .A2(new_n496_), .B(new_n1087_), .ZN(new_n1088_));
  AOI21_X1   g00830(.A1(new_n1088_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1089_));
  XNOR2_X1   g00831(.A1(new_n660_), .A2(new_n1089_), .ZN(new_n1090_));
  XOR2_X1    g00832(.A1(new_n1086_), .A2(new_n1090_), .Z(new_n1091_));
  OAI22_X1   g00833(.A1(new_n780_), .A2(new_n341_), .B1(new_n404_), .B2(new_n861_), .ZN(new_n1092_));
  OAI21_X1   g00834(.A1(new_n706_), .A2(new_n366_), .B(new_n1092_), .ZN(new_n1093_));
  AOI21_X1   g00835(.A1(new_n1093_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1094_));
  XNOR2_X1   g00836(.A1(new_n860_), .A2(new_n1094_), .ZN(new_n1095_));
  XOR2_X1    g00837(.A1(new_n1091_), .A2(new_n1095_), .Z(new_n1096_));
  NOR2_X1    g00838(.A1(new_n1096_), .A2(new_n1040_), .ZN(new_n1097_));
  XOR2_X1    g00839(.A1(new_n1091_), .A2(new_n1095_), .Z(new_n1098_));
  AOI21_X1   g00840(.A1(new_n1040_), .A2(new_n1098_), .B(new_n1097_), .ZN(new_n1099_));
  NOR2_X1    g00841(.A1(new_n1099_), .A2(new_n1012_), .ZN(new_n1100_));
  XOR2_X1    g00842(.A1(new_n1100_), .A2(new_n1009_), .Z(new_n1101_));
  XOR2_X1    g00843(.A1(new_n1101_), .A2(new_n958_), .Z(new_n1102_));
  NOR4_X1    g00844(.A1(new_n926_), .A2(new_n928_), .A3(\b[14] ), .A4(\b[15] ), .ZN(new_n1103_));
  NOR2_X1    g00845(.A1(new_n930_), .A2(new_n1017_), .ZN(new_n1104_));
  INV_X1     g00846(.I(new_n1104_), .ZN(new_n1105_));
  OAI22_X1   g00847(.A1(new_n1103_), .A2(new_n861_), .B1(new_n929_), .B2(new_n1105_), .ZN(new_n1106_));
  XNOR2_X1   g00848(.A1(\b[15] ), .A2(\b[16] ), .ZN(new_n1107_));
  INV_X1     g00849(.I(new_n1107_), .ZN(new_n1108_));
  INV_X1     g00850(.I(\b[16] ), .ZN(new_n1109_));
  NOR2_X1    g00851(.A1(new_n1017_), .A2(new_n1109_), .ZN(new_n1110_));
  INV_X1     g00852(.I(new_n1110_), .ZN(new_n1111_));
  NAND2_X1   g00853(.A1(new_n1017_), .A2(new_n1109_), .ZN(new_n1112_));
  AOI21_X1   g00854(.A1(new_n1111_), .A2(new_n1112_), .B(new_n1106_), .ZN(new_n1113_));
  AOI21_X1   g00855(.A1(new_n1106_), .A2(new_n1108_), .B(new_n1113_), .ZN(new_n1114_));
  OAI22_X1   g00856(.A1(new_n330_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n263_), .ZN(new_n1115_));
  OAI21_X1   g00857(.A1(new_n930_), .A2(new_n289_), .B(new_n1115_), .ZN(new_n1116_));
  AOI21_X1   g00858(.A1(new_n1116_), .A2(new_n260_), .B(new_n426_), .ZN(new_n1117_));
  XOR2_X1    g00859(.A1(new_n1114_), .A2(new_n1117_), .Z(new_n1118_));
  XOR2_X1    g00860(.A1(new_n1102_), .A2(new_n1118_), .Z(new_n1119_));
  NAND2_X1   g00861(.A1(new_n1036_), .A2(new_n1119_), .ZN(new_n1120_));
  XOR2_X1    g00862(.A1(new_n1102_), .A2(new_n1118_), .Z(new_n1121_));
  OAI21_X1   g00863(.A1(new_n1036_), .A2(new_n1121_), .B(new_n1120_), .ZN(\f[16] ));
  INV_X1     g00864(.I(new_n1118_), .ZN(new_n1123_));
  NAND2_X1   g00865(.A1(new_n1102_), .A2(new_n1123_), .ZN(new_n1124_));
  INV_X1     g00866(.I(new_n1095_), .ZN(new_n1125_));
  XOR2_X1    g00867(.A1(new_n1040_), .A2(new_n1091_), .Z(new_n1126_));
  NOR2_X1    g00868(.A1(new_n1126_), .A2(new_n1125_), .ZN(new_n1127_));
  OAI21_X1   g00869(.A1(new_n1099_), .A2(new_n1004_), .B(new_n1008_), .ZN(new_n1128_));
  NAND2_X1   g00870(.A1(new_n1099_), .A2(new_n1004_), .ZN(new_n1129_));
  NAND3_X1   g00871(.A1(new_n957_), .A2(new_n1128_), .A3(new_n1129_), .ZN(new_n1130_));
  INV_X1     g00872(.I(new_n1130_), .ZN(new_n1131_));
  NOR2_X1    g00873(.A1(new_n1086_), .A2(new_n1090_), .ZN(new_n1132_));
  NAND2_X1   g00874(.A1(new_n1076_), .A2(new_n1081_), .ZN(new_n1133_));
  OAI22_X1   g00875(.A1(new_n607_), .A2(new_n472_), .B1(new_n515_), .B2(new_n610_), .ZN(new_n1134_));
  OAI21_X1   g00876(.A1(new_n420_), .A2(new_n684_), .B(new_n1134_), .ZN(new_n1135_));
  AOI21_X1   g00877(.A1(new_n1135_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1136_));
  XOR2_X1    g00878(.A1(new_n700_), .A2(new_n1136_), .Z(new_n1137_));
  NAND2_X1   g00879(.A1(new_n1069_), .A2(new_n1070_), .ZN(new_n1138_));
  OAI21_X1   g00880(.A1(\b[1] ), .A2(new_n282_), .B(new_n1056_), .ZN(new_n1139_));
  OAI21_X1   g00881(.A1(new_n280_), .A2(new_n1061_), .B(new_n1139_), .ZN(new_n1140_));
  XOR2_X1    g00882(.A1(\a[14] ), .A2(\a[17] ), .Z(new_n1141_));
  AND3_X2    g00883(.A1(new_n1054_), .A2(new_n975_), .A3(new_n1141_), .Z(new_n1142_));
  NAND3_X1   g00884(.A1(new_n1140_), .A2(\b[0] ), .A3(new_n1142_), .ZN(new_n1143_));
  XOR2_X1    g00885(.A1(new_n1143_), .A2(\a[17] ), .Z(new_n1144_));
  XOR2_X1    g00886(.A1(new_n1144_), .A2(new_n1138_), .Z(new_n1145_));
  NAND2_X1   g00887(.A1(new_n1048_), .A2(new_n1073_), .ZN(new_n1146_));
  NAND2_X1   g00888(.A1(new_n1146_), .A2(new_n1074_), .ZN(new_n1147_));
  OAI22_X1   g00889(.A1(new_n970_), .A2(new_n325_), .B1(new_n419_), .B2(new_n820_), .ZN(new_n1148_));
  OAI21_X1   g00890(.A1(new_n298_), .A2(new_n894_), .B(new_n1148_), .ZN(new_n1149_));
  AOI21_X1   g00891(.A1(new_n378_), .A2(new_n817_), .B(new_n1149_), .ZN(new_n1150_));
  XOR2_X1    g00892(.A1(new_n1150_), .A2(new_n827_), .Z(new_n1151_));
  INV_X1     g00893(.I(new_n1151_), .ZN(new_n1152_));
  XOR2_X1    g00894(.A1(new_n1147_), .A2(new_n1152_), .Z(new_n1153_));
  XOR2_X1    g00895(.A1(new_n1153_), .A2(new_n1145_), .Z(new_n1154_));
  XOR2_X1    g00896(.A1(new_n1154_), .A2(new_n1137_), .Z(new_n1155_));
  NAND2_X1   g00897(.A1(new_n1155_), .A2(new_n1084_), .ZN(new_n1156_));
  XOR2_X1    g00898(.A1(new_n1156_), .A2(new_n1133_), .Z(new_n1157_));
  NAND2_X1   g00899(.A1(new_n1157_), .A2(new_n1044_), .ZN(new_n1158_));
  INV_X1     g00900(.I(new_n1044_), .ZN(new_n1159_));
  XNOR2_X1   g00901(.A1(new_n1156_), .A2(new_n1133_), .ZN(new_n1160_));
  NAND2_X1   g00902(.A1(new_n1160_), .A2(new_n1159_), .ZN(new_n1161_));
  OAI22_X1   g00903(.A1(new_n448_), .A2(new_n656_), .B1(new_n706_), .B2(new_n450_), .ZN(new_n1162_));
  OAI21_X1   g00904(.A1(new_n565_), .A2(new_n496_), .B(new_n1162_), .ZN(new_n1163_));
  AOI21_X1   g00905(.A1(new_n1163_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1164_));
  XNOR2_X1   g00906(.A1(new_n710_), .A2(new_n1164_), .ZN(new_n1165_));
  AOI21_X1   g00907(.A1(new_n1161_), .A2(new_n1158_), .B(new_n1165_), .ZN(new_n1166_));
  NOR2_X1    g00908(.A1(new_n1160_), .A2(new_n1159_), .ZN(new_n1167_));
  NOR2_X1    g00909(.A1(new_n1157_), .A2(new_n1044_), .ZN(new_n1168_));
  INV_X1     g00910(.I(new_n1165_), .ZN(new_n1169_));
  NOR3_X1    g00911(.A1(new_n1167_), .A2(new_n1168_), .A3(new_n1169_), .ZN(new_n1170_));
  NOR2_X1    g00912(.A1(new_n1170_), .A2(new_n1166_), .ZN(new_n1171_));
  XNOR2_X1   g00913(.A1(new_n1086_), .A2(new_n1090_), .ZN(new_n1172_));
  NOR3_X1    g00914(.A1(new_n1171_), .A2(new_n1132_), .A3(new_n1172_), .ZN(new_n1173_));
  NOR2_X1    g00915(.A1(new_n1086_), .A2(new_n1090_), .ZN(new_n1174_));
  NOR2_X1    g00916(.A1(new_n1173_), .A2(new_n1174_), .ZN(new_n1175_));
  NOR3_X1    g00917(.A1(new_n1175_), .A2(new_n1037_), .A3(new_n1039_), .ZN(new_n1176_));
  NOR3_X1    g00918(.A1(new_n1173_), .A2(new_n1040_), .A3(new_n1174_), .ZN(new_n1177_));
  NOR2_X1    g00919(.A1(new_n1176_), .A2(new_n1177_), .ZN(new_n1178_));
  OAI22_X1   g00920(.A1(new_n861_), .A2(new_n341_), .B1(new_n404_), .B2(new_n930_), .ZN(new_n1179_));
  OAI21_X1   g00921(.A1(new_n780_), .A2(new_n366_), .B(new_n1179_), .ZN(new_n1180_));
  AOI21_X1   g00922(.A1(new_n1180_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1181_));
  XNOR2_X1   g00923(.A1(new_n937_), .A2(new_n1181_), .ZN(new_n1182_));
  INV_X1     g00924(.I(new_n1182_), .ZN(new_n1183_));
  XOR2_X1    g00925(.A1(new_n1178_), .A2(new_n1183_), .Z(new_n1184_));
  NOR2_X1    g00926(.A1(\b[14] ), .A2(\b[15] ), .ZN(new_n1185_));
  AOI21_X1   g00927(.A1(new_n929_), .A2(new_n1185_), .B(new_n861_), .ZN(new_n1186_));
  NOR2_X1    g00928(.A1(new_n929_), .A2(new_n1105_), .ZN(new_n1187_));
  NOR2_X1    g00929(.A1(new_n1186_), .A2(new_n1187_), .ZN(new_n1188_));
  INV_X1     g00930(.I(\b[17] ), .ZN(new_n1189_));
  NOR2_X1    g00931(.A1(new_n1189_), .A2(\b[15] ), .ZN(new_n1190_));
  NOR2_X1    g00932(.A1(new_n1017_), .A2(\b[17] ), .ZN(new_n1191_));
  OAI21_X1   g00933(.A1(new_n1190_), .A2(new_n1191_), .B(new_n1108_), .ZN(new_n1192_));
  INV_X1     g00934(.I(new_n1192_), .ZN(new_n1193_));
  NAND2_X1   g00935(.A1(new_n1188_), .A2(new_n1193_), .ZN(new_n1194_));
  NAND2_X1   g00936(.A1(new_n1106_), .A2(new_n1192_), .ZN(new_n1195_));
  NAND2_X1   g00937(.A1(new_n1194_), .A2(new_n1195_), .ZN(new_n1196_));
  OAI22_X1   g00938(.A1(new_n330_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n263_), .ZN(new_n1197_));
  OAI21_X1   g00939(.A1(new_n1017_), .A2(new_n289_), .B(new_n1197_), .ZN(new_n1198_));
  AOI21_X1   g00940(.A1(new_n1198_), .A2(new_n260_), .B(new_n426_), .ZN(new_n1199_));
  XOR2_X1    g00941(.A1(new_n1196_), .A2(new_n1199_), .Z(new_n1200_));
  NAND2_X1   g00942(.A1(new_n1184_), .A2(new_n1200_), .ZN(new_n1201_));
  NOR2_X1    g00943(.A1(new_n1201_), .A2(new_n1131_), .ZN(new_n1202_));
  NAND2_X1   g00944(.A1(new_n1201_), .A2(new_n1131_), .ZN(new_n1203_));
  INV_X1     g00945(.I(new_n1203_), .ZN(new_n1204_));
  NOR2_X1    g00946(.A1(new_n1204_), .A2(new_n1202_), .ZN(new_n1205_));
  NOR2_X1    g00947(.A1(new_n1205_), .A2(new_n1127_), .ZN(new_n1206_));
  NOR4_X1    g00948(.A1(new_n1204_), .A2(new_n1125_), .A3(new_n1126_), .A4(new_n1202_), .ZN(new_n1207_));
  NOR2_X1    g00949(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1208_));
  NOR2_X1    g00950(.A1(new_n1208_), .A2(new_n1121_), .ZN(new_n1209_));
  XNOR2_X1   g00951(.A1(new_n1209_), .A2(new_n1124_), .ZN(new_n1210_));
  XOR2_X1    g00952(.A1(new_n1210_), .A2(new_n1036_), .Z(\f[17] ));
  OAI21_X1   g00953(.A1(new_n1176_), .A2(new_n1177_), .B(new_n1127_), .ZN(new_n1212_));
  NOR3_X1    g00954(.A1(new_n1176_), .A2(new_n1127_), .A3(new_n1177_), .ZN(new_n1213_));
  NAND4_X1   g00955(.A1(new_n957_), .A2(new_n1128_), .A3(new_n1129_), .A4(new_n1183_), .ZN(new_n1214_));
  OAI21_X1   g00956(.A1(new_n1214_), .A2(new_n1213_), .B(new_n1212_), .ZN(new_n1215_));
  INV_X1     g00957(.I(new_n1215_), .ZN(new_n1216_));
  AOI21_X1   g00958(.A1(new_n1161_), .A2(new_n1158_), .B(new_n1169_), .ZN(new_n1217_));
  INV_X1     g00959(.I(new_n1217_), .ZN(new_n1218_));
  OAI21_X1   g00960(.A1(new_n1171_), .A2(new_n1086_), .B(new_n1090_), .ZN(new_n1219_));
  AOI21_X1   g00961(.A1(new_n1171_), .A2(new_n1086_), .B(new_n1040_), .ZN(new_n1220_));
  XOR2_X1    g00962(.A1(new_n1147_), .A2(new_n1145_), .Z(new_n1221_));
  XOR2_X1    g00963(.A1(new_n1221_), .A2(new_n1152_), .Z(new_n1222_));
  NOR2_X1    g00964(.A1(new_n1222_), .A2(new_n1137_), .ZN(new_n1223_));
  AOI21_X1   g00965(.A1(new_n1155_), .A2(new_n1076_), .B(new_n1081_), .ZN(new_n1224_));
  OAI21_X1   g00966(.A1(new_n1155_), .A2(new_n1076_), .B(new_n1159_), .ZN(new_n1225_));
  OR2_X2     g00967(.A1(new_n1224_), .A2(new_n1225_), .Z(new_n1226_));
  XOR2_X1    g00968(.A1(\a[17] ), .A2(\a[18] ), .Z(new_n1227_));
  NAND2_X1   g00969(.A1(new_n1227_), .A2(\b[0] ), .ZN(new_n1228_));
  OAI22_X1   g00970(.A1(new_n280_), .A2(new_n1055_), .B1(new_n1061_), .B2(new_n298_), .ZN(new_n1229_));
  AOI21_X1   g00971(.A1(\b[1] ), .A2(new_n1142_), .B(new_n1229_), .ZN(new_n1230_));
  NOR3_X1    g00972(.A1(new_n1230_), .A2(new_n403_), .A3(new_n1055_), .ZN(new_n1231_));
  XOR2_X1    g00973(.A1(new_n1231_), .A2(new_n1057_), .Z(new_n1232_));
  INV_X1     g00974(.I(new_n1144_), .ZN(new_n1233_));
  NOR2_X1    g00975(.A1(new_n1233_), .A2(new_n1138_), .ZN(new_n1234_));
  INV_X1     g00976(.I(new_n820_), .ZN(new_n1235_));
  AOI22_X1   g00977(.A1(new_n1235_), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n817_), .ZN(new_n1236_));
  AOI21_X1   g00978(.A1(\b[4] ), .A2(new_n895_), .B(new_n1236_), .ZN(new_n1237_));
  OAI21_X1   g00979(.A1(new_n1237_), .A2(\a[14] ), .B(new_n817_), .ZN(new_n1238_));
  XOR2_X1    g00980(.A1(new_n556_), .A2(new_n1238_), .Z(new_n1239_));
  XNOR2_X1   g00981(.A1(new_n1234_), .A2(new_n1239_), .ZN(new_n1240_));
  XOR2_X1    g00982(.A1(new_n1240_), .A2(new_n1232_), .Z(new_n1241_));
  XOR2_X1    g00983(.A1(new_n1241_), .A2(new_n1228_), .Z(new_n1242_));
  NOR2_X1    g00984(.A1(new_n1145_), .A2(new_n1152_), .ZN(new_n1243_));
  INV_X1     g00985(.I(new_n1243_), .ZN(new_n1244_));
  INV_X1     g00986(.I(new_n1052_), .ZN(new_n1245_));
  XOR2_X1    g00987(.A1(new_n1138_), .A2(new_n1150_), .Z(new_n1246_));
  XOR2_X1    g00988(.A1(new_n1246_), .A2(new_n1144_), .Z(new_n1247_));
  XOR2_X1    g00989(.A1(new_n1247_), .A2(\a[14] ), .Z(new_n1248_));
  AOI21_X1   g00990(.A1(new_n1248_), .A2(new_n1071_), .B(new_n1245_), .ZN(new_n1249_));
  OAI21_X1   g00991(.A1(new_n1248_), .A2(new_n1071_), .B(new_n1048_), .ZN(new_n1250_));
  NOR2_X1    g00992(.A1(new_n1249_), .A2(new_n1250_), .ZN(new_n1251_));
  INV_X1     g00993(.I(new_n1251_), .ZN(new_n1252_));
  AOI21_X1   g00994(.A1(new_n1252_), .A2(new_n1244_), .B(new_n1242_), .ZN(new_n1253_));
  AND3_X2    g00995(.A1(new_n1252_), .A2(new_n1242_), .A3(new_n1244_), .Z(new_n1254_));
  NOR2_X1    g00996(.A1(new_n1254_), .A2(new_n1253_), .ZN(new_n1255_));
  OAI22_X1   g00997(.A1(new_n607_), .A2(new_n515_), .B1(new_n565_), .B2(new_n610_), .ZN(new_n1256_));
  OAI21_X1   g00998(.A1(new_n472_), .A2(new_n684_), .B(new_n1256_), .ZN(new_n1257_));
  AOI21_X1   g00999(.A1(new_n1257_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1258_));
  XOR2_X1    g01000(.A1(new_n759_), .A2(new_n1258_), .Z(new_n1259_));
  NOR2_X1    g01001(.A1(new_n1255_), .A2(new_n1259_), .ZN(new_n1260_));
  XOR2_X1    g01002(.A1(new_n1226_), .A2(new_n1260_), .Z(new_n1261_));
  NOR2_X1    g01003(.A1(new_n1261_), .A2(new_n1223_), .ZN(new_n1262_));
  INV_X1     g01004(.I(new_n1223_), .ZN(new_n1263_));
  XNOR2_X1   g01005(.A1(new_n1226_), .A2(new_n1260_), .ZN(new_n1264_));
  NOR2_X1    g01006(.A1(new_n1264_), .A2(new_n1263_), .ZN(new_n1265_));
  OAI22_X1   g01007(.A1(new_n448_), .A2(new_n706_), .B1(new_n780_), .B2(new_n450_), .ZN(new_n1266_));
  OAI21_X1   g01008(.A1(new_n656_), .A2(new_n496_), .B(new_n1266_), .ZN(new_n1267_));
  AOI21_X1   g01009(.A1(new_n1267_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1268_));
  XOR2_X1    g01010(.A1(new_n785_), .A2(new_n1268_), .Z(new_n1269_));
  INV_X1     g01011(.I(new_n1269_), .ZN(new_n1270_));
  OAI21_X1   g01012(.A1(new_n1265_), .A2(new_n1262_), .B(new_n1270_), .ZN(new_n1271_));
  AOI21_X1   g01013(.A1(new_n1220_), .A2(new_n1219_), .B(new_n1271_), .ZN(new_n1272_));
  AND3_X2    g01014(.A1(new_n1220_), .A2(new_n1219_), .A3(new_n1271_), .Z(new_n1273_));
  OAI21_X1   g01015(.A1(new_n1273_), .A2(new_n1272_), .B(new_n1218_), .ZN(new_n1274_));
  OR3_X2     g01016(.A1(new_n1273_), .A2(new_n1272_), .A3(new_n1218_), .Z(new_n1275_));
  OAI22_X1   g01017(.A1(new_n930_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1017_), .ZN(new_n1276_));
  OAI21_X1   g01018(.A1(new_n861_), .A2(new_n366_), .B(new_n1276_), .ZN(new_n1277_));
  AOI21_X1   g01019(.A1(new_n1277_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1278_));
  XOR2_X1    g01020(.A1(new_n1024_), .A2(new_n1278_), .Z(new_n1279_));
  AOI21_X1   g01021(.A1(new_n1275_), .A2(new_n1274_), .B(new_n1279_), .ZN(new_n1280_));
  NAND2_X1   g01022(.A1(new_n1275_), .A2(new_n1274_), .ZN(new_n1281_));
  INV_X1     g01023(.I(new_n1279_), .ZN(new_n1282_));
  NOR2_X1    g01024(.A1(new_n1281_), .A2(new_n1282_), .ZN(new_n1283_));
  NOR2_X1    g01025(.A1(new_n1283_), .A2(new_n1280_), .ZN(new_n1284_));
  NOR2_X1    g01026(.A1(\b[16] ), .A2(\b[17] ), .ZN(new_n1285_));
  NAND2_X1   g01027(.A1(new_n1188_), .A2(new_n1285_), .ZN(new_n1286_));
  NOR2_X1    g01028(.A1(new_n1109_), .A2(new_n1189_), .ZN(new_n1287_));
  AOI22_X1   g01029(.A1(new_n1286_), .A2(\b[15] ), .B1(new_n1106_), .B2(new_n1287_), .ZN(new_n1288_));
  XNOR2_X1   g01030(.A1(\b[17] ), .A2(\b[18] ), .ZN(new_n1289_));
  NOR2_X1    g01031(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_));
  NOR3_X1    g01032(.A1(new_n1106_), .A2(\b[16] ), .A3(\b[17] ), .ZN(new_n1291_));
  INV_X1     g01033(.I(new_n1287_), .ZN(new_n1292_));
  OAI22_X1   g01034(.A1(new_n1291_), .A2(new_n1017_), .B1(new_n1188_), .B2(new_n1292_), .ZN(new_n1293_));
  INV_X1     g01035(.I(\b[18] ), .ZN(new_n1294_));
  NOR2_X1    g01036(.A1(new_n1189_), .A2(new_n1294_), .ZN(new_n1295_));
  INV_X1     g01037(.I(new_n1295_), .ZN(new_n1296_));
  NAND2_X1   g01038(.A1(new_n1189_), .A2(new_n1294_), .ZN(new_n1297_));
  AOI21_X1   g01039(.A1(new_n1296_), .A2(new_n1297_), .B(new_n1293_), .ZN(new_n1298_));
  NOR2_X1    g01040(.A1(new_n1298_), .A2(new_n1290_), .ZN(new_n1299_));
  OAI22_X1   g01041(.A1(new_n330_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n263_), .ZN(new_n1300_));
  OAI21_X1   g01042(.A1(new_n1109_), .A2(new_n289_), .B(new_n1300_), .ZN(new_n1301_));
  AOI21_X1   g01043(.A1(new_n1301_), .A2(new_n260_), .B(new_n426_), .ZN(new_n1302_));
  XOR2_X1    g01044(.A1(new_n1299_), .A2(new_n1302_), .Z(new_n1303_));
  INV_X1     g01045(.I(new_n1303_), .ZN(new_n1304_));
  XOR2_X1    g01046(.A1(new_n1284_), .A2(new_n1304_), .Z(new_n1305_));
  OR2_X2     g01047(.A1(new_n1305_), .A2(new_n1216_), .Z(new_n1306_));
  XOR2_X1    g01048(.A1(new_n1284_), .A2(new_n1303_), .Z(new_n1307_));
  OAI21_X1   g01049(.A1(new_n1215_), .A2(new_n1307_), .B(new_n1306_), .ZN(new_n1308_));
  INV_X1     g01050(.I(new_n1308_), .ZN(new_n1309_));
  INV_X1     g01051(.I(new_n1208_), .ZN(new_n1310_));
  AOI21_X1   g01052(.A1(new_n1310_), .A2(new_n1102_), .B(new_n1123_), .ZN(new_n1311_));
  OAI21_X1   g01053(.A1(new_n1310_), .A2(new_n1102_), .B(new_n1036_), .ZN(new_n1312_));
  NOR2_X1    g01054(.A1(new_n1311_), .A2(new_n1312_), .ZN(new_n1313_));
  XOR2_X1    g01055(.A1(new_n1201_), .A2(new_n1127_), .Z(new_n1314_));
  NOR2_X1    g01056(.A1(new_n1314_), .A2(new_n1130_), .ZN(new_n1315_));
  NOR2_X1    g01057(.A1(new_n1313_), .A2(new_n1315_), .ZN(new_n1316_));
  OAI21_X1   g01058(.A1(new_n1130_), .A2(new_n1314_), .B(new_n1309_), .ZN(new_n1317_));
  OAI22_X1   g01059(.A1(new_n1316_), .A2(new_n1309_), .B1(new_n1313_), .B2(new_n1317_), .ZN(\f[18] ));
  INV_X1     g01060(.I(new_n1259_), .ZN(new_n1319_));
  NAND2_X1   g01061(.A1(new_n1255_), .A2(new_n1263_), .ZN(new_n1320_));
  NAND2_X1   g01062(.A1(new_n1320_), .A2(new_n1319_), .ZN(new_n1321_));
  OAI22_X1   g01063(.A1(new_n1226_), .A2(new_n1321_), .B1(new_n1263_), .B2(new_n1255_), .ZN(new_n1322_));
  INV_X1     g01064(.I(new_n1232_), .ZN(new_n1323_));
  XOR2_X1    g01065(.A1(new_n1234_), .A2(new_n1323_), .Z(new_n1324_));
  XOR2_X1    g01066(.A1(new_n1324_), .A2(new_n1228_), .Z(new_n1325_));
  NOR2_X1    g01067(.A1(new_n1325_), .A2(new_n1239_), .ZN(new_n1326_));
  NAND2_X1   g01068(.A1(new_n1242_), .A2(new_n1326_), .ZN(new_n1327_));
  AOI21_X1   g01069(.A1(new_n1327_), .A2(new_n1244_), .B(new_n1252_), .ZN(new_n1328_));
  NAND2_X1   g01070(.A1(new_n1233_), .A2(new_n1323_), .ZN(new_n1329_));
  NOR2_X1    g01071(.A1(new_n1138_), .A2(new_n1228_), .ZN(new_n1330_));
  OAI21_X1   g01072(.A1(new_n1233_), .A2(new_n1323_), .B(new_n1330_), .ZN(new_n1331_));
  INV_X1     g01073(.I(new_n1142_), .ZN(new_n1332_));
  OAI22_X1   g01074(.A1(new_n298_), .A2(new_n1055_), .B1(new_n1061_), .B2(new_n325_), .ZN(new_n1333_));
  OAI21_X1   g01075(.A1(new_n1332_), .A2(new_n280_), .B(new_n1333_), .ZN(new_n1334_));
  AOI21_X1   g01076(.A1(new_n1334_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n1335_));
  XOR2_X1    g01077(.A1(new_n1335_), .A2(new_n807_), .Z(new_n1336_));
  INV_X1     g01078(.I(new_n1336_), .ZN(new_n1337_));
  XOR2_X1    g01079(.A1(\a[18] ), .A2(\a[20] ), .Z(new_n1338_));
  XOR2_X1    g01080(.A1(\a[17] ), .A2(\a[19] ), .Z(new_n1339_));
  AND2_X2    g01081(.A1(new_n1338_), .A2(new_n1339_), .Z(new_n1340_));
  INV_X1     g01082(.I(\a[19] ), .ZN(new_n1341_));
  NOR3_X1    g01083(.A1(new_n1341_), .A2(\a[17] ), .A3(\a[18] ), .ZN(new_n1342_));
  AND3_X2    g01084(.A1(new_n1341_), .A2(\a[17] ), .A3(\a[18] ), .Z(new_n1343_));
  NOR2_X1    g01085(.A1(new_n1343_), .A2(new_n1342_), .ZN(new_n1344_));
  NOR2_X1    g01086(.A1(new_n1344_), .A2(new_n269_), .ZN(new_n1345_));
  INV_X1     g01087(.I(\a[20] ), .ZN(new_n1346_));
  NAND2_X1   g01088(.A1(new_n1339_), .A2(new_n1338_), .ZN(new_n1347_));
  OAI21_X1   g01089(.A1(new_n1347_), .A2(new_n258_), .B(new_n1346_), .ZN(new_n1348_));
  OAI21_X1   g01090(.A1(new_n1348_), .A2(new_n1345_), .B(new_n1340_), .ZN(new_n1349_));
  NOR2_X1    g01091(.A1(new_n1349_), .A2(new_n271_), .ZN(new_n1350_));
  AND2_X2    g01092(.A1(new_n1349_), .A2(new_n271_), .Z(new_n1351_));
  NOR2_X1    g01093(.A1(new_n1351_), .A2(new_n1350_), .ZN(new_n1352_));
  NAND2_X1   g01094(.A1(new_n1228_), .A2(\a[20] ), .ZN(new_n1353_));
  INV_X1     g01095(.I(new_n1353_), .ZN(new_n1354_));
  XOR2_X1    g01096(.A1(new_n1352_), .A2(new_n1354_), .Z(new_n1355_));
  XOR2_X1    g01097(.A1(new_n1355_), .A2(new_n1337_), .Z(new_n1356_));
  AOI21_X1   g01098(.A1(new_n1329_), .A2(new_n1331_), .B(new_n1356_), .ZN(new_n1357_));
  NAND2_X1   g01099(.A1(new_n1331_), .A2(new_n1329_), .ZN(new_n1358_));
  NAND2_X1   g01100(.A1(new_n1355_), .A2(new_n1336_), .ZN(new_n1359_));
  OR2_X2     g01101(.A1(new_n1355_), .A2(new_n1336_), .Z(new_n1360_));
  AOI21_X1   g01102(.A1(new_n1359_), .A2(new_n1360_), .B(new_n1358_), .ZN(new_n1361_));
  NOR2_X1    g01103(.A1(new_n1361_), .A2(new_n1357_), .ZN(new_n1362_));
  AOI22_X1   g01104(.A1(new_n1235_), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n817_), .ZN(new_n1363_));
  AOI21_X1   g01105(.A1(\b[5] ), .A2(new_n895_), .B(new_n1363_), .ZN(new_n1364_));
  OAI21_X1   g01106(.A1(new_n1364_), .A2(\a[14] ), .B(new_n817_), .ZN(new_n1365_));
  XNOR2_X1   g01107(.A1(new_n471_), .A2(new_n1365_), .ZN(new_n1366_));
  NOR2_X1    g01108(.A1(new_n1362_), .A2(new_n1366_), .ZN(new_n1367_));
  INV_X1     g01109(.I(new_n1362_), .ZN(new_n1368_));
  INV_X1     g01110(.I(new_n1366_), .ZN(new_n1369_));
  NOR2_X1    g01111(.A1(new_n1368_), .A2(new_n1369_), .ZN(new_n1370_));
  OAI21_X1   g01112(.A1(new_n1367_), .A2(new_n1370_), .B(new_n1328_), .ZN(new_n1371_));
  INV_X1     g01113(.I(new_n1328_), .ZN(new_n1372_));
  XOR2_X1    g01114(.A1(new_n1362_), .A2(new_n1366_), .Z(new_n1373_));
  NAND2_X1   g01115(.A1(new_n1372_), .A2(new_n1373_), .ZN(new_n1374_));
  NAND2_X1   g01116(.A1(new_n1374_), .A2(new_n1371_), .ZN(new_n1375_));
  INV_X1     g01117(.I(new_n1375_), .ZN(new_n1376_));
  OAI22_X1   g01118(.A1(new_n607_), .A2(new_n565_), .B1(new_n656_), .B2(new_n610_), .ZN(new_n1377_));
  OAI21_X1   g01119(.A1(new_n515_), .A2(new_n684_), .B(new_n1377_), .ZN(new_n1378_));
  AOI21_X1   g01120(.A1(new_n1378_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1379_));
  XNOR2_X1   g01121(.A1(new_n660_), .A2(new_n1379_), .ZN(new_n1380_));
  NOR2_X1    g01122(.A1(new_n1376_), .A2(new_n1380_), .ZN(new_n1381_));
  INV_X1     g01123(.I(new_n1380_), .ZN(new_n1382_));
  NOR2_X1    g01124(.A1(new_n1375_), .A2(new_n1382_), .ZN(new_n1383_));
  OAI21_X1   g01125(.A1(new_n1381_), .A2(new_n1383_), .B(new_n1322_), .ZN(new_n1384_));
  INV_X1     g01126(.I(new_n1322_), .ZN(new_n1385_));
  XOR2_X1    g01127(.A1(new_n1375_), .A2(new_n1382_), .Z(new_n1386_));
  NAND2_X1   g01128(.A1(new_n1385_), .A2(new_n1386_), .ZN(new_n1387_));
  NAND2_X1   g01129(.A1(new_n1387_), .A2(new_n1384_), .ZN(new_n1388_));
  INV_X1     g01130(.I(new_n1388_), .ZN(new_n1389_));
  OAI22_X1   g01131(.A1(new_n448_), .A2(new_n780_), .B1(new_n861_), .B2(new_n450_), .ZN(new_n1390_));
  OAI21_X1   g01132(.A1(new_n706_), .A2(new_n496_), .B(new_n1390_), .ZN(new_n1391_));
  AOI21_X1   g01133(.A1(new_n1391_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1392_));
  XNOR2_X1   g01134(.A1(new_n860_), .A2(new_n1392_), .ZN(new_n1393_));
  NOR2_X1    g01135(.A1(new_n1389_), .A2(new_n1393_), .ZN(new_n1394_));
  INV_X1     g01136(.I(new_n1394_), .ZN(new_n1395_));
  NAND2_X1   g01137(.A1(new_n1389_), .A2(new_n1393_), .ZN(new_n1396_));
  NAND2_X1   g01138(.A1(new_n1395_), .A2(new_n1396_), .ZN(new_n1397_));
  OAI21_X1   g01139(.A1(new_n1265_), .A2(new_n1262_), .B(new_n1217_), .ZN(new_n1398_));
  NOR3_X1    g01140(.A1(new_n1265_), .A2(new_n1262_), .A3(new_n1217_), .ZN(new_n1399_));
  NOR2_X1    g01141(.A1(new_n1399_), .A2(new_n1269_), .ZN(new_n1400_));
  NAND3_X1   g01142(.A1(new_n1400_), .A2(new_n1219_), .A3(new_n1220_), .ZN(new_n1401_));
  NAND2_X1   g01143(.A1(new_n1401_), .A2(new_n1398_), .ZN(new_n1402_));
  OAI22_X1   g01144(.A1(new_n1017_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1109_), .ZN(new_n1403_));
  OAI21_X1   g01145(.A1(new_n930_), .A2(new_n366_), .B(new_n1403_), .ZN(new_n1404_));
  AOI21_X1   g01146(.A1(new_n1404_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1405_));
  XOR2_X1    g01147(.A1(new_n1114_), .A2(new_n1405_), .Z(new_n1406_));
  NOR2_X1    g01148(.A1(new_n1402_), .A2(new_n1406_), .ZN(new_n1407_));
  INV_X1     g01149(.I(new_n1406_), .ZN(new_n1408_));
  AOI21_X1   g01150(.A1(new_n1401_), .A2(new_n1398_), .B(new_n1408_), .ZN(new_n1409_));
  OAI21_X1   g01151(.A1(new_n1407_), .A2(new_n1409_), .B(new_n1397_), .ZN(new_n1410_));
  INV_X1     g01152(.I(new_n1397_), .ZN(new_n1411_));
  AOI21_X1   g01153(.A1(new_n1401_), .A2(new_n1398_), .B(new_n1406_), .ZN(new_n1412_));
  NOR2_X1    g01154(.A1(new_n1402_), .A2(new_n1408_), .ZN(new_n1413_));
  OAI21_X1   g01155(.A1(new_n1413_), .A2(new_n1412_), .B(new_n1411_), .ZN(new_n1414_));
  XOR2_X1    g01156(.A1(new_n1281_), .A2(new_n1279_), .Z(new_n1415_));
  AOI21_X1   g01157(.A1(new_n1410_), .A2(new_n1414_), .B(new_n1415_), .ZN(new_n1416_));
  XOR2_X1    g01158(.A1(new_n1416_), .A2(new_n1280_), .Z(new_n1417_));
  XOR2_X1    g01159(.A1(new_n1417_), .A2(new_n1215_), .Z(new_n1418_));
  XNOR2_X1   g01160(.A1(\b[17] ), .A2(\b[19] ), .ZN(new_n1419_));
  NOR2_X1    g01161(.A1(new_n1419_), .A2(new_n1289_), .ZN(new_n1420_));
  XOR2_X1    g01162(.A1(new_n1293_), .A2(new_n1420_), .Z(new_n1421_));
  NAND2_X1   g01163(.A1(new_n286_), .A2(\b[18] ), .ZN(new_n1422_));
  AOI22_X1   g01164(.A1(new_n304_), .A2(\b[17] ), .B1(new_n262_), .B2(\b[19] ), .ZN(new_n1423_));
  AOI21_X1   g01165(.A1(new_n1422_), .A2(new_n1423_), .B(new_n426_), .ZN(new_n1424_));
  NAND2_X1   g01166(.A1(new_n1421_), .A2(new_n1424_), .ZN(new_n1425_));
  XOR2_X1    g01167(.A1(new_n1425_), .A2(new_n260_), .Z(new_n1426_));
  INV_X1     g01168(.I(new_n1426_), .ZN(new_n1427_));
  NAND2_X1   g01169(.A1(new_n1418_), .A2(new_n1427_), .ZN(new_n1428_));
  XOR2_X1    g01170(.A1(new_n1425_), .A2(\a[2] ), .Z(new_n1429_));
  OR2_X2     g01171(.A1(new_n1418_), .A2(new_n1429_), .Z(new_n1430_));
  NAND2_X1   g01172(.A1(new_n1430_), .A2(new_n1428_), .ZN(new_n1431_));
  XOR2_X1    g01173(.A1(new_n1284_), .A2(new_n1216_), .Z(new_n1432_));
  NOR2_X1    g01174(.A1(new_n1432_), .A2(new_n1304_), .ZN(new_n1433_));
  AOI21_X1   g01175(.A1(new_n1308_), .A2(new_n1433_), .B(new_n1315_), .ZN(new_n1434_));
  NOR3_X1    g01176(.A1(new_n1434_), .A2(new_n1311_), .A3(new_n1312_), .ZN(new_n1435_));
  XOR2_X1    g01177(.A1(new_n1431_), .A2(new_n1435_), .Z(\f[19] ));
  INV_X1     g01178(.I(new_n1398_), .ZN(new_n1437_));
  NAND2_X1   g01179(.A1(new_n1220_), .A2(new_n1219_), .ZN(new_n1438_));
  NOR3_X1    g01180(.A1(new_n1438_), .A2(new_n1269_), .A3(new_n1399_), .ZN(new_n1439_));
  NOR2_X1    g01181(.A1(new_n1439_), .A2(new_n1437_), .ZN(new_n1440_));
  NOR2_X1    g01182(.A1(new_n1440_), .A2(new_n1411_), .ZN(new_n1441_));
  NOR2_X1    g01183(.A1(new_n1402_), .A2(new_n1397_), .ZN(new_n1442_));
  OAI21_X1   g01184(.A1(new_n1441_), .A2(new_n1442_), .B(new_n1406_), .ZN(new_n1443_));
  NAND2_X1   g01185(.A1(new_n1410_), .A2(new_n1414_), .ZN(new_n1444_));
  AOI21_X1   g01186(.A1(new_n1444_), .A2(new_n1281_), .B(new_n1282_), .ZN(new_n1445_));
  OAI21_X1   g01187(.A1(new_n1444_), .A2(new_n1281_), .B(new_n1215_), .ZN(new_n1446_));
  NOR2_X1    g01188(.A1(new_n1445_), .A2(new_n1446_), .ZN(new_n1447_));
  INV_X1     g01189(.I(new_n1367_), .ZN(new_n1448_));
  OAI22_X1   g01190(.A1(new_n970_), .A2(new_n472_), .B1(new_n515_), .B2(new_n820_), .ZN(new_n1449_));
  OAI21_X1   g01191(.A1(new_n420_), .A2(new_n894_), .B(new_n1449_), .ZN(new_n1450_));
  AOI21_X1   g01192(.A1(new_n1450_), .A2(new_n827_), .B(new_n970_), .ZN(new_n1451_));
  XOR2_X1    g01193(.A1(new_n700_), .A2(new_n1451_), .Z(new_n1452_));
  NOR3_X1    g01194(.A1(new_n1351_), .A2(new_n1350_), .A3(new_n1353_), .ZN(new_n1453_));
  OAI21_X1   g01195(.A1(\b[1] ), .A2(new_n282_), .B(new_n1340_), .ZN(new_n1454_));
  OAI21_X1   g01196(.A1(new_n280_), .A2(new_n1344_), .B(new_n1454_), .ZN(new_n1455_));
  XOR2_X1    g01197(.A1(\a[17] ), .A2(\a[20] ), .Z(new_n1456_));
  NAND3_X1   g01198(.A1(new_n1339_), .A2(new_n1227_), .A3(new_n1456_), .ZN(new_n1457_));
  INV_X1     g01199(.I(new_n1457_), .ZN(new_n1458_));
  NAND3_X1   g01200(.A1(new_n1455_), .A2(\b[0] ), .A3(new_n1458_), .ZN(new_n1459_));
  XOR2_X1    g01201(.A1(new_n1459_), .A2(new_n1346_), .Z(new_n1460_));
  XOR2_X1    g01202(.A1(new_n1460_), .A2(new_n1453_), .Z(new_n1461_));
  NAND2_X1   g01203(.A1(new_n1358_), .A2(new_n1359_), .ZN(new_n1462_));
  NAND2_X1   g01204(.A1(new_n1462_), .A2(new_n1360_), .ZN(new_n1463_));
  OAI22_X1   g01205(.A1(new_n325_), .A2(new_n1055_), .B1(new_n1061_), .B2(new_n419_), .ZN(new_n1464_));
  OAI21_X1   g01206(.A1(new_n1332_), .A2(new_n298_), .B(new_n1464_), .ZN(new_n1465_));
  AOI21_X1   g01207(.A1(new_n378_), .A2(new_n1056_), .B(new_n1465_), .ZN(new_n1466_));
  XOR2_X1    g01208(.A1(new_n1466_), .A2(new_n1057_), .Z(new_n1467_));
  INV_X1     g01209(.I(new_n1467_), .ZN(new_n1468_));
  XOR2_X1    g01210(.A1(new_n1463_), .A2(new_n1468_), .Z(new_n1469_));
  XOR2_X1    g01211(.A1(new_n1469_), .A2(new_n1461_), .Z(new_n1470_));
  XOR2_X1    g01212(.A1(new_n1470_), .A2(new_n1452_), .Z(new_n1471_));
  NAND3_X1   g01213(.A1(new_n1471_), .A2(new_n1448_), .A3(new_n1373_), .ZN(new_n1472_));
  NOR2_X1    g01214(.A1(new_n1362_), .A2(new_n1366_), .ZN(new_n1473_));
  INV_X1     g01215(.I(new_n1473_), .ZN(new_n1474_));
  AOI21_X1   g01216(.A1(new_n1472_), .A2(new_n1474_), .B(new_n1328_), .ZN(new_n1475_));
  NAND3_X1   g01217(.A1(new_n1472_), .A2(new_n1328_), .A3(new_n1474_), .ZN(new_n1476_));
  INV_X1     g01218(.I(new_n1476_), .ZN(new_n1477_));
  OAI22_X1   g01219(.A1(new_n607_), .A2(new_n656_), .B1(new_n706_), .B2(new_n610_), .ZN(new_n1478_));
  OAI21_X1   g01220(.A1(new_n565_), .A2(new_n684_), .B(new_n1478_), .ZN(new_n1479_));
  AOI21_X1   g01221(.A1(new_n1479_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1480_));
  XNOR2_X1   g01222(.A1(new_n710_), .A2(new_n1480_), .ZN(new_n1481_));
  INV_X1     g01223(.I(new_n1481_), .ZN(new_n1482_));
  OAI21_X1   g01224(.A1(new_n1477_), .A2(new_n1475_), .B(new_n1482_), .ZN(new_n1483_));
  INV_X1     g01225(.I(new_n1475_), .ZN(new_n1484_));
  NAND3_X1   g01226(.A1(new_n1484_), .A2(new_n1476_), .A3(new_n1481_), .ZN(new_n1485_));
  NAND2_X1   g01227(.A1(new_n1485_), .A2(new_n1483_), .ZN(new_n1486_));
  NAND2_X1   g01228(.A1(new_n1486_), .A2(new_n1386_), .ZN(new_n1487_));
  NOR2_X1    g01229(.A1(new_n1487_), .A2(new_n1381_), .ZN(new_n1488_));
  NOR2_X1    g01230(.A1(new_n1376_), .A2(new_n1380_), .ZN(new_n1489_));
  OAI21_X1   g01231(.A1(new_n1488_), .A2(new_n1489_), .B(new_n1385_), .ZN(new_n1490_));
  INV_X1     g01232(.I(new_n1490_), .ZN(new_n1491_));
  NOR3_X1    g01233(.A1(new_n1488_), .A2(new_n1385_), .A3(new_n1489_), .ZN(new_n1492_));
  OAI22_X1   g01234(.A1(new_n448_), .A2(new_n861_), .B1(new_n930_), .B2(new_n450_), .ZN(new_n1493_));
  OAI21_X1   g01235(.A1(new_n780_), .A2(new_n496_), .B(new_n1493_), .ZN(new_n1494_));
  AOI21_X1   g01236(.A1(new_n1494_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1495_));
  XNOR2_X1   g01237(.A1(new_n937_), .A2(new_n1495_), .ZN(new_n1496_));
  NOR3_X1    g01238(.A1(new_n1491_), .A2(new_n1492_), .A3(new_n1496_), .ZN(new_n1497_));
  INV_X1     g01239(.I(new_n1492_), .ZN(new_n1498_));
  INV_X1     g01240(.I(new_n1496_), .ZN(new_n1499_));
  AOI21_X1   g01241(.A1(new_n1498_), .A2(new_n1490_), .B(new_n1499_), .ZN(new_n1500_));
  OR2_X2     g01242(.A1(new_n1500_), .A2(new_n1497_), .Z(new_n1501_));
  XNOR2_X1   g01243(.A1(new_n1388_), .A2(new_n1393_), .ZN(new_n1502_));
  NAND3_X1   g01244(.A1(new_n1501_), .A2(new_n1395_), .A3(new_n1502_), .ZN(new_n1503_));
  INV_X1     g01245(.I(new_n1503_), .ZN(new_n1504_));
  NOR2_X1    g01246(.A1(new_n1389_), .A2(new_n1393_), .ZN(new_n1506_));
  OAI21_X1   g01247(.A1(new_n1504_), .A2(new_n1506_), .B(new_n1440_), .ZN(new_n1507_));
  INV_X1     g01248(.I(new_n1506_), .ZN(new_n1508_));
  NAND3_X1   g01249(.A1(new_n1503_), .A2(new_n1402_), .A3(new_n1508_), .ZN(new_n1509_));
  NAND2_X1   g01250(.A1(new_n1507_), .A2(new_n1509_), .ZN(new_n1510_));
  OAI22_X1   g01251(.A1(new_n1109_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1189_), .ZN(new_n1511_));
  OAI21_X1   g01252(.A1(new_n1017_), .A2(new_n366_), .B(new_n1511_), .ZN(new_n1512_));
  AOI21_X1   g01253(.A1(new_n1512_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1513_));
  XNOR2_X1   g01254(.A1(new_n1196_), .A2(new_n1513_), .ZN(new_n1514_));
  XNOR2_X1   g01255(.A1(new_n1510_), .A2(new_n1514_), .ZN(new_n1515_));
  NOR2_X1    g01256(.A1(\b[18] ), .A2(\b[19] ), .ZN(new_n1516_));
  AOI21_X1   g01257(.A1(new_n1288_), .A2(new_n1516_), .B(new_n1189_), .ZN(new_n1517_));
  INV_X1     g01258(.I(\b[19] ), .ZN(new_n1518_));
  NOR2_X1    g01259(.A1(new_n1294_), .A2(new_n1518_), .ZN(new_n1519_));
  INV_X1     g01260(.I(new_n1519_), .ZN(new_n1520_));
  NOR2_X1    g01261(.A1(new_n1288_), .A2(new_n1520_), .ZN(new_n1521_));
  NOR2_X1    g01262(.A1(new_n1517_), .A2(new_n1521_), .ZN(new_n1522_));
  XNOR2_X1   g01263(.A1(\b[19] ), .A2(\b[20] ), .ZN(new_n1523_));
  NOR2_X1    g01264(.A1(new_n1522_), .A2(new_n1523_), .ZN(new_n1524_));
  INV_X1     g01265(.I(\b[20] ), .ZN(new_n1525_));
  NOR2_X1    g01266(.A1(new_n1518_), .A2(new_n1525_), .ZN(new_n1526_));
  INV_X1     g01267(.I(new_n1526_), .ZN(new_n1527_));
  NAND2_X1   g01268(.A1(new_n1518_), .A2(new_n1525_), .ZN(new_n1528_));
  NAND2_X1   g01269(.A1(new_n1527_), .A2(new_n1528_), .ZN(new_n1529_));
  AOI21_X1   g01270(.A1(new_n1522_), .A2(new_n1529_), .B(new_n1524_), .ZN(new_n1530_));
  OAI22_X1   g01271(.A1(new_n330_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n263_), .ZN(new_n1531_));
  OAI21_X1   g01272(.A1(new_n1294_), .A2(new_n289_), .B(new_n1531_), .ZN(new_n1532_));
  AOI21_X1   g01273(.A1(new_n1532_), .A2(new_n260_), .B(new_n426_), .ZN(new_n1533_));
  XOR2_X1    g01274(.A1(new_n1530_), .A2(new_n1533_), .Z(new_n1534_));
  INV_X1     g01275(.I(new_n1534_), .ZN(new_n1535_));
  NAND2_X1   g01276(.A1(new_n1515_), .A2(new_n1535_), .ZN(new_n1536_));
  OR2_X2     g01277(.A1(new_n1536_), .A2(new_n1447_), .Z(new_n1537_));
  NAND2_X1   g01278(.A1(new_n1536_), .A2(new_n1447_), .ZN(new_n1538_));
  NAND2_X1   g01279(.A1(new_n1537_), .A2(new_n1538_), .ZN(new_n1539_));
  NAND2_X1   g01280(.A1(new_n1539_), .A2(new_n1443_), .ZN(new_n1540_));
  INV_X1     g01281(.I(new_n1443_), .ZN(new_n1541_));
  NAND3_X1   g01282(.A1(new_n1537_), .A2(new_n1541_), .A3(new_n1538_), .ZN(new_n1542_));
  NAND3_X1   g01283(.A1(new_n1540_), .A2(new_n1428_), .A3(new_n1542_), .ZN(new_n1543_));
  NAND2_X1   g01284(.A1(new_n1543_), .A2(new_n1435_), .ZN(new_n1544_));
  XNOR2_X1   g01285(.A1(new_n1544_), .A2(new_n1431_), .ZN(\f[20] ));
  OAI21_X1   g01286(.A1(new_n1500_), .A2(new_n1497_), .B(new_n1388_), .ZN(new_n1546_));
  NAND2_X1   g01287(.A1(new_n1546_), .A2(new_n1393_), .ZN(new_n1547_));
  NOR3_X1    g01288(.A1(new_n1500_), .A2(new_n1497_), .A3(new_n1388_), .ZN(new_n1548_));
  NOR2_X1    g01289(.A1(new_n1440_), .A2(new_n1548_), .ZN(new_n1549_));
  AOI21_X1   g01290(.A1(new_n1484_), .A2(new_n1476_), .B(new_n1482_), .ZN(new_n1550_));
  AOI21_X1   g01291(.A1(new_n1486_), .A2(new_n1375_), .B(new_n1382_), .ZN(new_n1551_));
  OAI21_X1   g01292(.A1(new_n1486_), .A2(new_n1375_), .B(new_n1322_), .ZN(new_n1552_));
  NOR2_X1    g01293(.A1(new_n1551_), .A2(new_n1552_), .ZN(new_n1553_));
  INV_X1     g01294(.I(new_n1553_), .ZN(new_n1554_));
  XOR2_X1    g01295(.A1(new_n1463_), .A2(new_n1461_), .Z(new_n1555_));
  XOR2_X1    g01296(.A1(new_n1555_), .A2(new_n1468_), .Z(new_n1556_));
  NOR2_X1    g01297(.A1(new_n1556_), .A2(new_n1452_), .ZN(new_n1557_));
  AOI21_X1   g01298(.A1(new_n1471_), .A2(new_n1368_), .B(new_n1369_), .ZN(new_n1558_));
  OAI21_X1   g01299(.A1(new_n1471_), .A2(new_n1368_), .B(new_n1328_), .ZN(new_n1559_));
  NOR2_X1    g01300(.A1(new_n1558_), .A2(new_n1559_), .ZN(new_n1560_));
  XOR2_X1    g01301(.A1(\a[20] ), .A2(\a[21] ), .Z(new_n1561_));
  NAND2_X1   g01302(.A1(new_n1561_), .A2(\b[0] ), .ZN(new_n1562_));
  INV_X1     g01303(.I(new_n1562_), .ZN(new_n1563_));
  OAI22_X1   g01304(.A1(new_n1347_), .A2(new_n280_), .B1(new_n1344_), .B2(new_n298_), .ZN(new_n1564_));
  AOI21_X1   g01305(.A1(\b[1] ), .A2(new_n1458_), .B(new_n1564_), .ZN(new_n1565_));
  NOR3_X1    g01306(.A1(new_n1565_), .A2(new_n403_), .A3(new_n1347_), .ZN(new_n1566_));
  XOR2_X1    g01307(.A1(new_n1566_), .A2(\a[20] ), .Z(new_n1567_));
  INV_X1     g01308(.I(new_n1453_), .ZN(new_n1568_));
  NOR2_X1    g01309(.A1(new_n1460_), .A2(new_n1568_), .ZN(new_n1569_));
  INV_X1     g01310(.I(new_n1061_), .ZN(new_n1570_));
  AOI22_X1   g01311(.A1(new_n1056_), .A2(\b[5] ), .B1(new_n1570_), .B2(\b[6] ), .ZN(new_n1571_));
  AOI21_X1   g01312(.A1(\b[4] ), .A2(new_n1142_), .B(new_n1571_), .ZN(new_n1572_));
  OAI21_X1   g01313(.A1(new_n1572_), .A2(\a[17] ), .B(new_n1056_), .ZN(new_n1573_));
  XOR2_X1    g01314(.A1(new_n556_), .A2(new_n1573_), .Z(new_n1574_));
  XNOR2_X1   g01315(.A1(new_n1569_), .A2(new_n1574_), .ZN(new_n1575_));
  XOR2_X1    g01316(.A1(new_n1575_), .A2(new_n1567_), .Z(new_n1576_));
  XOR2_X1    g01317(.A1(new_n1576_), .A2(new_n1563_), .Z(new_n1577_));
  NOR2_X1    g01318(.A1(new_n1461_), .A2(new_n1468_), .ZN(new_n1578_));
  INV_X1     g01319(.I(new_n1578_), .ZN(new_n1579_));
  XOR2_X1    g01320(.A1(new_n1453_), .A2(new_n1466_), .Z(new_n1580_));
  XOR2_X1    g01321(.A1(new_n1580_), .A2(new_n1460_), .Z(new_n1581_));
  XOR2_X1    g01322(.A1(new_n1581_), .A2(\a[17] ), .Z(new_n1582_));
  AOI21_X1   g01323(.A1(new_n1582_), .A2(new_n1355_), .B(new_n1337_), .ZN(new_n1583_));
  OAI21_X1   g01324(.A1(new_n1582_), .A2(new_n1355_), .B(new_n1358_), .ZN(new_n1584_));
  NOR2_X1    g01325(.A1(new_n1583_), .A2(new_n1584_), .ZN(new_n1585_));
  INV_X1     g01326(.I(new_n1585_), .ZN(new_n1586_));
  AOI21_X1   g01327(.A1(new_n1586_), .A2(new_n1579_), .B(new_n1577_), .ZN(new_n1587_));
  AND3_X2    g01328(.A1(new_n1586_), .A2(new_n1577_), .A3(new_n1579_), .Z(new_n1588_));
  NOR2_X1    g01329(.A1(new_n1588_), .A2(new_n1587_), .ZN(new_n1589_));
  OAI22_X1   g01330(.A1(new_n970_), .A2(new_n515_), .B1(new_n565_), .B2(new_n820_), .ZN(new_n1590_));
  OAI21_X1   g01331(.A1(new_n472_), .A2(new_n894_), .B(new_n1590_), .ZN(new_n1591_));
  AOI21_X1   g01332(.A1(new_n1591_), .A2(new_n827_), .B(new_n970_), .ZN(new_n1592_));
  XOR2_X1    g01333(.A1(new_n759_), .A2(new_n1592_), .Z(new_n1593_));
  NOR2_X1    g01334(.A1(new_n1589_), .A2(new_n1593_), .ZN(new_n1594_));
  XOR2_X1    g01335(.A1(new_n1560_), .A2(new_n1594_), .Z(new_n1595_));
  XOR2_X1    g01336(.A1(new_n1595_), .A2(new_n1557_), .Z(new_n1596_));
  OAI22_X1   g01337(.A1(new_n607_), .A2(new_n706_), .B1(new_n780_), .B2(new_n610_), .ZN(new_n1597_));
  OAI21_X1   g01338(.A1(new_n656_), .A2(new_n684_), .B(new_n1597_), .ZN(new_n1598_));
  AOI21_X1   g01339(.A1(new_n1598_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1599_));
  XOR2_X1    g01340(.A1(new_n785_), .A2(new_n1599_), .Z(new_n1600_));
  INV_X1     g01341(.I(new_n1600_), .ZN(new_n1601_));
  NAND3_X1   g01342(.A1(new_n1554_), .A2(new_n1596_), .A3(new_n1601_), .ZN(new_n1602_));
  NAND2_X1   g01343(.A1(new_n1596_), .A2(new_n1601_), .ZN(new_n1603_));
  NAND2_X1   g01344(.A1(new_n1603_), .A2(new_n1553_), .ZN(new_n1604_));
  AOI21_X1   g01345(.A1(new_n1602_), .A2(new_n1604_), .B(new_n1550_), .ZN(new_n1605_));
  INV_X1     g01346(.I(new_n1605_), .ZN(new_n1606_));
  NAND3_X1   g01347(.A1(new_n1602_), .A2(new_n1604_), .A3(new_n1550_), .ZN(new_n1607_));
  NAND2_X1   g01348(.A1(new_n1606_), .A2(new_n1607_), .ZN(new_n1608_));
  OAI22_X1   g01349(.A1(new_n448_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n450_), .ZN(new_n1609_));
  OAI21_X1   g01350(.A1(new_n861_), .A2(new_n496_), .B(new_n1609_), .ZN(new_n1610_));
  AOI21_X1   g01351(.A1(new_n1610_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1611_));
  XOR2_X1    g01352(.A1(new_n1024_), .A2(new_n1611_), .Z(new_n1612_));
  INV_X1     g01353(.I(new_n1612_), .ZN(new_n1613_));
  NAND2_X1   g01354(.A1(new_n1608_), .A2(new_n1613_), .ZN(new_n1614_));
  AOI21_X1   g01355(.A1(new_n1547_), .A2(new_n1549_), .B(new_n1614_), .ZN(new_n1615_));
  INV_X1     g01356(.I(new_n1615_), .ZN(new_n1616_));
  NAND3_X1   g01357(.A1(new_n1614_), .A2(new_n1547_), .A3(new_n1549_), .ZN(new_n1617_));
  AOI21_X1   g01358(.A1(new_n1616_), .A2(new_n1617_), .B(new_n1500_), .ZN(new_n1618_));
  INV_X1     g01359(.I(new_n1500_), .ZN(new_n1619_));
  INV_X1     g01360(.I(new_n1617_), .ZN(new_n1620_));
  NOR3_X1    g01361(.A1(new_n1620_), .A2(new_n1615_), .A3(new_n1619_), .ZN(new_n1621_));
  NOR2_X1    g01362(.A1(new_n1618_), .A2(new_n1621_), .ZN(new_n1622_));
  OAI22_X1   g01363(.A1(new_n1189_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1294_), .ZN(new_n1623_));
  OAI21_X1   g01364(.A1(new_n1109_), .A2(new_n366_), .B(new_n1623_), .ZN(new_n1624_));
  AOI21_X1   g01365(.A1(new_n1624_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1625_));
  XOR2_X1    g01366(.A1(new_n1299_), .A2(new_n1625_), .Z(new_n1626_));
  INV_X1     g01367(.I(new_n1626_), .ZN(new_n1627_));
  XOR2_X1    g01368(.A1(new_n1622_), .A2(new_n1627_), .Z(new_n1628_));
  AOI21_X1   g01369(.A1(new_n1507_), .A2(new_n1509_), .B(new_n1443_), .ZN(new_n1629_));
  NAND3_X1   g01370(.A1(new_n1507_), .A2(new_n1443_), .A3(new_n1509_), .ZN(new_n1630_));
  NOR3_X1    g01371(.A1(new_n1445_), .A2(new_n1446_), .A3(new_n1514_), .ZN(new_n1631_));
  AOI21_X1   g01372(.A1(new_n1631_), .A2(new_n1630_), .B(new_n1629_), .ZN(new_n1632_));
  INV_X1     g01373(.I(new_n1523_), .ZN(new_n1633_));
  INV_X1     g01374(.I(\b[21] ), .ZN(new_n1634_));
  NOR2_X1    g01375(.A1(new_n1634_), .A2(\b[19] ), .ZN(new_n1635_));
  NOR2_X1    g01376(.A1(new_n1518_), .A2(\b[21] ), .ZN(new_n1636_));
  OAI21_X1   g01377(.A1(new_n1635_), .A2(new_n1636_), .B(new_n1633_), .ZN(new_n1637_));
  XOR2_X1    g01378(.A1(new_n1522_), .A2(new_n1637_), .Z(new_n1638_));
  NAND2_X1   g01379(.A1(new_n286_), .A2(\b[20] ), .ZN(new_n1639_));
  AOI22_X1   g01380(.A1(new_n304_), .A2(\b[19] ), .B1(new_n262_), .B2(\b[21] ), .ZN(new_n1640_));
  AOI21_X1   g01381(.A1(new_n1639_), .A2(new_n1640_), .B(new_n426_), .ZN(new_n1641_));
  NAND2_X1   g01382(.A1(new_n1638_), .A2(new_n1641_), .ZN(new_n1642_));
  XOR2_X1    g01383(.A1(new_n1642_), .A2(\a[2] ), .Z(new_n1643_));
  XOR2_X1    g01384(.A1(new_n1632_), .A2(new_n1643_), .Z(new_n1644_));
  NOR2_X1    g01385(.A1(new_n1644_), .A2(new_n1628_), .ZN(new_n1645_));
  INV_X1     g01386(.I(new_n1628_), .ZN(new_n1646_));
  INV_X1     g01387(.I(new_n1643_), .ZN(new_n1647_));
  XOR2_X1    g01388(.A1(new_n1632_), .A2(new_n1647_), .Z(new_n1648_));
  NOR2_X1    g01389(.A1(new_n1646_), .A2(new_n1648_), .ZN(new_n1649_));
  NOR2_X1    g01390(.A1(new_n1649_), .A2(new_n1645_), .ZN(new_n1650_));
  AOI21_X1   g01391(.A1(new_n1540_), .A2(new_n1542_), .B(new_n1428_), .ZN(new_n1651_));
  OAI21_X1   g01392(.A1(new_n1651_), .A2(new_n1435_), .B(new_n1431_), .ZN(new_n1652_));
  INV_X1     g01393(.I(new_n1652_), .ZN(new_n1653_));
  NOR2_X1    g01394(.A1(new_n1447_), .A2(new_n1541_), .ZN(new_n1654_));
  AND2_X2    g01395(.A1(new_n1515_), .A2(new_n1654_), .Z(new_n1655_));
  NOR2_X1    g01396(.A1(new_n1515_), .A2(new_n1654_), .ZN(new_n1656_));
  NOR3_X1    g01397(.A1(new_n1655_), .A2(new_n1535_), .A3(new_n1656_), .ZN(new_n1657_));
  NOR2_X1    g01398(.A1(new_n1653_), .A2(new_n1657_), .ZN(new_n1658_));
  INV_X1     g01399(.I(new_n1657_), .ZN(new_n1659_));
  NAND2_X1   g01400(.A1(new_n1650_), .A2(new_n1659_), .ZN(new_n1660_));
  OAI22_X1   g01401(.A1(new_n1658_), .A2(new_n1650_), .B1(new_n1653_), .B2(new_n1660_), .ZN(\f[21] ));
  INV_X1     g01402(.I(new_n1650_), .ZN(new_n1662_));
  INV_X1     g01403(.I(new_n1632_), .ZN(new_n1663_));
  NAND2_X1   g01404(.A1(new_n1628_), .A2(new_n1663_), .ZN(new_n1664_));
  NAND2_X1   g01405(.A1(new_n1646_), .A2(new_n1632_), .ZN(new_n1665_));
  AOI21_X1   g01406(.A1(new_n1665_), .A2(new_n1664_), .B(new_n1647_), .ZN(new_n1666_));
  AOI21_X1   g01407(.A1(new_n1662_), .A2(new_n1666_), .B(new_n1657_), .ZN(new_n1667_));
  NOR2_X1    g01408(.A1(new_n1652_), .A2(new_n1667_), .ZN(new_n1668_));
  NOR2_X1    g01409(.A1(new_n1622_), .A2(new_n1626_), .ZN(new_n1669_));
  INV_X1     g01410(.I(new_n1607_), .ZN(new_n1670_));
  NOR2_X1    g01411(.A1(new_n1670_), .A2(new_n1605_), .ZN(new_n1671_));
  NOR2_X1    g01412(.A1(new_n1671_), .A2(new_n1619_), .ZN(new_n1672_));
  INV_X1     g01413(.I(new_n1672_), .ZN(new_n1673_));
  NAND2_X1   g01414(.A1(new_n1671_), .A2(new_n1619_), .ZN(new_n1674_));
  NAND4_X1   g01415(.A1(new_n1674_), .A2(new_n1547_), .A3(new_n1549_), .A4(new_n1613_), .ZN(new_n1675_));
  XNOR2_X1   g01416(.A1(new_n1560_), .A2(new_n1594_), .ZN(new_n1676_));
  NOR2_X1    g01417(.A1(new_n1676_), .A2(new_n1557_), .ZN(new_n1677_));
  INV_X1     g01418(.I(new_n1557_), .ZN(new_n1678_));
  NOR2_X1    g01419(.A1(new_n1595_), .A2(new_n1678_), .ZN(new_n1679_));
  NOR3_X1    g01420(.A1(new_n1677_), .A2(new_n1679_), .A3(new_n1550_), .ZN(new_n1680_));
  NOR2_X1    g01421(.A1(new_n1680_), .A2(new_n1600_), .ZN(new_n1681_));
  AOI22_X1   g01422(.A1(new_n1681_), .A2(new_n1553_), .B1(new_n1550_), .B2(new_n1596_), .ZN(new_n1682_));
  INV_X1     g01423(.I(new_n1589_), .ZN(new_n1683_));
  AOI21_X1   g01424(.A1(new_n1678_), .A2(new_n1589_), .B(new_n1593_), .ZN(new_n1684_));
  AOI22_X1   g01425(.A1(new_n1560_), .A2(new_n1684_), .B1(new_n1557_), .B2(new_n1683_), .ZN(new_n1685_));
  XOR2_X1    g01426(.A1(new_n1569_), .A2(new_n1567_), .Z(new_n1686_));
  XOR2_X1    g01427(.A1(new_n1686_), .A2(new_n1562_), .Z(new_n1687_));
  NOR2_X1    g01428(.A1(new_n1687_), .A2(new_n1574_), .ZN(new_n1688_));
  NAND2_X1   g01429(.A1(new_n1577_), .A2(new_n1688_), .ZN(new_n1689_));
  AOI21_X1   g01430(.A1(new_n1689_), .A2(new_n1579_), .B(new_n1586_), .ZN(new_n1690_));
  NAND2_X1   g01431(.A1(new_n1460_), .A2(new_n1567_), .ZN(new_n1691_));
  NOR2_X1    g01432(.A1(new_n1460_), .A2(new_n1567_), .ZN(new_n1692_));
  NAND2_X1   g01433(.A1(new_n1453_), .A2(new_n1563_), .ZN(new_n1693_));
  OAI21_X1   g01434(.A1(new_n1692_), .A2(new_n1693_), .B(new_n1691_), .ZN(new_n1694_));
  OAI22_X1   g01435(.A1(new_n1347_), .A2(new_n298_), .B1(new_n1344_), .B2(new_n325_), .ZN(new_n1695_));
  OAI21_X1   g01436(.A1(new_n280_), .A2(new_n1457_), .B(new_n1695_), .ZN(new_n1696_));
  AOI21_X1   g01437(.A1(new_n1696_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n1697_));
  XOR2_X1    g01438(.A1(new_n1697_), .A2(new_n807_), .Z(new_n1698_));
  INV_X1     g01439(.I(new_n1698_), .ZN(new_n1699_));
  XNOR2_X1   g01440(.A1(\a[21] ), .A2(\a[23] ), .ZN(new_n1700_));
  XNOR2_X1   g01441(.A1(\a[20] ), .A2(\a[22] ), .ZN(new_n1701_));
  NOR2_X1    g01442(.A1(new_n1701_), .A2(new_n1700_), .ZN(new_n1702_));
  INV_X1     g01443(.I(\a[22] ), .ZN(new_n1703_));
  NOR3_X1    g01444(.A1(new_n1703_), .A2(\a[20] ), .A3(\a[21] ), .ZN(new_n1704_));
  INV_X1     g01445(.I(\a[21] ), .ZN(new_n1705_));
  NOR3_X1    g01446(.A1(new_n1346_), .A2(new_n1705_), .A3(\a[22] ), .ZN(new_n1706_));
  NOR2_X1    g01447(.A1(new_n1706_), .A2(new_n1704_), .ZN(new_n1707_));
  NOR2_X1    g01448(.A1(new_n1707_), .A2(new_n269_), .ZN(new_n1708_));
  INV_X1     g01449(.I(\a[23] ), .ZN(new_n1709_));
  XOR2_X1    g01450(.A1(\a[21] ), .A2(\a[23] ), .Z(new_n1710_));
  XOR2_X1    g01451(.A1(\a[20] ), .A2(\a[22] ), .Z(new_n1711_));
  NAND2_X1   g01452(.A1(new_n1711_), .A2(new_n1710_), .ZN(new_n1712_));
  OAI21_X1   g01453(.A1(new_n1712_), .A2(new_n258_), .B(new_n1709_), .ZN(new_n1713_));
  OAI21_X1   g01454(.A1(new_n1713_), .A2(new_n1708_), .B(new_n1702_), .ZN(new_n1714_));
  OR2_X2     g01455(.A1(new_n1714_), .A2(new_n271_), .Z(new_n1715_));
  NAND2_X1   g01456(.A1(new_n1714_), .A2(new_n271_), .ZN(new_n1716_));
  NAND2_X1   g01457(.A1(new_n1715_), .A2(new_n1716_), .ZN(new_n1717_));
  NOR2_X1    g01458(.A1(new_n1563_), .A2(new_n1709_), .ZN(new_n1718_));
  XOR2_X1    g01459(.A1(new_n1717_), .A2(new_n1718_), .Z(new_n1719_));
  XOR2_X1    g01460(.A1(new_n1719_), .A2(new_n1699_), .Z(new_n1720_));
  NAND2_X1   g01461(.A1(new_n1720_), .A2(new_n1694_), .ZN(new_n1721_));
  INV_X1     g01462(.I(new_n1694_), .ZN(new_n1722_));
  OR2_X2     g01463(.A1(new_n1719_), .A2(new_n1699_), .Z(new_n1723_));
  NAND2_X1   g01464(.A1(new_n1719_), .A2(new_n1699_), .ZN(new_n1724_));
  NAND2_X1   g01465(.A1(new_n1723_), .A2(new_n1724_), .ZN(new_n1725_));
  NAND2_X1   g01466(.A1(new_n1722_), .A2(new_n1725_), .ZN(new_n1726_));
  NAND2_X1   g01467(.A1(new_n1726_), .A2(new_n1721_), .ZN(new_n1727_));
  AOI22_X1   g01468(.A1(new_n1056_), .A2(\b[6] ), .B1(new_n1570_), .B2(\b[7] ), .ZN(new_n1728_));
  AOI21_X1   g01469(.A1(\b[5] ), .A2(new_n1142_), .B(new_n1728_), .ZN(new_n1729_));
  OAI21_X1   g01470(.A1(new_n1729_), .A2(\a[17] ), .B(new_n1056_), .ZN(new_n1730_));
  XNOR2_X1   g01471(.A1(new_n471_), .A2(new_n1730_), .ZN(new_n1731_));
  XOR2_X1    g01472(.A1(new_n1727_), .A2(new_n1731_), .Z(new_n1732_));
  INV_X1     g01473(.I(new_n1731_), .ZN(new_n1733_));
  XOR2_X1    g01474(.A1(new_n1727_), .A2(new_n1733_), .Z(new_n1734_));
  INV_X1     g01475(.I(new_n1734_), .ZN(new_n1735_));
  NOR2_X1    g01476(.A1(new_n1690_), .A2(new_n1735_), .ZN(new_n1736_));
  AOI21_X1   g01477(.A1(new_n1690_), .A2(new_n1732_), .B(new_n1736_), .ZN(new_n1737_));
  OAI22_X1   g01478(.A1(new_n970_), .A2(new_n565_), .B1(new_n656_), .B2(new_n820_), .ZN(new_n1738_));
  OAI21_X1   g01479(.A1(new_n515_), .A2(new_n894_), .B(new_n1738_), .ZN(new_n1739_));
  AOI21_X1   g01480(.A1(new_n1739_), .A2(new_n827_), .B(new_n970_), .ZN(new_n1740_));
  XNOR2_X1   g01481(.A1(new_n660_), .A2(new_n1740_), .ZN(new_n1741_));
  NOR2_X1    g01482(.A1(new_n1737_), .A2(new_n1741_), .ZN(new_n1742_));
  INV_X1     g01483(.I(new_n1742_), .ZN(new_n1743_));
  NAND2_X1   g01484(.A1(new_n1737_), .A2(new_n1741_), .ZN(new_n1744_));
  AOI21_X1   g01485(.A1(new_n1743_), .A2(new_n1744_), .B(new_n1685_), .ZN(new_n1745_));
  NAND2_X1   g01486(.A1(new_n1683_), .A2(new_n1557_), .ZN(new_n1746_));
  NAND2_X1   g01487(.A1(new_n1560_), .A2(new_n1684_), .ZN(new_n1747_));
  NAND2_X1   g01488(.A1(new_n1747_), .A2(new_n1746_), .ZN(new_n1748_));
  NAND2_X1   g01489(.A1(new_n1690_), .A2(new_n1732_), .ZN(new_n1749_));
  OAI21_X1   g01490(.A1(new_n1690_), .A2(new_n1735_), .B(new_n1749_), .ZN(new_n1750_));
  NOR2_X1    g01491(.A1(new_n1750_), .A2(new_n1741_), .ZN(new_n1751_));
  INV_X1     g01492(.I(new_n1741_), .ZN(new_n1752_));
  NOR2_X1    g01493(.A1(new_n1737_), .A2(new_n1752_), .ZN(new_n1753_));
  NOR2_X1    g01494(.A1(new_n1753_), .A2(new_n1751_), .ZN(new_n1754_));
  NOR2_X1    g01495(.A1(new_n1748_), .A2(new_n1754_), .ZN(new_n1755_));
  NOR2_X1    g01496(.A1(new_n1755_), .A2(new_n1745_), .ZN(new_n1756_));
  OAI22_X1   g01497(.A1(new_n607_), .A2(new_n780_), .B1(new_n861_), .B2(new_n610_), .ZN(new_n1757_));
  OAI21_X1   g01498(.A1(new_n706_), .A2(new_n684_), .B(new_n1757_), .ZN(new_n1758_));
  AOI21_X1   g01499(.A1(new_n1758_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1759_));
  XNOR2_X1   g01500(.A1(new_n860_), .A2(new_n1759_), .ZN(new_n1760_));
  XOR2_X1    g01501(.A1(new_n1756_), .A2(new_n1760_), .Z(new_n1761_));
  NOR2_X1    g01502(.A1(new_n1682_), .A2(new_n1761_), .ZN(new_n1762_));
  XOR2_X1    g01503(.A1(new_n1756_), .A2(new_n1760_), .Z(new_n1763_));
  AOI21_X1   g01504(.A1(new_n1682_), .A2(new_n1763_), .B(new_n1762_), .ZN(new_n1764_));
  OAI22_X1   g01505(.A1(new_n448_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n450_), .ZN(new_n1765_));
  OAI21_X1   g01506(.A1(new_n930_), .A2(new_n496_), .B(new_n1765_), .ZN(new_n1766_));
  AOI21_X1   g01507(.A1(new_n1766_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1767_));
  XOR2_X1    g01508(.A1(new_n1114_), .A2(new_n1767_), .Z(new_n1768_));
  NOR2_X1    g01509(.A1(new_n1764_), .A2(new_n1768_), .ZN(new_n1769_));
  NAND2_X1   g01510(.A1(new_n1764_), .A2(new_n1768_), .ZN(new_n1770_));
  INV_X1     g01511(.I(new_n1770_), .ZN(new_n1771_));
  NOR2_X1    g01512(.A1(new_n1771_), .A2(new_n1769_), .ZN(new_n1772_));
  OAI22_X1   g01513(.A1(new_n1294_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1518_), .ZN(new_n1773_));
  OAI21_X1   g01514(.A1(new_n1189_), .A2(new_n366_), .B(new_n1773_), .ZN(new_n1774_));
  AOI21_X1   g01515(.A1(new_n1774_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1775_));
  XNOR2_X1   g01516(.A1(new_n1421_), .A2(new_n1775_), .ZN(new_n1776_));
  INV_X1     g01517(.I(new_n1776_), .ZN(new_n1777_));
  NAND2_X1   g01518(.A1(new_n1772_), .A2(new_n1777_), .ZN(new_n1778_));
  OAI21_X1   g01519(.A1(new_n1771_), .A2(new_n1769_), .B(new_n1776_), .ZN(new_n1779_));
  AOI22_X1   g01520(.A1(new_n1778_), .A2(new_n1779_), .B1(new_n1675_), .B2(new_n1673_), .ZN(new_n1780_));
  NAND2_X1   g01521(.A1(new_n1675_), .A2(new_n1673_), .ZN(new_n1781_));
  INV_X1     g01522(.I(new_n1769_), .ZN(new_n1782_));
  AOI21_X1   g01523(.A1(new_n1782_), .A2(new_n1770_), .B(new_n1776_), .ZN(new_n1783_));
  NOR3_X1    g01524(.A1(new_n1771_), .A2(new_n1769_), .A3(new_n1777_), .ZN(new_n1784_));
  NOR2_X1    g01525(.A1(new_n1783_), .A2(new_n1784_), .ZN(new_n1785_));
  NOR2_X1    g01526(.A1(new_n1785_), .A2(new_n1781_), .ZN(new_n1786_));
  NOR2_X1    g01527(.A1(new_n1780_), .A2(new_n1786_), .ZN(new_n1787_));
  NOR3_X1    g01528(.A1(new_n1628_), .A2(new_n1669_), .A3(new_n1787_), .ZN(new_n1788_));
  NOR2_X1    g01529(.A1(new_n1622_), .A2(new_n1626_), .ZN(new_n1789_));
  OAI21_X1   g01530(.A1(new_n1788_), .A2(new_n1789_), .B(new_n1632_), .ZN(new_n1790_));
  NOR3_X1    g01531(.A1(new_n1788_), .A2(new_n1632_), .A3(new_n1789_), .ZN(new_n1791_));
  INV_X1     g01532(.I(new_n1791_), .ZN(new_n1792_));
  NAND2_X1   g01533(.A1(new_n1792_), .A2(new_n1790_), .ZN(new_n1793_));
  NOR2_X1    g01534(.A1(\b[20] ), .A2(\b[21] ), .ZN(new_n1794_));
  AOI21_X1   g01535(.A1(new_n1522_), .A2(new_n1794_), .B(new_n1518_), .ZN(new_n1795_));
  NOR2_X1    g01536(.A1(new_n1525_), .A2(new_n1634_), .ZN(new_n1796_));
  INV_X1     g01537(.I(new_n1796_), .ZN(new_n1797_));
  NOR2_X1    g01538(.A1(new_n1522_), .A2(new_n1797_), .ZN(new_n1798_));
  NOR2_X1    g01539(.A1(new_n1795_), .A2(new_n1798_), .ZN(new_n1799_));
  INV_X1     g01540(.I(new_n1799_), .ZN(new_n1800_));
  XNOR2_X1   g01541(.A1(\b[21] ), .A2(\b[22] ), .ZN(new_n1801_));
  INV_X1     g01542(.I(new_n1801_), .ZN(new_n1802_));
  INV_X1     g01543(.I(\b[22] ), .ZN(new_n1803_));
  NOR2_X1    g01544(.A1(new_n1634_), .A2(new_n1803_), .ZN(new_n1804_));
  INV_X1     g01545(.I(new_n1804_), .ZN(new_n1805_));
  NAND2_X1   g01546(.A1(new_n1634_), .A2(new_n1803_), .ZN(new_n1806_));
  AOI21_X1   g01547(.A1(new_n1805_), .A2(new_n1806_), .B(new_n1800_), .ZN(new_n1807_));
  AOI21_X1   g01548(.A1(new_n1800_), .A2(new_n1802_), .B(new_n1807_), .ZN(new_n1808_));
  OAI22_X1   g01549(.A1(new_n330_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n263_), .ZN(new_n1809_));
  OAI21_X1   g01550(.A1(new_n1525_), .A2(new_n289_), .B(new_n1809_), .ZN(new_n1810_));
  AOI21_X1   g01551(.A1(new_n1810_), .A2(new_n260_), .B(new_n426_), .ZN(new_n1811_));
  XOR2_X1    g01552(.A1(new_n1808_), .A2(new_n1811_), .Z(new_n1812_));
  INV_X1     g01553(.I(new_n1812_), .ZN(new_n1813_));
  NAND2_X1   g01554(.A1(new_n1793_), .A2(new_n1813_), .ZN(new_n1814_));
  INV_X1     g01555(.I(new_n1793_), .ZN(new_n1815_));
  NAND2_X1   g01556(.A1(new_n1815_), .A2(new_n1812_), .ZN(new_n1816_));
  NAND2_X1   g01557(.A1(new_n1816_), .A2(new_n1814_), .ZN(new_n1817_));
  NAND2_X1   g01558(.A1(new_n1668_), .A2(new_n1817_), .ZN(new_n1818_));
  XOR2_X1    g01559(.A1(new_n1793_), .A2(new_n1812_), .Z(new_n1819_));
  OAI21_X1   g01560(.A1(new_n1668_), .A2(new_n1819_), .B(new_n1818_), .ZN(\f[22] ));
  OAI21_X1   g01561(.A1(new_n1769_), .A2(new_n1771_), .B(new_n1781_), .ZN(new_n1821_));
  NAND2_X1   g01562(.A1(new_n1549_), .A2(new_n1547_), .ZN(new_n1822_));
  OAI21_X1   g01563(.A1(new_n1608_), .A2(new_n1500_), .B(new_n1613_), .ZN(new_n1823_));
  NOR2_X1    g01564(.A1(new_n1822_), .A2(new_n1823_), .ZN(new_n1824_));
  NOR2_X1    g01565(.A1(new_n1824_), .A2(new_n1672_), .ZN(new_n1825_));
  NAND2_X1   g01566(.A1(new_n1825_), .A2(new_n1772_), .ZN(new_n1826_));
  AOI21_X1   g01567(.A1(new_n1821_), .A2(new_n1826_), .B(new_n1777_), .ZN(new_n1827_));
  OAI21_X1   g01568(.A1(new_n1787_), .A2(new_n1622_), .B(new_n1626_), .ZN(new_n1828_));
  NOR4_X1    g01569(.A1(new_n1780_), .A2(new_n1786_), .A3(new_n1618_), .A4(new_n1621_), .ZN(new_n1829_));
  NOR2_X1    g01570(.A1(new_n1829_), .A2(new_n1632_), .ZN(new_n1830_));
  NAND2_X1   g01571(.A1(new_n1596_), .A2(new_n1550_), .ZN(new_n1831_));
  OAI21_X1   g01572(.A1(new_n1596_), .A2(new_n1550_), .B(new_n1601_), .ZN(new_n1832_));
  OAI21_X1   g01573(.A1(new_n1554_), .A2(new_n1832_), .B(new_n1831_), .ZN(new_n1833_));
  INV_X1     g01574(.I(new_n1756_), .ZN(new_n1834_));
  INV_X1     g01575(.I(new_n1760_), .ZN(new_n1835_));
  NAND2_X1   g01576(.A1(new_n1834_), .A2(new_n1835_), .ZN(new_n1836_));
  INV_X1     g01577(.I(new_n1754_), .ZN(new_n1837_));
  INV_X1     g01578(.I(new_n1690_), .ZN(new_n1838_));
  INV_X1     g01579(.I(new_n1727_), .ZN(new_n1839_));
  NOR2_X1    g01580(.A1(new_n1839_), .A2(new_n1731_), .ZN(new_n1840_));
  OAI22_X1   g01581(.A1(new_n1055_), .A2(new_n472_), .B1(new_n515_), .B2(new_n1061_), .ZN(new_n1841_));
  OAI21_X1   g01582(.A1(new_n420_), .A2(new_n1332_), .B(new_n1841_), .ZN(new_n1842_));
  AOI21_X1   g01583(.A1(new_n1842_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n1843_));
  XOR2_X1    g01584(.A1(new_n700_), .A2(new_n1843_), .Z(new_n1844_));
  INV_X1     g01585(.I(new_n1844_), .ZN(new_n1845_));
  NAND3_X1   g01586(.A1(new_n1715_), .A2(new_n1716_), .A3(new_n1718_), .ZN(new_n1846_));
  OAI21_X1   g01587(.A1(\b[1] ), .A2(new_n282_), .B(new_n1702_), .ZN(new_n1847_));
  OAI21_X1   g01588(.A1(new_n280_), .A2(new_n1707_), .B(new_n1847_), .ZN(new_n1848_));
  XOR2_X1    g01589(.A1(\a[20] ), .A2(\a[23] ), .Z(new_n1849_));
  NAND3_X1   g01590(.A1(new_n1711_), .A2(new_n1561_), .A3(new_n1849_), .ZN(new_n1850_));
  INV_X1     g01591(.I(new_n1850_), .ZN(new_n1851_));
  NAND3_X1   g01592(.A1(new_n1848_), .A2(\b[0] ), .A3(new_n1851_), .ZN(new_n1852_));
  XOR2_X1    g01593(.A1(new_n1852_), .A2(new_n1709_), .Z(new_n1853_));
  XNOR2_X1   g01594(.A1(new_n1853_), .A2(new_n1846_), .ZN(new_n1854_));
  INV_X1     g01595(.I(new_n1854_), .ZN(new_n1855_));
  NAND2_X1   g01596(.A1(new_n1694_), .A2(new_n1723_), .ZN(new_n1856_));
  NAND2_X1   g01597(.A1(new_n1856_), .A2(new_n1724_), .ZN(new_n1857_));
  OAI22_X1   g01598(.A1(new_n1347_), .A2(new_n325_), .B1(new_n1344_), .B2(new_n419_), .ZN(new_n1858_));
  OAI21_X1   g01599(.A1(new_n298_), .A2(new_n1457_), .B(new_n1858_), .ZN(new_n1859_));
  AOI21_X1   g01600(.A1(new_n378_), .A2(new_n1340_), .B(new_n1859_), .ZN(new_n1860_));
  XOR2_X1    g01601(.A1(new_n1860_), .A2(new_n1346_), .Z(new_n1861_));
  XOR2_X1    g01602(.A1(new_n1857_), .A2(new_n1861_), .Z(new_n1862_));
  NOR2_X1    g01603(.A1(new_n1862_), .A2(new_n1855_), .ZN(new_n1863_));
  INV_X1     g01604(.I(new_n1861_), .ZN(new_n1864_));
  XOR2_X1    g01605(.A1(new_n1857_), .A2(new_n1864_), .Z(new_n1865_));
  NOR2_X1    g01606(.A1(new_n1865_), .A2(new_n1854_), .ZN(new_n1866_));
  NOR2_X1    g01607(.A1(new_n1863_), .A2(new_n1866_), .ZN(new_n1867_));
  NOR2_X1    g01608(.A1(new_n1867_), .A2(new_n1845_), .ZN(new_n1868_));
  NOR3_X1    g01609(.A1(new_n1863_), .A2(new_n1866_), .A3(new_n1844_), .ZN(new_n1869_));
  NOR2_X1    g01610(.A1(new_n1868_), .A2(new_n1869_), .ZN(new_n1870_));
  NOR3_X1    g01611(.A1(new_n1870_), .A2(new_n1840_), .A3(new_n1735_), .ZN(new_n1871_));
  NOR2_X1    g01612(.A1(new_n1839_), .A2(new_n1731_), .ZN(new_n1872_));
  OAI21_X1   g01613(.A1(new_n1871_), .A2(new_n1872_), .B(new_n1838_), .ZN(new_n1873_));
  INV_X1     g01614(.I(new_n1873_), .ZN(new_n1874_));
  NOR3_X1    g01615(.A1(new_n1871_), .A2(new_n1838_), .A3(new_n1872_), .ZN(new_n1875_));
  OAI22_X1   g01616(.A1(new_n970_), .A2(new_n656_), .B1(new_n706_), .B2(new_n820_), .ZN(new_n1876_));
  OAI21_X1   g01617(.A1(new_n565_), .A2(new_n894_), .B(new_n1876_), .ZN(new_n1877_));
  AOI21_X1   g01618(.A1(new_n1877_), .A2(new_n827_), .B(new_n970_), .ZN(new_n1878_));
  XNOR2_X1   g01619(.A1(new_n710_), .A2(new_n1878_), .ZN(new_n1879_));
  INV_X1     g01620(.I(new_n1879_), .ZN(new_n1880_));
  OAI21_X1   g01621(.A1(new_n1874_), .A2(new_n1875_), .B(new_n1880_), .ZN(new_n1881_));
  OR3_X2     g01622(.A1(new_n1871_), .A2(new_n1838_), .A3(new_n1872_), .Z(new_n1882_));
  NAND3_X1   g01623(.A1(new_n1882_), .A2(new_n1873_), .A3(new_n1879_), .ZN(new_n1883_));
  NAND2_X1   g01624(.A1(new_n1881_), .A2(new_n1883_), .ZN(new_n1884_));
  NAND3_X1   g01625(.A1(new_n1884_), .A2(new_n1837_), .A3(new_n1743_), .ZN(new_n1885_));
  NOR2_X1    g01626(.A1(new_n1737_), .A2(new_n1741_), .ZN(new_n1887_));
  INV_X1     g01627(.I(new_n1887_), .ZN(new_n1888_));
  AOI21_X1   g01628(.A1(new_n1885_), .A2(new_n1888_), .B(new_n1748_), .ZN(new_n1889_));
  AOI21_X1   g01629(.A1(new_n1882_), .A2(new_n1873_), .B(new_n1879_), .ZN(new_n1890_));
  NOR3_X1    g01630(.A1(new_n1874_), .A2(new_n1875_), .A3(new_n1880_), .ZN(new_n1891_));
  OAI22_X1   g01631(.A1(new_n1891_), .A2(new_n1890_), .B1(new_n1751_), .B2(new_n1753_), .ZN(new_n1892_));
  NOR2_X1    g01632(.A1(new_n1892_), .A2(new_n1742_), .ZN(new_n1893_));
  NOR3_X1    g01633(.A1(new_n1893_), .A2(new_n1685_), .A3(new_n1887_), .ZN(new_n1894_));
  OAI22_X1   g01634(.A1(new_n607_), .A2(new_n861_), .B1(new_n930_), .B2(new_n610_), .ZN(new_n1895_));
  OAI21_X1   g01635(.A1(new_n780_), .A2(new_n684_), .B(new_n1895_), .ZN(new_n1896_));
  AOI21_X1   g01636(.A1(new_n1896_), .A2(new_n612_), .B(new_n607_), .ZN(new_n1897_));
  XNOR2_X1   g01637(.A1(new_n937_), .A2(new_n1897_), .ZN(new_n1898_));
  NOR3_X1    g01638(.A1(new_n1894_), .A2(new_n1889_), .A3(new_n1898_), .ZN(new_n1899_));
  OAI21_X1   g01639(.A1(new_n1893_), .A2(new_n1887_), .B(new_n1685_), .ZN(new_n1900_));
  NAND3_X1   g01640(.A1(new_n1885_), .A2(new_n1748_), .A3(new_n1888_), .ZN(new_n1901_));
  INV_X1     g01641(.I(new_n1898_), .ZN(new_n1902_));
  AOI21_X1   g01642(.A1(new_n1900_), .A2(new_n1901_), .B(new_n1902_), .ZN(new_n1903_));
  OR2_X2     g01643(.A1(new_n1899_), .A2(new_n1903_), .Z(new_n1904_));
  NAND3_X1   g01644(.A1(new_n1904_), .A2(new_n1836_), .A3(new_n1763_), .ZN(new_n1905_));
  NOR2_X1    g01645(.A1(new_n1756_), .A2(new_n1760_), .ZN(new_n1907_));
  INV_X1     g01646(.I(new_n1907_), .ZN(new_n1908_));
  AOI21_X1   g01647(.A1(new_n1905_), .A2(new_n1908_), .B(new_n1833_), .ZN(new_n1909_));
  INV_X1     g01648(.I(new_n1909_), .ZN(new_n1910_));
  NAND3_X1   g01649(.A1(new_n1905_), .A2(new_n1833_), .A3(new_n1908_), .ZN(new_n1911_));
  OAI22_X1   g01650(.A1(new_n448_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n450_), .ZN(new_n1912_));
  OAI21_X1   g01651(.A1(new_n1017_), .A2(new_n496_), .B(new_n1912_), .ZN(new_n1913_));
  AOI21_X1   g01652(.A1(new_n1913_), .A2(new_n452_), .B(new_n448_), .ZN(new_n1914_));
  XNOR2_X1   g01653(.A1(new_n1196_), .A2(new_n1914_), .ZN(new_n1915_));
  INV_X1     g01654(.I(new_n1915_), .ZN(new_n1916_));
  NAND3_X1   g01655(.A1(new_n1910_), .A2(new_n1911_), .A3(new_n1916_), .ZN(new_n1917_));
  INV_X1     g01656(.I(new_n1911_), .ZN(new_n1918_));
  OAI21_X1   g01657(.A1(new_n1918_), .A2(new_n1909_), .B(new_n1915_), .ZN(new_n1919_));
  NAND2_X1   g01658(.A1(new_n1917_), .A2(new_n1919_), .ZN(new_n1920_));
  XOR2_X1    g01659(.A1(new_n1764_), .A2(new_n1768_), .Z(new_n1921_));
  AND3_X2    g01660(.A1(new_n1921_), .A2(new_n1782_), .A3(new_n1920_), .Z(new_n1922_));
  NOR3_X1    g01661(.A1(new_n1918_), .A2(new_n1909_), .A3(new_n1915_), .ZN(new_n1923_));
  AOI21_X1   g01662(.A1(new_n1910_), .A2(new_n1911_), .B(new_n1916_), .ZN(new_n1924_));
  NOR2_X1    g01663(.A1(new_n1764_), .A2(new_n1768_), .ZN(new_n1925_));
  NOR2_X1    g01664(.A1(new_n1922_), .A2(new_n1925_), .ZN(new_n1926_));
  NOR2_X1    g01665(.A1(new_n1926_), .A2(new_n1781_), .ZN(new_n1927_));
  NOR3_X1    g01666(.A1(new_n1922_), .A2(new_n1825_), .A3(new_n1925_), .ZN(new_n1928_));
  NOR2_X1    g01667(.A1(new_n1927_), .A2(new_n1928_), .ZN(new_n1929_));
  OAI22_X1   g01668(.A1(new_n1518_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1525_), .ZN(new_n1930_));
  OAI21_X1   g01669(.A1(new_n1294_), .A2(new_n366_), .B(new_n1930_), .ZN(new_n1931_));
  AOI21_X1   g01670(.A1(new_n1931_), .A2(new_n334_), .B(new_n341_), .ZN(new_n1932_));
  XOR2_X1    g01671(.A1(new_n1530_), .A2(new_n1932_), .Z(new_n1933_));
  INV_X1     g01672(.I(new_n1933_), .ZN(new_n1934_));
  XOR2_X1    g01673(.A1(new_n1929_), .A2(new_n1934_), .Z(new_n1935_));
  INV_X1     g01674(.I(\b[23] ), .ZN(new_n1936_));
  NOR2_X1    g01675(.A1(new_n1936_), .A2(\b[21] ), .ZN(new_n1937_));
  NOR2_X1    g01676(.A1(new_n1634_), .A2(\b[23] ), .ZN(new_n1938_));
  OAI21_X1   g01677(.A1(new_n1937_), .A2(new_n1938_), .B(new_n1802_), .ZN(new_n1939_));
  XOR2_X1    g01678(.A1(new_n1799_), .A2(new_n1939_), .Z(new_n1940_));
  NAND2_X1   g01679(.A1(new_n286_), .A2(\b[22] ), .ZN(new_n1941_));
  AOI22_X1   g01680(.A1(new_n304_), .A2(\b[21] ), .B1(new_n262_), .B2(\b[23] ), .ZN(new_n1942_));
  AOI21_X1   g01681(.A1(new_n1941_), .A2(new_n1942_), .B(new_n426_), .ZN(new_n1943_));
  NAND2_X1   g01682(.A1(new_n1940_), .A2(new_n1943_), .ZN(new_n1944_));
  XOR2_X1    g01683(.A1(new_n1944_), .A2(\a[2] ), .Z(new_n1945_));
  INV_X1     g01684(.I(new_n1945_), .ZN(new_n1946_));
  NAND2_X1   g01685(.A1(new_n1935_), .A2(new_n1946_), .ZN(new_n1947_));
  AOI21_X1   g01686(.A1(new_n1828_), .A2(new_n1830_), .B(new_n1947_), .ZN(new_n1948_));
  NAND2_X1   g01687(.A1(new_n1830_), .A2(new_n1828_), .ZN(new_n1949_));
  AOI21_X1   g01688(.A1(new_n1935_), .A2(new_n1946_), .B(new_n1949_), .ZN(new_n1950_));
  NOR2_X1    g01689(.A1(new_n1948_), .A2(new_n1950_), .ZN(new_n1951_));
  NOR2_X1    g01690(.A1(new_n1951_), .A2(new_n1827_), .ZN(new_n1952_));
  INV_X1     g01691(.I(new_n1952_), .ZN(new_n1953_));
  NAND2_X1   g01692(.A1(new_n1951_), .A2(new_n1827_), .ZN(new_n1954_));
  AOI21_X1   g01693(.A1(new_n1953_), .A2(new_n1954_), .B(new_n1819_), .ZN(new_n1955_));
  XNOR2_X1   g01694(.A1(new_n1955_), .A2(new_n1814_), .ZN(new_n1956_));
  XOR2_X1    g01695(.A1(new_n1956_), .A2(new_n1668_), .Z(\f[23] ));
  INV_X1     g01696(.I(new_n1954_), .ZN(new_n1958_));
  OAI21_X1   g01697(.A1(new_n1958_), .A2(new_n1952_), .B(new_n1793_), .ZN(new_n1959_));
  NAND2_X1   g01698(.A1(new_n1959_), .A2(new_n1812_), .ZN(new_n1960_));
  NAND3_X1   g01699(.A1(new_n1953_), .A2(new_n1815_), .A3(new_n1954_), .ZN(new_n1961_));
  NAND3_X1   g01700(.A1(new_n1960_), .A2(new_n1668_), .A3(new_n1961_), .ZN(new_n1962_));
  INV_X1     g01701(.I(new_n1962_), .ZN(new_n1963_));
  OAI21_X1   g01702(.A1(new_n1927_), .A2(new_n1928_), .B(new_n1827_), .ZN(new_n1964_));
  NOR3_X1    g01703(.A1(new_n1927_), .A2(new_n1827_), .A3(new_n1928_), .ZN(new_n1965_));
  NAND3_X1   g01704(.A1(new_n1830_), .A2(new_n1828_), .A3(new_n1934_), .ZN(new_n1966_));
  OAI21_X1   g01705(.A1(new_n1966_), .A2(new_n1965_), .B(new_n1964_), .ZN(new_n1967_));
  INV_X1     g01706(.I(new_n1764_), .ZN(new_n1968_));
  INV_X1     g01707(.I(new_n1768_), .ZN(new_n1969_));
  AOI21_X1   g01708(.A1(new_n1920_), .A2(new_n1968_), .B(new_n1969_), .ZN(new_n1970_));
  NAND3_X1   g01709(.A1(new_n1917_), .A2(new_n1919_), .A3(new_n1764_), .ZN(new_n1971_));
  INV_X1     g01710(.I(new_n1971_), .ZN(new_n1972_));
  NOR3_X1    g01711(.A1(new_n1825_), .A2(new_n1970_), .A3(new_n1972_), .ZN(new_n1973_));
  INV_X1     g01712(.I(new_n1903_), .ZN(new_n1974_));
  OAI21_X1   g01713(.A1(new_n1899_), .A2(new_n1903_), .B(new_n1834_), .ZN(new_n1975_));
  NAND2_X1   g01714(.A1(new_n1975_), .A2(new_n1760_), .ZN(new_n1976_));
  OR3_X2     g01715(.A1(new_n1899_), .A2(new_n1903_), .A3(new_n1834_), .Z(new_n1977_));
  NAND3_X1   g01716(.A1(new_n1976_), .A2(new_n1833_), .A3(new_n1977_), .ZN(new_n1978_));
  INV_X1     g01717(.I(new_n1978_), .ZN(new_n1979_));
  OAI21_X1   g01718(.A1(new_n1874_), .A2(new_n1875_), .B(new_n1879_), .ZN(new_n1980_));
  INV_X1     g01719(.I(new_n1980_), .ZN(new_n1981_));
  OAI21_X1   g01720(.A1(new_n1891_), .A2(new_n1890_), .B(new_n1750_), .ZN(new_n1982_));
  NAND2_X1   g01721(.A1(new_n1982_), .A2(new_n1741_), .ZN(new_n1983_));
  NAND3_X1   g01722(.A1(new_n1881_), .A2(new_n1883_), .A3(new_n1737_), .ZN(new_n1984_));
  NAND3_X1   g01723(.A1(new_n1983_), .A2(new_n1748_), .A3(new_n1984_), .ZN(new_n1985_));
  XOR2_X1    g01724(.A1(new_n1857_), .A2(new_n1854_), .Z(new_n1986_));
  XOR2_X1    g01725(.A1(new_n1986_), .A2(new_n1864_), .Z(new_n1987_));
  NOR2_X1    g01726(.A1(new_n1987_), .A2(new_n1844_), .ZN(new_n1988_));
  INV_X1     g01727(.I(new_n1988_), .ZN(new_n1989_));
  OAI21_X1   g01728(.A1(new_n1870_), .A2(new_n1839_), .B(new_n1731_), .ZN(new_n1990_));
  AOI21_X1   g01729(.A1(new_n1870_), .A2(new_n1839_), .B(new_n1838_), .ZN(new_n1991_));
  XOR2_X1    g01730(.A1(\a[23] ), .A2(\a[24] ), .Z(new_n1992_));
  NAND2_X1   g01731(.A1(new_n1992_), .A2(\b[0] ), .ZN(new_n1993_));
  OAI22_X1   g01732(.A1(new_n1712_), .A2(new_n280_), .B1(new_n298_), .B2(new_n1707_), .ZN(new_n1994_));
  AOI21_X1   g01733(.A1(\b[1] ), .A2(new_n1851_), .B(new_n1994_), .ZN(new_n1995_));
  NOR3_X1    g01734(.A1(new_n1995_), .A2(new_n403_), .A3(new_n1712_), .ZN(new_n1996_));
  XOR2_X1    g01735(.A1(new_n1996_), .A2(\a[23] ), .Z(new_n1997_));
  NOR2_X1    g01736(.A1(new_n1853_), .A2(new_n1846_), .ZN(new_n1998_));
  INV_X1     g01737(.I(new_n1344_), .ZN(new_n1999_));
  AOI22_X1   g01738(.A1(\b[6] ), .A2(new_n1999_), .B1(new_n1340_), .B2(\b[5] ), .ZN(new_n2000_));
  AOI21_X1   g01739(.A1(\b[4] ), .A2(new_n1458_), .B(new_n2000_), .ZN(new_n2001_));
  OAI21_X1   g01740(.A1(new_n2001_), .A2(\a[20] ), .B(new_n1340_), .ZN(new_n2002_));
  XOR2_X1    g01741(.A1(new_n556_), .A2(new_n2002_), .Z(new_n2003_));
  XOR2_X1    g01742(.A1(new_n2003_), .A2(new_n1998_), .Z(new_n2004_));
  NOR2_X1    g01743(.A1(new_n2004_), .A2(new_n1997_), .ZN(new_n2005_));
  NAND2_X1   g01744(.A1(new_n2004_), .A2(new_n1997_), .ZN(new_n2006_));
  INV_X1     g01745(.I(new_n2006_), .ZN(new_n2007_));
  OAI21_X1   g01746(.A1(new_n2007_), .A2(new_n2005_), .B(new_n1993_), .ZN(new_n2008_));
  INV_X1     g01747(.I(new_n1993_), .ZN(new_n2009_));
  INV_X1     g01748(.I(new_n1997_), .ZN(new_n2010_));
  XNOR2_X1   g01749(.A1(new_n2003_), .A2(new_n1998_), .ZN(new_n2011_));
  NAND2_X1   g01750(.A1(new_n2011_), .A2(new_n2010_), .ZN(new_n2012_));
  NAND3_X1   g01751(.A1(new_n2012_), .A2(new_n2006_), .A3(new_n2009_), .ZN(new_n2013_));
  NOR2_X1    g01752(.A1(new_n1854_), .A2(new_n1864_), .ZN(new_n2014_));
  INV_X1     g01753(.I(new_n2014_), .ZN(new_n2015_));
  INV_X1     g01754(.I(new_n1853_), .ZN(new_n2016_));
  XOR2_X1    g01755(.A1(new_n1846_), .A2(new_n1860_), .Z(new_n2017_));
  XOR2_X1    g01756(.A1(new_n2017_), .A2(new_n2016_), .Z(new_n2018_));
  XOR2_X1    g01757(.A1(new_n2018_), .A2(new_n1346_), .Z(new_n2019_));
  OAI21_X1   g01758(.A1(new_n2019_), .A2(new_n1719_), .B(new_n1698_), .ZN(new_n2020_));
  NAND2_X1   g01759(.A1(new_n2019_), .A2(new_n1719_), .ZN(new_n2021_));
  NAND3_X1   g01760(.A1(new_n2020_), .A2(new_n2021_), .A3(new_n1694_), .ZN(new_n2022_));
  NAND2_X1   g01761(.A1(new_n2022_), .A2(new_n2015_), .ZN(new_n2023_));
  NAND3_X1   g01762(.A1(new_n2023_), .A2(new_n2008_), .A3(new_n2013_), .ZN(new_n2024_));
  NAND2_X1   g01763(.A1(new_n2008_), .A2(new_n2013_), .ZN(new_n2025_));
  NAND3_X1   g01764(.A1(new_n2022_), .A2(new_n2025_), .A3(new_n2015_), .ZN(new_n2026_));
  NAND2_X1   g01765(.A1(new_n2024_), .A2(new_n2026_), .ZN(new_n2027_));
  OAI22_X1   g01766(.A1(new_n1055_), .A2(new_n515_), .B1(new_n565_), .B2(new_n1061_), .ZN(new_n2028_));
  OAI21_X1   g01767(.A1(new_n472_), .A2(new_n1332_), .B(new_n2028_), .ZN(new_n2029_));
  AOI21_X1   g01768(.A1(new_n2029_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n2030_));
  XOR2_X1    g01769(.A1(new_n759_), .A2(new_n2030_), .Z(new_n2031_));
  INV_X1     g01770(.I(new_n2031_), .ZN(new_n2032_));
  NAND2_X1   g01771(.A1(new_n2027_), .A2(new_n2032_), .ZN(new_n2033_));
  AOI21_X1   g01772(.A1(new_n1991_), .A2(new_n1990_), .B(new_n2033_), .ZN(new_n2034_));
  NAND3_X1   g01773(.A1(new_n1991_), .A2(new_n1990_), .A3(new_n2033_), .ZN(new_n2035_));
  INV_X1     g01774(.I(new_n2035_), .ZN(new_n2036_));
  OAI21_X1   g01775(.A1(new_n2036_), .A2(new_n2034_), .B(new_n1989_), .ZN(new_n2037_));
  NAND2_X1   g01776(.A1(new_n1870_), .A2(new_n1839_), .ZN(new_n2038_));
  NAND3_X1   g01777(.A1(new_n1990_), .A2(new_n2038_), .A3(new_n1690_), .ZN(new_n2039_));
  INV_X1     g01778(.I(new_n2033_), .ZN(new_n2040_));
  NAND2_X1   g01779(.A1(new_n2039_), .A2(new_n2040_), .ZN(new_n2041_));
  NAND3_X1   g01780(.A1(new_n2041_), .A2(new_n2035_), .A3(new_n1988_), .ZN(new_n2042_));
  OAI22_X1   g01781(.A1(new_n970_), .A2(new_n706_), .B1(new_n780_), .B2(new_n820_), .ZN(new_n2043_));
  OAI21_X1   g01782(.A1(new_n656_), .A2(new_n894_), .B(new_n2043_), .ZN(new_n2044_));
  AOI21_X1   g01783(.A1(new_n2044_), .A2(new_n827_), .B(new_n970_), .ZN(new_n2045_));
  XOR2_X1    g01784(.A1(new_n785_), .A2(new_n2045_), .Z(new_n2046_));
  AOI21_X1   g01785(.A1(new_n2037_), .A2(new_n2042_), .B(new_n2046_), .ZN(new_n2047_));
  NAND2_X1   g01786(.A1(new_n1985_), .A2(new_n2047_), .ZN(new_n2048_));
  AOI21_X1   g01787(.A1(new_n1884_), .A2(new_n1750_), .B(new_n1752_), .ZN(new_n2049_));
  NAND2_X1   g01788(.A1(new_n1748_), .A2(new_n1984_), .ZN(new_n2050_));
  NOR2_X1    g01789(.A1(new_n2050_), .A2(new_n2049_), .ZN(new_n2051_));
  INV_X1     g01790(.I(new_n2047_), .ZN(new_n2052_));
  NAND2_X1   g01791(.A1(new_n2051_), .A2(new_n2052_), .ZN(new_n2053_));
  AOI21_X1   g01792(.A1(new_n2053_), .A2(new_n2048_), .B(new_n1981_), .ZN(new_n2054_));
  NOR2_X1    g01793(.A1(new_n2051_), .A2(new_n2052_), .ZN(new_n2055_));
  NOR2_X1    g01794(.A1(new_n1985_), .A2(new_n2047_), .ZN(new_n2056_));
  NOR3_X1    g01795(.A1(new_n2055_), .A2(new_n2056_), .A3(new_n1980_), .ZN(new_n2057_));
  NOR2_X1    g01796(.A1(new_n2054_), .A2(new_n2057_), .ZN(new_n2058_));
  OAI22_X1   g01797(.A1(new_n607_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n610_), .ZN(new_n2059_));
  OAI21_X1   g01798(.A1(new_n861_), .A2(new_n684_), .B(new_n2059_), .ZN(new_n2060_));
  AOI21_X1   g01799(.A1(new_n2060_), .A2(new_n612_), .B(new_n607_), .ZN(new_n2061_));
  XOR2_X1    g01800(.A1(new_n1024_), .A2(new_n2061_), .Z(new_n2062_));
  NOR3_X1    g01801(.A1(new_n1979_), .A2(new_n2058_), .A3(new_n2062_), .ZN(new_n2063_));
  OAI21_X1   g01802(.A1(new_n2055_), .A2(new_n2056_), .B(new_n1980_), .ZN(new_n2064_));
  NAND3_X1   g01803(.A1(new_n2053_), .A2(new_n2048_), .A3(new_n1981_), .ZN(new_n2065_));
  NAND2_X1   g01804(.A1(new_n2064_), .A2(new_n2065_), .ZN(new_n2066_));
  INV_X1     g01805(.I(new_n2062_), .ZN(new_n2067_));
  AOI21_X1   g01806(.A1(new_n2066_), .A2(new_n2067_), .B(new_n1978_), .ZN(new_n2068_));
  OAI21_X1   g01807(.A1(new_n2063_), .A2(new_n2068_), .B(new_n1974_), .ZN(new_n2069_));
  INV_X1     g01808(.I(new_n2069_), .ZN(new_n2070_));
  NOR3_X1    g01809(.A1(new_n2063_), .A2(new_n1974_), .A3(new_n2068_), .ZN(new_n2071_));
  NOR2_X1    g01810(.A1(new_n2070_), .A2(new_n2071_), .ZN(new_n2072_));
  OAI22_X1   g01811(.A1(new_n448_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n450_), .ZN(new_n2073_));
  OAI21_X1   g01812(.A1(new_n1109_), .A2(new_n496_), .B(new_n2073_), .ZN(new_n2074_));
  AOI21_X1   g01813(.A1(new_n2074_), .A2(new_n452_), .B(new_n448_), .ZN(new_n2075_));
  XOR2_X1    g01814(.A1(new_n1299_), .A2(new_n2075_), .Z(new_n2076_));
  NOR3_X1    g01815(.A1(new_n1973_), .A2(new_n2072_), .A3(new_n2076_), .ZN(new_n2077_));
  OAI21_X1   g01816(.A1(new_n1924_), .A2(new_n1923_), .B(new_n1968_), .ZN(new_n2078_));
  NAND2_X1   g01817(.A1(new_n2078_), .A2(new_n1768_), .ZN(new_n2079_));
  NAND3_X1   g01818(.A1(new_n2079_), .A2(new_n1781_), .A3(new_n1971_), .ZN(new_n2080_));
  NOR2_X1    g01819(.A1(new_n2072_), .A2(new_n2076_), .ZN(new_n2081_));
  NOR2_X1    g01820(.A1(new_n2080_), .A2(new_n2081_), .ZN(new_n2082_));
  OAI21_X1   g01821(.A1(new_n2077_), .A2(new_n2082_), .B(new_n1919_), .ZN(new_n2083_));
  OR3_X2     g01822(.A1(new_n2077_), .A2(new_n1919_), .A3(new_n2082_), .Z(new_n2084_));
  NAND2_X1   g01823(.A1(new_n2084_), .A2(new_n2083_), .ZN(new_n2085_));
  OAI22_X1   g01824(.A1(new_n1525_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1634_), .ZN(new_n2086_));
  OAI21_X1   g01825(.A1(new_n1518_), .A2(new_n366_), .B(new_n2086_), .ZN(new_n2087_));
  AOI21_X1   g01826(.A1(new_n2087_), .A2(new_n334_), .B(new_n341_), .ZN(new_n2088_));
  XNOR2_X1   g01827(.A1(new_n1638_), .A2(new_n2088_), .ZN(new_n2089_));
  NOR2_X1    g01828(.A1(new_n2085_), .A2(new_n2089_), .ZN(new_n2090_));
  NAND2_X1   g01829(.A1(new_n2085_), .A2(new_n2089_), .ZN(new_n2091_));
  INV_X1     g01830(.I(new_n2091_), .ZN(new_n2092_));
  NOR2_X1    g01831(.A1(new_n2092_), .A2(new_n2090_), .ZN(new_n2093_));
  NOR2_X1    g01832(.A1(\b[22] ), .A2(\b[23] ), .ZN(new_n2094_));
  AOI21_X1   g01833(.A1(new_n1799_), .A2(new_n2094_), .B(new_n1634_), .ZN(new_n2095_));
  NOR2_X1    g01834(.A1(new_n1803_), .A2(new_n1936_), .ZN(new_n2096_));
  INV_X1     g01835(.I(new_n2096_), .ZN(new_n2097_));
  NOR2_X1    g01836(.A1(new_n1799_), .A2(new_n2097_), .ZN(new_n2098_));
  NOR2_X1    g01837(.A1(new_n2095_), .A2(new_n2098_), .ZN(new_n2099_));
  XNOR2_X1   g01838(.A1(\b[23] ), .A2(\b[24] ), .ZN(new_n2100_));
  NOR2_X1    g01839(.A1(new_n2099_), .A2(new_n2100_), .ZN(new_n2101_));
  INV_X1     g01840(.I(\b[24] ), .ZN(new_n2102_));
  NOR2_X1    g01841(.A1(new_n1936_), .A2(new_n2102_), .ZN(new_n2103_));
  NOR2_X1    g01842(.A1(\b[23] ), .A2(\b[24] ), .ZN(new_n2104_));
  OR2_X2     g01843(.A1(new_n2103_), .A2(new_n2104_), .Z(new_n2105_));
  AOI21_X1   g01844(.A1(new_n2099_), .A2(new_n2105_), .B(new_n2101_), .ZN(new_n2106_));
  OAI22_X1   g01845(.A1(new_n330_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n263_), .ZN(new_n2107_));
  OAI21_X1   g01846(.A1(new_n1803_), .A2(new_n289_), .B(new_n2107_), .ZN(new_n2108_));
  AOI21_X1   g01847(.A1(new_n2108_), .A2(new_n260_), .B(new_n426_), .ZN(new_n2109_));
  XOR2_X1    g01848(.A1(new_n2106_), .A2(new_n2109_), .Z(new_n2110_));
  NOR2_X1    g01849(.A1(new_n2093_), .A2(new_n2110_), .ZN(new_n2111_));
  INV_X1     g01850(.I(new_n2093_), .ZN(new_n2112_));
  INV_X1     g01851(.I(new_n2110_), .ZN(new_n2113_));
  NOR2_X1    g01852(.A1(new_n2112_), .A2(new_n2113_), .ZN(new_n2114_));
  OAI21_X1   g01853(.A1(new_n2114_), .A2(new_n2111_), .B(new_n1967_), .ZN(new_n2115_));
  INV_X1     g01854(.I(new_n1967_), .ZN(new_n2116_));
  NOR2_X1    g01855(.A1(new_n2112_), .A2(new_n2110_), .ZN(new_n2117_));
  NOR2_X1    g01856(.A1(new_n2093_), .A2(new_n2113_), .ZN(new_n2118_));
  OAI21_X1   g01857(.A1(new_n2117_), .A2(new_n2118_), .B(new_n2116_), .ZN(new_n2119_));
  NAND2_X1   g01858(.A1(new_n2115_), .A2(new_n2119_), .ZN(new_n2120_));
  NOR2_X1    g01859(.A1(new_n1947_), .A2(new_n1827_), .ZN(new_n2121_));
  INV_X1     g01860(.I(new_n2121_), .ZN(new_n2122_));
  NAND2_X1   g01861(.A1(new_n1947_), .A2(new_n1827_), .ZN(new_n2123_));
  AOI21_X1   g01862(.A1(new_n2122_), .A2(new_n2123_), .B(new_n1949_), .ZN(new_n2124_));
  OAI21_X1   g01863(.A1(new_n1963_), .A2(new_n2124_), .B(new_n2120_), .ZN(new_n2125_));
  OR2_X2     g01864(.A1(new_n2120_), .A2(new_n2124_), .Z(new_n2126_));
  OAI21_X1   g01865(.A1(new_n1963_), .A2(new_n2126_), .B(new_n2125_), .ZN(\f[24] ));
  NAND2_X1   g01866(.A1(new_n2112_), .A2(new_n2116_), .ZN(new_n2128_));
  NAND2_X1   g01867(.A1(new_n2093_), .A2(new_n1967_), .ZN(new_n2129_));
  AOI21_X1   g01868(.A1(new_n2128_), .A2(new_n2129_), .B(new_n2113_), .ZN(new_n2130_));
  AOI21_X1   g01869(.A1(new_n2120_), .A2(new_n2130_), .B(new_n2124_), .ZN(new_n2131_));
  NOR2_X1    g01870(.A1(new_n1962_), .A2(new_n2131_), .ZN(new_n2132_));
  INV_X1     g01871(.I(new_n2085_), .ZN(new_n2133_));
  INV_X1     g01872(.I(new_n2071_), .ZN(new_n2134_));
  NAND2_X1   g01873(.A1(new_n2134_), .A2(new_n2069_), .ZN(new_n2135_));
  INV_X1     g01874(.I(new_n2076_), .ZN(new_n2136_));
  OAI21_X1   g01875(.A1(new_n2135_), .A2(new_n1924_), .B(new_n2136_), .ZN(new_n2137_));
  OAI22_X1   g01876(.A1(new_n2137_), .A2(new_n2080_), .B1(new_n1919_), .B2(new_n2072_), .ZN(new_n2138_));
  NAND2_X1   g01877(.A1(new_n2066_), .A2(new_n1903_), .ZN(new_n2139_));
  OAI21_X1   g01878(.A1(new_n2066_), .A2(new_n1903_), .B(new_n2067_), .ZN(new_n2140_));
  OAI21_X1   g01879(.A1(new_n1978_), .A2(new_n2140_), .B(new_n2139_), .ZN(new_n2141_));
  INV_X1     g01880(.I(new_n2141_), .ZN(new_n2142_));
  INV_X1     g01881(.I(new_n2027_), .ZN(new_n2143_));
  OAI21_X1   g01882(.A1(new_n2027_), .A2(new_n1988_), .B(new_n2032_), .ZN(new_n2144_));
  OAI22_X1   g01883(.A1(new_n2039_), .A2(new_n2144_), .B1(new_n1989_), .B2(new_n2143_), .ZN(new_n2145_));
  XOR2_X1    g01884(.A1(new_n1998_), .A2(new_n1997_), .Z(new_n2146_));
  XOR2_X1    g01885(.A1(new_n2146_), .A2(new_n1993_), .Z(new_n2147_));
  NOR2_X1    g01886(.A1(new_n2147_), .A2(new_n2003_), .ZN(new_n2148_));
  AOI21_X1   g01887(.A1(new_n2025_), .A2(new_n2148_), .B(new_n2014_), .ZN(new_n2149_));
  NOR2_X1    g01888(.A1(new_n2149_), .A2(new_n2022_), .ZN(new_n2150_));
  NAND2_X1   g01889(.A1(new_n1853_), .A2(new_n1997_), .ZN(new_n2151_));
  NOR2_X1    g01890(.A1(new_n1846_), .A2(new_n1993_), .ZN(new_n2152_));
  OAI21_X1   g01891(.A1(new_n1853_), .A2(new_n1997_), .B(new_n2152_), .ZN(new_n2153_));
  NAND2_X1   g01892(.A1(new_n2153_), .A2(new_n2151_), .ZN(new_n2154_));
  OAI22_X1   g01893(.A1(new_n1712_), .A2(new_n298_), .B1(new_n325_), .B2(new_n1707_), .ZN(new_n2155_));
  OAI21_X1   g01894(.A1(new_n280_), .A2(new_n1850_), .B(new_n2155_), .ZN(new_n2156_));
  AOI21_X1   g01895(.A1(new_n2156_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n2157_));
  XOR2_X1    g01896(.A1(new_n2157_), .A2(new_n807_), .Z(new_n2158_));
  XNOR2_X1   g01897(.A1(\a[24] ), .A2(\a[26] ), .ZN(new_n2159_));
  XNOR2_X1   g01898(.A1(\a[23] ), .A2(\a[25] ), .ZN(new_n2160_));
  NOR2_X1    g01899(.A1(new_n2160_), .A2(new_n2159_), .ZN(new_n2161_));
  INV_X1     g01900(.I(\a[25] ), .ZN(new_n2162_));
  NOR3_X1    g01901(.A1(new_n2162_), .A2(\a[23] ), .A3(\a[24] ), .ZN(new_n2163_));
  INV_X1     g01902(.I(\a[24] ), .ZN(new_n2164_));
  NOR3_X1    g01903(.A1(new_n1709_), .A2(new_n2164_), .A3(\a[25] ), .ZN(new_n2165_));
  NOR2_X1    g01904(.A1(new_n2165_), .A2(new_n2163_), .ZN(new_n2166_));
  NOR2_X1    g01905(.A1(new_n2166_), .A2(new_n269_), .ZN(new_n2167_));
  INV_X1     g01906(.I(\a[26] ), .ZN(new_n2168_));
  XOR2_X1    g01907(.A1(\a[24] ), .A2(\a[26] ), .Z(new_n2169_));
  XOR2_X1    g01908(.A1(\a[23] ), .A2(\a[25] ), .Z(new_n2170_));
  NAND2_X1   g01909(.A1(new_n2170_), .A2(new_n2169_), .ZN(new_n2171_));
  OAI21_X1   g01910(.A1(new_n2171_), .A2(new_n258_), .B(new_n2168_), .ZN(new_n2172_));
  OAI21_X1   g01911(.A1(new_n2172_), .A2(new_n2167_), .B(new_n2161_), .ZN(new_n2173_));
  NOR2_X1    g01912(.A1(new_n2173_), .A2(new_n271_), .ZN(new_n2174_));
  INV_X1     g01913(.I(new_n2174_), .ZN(new_n2175_));
  NAND2_X1   g01914(.A1(new_n2173_), .A2(new_n271_), .ZN(new_n2176_));
  NAND2_X1   g01915(.A1(new_n2175_), .A2(new_n2176_), .ZN(new_n2177_));
  NOR2_X1    g01916(.A1(new_n2009_), .A2(new_n2168_), .ZN(new_n2178_));
  INV_X1     g01917(.I(new_n2178_), .ZN(new_n2179_));
  XOR2_X1    g01918(.A1(new_n2177_), .A2(new_n2179_), .Z(new_n2180_));
  XOR2_X1    g01919(.A1(new_n2180_), .A2(new_n2158_), .Z(new_n2181_));
  NAND2_X1   g01920(.A1(new_n2181_), .A2(new_n2154_), .ZN(new_n2182_));
  INV_X1     g01921(.I(new_n2154_), .ZN(new_n2183_));
  INV_X1     g01922(.I(new_n2158_), .ZN(new_n2184_));
  INV_X1     g01923(.I(new_n2180_), .ZN(new_n2185_));
  NOR2_X1    g01924(.A1(new_n2185_), .A2(new_n2184_), .ZN(new_n2186_));
  NOR2_X1    g01925(.A1(new_n2180_), .A2(new_n2158_), .ZN(new_n2187_));
  OAI21_X1   g01926(.A1(new_n2186_), .A2(new_n2187_), .B(new_n2183_), .ZN(new_n2188_));
  NAND2_X1   g01927(.A1(new_n2188_), .A2(new_n2182_), .ZN(new_n2189_));
  INV_X1     g01928(.I(new_n2189_), .ZN(new_n2190_));
  AOI22_X1   g01929(.A1(\b[7] ), .A2(new_n1999_), .B1(new_n1340_), .B2(\b[6] ), .ZN(new_n2191_));
  AOI21_X1   g01930(.A1(\b[5] ), .A2(new_n1458_), .B(new_n2191_), .ZN(new_n2192_));
  OAI21_X1   g01931(.A1(new_n2192_), .A2(\a[20] ), .B(new_n1340_), .ZN(new_n2193_));
  XNOR2_X1   g01932(.A1(new_n471_), .A2(new_n2193_), .ZN(new_n2194_));
  NOR2_X1    g01933(.A1(new_n2190_), .A2(new_n2194_), .ZN(new_n2195_));
  INV_X1     g01934(.I(new_n2194_), .ZN(new_n2196_));
  NOR2_X1    g01935(.A1(new_n2189_), .A2(new_n2196_), .ZN(new_n2197_));
  OAI21_X1   g01936(.A1(new_n2195_), .A2(new_n2197_), .B(new_n2150_), .ZN(new_n2198_));
  INV_X1     g01937(.I(new_n2150_), .ZN(new_n2199_));
  XOR2_X1    g01938(.A1(new_n2189_), .A2(new_n2196_), .Z(new_n2200_));
  NAND2_X1   g01939(.A1(new_n2199_), .A2(new_n2200_), .ZN(new_n2201_));
  NAND2_X1   g01940(.A1(new_n2201_), .A2(new_n2198_), .ZN(new_n2202_));
  OAI22_X1   g01941(.A1(new_n1055_), .A2(new_n565_), .B1(new_n656_), .B2(new_n1061_), .ZN(new_n2203_));
  OAI21_X1   g01942(.A1(new_n515_), .A2(new_n1332_), .B(new_n2203_), .ZN(new_n2204_));
  AOI21_X1   g01943(.A1(new_n2204_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n2205_));
  XNOR2_X1   g01944(.A1(new_n660_), .A2(new_n2205_), .ZN(new_n2206_));
  XOR2_X1    g01945(.A1(new_n2202_), .A2(new_n2206_), .Z(new_n2207_));
  NAND2_X1   g01946(.A1(new_n2145_), .A2(new_n2207_), .ZN(new_n2208_));
  INV_X1     g01947(.I(new_n2145_), .ZN(new_n2209_));
  INV_X1     g01948(.I(new_n2206_), .ZN(new_n2210_));
  XOR2_X1    g01949(.A1(new_n2202_), .A2(new_n2210_), .Z(new_n2211_));
  NAND2_X1   g01950(.A1(new_n2209_), .A2(new_n2211_), .ZN(new_n2212_));
  NAND2_X1   g01951(.A1(new_n2212_), .A2(new_n2208_), .ZN(new_n2213_));
  OAI22_X1   g01952(.A1(new_n970_), .A2(new_n780_), .B1(new_n861_), .B2(new_n820_), .ZN(new_n2214_));
  OAI21_X1   g01953(.A1(new_n706_), .A2(new_n894_), .B(new_n2214_), .ZN(new_n2215_));
  AOI21_X1   g01954(.A1(new_n2215_), .A2(new_n827_), .B(new_n970_), .ZN(new_n2216_));
  XNOR2_X1   g01955(.A1(new_n860_), .A2(new_n2216_), .ZN(new_n2217_));
  INV_X1     g01956(.I(new_n2217_), .ZN(new_n2218_));
  XOR2_X1    g01957(.A1(new_n2213_), .A2(new_n2218_), .Z(new_n2219_));
  INV_X1     g01958(.I(new_n2037_), .ZN(new_n2220_));
  INV_X1     g01959(.I(new_n2042_), .ZN(new_n2221_));
  NOR2_X1    g01960(.A1(new_n2220_), .A2(new_n2221_), .ZN(new_n2222_));
  NOR2_X1    g01961(.A1(new_n2222_), .A2(new_n1980_), .ZN(new_n2223_));
  INV_X1     g01962(.I(new_n2046_), .ZN(new_n2224_));
  NAND3_X1   g01963(.A1(new_n2037_), .A2(new_n2042_), .A3(new_n1980_), .ZN(new_n2225_));
  NAND2_X1   g01964(.A1(new_n2225_), .A2(new_n2224_), .ZN(new_n2226_));
  INV_X1     g01965(.I(new_n2226_), .ZN(new_n2227_));
  AOI21_X1   g01966(.A1(new_n2227_), .A2(new_n2051_), .B(new_n2223_), .ZN(new_n2228_));
  OAI22_X1   g01967(.A1(new_n607_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n610_), .ZN(new_n2229_));
  OAI21_X1   g01968(.A1(new_n930_), .A2(new_n684_), .B(new_n2229_), .ZN(new_n2230_));
  AOI21_X1   g01969(.A1(new_n2230_), .A2(new_n612_), .B(new_n607_), .ZN(new_n2231_));
  XOR2_X1    g01970(.A1(new_n1114_), .A2(new_n2231_), .Z(new_n2232_));
  INV_X1     g01971(.I(new_n2232_), .ZN(new_n2233_));
  NAND2_X1   g01972(.A1(new_n2228_), .A2(new_n2233_), .ZN(new_n2234_));
  OAI22_X1   g01973(.A1(new_n1985_), .A2(new_n2226_), .B1(new_n1980_), .B2(new_n2222_), .ZN(new_n2235_));
  NAND2_X1   g01974(.A1(new_n2235_), .A2(new_n2232_), .ZN(new_n2236_));
  AOI21_X1   g01975(.A1(new_n2234_), .A2(new_n2236_), .B(new_n2219_), .ZN(new_n2237_));
  XOR2_X1    g01976(.A1(new_n2213_), .A2(new_n2217_), .Z(new_n2238_));
  NAND2_X1   g01977(.A1(new_n2235_), .A2(new_n2233_), .ZN(new_n2239_));
  NAND2_X1   g01978(.A1(new_n2228_), .A2(new_n2232_), .ZN(new_n2240_));
  AOI21_X1   g01979(.A1(new_n2240_), .A2(new_n2239_), .B(new_n2238_), .ZN(new_n2241_));
  NOR2_X1    g01980(.A1(new_n2237_), .A2(new_n2241_), .ZN(new_n2242_));
  OAI22_X1   g01981(.A1(new_n448_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n450_), .ZN(new_n2243_));
  OAI21_X1   g01982(.A1(new_n1189_), .A2(new_n496_), .B(new_n2243_), .ZN(new_n2244_));
  AOI21_X1   g01983(.A1(new_n2244_), .A2(new_n452_), .B(new_n448_), .ZN(new_n2245_));
  XNOR2_X1   g01984(.A1(new_n1421_), .A2(new_n2245_), .ZN(new_n2246_));
  XOR2_X1    g01985(.A1(new_n2242_), .A2(new_n2246_), .Z(new_n2247_));
  NOR2_X1    g01986(.A1(new_n2247_), .A2(new_n2142_), .ZN(new_n2248_));
  INV_X1     g01987(.I(new_n2246_), .ZN(new_n2249_));
  XOR2_X1    g01988(.A1(new_n2242_), .A2(new_n2249_), .Z(new_n2250_));
  NOR2_X1    g01989(.A1(new_n2250_), .A2(new_n2141_), .ZN(new_n2251_));
  NOR2_X1    g01990(.A1(new_n2248_), .A2(new_n2251_), .ZN(new_n2252_));
  OAI22_X1   g01991(.A1(new_n1634_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1803_), .ZN(new_n2253_));
  OAI21_X1   g01992(.A1(new_n1525_), .A2(new_n366_), .B(new_n2253_), .ZN(new_n2254_));
  AOI21_X1   g01993(.A1(new_n2254_), .A2(new_n334_), .B(new_n341_), .ZN(new_n2255_));
  XOR2_X1    g01994(.A1(new_n1808_), .A2(new_n2255_), .Z(new_n2256_));
  NOR2_X1    g01995(.A1(new_n2252_), .A2(new_n2256_), .ZN(new_n2257_));
  INV_X1     g01996(.I(new_n2252_), .ZN(new_n2258_));
  INV_X1     g01997(.I(new_n2256_), .ZN(new_n2259_));
  NOR2_X1    g01998(.A1(new_n2258_), .A2(new_n2259_), .ZN(new_n2260_));
  OAI21_X1   g01999(.A1(new_n2257_), .A2(new_n2260_), .B(new_n2138_), .ZN(new_n2261_));
  AOI21_X1   g02000(.A1(new_n2072_), .A2(new_n1919_), .B(new_n2076_), .ZN(new_n2262_));
  AOI22_X1   g02001(.A1(new_n1973_), .A2(new_n2262_), .B1(new_n1924_), .B2(new_n2135_), .ZN(new_n2263_));
  NOR2_X1    g02002(.A1(new_n2258_), .A2(new_n2256_), .ZN(new_n2264_));
  NOR2_X1    g02003(.A1(new_n2252_), .A2(new_n2259_), .ZN(new_n2265_));
  OAI21_X1   g02004(.A1(new_n2264_), .A2(new_n2265_), .B(new_n2263_), .ZN(new_n2266_));
  NAND2_X1   g02005(.A1(new_n2266_), .A2(new_n2261_), .ZN(new_n2267_));
  INV_X1     g02006(.I(new_n2267_), .ZN(new_n2268_));
  NOR2_X1    g02007(.A1(new_n2093_), .A2(new_n2268_), .ZN(new_n2269_));
  OAI21_X1   g02008(.A1(new_n2133_), .A2(new_n2089_), .B(new_n2269_), .ZN(new_n2270_));
  NOR2_X1    g02009(.A1(new_n2133_), .A2(new_n2089_), .ZN(new_n2271_));
  INV_X1     g02010(.I(new_n2271_), .ZN(new_n2272_));
  AOI21_X1   g02011(.A1(new_n2270_), .A2(new_n2272_), .B(new_n1967_), .ZN(new_n2273_));
  AND3_X2    g02012(.A1(new_n2270_), .A2(new_n1967_), .A3(new_n2272_), .Z(new_n2274_));
  NOR2_X1    g02013(.A1(new_n2274_), .A2(new_n2273_), .ZN(new_n2275_));
  XNOR2_X1   g02014(.A1(\b[23] ), .A2(\b[25] ), .ZN(new_n2276_));
  NOR2_X1    g02015(.A1(new_n2276_), .A2(new_n2100_), .ZN(new_n2277_));
  NAND2_X1   g02016(.A1(new_n2099_), .A2(new_n2277_), .ZN(new_n2278_));
  OAI22_X1   g02017(.A1(new_n2095_), .A2(new_n2098_), .B1(new_n2100_), .B2(new_n2276_), .ZN(new_n2279_));
  NAND2_X1   g02018(.A1(new_n2278_), .A2(new_n2279_), .ZN(new_n2280_));
  INV_X1     g02019(.I(\b[25] ), .ZN(new_n2281_));
  OAI22_X1   g02020(.A1(new_n330_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n263_), .ZN(new_n2282_));
  OAI21_X1   g02021(.A1(new_n1936_), .A2(new_n289_), .B(new_n2282_), .ZN(new_n2283_));
  AOI21_X1   g02022(.A1(new_n2283_), .A2(new_n260_), .B(new_n426_), .ZN(new_n2284_));
  XNOR2_X1   g02023(.A1(new_n2280_), .A2(new_n2284_), .ZN(new_n2285_));
  OR2_X2     g02024(.A1(new_n2275_), .A2(new_n2285_), .Z(new_n2286_));
  NAND2_X1   g02025(.A1(new_n2275_), .A2(new_n2285_), .ZN(new_n2287_));
  NAND2_X1   g02026(.A1(new_n2286_), .A2(new_n2287_), .ZN(new_n2288_));
  XOR2_X1    g02027(.A1(new_n2275_), .A2(new_n2285_), .Z(new_n2289_));
  MUX2_X1    g02028(.I0(new_n2289_), .I1(new_n2288_), .S(new_n2132_), .Z(\f[25] ));
  XOR2_X1    g02029(.A1(new_n2138_), .A2(new_n2258_), .Z(new_n2291_));
  NAND2_X1   g02030(.A1(new_n2291_), .A2(new_n2256_), .ZN(new_n2292_));
  INV_X1     g02031(.I(new_n2292_), .ZN(new_n2293_));
  INV_X1     g02032(.I(new_n2089_), .ZN(new_n2294_));
  AOI21_X1   g02033(.A1(new_n2085_), .A2(new_n2267_), .B(new_n2294_), .ZN(new_n2295_));
  NAND4_X1   g02034(.A1(new_n2084_), .A2(new_n2266_), .A3(new_n2261_), .A4(new_n2083_), .ZN(new_n2296_));
  NAND2_X1   g02035(.A1(new_n1967_), .A2(new_n2296_), .ZN(new_n2297_));
  NOR2_X1    g02036(.A1(new_n2297_), .A2(new_n2295_), .ZN(new_n2298_));
  OAI21_X1   g02037(.A1(new_n2237_), .A2(new_n2241_), .B(new_n2142_), .ZN(new_n2299_));
  NAND2_X1   g02038(.A1(new_n2141_), .A2(new_n2242_), .ZN(new_n2300_));
  AOI21_X1   g02039(.A1(new_n2299_), .A2(new_n2300_), .B(new_n2249_), .ZN(new_n2301_));
  INV_X1     g02040(.I(new_n2301_), .ZN(new_n2302_));
  NAND2_X1   g02041(.A1(new_n2235_), .A2(new_n2238_), .ZN(new_n2303_));
  NAND2_X1   g02042(.A1(new_n2228_), .A2(new_n2219_), .ZN(new_n2304_));
  AOI21_X1   g02043(.A1(new_n2304_), .A2(new_n2303_), .B(new_n2233_), .ZN(new_n2305_));
  NOR2_X1    g02044(.A1(new_n2213_), .A2(new_n2217_), .ZN(new_n2306_));
  INV_X1     g02045(.I(new_n2213_), .ZN(new_n2307_));
  NOR2_X1    g02046(.A1(new_n2307_), .A2(new_n2218_), .ZN(new_n2308_));
  INV_X1     g02047(.I(new_n2308_), .ZN(new_n2309_));
  AOI21_X1   g02048(.A1(new_n2235_), .A2(new_n2309_), .B(new_n2306_), .ZN(new_n2310_));
  NAND2_X1   g02049(.A1(new_n2202_), .A2(new_n2210_), .ZN(new_n2311_));
  OAI22_X1   g02050(.A1(new_n1347_), .A2(new_n472_), .B1(new_n515_), .B2(new_n1344_), .ZN(new_n2312_));
  OAI21_X1   g02051(.A1(new_n420_), .A2(new_n1457_), .B(new_n2312_), .ZN(new_n2313_));
  AOI21_X1   g02052(.A1(new_n2313_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n2314_));
  XOR2_X1    g02053(.A1(new_n700_), .A2(new_n2314_), .Z(new_n2315_));
  INV_X1     g02054(.I(new_n2315_), .ZN(new_n2316_));
  NAND3_X1   g02055(.A1(new_n2175_), .A2(new_n2176_), .A3(new_n2178_), .ZN(new_n2317_));
  NOR2_X1    g02056(.A1(new_n2166_), .A2(new_n280_), .ZN(new_n2318_));
  AOI21_X1   g02057(.A1(new_n269_), .A2(new_n490_), .B(new_n2171_), .ZN(new_n2319_));
  NOR2_X1    g02058(.A1(new_n2319_), .A2(new_n2318_), .ZN(new_n2320_));
  XOR2_X1    g02059(.A1(\a[23] ), .A2(\a[26] ), .Z(new_n2321_));
  NAND3_X1   g02060(.A1(new_n2170_), .A2(new_n1992_), .A3(new_n2321_), .ZN(new_n2322_));
  NOR3_X1    g02061(.A1(new_n2320_), .A2(new_n258_), .A3(new_n2322_), .ZN(new_n2323_));
  NOR2_X1    g02062(.A1(new_n2323_), .A2(new_n2168_), .ZN(new_n2324_));
  NAND2_X1   g02063(.A1(new_n2323_), .A2(new_n2168_), .ZN(new_n2325_));
  INV_X1     g02064(.I(new_n2325_), .ZN(new_n2326_));
  NOR2_X1    g02065(.A1(new_n2326_), .A2(new_n2324_), .ZN(new_n2327_));
  XOR2_X1    g02066(.A1(new_n2327_), .A2(new_n2317_), .Z(new_n2328_));
  INV_X1     g02067(.I(new_n2187_), .ZN(new_n2329_));
  OAI21_X1   g02068(.A1(new_n2184_), .A2(new_n2185_), .B(new_n2154_), .ZN(new_n2330_));
  NOR4_X1    g02069(.A1(new_n322_), .A2(new_n319_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n2331_));
  AOI22_X1   g02070(.A1(new_n317_), .A2(new_n268_), .B1(new_n323_), .B2(new_n373_), .ZN(new_n2332_));
  NOR2_X1    g02071(.A1(new_n2332_), .A2(new_n2331_), .ZN(new_n2333_));
  NOR2_X1    g02072(.A1(new_n2333_), .A2(new_n1712_), .ZN(new_n2334_));
  OAI22_X1   g02073(.A1(new_n1712_), .A2(new_n325_), .B1(new_n419_), .B2(new_n1707_), .ZN(new_n2335_));
  OAI21_X1   g02074(.A1(new_n298_), .A2(new_n1850_), .B(new_n2335_), .ZN(new_n2336_));
  NOR2_X1    g02075(.A1(new_n2334_), .A2(new_n2336_), .ZN(new_n2337_));
  XOR2_X1    g02076(.A1(new_n2337_), .A2(new_n1709_), .Z(new_n2338_));
  INV_X1     g02077(.I(new_n2338_), .ZN(new_n2339_));
  NAND3_X1   g02078(.A1(new_n2330_), .A2(new_n2329_), .A3(new_n2339_), .ZN(new_n2340_));
  INV_X1     g02079(.I(new_n2340_), .ZN(new_n2341_));
  AOI21_X1   g02080(.A1(new_n2330_), .A2(new_n2329_), .B(new_n2339_), .ZN(new_n2342_));
  OAI21_X1   g02081(.A1(new_n2341_), .A2(new_n2342_), .B(new_n2328_), .ZN(new_n2343_));
  INV_X1     g02082(.I(new_n2328_), .ZN(new_n2344_));
  INV_X1     g02083(.I(new_n2342_), .ZN(new_n2345_));
  NAND3_X1   g02084(.A1(new_n2345_), .A2(new_n2344_), .A3(new_n2340_), .ZN(new_n2346_));
  AOI21_X1   g02085(.A1(new_n2346_), .A2(new_n2343_), .B(new_n2316_), .ZN(new_n2347_));
  NAND3_X1   g02086(.A1(new_n2346_), .A2(new_n2343_), .A3(new_n2316_), .ZN(new_n2348_));
  INV_X1     g02087(.I(new_n2348_), .ZN(new_n2349_));
  OAI21_X1   g02088(.A1(new_n2349_), .A2(new_n2347_), .B(new_n2200_), .ZN(new_n2350_));
  NOR2_X1    g02089(.A1(new_n2350_), .A2(new_n2195_), .ZN(new_n2351_));
  INV_X1     g02090(.I(new_n2343_), .ZN(new_n2352_));
  NOR3_X1    g02091(.A1(new_n2341_), .A2(new_n2328_), .A3(new_n2342_), .ZN(new_n2353_));
  OAI21_X1   g02092(.A1(new_n2352_), .A2(new_n2353_), .B(new_n2315_), .ZN(new_n2354_));
  NAND2_X1   g02093(.A1(new_n2354_), .A2(new_n2348_), .ZN(new_n2355_));
  NOR2_X1    g02094(.A1(new_n2190_), .A2(new_n2194_), .ZN(new_n2357_));
  OAI21_X1   g02095(.A1(new_n2351_), .A2(new_n2357_), .B(new_n2199_), .ZN(new_n2358_));
  INV_X1     g02096(.I(new_n2195_), .ZN(new_n2359_));
  NAND3_X1   g02097(.A1(new_n2355_), .A2(new_n2359_), .A3(new_n2200_), .ZN(new_n2360_));
  INV_X1     g02098(.I(new_n2357_), .ZN(new_n2361_));
  NAND3_X1   g02099(.A1(new_n2360_), .A2(new_n2150_), .A3(new_n2361_), .ZN(new_n2362_));
  OAI22_X1   g02100(.A1(new_n1055_), .A2(new_n656_), .B1(new_n706_), .B2(new_n1061_), .ZN(new_n2363_));
  OAI21_X1   g02101(.A1(new_n565_), .A2(new_n1332_), .B(new_n2363_), .ZN(new_n2364_));
  AOI21_X1   g02102(.A1(new_n2364_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n2365_));
  XNOR2_X1   g02103(.A1(new_n710_), .A2(new_n2365_), .ZN(new_n2366_));
  AOI21_X1   g02104(.A1(new_n2358_), .A2(new_n2362_), .B(new_n2366_), .ZN(new_n2367_));
  AOI21_X1   g02105(.A1(new_n2360_), .A2(new_n2361_), .B(new_n2150_), .ZN(new_n2368_));
  NOR3_X1    g02106(.A1(new_n2351_), .A2(new_n2199_), .A3(new_n2357_), .ZN(new_n2369_));
  INV_X1     g02107(.I(new_n2366_), .ZN(new_n2370_));
  NOR3_X1    g02108(.A1(new_n2369_), .A2(new_n2368_), .A3(new_n2370_), .ZN(new_n2371_));
  OR2_X2     g02109(.A1(new_n2371_), .A2(new_n2367_), .Z(new_n2372_));
  NAND3_X1   g02110(.A1(new_n2372_), .A2(new_n2211_), .A3(new_n2311_), .ZN(new_n2373_));
  NAND2_X1   g02111(.A1(new_n2202_), .A2(new_n2210_), .ZN(new_n2375_));
  AOI21_X1   g02112(.A1(new_n2373_), .A2(new_n2375_), .B(new_n2145_), .ZN(new_n2376_));
  NAND3_X1   g02113(.A1(new_n2373_), .A2(new_n2145_), .A3(new_n2375_), .ZN(new_n2377_));
  INV_X1     g02114(.I(new_n2377_), .ZN(new_n2378_));
  OAI22_X1   g02115(.A1(new_n970_), .A2(new_n861_), .B1(new_n930_), .B2(new_n820_), .ZN(new_n2379_));
  OAI21_X1   g02116(.A1(new_n780_), .A2(new_n894_), .B(new_n2379_), .ZN(new_n2380_));
  AOI21_X1   g02117(.A1(new_n2380_), .A2(new_n827_), .B(new_n970_), .ZN(new_n2381_));
  XNOR2_X1   g02118(.A1(new_n937_), .A2(new_n2381_), .ZN(new_n2382_));
  NOR3_X1    g02119(.A1(new_n2378_), .A2(new_n2376_), .A3(new_n2382_), .ZN(new_n2383_));
  AND3_X2    g02120(.A1(new_n2372_), .A2(new_n2211_), .A3(new_n2311_), .Z(new_n2384_));
  INV_X1     g02121(.I(new_n2375_), .ZN(new_n2385_));
  OAI21_X1   g02122(.A1(new_n2384_), .A2(new_n2385_), .B(new_n2209_), .ZN(new_n2386_));
  INV_X1     g02123(.I(new_n2382_), .ZN(new_n2387_));
  AOI21_X1   g02124(.A1(new_n2386_), .A2(new_n2377_), .B(new_n2387_), .ZN(new_n2388_));
  NOR2_X1    g02125(.A1(new_n2383_), .A2(new_n2388_), .ZN(new_n2389_));
  OAI22_X1   g02126(.A1(new_n607_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n610_), .ZN(new_n2390_));
  OAI21_X1   g02127(.A1(new_n1017_), .A2(new_n684_), .B(new_n2390_), .ZN(new_n2391_));
  AOI21_X1   g02128(.A1(new_n2391_), .A2(new_n612_), .B(new_n607_), .ZN(new_n2392_));
  XNOR2_X1   g02129(.A1(new_n1196_), .A2(new_n2392_), .ZN(new_n2393_));
  INV_X1     g02130(.I(new_n2393_), .ZN(new_n2394_));
  NAND2_X1   g02131(.A1(new_n2389_), .A2(new_n2394_), .ZN(new_n2395_));
  NAND3_X1   g02132(.A1(new_n2386_), .A2(new_n2377_), .A3(new_n2387_), .ZN(new_n2396_));
  OAI21_X1   g02133(.A1(new_n2378_), .A2(new_n2376_), .B(new_n2382_), .ZN(new_n2397_));
  NAND2_X1   g02134(.A1(new_n2397_), .A2(new_n2396_), .ZN(new_n2398_));
  NAND2_X1   g02135(.A1(new_n2398_), .A2(new_n2393_), .ZN(new_n2399_));
  AOI21_X1   g02136(.A1(new_n2395_), .A2(new_n2399_), .B(new_n2310_), .ZN(new_n2400_));
  INV_X1     g02137(.I(new_n2306_), .ZN(new_n2401_));
  OAI21_X1   g02138(.A1(new_n2228_), .A2(new_n2308_), .B(new_n2401_), .ZN(new_n2402_));
  NAND2_X1   g02139(.A1(new_n2398_), .A2(new_n2394_), .ZN(new_n2403_));
  NAND2_X1   g02140(.A1(new_n2389_), .A2(new_n2393_), .ZN(new_n2404_));
  AOI21_X1   g02141(.A1(new_n2404_), .A2(new_n2403_), .B(new_n2402_), .ZN(new_n2405_));
  NOR3_X1    g02142(.A1(new_n2400_), .A2(new_n2405_), .A3(new_n2305_), .ZN(new_n2406_));
  NOR2_X1    g02143(.A1(new_n2406_), .A2(new_n2242_), .ZN(new_n2407_));
  NAND2_X1   g02144(.A1(new_n2142_), .A2(new_n2407_), .ZN(new_n2408_));
  NOR2_X1    g02145(.A1(new_n2142_), .A2(new_n2407_), .ZN(new_n2409_));
  INV_X1     g02146(.I(new_n2409_), .ZN(new_n2410_));
  OAI22_X1   g02147(.A1(new_n448_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n450_), .ZN(new_n2411_));
  OAI21_X1   g02148(.A1(new_n1294_), .A2(new_n496_), .B(new_n2411_), .ZN(new_n2412_));
  AOI21_X1   g02149(.A1(new_n2412_), .A2(new_n452_), .B(new_n448_), .ZN(new_n2413_));
  XOR2_X1    g02150(.A1(new_n1530_), .A2(new_n2413_), .Z(new_n2414_));
  INV_X1     g02151(.I(new_n2414_), .ZN(new_n2415_));
  NAND3_X1   g02152(.A1(new_n2410_), .A2(new_n2408_), .A3(new_n2415_), .ZN(new_n2416_));
  INV_X1     g02153(.I(new_n2408_), .ZN(new_n2417_));
  OAI21_X1   g02154(.A1(new_n2417_), .A2(new_n2409_), .B(new_n2414_), .ZN(new_n2418_));
  NAND2_X1   g02155(.A1(new_n2418_), .A2(new_n2416_), .ZN(new_n2419_));
  INV_X1     g02156(.I(new_n2419_), .ZN(new_n2420_));
  AOI21_X1   g02157(.A1(new_n2420_), .A2(new_n2302_), .B(new_n2252_), .ZN(new_n2421_));
  AND2_X2    g02158(.A1(new_n2421_), .A2(new_n2263_), .Z(new_n2422_));
  NOR2_X1    g02159(.A1(new_n2421_), .A2(new_n2263_), .ZN(new_n2423_));
  NOR2_X1    g02160(.A1(new_n2422_), .A2(new_n2423_), .ZN(new_n2424_));
  OAI22_X1   g02161(.A1(new_n1803_), .A2(new_n341_), .B1(new_n404_), .B2(new_n1936_), .ZN(new_n2425_));
  OAI21_X1   g02162(.A1(new_n1634_), .A2(new_n366_), .B(new_n2425_), .ZN(new_n2426_));
  AOI21_X1   g02163(.A1(new_n2426_), .A2(new_n334_), .B(new_n341_), .ZN(new_n2427_));
  XNOR2_X1   g02164(.A1(new_n1940_), .A2(new_n2427_), .ZN(new_n2428_));
  INV_X1     g02165(.I(new_n2428_), .ZN(new_n2429_));
  NAND2_X1   g02166(.A1(new_n2424_), .A2(new_n2429_), .ZN(new_n2430_));
  OAI21_X1   g02167(.A1(new_n2422_), .A2(new_n2423_), .B(new_n2428_), .ZN(new_n2431_));
  NOR2_X1    g02168(.A1(\b[24] ), .A2(\b[25] ), .ZN(new_n2432_));
  AOI21_X1   g02169(.A1(new_n2099_), .A2(new_n2432_), .B(new_n1936_), .ZN(new_n2433_));
  NOR2_X1    g02170(.A1(new_n2102_), .A2(new_n2281_), .ZN(new_n2434_));
  INV_X1     g02171(.I(new_n2434_), .ZN(new_n2435_));
  NOR2_X1    g02172(.A1(new_n2099_), .A2(new_n2435_), .ZN(new_n2436_));
  NOR2_X1    g02173(.A1(new_n2433_), .A2(new_n2436_), .ZN(new_n2437_));
  XNOR2_X1   g02174(.A1(\b[25] ), .A2(\b[26] ), .ZN(new_n2438_));
  INV_X1     g02175(.I(\b[26] ), .ZN(new_n2439_));
  NOR2_X1    g02176(.A1(new_n2281_), .A2(new_n2439_), .ZN(new_n2440_));
  NOR2_X1    g02177(.A1(\b[25] ), .A2(\b[26] ), .ZN(new_n2441_));
  OAI21_X1   g02178(.A1(new_n2440_), .A2(new_n2441_), .B(new_n2437_), .ZN(new_n2442_));
  OAI21_X1   g02179(.A1(new_n2437_), .A2(new_n2438_), .B(new_n2442_), .ZN(new_n2443_));
  OAI22_X1   g02180(.A1(new_n330_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n263_), .ZN(new_n2444_));
  OAI21_X1   g02181(.A1(new_n2102_), .A2(new_n289_), .B(new_n2444_), .ZN(new_n2445_));
  AOI21_X1   g02182(.A1(new_n2445_), .A2(new_n260_), .B(new_n426_), .ZN(new_n2446_));
  XNOR2_X1   g02183(.A1(new_n2443_), .A2(new_n2446_), .ZN(new_n2447_));
  AOI21_X1   g02184(.A1(new_n2430_), .A2(new_n2431_), .B(new_n2447_), .ZN(new_n2448_));
  INV_X1     g02185(.I(new_n2448_), .ZN(new_n2449_));
  NOR2_X1    g02186(.A1(new_n2449_), .A2(new_n2298_), .ZN(new_n2450_));
  NAND2_X1   g02187(.A1(new_n2449_), .A2(new_n2298_), .ZN(new_n2451_));
  INV_X1     g02188(.I(new_n2451_), .ZN(new_n2452_));
  NOR2_X1    g02189(.A1(new_n2452_), .A2(new_n2450_), .ZN(new_n2453_));
  NOR2_X1    g02190(.A1(new_n2453_), .A2(new_n2293_), .ZN(new_n2454_));
  NOR3_X1    g02191(.A1(new_n2452_), .A2(new_n2292_), .A3(new_n2450_), .ZN(new_n2455_));
  NOR2_X1    g02192(.A1(new_n2454_), .A2(new_n2455_), .ZN(new_n2456_));
  INV_X1     g02193(.I(new_n2456_), .ZN(new_n2457_));
  NAND2_X1   g02194(.A1(new_n2289_), .A2(new_n2457_), .ZN(new_n2458_));
  XOR2_X1    g02195(.A1(new_n2458_), .A2(new_n2286_), .Z(new_n2459_));
  XOR2_X1    g02196(.A1(new_n2459_), .A2(new_n2132_), .Z(\f[26] ));
  XOR2_X1    g02197(.A1(new_n2448_), .A2(new_n2293_), .Z(new_n2461_));
  NAND2_X1   g02198(.A1(new_n2461_), .A2(new_n2298_), .ZN(new_n2462_));
  OAI21_X1   g02199(.A1(new_n2456_), .A2(new_n2275_), .B(new_n2285_), .ZN(new_n2463_));
  NAND2_X1   g02200(.A1(new_n2456_), .A2(new_n2275_), .ZN(new_n2464_));
  INV_X1     g02201(.I(new_n2464_), .ZN(new_n2465_));
  NOR3_X1    g02202(.A1(new_n2465_), .A2(new_n1962_), .A3(new_n2131_), .ZN(new_n2466_));
  NAND2_X1   g02203(.A1(new_n2466_), .A2(new_n2463_), .ZN(new_n2467_));
  NOR2_X1    g02204(.A1(new_n2292_), .A2(new_n2424_), .ZN(new_n2468_));
  AOI21_X1   g02205(.A1(new_n2292_), .A2(new_n2424_), .B(new_n2428_), .ZN(new_n2469_));
  AOI21_X1   g02206(.A1(new_n2298_), .A2(new_n2469_), .B(new_n2468_), .ZN(new_n2470_));
  INV_X1     g02207(.I(new_n2470_), .ZN(new_n2471_));
  AOI21_X1   g02208(.A1(new_n2419_), .A2(new_n2301_), .B(new_n2258_), .ZN(new_n2472_));
  XOR2_X1    g02209(.A1(new_n2310_), .A2(new_n2398_), .Z(new_n2473_));
  NOR2_X1    g02210(.A1(new_n2473_), .A2(new_n2394_), .ZN(new_n2474_));
  AOI21_X1   g02211(.A1(new_n2058_), .A2(new_n1974_), .B(new_n2062_), .ZN(new_n2475_));
  NAND4_X1   g02212(.A1(new_n2475_), .A2(new_n1833_), .A3(new_n1976_), .A4(new_n1977_), .ZN(new_n2476_));
  OAI21_X1   g02213(.A1(new_n2405_), .A2(new_n2400_), .B(new_n2305_), .ZN(new_n2477_));
  AOI22_X1   g02214(.A1(new_n2476_), .A2(new_n2139_), .B1(new_n2477_), .B2(new_n2242_), .ZN(new_n2478_));
  OAI21_X1   g02215(.A1(new_n2389_), .A2(new_n2307_), .B(new_n2217_), .ZN(new_n2479_));
  NAND2_X1   g02216(.A1(new_n2389_), .A2(new_n2307_), .ZN(new_n2480_));
  NAND3_X1   g02217(.A1(new_n2479_), .A2(new_n2480_), .A3(new_n2235_), .ZN(new_n2481_));
  AOI21_X1   g02218(.A1(new_n2358_), .A2(new_n2362_), .B(new_n2370_), .ZN(new_n2482_));
  INV_X1     g02219(.I(new_n2482_), .ZN(new_n2483_));
  OAI21_X1   g02220(.A1(new_n2371_), .A2(new_n2367_), .B(new_n2202_), .ZN(new_n2484_));
  NAND2_X1   g02221(.A1(new_n2484_), .A2(new_n2206_), .ZN(new_n2485_));
  OR3_X2     g02222(.A1(new_n2371_), .A2(new_n2367_), .A3(new_n2202_), .Z(new_n2486_));
  NAND3_X1   g02223(.A1(new_n2485_), .A2(new_n2486_), .A3(new_n2145_), .ZN(new_n2487_));
  NAND2_X1   g02224(.A1(new_n2330_), .A2(new_n2329_), .ZN(new_n2488_));
  XOR2_X1    g02225(.A1(new_n2488_), .A2(new_n2328_), .Z(new_n2489_));
  OR2_X2     g02226(.A1(new_n2489_), .A2(new_n2339_), .Z(new_n2490_));
  NAND2_X1   g02227(.A1(new_n2489_), .A2(new_n2339_), .ZN(new_n2491_));
  AOI21_X1   g02228(.A1(new_n2490_), .A2(new_n2491_), .B(new_n2315_), .ZN(new_n2492_));
  INV_X1     g02229(.I(new_n2492_), .ZN(new_n2493_));
  OAI21_X1   g02230(.A1(new_n2349_), .A2(new_n2347_), .B(new_n2189_), .ZN(new_n2494_));
  NAND2_X1   g02231(.A1(new_n2494_), .A2(new_n2194_), .ZN(new_n2495_));
  NAND3_X1   g02232(.A1(new_n2354_), .A2(new_n2348_), .A3(new_n2190_), .ZN(new_n2496_));
  AND2_X2    g02233(.A1(new_n2496_), .A2(new_n2150_), .Z(new_n2497_));
  XOR2_X1    g02234(.A1(\a[26] ), .A2(\a[27] ), .Z(new_n2498_));
  NAND2_X1   g02235(.A1(new_n2498_), .A2(\b[0] ), .ZN(new_n2499_));
  INV_X1     g02236(.I(new_n2499_), .ZN(new_n2500_));
  NOR2_X1    g02237(.A1(new_n2322_), .A2(new_n269_), .ZN(new_n2501_));
  OAI22_X1   g02238(.A1(new_n2171_), .A2(new_n280_), .B1(new_n298_), .B2(new_n2166_), .ZN(new_n2502_));
  NOR2_X1    g02239(.A1(new_n2502_), .A2(new_n2501_), .ZN(new_n2503_));
  NOR3_X1    g02240(.A1(new_n2503_), .A2(new_n403_), .A3(new_n2171_), .ZN(new_n2504_));
  NOR2_X1    g02241(.A1(new_n2504_), .A2(new_n2168_), .ZN(new_n2505_));
  NAND2_X1   g02242(.A1(new_n2504_), .A2(new_n2168_), .ZN(new_n2506_));
  INV_X1     g02243(.I(new_n2506_), .ZN(new_n2507_));
  NOR2_X1    g02244(.A1(new_n2507_), .A2(new_n2505_), .ZN(new_n2508_));
  INV_X1     g02245(.I(new_n2317_), .ZN(new_n2509_));
  OAI22_X1   g02246(.A1(new_n1712_), .A2(new_n419_), .B1(new_n420_), .B2(new_n1707_), .ZN(new_n2510_));
  OAI21_X1   g02247(.A1(new_n325_), .A2(new_n1850_), .B(new_n2510_), .ZN(new_n2511_));
  AOI21_X1   g02248(.A1(new_n2511_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n2512_));
  INV_X1     g02249(.I(new_n2512_), .ZN(new_n2513_));
  NOR2_X1    g02250(.A1(new_n556_), .A2(new_n2513_), .ZN(new_n2514_));
  INV_X1     g02251(.I(new_n2514_), .ZN(new_n2515_));
  NAND2_X1   g02252(.A1(new_n556_), .A2(new_n2513_), .ZN(new_n2516_));
  AOI22_X1   g02253(.A1(new_n2515_), .A2(new_n2516_), .B1(new_n2327_), .B2(new_n2509_), .ZN(new_n2517_));
  INV_X1     g02254(.I(new_n2324_), .ZN(new_n2518_));
  NAND2_X1   g02255(.A1(new_n2518_), .A2(new_n2325_), .ZN(new_n2519_));
  INV_X1     g02256(.I(new_n2516_), .ZN(new_n2520_));
  NOR4_X1    g02257(.A1(new_n2520_), .A2(new_n2514_), .A3(new_n2519_), .A4(new_n2317_), .ZN(new_n2521_));
  OAI21_X1   g02258(.A1(new_n2517_), .A2(new_n2521_), .B(new_n2508_), .ZN(new_n2522_));
  INV_X1     g02259(.I(new_n2505_), .ZN(new_n2523_));
  NAND2_X1   g02260(.A1(new_n2523_), .A2(new_n2506_), .ZN(new_n2524_));
  OAI22_X1   g02261(.A1(new_n2520_), .A2(new_n2514_), .B1(new_n2519_), .B2(new_n2317_), .ZN(new_n2525_));
  NAND4_X1   g02262(.A1(new_n2515_), .A2(new_n2516_), .A3(new_n2327_), .A4(new_n2509_), .ZN(new_n2526_));
  NAND3_X1   g02263(.A1(new_n2525_), .A2(new_n2526_), .A3(new_n2524_), .ZN(new_n2527_));
  AOI21_X1   g02264(.A1(new_n2522_), .A2(new_n2527_), .B(new_n2500_), .ZN(new_n2528_));
  AOI21_X1   g02265(.A1(new_n2525_), .A2(new_n2526_), .B(new_n2524_), .ZN(new_n2529_));
  NOR3_X1    g02266(.A1(new_n2517_), .A2(new_n2521_), .A3(new_n2508_), .ZN(new_n2530_));
  NOR3_X1    g02267(.A1(new_n2530_), .A2(new_n2529_), .A3(new_n2499_), .ZN(new_n2531_));
  OR2_X2     g02268(.A1(new_n2531_), .A2(new_n2528_), .Z(new_n2532_));
  INV_X1     g02269(.I(new_n2532_), .ZN(new_n2533_));
  NAND2_X1   g02270(.A1(new_n2344_), .A2(new_n2338_), .ZN(new_n2534_));
  NAND2_X1   g02271(.A1(new_n2317_), .A2(new_n2337_), .ZN(new_n2535_));
  NOR2_X1    g02272(.A1(new_n2317_), .A2(new_n2337_), .ZN(new_n2536_));
  INV_X1     g02273(.I(new_n2536_), .ZN(new_n2537_));
  AOI21_X1   g02274(.A1(new_n2537_), .A2(new_n2535_), .B(new_n2519_), .ZN(new_n2538_));
  INV_X1     g02275(.I(new_n2535_), .ZN(new_n2539_));
  NOR3_X1    g02276(.A1(new_n2539_), .A2(new_n2536_), .A3(new_n2327_), .ZN(new_n2540_));
  OAI21_X1   g02277(.A1(new_n2538_), .A2(new_n2540_), .B(new_n1709_), .ZN(new_n2541_));
  OAI21_X1   g02278(.A1(new_n2539_), .A2(new_n2536_), .B(new_n2327_), .ZN(new_n2542_));
  NAND3_X1   g02279(.A1(new_n2537_), .A2(new_n2535_), .A3(new_n2519_), .ZN(new_n2543_));
  NAND3_X1   g02280(.A1(new_n2542_), .A2(new_n2543_), .A3(\a[23] ), .ZN(new_n2544_));
  NAND2_X1   g02281(.A1(new_n2541_), .A2(new_n2544_), .ZN(new_n2545_));
  AOI21_X1   g02282(.A1(new_n2545_), .A2(new_n2180_), .B(new_n2184_), .ZN(new_n2546_));
  OAI21_X1   g02283(.A1(new_n2545_), .A2(new_n2180_), .B(new_n2154_), .ZN(new_n2547_));
  OR2_X2     g02284(.A1(new_n2546_), .A2(new_n2547_), .Z(new_n2548_));
  NAND2_X1   g02285(.A1(new_n2548_), .A2(new_n2534_), .ZN(new_n2549_));
  NAND2_X1   g02286(.A1(new_n2549_), .A2(new_n2533_), .ZN(new_n2550_));
  NAND3_X1   g02287(.A1(new_n2548_), .A2(new_n2532_), .A3(new_n2534_), .ZN(new_n2551_));
  NAND2_X1   g02288(.A1(new_n2550_), .A2(new_n2551_), .ZN(new_n2552_));
  OAI22_X1   g02289(.A1(new_n1347_), .A2(new_n515_), .B1(new_n565_), .B2(new_n1344_), .ZN(new_n2553_));
  OAI21_X1   g02290(.A1(new_n472_), .A2(new_n1457_), .B(new_n2553_), .ZN(new_n2554_));
  AOI21_X1   g02291(.A1(new_n2554_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n2555_));
  XOR2_X1    g02292(.A1(new_n759_), .A2(new_n2555_), .Z(new_n2556_));
  INV_X1     g02293(.I(new_n2556_), .ZN(new_n2557_));
  NAND2_X1   g02294(.A1(new_n2552_), .A2(new_n2557_), .ZN(new_n2558_));
  AOI21_X1   g02295(.A1(new_n2497_), .A2(new_n2495_), .B(new_n2558_), .ZN(new_n2559_));
  NAND3_X1   g02296(.A1(new_n2495_), .A2(new_n2150_), .A3(new_n2496_), .ZN(new_n2560_));
  INV_X1     g02297(.I(new_n2558_), .ZN(new_n2561_));
  NOR2_X1    g02298(.A1(new_n2560_), .A2(new_n2561_), .ZN(new_n2562_));
  OAI21_X1   g02299(.A1(new_n2562_), .A2(new_n2559_), .B(new_n2493_), .ZN(new_n2563_));
  NAND2_X1   g02300(.A1(new_n2560_), .A2(new_n2561_), .ZN(new_n2564_));
  NAND3_X1   g02301(.A1(new_n2497_), .A2(new_n2495_), .A3(new_n2558_), .ZN(new_n2565_));
  NAND3_X1   g02302(.A1(new_n2564_), .A2(new_n2565_), .A3(new_n2492_), .ZN(new_n2566_));
  NAND2_X1   g02303(.A1(new_n2563_), .A2(new_n2566_), .ZN(new_n2567_));
  OAI22_X1   g02304(.A1(new_n1055_), .A2(new_n706_), .B1(new_n780_), .B2(new_n1061_), .ZN(new_n2568_));
  OAI21_X1   g02305(.A1(new_n656_), .A2(new_n1332_), .B(new_n2568_), .ZN(new_n2569_));
  AOI21_X1   g02306(.A1(new_n2569_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n2570_));
  XOR2_X1    g02307(.A1(new_n785_), .A2(new_n2570_), .Z(new_n2571_));
  INV_X1     g02308(.I(new_n2571_), .ZN(new_n2572_));
  NAND3_X1   g02309(.A1(new_n2487_), .A2(new_n2567_), .A3(new_n2572_), .ZN(new_n2573_));
  INV_X1     g02310(.I(new_n2573_), .ZN(new_n2574_));
  AOI21_X1   g02311(.A1(new_n2567_), .A2(new_n2572_), .B(new_n2487_), .ZN(new_n2575_));
  OAI21_X1   g02312(.A1(new_n2574_), .A2(new_n2575_), .B(new_n2483_), .ZN(new_n2576_));
  INV_X1     g02313(.I(new_n2575_), .ZN(new_n2577_));
  NAND3_X1   g02314(.A1(new_n2577_), .A2(new_n2482_), .A3(new_n2573_), .ZN(new_n2578_));
  OAI22_X1   g02315(.A1(new_n970_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n820_), .ZN(new_n2579_));
  OAI21_X1   g02316(.A1(new_n861_), .A2(new_n894_), .B(new_n2579_), .ZN(new_n2580_));
  AOI21_X1   g02317(.A1(new_n2580_), .A2(new_n827_), .B(new_n970_), .ZN(new_n2581_));
  XOR2_X1    g02318(.A1(new_n1024_), .A2(new_n2581_), .Z(new_n2582_));
  AOI21_X1   g02319(.A1(new_n2578_), .A2(new_n2576_), .B(new_n2582_), .ZN(new_n2583_));
  NAND2_X1   g02320(.A1(new_n2481_), .A2(new_n2583_), .ZN(new_n2584_));
  AOI21_X1   g02321(.A1(new_n2398_), .A2(new_n2213_), .B(new_n2218_), .ZN(new_n2585_));
  NOR2_X1    g02322(.A1(new_n2398_), .A2(new_n2213_), .ZN(new_n2586_));
  NOR3_X1    g02323(.A1(new_n2585_), .A2(new_n2586_), .A3(new_n2228_), .ZN(new_n2587_));
  INV_X1     g02324(.I(new_n2583_), .ZN(new_n2588_));
  NAND2_X1   g02325(.A1(new_n2587_), .A2(new_n2588_), .ZN(new_n2589_));
  AOI21_X1   g02326(.A1(new_n2584_), .A2(new_n2589_), .B(new_n2388_), .ZN(new_n2590_));
  NOR2_X1    g02327(.A1(new_n2587_), .A2(new_n2588_), .ZN(new_n2591_));
  NOR2_X1    g02328(.A1(new_n2481_), .A2(new_n2583_), .ZN(new_n2592_));
  NOR3_X1    g02329(.A1(new_n2592_), .A2(new_n2591_), .A3(new_n2397_), .ZN(new_n2593_));
  NOR2_X1    g02330(.A1(new_n2590_), .A2(new_n2593_), .ZN(new_n2594_));
  OAI22_X1   g02331(.A1(new_n607_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n610_), .ZN(new_n2595_));
  OAI21_X1   g02332(.A1(new_n1109_), .A2(new_n684_), .B(new_n2595_), .ZN(new_n2596_));
  AOI21_X1   g02333(.A1(new_n2596_), .A2(new_n612_), .B(new_n607_), .ZN(new_n2597_));
  XOR2_X1    g02334(.A1(new_n1299_), .A2(new_n2597_), .Z(new_n2598_));
  NOR3_X1    g02335(.A1(new_n2478_), .A2(new_n2594_), .A3(new_n2598_), .ZN(new_n2599_));
  INV_X1     g02336(.I(new_n2599_), .ZN(new_n2600_));
  NAND2_X1   g02337(.A1(new_n2477_), .A2(new_n2242_), .ZN(new_n2601_));
  NAND2_X1   g02338(.A1(new_n2601_), .A2(new_n2141_), .ZN(new_n2602_));
  OAI21_X1   g02339(.A1(new_n2592_), .A2(new_n2591_), .B(new_n2397_), .ZN(new_n2603_));
  NAND3_X1   g02340(.A1(new_n2584_), .A2(new_n2589_), .A3(new_n2388_), .ZN(new_n2604_));
  NAND2_X1   g02341(.A1(new_n2603_), .A2(new_n2604_), .ZN(new_n2605_));
  INV_X1     g02342(.I(new_n2598_), .ZN(new_n2606_));
  AOI21_X1   g02343(.A1(new_n2605_), .A2(new_n2606_), .B(new_n2602_), .ZN(new_n2607_));
  INV_X1     g02344(.I(new_n2607_), .ZN(new_n2608_));
  AOI21_X1   g02345(.A1(new_n2608_), .A2(new_n2600_), .B(new_n2474_), .ZN(new_n2609_));
  XOR2_X1    g02346(.A1(new_n2310_), .A2(new_n2389_), .Z(new_n2610_));
  NAND2_X1   g02347(.A1(new_n2610_), .A2(new_n2393_), .ZN(new_n2611_));
  NOR3_X1    g02348(.A1(new_n2607_), .A2(new_n2599_), .A3(new_n2611_), .ZN(new_n2612_));
  OAI22_X1   g02349(.A1(new_n448_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n450_), .ZN(new_n2613_));
  OAI21_X1   g02350(.A1(new_n1518_), .A2(new_n496_), .B(new_n2613_), .ZN(new_n2614_));
  AOI21_X1   g02351(.A1(new_n2614_), .A2(new_n452_), .B(new_n448_), .ZN(new_n2615_));
  XNOR2_X1   g02352(.A1(new_n1638_), .A2(new_n2615_), .ZN(new_n2616_));
  INV_X1     g02353(.I(new_n2616_), .ZN(new_n2617_));
  OAI21_X1   g02354(.A1(new_n2609_), .A2(new_n2612_), .B(new_n2617_), .ZN(new_n2618_));
  INV_X1     g02355(.I(new_n2618_), .ZN(new_n2619_));
  OAI21_X1   g02356(.A1(new_n2263_), .A2(new_n2472_), .B(new_n2619_), .ZN(new_n2620_));
  NOR3_X1    g02357(.A1(new_n2417_), .A2(new_n2409_), .A3(new_n2414_), .ZN(new_n2621_));
  AOI21_X1   g02358(.A1(new_n2410_), .A2(new_n2408_), .B(new_n2415_), .ZN(new_n2622_));
  OAI21_X1   g02359(.A1(new_n2622_), .A2(new_n2621_), .B(new_n2301_), .ZN(new_n2623_));
  NAND2_X1   g02360(.A1(new_n2623_), .A2(new_n2252_), .ZN(new_n2624_));
  NAND3_X1   g02361(.A1(new_n2138_), .A2(new_n2624_), .A3(new_n2618_), .ZN(new_n2625_));
  NAND2_X1   g02362(.A1(new_n2620_), .A2(new_n2625_), .ZN(new_n2626_));
  NAND2_X1   g02363(.A1(new_n2626_), .A2(new_n2418_), .ZN(new_n2627_));
  NAND3_X1   g02364(.A1(new_n2620_), .A2(new_n2625_), .A3(new_n2622_), .ZN(new_n2628_));
  NAND2_X1   g02365(.A1(new_n2627_), .A2(new_n2628_), .ZN(new_n2629_));
  INV_X1     g02366(.I(new_n2629_), .ZN(new_n2630_));
  OAI22_X1   g02367(.A1(new_n1936_), .A2(new_n341_), .B1(new_n404_), .B2(new_n2102_), .ZN(new_n2631_));
  OAI21_X1   g02368(.A1(new_n1803_), .A2(new_n366_), .B(new_n2631_), .ZN(new_n2632_));
  AOI21_X1   g02369(.A1(new_n2632_), .A2(new_n334_), .B(new_n341_), .ZN(new_n2633_));
  XOR2_X1    g02370(.A1(new_n2106_), .A2(new_n2633_), .Z(new_n2634_));
  NOR2_X1    g02371(.A1(new_n2630_), .A2(new_n2634_), .ZN(new_n2635_));
  INV_X1     g02372(.I(new_n2634_), .ZN(new_n2636_));
  NOR2_X1    g02373(.A1(new_n2629_), .A2(new_n2636_), .ZN(new_n2637_));
  OAI21_X1   g02374(.A1(new_n2635_), .A2(new_n2637_), .B(new_n2471_), .ZN(new_n2638_));
  XOR2_X1    g02375(.A1(new_n2629_), .A2(new_n2634_), .Z(new_n2639_));
  OAI21_X1   g02376(.A1(new_n2471_), .A2(new_n2639_), .B(new_n2638_), .ZN(new_n2640_));
  INV_X1     g02377(.I(new_n2640_), .ZN(new_n2641_));
  INV_X1     g02378(.I(new_n2438_), .ZN(new_n2642_));
  INV_X1     g02379(.I(\b[27] ), .ZN(new_n2643_));
  NOR2_X1    g02380(.A1(new_n2643_), .A2(\b[25] ), .ZN(new_n2644_));
  NOR2_X1    g02381(.A1(new_n2281_), .A2(\b[27] ), .ZN(new_n2645_));
  OAI21_X1   g02382(.A1(new_n2644_), .A2(new_n2645_), .B(new_n2642_), .ZN(new_n2646_));
  XOR2_X1    g02383(.A1(new_n2437_), .A2(new_n2646_), .Z(new_n2647_));
  OAI22_X1   g02384(.A1(new_n330_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n263_), .ZN(new_n2648_));
  OAI21_X1   g02385(.A1(new_n2281_), .A2(new_n289_), .B(new_n2648_), .ZN(new_n2649_));
  AOI21_X1   g02386(.A1(new_n2649_), .A2(new_n260_), .B(new_n426_), .ZN(new_n2650_));
  XNOR2_X1   g02387(.A1(new_n2647_), .A2(new_n2650_), .ZN(new_n2651_));
  NOR2_X1    g02388(.A1(new_n2641_), .A2(new_n2651_), .ZN(new_n2652_));
  XOR2_X1    g02389(.A1(new_n2467_), .A2(new_n2652_), .Z(new_n2653_));
  XOR2_X1    g02390(.A1(new_n2653_), .A2(new_n2462_), .Z(\f[27] ));
  NAND3_X1   g02391(.A1(new_n2466_), .A2(new_n2463_), .A3(new_n2640_), .ZN(new_n2655_));
  AOI21_X1   g02392(.A1(new_n2466_), .A2(new_n2463_), .B(new_n2640_), .ZN(new_n2656_));
  NOR2_X1    g02393(.A1(new_n2462_), .A2(new_n2651_), .ZN(new_n2657_));
  INV_X1     g02394(.I(new_n2657_), .ZN(new_n2658_));
  OAI21_X1   g02395(.A1(new_n2656_), .A2(new_n2658_), .B(new_n2655_), .ZN(new_n2659_));
  NOR2_X1    g02396(.A1(new_n2594_), .A2(new_n2611_), .ZN(new_n2660_));
  NOR3_X1    g02397(.A1(new_n2474_), .A2(new_n2590_), .A3(new_n2593_), .ZN(new_n2661_));
  NOR3_X1    g02398(.A1(new_n2661_), .A2(new_n2602_), .A3(new_n2598_), .ZN(new_n2662_));
  NOR2_X1    g02399(.A1(new_n2662_), .A2(new_n2660_), .ZN(new_n2663_));
  NAND2_X1   g02400(.A1(new_n2578_), .A2(new_n2576_), .ZN(new_n2664_));
  NAND2_X1   g02401(.A1(new_n2664_), .A2(new_n2388_), .ZN(new_n2665_));
  INV_X1     g02402(.I(new_n2582_), .ZN(new_n2666_));
  OAI21_X1   g02403(.A1(new_n2664_), .A2(new_n2388_), .B(new_n2666_), .ZN(new_n2667_));
  OAI21_X1   g02404(.A1(new_n2481_), .A2(new_n2667_), .B(new_n2665_), .ZN(new_n2668_));
  INV_X1     g02405(.I(new_n2552_), .ZN(new_n2669_));
  OAI21_X1   g02406(.A1(new_n2492_), .A2(new_n2552_), .B(new_n2557_), .ZN(new_n2670_));
  OAI22_X1   g02407(.A1(new_n2560_), .A2(new_n2670_), .B1(new_n2669_), .B2(new_n2493_), .ZN(new_n2671_));
  NOR2_X1    g02408(.A1(new_n2546_), .A2(new_n2547_), .ZN(new_n2672_));
  AOI21_X1   g02409(.A1(new_n2327_), .A2(new_n2509_), .B(new_n2508_), .ZN(new_n2673_));
  NOR3_X1    g02410(.A1(new_n2519_), .A2(new_n2524_), .A3(new_n2317_), .ZN(new_n2674_));
  OAI21_X1   g02411(.A1(new_n2673_), .A2(new_n2674_), .B(new_n2499_), .ZN(new_n2675_));
  OAI21_X1   g02412(.A1(new_n2519_), .A2(new_n2317_), .B(new_n2524_), .ZN(new_n2676_));
  INV_X1     g02413(.I(new_n2674_), .ZN(new_n2677_));
  NAND3_X1   g02414(.A1(new_n2677_), .A2(new_n2676_), .A3(new_n2500_), .ZN(new_n2678_));
  AOI22_X1   g02415(.A1(new_n2678_), .A2(new_n2675_), .B1(new_n2515_), .B2(new_n2516_), .ZN(new_n2679_));
  OAI21_X1   g02416(.A1(new_n2531_), .A2(new_n2528_), .B(new_n2679_), .ZN(new_n2680_));
  NAND2_X1   g02417(.A1(new_n2680_), .A2(new_n2534_), .ZN(new_n2681_));
  NAND2_X1   g02418(.A1(new_n2681_), .A2(new_n2672_), .ZN(new_n2682_));
  NOR2_X1    g02419(.A1(new_n2327_), .A2(new_n2508_), .ZN(new_n2683_));
  NAND4_X1   g02420(.A1(new_n2175_), .A2(new_n2176_), .A3(new_n2178_), .A4(new_n2500_), .ZN(new_n2684_));
  AOI21_X1   g02421(.A1(new_n2327_), .A2(new_n2508_), .B(new_n2684_), .ZN(new_n2685_));
  NOR2_X1    g02422(.A1(new_n2685_), .A2(new_n2683_), .ZN(new_n2686_));
  INV_X1     g02423(.I(new_n2686_), .ZN(new_n2687_));
  OAI22_X1   g02424(.A1(new_n2171_), .A2(new_n298_), .B1(new_n325_), .B2(new_n2166_), .ZN(new_n2688_));
  OAI21_X1   g02425(.A1(new_n280_), .A2(new_n2322_), .B(new_n2688_), .ZN(new_n2689_));
  AOI21_X1   g02426(.A1(new_n2689_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n2690_));
  XOR2_X1    g02427(.A1(new_n2690_), .A2(new_n329_), .Z(new_n2691_));
  XNOR2_X1   g02428(.A1(\a[27] ), .A2(\a[29] ), .ZN(new_n2692_));
  XNOR2_X1   g02429(.A1(\a[26] ), .A2(\a[28] ), .ZN(new_n2693_));
  NOR2_X1    g02430(.A1(new_n2693_), .A2(new_n2692_), .ZN(new_n2694_));
  INV_X1     g02431(.I(\a[27] ), .ZN(new_n2695_));
  NAND3_X1   g02432(.A1(new_n2168_), .A2(new_n2695_), .A3(\a[28] ), .ZN(new_n2696_));
  INV_X1     g02433(.I(\a[28] ), .ZN(new_n2697_));
  NAND3_X1   g02434(.A1(new_n2697_), .A2(\a[26] ), .A3(\a[27] ), .ZN(new_n2698_));
  NAND2_X1   g02435(.A1(new_n2696_), .A2(new_n2698_), .ZN(new_n2699_));
  INV_X1     g02436(.I(new_n2699_), .ZN(new_n2700_));
  NOR2_X1    g02437(.A1(new_n2700_), .A2(new_n269_), .ZN(new_n2701_));
  INV_X1     g02438(.I(\a[29] ), .ZN(new_n2702_));
  XOR2_X1    g02439(.A1(\a[27] ), .A2(\a[29] ), .Z(new_n2703_));
  XOR2_X1    g02440(.A1(\a[26] ), .A2(\a[28] ), .Z(new_n2704_));
  NAND2_X1   g02441(.A1(new_n2704_), .A2(new_n2703_), .ZN(new_n2705_));
  OAI21_X1   g02442(.A1(new_n2705_), .A2(new_n258_), .B(new_n2702_), .ZN(new_n2706_));
  OAI21_X1   g02443(.A1(new_n2706_), .A2(new_n2701_), .B(new_n2694_), .ZN(new_n2707_));
  NOR2_X1    g02444(.A1(new_n2707_), .A2(new_n271_), .ZN(new_n2708_));
  NAND2_X1   g02445(.A1(new_n2707_), .A2(new_n271_), .ZN(new_n2709_));
  INV_X1     g02446(.I(new_n2709_), .ZN(new_n2710_));
  NOR2_X1    g02447(.A1(new_n2500_), .A2(new_n2702_), .ZN(new_n2711_));
  NOR3_X1    g02448(.A1(new_n2710_), .A2(new_n2708_), .A3(new_n2711_), .ZN(new_n2712_));
  INV_X1     g02449(.I(new_n2708_), .ZN(new_n2713_));
  INV_X1     g02450(.I(new_n2711_), .ZN(new_n2714_));
  AOI21_X1   g02451(.A1(new_n2713_), .A2(new_n2709_), .B(new_n2714_), .ZN(new_n2715_));
  NOR2_X1    g02452(.A1(new_n2715_), .A2(new_n2712_), .ZN(new_n2716_));
  XOR2_X1    g02453(.A1(new_n2716_), .A2(new_n2691_), .Z(new_n2717_));
  NAND2_X1   g02454(.A1(new_n2687_), .A2(new_n2717_), .ZN(new_n2718_));
  NOR2_X1    g02455(.A1(new_n2716_), .A2(new_n2691_), .ZN(new_n2719_));
  XOR2_X1    g02456(.A1(new_n2690_), .A2(new_n807_), .Z(new_n2720_));
  INV_X1     g02457(.I(new_n2716_), .ZN(new_n2721_));
  NOR2_X1    g02458(.A1(new_n2721_), .A2(new_n2720_), .ZN(new_n2722_));
  OAI21_X1   g02459(.A1(new_n2719_), .A2(new_n2722_), .B(new_n2686_), .ZN(new_n2723_));
  NAND2_X1   g02460(.A1(new_n2718_), .A2(new_n2723_), .ZN(new_n2724_));
  INV_X1     g02461(.I(new_n1707_), .ZN(new_n2725_));
  AOI22_X1   g02462(.A1(\b[7] ), .A2(new_n2725_), .B1(new_n1702_), .B2(\b[6] ), .ZN(new_n2726_));
  AOI21_X1   g02463(.A1(\b[5] ), .A2(new_n1851_), .B(new_n2726_), .ZN(new_n2727_));
  OAI21_X1   g02464(.A1(new_n2727_), .A2(\a[23] ), .B(new_n1702_), .ZN(new_n2728_));
  XNOR2_X1   g02465(.A1(new_n471_), .A2(new_n2728_), .ZN(new_n2729_));
  INV_X1     g02466(.I(new_n2729_), .ZN(new_n2730_));
  NAND2_X1   g02467(.A1(new_n2724_), .A2(new_n2730_), .ZN(new_n2731_));
  INV_X1     g02468(.I(new_n2724_), .ZN(new_n2732_));
  NAND2_X1   g02469(.A1(new_n2732_), .A2(new_n2729_), .ZN(new_n2733_));
  AOI21_X1   g02470(.A1(new_n2731_), .A2(new_n2733_), .B(new_n2682_), .ZN(new_n2734_));
  NAND3_X1   g02471(.A1(new_n2718_), .A2(new_n2723_), .A3(new_n2730_), .ZN(new_n2735_));
  NAND2_X1   g02472(.A1(new_n2724_), .A2(new_n2729_), .ZN(new_n2736_));
  AOI22_X1   g02473(.A1(new_n2672_), .A2(new_n2681_), .B1(new_n2736_), .B2(new_n2735_), .ZN(new_n2737_));
  NOR2_X1    g02474(.A1(new_n2734_), .A2(new_n2737_), .ZN(new_n2738_));
  INV_X1     g02475(.I(new_n2738_), .ZN(new_n2739_));
  OAI22_X1   g02476(.A1(new_n1347_), .A2(new_n565_), .B1(new_n656_), .B2(new_n1344_), .ZN(new_n2740_));
  OAI21_X1   g02477(.A1(new_n515_), .A2(new_n1457_), .B(new_n2740_), .ZN(new_n2741_));
  AOI21_X1   g02478(.A1(new_n2741_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n2742_));
  XNOR2_X1   g02479(.A1(new_n660_), .A2(new_n2742_), .ZN(new_n2743_));
  INV_X1     g02480(.I(new_n2743_), .ZN(new_n2744_));
  NAND2_X1   g02481(.A1(new_n2739_), .A2(new_n2744_), .ZN(new_n2745_));
  NAND2_X1   g02482(.A1(new_n2738_), .A2(new_n2743_), .ZN(new_n2746_));
  NAND2_X1   g02483(.A1(new_n2745_), .A2(new_n2746_), .ZN(new_n2747_));
  NAND2_X1   g02484(.A1(new_n2671_), .A2(new_n2747_), .ZN(new_n2748_));
  INV_X1     g02485(.I(new_n2671_), .ZN(new_n2749_));
  AOI21_X1   g02486(.A1(new_n2534_), .A2(new_n2680_), .B(new_n2548_), .ZN(new_n2750_));
  NAND2_X1   g02487(.A1(new_n2733_), .A2(new_n2731_), .ZN(new_n2751_));
  NAND2_X1   g02488(.A1(new_n2750_), .A2(new_n2751_), .ZN(new_n2752_));
  INV_X1     g02489(.I(new_n2737_), .ZN(new_n2753_));
  NAND3_X1   g02490(.A1(new_n2752_), .A2(new_n2753_), .A3(new_n2744_), .ZN(new_n2754_));
  OAI21_X1   g02491(.A1(new_n2734_), .A2(new_n2737_), .B(new_n2743_), .ZN(new_n2755_));
  NAND2_X1   g02492(.A1(new_n2754_), .A2(new_n2755_), .ZN(new_n2756_));
  NAND2_X1   g02493(.A1(new_n2749_), .A2(new_n2756_), .ZN(new_n2757_));
  OAI22_X1   g02494(.A1(new_n1055_), .A2(new_n780_), .B1(new_n861_), .B2(new_n1061_), .ZN(new_n2758_));
  OAI21_X1   g02495(.A1(new_n706_), .A2(new_n1332_), .B(new_n2758_), .ZN(new_n2759_));
  AOI21_X1   g02496(.A1(new_n2759_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n2760_));
  XNOR2_X1   g02497(.A1(new_n860_), .A2(new_n2760_), .ZN(new_n2761_));
  INV_X1     g02498(.I(new_n2761_), .ZN(new_n2762_));
  NAND3_X1   g02499(.A1(new_n2757_), .A2(new_n2748_), .A3(new_n2762_), .ZN(new_n2763_));
  NAND2_X1   g02500(.A1(new_n2757_), .A2(new_n2748_), .ZN(new_n2764_));
  NAND2_X1   g02501(.A1(new_n2764_), .A2(new_n2761_), .ZN(new_n2765_));
  NAND2_X1   g02502(.A1(new_n2765_), .A2(new_n2763_), .ZN(new_n2766_));
  INV_X1     g02503(.I(new_n2766_), .ZN(new_n2767_));
  NAND2_X1   g02504(.A1(new_n2567_), .A2(new_n2482_), .ZN(new_n2768_));
  OAI21_X1   g02505(.A1(new_n2567_), .A2(new_n2482_), .B(new_n2572_), .ZN(new_n2769_));
  OAI21_X1   g02506(.A1(new_n2487_), .A2(new_n2769_), .B(new_n2768_), .ZN(new_n2770_));
  OAI22_X1   g02507(.A1(new_n970_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n820_), .ZN(new_n2771_));
  OAI21_X1   g02508(.A1(new_n930_), .A2(new_n894_), .B(new_n2771_), .ZN(new_n2772_));
  AOI21_X1   g02509(.A1(new_n2772_), .A2(new_n827_), .B(new_n970_), .ZN(new_n2773_));
  XOR2_X1    g02510(.A1(new_n1114_), .A2(new_n2773_), .Z(new_n2774_));
  INV_X1     g02511(.I(new_n2774_), .ZN(new_n2775_));
  XOR2_X1    g02512(.A1(new_n2770_), .A2(new_n2775_), .Z(new_n2776_));
  NOR2_X1    g02513(.A1(new_n2776_), .A2(new_n2767_), .ZN(new_n2777_));
  INV_X1     g02514(.I(new_n2770_), .ZN(new_n2778_));
  NAND2_X1   g02515(.A1(new_n2778_), .A2(new_n2775_), .ZN(new_n2779_));
  NAND2_X1   g02516(.A1(new_n2770_), .A2(new_n2774_), .ZN(new_n2780_));
  AOI21_X1   g02517(.A1(new_n2779_), .A2(new_n2780_), .B(new_n2766_), .ZN(new_n2781_));
  NOR2_X1    g02518(.A1(new_n2777_), .A2(new_n2781_), .ZN(new_n2782_));
  OAI22_X1   g02519(.A1(new_n607_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n610_), .ZN(new_n2783_));
  OAI21_X1   g02520(.A1(new_n1189_), .A2(new_n684_), .B(new_n2783_), .ZN(new_n2784_));
  AOI21_X1   g02521(.A1(new_n2784_), .A2(new_n612_), .B(new_n607_), .ZN(new_n2785_));
  XNOR2_X1   g02522(.A1(new_n1421_), .A2(new_n2785_), .ZN(new_n2786_));
  INV_X1     g02523(.I(new_n2786_), .ZN(new_n2787_));
  XOR2_X1    g02524(.A1(new_n2782_), .A2(new_n2787_), .Z(new_n2788_));
  NAND2_X1   g02525(.A1(new_n2788_), .A2(new_n2668_), .ZN(new_n2789_));
  NAND2_X1   g02526(.A1(new_n2782_), .A2(new_n2787_), .ZN(new_n2790_));
  INV_X1     g02527(.I(new_n2782_), .ZN(new_n2791_));
  NAND2_X1   g02528(.A1(new_n2791_), .A2(new_n2786_), .ZN(new_n2792_));
  AOI21_X1   g02529(.A1(new_n2792_), .A2(new_n2790_), .B(new_n2668_), .ZN(new_n2793_));
  INV_X1     g02530(.I(new_n2793_), .ZN(new_n2794_));
  NAND2_X1   g02531(.A1(new_n2794_), .A2(new_n2789_), .ZN(new_n2795_));
  XOR2_X1    g02532(.A1(new_n2663_), .A2(new_n2795_), .Z(new_n2796_));
  OAI22_X1   g02533(.A1(new_n448_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n450_), .ZN(new_n2797_));
  OAI21_X1   g02534(.A1(new_n1525_), .A2(new_n496_), .B(new_n2797_), .ZN(new_n2798_));
  AOI21_X1   g02535(.A1(new_n2798_), .A2(new_n452_), .B(new_n448_), .ZN(new_n2799_));
  XOR2_X1    g02536(.A1(new_n1808_), .A2(new_n2799_), .Z(new_n2800_));
  NOR2_X1    g02537(.A1(new_n2796_), .A2(new_n2800_), .ZN(new_n2801_));
  INV_X1     g02538(.I(new_n2801_), .ZN(new_n2802_));
  NAND2_X1   g02539(.A1(new_n2796_), .A2(new_n2800_), .ZN(new_n2803_));
  NAND2_X1   g02540(.A1(new_n2802_), .A2(new_n2803_), .ZN(new_n2804_));
  INV_X1     g02541(.I(new_n2804_), .ZN(new_n2805_));
  INV_X1     g02542(.I(new_n2609_), .ZN(new_n2806_));
  INV_X1     g02543(.I(new_n2612_), .ZN(new_n2807_));
  AOI21_X1   g02544(.A1(new_n2806_), .A2(new_n2807_), .B(new_n2418_), .ZN(new_n2808_));
  NOR3_X1    g02545(.A1(new_n2609_), .A2(new_n2612_), .A3(new_n2622_), .ZN(new_n2809_));
  INV_X1     g02546(.I(new_n2809_), .ZN(new_n2810_));
  NOR3_X1    g02547(.A1(new_n2263_), .A2(new_n2472_), .A3(new_n2616_), .ZN(new_n2811_));
  AOI21_X1   g02548(.A1(new_n2811_), .A2(new_n2810_), .B(new_n2808_), .ZN(new_n2812_));
  OAI22_X1   g02549(.A1(new_n2102_), .A2(new_n341_), .B1(new_n404_), .B2(new_n2281_), .ZN(new_n2813_));
  OAI21_X1   g02550(.A1(new_n1936_), .A2(new_n366_), .B(new_n2813_), .ZN(new_n2814_));
  AOI21_X1   g02551(.A1(new_n2814_), .A2(new_n334_), .B(new_n341_), .ZN(new_n2815_));
  XNOR2_X1   g02552(.A1(new_n2280_), .A2(new_n2815_), .ZN(new_n2816_));
  INV_X1     g02553(.I(new_n2816_), .ZN(new_n2817_));
  NAND2_X1   g02554(.A1(new_n2812_), .A2(new_n2817_), .ZN(new_n2818_));
  INV_X1     g02555(.I(new_n2808_), .ZN(new_n2819_));
  NAND3_X1   g02556(.A1(new_n2138_), .A2(new_n2624_), .A3(new_n2617_), .ZN(new_n2820_));
  OAI21_X1   g02557(.A1(new_n2820_), .A2(new_n2809_), .B(new_n2819_), .ZN(new_n2821_));
  NAND2_X1   g02558(.A1(new_n2821_), .A2(new_n2816_), .ZN(new_n2822_));
  AOI21_X1   g02559(.A1(new_n2818_), .A2(new_n2822_), .B(new_n2805_), .ZN(new_n2823_));
  NAND2_X1   g02560(.A1(new_n2821_), .A2(new_n2817_), .ZN(new_n2824_));
  NAND2_X1   g02561(.A1(new_n2812_), .A2(new_n2816_), .ZN(new_n2825_));
  AOI21_X1   g02562(.A1(new_n2825_), .A2(new_n2824_), .B(new_n2804_), .ZN(new_n2826_));
  NOR2_X1    g02563(.A1(new_n2823_), .A2(new_n2826_), .ZN(new_n2827_));
  NOR3_X1    g02564(.A1(new_n2639_), .A2(new_n2635_), .A3(new_n2827_), .ZN(new_n2828_));
  NOR2_X1    g02565(.A1(new_n2630_), .A2(new_n2634_), .ZN(new_n2829_));
  OAI21_X1   g02566(.A1(new_n2828_), .A2(new_n2829_), .B(new_n2470_), .ZN(new_n2830_));
  INV_X1     g02567(.I(new_n2830_), .ZN(new_n2831_));
  NOR3_X1    g02568(.A1(new_n2828_), .A2(new_n2470_), .A3(new_n2829_), .ZN(new_n2832_));
  NOR2_X1    g02569(.A1(new_n2831_), .A2(new_n2832_), .ZN(new_n2833_));
  INV_X1     g02570(.I(new_n2833_), .ZN(new_n2834_));
  NOR2_X1    g02571(.A1(\b[26] ), .A2(\b[27] ), .ZN(new_n2835_));
  AOI21_X1   g02572(.A1(new_n2437_), .A2(new_n2835_), .B(new_n2281_), .ZN(new_n2836_));
  NOR2_X1    g02573(.A1(new_n2439_), .A2(new_n2643_), .ZN(new_n2837_));
  INV_X1     g02574(.I(new_n2837_), .ZN(new_n2838_));
  NOR2_X1    g02575(.A1(new_n2437_), .A2(new_n2838_), .ZN(new_n2839_));
  NOR2_X1    g02576(.A1(new_n2836_), .A2(new_n2839_), .ZN(new_n2840_));
  XNOR2_X1   g02577(.A1(\b[27] ), .A2(\b[28] ), .ZN(new_n2841_));
  INV_X1     g02578(.I(\b[28] ), .ZN(new_n2842_));
  NOR2_X1    g02579(.A1(new_n2643_), .A2(new_n2842_), .ZN(new_n2843_));
  NOR2_X1    g02580(.A1(\b[27] ), .A2(\b[28] ), .ZN(new_n2844_));
  OAI21_X1   g02581(.A1(new_n2843_), .A2(new_n2844_), .B(new_n2840_), .ZN(new_n2845_));
  OAI21_X1   g02582(.A1(new_n2840_), .A2(new_n2841_), .B(new_n2845_), .ZN(new_n2846_));
  OAI22_X1   g02583(.A1(new_n330_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n263_), .ZN(new_n2847_));
  OAI21_X1   g02584(.A1(new_n2439_), .A2(new_n289_), .B(new_n2847_), .ZN(new_n2848_));
  AOI21_X1   g02585(.A1(new_n2848_), .A2(new_n260_), .B(new_n426_), .ZN(new_n2849_));
  XNOR2_X1   g02586(.A1(new_n2846_), .A2(new_n2849_), .ZN(new_n2850_));
  INV_X1     g02587(.I(new_n2850_), .ZN(new_n2851_));
  NAND2_X1   g02588(.A1(new_n2834_), .A2(new_n2851_), .ZN(new_n2852_));
  NAND2_X1   g02589(.A1(new_n2833_), .A2(new_n2850_), .ZN(new_n2853_));
  NAND2_X1   g02590(.A1(new_n2852_), .A2(new_n2853_), .ZN(new_n2854_));
  NAND2_X1   g02591(.A1(new_n2659_), .A2(new_n2854_), .ZN(new_n2855_));
  XOR2_X1    g02592(.A1(new_n2833_), .A2(new_n2851_), .Z(new_n2856_));
  OAI21_X1   g02593(.A1(new_n2659_), .A2(new_n2856_), .B(new_n2855_), .ZN(\f[28] ));
  XOR2_X1    g02594(.A1(new_n2821_), .A2(new_n2804_), .Z(new_n2858_));
  NOR2_X1    g02595(.A1(new_n2858_), .A2(new_n2817_), .ZN(new_n2859_));
  OAI21_X1   g02596(.A1(new_n2827_), .A2(new_n2630_), .B(new_n2634_), .ZN(new_n2860_));
  INV_X1     g02597(.I(new_n2860_), .ZN(new_n2861_));
  NOR3_X1    g02598(.A1(new_n2823_), .A2(new_n2826_), .A3(new_n2629_), .ZN(new_n2862_));
  NOR2_X1    g02599(.A1(new_n2470_), .A2(new_n2862_), .ZN(new_n2863_));
  INV_X1     g02600(.I(new_n2863_), .ZN(new_n2864_));
  NOR2_X1    g02601(.A1(new_n2864_), .A2(new_n2861_), .ZN(new_n2865_));
  OAI22_X1   g02602(.A1(new_n607_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n610_), .ZN(new_n2866_));
  OAI21_X1   g02603(.A1(new_n1294_), .A2(new_n684_), .B(new_n2866_), .ZN(new_n2867_));
  AOI21_X1   g02604(.A1(new_n2867_), .A2(new_n612_), .B(new_n607_), .ZN(new_n2868_));
  XOR2_X1    g02605(.A1(new_n1530_), .A2(new_n2868_), .Z(new_n2869_));
  INV_X1     g02606(.I(new_n2668_), .ZN(new_n2870_));
  XNOR2_X1   g02607(.A1(new_n2766_), .A2(new_n2770_), .ZN(new_n2871_));
  NOR2_X1    g02608(.A1(new_n2871_), .A2(new_n2775_), .ZN(new_n2872_));
  INV_X1     g02609(.I(new_n2872_), .ZN(new_n2873_));
  NAND2_X1   g02610(.A1(new_n2764_), .A2(new_n2762_), .ZN(new_n2874_));
  NAND2_X1   g02611(.A1(new_n2736_), .A2(new_n2735_), .ZN(new_n2875_));
  OAI22_X1   g02612(.A1(new_n1712_), .A2(new_n472_), .B1(new_n515_), .B2(new_n1707_), .ZN(new_n2876_));
  OAI21_X1   g02613(.A1(new_n420_), .A2(new_n1850_), .B(new_n2876_), .ZN(new_n2877_));
  AOI21_X1   g02614(.A1(new_n2877_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n2878_));
  XOR2_X1    g02615(.A1(new_n700_), .A2(new_n2878_), .Z(new_n2879_));
  NAND3_X1   g02616(.A1(new_n2713_), .A2(new_n2709_), .A3(new_n2711_), .ZN(new_n2880_));
  OAI21_X1   g02617(.A1(\b[1] ), .A2(new_n282_), .B(new_n2694_), .ZN(new_n2881_));
  OAI21_X1   g02618(.A1(new_n280_), .A2(new_n2700_), .B(new_n2881_), .ZN(new_n2882_));
  XOR2_X1    g02619(.A1(\a[26] ), .A2(\a[29] ), .Z(new_n2883_));
  NAND3_X1   g02620(.A1(new_n2704_), .A2(new_n2498_), .A3(new_n2883_), .ZN(new_n2884_));
  NOR2_X1    g02621(.A1(new_n2884_), .A2(new_n258_), .ZN(new_n2885_));
  AOI21_X1   g02622(.A1(new_n2882_), .A2(new_n2885_), .B(new_n2702_), .ZN(new_n2886_));
  NAND3_X1   g02623(.A1(new_n2882_), .A2(new_n2702_), .A3(new_n2885_), .ZN(new_n2887_));
  INV_X1     g02624(.I(new_n2887_), .ZN(new_n2888_));
  NOR2_X1    g02625(.A1(new_n2888_), .A2(new_n2886_), .ZN(new_n2889_));
  XOR2_X1    g02626(.A1(new_n2889_), .A2(new_n2880_), .Z(new_n2890_));
  INV_X1     g02627(.I(new_n2890_), .ZN(new_n2891_));
  INV_X1     g02628(.I(new_n2722_), .ZN(new_n2892_));
  OAI22_X1   g02629(.A1(new_n2685_), .A2(new_n2683_), .B1(new_n2691_), .B2(new_n2716_), .ZN(new_n2893_));
  NAND2_X1   g02630(.A1(new_n378_), .A2(new_n2161_), .ZN(new_n2894_));
  INV_X1     g02631(.I(new_n2322_), .ZN(new_n2895_));
  INV_X1     g02632(.I(new_n2166_), .ZN(new_n2896_));
  AOI22_X1   g02633(.A1(new_n2161_), .A2(\b[4] ), .B1(\b[5] ), .B2(new_n2896_), .ZN(new_n2897_));
  AOI21_X1   g02634(.A1(\b[3] ), .A2(new_n2895_), .B(new_n2897_), .ZN(new_n2898_));
  NAND2_X1   g02635(.A1(new_n2898_), .A2(new_n2894_), .ZN(new_n2899_));
  XOR2_X1    g02636(.A1(new_n2899_), .A2(\a[26] ), .Z(new_n2900_));
  INV_X1     g02637(.I(new_n2900_), .ZN(new_n2901_));
  NAND3_X1   g02638(.A1(new_n2893_), .A2(new_n2892_), .A3(new_n2901_), .ZN(new_n2902_));
  NAND2_X1   g02639(.A1(new_n2519_), .A2(new_n2524_), .ZN(new_n2903_));
  NOR2_X1    g02640(.A1(new_n2317_), .A2(new_n2499_), .ZN(new_n2904_));
  OAI21_X1   g02641(.A1(new_n2519_), .A2(new_n2524_), .B(new_n2904_), .ZN(new_n2905_));
  AOI21_X1   g02642(.A1(new_n2903_), .A2(new_n2905_), .B(new_n2719_), .ZN(new_n2906_));
  OAI21_X1   g02643(.A1(new_n2906_), .A2(new_n2722_), .B(new_n2900_), .ZN(new_n2907_));
  AOI21_X1   g02644(.A1(new_n2902_), .A2(new_n2907_), .B(new_n2891_), .ZN(new_n2908_));
  NOR3_X1    g02645(.A1(new_n2906_), .A2(new_n2722_), .A3(new_n2900_), .ZN(new_n2909_));
  AOI21_X1   g02646(.A1(new_n2893_), .A2(new_n2892_), .B(new_n2901_), .ZN(new_n2910_));
  NOR3_X1    g02647(.A1(new_n2910_), .A2(new_n2909_), .A3(new_n2890_), .ZN(new_n2911_));
  OAI21_X1   g02648(.A1(new_n2908_), .A2(new_n2911_), .B(new_n2879_), .ZN(new_n2912_));
  INV_X1     g02649(.I(new_n2879_), .ZN(new_n2913_));
  OAI21_X1   g02650(.A1(new_n2910_), .A2(new_n2909_), .B(new_n2890_), .ZN(new_n2914_));
  NAND3_X1   g02651(.A1(new_n2902_), .A2(new_n2907_), .A3(new_n2891_), .ZN(new_n2915_));
  NAND3_X1   g02652(.A1(new_n2914_), .A2(new_n2915_), .A3(new_n2913_), .ZN(new_n2916_));
  NAND2_X1   g02653(.A1(new_n2912_), .A2(new_n2916_), .ZN(new_n2917_));
  NAND3_X1   g02654(.A1(new_n2917_), .A2(new_n2875_), .A3(new_n2731_), .ZN(new_n2918_));
  INV_X1     g02655(.I(new_n2918_), .ZN(new_n2919_));
  NOR2_X1    g02656(.A1(new_n2732_), .A2(new_n2729_), .ZN(new_n2921_));
  OAI21_X1   g02657(.A1(new_n2919_), .A2(new_n2921_), .B(new_n2682_), .ZN(new_n2922_));
  INV_X1     g02658(.I(new_n2921_), .ZN(new_n2923_));
  NAND3_X1   g02659(.A1(new_n2918_), .A2(new_n2750_), .A3(new_n2923_), .ZN(new_n2924_));
  OAI22_X1   g02660(.A1(new_n1347_), .A2(new_n656_), .B1(new_n706_), .B2(new_n1344_), .ZN(new_n2925_));
  OAI21_X1   g02661(.A1(new_n565_), .A2(new_n1457_), .B(new_n2925_), .ZN(new_n2926_));
  AOI21_X1   g02662(.A1(new_n2926_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n2927_));
  XNOR2_X1   g02663(.A1(new_n710_), .A2(new_n2927_), .ZN(new_n2928_));
  AOI21_X1   g02664(.A1(new_n2922_), .A2(new_n2924_), .B(new_n2928_), .ZN(new_n2929_));
  AOI21_X1   g02665(.A1(new_n2918_), .A2(new_n2923_), .B(new_n2750_), .ZN(new_n2930_));
  INV_X1     g02666(.I(new_n2924_), .ZN(new_n2931_));
  INV_X1     g02667(.I(new_n2928_), .ZN(new_n2932_));
  NOR3_X1    g02668(.A1(new_n2931_), .A2(new_n2930_), .A3(new_n2932_), .ZN(new_n2933_));
  OAI21_X1   g02669(.A1(new_n2933_), .A2(new_n2929_), .B(new_n2756_), .ZN(new_n2934_));
  AOI21_X1   g02670(.A1(new_n2739_), .A2(new_n2744_), .B(new_n2934_), .ZN(new_n2935_));
  OAI21_X1   g02671(.A1(new_n2931_), .A2(new_n2930_), .B(new_n2932_), .ZN(new_n2936_));
  NAND3_X1   g02672(.A1(new_n2922_), .A2(new_n2924_), .A3(new_n2928_), .ZN(new_n2937_));
  NAND2_X1   g02673(.A1(new_n2936_), .A2(new_n2937_), .ZN(new_n2938_));
  NAND2_X1   g02674(.A1(new_n2739_), .A2(new_n2744_), .ZN(new_n2940_));
  INV_X1     g02675(.I(new_n2940_), .ZN(new_n2941_));
  OAI21_X1   g02676(.A1(new_n2935_), .A2(new_n2941_), .B(new_n2749_), .ZN(new_n2942_));
  NAND3_X1   g02677(.A1(new_n2938_), .A2(new_n2745_), .A3(new_n2756_), .ZN(new_n2943_));
  NAND3_X1   g02678(.A1(new_n2943_), .A2(new_n2671_), .A3(new_n2940_), .ZN(new_n2944_));
  OAI22_X1   g02679(.A1(new_n1055_), .A2(new_n861_), .B1(new_n930_), .B2(new_n1061_), .ZN(new_n2945_));
  OAI21_X1   g02680(.A1(new_n780_), .A2(new_n1332_), .B(new_n2945_), .ZN(new_n2946_));
  AOI21_X1   g02681(.A1(new_n2946_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n2947_));
  XNOR2_X1   g02682(.A1(new_n937_), .A2(new_n2947_), .ZN(new_n2948_));
  INV_X1     g02683(.I(new_n2948_), .ZN(new_n2949_));
  NAND3_X1   g02684(.A1(new_n2942_), .A2(new_n2944_), .A3(new_n2949_), .ZN(new_n2950_));
  AOI21_X1   g02685(.A1(new_n2943_), .A2(new_n2940_), .B(new_n2671_), .ZN(new_n2951_));
  INV_X1     g02686(.I(new_n2944_), .ZN(new_n2952_));
  OAI21_X1   g02687(.A1(new_n2952_), .A2(new_n2951_), .B(new_n2948_), .ZN(new_n2953_));
  NAND2_X1   g02688(.A1(new_n2953_), .A2(new_n2950_), .ZN(new_n2954_));
  NAND3_X1   g02689(.A1(new_n2766_), .A2(new_n2954_), .A3(new_n2874_), .ZN(new_n2955_));
  NAND2_X1   g02690(.A1(new_n2764_), .A2(new_n2762_), .ZN(new_n2957_));
  AOI21_X1   g02691(.A1(new_n2955_), .A2(new_n2957_), .B(new_n2770_), .ZN(new_n2958_));
  INV_X1     g02692(.I(new_n2958_), .ZN(new_n2959_));
  NAND3_X1   g02693(.A1(new_n2955_), .A2(new_n2770_), .A3(new_n2957_), .ZN(new_n2960_));
  OAI22_X1   g02694(.A1(new_n970_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n820_), .ZN(new_n2961_));
  OAI21_X1   g02695(.A1(new_n1017_), .A2(new_n894_), .B(new_n2961_), .ZN(new_n2962_));
  AOI21_X1   g02696(.A1(new_n2962_), .A2(new_n827_), .B(new_n970_), .ZN(new_n2963_));
  XNOR2_X1   g02697(.A1(new_n1196_), .A2(new_n2963_), .ZN(new_n2964_));
  INV_X1     g02698(.I(new_n2964_), .ZN(new_n2965_));
  NAND3_X1   g02699(.A1(new_n2959_), .A2(new_n2960_), .A3(new_n2965_), .ZN(new_n2966_));
  INV_X1     g02700(.I(new_n2960_), .ZN(new_n2967_));
  OAI21_X1   g02701(.A1(new_n2967_), .A2(new_n2958_), .B(new_n2964_), .ZN(new_n2968_));
  NAND3_X1   g02702(.A1(new_n2873_), .A2(new_n2966_), .A3(new_n2968_), .ZN(new_n2969_));
  NAND3_X1   g02703(.A1(new_n2870_), .A2(new_n2791_), .A3(new_n2969_), .ZN(new_n2970_));
  NAND2_X1   g02704(.A1(new_n2969_), .A2(new_n2791_), .ZN(new_n2971_));
  NAND2_X1   g02705(.A1(new_n2971_), .A2(new_n2668_), .ZN(new_n2972_));
  NAND2_X1   g02706(.A1(new_n2970_), .A2(new_n2972_), .ZN(new_n2973_));
  XOR2_X1    g02707(.A1(new_n2668_), .A2(new_n2782_), .Z(new_n2974_));
  NOR2_X1    g02708(.A1(new_n2974_), .A2(new_n2787_), .ZN(new_n2975_));
  NOR3_X1    g02709(.A1(new_n2662_), .A2(new_n2660_), .A3(new_n2795_), .ZN(new_n2976_));
  OAI22_X1   g02710(.A1(new_n448_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n450_), .ZN(new_n2977_));
  OAI21_X1   g02711(.A1(new_n1634_), .A2(new_n496_), .B(new_n2977_), .ZN(new_n2978_));
  AOI21_X1   g02712(.A1(new_n2978_), .A2(new_n452_), .B(new_n448_), .ZN(new_n2979_));
  XNOR2_X1   g02713(.A1(new_n1940_), .A2(new_n2979_), .ZN(new_n2980_));
  INV_X1     g02714(.I(new_n2980_), .ZN(new_n2981_));
  OAI21_X1   g02715(.A1(new_n2976_), .A2(new_n2975_), .B(new_n2981_), .ZN(new_n2982_));
  INV_X1     g02716(.I(new_n2975_), .ZN(new_n2983_));
  NAND2_X1   g02717(.A1(new_n2605_), .A2(new_n2474_), .ZN(new_n2984_));
  NAND3_X1   g02718(.A1(new_n2611_), .A2(new_n2603_), .A3(new_n2604_), .ZN(new_n2985_));
  NAND3_X1   g02719(.A1(new_n2478_), .A2(new_n2985_), .A3(new_n2606_), .ZN(new_n2986_));
  AOI21_X1   g02720(.A1(new_n2668_), .A2(new_n2788_), .B(new_n2793_), .ZN(new_n2987_));
  NAND3_X1   g02721(.A1(new_n2986_), .A2(new_n2984_), .A3(new_n2987_), .ZN(new_n2988_));
  NAND3_X1   g02722(.A1(new_n2988_), .A2(new_n2983_), .A3(new_n2980_), .ZN(new_n2989_));
  AOI21_X1   g02723(.A1(new_n2982_), .A2(new_n2989_), .B(new_n2973_), .ZN(new_n2990_));
  XOR2_X1    g02724(.A1(new_n2971_), .A2(new_n2668_), .Z(new_n2991_));
  AOI21_X1   g02725(.A1(new_n2988_), .A2(new_n2983_), .B(new_n2980_), .ZN(new_n2992_));
  NOR3_X1    g02726(.A1(new_n2976_), .A2(new_n2975_), .A3(new_n2981_), .ZN(new_n2993_));
  NOR3_X1    g02727(.A1(new_n2993_), .A2(new_n2992_), .A3(new_n2991_), .ZN(new_n2994_));
  OAI21_X1   g02728(.A1(new_n2994_), .A2(new_n2990_), .B(new_n2869_), .ZN(new_n2995_));
  INV_X1     g02729(.I(new_n2869_), .ZN(new_n2996_));
  OAI21_X1   g02730(.A1(new_n2993_), .A2(new_n2992_), .B(new_n2991_), .ZN(new_n2997_));
  NAND3_X1   g02731(.A1(new_n2982_), .A2(new_n2989_), .A3(new_n2973_), .ZN(new_n2998_));
  NAND3_X1   g02732(.A1(new_n2997_), .A2(new_n2998_), .A3(new_n2996_), .ZN(new_n2999_));
  NAND2_X1   g02733(.A1(new_n2995_), .A2(new_n2999_), .ZN(new_n3000_));
  XOR2_X1    g02734(.A1(new_n2663_), .A2(new_n2987_), .Z(new_n3001_));
  INV_X1     g02735(.I(new_n2800_), .ZN(new_n3002_));
  XOR2_X1    g02736(.A1(new_n3001_), .A2(new_n3002_), .Z(new_n3003_));
  AND3_X2    g02737(.A1(new_n3000_), .A2(new_n3003_), .A3(new_n2802_), .Z(new_n3004_));
  AOI21_X1   g02738(.A1(new_n2997_), .A2(new_n2998_), .B(new_n2996_), .ZN(new_n3005_));
  NOR3_X1    g02739(.A1(new_n2994_), .A2(new_n2990_), .A3(new_n2869_), .ZN(new_n3006_));
  NOR2_X1    g02740(.A1(new_n2796_), .A2(new_n2800_), .ZN(new_n3007_));
  NOR2_X1    g02741(.A1(new_n3004_), .A2(new_n3007_), .ZN(new_n3008_));
  NOR2_X1    g02742(.A1(new_n3008_), .A2(new_n2821_), .ZN(new_n3009_));
  NOR3_X1    g02743(.A1(new_n3004_), .A2(new_n2812_), .A3(new_n3007_), .ZN(new_n3010_));
  NOR2_X1    g02744(.A1(new_n3009_), .A2(new_n3010_), .ZN(new_n3011_));
  OAI22_X1   g02745(.A1(new_n2281_), .A2(new_n341_), .B1(new_n404_), .B2(new_n2439_), .ZN(new_n3012_));
  OAI21_X1   g02746(.A1(new_n2102_), .A2(new_n366_), .B(new_n3012_), .ZN(new_n3013_));
  AOI21_X1   g02747(.A1(new_n3013_), .A2(new_n334_), .B(new_n341_), .ZN(new_n3014_));
  XNOR2_X1   g02748(.A1(new_n2443_), .A2(new_n3014_), .ZN(new_n3015_));
  XOR2_X1    g02749(.A1(new_n3011_), .A2(new_n3015_), .Z(new_n3016_));
  INV_X1     g02750(.I(new_n2841_), .ZN(new_n3017_));
  INV_X1     g02751(.I(\b[29] ), .ZN(new_n3018_));
  NOR2_X1    g02752(.A1(new_n3018_), .A2(\b[27] ), .ZN(new_n3019_));
  NOR2_X1    g02753(.A1(new_n2643_), .A2(\b[29] ), .ZN(new_n3020_));
  OAI21_X1   g02754(.A1(new_n3019_), .A2(new_n3020_), .B(new_n3017_), .ZN(new_n3021_));
  XOR2_X1    g02755(.A1(new_n2840_), .A2(new_n3021_), .Z(new_n3022_));
  NAND2_X1   g02756(.A1(new_n286_), .A2(\b[28] ), .ZN(new_n3023_));
  AOI22_X1   g02757(.A1(new_n304_), .A2(\b[27] ), .B1(new_n262_), .B2(\b[29] ), .ZN(new_n3024_));
  AOI21_X1   g02758(.A1(new_n3023_), .A2(new_n3024_), .B(new_n426_), .ZN(new_n3025_));
  NAND2_X1   g02759(.A1(new_n3022_), .A2(new_n3025_), .ZN(new_n3026_));
  XOR2_X1    g02760(.A1(new_n3026_), .A2(\a[2] ), .Z(new_n3027_));
  INV_X1     g02761(.I(new_n3027_), .ZN(new_n3028_));
  NAND2_X1   g02762(.A1(new_n3016_), .A2(new_n3028_), .ZN(new_n3029_));
  NOR2_X1    g02763(.A1(new_n3029_), .A2(new_n2865_), .ZN(new_n3030_));
  INV_X1     g02764(.I(new_n3030_), .ZN(new_n3031_));
  NAND2_X1   g02765(.A1(new_n3029_), .A2(new_n2865_), .ZN(new_n3032_));
  AOI21_X1   g02766(.A1(new_n3031_), .A2(new_n3032_), .B(new_n2859_), .ZN(new_n3033_));
  INV_X1     g02767(.I(new_n3033_), .ZN(new_n3034_));
  NAND3_X1   g02768(.A1(new_n3031_), .A2(new_n2859_), .A3(new_n3032_), .ZN(new_n3035_));
  AOI21_X1   g02769(.A1(new_n3034_), .A2(new_n3035_), .B(new_n2856_), .ZN(new_n3036_));
  XOR2_X1    g02770(.A1(new_n3036_), .A2(new_n2852_), .Z(new_n3037_));
  XNOR2_X1   g02771(.A1(new_n3037_), .A2(new_n2659_), .ZN(\f[29] ));
  NAND2_X1   g02772(.A1(new_n2988_), .A2(new_n2983_), .ZN(new_n3039_));
  NAND2_X1   g02773(.A1(new_n3039_), .A2(new_n2973_), .ZN(new_n3040_));
  NAND3_X1   g02774(.A1(new_n2988_), .A2(new_n2991_), .A3(new_n2983_), .ZN(new_n3041_));
  NAND2_X1   g02775(.A1(new_n3040_), .A2(new_n3041_), .ZN(new_n3042_));
  NAND2_X1   g02776(.A1(new_n3042_), .A2(new_n2869_), .ZN(new_n3043_));
  NAND3_X1   g02777(.A1(new_n3040_), .A2(new_n2996_), .A3(new_n3041_), .ZN(new_n3044_));
  AOI21_X1   g02778(.A1(new_n3043_), .A2(new_n3044_), .B(new_n2980_), .ZN(new_n3045_));
  AOI21_X1   g02779(.A1(new_n3000_), .A2(new_n3001_), .B(new_n3002_), .ZN(new_n3046_));
  NAND3_X1   g02780(.A1(new_n2995_), .A2(new_n2999_), .A3(new_n2796_), .ZN(new_n3047_));
  NAND2_X1   g02781(.A1(new_n2821_), .A2(new_n3047_), .ZN(new_n3048_));
  NOR2_X1    g02782(.A1(new_n2991_), .A2(new_n2996_), .ZN(new_n3049_));
  INV_X1     g02783(.I(new_n3049_), .ZN(new_n3050_));
  NAND2_X1   g02784(.A1(new_n2973_), .A2(new_n2996_), .ZN(new_n3051_));
  NAND2_X1   g02785(.A1(new_n2991_), .A2(new_n2869_), .ZN(new_n3052_));
  AOI21_X1   g02786(.A1(new_n3051_), .A2(new_n3052_), .B(new_n2983_), .ZN(new_n3053_));
  OAI22_X1   g02787(.A1(new_n3053_), .A2(new_n2795_), .B1(new_n2660_), .B2(new_n2662_), .ZN(new_n3054_));
  AOI21_X1   g02788(.A1(new_n2966_), .A2(new_n2968_), .B(new_n2873_), .ZN(new_n3055_));
  OAI21_X1   g02789(.A1(new_n3055_), .A2(new_n2791_), .B(new_n2668_), .ZN(new_n3056_));
  AOI21_X1   g02790(.A1(new_n2942_), .A2(new_n2944_), .B(new_n2949_), .ZN(new_n3057_));
  NOR3_X1    g02791(.A1(new_n2952_), .A2(new_n2951_), .A3(new_n2948_), .ZN(new_n3058_));
  OAI21_X1   g02792(.A1(new_n3058_), .A2(new_n3057_), .B(new_n2764_), .ZN(new_n3059_));
  NAND2_X1   g02793(.A1(new_n3059_), .A2(new_n2761_), .ZN(new_n3060_));
  INV_X1     g02794(.I(new_n2748_), .ZN(new_n3061_));
  AOI21_X1   g02795(.A1(new_n2749_), .A2(new_n2756_), .B(new_n3061_), .ZN(new_n3062_));
  NAND3_X1   g02796(.A1(new_n2953_), .A2(new_n2950_), .A3(new_n3062_), .ZN(new_n3063_));
  NAND3_X1   g02797(.A1(new_n3060_), .A2(new_n2770_), .A3(new_n3063_), .ZN(new_n3064_));
  AOI21_X1   g02798(.A1(new_n2922_), .A2(new_n2924_), .B(new_n2932_), .ZN(new_n3065_));
  INV_X1     g02799(.I(new_n3065_), .ZN(new_n3066_));
  AOI21_X1   g02800(.A1(new_n2938_), .A2(new_n2739_), .B(new_n2744_), .ZN(new_n3067_));
  NAND3_X1   g02801(.A1(new_n2936_), .A2(new_n2937_), .A3(new_n2738_), .ZN(new_n3068_));
  NAND2_X1   g02802(.A1(new_n2671_), .A2(new_n3068_), .ZN(new_n3069_));
  NOR2_X1    g02803(.A1(new_n3069_), .A2(new_n3067_), .ZN(new_n3070_));
  NAND3_X1   g02804(.A1(new_n2893_), .A2(new_n2891_), .A3(new_n2892_), .ZN(new_n3071_));
  OAI21_X1   g02805(.A1(new_n2906_), .A2(new_n2722_), .B(new_n2890_), .ZN(new_n3072_));
  AOI21_X1   g02806(.A1(new_n3071_), .A2(new_n3072_), .B(new_n2901_), .ZN(new_n3073_));
  NAND3_X1   g02807(.A1(new_n3071_), .A2(new_n3072_), .A3(new_n2901_), .ZN(new_n3074_));
  INV_X1     g02808(.I(new_n3074_), .ZN(new_n3075_));
  OAI21_X1   g02809(.A1(new_n3075_), .A2(new_n3073_), .B(new_n2913_), .ZN(new_n3076_));
  AOI21_X1   g02810(.A1(new_n2914_), .A2(new_n2915_), .B(new_n2913_), .ZN(new_n3077_));
  NOR3_X1    g02811(.A1(new_n2908_), .A2(new_n2911_), .A3(new_n2879_), .ZN(new_n3078_));
  OAI21_X1   g02812(.A1(new_n3078_), .A2(new_n3077_), .B(new_n2724_), .ZN(new_n3079_));
  NAND2_X1   g02813(.A1(new_n3079_), .A2(new_n2729_), .ZN(new_n3080_));
  NOR3_X1    g02814(.A1(new_n3078_), .A2(new_n3077_), .A3(new_n2724_), .ZN(new_n3081_));
  NOR2_X1    g02815(.A1(new_n2682_), .A2(new_n3081_), .ZN(new_n3082_));
  NAND2_X1   g02816(.A1(new_n3082_), .A2(new_n3080_), .ZN(new_n3083_));
  XOR2_X1    g02817(.A1(\a[29] ), .A2(\a[30] ), .Z(new_n3084_));
  NAND2_X1   g02818(.A1(new_n3084_), .A2(\b[0] ), .ZN(new_n3085_));
  AOI22_X1   g02819(.A1(new_n2694_), .A2(\b[2] ), .B1(\b[3] ), .B2(new_n2699_), .ZN(new_n3086_));
  OAI21_X1   g02820(.A1(new_n269_), .A2(new_n2884_), .B(new_n3086_), .ZN(new_n3087_));
  NOR2_X1    g02821(.A1(new_n403_), .A2(new_n2705_), .ZN(new_n3088_));
  AOI21_X1   g02822(.A1(new_n3087_), .A2(new_n3088_), .B(new_n2702_), .ZN(new_n3089_));
  INV_X1     g02823(.I(new_n3089_), .ZN(new_n3090_));
  NAND3_X1   g02824(.A1(new_n3087_), .A2(new_n3088_), .A3(new_n2702_), .ZN(new_n3091_));
  NAND2_X1   g02825(.A1(new_n3090_), .A2(new_n3091_), .ZN(new_n3092_));
  NOR3_X1    g02826(.A1(new_n2710_), .A2(new_n2708_), .A3(new_n2714_), .ZN(new_n3093_));
  NAND2_X1   g02827(.A1(new_n2889_), .A2(new_n3093_), .ZN(new_n3094_));
  OAI22_X1   g02828(.A1(new_n2171_), .A2(new_n419_), .B1(new_n420_), .B2(new_n2166_), .ZN(new_n3095_));
  OAI21_X1   g02829(.A1(new_n325_), .A2(new_n2322_), .B(new_n3095_), .ZN(new_n3096_));
  AOI21_X1   g02830(.A1(new_n3096_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n3097_));
  INV_X1     g02831(.I(new_n3097_), .ZN(new_n3098_));
  NOR2_X1    g02832(.A1(new_n556_), .A2(new_n3098_), .ZN(new_n3099_));
  NOR2_X1    g02833(.A1(new_n425_), .A2(new_n3097_), .ZN(new_n3100_));
  OAI21_X1   g02834(.A1(new_n3099_), .A2(new_n3100_), .B(new_n3094_), .ZN(new_n3101_));
  INV_X1     g02835(.I(new_n2886_), .ZN(new_n3102_));
  NAND2_X1   g02836(.A1(new_n3102_), .A2(new_n2887_), .ZN(new_n3103_));
  NOR2_X1    g02837(.A1(new_n3103_), .A2(new_n2880_), .ZN(new_n3104_));
  NAND2_X1   g02838(.A1(new_n425_), .A2(new_n3097_), .ZN(new_n3105_));
  NAND2_X1   g02839(.A1(new_n556_), .A2(new_n3098_), .ZN(new_n3106_));
  NAND3_X1   g02840(.A1(new_n3104_), .A2(new_n3105_), .A3(new_n3106_), .ZN(new_n3107_));
  AOI21_X1   g02841(.A1(new_n3101_), .A2(new_n3107_), .B(new_n3092_), .ZN(new_n3108_));
  INV_X1     g02842(.I(new_n3091_), .ZN(new_n3109_));
  NOR2_X1    g02843(.A1(new_n3109_), .A2(new_n3089_), .ZN(new_n3110_));
  AOI21_X1   g02844(.A1(new_n3105_), .A2(new_n3106_), .B(new_n3104_), .ZN(new_n3111_));
  NOR3_X1    g02845(.A1(new_n3094_), .A2(new_n3099_), .A3(new_n3100_), .ZN(new_n3112_));
  NOR3_X1    g02846(.A1(new_n3111_), .A2(new_n3110_), .A3(new_n3112_), .ZN(new_n3113_));
  OAI21_X1   g02847(.A1(new_n3113_), .A2(new_n3108_), .B(new_n3085_), .ZN(new_n3114_));
  INV_X1     g02848(.I(new_n3085_), .ZN(new_n3115_));
  OAI21_X1   g02849(.A1(new_n3111_), .A2(new_n3112_), .B(new_n3110_), .ZN(new_n3116_));
  NAND3_X1   g02850(.A1(new_n3101_), .A2(new_n3107_), .A3(new_n3092_), .ZN(new_n3117_));
  NAND3_X1   g02851(.A1(new_n3116_), .A2(new_n3117_), .A3(new_n3115_), .ZN(new_n3118_));
  NAND2_X1   g02852(.A1(new_n3114_), .A2(new_n3118_), .ZN(new_n3119_));
  NOR2_X1    g02853(.A1(new_n2890_), .A2(new_n2901_), .ZN(new_n3120_));
  INV_X1     g02854(.I(new_n3120_), .ZN(new_n3121_));
  INV_X1     g02855(.I(new_n2899_), .ZN(new_n3122_));
  NAND2_X1   g02856(.A1(new_n2880_), .A2(new_n3122_), .ZN(new_n3123_));
  NAND2_X1   g02857(.A1(new_n3093_), .A2(new_n2899_), .ZN(new_n3124_));
  AOI21_X1   g02858(.A1(new_n3124_), .A2(new_n3123_), .B(new_n3103_), .ZN(new_n3125_));
  NOR2_X1    g02859(.A1(new_n3093_), .A2(new_n2899_), .ZN(new_n3126_));
  NOR2_X1    g02860(.A1(new_n2880_), .A2(new_n3122_), .ZN(new_n3127_));
  NOR3_X1    g02861(.A1(new_n3126_), .A2(new_n3127_), .A3(new_n2889_), .ZN(new_n3128_));
  OAI21_X1   g02862(.A1(new_n3125_), .A2(new_n3128_), .B(new_n2168_), .ZN(new_n3129_));
  OAI21_X1   g02863(.A1(new_n3126_), .A2(new_n3127_), .B(new_n2889_), .ZN(new_n3130_));
  NAND3_X1   g02864(.A1(new_n3124_), .A2(new_n3123_), .A3(new_n3103_), .ZN(new_n3131_));
  NAND3_X1   g02865(.A1(new_n3130_), .A2(new_n3131_), .A3(\a[26] ), .ZN(new_n3132_));
  NAND2_X1   g02866(.A1(new_n3129_), .A2(new_n3132_), .ZN(new_n3133_));
  AOI21_X1   g02867(.A1(new_n3133_), .A2(new_n2721_), .B(new_n2691_), .ZN(new_n3134_));
  NAND3_X1   g02868(.A1(new_n3129_), .A2(new_n3132_), .A3(new_n2716_), .ZN(new_n3135_));
  NAND2_X1   g02869(.A1(new_n3135_), .A2(new_n2687_), .ZN(new_n3136_));
  OR2_X2     g02870(.A1(new_n3134_), .A2(new_n3136_), .Z(new_n3137_));
  AOI21_X1   g02871(.A1(new_n3137_), .A2(new_n3121_), .B(new_n3119_), .ZN(new_n3138_));
  AND2_X2    g02872(.A1(new_n3114_), .A2(new_n3118_), .Z(new_n3139_));
  NOR2_X1    g02873(.A1(new_n3134_), .A2(new_n3136_), .ZN(new_n3140_));
  NOR3_X1    g02874(.A1(new_n3139_), .A2(new_n3120_), .A3(new_n3140_), .ZN(new_n3141_));
  NOR2_X1    g02875(.A1(new_n3138_), .A2(new_n3141_), .ZN(new_n3142_));
  OAI22_X1   g02876(.A1(new_n1712_), .A2(new_n515_), .B1(new_n565_), .B2(new_n1707_), .ZN(new_n3143_));
  OAI21_X1   g02877(.A1(new_n472_), .A2(new_n1850_), .B(new_n3143_), .ZN(new_n3144_));
  AOI21_X1   g02878(.A1(new_n3144_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n3145_));
  XOR2_X1    g02879(.A1(new_n759_), .A2(new_n3145_), .Z(new_n3146_));
  NOR2_X1    g02880(.A1(new_n3142_), .A2(new_n3146_), .ZN(new_n3147_));
  NAND2_X1   g02881(.A1(new_n3083_), .A2(new_n3147_), .ZN(new_n3148_));
  AOI21_X1   g02882(.A1(new_n2917_), .A2(new_n2724_), .B(new_n2730_), .ZN(new_n3149_));
  NAND3_X1   g02883(.A1(new_n2912_), .A2(new_n2916_), .A3(new_n2732_), .ZN(new_n3150_));
  NAND3_X1   g02884(.A1(new_n3150_), .A2(new_n2672_), .A3(new_n2681_), .ZN(new_n3151_));
  NOR2_X1    g02885(.A1(new_n3151_), .A2(new_n3149_), .ZN(new_n3152_));
  OAI21_X1   g02886(.A1(new_n3140_), .A2(new_n3120_), .B(new_n3139_), .ZN(new_n3153_));
  NAND3_X1   g02887(.A1(new_n3137_), .A2(new_n3119_), .A3(new_n3121_), .ZN(new_n3154_));
  NAND2_X1   g02888(.A1(new_n3154_), .A2(new_n3153_), .ZN(new_n3155_));
  INV_X1     g02889(.I(new_n3146_), .ZN(new_n3156_));
  NAND2_X1   g02890(.A1(new_n3155_), .A2(new_n3156_), .ZN(new_n3157_));
  NAND2_X1   g02891(.A1(new_n3152_), .A2(new_n3157_), .ZN(new_n3158_));
  NAND2_X1   g02892(.A1(new_n3148_), .A2(new_n3158_), .ZN(new_n3159_));
  NAND2_X1   g02893(.A1(new_n3159_), .A2(new_n3076_), .ZN(new_n3160_));
  INV_X1     g02894(.I(new_n3073_), .ZN(new_n3161_));
  AOI21_X1   g02895(.A1(new_n3161_), .A2(new_n3074_), .B(new_n2879_), .ZN(new_n3162_));
  XOR2_X1    g02896(.A1(new_n3152_), .A2(new_n3157_), .Z(new_n3163_));
  NAND2_X1   g02897(.A1(new_n3163_), .A2(new_n3162_), .ZN(new_n3164_));
  NAND2_X1   g02898(.A1(new_n3164_), .A2(new_n3160_), .ZN(new_n3165_));
  OAI22_X1   g02899(.A1(new_n1347_), .A2(new_n706_), .B1(new_n780_), .B2(new_n1344_), .ZN(new_n3166_));
  OAI21_X1   g02900(.A1(new_n656_), .A2(new_n1457_), .B(new_n3166_), .ZN(new_n3167_));
  AOI21_X1   g02901(.A1(new_n3167_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n3168_));
  XOR2_X1    g02902(.A1(new_n785_), .A2(new_n3168_), .Z(new_n3169_));
  INV_X1     g02903(.I(new_n3169_), .ZN(new_n3170_));
  NAND2_X1   g02904(.A1(new_n3165_), .A2(new_n3170_), .ZN(new_n3171_));
  NOR2_X1    g02905(.A1(new_n3070_), .A2(new_n3171_), .ZN(new_n3172_));
  OAI21_X1   g02906(.A1(new_n2933_), .A2(new_n2929_), .B(new_n2739_), .ZN(new_n3173_));
  NAND2_X1   g02907(.A1(new_n3173_), .A2(new_n2743_), .ZN(new_n3174_));
  NAND3_X1   g02908(.A1(new_n3174_), .A2(new_n2671_), .A3(new_n3068_), .ZN(new_n3175_));
  NOR2_X1    g02909(.A1(new_n3163_), .A2(new_n3162_), .ZN(new_n3176_));
  NOR2_X1    g02910(.A1(new_n3159_), .A2(new_n3076_), .ZN(new_n3177_));
  NOR2_X1    g02911(.A1(new_n3176_), .A2(new_n3177_), .ZN(new_n3178_));
  NOR2_X1    g02912(.A1(new_n3178_), .A2(new_n3169_), .ZN(new_n3179_));
  NOR2_X1    g02913(.A1(new_n3179_), .A2(new_n3175_), .ZN(new_n3180_));
  OAI21_X1   g02914(.A1(new_n3172_), .A2(new_n3180_), .B(new_n3066_), .ZN(new_n3181_));
  NAND2_X1   g02915(.A1(new_n3179_), .A2(new_n3175_), .ZN(new_n3182_));
  NAND2_X1   g02916(.A1(new_n3070_), .A2(new_n3171_), .ZN(new_n3183_));
  NAND3_X1   g02917(.A1(new_n3183_), .A2(new_n3182_), .A3(new_n3065_), .ZN(new_n3184_));
  NAND2_X1   g02918(.A1(new_n3181_), .A2(new_n3184_), .ZN(new_n3185_));
  OAI22_X1   g02919(.A1(new_n1055_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n1061_), .ZN(new_n3186_));
  OAI21_X1   g02920(.A1(new_n861_), .A2(new_n1332_), .B(new_n3186_), .ZN(new_n3187_));
  AOI21_X1   g02921(.A1(new_n3187_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n3188_));
  XOR2_X1    g02922(.A1(new_n1024_), .A2(new_n3188_), .Z(new_n3189_));
  INV_X1     g02923(.I(new_n3189_), .ZN(new_n3190_));
  NAND2_X1   g02924(.A1(new_n3185_), .A2(new_n3190_), .ZN(new_n3191_));
  INV_X1     g02925(.I(new_n3191_), .ZN(new_n3192_));
  NAND2_X1   g02926(.A1(new_n3192_), .A2(new_n3064_), .ZN(new_n3193_));
  AOI21_X1   g02927(.A1(new_n2954_), .A2(new_n2764_), .B(new_n2762_), .ZN(new_n3194_));
  NAND2_X1   g02928(.A1(new_n3063_), .A2(new_n2770_), .ZN(new_n3195_));
  NOR2_X1    g02929(.A1(new_n3194_), .A2(new_n3195_), .ZN(new_n3196_));
  NAND2_X1   g02930(.A1(new_n3196_), .A2(new_n3191_), .ZN(new_n3197_));
  AOI21_X1   g02931(.A1(new_n3193_), .A2(new_n3197_), .B(new_n3057_), .ZN(new_n3198_));
  NOR2_X1    g02932(.A1(new_n3196_), .A2(new_n3191_), .ZN(new_n3199_));
  NOR2_X1    g02933(.A1(new_n3192_), .A2(new_n3064_), .ZN(new_n3200_));
  NOR3_X1    g02934(.A1(new_n3200_), .A2(new_n3199_), .A3(new_n2953_), .ZN(new_n3201_));
  NOR2_X1    g02935(.A1(new_n3201_), .A2(new_n3198_), .ZN(new_n3202_));
  OAI22_X1   g02936(.A1(new_n970_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n820_), .ZN(new_n3203_));
  OAI21_X1   g02937(.A1(new_n1109_), .A2(new_n894_), .B(new_n3203_), .ZN(new_n3204_));
  AOI21_X1   g02938(.A1(new_n3204_), .A2(new_n827_), .B(new_n970_), .ZN(new_n3205_));
  XOR2_X1    g02939(.A1(new_n1299_), .A2(new_n3205_), .Z(new_n3206_));
  NOR2_X1    g02940(.A1(new_n3202_), .A2(new_n3206_), .ZN(new_n3207_));
  NAND2_X1   g02941(.A1(new_n3056_), .A2(new_n3207_), .ZN(new_n3208_));
  INV_X1     g02942(.I(new_n3208_), .ZN(new_n3209_));
  NOR2_X1    g02943(.A1(new_n3056_), .A2(new_n3207_), .ZN(new_n3210_));
  OAI21_X1   g02944(.A1(new_n3209_), .A2(new_n3210_), .B(new_n2968_), .ZN(new_n3211_));
  INV_X1     g02945(.I(new_n2968_), .ZN(new_n3212_));
  INV_X1     g02946(.I(new_n3210_), .ZN(new_n3213_));
  NAND3_X1   g02947(.A1(new_n3213_), .A2(new_n3212_), .A3(new_n3208_), .ZN(new_n3214_));
  NAND2_X1   g02948(.A1(new_n3211_), .A2(new_n3214_), .ZN(new_n3215_));
  OAI22_X1   g02949(.A1(new_n607_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n610_), .ZN(new_n3216_));
  OAI21_X1   g02950(.A1(new_n1518_), .A2(new_n684_), .B(new_n3216_), .ZN(new_n3217_));
  AOI21_X1   g02951(.A1(new_n3217_), .A2(new_n612_), .B(new_n607_), .ZN(new_n3218_));
  XNOR2_X1   g02952(.A1(new_n1638_), .A2(new_n3218_), .ZN(new_n3219_));
  INV_X1     g02953(.I(new_n3219_), .ZN(new_n3220_));
  NAND2_X1   g02954(.A1(new_n3215_), .A2(new_n3220_), .ZN(new_n3221_));
  XOR2_X1    g02955(.A1(new_n3054_), .A2(new_n3221_), .Z(new_n3222_));
  NAND2_X1   g02956(.A1(new_n3222_), .A2(new_n3050_), .ZN(new_n3223_));
  NAND2_X1   g02957(.A1(new_n3052_), .A2(new_n3051_), .ZN(new_n3224_));
  NAND2_X1   g02958(.A1(new_n3224_), .A2(new_n2975_), .ZN(new_n3225_));
  AOI21_X1   g02959(.A1(new_n3225_), .A2(new_n2987_), .B(new_n2663_), .ZN(new_n3226_));
  NOR2_X1    g02960(.A1(new_n3226_), .A2(new_n3221_), .ZN(new_n3227_));
  INV_X1     g02961(.I(new_n3221_), .ZN(new_n3228_));
  NOR2_X1    g02962(.A1(new_n3228_), .A2(new_n3054_), .ZN(new_n3229_));
  NOR2_X1    g02963(.A1(new_n3227_), .A2(new_n3229_), .ZN(new_n3230_));
  NAND2_X1   g02964(.A1(new_n3230_), .A2(new_n3049_), .ZN(new_n3231_));
  OAI22_X1   g02965(.A1(new_n448_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n450_), .ZN(new_n3232_));
  OAI21_X1   g02966(.A1(new_n1803_), .A2(new_n496_), .B(new_n3232_), .ZN(new_n3233_));
  AOI21_X1   g02967(.A1(new_n3233_), .A2(new_n452_), .B(new_n448_), .ZN(new_n3234_));
  XOR2_X1    g02968(.A1(new_n2106_), .A2(new_n3234_), .Z(new_n3235_));
  AOI21_X1   g02969(.A1(new_n3231_), .A2(new_n3223_), .B(new_n3235_), .ZN(new_n3236_));
  OAI21_X1   g02970(.A1(new_n3046_), .A2(new_n3048_), .B(new_n3236_), .ZN(new_n3237_));
  NOR2_X1    g02971(.A1(new_n3048_), .A2(new_n3046_), .ZN(new_n3238_));
  INV_X1     g02972(.I(new_n3236_), .ZN(new_n3239_));
  NAND2_X1   g02973(.A1(new_n3239_), .A2(new_n3238_), .ZN(new_n3240_));
  NAND2_X1   g02974(.A1(new_n3240_), .A2(new_n3237_), .ZN(new_n3241_));
  XOR2_X1    g02975(.A1(new_n3241_), .A2(new_n3045_), .Z(new_n3242_));
  OAI22_X1   g02976(.A1(new_n2439_), .A2(new_n341_), .B1(new_n404_), .B2(new_n2643_), .ZN(new_n3243_));
  OAI21_X1   g02977(.A1(new_n2281_), .A2(new_n366_), .B(new_n3243_), .ZN(new_n3244_));
  AOI21_X1   g02978(.A1(new_n3244_), .A2(new_n334_), .B(new_n341_), .ZN(new_n3245_));
  XNOR2_X1   g02979(.A1(new_n2647_), .A2(new_n3245_), .ZN(new_n3246_));
  XOR2_X1    g02980(.A1(new_n3242_), .A2(new_n3246_), .Z(new_n3247_));
  OAI21_X1   g02981(.A1(new_n3009_), .A2(new_n3010_), .B(new_n2859_), .ZN(new_n3248_));
  NOR3_X1    g02982(.A1(new_n3009_), .A2(new_n2859_), .A3(new_n3010_), .ZN(new_n3249_));
  INV_X1     g02983(.I(new_n3015_), .ZN(new_n3250_));
  NAND3_X1   g02984(.A1(new_n2863_), .A2(new_n2860_), .A3(new_n3250_), .ZN(new_n3251_));
  OAI21_X1   g02985(.A1(new_n3251_), .A2(new_n3249_), .B(new_n3248_), .ZN(new_n3252_));
  NOR2_X1    g02986(.A1(\b[28] ), .A2(\b[29] ), .ZN(new_n3253_));
  AOI21_X1   g02987(.A1(new_n2840_), .A2(new_n3253_), .B(new_n2643_), .ZN(new_n3254_));
  NOR2_X1    g02988(.A1(new_n2842_), .A2(new_n3018_), .ZN(new_n3255_));
  INV_X1     g02989(.I(new_n3255_), .ZN(new_n3256_));
  NOR2_X1    g02990(.A1(new_n2840_), .A2(new_n3256_), .ZN(new_n3257_));
  NOR2_X1    g02991(.A1(new_n3254_), .A2(new_n3257_), .ZN(new_n3258_));
  XNOR2_X1   g02992(.A1(\b[29] ), .A2(\b[30] ), .ZN(new_n3259_));
  INV_X1     g02993(.I(\b[30] ), .ZN(new_n3260_));
  NOR2_X1    g02994(.A1(new_n3018_), .A2(new_n3260_), .ZN(new_n3261_));
  NOR2_X1    g02995(.A1(\b[29] ), .A2(\b[30] ), .ZN(new_n3262_));
  OAI21_X1   g02996(.A1(new_n3261_), .A2(new_n3262_), .B(new_n3258_), .ZN(new_n3263_));
  OAI21_X1   g02997(.A1(new_n3258_), .A2(new_n3259_), .B(new_n3263_), .ZN(new_n3264_));
  OAI22_X1   g02998(.A1(new_n330_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n263_), .ZN(new_n3265_));
  OAI21_X1   g02999(.A1(new_n2842_), .A2(new_n289_), .B(new_n3265_), .ZN(new_n3266_));
  AOI21_X1   g03000(.A1(new_n3266_), .A2(new_n260_), .B(new_n426_), .ZN(new_n3267_));
  XNOR2_X1   g03001(.A1(new_n3264_), .A2(new_n3267_), .ZN(new_n3268_));
  INV_X1     g03002(.I(new_n3268_), .ZN(new_n3269_));
  NAND2_X1   g03003(.A1(new_n3252_), .A2(new_n3269_), .ZN(new_n3270_));
  NOR2_X1    g03004(.A1(new_n3252_), .A2(new_n3269_), .ZN(new_n3271_));
  INV_X1     g03005(.I(new_n3271_), .ZN(new_n3272_));
  AOI21_X1   g03006(.A1(new_n3270_), .A2(new_n3272_), .B(new_n3247_), .ZN(new_n3273_));
  INV_X1     g03007(.I(new_n3247_), .ZN(new_n3274_));
  INV_X1     g03008(.I(new_n3252_), .ZN(new_n3275_));
  NAND2_X1   g03009(.A1(new_n3275_), .A2(new_n3269_), .ZN(new_n3276_));
  NAND2_X1   g03010(.A1(new_n3252_), .A2(new_n3268_), .ZN(new_n3277_));
  AOI21_X1   g03011(.A1(new_n3277_), .A2(new_n3276_), .B(new_n3274_), .ZN(new_n3278_));
  NOR2_X1    g03012(.A1(new_n3278_), .A2(new_n3273_), .ZN(new_n3279_));
  INV_X1     g03013(.I(new_n3035_), .ZN(new_n3280_));
  OAI21_X1   g03014(.A1(new_n3280_), .A2(new_n3033_), .B(new_n2834_), .ZN(new_n3281_));
  NAND2_X1   g03015(.A1(new_n3281_), .A2(new_n2850_), .ZN(new_n3282_));
  NAND3_X1   g03016(.A1(new_n3034_), .A2(new_n3035_), .A3(new_n2833_), .ZN(new_n3283_));
  NAND3_X1   g03017(.A1(new_n2659_), .A2(new_n3282_), .A3(new_n3283_), .ZN(new_n3284_));
  INV_X1     g03018(.I(new_n3284_), .ZN(new_n3285_));
  OR2_X2     g03019(.A1(new_n3029_), .A2(new_n2859_), .Z(new_n3286_));
  NAND2_X1   g03020(.A1(new_n3029_), .A2(new_n2859_), .ZN(new_n3287_));
  NAND2_X1   g03021(.A1(new_n3286_), .A2(new_n3287_), .ZN(new_n3288_));
  AND2_X2    g03022(.A1(new_n3288_), .A2(new_n2865_), .Z(new_n3289_));
  NOR2_X1    g03023(.A1(new_n3285_), .A2(new_n3289_), .ZN(new_n3290_));
  INV_X1     g03024(.I(new_n3289_), .ZN(new_n3291_));
  NAND2_X1   g03025(.A1(new_n3291_), .A2(new_n3279_), .ZN(new_n3292_));
  OAI22_X1   g03026(.A1(new_n3290_), .A2(new_n3279_), .B1(new_n3285_), .B2(new_n3292_), .ZN(\f[30] ));
  INV_X1     g03027(.I(new_n3242_), .ZN(new_n3294_));
  NOR2_X1    g03028(.A1(new_n3294_), .A2(new_n3246_), .ZN(new_n3295_));
  NOR2_X1    g03029(.A1(new_n3230_), .A2(new_n3049_), .ZN(new_n3296_));
  NOR2_X1    g03030(.A1(new_n3222_), .A2(new_n3050_), .ZN(new_n3297_));
  OAI21_X1   g03031(.A1(new_n3297_), .A2(new_n3296_), .B(new_n3045_), .ZN(new_n3298_));
  NOR3_X1    g03032(.A1(new_n3297_), .A2(new_n3296_), .A3(new_n3045_), .ZN(new_n3299_));
  OAI21_X1   g03033(.A1(new_n3006_), .A2(new_n3005_), .B(new_n3001_), .ZN(new_n3300_));
  NAND2_X1   g03034(.A1(new_n3300_), .A2(new_n2800_), .ZN(new_n3301_));
  INV_X1     g03035(.I(new_n3235_), .ZN(new_n3302_));
  NAND4_X1   g03036(.A1(new_n3301_), .A2(new_n2821_), .A3(new_n3047_), .A4(new_n3302_), .ZN(new_n3303_));
  OAI21_X1   g03037(.A1(new_n3303_), .A2(new_n3299_), .B(new_n3298_), .ZN(new_n3304_));
  AND2_X2    g03038(.A1(new_n3211_), .A2(new_n3214_), .Z(new_n3305_));
  NOR2_X1    g03039(.A1(new_n3305_), .A2(new_n3050_), .ZN(new_n3306_));
  AOI21_X1   g03040(.A1(new_n3305_), .A2(new_n3050_), .B(new_n3219_), .ZN(new_n3307_));
  AOI21_X1   g03041(.A1(new_n3307_), .A2(new_n3226_), .B(new_n3306_), .ZN(new_n3308_));
  OAI21_X1   g03042(.A1(new_n3200_), .A2(new_n3199_), .B(new_n2953_), .ZN(new_n3309_));
  NAND3_X1   g03043(.A1(new_n3193_), .A2(new_n3197_), .A3(new_n3057_), .ZN(new_n3310_));
  NAND2_X1   g03044(.A1(new_n3309_), .A2(new_n3310_), .ZN(new_n3311_));
  NAND2_X1   g03045(.A1(new_n3311_), .A2(new_n3212_), .ZN(new_n3312_));
  NAND2_X1   g03046(.A1(new_n2966_), .A2(new_n2968_), .ZN(new_n3313_));
  NAND2_X1   g03047(.A1(new_n3313_), .A2(new_n2872_), .ZN(new_n3314_));
  NAND2_X1   g03048(.A1(new_n3314_), .A2(new_n2782_), .ZN(new_n3315_));
  AOI21_X1   g03049(.A1(new_n3202_), .A2(new_n2968_), .B(new_n3206_), .ZN(new_n3316_));
  NAND3_X1   g03050(.A1(new_n3315_), .A2(new_n3316_), .A3(new_n2668_), .ZN(new_n3317_));
  AOI21_X1   g03051(.A1(new_n3183_), .A2(new_n3182_), .B(new_n3065_), .ZN(new_n3318_));
  NOR3_X1    g03052(.A1(new_n3172_), .A2(new_n3180_), .A3(new_n3066_), .ZN(new_n3319_));
  NOR2_X1    g03053(.A1(new_n3318_), .A2(new_n3319_), .ZN(new_n3320_));
  NOR2_X1    g03054(.A1(new_n3320_), .A2(new_n2953_), .ZN(new_n3321_));
  AOI21_X1   g03055(.A1(new_n3320_), .A2(new_n2953_), .B(new_n3189_), .ZN(new_n3322_));
  AOI21_X1   g03056(.A1(new_n3196_), .A2(new_n3322_), .B(new_n3321_), .ZN(new_n3323_));
  NAND2_X1   g03057(.A1(new_n3155_), .A2(new_n3162_), .ZN(new_n3324_));
  NAND3_X1   g03058(.A1(new_n3154_), .A2(new_n3153_), .A3(new_n3076_), .ZN(new_n3325_));
  NAND4_X1   g03059(.A1(new_n3082_), .A2(new_n3325_), .A3(new_n3080_), .A4(new_n3156_), .ZN(new_n3326_));
  NAND2_X1   g03060(.A1(new_n3326_), .A2(new_n3324_), .ZN(new_n3327_));
  NAND2_X1   g03061(.A1(new_n3094_), .A2(new_n3092_), .ZN(new_n3328_));
  NAND2_X1   g03062(.A1(new_n3104_), .A2(new_n3110_), .ZN(new_n3329_));
  NAND2_X1   g03063(.A1(new_n3329_), .A2(new_n3328_), .ZN(new_n3330_));
  NAND2_X1   g03064(.A1(new_n3330_), .A2(new_n3085_), .ZN(new_n3331_));
  NAND3_X1   g03065(.A1(new_n3329_), .A2(new_n3328_), .A3(new_n3115_), .ZN(new_n3332_));
  AOI22_X1   g03066(.A1(new_n3331_), .A2(new_n3332_), .B1(new_n3105_), .B2(new_n3106_), .ZN(new_n3333_));
  AOI21_X1   g03067(.A1(new_n3119_), .A2(new_n3333_), .B(new_n3120_), .ZN(new_n3334_));
  NOR2_X1    g03068(.A1(new_n3334_), .A2(new_n3137_), .ZN(new_n3335_));
  NAND2_X1   g03069(.A1(new_n3103_), .A2(new_n3092_), .ZN(new_n3336_));
  NOR2_X1    g03070(.A1(new_n2880_), .A2(new_n3085_), .ZN(new_n3337_));
  OAI21_X1   g03071(.A1(new_n3103_), .A2(new_n3092_), .B(new_n3337_), .ZN(new_n3338_));
  NAND2_X1   g03072(.A1(new_n3338_), .A2(new_n3336_), .ZN(new_n3339_));
  OAI22_X1   g03073(.A1(new_n325_), .A2(new_n2700_), .B1(new_n2705_), .B2(new_n298_), .ZN(new_n3340_));
  OAI21_X1   g03074(.A1(new_n280_), .A2(new_n2884_), .B(new_n3340_), .ZN(new_n3341_));
  AOI21_X1   g03075(.A1(new_n3341_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n3342_));
  XOR2_X1    g03076(.A1(new_n3342_), .A2(new_n807_), .Z(new_n3343_));
  XNOR2_X1   g03077(.A1(\a[30] ), .A2(\a[32] ), .ZN(new_n3344_));
  XNOR2_X1   g03078(.A1(\a[29] ), .A2(\a[31] ), .ZN(new_n3345_));
  NOR2_X1    g03079(.A1(new_n3345_), .A2(new_n3344_), .ZN(new_n3346_));
  INV_X1     g03080(.I(\a[30] ), .ZN(new_n3347_));
  NAND3_X1   g03081(.A1(new_n2702_), .A2(new_n3347_), .A3(\a[31] ), .ZN(new_n3348_));
  INV_X1     g03082(.I(\a[31] ), .ZN(new_n3349_));
  NAND3_X1   g03083(.A1(new_n3349_), .A2(\a[29] ), .A3(\a[30] ), .ZN(new_n3350_));
  NAND2_X1   g03084(.A1(new_n3348_), .A2(new_n3350_), .ZN(new_n3351_));
  INV_X1     g03085(.I(new_n3351_), .ZN(new_n3352_));
  NOR2_X1    g03086(.A1(new_n3352_), .A2(new_n269_), .ZN(new_n3353_));
  INV_X1     g03087(.I(\a[32] ), .ZN(new_n3354_));
  XOR2_X1    g03088(.A1(\a[30] ), .A2(\a[32] ), .Z(new_n3355_));
  XOR2_X1    g03089(.A1(\a[29] ), .A2(\a[31] ), .Z(new_n3356_));
  NAND2_X1   g03090(.A1(new_n3356_), .A2(new_n3355_), .ZN(new_n3357_));
  OAI21_X1   g03091(.A1(new_n3357_), .A2(new_n258_), .B(new_n3354_), .ZN(new_n3358_));
  OAI21_X1   g03092(.A1(new_n3358_), .A2(new_n3353_), .B(new_n3346_), .ZN(new_n3359_));
  NOR2_X1    g03093(.A1(new_n3359_), .A2(new_n271_), .ZN(new_n3360_));
  INV_X1     g03094(.I(new_n3360_), .ZN(new_n3361_));
  NAND2_X1   g03095(.A1(new_n3359_), .A2(new_n271_), .ZN(new_n3362_));
  NAND2_X1   g03096(.A1(new_n3085_), .A2(\a[32] ), .ZN(new_n3363_));
  NAND3_X1   g03097(.A1(new_n3361_), .A2(new_n3362_), .A3(new_n3363_), .ZN(new_n3364_));
  INV_X1     g03098(.I(new_n3364_), .ZN(new_n3365_));
  INV_X1     g03099(.I(new_n3362_), .ZN(new_n3366_));
  NOR2_X1    g03100(.A1(new_n3366_), .A2(new_n3360_), .ZN(new_n3367_));
  NOR2_X1    g03101(.A1(new_n3367_), .A2(new_n3363_), .ZN(new_n3368_));
  NOR2_X1    g03102(.A1(new_n3368_), .A2(new_n3365_), .ZN(new_n3369_));
  NOR2_X1    g03103(.A1(new_n3369_), .A2(new_n3343_), .ZN(new_n3370_));
  XOR2_X1    g03104(.A1(new_n3342_), .A2(new_n329_), .Z(new_n3371_));
  NAND2_X1   g03105(.A1(new_n3361_), .A2(new_n3362_), .ZN(new_n3372_));
  INV_X1     g03106(.I(new_n3363_), .ZN(new_n3373_));
  NAND2_X1   g03107(.A1(new_n3372_), .A2(new_n3373_), .ZN(new_n3374_));
  NAND2_X1   g03108(.A1(new_n3374_), .A2(new_n3364_), .ZN(new_n3375_));
  NOR2_X1    g03109(.A1(new_n3375_), .A2(new_n3371_), .ZN(new_n3376_));
  OAI21_X1   g03110(.A1(new_n3370_), .A2(new_n3376_), .B(new_n3339_), .ZN(new_n3377_));
  NOR2_X1    g03111(.A1(new_n2889_), .A2(new_n3110_), .ZN(new_n3378_));
  NAND4_X1   g03112(.A1(new_n2713_), .A2(new_n2709_), .A3(new_n2711_), .A4(new_n3115_), .ZN(new_n3379_));
  AOI21_X1   g03113(.A1(new_n2889_), .A2(new_n3110_), .B(new_n3379_), .ZN(new_n3380_));
  NOR2_X1    g03114(.A1(new_n3380_), .A2(new_n3378_), .ZN(new_n3381_));
  NOR2_X1    g03115(.A1(new_n3369_), .A2(new_n3371_), .ZN(new_n3382_));
  NOR2_X1    g03116(.A1(new_n3375_), .A2(new_n3343_), .ZN(new_n3383_));
  OAI21_X1   g03117(.A1(new_n3382_), .A2(new_n3383_), .B(new_n3381_), .ZN(new_n3384_));
  NAND2_X1   g03118(.A1(new_n3377_), .A2(new_n3384_), .ZN(new_n3385_));
  AOI22_X1   g03119(.A1(\b[7] ), .A2(new_n2896_), .B1(new_n2161_), .B2(\b[6] ), .ZN(new_n3386_));
  AOI21_X1   g03120(.A1(\b[5] ), .A2(new_n2895_), .B(new_n3386_), .ZN(new_n3387_));
  OAI21_X1   g03121(.A1(new_n3387_), .A2(\a[26] ), .B(new_n2161_), .ZN(new_n3388_));
  XNOR2_X1   g03122(.A1(new_n471_), .A2(new_n3388_), .ZN(new_n3389_));
  INV_X1     g03123(.I(new_n3389_), .ZN(new_n3390_));
  NAND2_X1   g03124(.A1(new_n3385_), .A2(new_n3390_), .ZN(new_n3391_));
  NOR2_X1    g03125(.A1(new_n3370_), .A2(new_n3376_), .ZN(new_n3392_));
  NOR2_X1    g03126(.A1(new_n3392_), .A2(new_n3381_), .ZN(new_n3393_));
  INV_X1     g03127(.I(new_n3384_), .ZN(new_n3394_));
  NOR2_X1    g03128(.A1(new_n3394_), .A2(new_n3393_), .ZN(new_n3395_));
  NAND2_X1   g03129(.A1(new_n3395_), .A2(new_n3389_), .ZN(new_n3396_));
  NAND2_X1   g03130(.A1(new_n3396_), .A2(new_n3391_), .ZN(new_n3397_));
  NAND2_X1   g03131(.A1(new_n3335_), .A2(new_n3397_), .ZN(new_n3398_));
  NAND3_X1   g03132(.A1(new_n3377_), .A2(new_n3384_), .A3(new_n3390_), .ZN(new_n3399_));
  OAI21_X1   g03133(.A1(new_n3394_), .A2(new_n3393_), .B(new_n3389_), .ZN(new_n3400_));
  NAND2_X1   g03134(.A1(new_n3400_), .A2(new_n3399_), .ZN(new_n3401_));
  OAI21_X1   g03135(.A1(new_n3334_), .A2(new_n3137_), .B(new_n3401_), .ZN(new_n3402_));
  NAND2_X1   g03136(.A1(new_n3398_), .A2(new_n3402_), .ZN(new_n3403_));
  OAI22_X1   g03137(.A1(new_n1712_), .A2(new_n565_), .B1(new_n656_), .B2(new_n1707_), .ZN(new_n3404_));
  OAI21_X1   g03138(.A1(new_n515_), .A2(new_n1850_), .B(new_n3404_), .ZN(new_n3405_));
  AOI21_X1   g03139(.A1(new_n3405_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n3406_));
  XNOR2_X1   g03140(.A1(new_n660_), .A2(new_n3406_), .ZN(new_n3407_));
  INV_X1     g03141(.I(new_n3407_), .ZN(new_n3408_));
  NAND2_X1   g03142(.A1(new_n3403_), .A2(new_n3408_), .ZN(new_n3409_));
  AND2_X2    g03143(.A1(new_n3396_), .A2(new_n3391_), .Z(new_n3410_));
  NOR3_X1    g03144(.A1(new_n3410_), .A2(new_n3137_), .A3(new_n3334_), .ZN(new_n3411_));
  INV_X1     g03145(.I(new_n3402_), .ZN(new_n3412_));
  NOR2_X1    g03146(.A1(new_n3411_), .A2(new_n3412_), .ZN(new_n3413_));
  NAND2_X1   g03147(.A1(new_n3413_), .A2(new_n3407_), .ZN(new_n3414_));
  NAND2_X1   g03148(.A1(new_n3414_), .A2(new_n3409_), .ZN(new_n3415_));
  NAND2_X1   g03149(.A1(new_n3415_), .A2(new_n3327_), .ZN(new_n3416_));
  NOR2_X1    g03150(.A1(new_n3142_), .A2(new_n3076_), .ZN(new_n3417_));
  NOR3_X1    g03151(.A1(new_n3138_), .A2(new_n3141_), .A3(new_n3162_), .ZN(new_n3418_));
  NOR4_X1    g03152(.A1(new_n3151_), .A2(new_n3418_), .A3(new_n3149_), .A4(new_n3146_), .ZN(new_n3419_));
  NOR2_X1    g03153(.A1(new_n3419_), .A2(new_n3417_), .ZN(new_n3420_));
  NOR2_X1    g03154(.A1(new_n3403_), .A2(new_n3407_), .ZN(new_n3421_));
  AOI21_X1   g03155(.A1(new_n3398_), .A2(new_n3402_), .B(new_n3408_), .ZN(new_n3422_));
  OAI21_X1   g03156(.A1(new_n3421_), .A2(new_n3422_), .B(new_n3420_), .ZN(new_n3423_));
  NAND2_X1   g03157(.A1(new_n3423_), .A2(new_n3416_), .ZN(new_n3424_));
  OAI22_X1   g03158(.A1(new_n1347_), .A2(new_n780_), .B1(new_n861_), .B2(new_n1344_), .ZN(new_n3425_));
  OAI21_X1   g03159(.A1(new_n706_), .A2(new_n1457_), .B(new_n3425_), .ZN(new_n3426_));
  AOI21_X1   g03160(.A1(new_n3426_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n3427_));
  XNOR2_X1   g03161(.A1(new_n860_), .A2(new_n3427_), .ZN(new_n3428_));
  INV_X1     g03162(.I(new_n3428_), .ZN(new_n3429_));
  NAND2_X1   g03163(.A1(new_n3424_), .A2(new_n3429_), .ZN(new_n3430_));
  AOI21_X1   g03164(.A1(new_n3409_), .A2(new_n3414_), .B(new_n3420_), .ZN(new_n3431_));
  INV_X1     g03165(.I(new_n3421_), .ZN(new_n3432_));
  OAI21_X1   g03166(.A1(new_n3411_), .A2(new_n3412_), .B(new_n3407_), .ZN(new_n3433_));
  AOI21_X1   g03167(.A1(new_n3432_), .A2(new_n3433_), .B(new_n3327_), .ZN(new_n3434_));
  NOR2_X1    g03168(.A1(new_n3431_), .A2(new_n3434_), .ZN(new_n3435_));
  NAND2_X1   g03169(.A1(new_n3435_), .A2(new_n3428_), .ZN(new_n3436_));
  NAND2_X1   g03170(.A1(new_n3436_), .A2(new_n3430_), .ZN(new_n3437_));
  OAI21_X1   g03171(.A1(new_n3165_), .A2(new_n3065_), .B(new_n3170_), .ZN(new_n3438_));
  OAI22_X1   g03172(.A1(new_n3438_), .A2(new_n3175_), .B1(new_n3066_), .B2(new_n3178_), .ZN(new_n3439_));
  OAI22_X1   g03173(.A1(new_n1055_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n1061_), .ZN(new_n3440_));
  OAI21_X1   g03174(.A1(new_n930_), .A2(new_n1332_), .B(new_n3440_), .ZN(new_n3441_));
  AOI21_X1   g03175(.A1(new_n3441_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n3442_));
  XOR2_X1    g03176(.A1(new_n1114_), .A2(new_n3442_), .Z(new_n3443_));
  INV_X1     g03177(.I(new_n3443_), .ZN(new_n3444_));
  XOR2_X1    g03178(.A1(new_n3439_), .A2(new_n3444_), .Z(new_n3445_));
  NAND2_X1   g03179(.A1(new_n3445_), .A2(new_n3437_), .ZN(new_n3446_));
  XOR2_X1    g03180(.A1(new_n3439_), .A2(new_n3444_), .Z(new_n3447_));
  OAI21_X1   g03181(.A1(new_n3437_), .A2(new_n3447_), .B(new_n3446_), .ZN(new_n3448_));
  OAI22_X1   g03182(.A1(new_n970_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n820_), .ZN(new_n3449_));
  OAI21_X1   g03183(.A1(new_n1189_), .A2(new_n894_), .B(new_n3449_), .ZN(new_n3450_));
  AOI21_X1   g03184(.A1(new_n3450_), .A2(new_n827_), .B(new_n970_), .ZN(new_n3451_));
  XNOR2_X1   g03185(.A1(new_n1421_), .A2(new_n3451_), .ZN(new_n3452_));
  INV_X1     g03186(.I(new_n3452_), .ZN(new_n3453_));
  XOR2_X1    g03187(.A1(new_n3448_), .A2(new_n3453_), .Z(new_n3454_));
  NOR2_X1    g03188(.A1(new_n3454_), .A2(new_n3323_), .ZN(new_n3455_));
  NAND2_X1   g03189(.A1(new_n3185_), .A2(new_n3057_), .ZN(new_n3456_));
  OAI21_X1   g03190(.A1(new_n3185_), .A2(new_n3057_), .B(new_n3190_), .ZN(new_n3457_));
  OAI21_X1   g03191(.A1(new_n3064_), .A2(new_n3457_), .B(new_n3456_), .ZN(new_n3458_));
  XOR2_X1    g03192(.A1(new_n3448_), .A2(new_n3452_), .Z(new_n3459_));
  NOR2_X1    g03193(.A1(new_n3459_), .A2(new_n3458_), .ZN(new_n3460_));
  NOR2_X1    g03194(.A1(new_n3455_), .A2(new_n3460_), .ZN(new_n3461_));
  OAI22_X1   g03195(.A1(new_n607_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n610_), .ZN(new_n3462_));
  OAI21_X1   g03196(.A1(new_n1525_), .A2(new_n684_), .B(new_n3462_), .ZN(new_n3463_));
  AOI21_X1   g03197(.A1(new_n3463_), .A2(new_n612_), .B(new_n607_), .ZN(new_n3464_));
  XOR2_X1    g03198(.A1(new_n1808_), .A2(new_n3464_), .Z(new_n3465_));
  XOR2_X1    g03199(.A1(new_n3461_), .A2(new_n3465_), .Z(new_n3466_));
  AOI21_X1   g03200(.A1(new_n3312_), .A2(new_n3317_), .B(new_n3466_), .ZN(new_n3467_));
  INV_X1     g03201(.I(new_n3206_), .ZN(new_n3468_));
  OAI21_X1   g03202(.A1(new_n3311_), .A2(new_n3212_), .B(new_n3468_), .ZN(new_n3469_));
  OAI21_X1   g03203(.A1(new_n3056_), .A2(new_n3469_), .B(new_n3312_), .ZN(new_n3470_));
  INV_X1     g03204(.I(new_n3465_), .ZN(new_n3471_));
  XOR2_X1    g03205(.A1(new_n3461_), .A2(new_n3471_), .Z(new_n3472_));
  NOR2_X1    g03206(.A1(new_n3472_), .A2(new_n3470_), .ZN(new_n3473_));
  NOR2_X1    g03207(.A1(new_n3467_), .A2(new_n3473_), .ZN(new_n3474_));
  OAI22_X1   g03208(.A1(new_n448_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n450_), .ZN(new_n3475_));
  OAI21_X1   g03209(.A1(new_n1936_), .A2(new_n496_), .B(new_n3475_), .ZN(new_n3476_));
  AOI21_X1   g03210(.A1(new_n3476_), .A2(new_n452_), .B(new_n448_), .ZN(new_n3477_));
  XNOR2_X1   g03211(.A1(new_n2280_), .A2(new_n3477_), .ZN(new_n3478_));
  XOR2_X1    g03212(.A1(new_n3474_), .A2(new_n3478_), .Z(new_n3479_));
  NOR2_X1    g03213(.A1(new_n3479_), .A2(new_n3308_), .ZN(new_n3480_));
  OAI21_X1   g03214(.A1(new_n3215_), .A2(new_n3049_), .B(new_n3220_), .ZN(new_n3481_));
  OAI22_X1   g03215(.A1(new_n3054_), .A2(new_n3481_), .B1(new_n3050_), .B2(new_n3305_), .ZN(new_n3482_));
  INV_X1     g03216(.I(new_n3478_), .ZN(new_n3483_));
  XOR2_X1    g03217(.A1(new_n3474_), .A2(new_n3483_), .Z(new_n3484_));
  NOR2_X1    g03218(.A1(new_n3484_), .A2(new_n3482_), .ZN(new_n3485_));
  NOR2_X1    g03219(.A1(new_n3480_), .A2(new_n3485_), .ZN(new_n3486_));
  OAI22_X1   g03220(.A1(new_n2643_), .A2(new_n341_), .B1(new_n404_), .B2(new_n2842_), .ZN(new_n3487_));
  OAI21_X1   g03221(.A1(new_n2439_), .A2(new_n366_), .B(new_n3487_), .ZN(new_n3488_));
  AOI21_X1   g03222(.A1(new_n3488_), .A2(new_n334_), .B(new_n341_), .ZN(new_n3489_));
  XNOR2_X1   g03223(.A1(new_n2846_), .A2(new_n3489_), .ZN(new_n3490_));
  NOR2_X1    g03224(.A1(new_n3486_), .A2(new_n3490_), .ZN(new_n3491_));
  INV_X1     g03225(.I(new_n3486_), .ZN(new_n3492_));
  INV_X1     g03226(.I(new_n3490_), .ZN(new_n3493_));
  NOR2_X1    g03227(.A1(new_n3492_), .A2(new_n3493_), .ZN(new_n3494_));
  OAI21_X1   g03228(.A1(new_n3494_), .A2(new_n3491_), .B(new_n3304_), .ZN(new_n3495_));
  INV_X1     g03229(.I(new_n3045_), .ZN(new_n3496_));
  AOI21_X1   g03230(.A1(new_n3223_), .A2(new_n3231_), .B(new_n3496_), .ZN(new_n3497_));
  NAND3_X1   g03231(.A1(new_n3496_), .A2(new_n3223_), .A3(new_n3231_), .ZN(new_n3498_));
  NOR3_X1    g03232(.A1(new_n3048_), .A2(new_n3046_), .A3(new_n3235_), .ZN(new_n3499_));
  AOI21_X1   g03233(.A1(new_n3499_), .A2(new_n3498_), .B(new_n3497_), .ZN(new_n3500_));
  NOR2_X1    g03234(.A1(new_n3492_), .A2(new_n3490_), .ZN(new_n3501_));
  NOR2_X1    g03235(.A1(new_n3486_), .A2(new_n3493_), .ZN(new_n3502_));
  OAI21_X1   g03236(.A1(new_n3501_), .A2(new_n3502_), .B(new_n3500_), .ZN(new_n3503_));
  NAND2_X1   g03237(.A1(new_n3503_), .A2(new_n3495_), .ZN(new_n3504_));
  INV_X1     g03238(.I(new_n3504_), .ZN(new_n3505_));
  NOR3_X1    g03239(.A1(new_n3247_), .A2(new_n3295_), .A3(new_n3505_), .ZN(new_n3506_));
  NOR2_X1    g03240(.A1(new_n3294_), .A2(new_n3246_), .ZN(new_n3507_));
  NOR2_X1    g03241(.A1(new_n3506_), .A2(new_n3507_), .ZN(new_n3508_));
  NOR2_X1    g03242(.A1(new_n3508_), .A2(new_n3252_), .ZN(new_n3509_));
  NOR3_X1    g03243(.A1(new_n3506_), .A2(new_n3275_), .A3(new_n3507_), .ZN(new_n3510_));
  NOR2_X1    g03244(.A1(new_n3509_), .A2(new_n3510_), .ZN(new_n3511_));
  XNOR2_X1   g03245(.A1(\b[29] ), .A2(\b[31] ), .ZN(new_n3512_));
  NOR2_X1    g03246(.A1(new_n3512_), .A2(new_n3259_), .ZN(new_n3513_));
  XNOR2_X1   g03247(.A1(new_n3258_), .A2(new_n3513_), .ZN(new_n3514_));
  NAND2_X1   g03248(.A1(new_n286_), .A2(\b[30] ), .ZN(new_n3515_));
  AOI22_X1   g03249(.A1(new_n304_), .A2(\b[29] ), .B1(new_n262_), .B2(\b[31] ), .ZN(new_n3516_));
  AOI21_X1   g03250(.A1(new_n3515_), .A2(new_n3516_), .B(new_n426_), .ZN(new_n3517_));
  NAND2_X1   g03251(.A1(new_n3514_), .A2(new_n3517_), .ZN(new_n3518_));
  XOR2_X1    g03252(.A1(new_n3518_), .A2(new_n260_), .Z(new_n3519_));
  XOR2_X1    g03253(.A1(new_n3518_), .A2(\a[2] ), .Z(new_n3520_));
  INV_X1     g03254(.I(new_n3520_), .ZN(new_n3521_));
  NAND2_X1   g03255(.A1(new_n3511_), .A2(new_n3521_), .ZN(new_n3522_));
  OAI21_X1   g03256(.A1(new_n3511_), .A2(new_n3519_), .B(new_n3522_), .ZN(new_n3523_));
  INV_X1     g03257(.I(new_n3279_), .ZN(new_n3524_));
  NAND2_X1   g03258(.A1(new_n3247_), .A2(new_n3252_), .ZN(new_n3525_));
  NAND2_X1   g03259(.A1(new_n3274_), .A2(new_n3275_), .ZN(new_n3526_));
  AOI21_X1   g03260(.A1(new_n3526_), .A2(new_n3525_), .B(new_n3269_), .ZN(new_n3527_));
  AOI21_X1   g03261(.A1(new_n3524_), .A2(new_n3527_), .B(new_n3289_), .ZN(new_n3528_));
  NOR2_X1    g03262(.A1(new_n3284_), .A2(new_n3528_), .ZN(new_n3529_));
  XOR2_X1    g03263(.A1(new_n3529_), .A2(new_n3523_), .Z(\f[31] ));
  NOR3_X1    g03264(.A1(new_n3284_), .A2(new_n3511_), .A3(new_n3528_), .ZN(new_n3531_));
  OAI21_X1   g03265(.A1(new_n3284_), .A2(new_n3528_), .B(new_n3511_), .ZN(new_n3532_));
  AOI21_X1   g03266(.A1(new_n3532_), .A2(new_n3521_), .B(new_n3531_), .ZN(new_n3533_));
  XOR2_X1    g03267(.A1(new_n3304_), .A2(new_n3492_), .Z(new_n3534_));
  NAND2_X1   g03268(.A1(new_n3534_), .A2(new_n3490_), .ZN(new_n3535_));
  INV_X1     g03269(.I(new_n3535_), .ZN(new_n3536_));
  INV_X1     g03270(.I(new_n3246_), .ZN(new_n3537_));
  AOI21_X1   g03271(.A1(new_n3242_), .A2(new_n3504_), .B(new_n3537_), .ZN(new_n3538_));
  OAI21_X1   g03272(.A1(new_n3242_), .A2(new_n3504_), .B(new_n3252_), .ZN(new_n3539_));
  NOR2_X1    g03273(.A1(new_n3539_), .A2(new_n3538_), .ZN(new_n3540_));
  XOR2_X1    g03274(.A1(new_n3482_), .A2(new_n3474_), .Z(new_n3541_));
  NOR2_X1    g03275(.A1(new_n3541_), .A2(new_n3483_), .ZN(new_n3542_));
  XOR2_X1    g03276(.A1(new_n3470_), .A2(new_n3461_), .Z(new_n3543_));
  NOR2_X1    g03277(.A1(new_n3543_), .A2(new_n3471_), .ZN(new_n3544_));
  OAI22_X1   g03278(.A1(new_n970_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n820_), .ZN(new_n3545_));
  OAI21_X1   g03279(.A1(new_n1294_), .A2(new_n894_), .B(new_n3545_), .ZN(new_n3546_));
  AOI21_X1   g03280(.A1(new_n3546_), .A2(new_n827_), .B(new_n970_), .ZN(new_n3547_));
  XOR2_X1    g03281(.A1(new_n1530_), .A2(new_n3547_), .Z(new_n3548_));
  INV_X1     g03282(.I(new_n3548_), .ZN(new_n3549_));
  XNOR2_X1   g03283(.A1(new_n3439_), .A2(new_n3437_), .ZN(new_n3550_));
  NAND2_X1   g03284(.A1(new_n3550_), .A2(new_n3443_), .ZN(new_n3551_));
  AOI21_X1   g03285(.A1(new_n3178_), .A2(new_n3066_), .B(new_n3169_), .ZN(new_n3552_));
  AOI22_X1   g03286(.A1(new_n3070_), .A2(new_n3552_), .B1(new_n3065_), .B2(new_n3165_), .ZN(new_n3553_));
  OAI22_X1   g03287(.A1(new_n1712_), .A2(new_n656_), .B1(new_n706_), .B2(new_n1707_), .ZN(new_n3554_));
  OAI21_X1   g03288(.A1(new_n565_), .A2(new_n1850_), .B(new_n3554_), .ZN(new_n3555_));
  AOI21_X1   g03289(.A1(new_n3555_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n3556_));
  XNOR2_X1   g03290(.A1(new_n710_), .A2(new_n3556_), .ZN(new_n3557_));
  INV_X1     g03291(.I(new_n3335_), .ZN(new_n3558_));
  INV_X1     g03292(.I(new_n3391_), .ZN(new_n3559_));
  OAI22_X1   g03293(.A1(new_n2171_), .A2(new_n472_), .B1(new_n515_), .B2(new_n2166_), .ZN(new_n3560_));
  OAI21_X1   g03294(.A1(new_n420_), .A2(new_n2322_), .B(new_n3560_), .ZN(new_n3561_));
  AOI21_X1   g03295(.A1(new_n3561_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n3562_));
  XOR2_X1    g03296(.A1(new_n700_), .A2(new_n3562_), .Z(new_n3563_));
  INV_X1     g03297(.I(new_n3563_), .ZN(new_n3564_));
  NAND2_X1   g03298(.A1(new_n3367_), .A2(new_n3373_), .ZN(new_n3565_));
  OAI21_X1   g03299(.A1(\b[1] ), .A2(new_n282_), .B(new_n3346_), .ZN(new_n3566_));
  OAI21_X1   g03300(.A1(new_n280_), .A2(new_n3352_), .B(new_n3566_), .ZN(new_n3567_));
  XOR2_X1    g03301(.A1(\a[29] ), .A2(\a[32] ), .Z(new_n3568_));
  NAND3_X1   g03302(.A1(new_n3356_), .A2(new_n3084_), .A3(new_n3568_), .ZN(new_n3569_));
  NOR2_X1    g03303(.A1(new_n3569_), .A2(new_n258_), .ZN(new_n3570_));
  AOI21_X1   g03304(.A1(new_n3567_), .A2(new_n3570_), .B(new_n3354_), .ZN(new_n3571_));
  NAND3_X1   g03305(.A1(new_n3567_), .A2(new_n3354_), .A3(new_n3570_), .ZN(new_n3572_));
  INV_X1     g03306(.I(new_n3572_), .ZN(new_n3573_));
  NOR2_X1    g03307(.A1(new_n3573_), .A2(new_n3571_), .ZN(new_n3574_));
  XOR2_X1    g03308(.A1(new_n3565_), .A2(new_n3574_), .Z(new_n3575_));
  AOI22_X1   g03309(.A1(new_n3338_), .A2(new_n3336_), .B1(new_n3343_), .B2(new_n3375_), .ZN(new_n3576_));
  NOR2_X1    g03310(.A1(new_n2333_), .A2(new_n2705_), .ZN(new_n3577_));
  OAI22_X1   g03311(.A1(new_n325_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n419_), .ZN(new_n3578_));
  OAI21_X1   g03312(.A1(new_n298_), .A2(new_n2884_), .B(new_n3578_), .ZN(new_n3579_));
  NOR2_X1    g03313(.A1(new_n3579_), .A2(new_n3577_), .ZN(new_n3580_));
  XOR2_X1    g03314(.A1(new_n3580_), .A2(new_n2702_), .Z(new_n3581_));
  NOR3_X1    g03315(.A1(new_n3576_), .A2(new_n3383_), .A3(new_n3581_), .ZN(new_n3582_));
  INV_X1     g03316(.I(new_n3383_), .ZN(new_n3583_));
  OAI22_X1   g03317(.A1(new_n3371_), .A2(new_n3369_), .B1(new_n3380_), .B2(new_n3378_), .ZN(new_n3584_));
  INV_X1     g03318(.I(new_n3581_), .ZN(new_n3585_));
  AOI21_X1   g03319(.A1(new_n3584_), .A2(new_n3583_), .B(new_n3585_), .ZN(new_n3586_));
  OAI21_X1   g03320(.A1(new_n3582_), .A2(new_n3586_), .B(new_n3575_), .ZN(new_n3587_));
  INV_X1     g03321(.I(new_n3575_), .ZN(new_n3588_));
  NAND3_X1   g03322(.A1(new_n3584_), .A2(new_n3583_), .A3(new_n3585_), .ZN(new_n3589_));
  OAI21_X1   g03323(.A1(new_n3576_), .A2(new_n3383_), .B(new_n3581_), .ZN(new_n3590_));
  NAND3_X1   g03324(.A1(new_n3590_), .A2(new_n3589_), .A3(new_n3588_), .ZN(new_n3591_));
  AOI21_X1   g03325(.A1(new_n3587_), .A2(new_n3591_), .B(new_n3564_), .ZN(new_n3592_));
  AOI21_X1   g03326(.A1(new_n3590_), .A2(new_n3589_), .B(new_n3588_), .ZN(new_n3593_));
  NOR3_X1    g03327(.A1(new_n3582_), .A2(new_n3586_), .A3(new_n3575_), .ZN(new_n3594_));
  NOR3_X1    g03328(.A1(new_n3594_), .A2(new_n3593_), .A3(new_n3563_), .ZN(new_n3595_));
  OAI21_X1   g03329(.A1(new_n3595_), .A2(new_n3592_), .B(new_n3401_), .ZN(new_n3596_));
  NOR2_X1    g03330(.A1(new_n3596_), .A2(new_n3559_), .ZN(new_n3597_));
  OAI21_X1   g03331(.A1(new_n3594_), .A2(new_n3593_), .B(new_n3563_), .ZN(new_n3598_));
  NAND3_X1   g03332(.A1(new_n3587_), .A2(new_n3591_), .A3(new_n3564_), .ZN(new_n3599_));
  NAND2_X1   g03333(.A1(new_n3598_), .A2(new_n3599_), .ZN(new_n3600_));
  INV_X1     g03334(.I(new_n3600_), .ZN(new_n3601_));
  NOR2_X1    g03335(.A1(new_n3395_), .A2(new_n3389_), .ZN(new_n3602_));
  OAI21_X1   g03336(.A1(new_n3597_), .A2(new_n3602_), .B(new_n3558_), .ZN(new_n3603_));
  NAND3_X1   g03337(.A1(new_n3600_), .A2(new_n3391_), .A3(new_n3401_), .ZN(new_n3604_));
  INV_X1     g03338(.I(new_n3602_), .ZN(new_n3605_));
  NAND3_X1   g03339(.A1(new_n3604_), .A2(new_n3335_), .A3(new_n3605_), .ZN(new_n3606_));
  NAND2_X1   g03340(.A1(new_n3603_), .A2(new_n3606_), .ZN(new_n3607_));
  OAI21_X1   g03341(.A1(new_n3419_), .A2(new_n3417_), .B(new_n3433_), .ZN(new_n3608_));
  OAI22_X1   g03342(.A1(new_n1347_), .A2(new_n861_), .B1(new_n930_), .B2(new_n1344_), .ZN(new_n3609_));
  OAI21_X1   g03343(.A1(new_n780_), .A2(new_n1457_), .B(new_n3609_), .ZN(new_n3610_));
  AOI21_X1   g03344(.A1(new_n3610_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n3611_));
  XNOR2_X1   g03345(.A1(new_n937_), .A2(new_n3611_), .ZN(new_n3612_));
  INV_X1     g03346(.I(new_n3612_), .ZN(new_n3613_));
  NAND3_X1   g03347(.A1(new_n3608_), .A2(new_n3432_), .A3(new_n3613_), .ZN(new_n3614_));
  AOI21_X1   g03348(.A1(new_n3326_), .A2(new_n3324_), .B(new_n3422_), .ZN(new_n3615_));
  OAI21_X1   g03349(.A1(new_n3615_), .A2(new_n3421_), .B(new_n3612_), .ZN(new_n3616_));
  AOI21_X1   g03350(.A1(new_n3616_), .A2(new_n3614_), .B(new_n3607_), .ZN(new_n3617_));
  AOI21_X1   g03351(.A1(new_n3604_), .A2(new_n3605_), .B(new_n3335_), .ZN(new_n3618_));
  NOR3_X1    g03352(.A1(new_n3597_), .A2(new_n3558_), .A3(new_n3602_), .ZN(new_n3619_));
  NOR2_X1    g03353(.A1(new_n3619_), .A2(new_n3618_), .ZN(new_n3620_));
  NOR3_X1    g03354(.A1(new_n3615_), .A2(new_n3421_), .A3(new_n3612_), .ZN(new_n3621_));
  AOI21_X1   g03355(.A1(new_n3608_), .A2(new_n3432_), .B(new_n3613_), .ZN(new_n3622_));
  NOR3_X1    g03356(.A1(new_n3621_), .A2(new_n3622_), .A3(new_n3620_), .ZN(new_n3623_));
  OAI21_X1   g03357(.A1(new_n3623_), .A2(new_n3617_), .B(new_n3557_), .ZN(new_n3624_));
  INV_X1     g03358(.I(new_n3557_), .ZN(new_n3625_));
  OAI21_X1   g03359(.A1(new_n3621_), .A2(new_n3622_), .B(new_n3620_), .ZN(new_n3626_));
  NAND3_X1   g03360(.A1(new_n3616_), .A2(new_n3614_), .A3(new_n3607_), .ZN(new_n3627_));
  NAND3_X1   g03361(.A1(new_n3626_), .A2(new_n3627_), .A3(new_n3625_), .ZN(new_n3628_));
  NAND2_X1   g03362(.A1(new_n3624_), .A2(new_n3628_), .ZN(new_n3629_));
  OAI21_X1   g03363(.A1(new_n3431_), .A2(new_n3434_), .B(new_n3428_), .ZN(new_n3630_));
  NAND3_X1   g03364(.A1(new_n3423_), .A2(new_n3416_), .A3(new_n3429_), .ZN(new_n3631_));
  NAND2_X1   g03365(.A1(new_n3630_), .A2(new_n3631_), .ZN(new_n3632_));
  AND3_X2    g03366(.A1(new_n3629_), .A2(new_n3430_), .A3(new_n3632_), .Z(new_n3633_));
  NAND2_X1   g03367(.A1(new_n3424_), .A2(new_n3429_), .ZN(new_n3635_));
  INV_X1     g03368(.I(new_n3635_), .ZN(new_n3636_));
  OAI21_X1   g03369(.A1(new_n3633_), .A2(new_n3636_), .B(new_n3553_), .ZN(new_n3637_));
  NAND3_X1   g03370(.A1(new_n3629_), .A2(new_n3430_), .A3(new_n3632_), .ZN(new_n3638_));
  NAND3_X1   g03371(.A1(new_n3638_), .A2(new_n3439_), .A3(new_n3635_), .ZN(new_n3639_));
  OAI22_X1   g03372(.A1(new_n1055_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n1061_), .ZN(new_n3640_));
  OAI21_X1   g03373(.A1(new_n1017_), .A2(new_n1332_), .B(new_n3640_), .ZN(new_n3641_));
  AOI21_X1   g03374(.A1(new_n3641_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n3642_));
  XNOR2_X1   g03375(.A1(new_n1196_), .A2(new_n3642_), .ZN(new_n3643_));
  INV_X1     g03376(.I(new_n3643_), .ZN(new_n3644_));
  NAND3_X1   g03377(.A1(new_n3637_), .A2(new_n3639_), .A3(new_n3644_), .ZN(new_n3645_));
  AOI21_X1   g03378(.A1(new_n3638_), .A2(new_n3635_), .B(new_n3439_), .ZN(new_n3646_));
  INV_X1     g03379(.I(new_n3639_), .ZN(new_n3647_));
  OAI21_X1   g03380(.A1(new_n3647_), .A2(new_n3646_), .B(new_n3643_), .ZN(new_n3648_));
  NAND3_X1   g03381(.A1(new_n3648_), .A2(new_n3645_), .A3(new_n3551_), .ZN(new_n3649_));
  NAND2_X1   g03382(.A1(new_n3649_), .A2(new_n3448_), .ZN(new_n3650_));
  NOR2_X1    g03383(.A1(new_n3650_), .A2(new_n3458_), .ZN(new_n3651_));
  AOI21_X1   g03384(.A1(new_n3649_), .A2(new_n3448_), .B(new_n3323_), .ZN(new_n3652_));
  NOR2_X1    g03385(.A1(new_n3651_), .A2(new_n3652_), .ZN(new_n3653_));
  XOR2_X1    g03386(.A1(new_n3448_), .A2(new_n3323_), .Z(new_n3654_));
  NOR2_X1    g03387(.A1(new_n3654_), .A2(new_n3453_), .ZN(new_n3655_));
  INV_X1     g03388(.I(new_n3655_), .ZN(new_n3656_));
  NAND3_X1   g03389(.A1(new_n3317_), .A2(new_n3461_), .A3(new_n3312_), .ZN(new_n3657_));
  OAI22_X1   g03390(.A1(new_n607_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n610_), .ZN(new_n3658_));
  OAI21_X1   g03391(.A1(new_n1634_), .A2(new_n684_), .B(new_n3658_), .ZN(new_n3659_));
  AOI21_X1   g03392(.A1(new_n3659_), .A2(new_n612_), .B(new_n607_), .ZN(new_n3660_));
  XNOR2_X1   g03393(.A1(new_n1940_), .A2(new_n3660_), .ZN(new_n3661_));
  AOI21_X1   g03394(.A1(new_n3657_), .A2(new_n3656_), .B(new_n3661_), .ZN(new_n3662_));
  XOR2_X1    g03395(.A1(new_n3448_), .A2(new_n3452_), .Z(new_n3663_));
  NAND2_X1   g03396(.A1(new_n3663_), .A2(new_n3458_), .ZN(new_n3664_));
  OAI21_X1   g03397(.A1(new_n3458_), .A2(new_n3459_), .B(new_n3664_), .ZN(new_n3665_));
  OAI21_X1   g03398(.A1(new_n3470_), .A2(new_n3665_), .B(new_n3656_), .ZN(new_n3666_));
  INV_X1     g03399(.I(new_n3661_), .ZN(new_n3667_));
  NOR2_X1    g03400(.A1(new_n3666_), .A2(new_n3667_), .ZN(new_n3668_));
  OAI21_X1   g03401(.A1(new_n3662_), .A2(new_n3668_), .B(new_n3653_), .ZN(new_n3669_));
  INV_X1     g03402(.I(new_n3653_), .ZN(new_n3670_));
  NAND2_X1   g03403(.A1(new_n3666_), .A2(new_n3667_), .ZN(new_n3671_));
  NAND3_X1   g03404(.A1(new_n3657_), .A2(new_n3656_), .A3(new_n3661_), .ZN(new_n3672_));
  NAND3_X1   g03405(.A1(new_n3672_), .A2(new_n3671_), .A3(new_n3670_), .ZN(new_n3673_));
  AOI21_X1   g03406(.A1(new_n3669_), .A2(new_n3673_), .B(new_n3549_), .ZN(new_n3674_));
  AOI21_X1   g03407(.A1(new_n3672_), .A2(new_n3671_), .B(new_n3670_), .ZN(new_n3675_));
  NOR3_X1    g03408(.A1(new_n3662_), .A2(new_n3668_), .A3(new_n3653_), .ZN(new_n3676_));
  NOR3_X1    g03409(.A1(new_n3675_), .A2(new_n3676_), .A3(new_n3548_), .ZN(new_n3677_));
  NOR3_X1    g03410(.A1(new_n3677_), .A2(new_n3674_), .A3(new_n3544_), .ZN(new_n3678_));
  NOR3_X1    g03411(.A1(new_n3678_), .A2(new_n3482_), .A3(new_n3474_), .ZN(new_n3679_));
  INV_X1     g03412(.I(new_n3679_), .ZN(new_n3680_));
  OAI21_X1   g03413(.A1(new_n3678_), .A2(new_n3474_), .B(new_n3482_), .ZN(new_n3681_));
  OAI22_X1   g03414(.A1(new_n448_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n450_), .ZN(new_n3682_));
  OAI21_X1   g03415(.A1(new_n2102_), .A2(new_n496_), .B(new_n3682_), .ZN(new_n3683_));
  AOI21_X1   g03416(.A1(new_n3683_), .A2(new_n452_), .B(new_n448_), .ZN(new_n3684_));
  XNOR2_X1   g03417(.A1(new_n2443_), .A2(new_n3684_), .ZN(new_n3685_));
  INV_X1     g03418(.I(new_n3685_), .ZN(new_n3686_));
  NAND3_X1   g03419(.A1(new_n3680_), .A2(new_n3681_), .A3(new_n3686_), .ZN(new_n3687_));
  INV_X1     g03420(.I(new_n3687_), .ZN(new_n3688_));
  AOI21_X1   g03421(.A1(new_n3680_), .A2(new_n3681_), .B(new_n3686_), .ZN(new_n3689_));
  NOR3_X1    g03422(.A1(new_n3542_), .A2(new_n3688_), .A3(new_n3689_), .ZN(new_n3690_));
  NOR2_X1    g03423(.A1(new_n3690_), .A2(new_n3486_), .ZN(new_n3691_));
  NAND2_X1   g03424(.A1(new_n3691_), .A2(new_n3500_), .ZN(new_n3692_));
  OAI21_X1   g03425(.A1(new_n3690_), .A2(new_n3486_), .B(new_n3304_), .ZN(new_n3693_));
  OAI22_X1   g03426(.A1(new_n2842_), .A2(new_n341_), .B1(new_n404_), .B2(new_n3018_), .ZN(new_n3694_));
  OAI21_X1   g03427(.A1(new_n2643_), .A2(new_n366_), .B(new_n3694_), .ZN(new_n3695_));
  AOI21_X1   g03428(.A1(new_n3695_), .A2(new_n334_), .B(new_n341_), .ZN(new_n3696_));
  XNOR2_X1   g03429(.A1(new_n3022_), .A2(new_n3696_), .ZN(new_n3697_));
  AOI21_X1   g03430(.A1(new_n3692_), .A2(new_n3693_), .B(new_n3697_), .ZN(new_n3698_));
  INV_X1     g03431(.I(new_n3698_), .ZN(new_n3699_));
  NOR2_X1    g03432(.A1(new_n3540_), .A2(new_n3699_), .ZN(new_n3700_));
  INV_X1     g03433(.I(new_n3700_), .ZN(new_n3701_));
  NAND2_X1   g03434(.A1(new_n3540_), .A2(new_n3699_), .ZN(new_n3702_));
  AOI21_X1   g03435(.A1(new_n3701_), .A2(new_n3702_), .B(new_n3536_), .ZN(new_n3703_));
  NAND3_X1   g03436(.A1(new_n3701_), .A2(new_n3702_), .A3(new_n3536_), .ZN(new_n3704_));
  INV_X1     g03437(.I(new_n3704_), .ZN(new_n3705_));
  NOR2_X1    g03438(.A1(new_n3705_), .A2(new_n3703_), .ZN(new_n3706_));
  NOR2_X1    g03439(.A1(\b[30] ), .A2(\b[31] ), .ZN(new_n3707_));
  AOI21_X1   g03440(.A1(new_n3258_), .A2(new_n3707_), .B(new_n3018_), .ZN(new_n3708_));
  INV_X1     g03441(.I(\b[31] ), .ZN(new_n3709_));
  NOR2_X1    g03442(.A1(new_n3260_), .A2(new_n3709_), .ZN(new_n3710_));
  INV_X1     g03443(.I(new_n3710_), .ZN(new_n3711_));
  NOR2_X1    g03444(.A1(new_n3258_), .A2(new_n3711_), .ZN(new_n3712_));
  NOR2_X1    g03445(.A1(new_n3708_), .A2(new_n3712_), .ZN(new_n3713_));
  INV_X1     g03446(.I(new_n3713_), .ZN(new_n3714_));
  XNOR2_X1   g03447(.A1(\b[31] ), .A2(\b[32] ), .ZN(new_n3715_));
  INV_X1     g03448(.I(new_n3715_), .ZN(new_n3716_));
  INV_X1     g03449(.I(\b[32] ), .ZN(new_n3717_));
  NOR2_X1    g03450(.A1(new_n3709_), .A2(new_n3717_), .ZN(new_n3718_));
  INV_X1     g03451(.I(new_n3718_), .ZN(new_n3719_));
  NAND2_X1   g03452(.A1(new_n3709_), .A2(new_n3717_), .ZN(new_n3720_));
  AOI21_X1   g03453(.A1(new_n3719_), .A2(new_n3720_), .B(new_n3714_), .ZN(new_n3721_));
  AOI21_X1   g03454(.A1(new_n3714_), .A2(new_n3716_), .B(new_n3721_), .ZN(new_n3722_));
  OAI22_X1   g03455(.A1(new_n330_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n263_), .ZN(new_n3723_));
  OAI21_X1   g03456(.A1(new_n3260_), .A2(new_n289_), .B(new_n3723_), .ZN(new_n3724_));
  AOI21_X1   g03457(.A1(new_n3724_), .A2(new_n260_), .B(new_n426_), .ZN(new_n3725_));
  XOR2_X1    g03458(.A1(new_n3722_), .A2(new_n3725_), .Z(new_n3726_));
  INV_X1     g03459(.I(new_n3726_), .ZN(new_n3727_));
  XOR2_X1    g03460(.A1(new_n3706_), .A2(new_n3727_), .Z(new_n3728_));
  INV_X1     g03461(.I(new_n3706_), .ZN(new_n3729_));
  NAND2_X1   g03462(.A1(new_n3729_), .A2(new_n3727_), .ZN(new_n3730_));
  NAND2_X1   g03463(.A1(new_n3706_), .A2(new_n3726_), .ZN(new_n3731_));
  NAND2_X1   g03464(.A1(new_n3730_), .A2(new_n3731_), .ZN(new_n3732_));
  NAND2_X1   g03465(.A1(new_n3533_), .A2(new_n3732_), .ZN(new_n3733_));
  OAI21_X1   g03466(.A1(new_n3533_), .A2(new_n3728_), .B(new_n3733_), .ZN(\f[32] ));
  AOI21_X1   g03467(.A1(new_n3693_), .A2(new_n3692_), .B(new_n3535_), .ZN(new_n3735_));
  NAND3_X1   g03468(.A1(new_n3535_), .A2(new_n3692_), .A3(new_n3693_), .ZN(new_n3736_));
  NOR3_X1    g03469(.A1(new_n3539_), .A2(new_n3538_), .A3(new_n3697_), .ZN(new_n3737_));
  AOI21_X1   g03470(.A1(new_n3737_), .A2(new_n3736_), .B(new_n3735_), .ZN(new_n3738_));
  INV_X1     g03471(.I(new_n3738_), .ZN(new_n3739_));
  INV_X1     g03472(.I(new_n3681_), .ZN(new_n3740_));
  OAI21_X1   g03473(.A1(new_n3740_), .A2(new_n3679_), .B(new_n3685_), .ZN(new_n3741_));
  OAI21_X1   g03474(.A1(new_n3688_), .A2(new_n3689_), .B(new_n3542_), .ZN(new_n3742_));
  AOI21_X1   g03475(.A1(new_n3742_), .A2(new_n3486_), .B(new_n3500_), .ZN(new_n3743_));
  AOI21_X1   g03476(.A1(new_n3657_), .A2(new_n3656_), .B(new_n3653_), .ZN(new_n3744_));
  NOR2_X1    g03477(.A1(new_n3666_), .A2(new_n3670_), .ZN(new_n3745_));
  OAI21_X1   g03478(.A1(new_n3744_), .A2(new_n3745_), .B(new_n3548_), .ZN(new_n3746_));
  NOR3_X1    g03479(.A1(new_n3744_), .A2(new_n3745_), .A3(new_n3548_), .ZN(new_n3747_));
  INV_X1     g03480(.I(new_n3747_), .ZN(new_n3748_));
  AOI21_X1   g03481(.A1(new_n3748_), .A2(new_n3746_), .B(new_n3661_), .ZN(new_n3749_));
  INV_X1     g03482(.I(new_n3749_), .ZN(new_n3750_));
  OAI21_X1   g03483(.A1(new_n3677_), .A2(new_n3674_), .B(new_n3544_), .ZN(new_n3751_));
  AOI21_X1   g03484(.A1(new_n3751_), .A2(new_n3474_), .B(new_n3308_), .ZN(new_n3752_));
  NOR2_X1    g03485(.A1(new_n3653_), .A2(new_n3549_), .ZN(new_n3753_));
  OAI21_X1   g03486(.A1(new_n3651_), .A2(new_n3652_), .B(new_n3549_), .ZN(new_n3754_));
  NOR3_X1    g03487(.A1(new_n3651_), .A2(new_n3549_), .A3(new_n3652_), .ZN(new_n3755_));
  INV_X1     g03488(.I(new_n3755_), .ZN(new_n3756_));
  AOI21_X1   g03489(.A1(new_n3754_), .A2(new_n3756_), .B(new_n3656_), .ZN(new_n3757_));
  OAI21_X1   g03490(.A1(new_n3757_), .A2(new_n3665_), .B(new_n3470_), .ZN(new_n3758_));
  AOI21_X1   g03491(.A1(new_n3648_), .A2(new_n3645_), .B(new_n3551_), .ZN(new_n3759_));
  OAI21_X1   g03492(.A1(new_n3759_), .A2(new_n3448_), .B(new_n3458_), .ZN(new_n3760_));
  NOR2_X1    g03493(.A1(new_n3615_), .A2(new_n3421_), .ZN(new_n3761_));
  NAND2_X1   g03494(.A1(new_n3761_), .A2(new_n3607_), .ZN(new_n3762_));
  NAND2_X1   g03495(.A1(new_n3608_), .A2(new_n3432_), .ZN(new_n3763_));
  NAND2_X1   g03496(.A1(new_n3763_), .A2(new_n3620_), .ZN(new_n3764_));
  AOI21_X1   g03497(.A1(new_n3762_), .A2(new_n3764_), .B(new_n3625_), .ZN(new_n3765_));
  NOR2_X1    g03498(.A1(new_n3763_), .A2(new_n3620_), .ZN(new_n3766_));
  NOR2_X1    g03499(.A1(new_n3761_), .A2(new_n3607_), .ZN(new_n3767_));
  NOR3_X1    g03500(.A1(new_n3767_), .A2(new_n3766_), .A3(new_n3557_), .ZN(new_n3768_));
  OAI21_X1   g03501(.A1(new_n3765_), .A2(new_n3768_), .B(new_n3613_), .ZN(new_n3769_));
  AOI21_X1   g03502(.A1(new_n3626_), .A2(new_n3627_), .B(new_n3625_), .ZN(new_n3770_));
  NOR3_X1    g03503(.A1(new_n3623_), .A2(new_n3617_), .A3(new_n3557_), .ZN(new_n3771_));
  OAI21_X1   g03504(.A1(new_n3771_), .A2(new_n3770_), .B(new_n3424_), .ZN(new_n3772_));
  NAND2_X1   g03505(.A1(new_n3772_), .A2(new_n3428_), .ZN(new_n3773_));
  NOR3_X1    g03506(.A1(new_n3771_), .A2(new_n3770_), .A3(new_n3424_), .ZN(new_n3774_));
  NOR2_X1    g03507(.A1(new_n3553_), .A2(new_n3774_), .ZN(new_n3775_));
  NOR2_X1    g03508(.A1(new_n3620_), .A2(new_n3625_), .ZN(new_n3776_));
  OAI21_X1   g03509(.A1(new_n3619_), .A2(new_n3618_), .B(new_n3625_), .ZN(new_n3777_));
  NAND3_X1   g03510(.A1(new_n3603_), .A2(new_n3606_), .A3(new_n3557_), .ZN(new_n3778_));
  NAND2_X1   g03511(.A1(new_n3777_), .A2(new_n3778_), .ZN(new_n3779_));
  AOI21_X1   g03512(.A1(new_n3779_), .A2(new_n3403_), .B(new_n3408_), .ZN(new_n3780_));
  NAND3_X1   g03513(.A1(new_n3777_), .A2(new_n3778_), .A3(new_n3413_), .ZN(new_n3781_));
  NAND2_X1   g03514(.A1(new_n3781_), .A2(new_n3327_), .ZN(new_n3782_));
  NAND2_X1   g03515(.A1(new_n3584_), .A2(new_n3583_), .ZN(new_n3783_));
  XOR2_X1    g03516(.A1(new_n3783_), .A2(new_n3588_), .Z(new_n3784_));
  NAND2_X1   g03517(.A1(new_n3784_), .A2(new_n3581_), .ZN(new_n3785_));
  XOR2_X1    g03518(.A1(new_n3783_), .A2(new_n3575_), .Z(new_n3786_));
  NAND2_X1   g03519(.A1(new_n3786_), .A2(new_n3585_), .ZN(new_n3787_));
  AOI21_X1   g03520(.A1(new_n3785_), .A2(new_n3787_), .B(new_n3563_), .ZN(new_n3788_));
  INV_X1     g03521(.I(new_n3788_), .ZN(new_n3789_));
  AOI21_X1   g03522(.A1(new_n3600_), .A2(new_n3385_), .B(new_n3390_), .ZN(new_n3790_));
  OAI21_X1   g03523(.A1(new_n3385_), .A2(new_n3600_), .B(new_n3335_), .ZN(new_n3791_));
  NOR2_X1    g03524(.A1(new_n3791_), .A2(new_n3790_), .ZN(new_n3792_));
  XOR2_X1    g03525(.A1(\a[32] ), .A2(\a[33] ), .Z(new_n3793_));
  NAND2_X1   g03526(.A1(new_n3793_), .A2(\b[0] ), .ZN(new_n3794_));
  NOR2_X1    g03527(.A1(new_n3569_), .A2(new_n269_), .ZN(new_n3795_));
  OAI22_X1   g03528(.A1(new_n298_), .A2(new_n3352_), .B1(new_n3357_), .B2(new_n280_), .ZN(new_n3796_));
  NOR2_X1    g03529(.A1(new_n3796_), .A2(new_n3795_), .ZN(new_n3797_));
  NAND2_X1   g03530(.A1(new_n301_), .A2(new_n3346_), .ZN(new_n3798_));
  OAI21_X1   g03531(.A1(new_n3797_), .A2(new_n3798_), .B(\a[32] ), .ZN(new_n3799_));
  NOR3_X1    g03532(.A1(new_n3797_), .A2(\a[32] ), .A3(new_n3798_), .ZN(new_n3800_));
  INV_X1     g03533(.I(new_n3800_), .ZN(new_n3801_));
  NAND2_X1   g03534(.A1(new_n3801_), .A2(new_n3799_), .ZN(new_n3802_));
  NOR2_X1    g03535(.A1(new_n3372_), .A2(new_n3363_), .ZN(new_n3803_));
  NAND2_X1   g03536(.A1(new_n3803_), .A2(new_n3574_), .ZN(new_n3804_));
  OAI22_X1   g03537(.A1(new_n420_), .A2(new_n2700_), .B1(new_n2705_), .B2(new_n419_), .ZN(new_n3805_));
  OAI21_X1   g03538(.A1(new_n325_), .A2(new_n2884_), .B(new_n3805_), .ZN(new_n3806_));
  AOI21_X1   g03539(.A1(new_n3806_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n3807_));
  INV_X1     g03540(.I(new_n3807_), .ZN(new_n3808_));
  NOR2_X1    g03541(.A1(new_n556_), .A2(new_n3808_), .ZN(new_n3809_));
  NOR2_X1    g03542(.A1(new_n425_), .A2(new_n3807_), .ZN(new_n3810_));
  OAI21_X1   g03543(.A1(new_n3809_), .A2(new_n3810_), .B(new_n3804_), .ZN(new_n3811_));
  INV_X1     g03544(.I(new_n3571_), .ZN(new_n3812_));
  NAND2_X1   g03545(.A1(new_n3812_), .A2(new_n3572_), .ZN(new_n3813_));
  NOR2_X1    g03546(.A1(new_n3565_), .A2(new_n3813_), .ZN(new_n3814_));
  NOR2_X1    g03547(.A1(new_n3810_), .A2(new_n3809_), .ZN(new_n3815_));
  NAND2_X1   g03548(.A1(new_n3815_), .A2(new_n3814_), .ZN(new_n3816_));
  AOI21_X1   g03549(.A1(new_n3816_), .A2(new_n3811_), .B(new_n3802_), .ZN(new_n3817_));
  INV_X1     g03550(.I(new_n3799_), .ZN(new_n3818_));
  NOR2_X1    g03551(.A1(new_n3818_), .A2(new_n3800_), .ZN(new_n3819_));
  NOR2_X1    g03552(.A1(new_n3815_), .A2(new_n3814_), .ZN(new_n3820_));
  NOR3_X1    g03553(.A1(new_n3804_), .A2(new_n3809_), .A3(new_n3810_), .ZN(new_n3821_));
  NOR3_X1    g03554(.A1(new_n3820_), .A2(new_n3821_), .A3(new_n3819_), .ZN(new_n3822_));
  OAI21_X1   g03555(.A1(new_n3817_), .A2(new_n3822_), .B(new_n3794_), .ZN(new_n3823_));
  INV_X1     g03556(.I(new_n3794_), .ZN(new_n3824_));
  OAI21_X1   g03557(.A1(new_n3820_), .A2(new_n3821_), .B(new_n3819_), .ZN(new_n3825_));
  NAND3_X1   g03558(.A1(new_n3816_), .A2(new_n3811_), .A3(new_n3802_), .ZN(new_n3826_));
  NAND3_X1   g03559(.A1(new_n3826_), .A2(new_n3825_), .A3(new_n3824_), .ZN(new_n3827_));
  NAND2_X1   g03560(.A1(new_n3823_), .A2(new_n3827_), .ZN(new_n3828_));
  NOR2_X1    g03561(.A1(new_n3575_), .A2(new_n3585_), .ZN(new_n3829_));
  INV_X1     g03562(.I(new_n3829_), .ZN(new_n3830_));
  INV_X1     g03563(.I(new_n3580_), .ZN(new_n3831_));
  NOR2_X1    g03564(.A1(new_n3803_), .A2(new_n3831_), .ZN(new_n3832_));
  NOR2_X1    g03565(.A1(new_n3565_), .A2(new_n3580_), .ZN(new_n3833_));
  OAI21_X1   g03566(.A1(new_n3832_), .A2(new_n3833_), .B(new_n3574_), .ZN(new_n3834_));
  NAND2_X1   g03567(.A1(new_n3565_), .A2(new_n3580_), .ZN(new_n3835_));
  NAND2_X1   g03568(.A1(new_n3803_), .A2(new_n3831_), .ZN(new_n3836_));
  NAND3_X1   g03569(.A1(new_n3836_), .A2(new_n3835_), .A3(new_n3813_), .ZN(new_n3837_));
  AOI21_X1   g03570(.A1(new_n3834_), .A2(new_n3837_), .B(\a[29] ), .ZN(new_n3838_));
  AOI21_X1   g03571(.A1(new_n3836_), .A2(new_n3835_), .B(new_n3813_), .ZN(new_n3839_));
  NOR3_X1    g03572(.A1(new_n3832_), .A2(new_n3833_), .A3(new_n3574_), .ZN(new_n3840_));
  NOR3_X1    g03573(.A1(new_n3839_), .A2(new_n3840_), .A3(new_n2702_), .ZN(new_n3841_));
  OAI21_X1   g03574(.A1(new_n3841_), .A2(new_n3838_), .B(new_n3375_), .ZN(new_n3842_));
  NAND2_X1   g03575(.A1(new_n3842_), .A2(new_n3343_), .ZN(new_n3843_));
  OAI21_X1   g03576(.A1(new_n3839_), .A2(new_n3840_), .B(new_n2702_), .ZN(new_n3844_));
  NAND3_X1   g03577(.A1(new_n3834_), .A2(new_n3837_), .A3(\a[29] ), .ZN(new_n3845_));
  NAND3_X1   g03578(.A1(new_n3844_), .A2(new_n3845_), .A3(new_n3369_), .ZN(new_n3846_));
  NAND3_X1   g03579(.A1(new_n3843_), .A2(new_n3339_), .A3(new_n3846_), .ZN(new_n3847_));
  AOI21_X1   g03580(.A1(new_n3847_), .A2(new_n3830_), .B(new_n3828_), .ZN(new_n3848_));
  INV_X1     g03581(.I(new_n3828_), .ZN(new_n3849_));
  NAND2_X1   g03582(.A1(new_n3844_), .A2(new_n3845_), .ZN(new_n3850_));
  AOI21_X1   g03583(.A1(new_n3850_), .A2(new_n3375_), .B(new_n3371_), .ZN(new_n3851_));
  NAND2_X1   g03584(.A1(new_n3846_), .A2(new_n3339_), .ZN(new_n3852_));
  NOR2_X1    g03585(.A1(new_n3851_), .A2(new_n3852_), .ZN(new_n3853_));
  NOR3_X1    g03586(.A1(new_n3853_), .A2(new_n3849_), .A3(new_n3829_), .ZN(new_n3854_));
  OAI22_X1   g03587(.A1(new_n2171_), .A2(new_n515_), .B1(new_n565_), .B2(new_n2166_), .ZN(new_n3855_));
  OAI21_X1   g03588(.A1(new_n472_), .A2(new_n2322_), .B(new_n3855_), .ZN(new_n3856_));
  AOI21_X1   g03589(.A1(new_n3856_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n3857_));
  XOR2_X1    g03590(.A1(new_n759_), .A2(new_n3857_), .Z(new_n3858_));
  INV_X1     g03591(.I(new_n3858_), .ZN(new_n3859_));
  OAI21_X1   g03592(.A1(new_n3848_), .A2(new_n3854_), .B(new_n3859_), .ZN(new_n3860_));
  NOR2_X1    g03593(.A1(new_n3792_), .A2(new_n3860_), .ZN(new_n3861_));
  OAI21_X1   g03594(.A1(new_n3853_), .A2(new_n3829_), .B(new_n3849_), .ZN(new_n3862_));
  NAND3_X1   g03595(.A1(new_n3847_), .A2(new_n3828_), .A3(new_n3830_), .ZN(new_n3863_));
  AOI21_X1   g03596(.A1(new_n3862_), .A2(new_n3863_), .B(new_n3858_), .ZN(new_n3864_));
  NOR3_X1    g03597(.A1(new_n3864_), .A2(new_n3791_), .A3(new_n3790_), .ZN(new_n3865_));
  OAI21_X1   g03598(.A1(new_n3861_), .A2(new_n3865_), .B(new_n3789_), .ZN(new_n3866_));
  OAI21_X1   g03599(.A1(new_n3790_), .A2(new_n3791_), .B(new_n3864_), .ZN(new_n3867_));
  INV_X1     g03600(.I(new_n3790_), .ZN(new_n3868_));
  NAND2_X1   g03601(.A1(new_n3601_), .A2(new_n3395_), .ZN(new_n3869_));
  NAND4_X1   g03602(.A1(new_n3860_), .A2(new_n3868_), .A3(new_n3869_), .A4(new_n3335_), .ZN(new_n3870_));
  NAND3_X1   g03603(.A1(new_n3870_), .A2(new_n3867_), .A3(new_n3788_), .ZN(new_n3871_));
  OAI22_X1   g03604(.A1(new_n1712_), .A2(new_n706_), .B1(new_n780_), .B2(new_n1707_), .ZN(new_n3872_));
  OAI21_X1   g03605(.A1(new_n656_), .A2(new_n1850_), .B(new_n3872_), .ZN(new_n3873_));
  AOI21_X1   g03606(.A1(new_n3873_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n3874_));
  XOR2_X1    g03607(.A1(new_n785_), .A2(new_n3874_), .Z(new_n3875_));
  AOI21_X1   g03608(.A1(new_n3866_), .A2(new_n3871_), .B(new_n3875_), .ZN(new_n3876_));
  OAI21_X1   g03609(.A1(new_n3780_), .A2(new_n3782_), .B(new_n3876_), .ZN(new_n3877_));
  AOI21_X1   g03610(.A1(new_n3603_), .A2(new_n3606_), .B(new_n3557_), .ZN(new_n3878_));
  NOR3_X1    g03611(.A1(new_n3619_), .A2(new_n3618_), .A3(new_n3625_), .ZN(new_n3879_));
  OAI21_X1   g03612(.A1(new_n3879_), .A2(new_n3878_), .B(new_n3403_), .ZN(new_n3880_));
  NAND2_X1   g03613(.A1(new_n3880_), .A2(new_n3407_), .ZN(new_n3881_));
  AOI21_X1   g03614(.A1(new_n3870_), .A2(new_n3867_), .B(new_n3788_), .ZN(new_n3882_));
  NOR3_X1    g03615(.A1(new_n3861_), .A2(new_n3789_), .A3(new_n3865_), .ZN(new_n3883_));
  INV_X1     g03616(.I(new_n3875_), .ZN(new_n3884_));
  OAI21_X1   g03617(.A1(new_n3883_), .A2(new_n3882_), .B(new_n3884_), .ZN(new_n3885_));
  NAND4_X1   g03618(.A1(new_n3881_), .A2(new_n3885_), .A3(new_n3327_), .A4(new_n3781_), .ZN(new_n3886_));
  AOI21_X1   g03619(.A1(new_n3886_), .A2(new_n3877_), .B(new_n3776_), .ZN(new_n3887_));
  NAND2_X1   g03620(.A1(new_n3607_), .A2(new_n3557_), .ZN(new_n3888_));
  NOR2_X1    g03621(.A1(new_n3780_), .A2(new_n3782_), .ZN(new_n3889_));
  NOR2_X1    g03622(.A1(new_n3889_), .A2(new_n3885_), .ZN(new_n3890_));
  NOR3_X1    g03623(.A1(new_n3780_), .A2(new_n3876_), .A3(new_n3782_), .ZN(new_n3891_));
  NOR3_X1    g03624(.A1(new_n3890_), .A2(new_n3888_), .A3(new_n3891_), .ZN(new_n3892_));
  OAI22_X1   g03625(.A1(new_n1347_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n1344_), .ZN(new_n3893_));
  OAI21_X1   g03626(.A1(new_n861_), .A2(new_n1457_), .B(new_n3893_), .ZN(new_n3894_));
  AOI21_X1   g03627(.A1(new_n3894_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n3895_));
  XOR2_X1    g03628(.A1(new_n1024_), .A2(new_n3895_), .Z(new_n3896_));
  INV_X1     g03629(.I(new_n3896_), .ZN(new_n3897_));
  OAI21_X1   g03630(.A1(new_n3892_), .A2(new_n3887_), .B(new_n3897_), .ZN(new_n3898_));
  AOI21_X1   g03631(.A1(new_n3775_), .A2(new_n3773_), .B(new_n3898_), .ZN(new_n3899_));
  AOI21_X1   g03632(.A1(new_n3629_), .A2(new_n3424_), .B(new_n3429_), .ZN(new_n3900_));
  NAND3_X1   g03633(.A1(new_n3624_), .A2(new_n3628_), .A3(new_n3435_), .ZN(new_n3901_));
  NAND2_X1   g03634(.A1(new_n3439_), .A2(new_n3901_), .ZN(new_n3902_));
  OAI21_X1   g03635(.A1(new_n3890_), .A2(new_n3891_), .B(new_n3888_), .ZN(new_n3903_));
  NAND3_X1   g03636(.A1(new_n3886_), .A2(new_n3877_), .A3(new_n3776_), .ZN(new_n3904_));
  AOI21_X1   g03637(.A1(new_n3903_), .A2(new_n3904_), .B(new_n3896_), .ZN(new_n3905_));
  NOR3_X1    g03638(.A1(new_n3902_), .A2(new_n3905_), .A3(new_n3900_), .ZN(new_n3906_));
  OAI21_X1   g03639(.A1(new_n3899_), .A2(new_n3906_), .B(new_n3769_), .ZN(new_n3907_));
  INV_X1     g03640(.I(new_n3769_), .ZN(new_n3908_));
  OAI21_X1   g03641(.A1(new_n3902_), .A2(new_n3900_), .B(new_n3905_), .ZN(new_n3909_));
  NAND3_X1   g03642(.A1(new_n3775_), .A2(new_n3898_), .A3(new_n3773_), .ZN(new_n3910_));
  NAND3_X1   g03643(.A1(new_n3910_), .A2(new_n3909_), .A3(new_n3908_), .ZN(new_n3911_));
  NAND2_X1   g03644(.A1(new_n3911_), .A2(new_n3907_), .ZN(new_n3912_));
  OAI22_X1   g03645(.A1(new_n1055_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n1061_), .ZN(new_n3913_));
  OAI21_X1   g03646(.A1(new_n1109_), .A2(new_n1332_), .B(new_n3913_), .ZN(new_n3914_));
  AOI21_X1   g03647(.A1(new_n3914_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n3915_));
  XOR2_X1    g03648(.A1(new_n1299_), .A2(new_n3915_), .Z(new_n3916_));
  INV_X1     g03649(.I(new_n3916_), .ZN(new_n3917_));
  NAND2_X1   g03650(.A1(new_n3912_), .A2(new_n3917_), .ZN(new_n3918_));
  XOR2_X1    g03651(.A1(new_n3760_), .A2(new_n3918_), .Z(new_n3919_));
  NAND2_X1   g03652(.A1(new_n3919_), .A2(new_n3648_), .ZN(new_n3920_));
  AOI21_X1   g03653(.A1(new_n3637_), .A2(new_n3639_), .B(new_n3644_), .ZN(new_n3921_));
  NOR2_X1    g03654(.A1(new_n3447_), .A2(new_n3437_), .ZN(new_n3922_));
  AOI21_X1   g03655(.A1(new_n3437_), .A2(new_n3445_), .B(new_n3922_), .ZN(new_n3923_));
  XOR2_X1    g03656(.A1(new_n3439_), .A2(new_n3437_), .Z(new_n3924_));
  NOR2_X1    g03657(.A1(new_n3924_), .A2(new_n3444_), .ZN(new_n3925_));
  NOR3_X1    g03658(.A1(new_n3647_), .A2(new_n3646_), .A3(new_n3643_), .ZN(new_n3926_));
  OAI21_X1   g03659(.A1(new_n3926_), .A2(new_n3921_), .B(new_n3925_), .ZN(new_n3927_));
  AOI21_X1   g03660(.A1(new_n3927_), .A2(new_n3923_), .B(new_n3323_), .ZN(new_n3928_));
  XOR2_X1    g03661(.A1(new_n3928_), .A2(new_n3918_), .Z(new_n3929_));
  NAND2_X1   g03662(.A1(new_n3929_), .A2(new_n3921_), .ZN(new_n3930_));
  OAI22_X1   g03663(.A1(new_n970_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n820_), .ZN(new_n3931_));
  OAI21_X1   g03664(.A1(new_n1518_), .A2(new_n894_), .B(new_n3931_), .ZN(new_n3932_));
  AOI21_X1   g03665(.A1(new_n3932_), .A2(new_n827_), .B(new_n970_), .ZN(new_n3933_));
  XNOR2_X1   g03666(.A1(new_n1638_), .A2(new_n3933_), .ZN(new_n3934_));
  AOI21_X1   g03667(.A1(new_n3930_), .A2(new_n3920_), .B(new_n3934_), .ZN(new_n3935_));
  NAND2_X1   g03668(.A1(new_n3758_), .A2(new_n3935_), .ZN(new_n3936_));
  INV_X1     g03669(.I(new_n3754_), .ZN(new_n3937_));
  OAI21_X1   g03670(.A1(new_n3937_), .A2(new_n3755_), .B(new_n3655_), .ZN(new_n3938_));
  AOI22_X1   g03671(.A1(new_n3938_), .A2(new_n3461_), .B1(new_n3317_), .B2(new_n3312_), .ZN(new_n3939_));
  INV_X1     g03672(.I(new_n3935_), .ZN(new_n3940_));
  NAND2_X1   g03673(.A1(new_n3940_), .A2(new_n3939_), .ZN(new_n3941_));
  AOI21_X1   g03674(.A1(new_n3941_), .A2(new_n3936_), .B(new_n3753_), .ZN(new_n3942_));
  INV_X1     g03675(.I(new_n3753_), .ZN(new_n3943_));
  NOR2_X1    g03676(.A1(new_n3940_), .A2(new_n3939_), .ZN(new_n3944_));
  NOR2_X1    g03677(.A1(new_n3758_), .A2(new_n3935_), .ZN(new_n3945_));
  NOR3_X1    g03678(.A1(new_n3944_), .A2(new_n3945_), .A3(new_n3943_), .ZN(new_n3946_));
  NOR2_X1    g03679(.A1(new_n3942_), .A2(new_n3946_), .ZN(new_n3947_));
  OAI22_X1   g03680(.A1(new_n607_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n610_), .ZN(new_n3948_));
  OAI21_X1   g03681(.A1(new_n1803_), .A2(new_n684_), .B(new_n3948_), .ZN(new_n3949_));
  AOI21_X1   g03682(.A1(new_n3949_), .A2(new_n612_), .B(new_n607_), .ZN(new_n3950_));
  XOR2_X1    g03683(.A1(new_n2106_), .A2(new_n3950_), .Z(new_n3951_));
  NOR2_X1    g03684(.A1(new_n3947_), .A2(new_n3951_), .ZN(new_n3952_));
  INV_X1     g03685(.I(new_n3952_), .ZN(new_n3953_));
  NOR2_X1    g03686(.A1(new_n3752_), .A2(new_n3953_), .ZN(new_n3954_));
  INV_X1     g03687(.I(new_n3474_), .ZN(new_n3955_));
  INV_X1     g03688(.I(new_n3544_), .ZN(new_n3956_));
  OAI21_X1   g03689(.A1(new_n3675_), .A2(new_n3676_), .B(new_n3548_), .ZN(new_n3957_));
  NAND3_X1   g03690(.A1(new_n3669_), .A2(new_n3673_), .A3(new_n3549_), .ZN(new_n3958_));
  AOI21_X1   g03691(.A1(new_n3957_), .A2(new_n3958_), .B(new_n3956_), .ZN(new_n3959_));
  OAI21_X1   g03692(.A1(new_n3959_), .A2(new_n3955_), .B(new_n3482_), .ZN(new_n3960_));
  NOR2_X1    g03693(.A1(new_n3960_), .A2(new_n3952_), .ZN(new_n3961_));
  OAI21_X1   g03694(.A1(new_n3954_), .A2(new_n3961_), .B(new_n3750_), .ZN(new_n3962_));
  NAND2_X1   g03695(.A1(new_n3960_), .A2(new_n3952_), .ZN(new_n3963_));
  NAND2_X1   g03696(.A1(new_n3752_), .A2(new_n3953_), .ZN(new_n3964_));
  NAND3_X1   g03697(.A1(new_n3964_), .A2(new_n3963_), .A3(new_n3749_), .ZN(new_n3965_));
  NAND2_X1   g03698(.A1(new_n3962_), .A2(new_n3965_), .ZN(new_n3966_));
  OAI22_X1   g03699(.A1(new_n448_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n450_), .ZN(new_n3967_));
  OAI21_X1   g03700(.A1(new_n2281_), .A2(new_n496_), .B(new_n3967_), .ZN(new_n3968_));
  AOI21_X1   g03701(.A1(new_n3968_), .A2(new_n452_), .B(new_n448_), .ZN(new_n3969_));
  XNOR2_X1   g03702(.A1(new_n2647_), .A2(new_n3969_), .ZN(new_n3970_));
  INV_X1     g03703(.I(new_n3970_), .ZN(new_n3971_));
  NAND2_X1   g03704(.A1(new_n3966_), .A2(new_n3971_), .ZN(new_n3972_));
  NOR2_X1    g03705(.A1(new_n3743_), .A2(new_n3972_), .ZN(new_n3973_));
  XOR2_X1    g03706(.A1(new_n3482_), .A2(new_n3955_), .Z(new_n3974_));
  NAND2_X1   g03707(.A1(new_n3974_), .A2(new_n3478_), .ZN(new_n3975_));
  AOI21_X1   g03708(.A1(new_n3687_), .A2(new_n3741_), .B(new_n3975_), .ZN(new_n3976_));
  OAI21_X1   g03709(.A1(new_n3492_), .A2(new_n3976_), .B(new_n3304_), .ZN(new_n3977_));
  AOI21_X1   g03710(.A1(new_n3966_), .A2(new_n3971_), .B(new_n3977_), .ZN(new_n3978_));
  OAI21_X1   g03711(.A1(new_n3978_), .A2(new_n3973_), .B(new_n3741_), .ZN(new_n3979_));
  OR3_X2     g03712(.A1(new_n3978_), .A2(new_n3741_), .A3(new_n3973_), .Z(new_n3980_));
  NAND2_X1   g03713(.A1(new_n3980_), .A2(new_n3979_), .ZN(new_n3981_));
  OAI22_X1   g03714(.A1(new_n3018_), .A2(new_n341_), .B1(new_n404_), .B2(new_n3260_), .ZN(new_n3982_));
  OAI21_X1   g03715(.A1(new_n2842_), .A2(new_n366_), .B(new_n3982_), .ZN(new_n3983_));
  AOI21_X1   g03716(.A1(new_n3983_), .A2(new_n334_), .B(new_n341_), .ZN(new_n3984_));
  XNOR2_X1   g03717(.A1(new_n3264_), .A2(new_n3984_), .ZN(new_n3985_));
  OR2_X2     g03718(.A1(new_n3981_), .A2(new_n3985_), .Z(new_n3986_));
  NAND2_X1   g03719(.A1(new_n3981_), .A2(new_n3985_), .ZN(new_n3987_));
  NAND2_X1   g03720(.A1(new_n3986_), .A2(new_n3987_), .ZN(new_n3988_));
  INV_X1     g03721(.I(\b[33] ), .ZN(new_n3989_));
  NOR2_X1    g03722(.A1(new_n3989_), .A2(\b[31] ), .ZN(new_n3990_));
  NOR2_X1    g03723(.A1(new_n3709_), .A2(\b[33] ), .ZN(new_n3991_));
  OAI21_X1   g03724(.A1(new_n3990_), .A2(new_n3991_), .B(new_n3716_), .ZN(new_n3992_));
  XOR2_X1    g03725(.A1(new_n3713_), .A2(new_n3992_), .Z(new_n3993_));
  NAND2_X1   g03726(.A1(new_n286_), .A2(\b[32] ), .ZN(new_n3994_));
  AOI22_X1   g03727(.A1(new_n304_), .A2(\b[31] ), .B1(new_n262_), .B2(\b[33] ), .ZN(new_n3995_));
  AOI21_X1   g03728(.A1(new_n3994_), .A2(new_n3995_), .B(new_n426_), .ZN(new_n3996_));
  NAND2_X1   g03729(.A1(new_n3993_), .A2(new_n3996_), .ZN(new_n3997_));
  XOR2_X1    g03730(.A1(new_n3997_), .A2(\a[2] ), .Z(new_n3998_));
  NOR2_X1    g03731(.A1(new_n3988_), .A2(new_n3998_), .ZN(new_n3999_));
  INV_X1     g03732(.I(new_n3998_), .ZN(new_n4000_));
  AOI21_X1   g03733(.A1(new_n3986_), .A2(new_n3987_), .B(new_n4000_), .ZN(new_n4001_));
  OAI21_X1   g03734(.A1(new_n3999_), .A2(new_n4001_), .B(new_n3739_), .ZN(new_n4002_));
  AOI21_X1   g03735(.A1(new_n3986_), .A2(new_n3987_), .B(new_n3998_), .ZN(new_n4003_));
  NOR2_X1    g03736(.A1(new_n3988_), .A2(new_n4000_), .ZN(new_n4004_));
  OAI21_X1   g03737(.A1(new_n4004_), .A2(new_n4003_), .B(new_n3738_), .ZN(new_n4005_));
  AOI21_X1   g03738(.A1(new_n4002_), .A2(new_n4005_), .B(new_n3728_), .ZN(new_n4006_));
  XOR2_X1    g03739(.A1(new_n4006_), .A2(new_n3730_), .Z(new_n4007_));
  XOR2_X1    g03740(.A1(new_n4007_), .A2(new_n3533_), .Z(\f[33] ));
  XNOR2_X1   g03741(.A1(new_n3988_), .A2(new_n3738_), .ZN(new_n4009_));
  NAND2_X1   g03742(.A1(new_n4009_), .A2(new_n3998_), .ZN(new_n4010_));
  NAND2_X1   g03743(.A1(new_n4002_), .A2(new_n4005_), .ZN(new_n4011_));
  AOI21_X1   g03744(.A1(new_n4011_), .A2(new_n3727_), .B(new_n3729_), .ZN(new_n4012_));
  INV_X1     g03745(.I(new_n4012_), .ZN(new_n4013_));
  NOR2_X1    g03746(.A1(new_n4011_), .A2(new_n3727_), .ZN(new_n4014_));
  NOR2_X1    g03747(.A1(new_n3533_), .A2(new_n4014_), .ZN(new_n4015_));
  NAND2_X1   g03748(.A1(new_n4015_), .A2(new_n4013_), .ZN(new_n4016_));
  NAND2_X1   g03749(.A1(new_n3739_), .A2(new_n3987_), .ZN(new_n4017_));
  NAND2_X1   g03750(.A1(new_n4017_), .A2(new_n3986_), .ZN(new_n4018_));
  OR2_X2     g03751(.A1(new_n3942_), .A2(new_n3946_), .Z(new_n4019_));
  NAND2_X1   g03752(.A1(new_n4019_), .A2(new_n3749_), .ZN(new_n4020_));
  INV_X1     g03753(.I(new_n3951_), .ZN(new_n4021_));
  OAI21_X1   g03754(.A1(new_n4019_), .A2(new_n3749_), .B(new_n4021_), .ZN(new_n4022_));
  OAI21_X1   g03755(.A1(new_n3960_), .A2(new_n4022_), .B(new_n4020_), .ZN(new_n4023_));
  NAND2_X1   g03756(.A1(new_n3930_), .A2(new_n3920_), .ZN(new_n4024_));
  NAND2_X1   g03757(.A1(new_n4024_), .A2(new_n3753_), .ZN(new_n4025_));
  INV_X1     g03758(.I(new_n3934_), .ZN(new_n4026_));
  OAI21_X1   g03759(.A1(new_n4024_), .A2(new_n3753_), .B(new_n4026_), .ZN(new_n4027_));
  OAI21_X1   g03760(.A1(new_n4027_), .A2(new_n3758_), .B(new_n4025_), .ZN(new_n4028_));
  AOI21_X1   g03761(.A1(new_n3910_), .A2(new_n3909_), .B(new_n3908_), .ZN(new_n4029_));
  NOR3_X1    g03762(.A1(new_n3899_), .A2(new_n3906_), .A3(new_n3769_), .ZN(new_n4030_));
  NOR2_X1    g03763(.A1(new_n4029_), .A2(new_n4030_), .ZN(new_n4031_));
  NOR2_X1    g03764(.A1(new_n4031_), .A2(new_n3648_), .ZN(new_n4032_));
  AOI21_X1   g03765(.A1(new_n4031_), .A2(new_n3648_), .B(new_n3916_), .ZN(new_n4033_));
  AOI21_X1   g03766(.A1(new_n3928_), .A2(new_n4033_), .B(new_n4032_), .ZN(new_n4034_));
  NAND3_X1   g03767(.A1(new_n3881_), .A2(new_n3327_), .A3(new_n3781_), .ZN(new_n4035_));
  NOR2_X1    g03768(.A1(new_n3883_), .A2(new_n3882_), .ZN(new_n4036_));
  NAND3_X1   g03769(.A1(new_n3866_), .A2(new_n3871_), .A3(new_n3888_), .ZN(new_n4037_));
  NAND2_X1   g03770(.A1(new_n4037_), .A2(new_n3884_), .ZN(new_n4038_));
  OAI22_X1   g03771(.A1(new_n4035_), .A2(new_n4038_), .B1(new_n3888_), .B2(new_n4036_), .ZN(new_n4039_));
  NOR2_X1    g03772(.A1(new_n3848_), .A2(new_n3854_), .ZN(new_n4040_));
  NOR2_X1    g03773(.A1(new_n3789_), .A2(new_n4040_), .ZN(new_n4041_));
  NOR3_X1    g03774(.A1(new_n3788_), .A2(new_n3848_), .A3(new_n3854_), .ZN(new_n4042_));
  NOR4_X1    g03775(.A1(new_n4042_), .A2(new_n3790_), .A3(new_n3791_), .A4(new_n3858_), .ZN(new_n4043_));
  NAND2_X1   g03776(.A1(new_n3804_), .A2(new_n3802_), .ZN(new_n4044_));
  INV_X1     g03777(.I(new_n4044_), .ZN(new_n4045_));
  NOR2_X1    g03778(.A1(new_n3804_), .A2(new_n3802_), .ZN(new_n4046_));
  OAI21_X1   g03779(.A1(new_n4045_), .A2(new_n4046_), .B(new_n3794_), .ZN(new_n4047_));
  NAND2_X1   g03780(.A1(new_n3814_), .A2(new_n3819_), .ZN(new_n4048_));
  NAND3_X1   g03781(.A1(new_n4048_), .A2(new_n4044_), .A3(new_n3824_), .ZN(new_n4049_));
  AOI21_X1   g03782(.A1(new_n4047_), .A2(new_n4049_), .B(new_n3815_), .ZN(new_n4050_));
  AOI21_X1   g03783(.A1(new_n3828_), .A2(new_n4050_), .B(new_n3829_), .ZN(new_n4051_));
  NOR2_X1    g03784(.A1(new_n3574_), .A2(new_n3819_), .ZN(new_n4052_));
  NAND4_X1   g03785(.A1(new_n3361_), .A2(new_n3362_), .A3(new_n3373_), .A4(new_n3824_), .ZN(new_n4053_));
  AOI21_X1   g03786(.A1(new_n3574_), .A2(new_n3819_), .B(new_n4053_), .ZN(new_n4054_));
  NOR2_X1    g03787(.A1(new_n4054_), .A2(new_n4052_), .ZN(new_n4055_));
  OAI22_X1   g03788(.A1(new_n325_), .A2(new_n3352_), .B1(new_n3357_), .B2(new_n298_), .ZN(new_n4056_));
  OAI21_X1   g03789(.A1(new_n280_), .A2(new_n3569_), .B(new_n4056_), .ZN(new_n4057_));
  AOI21_X1   g03790(.A1(new_n4057_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n4058_));
  XOR2_X1    g03791(.A1(new_n4058_), .A2(new_n329_), .Z(new_n4059_));
  XNOR2_X1   g03792(.A1(\a[33] ), .A2(\a[35] ), .ZN(new_n4060_));
  XNOR2_X1   g03793(.A1(\a[32] ), .A2(\a[34] ), .ZN(new_n4061_));
  NOR2_X1    g03794(.A1(new_n4061_), .A2(new_n4060_), .ZN(new_n4062_));
  INV_X1     g03795(.I(\a[34] ), .ZN(new_n4063_));
  NOR3_X1    g03796(.A1(new_n4063_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n4064_));
  NAND3_X1   g03797(.A1(new_n4063_), .A2(\a[32] ), .A3(\a[33] ), .ZN(new_n4065_));
  INV_X1     g03798(.I(new_n4065_), .ZN(new_n4066_));
  NOR2_X1    g03799(.A1(new_n4066_), .A2(new_n4064_), .ZN(new_n4067_));
  NOR2_X1    g03800(.A1(new_n4067_), .A2(new_n269_), .ZN(new_n4068_));
  INV_X1     g03801(.I(\a[35] ), .ZN(new_n4069_));
  XOR2_X1    g03802(.A1(\a[33] ), .A2(\a[35] ), .Z(new_n4070_));
  XOR2_X1    g03803(.A1(\a[32] ), .A2(\a[34] ), .Z(new_n4071_));
  NAND2_X1   g03804(.A1(new_n4071_), .A2(new_n4070_), .ZN(new_n4072_));
  OAI21_X1   g03805(.A1(new_n4072_), .A2(new_n258_), .B(new_n4069_), .ZN(new_n4073_));
  OAI21_X1   g03806(.A1(new_n4073_), .A2(new_n4068_), .B(new_n4062_), .ZN(new_n4074_));
  NOR2_X1    g03807(.A1(new_n4074_), .A2(new_n271_), .ZN(new_n4075_));
  NAND2_X1   g03808(.A1(new_n4074_), .A2(new_n271_), .ZN(new_n4076_));
  INV_X1     g03809(.I(new_n4076_), .ZN(new_n4077_));
  NAND2_X1   g03810(.A1(new_n3794_), .A2(\a[35] ), .ZN(new_n4078_));
  INV_X1     g03811(.I(new_n4078_), .ZN(new_n4079_));
  NOR3_X1    g03812(.A1(new_n4077_), .A2(new_n4075_), .A3(new_n4079_), .ZN(new_n4080_));
  INV_X1     g03813(.I(new_n4075_), .ZN(new_n4081_));
  AOI21_X1   g03814(.A1(new_n4081_), .A2(new_n4076_), .B(new_n4078_), .ZN(new_n4082_));
  OR2_X2     g03815(.A1(new_n4082_), .A2(new_n4080_), .Z(new_n4083_));
  NAND2_X1   g03816(.A1(new_n4083_), .A2(new_n4059_), .ZN(new_n4084_));
  XOR2_X1    g03817(.A1(new_n4058_), .A2(new_n807_), .Z(new_n4085_));
  NOR2_X1    g03818(.A1(new_n4082_), .A2(new_n4080_), .ZN(new_n4086_));
  NAND2_X1   g03819(.A1(new_n4085_), .A2(new_n4086_), .ZN(new_n4087_));
  AOI21_X1   g03820(.A1(new_n4084_), .A2(new_n4087_), .B(new_n4055_), .ZN(new_n4088_));
  NOR2_X1    g03821(.A1(new_n4059_), .A2(new_n4086_), .ZN(new_n4089_));
  NOR2_X1    g03822(.A1(new_n4083_), .A2(new_n4085_), .ZN(new_n4090_));
  OAI21_X1   g03823(.A1(new_n4089_), .A2(new_n4090_), .B(new_n4055_), .ZN(new_n4091_));
  INV_X1     g03824(.I(new_n4091_), .ZN(new_n4092_));
  NOR2_X1    g03825(.A1(new_n4092_), .A2(new_n4088_), .ZN(new_n4093_));
  INV_X1     g03826(.I(new_n2884_), .ZN(new_n4094_));
  AOI22_X1   g03827(.A1(new_n2694_), .A2(\b[6] ), .B1(\b[7] ), .B2(new_n2699_), .ZN(new_n4095_));
  AOI21_X1   g03828(.A1(\b[5] ), .A2(new_n4094_), .B(new_n4095_), .ZN(new_n4096_));
  OAI21_X1   g03829(.A1(new_n4096_), .A2(\a[29] ), .B(new_n2694_), .ZN(new_n4097_));
  XNOR2_X1   g03830(.A1(new_n471_), .A2(new_n4097_), .ZN(new_n4098_));
  NOR2_X1    g03831(.A1(new_n4093_), .A2(new_n4098_), .ZN(new_n4099_));
  INV_X1     g03832(.I(new_n4055_), .ZN(new_n4100_));
  NAND2_X1   g03833(.A1(new_n4084_), .A2(new_n4087_), .ZN(new_n4101_));
  NAND2_X1   g03834(.A1(new_n4101_), .A2(new_n4100_), .ZN(new_n4102_));
  NAND2_X1   g03835(.A1(new_n4102_), .A2(new_n4091_), .ZN(new_n4103_));
  INV_X1     g03836(.I(new_n4098_), .ZN(new_n4104_));
  NOR2_X1    g03837(.A1(new_n4103_), .A2(new_n4104_), .ZN(new_n4105_));
  NOR2_X1    g03838(.A1(new_n4099_), .A2(new_n4105_), .ZN(new_n4106_));
  NOR3_X1    g03839(.A1(new_n4051_), .A2(new_n4106_), .A3(new_n3847_), .ZN(new_n4107_));
  AOI21_X1   g03840(.A1(new_n3826_), .A2(new_n3825_), .B(new_n3824_), .ZN(new_n4108_));
  NOR3_X1    g03841(.A1(new_n3817_), .A2(new_n3822_), .A3(new_n3794_), .ZN(new_n4109_));
  OAI21_X1   g03842(.A1(new_n4108_), .A2(new_n4109_), .B(new_n4050_), .ZN(new_n4110_));
  NAND2_X1   g03843(.A1(new_n4110_), .A2(new_n3830_), .ZN(new_n4111_));
  NAND3_X1   g03844(.A1(new_n4102_), .A2(new_n4091_), .A3(new_n4104_), .ZN(new_n4112_));
  OAI21_X1   g03845(.A1(new_n4092_), .A2(new_n4088_), .B(new_n4098_), .ZN(new_n4113_));
  NAND2_X1   g03846(.A1(new_n4113_), .A2(new_n4112_), .ZN(new_n4114_));
  INV_X1     g03847(.I(new_n4114_), .ZN(new_n4115_));
  AOI21_X1   g03848(.A1(new_n4111_), .A2(new_n3853_), .B(new_n4115_), .ZN(new_n4116_));
  NOR2_X1    g03849(.A1(new_n4116_), .A2(new_n4107_), .ZN(new_n4117_));
  OAI22_X1   g03850(.A1(new_n2171_), .A2(new_n565_), .B1(new_n656_), .B2(new_n2166_), .ZN(new_n4118_));
  OAI21_X1   g03851(.A1(new_n515_), .A2(new_n2322_), .B(new_n4118_), .ZN(new_n4119_));
  AOI21_X1   g03852(.A1(new_n4119_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n4120_));
  XNOR2_X1   g03853(.A1(new_n660_), .A2(new_n4120_), .ZN(new_n4121_));
  NOR2_X1    g03854(.A1(new_n4117_), .A2(new_n4121_), .ZN(new_n4122_));
  INV_X1     g03855(.I(new_n4106_), .ZN(new_n4123_));
  NAND3_X1   g03856(.A1(new_n4123_), .A2(new_n4111_), .A3(new_n3853_), .ZN(new_n4124_));
  OAI21_X1   g03857(.A1(new_n4051_), .A2(new_n3847_), .B(new_n4114_), .ZN(new_n4125_));
  NAND2_X1   g03858(.A1(new_n4124_), .A2(new_n4125_), .ZN(new_n4126_));
  INV_X1     g03859(.I(new_n4121_), .ZN(new_n4127_));
  NOR2_X1    g03860(.A1(new_n4126_), .A2(new_n4127_), .ZN(new_n4128_));
  OAI22_X1   g03861(.A1(new_n4043_), .A2(new_n4041_), .B1(new_n4128_), .B2(new_n4122_), .ZN(new_n4129_));
  NOR2_X1    g03862(.A1(new_n4043_), .A2(new_n4041_), .ZN(new_n4130_));
  NAND3_X1   g03863(.A1(new_n4124_), .A2(new_n4125_), .A3(new_n4127_), .ZN(new_n4131_));
  OAI21_X1   g03864(.A1(new_n4116_), .A2(new_n4107_), .B(new_n4121_), .ZN(new_n4132_));
  NAND2_X1   g03865(.A1(new_n4131_), .A2(new_n4132_), .ZN(new_n4133_));
  NAND2_X1   g03866(.A1(new_n4130_), .A2(new_n4133_), .ZN(new_n4134_));
  OAI22_X1   g03867(.A1(new_n1712_), .A2(new_n780_), .B1(new_n861_), .B2(new_n1707_), .ZN(new_n4135_));
  OAI21_X1   g03868(.A1(new_n706_), .A2(new_n1850_), .B(new_n4135_), .ZN(new_n4136_));
  AOI21_X1   g03869(.A1(new_n4136_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n4137_));
  XNOR2_X1   g03870(.A1(new_n860_), .A2(new_n4137_), .ZN(new_n4138_));
  INV_X1     g03871(.I(new_n4138_), .ZN(new_n4139_));
  NAND3_X1   g03872(.A1(new_n4134_), .A2(new_n4129_), .A3(new_n4139_), .ZN(new_n4140_));
  AOI21_X1   g03873(.A1(new_n4134_), .A2(new_n4129_), .B(new_n4139_), .ZN(new_n4141_));
  INV_X1     g03874(.I(new_n4141_), .ZN(new_n4142_));
  NAND2_X1   g03875(.A1(new_n4142_), .A2(new_n4140_), .ZN(new_n4143_));
  NAND2_X1   g03876(.A1(new_n4039_), .A2(new_n4143_), .ZN(new_n4144_));
  NOR2_X1    g03877(.A1(new_n4036_), .A2(new_n3888_), .ZN(new_n4145_));
  AOI21_X1   g03878(.A1(new_n4036_), .A2(new_n3888_), .B(new_n3875_), .ZN(new_n4146_));
  AOI21_X1   g03879(.A1(new_n3889_), .A2(new_n4146_), .B(new_n4145_), .ZN(new_n4147_));
  INV_X1     g03880(.I(new_n4129_), .ZN(new_n4148_));
  INV_X1     g03881(.I(new_n4133_), .ZN(new_n4149_));
  NOR3_X1    g03882(.A1(new_n4149_), .A2(new_n4041_), .A3(new_n4043_), .ZN(new_n4150_));
  OAI21_X1   g03883(.A1(new_n4148_), .A2(new_n4150_), .B(new_n4139_), .ZN(new_n4151_));
  NAND3_X1   g03884(.A1(new_n4134_), .A2(new_n4129_), .A3(new_n4138_), .ZN(new_n4152_));
  NAND2_X1   g03885(.A1(new_n4151_), .A2(new_n4152_), .ZN(new_n4153_));
  NAND2_X1   g03886(.A1(new_n4147_), .A2(new_n4153_), .ZN(new_n4154_));
  NAND2_X1   g03887(.A1(new_n4144_), .A2(new_n4154_), .ZN(new_n4155_));
  OAI22_X1   g03888(.A1(new_n1347_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n1344_), .ZN(new_n4156_));
  OAI21_X1   g03889(.A1(new_n930_), .A2(new_n1457_), .B(new_n4156_), .ZN(new_n4157_));
  AOI21_X1   g03890(.A1(new_n4157_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n4158_));
  XOR2_X1    g03891(.A1(new_n1114_), .A2(new_n4158_), .Z(new_n4159_));
  INV_X1     g03892(.I(new_n4159_), .ZN(new_n4160_));
  NAND2_X1   g03893(.A1(new_n4155_), .A2(new_n4160_), .ZN(new_n4161_));
  INV_X1     g03894(.I(new_n4140_), .ZN(new_n4162_));
  NOR2_X1    g03895(.A1(new_n4162_), .A2(new_n4141_), .ZN(new_n4163_));
  NOR2_X1    g03896(.A1(new_n4163_), .A2(new_n4147_), .ZN(new_n4164_));
  INV_X1     g03897(.I(new_n4153_), .ZN(new_n4165_));
  NOR2_X1    g03898(.A1(new_n4165_), .A2(new_n4039_), .ZN(new_n4166_));
  NOR2_X1    g03899(.A1(new_n4166_), .A2(new_n4164_), .ZN(new_n4167_));
  NAND2_X1   g03900(.A1(new_n4167_), .A2(new_n4159_), .ZN(new_n4168_));
  NAND2_X1   g03901(.A1(new_n4168_), .A2(new_n4161_), .ZN(new_n4169_));
  INV_X1     g03902(.I(new_n4169_), .ZN(new_n4170_));
  NAND3_X1   g03903(.A1(new_n3773_), .A2(new_n3439_), .A3(new_n3901_), .ZN(new_n4171_));
  OAI21_X1   g03904(.A1(new_n3887_), .A2(new_n3892_), .B(new_n3908_), .ZN(new_n4172_));
  NAND3_X1   g03905(.A1(new_n3903_), .A2(new_n3904_), .A3(new_n3769_), .ZN(new_n4173_));
  NAND2_X1   g03906(.A1(new_n4173_), .A2(new_n3897_), .ZN(new_n4174_));
  OAI21_X1   g03907(.A1(new_n4171_), .A2(new_n4174_), .B(new_n4172_), .ZN(new_n4175_));
  OAI22_X1   g03908(.A1(new_n1055_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n1061_), .ZN(new_n4176_));
  OAI21_X1   g03909(.A1(new_n1189_), .A2(new_n1332_), .B(new_n4176_), .ZN(new_n4177_));
  AOI21_X1   g03910(.A1(new_n4177_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n4178_));
  XNOR2_X1   g03911(.A1(new_n1421_), .A2(new_n4178_), .ZN(new_n4179_));
  INV_X1     g03912(.I(new_n4179_), .ZN(new_n4180_));
  NAND2_X1   g03913(.A1(new_n4175_), .A2(new_n4180_), .ZN(new_n4181_));
  NOR2_X1    g03914(.A1(new_n3902_), .A2(new_n3900_), .ZN(new_n4182_));
  NOR2_X1    g03915(.A1(new_n3892_), .A2(new_n3887_), .ZN(new_n4183_));
  INV_X1     g03916(.I(new_n4183_), .ZN(new_n4184_));
  AOI21_X1   g03917(.A1(new_n4183_), .A2(new_n3769_), .B(new_n3896_), .ZN(new_n4185_));
  AOI22_X1   g03918(.A1(new_n4182_), .A2(new_n4185_), .B1(new_n3908_), .B2(new_n4184_), .ZN(new_n4186_));
  NAND2_X1   g03919(.A1(new_n4186_), .A2(new_n4179_), .ZN(new_n4187_));
  AOI21_X1   g03920(.A1(new_n4187_), .A2(new_n4181_), .B(new_n4170_), .ZN(new_n4188_));
  NAND2_X1   g03921(.A1(new_n4186_), .A2(new_n4180_), .ZN(new_n4189_));
  NAND2_X1   g03922(.A1(new_n4175_), .A2(new_n4179_), .ZN(new_n4190_));
  AOI21_X1   g03923(.A1(new_n4189_), .A2(new_n4190_), .B(new_n4169_), .ZN(new_n4191_));
  NOR2_X1    g03924(.A1(new_n4188_), .A2(new_n4191_), .ZN(new_n4192_));
  OAI22_X1   g03925(.A1(new_n970_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n820_), .ZN(new_n4193_));
  OAI21_X1   g03926(.A1(new_n1525_), .A2(new_n894_), .B(new_n4193_), .ZN(new_n4194_));
  AOI21_X1   g03927(.A1(new_n4194_), .A2(new_n827_), .B(new_n970_), .ZN(new_n4195_));
  XOR2_X1    g03928(.A1(new_n1808_), .A2(new_n4195_), .Z(new_n4196_));
  XOR2_X1    g03929(.A1(new_n4192_), .A2(new_n4196_), .Z(new_n4197_));
  NOR2_X1    g03930(.A1(new_n4197_), .A2(new_n4034_), .ZN(new_n4198_));
  NAND2_X1   g03931(.A1(new_n3912_), .A2(new_n3921_), .ZN(new_n4199_));
  OAI21_X1   g03932(.A1(new_n3912_), .A2(new_n3921_), .B(new_n3917_), .ZN(new_n4200_));
  OAI21_X1   g03933(.A1(new_n3760_), .A2(new_n4200_), .B(new_n4199_), .ZN(new_n4201_));
  INV_X1     g03934(.I(new_n4196_), .ZN(new_n4202_));
  XOR2_X1    g03935(.A1(new_n4192_), .A2(new_n4202_), .Z(new_n4203_));
  NOR2_X1    g03936(.A1(new_n4203_), .A2(new_n4201_), .ZN(new_n4204_));
  NOR2_X1    g03937(.A1(new_n4198_), .A2(new_n4204_), .ZN(new_n4205_));
  XOR2_X1    g03938(.A1(new_n4028_), .A2(new_n4205_), .Z(new_n4206_));
  OAI22_X1   g03939(.A1(new_n607_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n610_), .ZN(new_n4207_));
  OAI21_X1   g03940(.A1(new_n1936_), .A2(new_n684_), .B(new_n4207_), .ZN(new_n4208_));
  AOI21_X1   g03941(.A1(new_n4208_), .A2(new_n612_), .B(new_n607_), .ZN(new_n4209_));
  XNOR2_X1   g03942(.A1(new_n2280_), .A2(new_n4209_), .ZN(new_n4210_));
  INV_X1     g03943(.I(new_n4210_), .ZN(new_n4211_));
  NAND2_X1   g03944(.A1(new_n4206_), .A2(new_n4211_), .ZN(new_n4212_));
  NOR2_X1    g03945(.A1(new_n4206_), .A2(new_n4211_), .ZN(new_n4213_));
  INV_X1     g03946(.I(new_n4213_), .ZN(new_n4214_));
  NAND2_X1   g03947(.A1(new_n4214_), .A2(new_n4212_), .ZN(new_n4215_));
  NAND2_X1   g03948(.A1(new_n4215_), .A2(new_n4023_), .ZN(new_n4216_));
  XOR2_X1    g03949(.A1(new_n4206_), .A2(new_n4210_), .Z(new_n4217_));
  OAI21_X1   g03950(.A1(new_n4023_), .A2(new_n4217_), .B(new_n4216_), .ZN(new_n4218_));
  INV_X1     g03951(.I(new_n4218_), .ZN(new_n4219_));
  OAI22_X1   g03952(.A1(new_n448_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n450_), .ZN(new_n4220_));
  OAI21_X1   g03953(.A1(new_n2439_), .A2(new_n496_), .B(new_n4220_), .ZN(new_n4221_));
  AOI21_X1   g03954(.A1(new_n4221_), .A2(new_n452_), .B(new_n448_), .ZN(new_n4222_));
  XNOR2_X1   g03955(.A1(new_n2846_), .A2(new_n4222_), .ZN(new_n4223_));
  NOR2_X1    g03956(.A1(new_n4219_), .A2(new_n4223_), .ZN(new_n4224_));
  INV_X1     g03957(.I(new_n4224_), .ZN(new_n4225_));
  NAND2_X1   g03958(.A1(new_n4219_), .A2(new_n4223_), .ZN(new_n4226_));
  NAND2_X1   g03959(.A1(new_n4225_), .A2(new_n4226_), .ZN(new_n4227_));
  AOI21_X1   g03960(.A1(new_n3962_), .A2(new_n3965_), .B(new_n3741_), .ZN(new_n4228_));
  INV_X1     g03961(.I(new_n4228_), .ZN(new_n4229_));
  OAI21_X1   g03962(.A1(new_n3966_), .A2(new_n3689_), .B(new_n3971_), .ZN(new_n4230_));
  OAI21_X1   g03963(.A1(new_n3977_), .A2(new_n4230_), .B(new_n4229_), .ZN(new_n4231_));
  XOR2_X1    g03964(.A1(new_n4227_), .A2(new_n4231_), .Z(new_n4232_));
  OAI22_X1   g03965(.A1(new_n3260_), .A2(new_n341_), .B1(new_n404_), .B2(new_n3709_), .ZN(new_n4233_));
  OAI21_X1   g03966(.A1(new_n3018_), .A2(new_n366_), .B(new_n4233_), .ZN(new_n4234_));
  AOI21_X1   g03967(.A1(new_n4234_), .A2(new_n334_), .B(new_n341_), .ZN(new_n4235_));
  XNOR2_X1   g03968(.A1(new_n3514_), .A2(new_n4235_), .ZN(new_n4236_));
  NOR2_X1    g03969(.A1(new_n4232_), .A2(new_n4236_), .ZN(new_n4237_));
  NAND2_X1   g03970(.A1(new_n4232_), .A2(new_n4236_), .ZN(new_n4238_));
  INV_X1     g03971(.I(new_n4238_), .ZN(new_n4239_));
  NOR2_X1    g03972(.A1(new_n4239_), .A2(new_n4237_), .ZN(new_n4240_));
  INV_X1     g03973(.I(new_n4240_), .ZN(new_n4241_));
  INV_X1     g03974(.I(new_n4236_), .ZN(new_n4242_));
  XOR2_X1    g03975(.A1(new_n4232_), .A2(new_n4242_), .Z(new_n4243_));
  NOR2_X1    g03976(.A1(new_n4018_), .A2(new_n4243_), .ZN(new_n4244_));
  AOI21_X1   g03977(.A1(new_n4018_), .A2(new_n4241_), .B(new_n4244_), .ZN(new_n4245_));
  NOR2_X1    g03978(.A1(\b[32] ), .A2(\b[33] ), .ZN(new_n4246_));
  AOI21_X1   g03979(.A1(new_n3713_), .A2(new_n4246_), .B(new_n3709_), .ZN(new_n4247_));
  NOR2_X1    g03980(.A1(new_n3717_), .A2(new_n3989_), .ZN(new_n4248_));
  INV_X1     g03981(.I(new_n4248_), .ZN(new_n4249_));
  NOR2_X1    g03982(.A1(new_n3713_), .A2(new_n4249_), .ZN(new_n4250_));
  NOR2_X1    g03983(.A1(new_n4247_), .A2(new_n4250_), .ZN(new_n4251_));
  XNOR2_X1   g03984(.A1(\b[33] ), .A2(\b[34] ), .ZN(new_n4252_));
  INV_X1     g03985(.I(\b[34] ), .ZN(new_n4253_));
  NOR2_X1    g03986(.A1(new_n3989_), .A2(new_n4253_), .ZN(new_n4254_));
  NOR2_X1    g03987(.A1(\b[33] ), .A2(\b[34] ), .ZN(new_n4255_));
  OAI21_X1   g03988(.A1(new_n4254_), .A2(new_n4255_), .B(new_n4251_), .ZN(new_n4256_));
  OAI21_X1   g03989(.A1(new_n4251_), .A2(new_n4252_), .B(new_n4256_), .ZN(new_n4257_));
  OAI22_X1   g03990(.A1(new_n330_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n263_), .ZN(new_n4258_));
  OAI21_X1   g03991(.A1(new_n3717_), .A2(new_n289_), .B(new_n4258_), .ZN(new_n4259_));
  AOI21_X1   g03992(.A1(new_n4259_), .A2(new_n260_), .B(new_n426_), .ZN(new_n4260_));
  XNOR2_X1   g03993(.A1(new_n4257_), .A2(new_n4260_), .ZN(new_n4261_));
  NOR2_X1    g03994(.A1(new_n4245_), .A2(new_n4261_), .ZN(new_n4262_));
  XOR2_X1    g03995(.A1(new_n4016_), .A2(new_n4262_), .Z(new_n4263_));
  XOR2_X1    g03996(.A1(new_n4263_), .A2(new_n4010_), .Z(\f[34] ));
  NOR2_X1    g03997(.A1(new_n4016_), .A2(new_n4245_), .ZN(new_n4265_));
  NOR2_X1    g03998(.A1(new_n4010_), .A2(new_n4261_), .ZN(new_n4266_));
  INV_X1     g03999(.I(new_n4266_), .ZN(new_n4267_));
  AOI21_X1   g04000(.A1(new_n4016_), .A2(new_n4245_), .B(new_n4267_), .ZN(new_n4268_));
  NOR2_X1    g04001(.A1(new_n4268_), .A2(new_n4265_), .ZN(new_n4269_));
  AOI21_X1   g04002(.A1(new_n3964_), .A2(new_n3963_), .B(new_n3749_), .ZN(new_n4270_));
  NOR3_X1    g04003(.A1(new_n3954_), .A2(new_n3961_), .A3(new_n3750_), .ZN(new_n4271_));
  NOR3_X1    g04004(.A1(new_n4271_), .A2(new_n4270_), .A3(new_n3689_), .ZN(new_n4272_));
  NOR2_X1    g04005(.A1(new_n4272_), .A2(new_n3970_), .ZN(new_n4273_));
  AOI21_X1   g04006(.A1(new_n3743_), .A2(new_n4273_), .B(new_n4228_), .ZN(new_n4274_));
  NAND2_X1   g04007(.A1(new_n4274_), .A2(new_n4242_), .ZN(new_n4275_));
  NAND2_X1   g04008(.A1(new_n4231_), .A2(new_n4236_), .ZN(new_n4276_));
  AOI22_X1   g04009(.A1(new_n4276_), .A2(new_n4275_), .B1(new_n4225_), .B2(new_n4226_), .ZN(new_n4277_));
  NAND2_X1   g04010(.A1(new_n4231_), .A2(new_n4242_), .ZN(new_n4278_));
  NAND2_X1   g04011(.A1(new_n4274_), .A2(new_n4236_), .ZN(new_n4279_));
  AOI21_X1   g04012(.A1(new_n4278_), .A2(new_n4279_), .B(new_n4227_), .ZN(new_n4280_));
  OAI21_X1   g04013(.A1(new_n4277_), .A2(new_n4280_), .B(new_n3981_), .ZN(new_n4281_));
  NAND2_X1   g04014(.A1(new_n4281_), .A2(new_n3985_), .ZN(new_n4282_));
  NOR3_X1    g04015(.A1(new_n3981_), .A2(new_n4277_), .A3(new_n4280_), .ZN(new_n4283_));
  NOR2_X1    g04016(.A1(new_n3738_), .A2(new_n4283_), .ZN(new_n4284_));
  NAND2_X1   g04017(.A1(new_n4284_), .A2(new_n4282_), .ZN(new_n4285_));
  INV_X1     g04018(.I(new_n4212_), .ZN(new_n4286_));
  AOI21_X1   g04019(.A1(new_n4023_), .A2(new_n4214_), .B(new_n4286_), .ZN(new_n4287_));
  NOR2_X1    g04020(.A1(new_n3929_), .A2(new_n3921_), .ZN(new_n4288_));
  NOR2_X1    g04021(.A1(new_n3919_), .A2(new_n3648_), .ZN(new_n4289_));
  NOR3_X1    g04022(.A1(new_n4288_), .A2(new_n4289_), .A3(new_n3753_), .ZN(new_n4290_));
  NOR2_X1    g04023(.A1(new_n4290_), .A2(new_n3934_), .ZN(new_n4291_));
  AOI22_X1   g04024(.A1(new_n4291_), .A2(new_n3939_), .B1(new_n3753_), .B2(new_n4024_), .ZN(new_n4292_));
  INV_X1     g04025(.I(new_n4205_), .ZN(new_n4293_));
  XOR2_X1    g04026(.A1(new_n4201_), .A2(new_n4192_), .Z(new_n4294_));
  NOR2_X1    g04027(.A1(new_n4294_), .A2(new_n4202_), .ZN(new_n4295_));
  INV_X1     g04028(.I(new_n4295_), .ZN(new_n4296_));
  OAI22_X1   g04029(.A1(new_n1055_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n1061_), .ZN(new_n4297_));
  OAI21_X1   g04030(.A1(new_n1294_), .A2(new_n1332_), .B(new_n4297_), .ZN(new_n4298_));
  AOI21_X1   g04031(.A1(new_n4298_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n4299_));
  XOR2_X1    g04032(.A1(new_n1530_), .A2(new_n4299_), .Z(new_n4300_));
  OAI21_X1   g04033(.A1(new_n4147_), .A2(new_n4141_), .B(new_n4140_), .ZN(new_n4301_));
  INV_X1     g04034(.I(new_n4041_), .ZN(new_n4302_));
  NOR2_X1    g04035(.A1(new_n4042_), .A2(new_n3858_), .ZN(new_n4303_));
  NAND2_X1   g04036(.A1(new_n4303_), .A2(new_n3792_), .ZN(new_n4304_));
  NAND2_X1   g04037(.A1(new_n4304_), .A2(new_n4302_), .ZN(new_n4305_));
  INV_X1     g04038(.I(new_n4122_), .ZN(new_n4306_));
  NAND2_X1   g04039(.A1(new_n4111_), .A2(new_n3853_), .ZN(new_n4307_));
  OAI22_X1   g04040(.A1(new_n472_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n515_), .ZN(new_n4308_));
  OAI21_X1   g04041(.A1(new_n420_), .A2(new_n2884_), .B(new_n4308_), .ZN(new_n4309_));
  AOI21_X1   g04042(.A1(new_n4309_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n4310_));
  XOR2_X1    g04043(.A1(new_n700_), .A2(new_n4310_), .Z(new_n4311_));
  INV_X1     g04044(.I(new_n4311_), .ZN(new_n4312_));
  NAND3_X1   g04045(.A1(new_n4081_), .A2(new_n4076_), .A3(new_n4079_), .ZN(new_n4313_));
  NOR2_X1    g04046(.A1(new_n4067_), .A2(new_n280_), .ZN(new_n4314_));
  AOI21_X1   g04047(.A1(new_n269_), .A2(new_n490_), .B(new_n4072_), .ZN(new_n4315_));
  NOR2_X1    g04048(.A1(new_n4315_), .A2(new_n4314_), .ZN(new_n4316_));
  XOR2_X1    g04049(.A1(\a[32] ), .A2(\a[35] ), .Z(new_n4317_));
  NAND3_X1   g04050(.A1(new_n4071_), .A2(new_n3793_), .A3(new_n4317_), .ZN(new_n4318_));
  INV_X1     g04051(.I(new_n4318_), .ZN(new_n4319_));
  NAND2_X1   g04052(.A1(new_n4319_), .A2(\b[0] ), .ZN(new_n4320_));
  OAI21_X1   g04053(.A1(new_n4316_), .A2(new_n4320_), .B(\a[35] ), .ZN(new_n4321_));
  INV_X1     g04054(.I(new_n4321_), .ZN(new_n4322_));
  NOR3_X1    g04055(.A1(new_n4316_), .A2(\a[35] ), .A3(new_n4320_), .ZN(new_n4323_));
  NOR2_X1    g04056(.A1(new_n4322_), .A2(new_n4323_), .ZN(new_n4324_));
  XOR2_X1    g04057(.A1(new_n4324_), .A2(new_n4313_), .Z(new_n4325_));
  NAND2_X1   g04058(.A1(new_n3813_), .A2(new_n3802_), .ZN(new_n4326_));
  NOR4_X1    g04059(.A1(new_n3366_), .A2(new_n3360_), .A3(new_n3363_), .A4(new_n3794_), .ZN(new_n4327_));
  OAI21_X1   g04060(.A1(new_n3813_), .A2(new_n3802_), .B(new_n4327_), .ZN(new_n4328_));
  AOI22_X1   g04061(.A1(new_n4326_), .A2(new_n4328_), .B1(new_n4083_), .B2(new_n4085_), .ZN(new_n4329_));
  NAND2_X1   g04062(.A1(new_n378_), .A2(new_n3346_), .ZN(new_n4330_));
  INV_X1     g04063(.I(new_n3569_), .ZN(new_n4331_));
  AOI22_X1   g04064(.A1(new_n3346_), .A2(\b[4] ), .B1(\b[5] ), .B2(new_n3351_), .ZN(new_n4332_));
  AOI21_X1   g04065(.A1(\b[3] ), .A2(new_n4331_), .B(new_n4332_), .ZN(new_n4333_));
  NAND2_X1   g04066(.A1(new_n4330_), .A2(new_n4333_), .ZN(new_n4334_));
  XOR2_X1    g04067(.A1(new_n4334_), .A2(\a[32] ), .Z(new_n4335_));
  NOR3_X1    g04068(.A1(new_n4329_), .A2(new_n4090_), .A3(new_n4335_), .ZN(new_n4336_));
  NAND2_X1   g04069(.A1(new_n4059_), .A2(new_n4086_), .ZN(new_n4337_));
  OAI22_X1   g04070(.A1(new_n4054_), .A2(new_n4052_), .B1(new_n4059_), .B2(new_n4086_), .ZN(new_n4338_));
  INV_X1     g04071(.I(new_n4335_), .ZN(new_n4339_));
  AOI21_X1   g04072(.A1(new_n4338_), .A2(new_n4337_), .B(new_n4339_), .ZN(new_n4340_));
  OAI21_X1   g04073(.A1(new_n4336_), .A2(new_n4340_), .B(new_n4325_), .ZN(new_n4341_));
  INV_X1     g04074(.I(new_n4325_), .ZN(new_n4342_));
  NAND3_X1   g04075(.A1(new_n4338_), .A2(new_n4337_), .A3(new_n4339_), .ZN(new_n4343_));
  OAI21_X1   g04076(.A1(new_n4329_), .A2(new_n4090_), .B(new_n4335_), .ZN(new_n4344_));
  NAND3_X1   g04077(.A1(new_n4344_), .A2(new_n4343_), .A3(new_n4342_), .ZN(new_n4345_));
  AOI21_X1   g04078(.A1(new_n4341_), .A2(new_n4345_), .B(new_n4312_), .ZN(new_n4346_));
  AOI21_X1   g04079(.A1(new_n4344_), .A2(new_n4343_), .B(new_n4342_), .ZN(new_n4347_));
  NOR3_X1    g04080(.A1(new_n4336_), .A2(new_n4340_), .A3(new_n4325_), .ZN(new_n4348_));
  NOR3_X1    g04081(.A1(new_n4348_), .A2(new_n4347_), .A3(new_n4311_), .ZN(new_n4349_));
  OAI21_X1   g04082(.A1(new_n4349_), .A2(new_n4346_), .B(new_n4114_), .ZN(new_n4350_));
  NOR2_X1    g04083(.A1(new_n4350_), .A2(new_n4099_), .ZN(new_n4351_));
  OAI21_X1   g04084(.A1(new_n4348_), .A2(new_n4347_), .B(new_n4311_), .ZN(new_n4352_));
  NAND3_X1   g04085(.A1(new_n4341_), .A2(new_n4345_), .A3(new_n4312_), .ZN(new_n4353_));
  NAND2_X1   g04086(.A1(new_n4352_), .A2(new_n4353_), .ZN(new_n4354_));
  NOR2_X1    g04087(.A1(new_n4093_), .A2(new_n4098_), .ZN(new_n4356_));
  OAI21_X1   g04088(.A1(new_n4351_), .A2(new_n4356_), .B(new_n4307_), .ZN(new_n4357_));
  NOR2_X1    g04089(.A1(new_n4051_), .A2(new_n3847_), .ZN(new_n4358_));
  INV_X1     g04090(.I(new_n4099_), .ZN(new_n4359_));
  NAND3_X1   g04091(.A1(new_n4354_), .A2(new_n4359_), .A3(new_n4114_), .ZN(new_n4360_));
  INV_X1     g04092(.I(new_n4356_), .ZN(new_n4361_));
  NAND3_X1   g04093(.A1(new_n4360_), .A2(new_n4358_), .A3(new_n4361_), .ZN(new_n4362_));
  OAI22_X1   g04094(.A1(new_n2171_), .A2(new_n656_), .B1(new_n706_), .B2(new_n2166_), .ZN(new_n4363_));
  OAI21_X1   g04095(.A1(new_n565_), .A2(new_n2322_), .B(new_n4363_), .ZN(new_n4364_));
  AOI21_X1   g04096(.A1(new_n4364_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n4365_));
  XNOR2_X1   g04097(.A1(new_n710_), .A2(new_n4365_), .ZN(new_n4366_));
  INV_X1     g04098(.I(new_n4366_), .ZN(new_n4367_));
  NAND3_X1   g04099(.A1(new_n4357_), .A2(new_n4362_), .A3(new_n4367_), .ZN(new_n4368_));
  AOI21_X1   g04100(.A1(new_n4360_), .A2(new_n4361_), .B(new_n4358_), .ZN(new_n4369_));
  NOR3_X1    g04101(.A1(new_n4351_), .A2(new_n4307_), .A3(new_n4356_), .ZN(new_n4370_));
  OAI21_X1   g04102(.A1(new_n4370_), .A2(new_n4369_), .B(new_n4366_), .ZN(new_n4371_));
  NAND2_X1   g04103(.A1(new_n4371_), .A2(new_n4368_), .ZN(new_n4372_));
  NAND3_X1   g04104(.A1(new_n4372_), .A2(new_n4306_), .A3(new_n4133_), .ZN(new_n4373_));
  NOR2_X1    g04105(.A1(new_n4117_), .A2(new_n4121_), .ZN(new_n4375_));
  INV_X1     g04106(.I(new_n4375_), .ZN(new_n4376_));
  AOI21_X1   g04107(.A1(new_n4373_), .A2(new_n4376_), .B(new_n4305_), .ZN(new_n4377_));
  NOR3_X1    g04108(.A1(new_n4370_), .A2(new_n4369_), .A3(new_n4366_), .ZN(new_n4378_));
  AOI21_X1   g04109(.A1(new_n4357_), .A2(new_n4362_), .B(new_n4367_), .ZN(new_n4379_));
  OAI21_X1   g04110(.A1(new_n4378_), .A2(new_n4379_), .B(new_n4133_), .ZN(new_n4380_));
  NOR2_X1    g04111(.A1(new_n4380_), .A2(new_n4122_), .ZN(new_n4381_));
  NOR3_X1    g04112(.A1(new_n4381_), .A2(new_n4130_), .A3(new_n4375_), .ZN(new_n4382_));
  OAI22_X1   g04113(.A1(new_n1712_), .A2(new_n861_), .B1(new_n930_), .B2(new_n1707_), .ZN(new_n4383_));
  OAI21_X1   g04114(.A1(new_n780_), .A2(new_n1850_), .B(new_n4383_), .ZN(new_n4384_));
  AOI21_X1   g04115(.A1(new_n4384_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n4385_));
  XNOR2_X1   g04116(.A1(new_n937_), .A2(new_n4385_), .ZN(new_n4386_));
  NOR3_X1    g04117(.A1(new_n4382_), .A2(new_n4377_), .A3(new_n4386_), .ZN(new_n4387_));
  OAI21_X1   g04118(.A1(new_n4381_), .A2(new_n4375_), .B(new_n4130_), .ZN(new_n4388_));
  NAND3_X1   g04119(.A1(new_n4373_), .A2(new_n4305_), .A3(new_n4376_), .ZN(new_n4389_));
  INV_X1     g04120(.I(new_n4386_), .ZN(new_n4390_));
  AOI21_X1   g04121(.A1(new_n4388_), .A2(new_n4389_), .B(new_n4390_), .ZN(new_n4391_));
  OAI22_X1   g04122(.A1(new_n1347_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n1344_), .ZN(new_n4392_));
  OAI21_X1   g04123(.A1(new_n1017_), .A2(new_n1457_), .B(new_n4392_), .ZN(new_n4393_));
  AOI21_X1   g04124(.A1(new_n4393_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n4394_));
  XNOR2_X1   g04125(.A1(new_n1196_), .A2(new_n4394_), .ZN(new_n4395_));
  NOR3_X1    g04126(.A1(new_n4387_), .A2(new_n4391_), .A3(new_n4395_), .ZN(new_n4396_));
  NAND3_X1   g04127(.A1(new_n4388_), .A2(new_n4389_), .A3(new_n4390_), .ZN(new_n4397_));
  OAI21_X1   g04128(.A1(new_n4382_), .A2(new_n4377_), .B(new_n4386_), .ZN(new_n4398_));
  INV_X1     g04129(.I(new_n4395_), .ZN(new_n4399_));
  AOI21_X1   g04130(.A1(new_n4398_), .A2(new_n4397_), .B(new_n4399_), .ZN(new_n4400_));
  OAI21_X1   g04131(.A1(new_n4396_), .A2(new_n4400_), .B(new_n4301_), .ZN(new_n4401_));
  AOI21_X1   g04132(.A1(new_n4039_), .A2(new_n4142_), .B(new_n4162_), .ZN(new_n4402_));
  AOI21_X1   g04133(.A1(new_n4398_), .A2(new_n4397_), .B(new_n4395_), .ZN(new_n4403_));
  NOR3_X1    g04134(.A1(new_n4387_), .A2(new_n4391_), .A3(new_n4399_), .ZN(new_n4404_));
  OAI21_X1   g04135(.A1(new_n4404_), .A2(new_n4403_), .B(new_n4402_), .ZN(new_n4405_));
  NAND2_X1   g04136(.A1(new_n4405_), .A2(new_n4401_), .ZN(new_n4406_));
  NAND3_X1   g04137(.A1(new_n4144_), .A2(new_n4154_), .A3(new_n4160_), .ZN(new_n4407_));
  OAI21_X1   g04138(.A1(new_n4166_), .A2(new_n4164_), .B(new_n4159_), .ZN(new_n4408_));
  NAND2_X1   g04139(.A1(new_n4408_), .A2(new_n4407_), .ZN(new_n4409_));
  NAND3_X1   g04140(.A1(new_n4406_), .A2(new_n4409_), .A3(new_n4161_), .ZN(new_n4410_));
  NAND2_X1   g04141(.A1(new_n4398_), .A2(new_n4397_), .ZN(new_n4411_));
  INV_X1     g04142(.I(new_n4411_), .ZN(new_n4412_));
  NOR2_X1    g04143(.A1(new_n4167_), .A2(new_n4159_), .ZN(new_n4413_));
  INV_X1     g04144(.I(new_n4413_), .ZN(new_n4414_));
  AOI21_X1   g04145(.A1(new_n4410_), .A2(new_n4414_), .B(new_n4175_), .ZN(new_n4415_));
  NOR2_X1    g04146(.A1(new_n4167_), .A2(new_n4159_), .ZN(new_n4416_));
  NAND3_X1   g04147(.A1(new_n4398_), .A2(new_n4397_), .A3(new_n4399_), .ZN(new_n4417_));
  OAI21_X1   g04148(.A1(new_n4387_), .A2(new_n4391_), .B(new_n4395_), .ZN(new_n4418_));
  AOI21_X1   g04149(.A1(new_n4418_), .A2(new_n4417_), .B(new_n4402_), .ZN(new_n4419_));
  OAI21_X1   g04150(.A1(new_n4387_), .A2(new_n4391_), .B(new_n4399_), .ZN(new_n4420_));
  NAND3_X1   g04151(.A1(new_n4398_), .A2(new_n4397_), .A3(new_n4395_), .ZN(new_n4421_));
  AOI21_X1   g04152(.A1(new_n4420_), .A2(new_n4421_), .B(new_n4301_), .ZN(new_n4422_));
  NOR2_X1    g04153(.A1(new_n4419_), .A2(new_n4422_), .ZN(new_n4423_));
  NOR3_X1    g04154(.A1(new_n4166_), .A2(new_n4164_), .A3(new_n4159_), .ZN(new_n4424_));
  AOI21_X1   g04155(.A1(new_n4144_), .A2(new_n4154_), .B(new_n4160_), .ZN(new_n4425_));
  NOR2_X1    g04156(.A1(new_n4424_), .A2(new_n4425_), .ZN(new_n4426_));
  NOR3_X1    g04157(.A1(new_n4423_), .A2(new_n4426_), .A3(new_n4416_), .ZN(new_n4427_));
  NOR3_X1    g04158(.A1(new_n4427_), .A2(new_n4186_), .A3(new_n4413_), .ZN(new_n4428_));
  NOR2_X1    g04159(.A1(new_n4428_), .A2(new_n4415_), .ZN(new_n4429_));
  INV_X1     g04160(.I(new_n4429_), .ZN(new_n4430_));
  OR2_X2     g04161(.A1(new_n4188_), .A2(new_n4191_), .Z(new_n4431_));
  NOR2_X1    g04162(.A1(new_n4186_), .A2(new_n4169_), .ZN(new_n4432_));
  NOR2_X1    g04163(.A1(new_n4170_), .A2(new_n4175_), .ZN(new_n4433_));
  OAI21_X1   g04164(.A1(new_n4433_), .A2(new_n4432_), .B(new_n4179_), .ZN(new_n4434_));
  OAI21_X1   g04165(.A1(new_n4201_), .A2(new_n4431_), .B(new_n4434_), .ZN(new_n4435_));
  OAI22_X1   g04166(.A1(new_n970_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n820_), .ZN(new_n4436_));
  OAI21_X1   g04167(.A1(new_n1634_), .A2(new_n894_), .B(new_n4436_), .ZN(new_n4437_));
  AOI21_X1   g04168(.A1(new_n4437_), .A2(new_n827_), .B(new_n970_), .ZN(new_n4438_));
  XNOR2_X1   g04169(.A1(new_n1940_), .A2(new_n4438_), .ZN(new_n4439_));
  INV_X1     g04170(.I(new_n4439_), .ZN(new_n4440_));
  NAND2_X1   g04171(.A1(new_n4435_), .A2(new_n4440_), .ZN(new_n4441_));
  NAND2_X1   g04172(.A1(new_n4034_), .A2(new_n4192_), .ZN(new_n4442_));
  NAND3_X1   g04173(.A1(new_n4442_), .A2(new_n4434_), .A3(new_n4439_), .ZN(new_n4443_));
  AOI21_X1   g04174(.A1(new_n4441_), .A2(new_n4443_), .B(new_n4430_), .ZN(new_n4444_));
  AOI21_X1   g04175(.A1(new_n4442_), .A2(new_n4434_), .B(new_n4439_), .ZN(new_n4445_));
  NOR2_X1    g04176(.A1(new_n4435_), .A2(new_n4440_), .ZN(new_n4446_));
  NOR3_X1    g04177(.A1(new_n4446_), .A2(new_n4445_), .A3(new_n4429_), .ZN(new_n4447_));
  OAI21_X1   g04178(.A1(new_n4447_), .A2(new_n4444_), .B(new_n4300_), .ZN(new_n4448_));
  INV_X1     g04179(.I(new_n4300_), .ZN(new_n4449_));
  OAI21_X1   g04180(.A1(new_n4446_), .A2(new_n4445_), .B(new_n4429_), .ZN(new_n4450_));
  NAND3_X1   g04181(.A1(new_n4441_), .A2(new_n4443_), .A3(new_n4430_), .ZN(new_n4451_));
  NAND3_X1   g04182(.A1(new_n4450_), .A2(new_n4451_), .A3(new_n4449_), .ZN(new_n4452_));
  NAND3_X1   g04183(.A1(new_n4448_), .A2(new_n4452_), .A3(new_n4296_), .ZN(new_n4453_));
  NAND3_X1   g04184(.A1(new_n4292_), .A2(new_n4453_), .A3(new_n4293_), .ZN(new_n4454_));
  AOI21_X1   g04185(.A1(new_n4450_), .A2(new_n4451_), .B(new_n4449_), .ZN(new_n4455_));
  NOR3_X1    g04186(.A1(new_n4447_), .A2(new_n4444_), .A3(new_n4300_), .ZN(new_n4456_));
  NOR3_X1    g04187(.A1(new_n4456_), .A2(new_n4455_), .A3(new_n4295_), .ZN(new_n4457_));
  OAI21_X1   g04188(.A1(new_n4457_), .A2(new_n4205_), .B(new_n4028_), .ZN(new_n4458_));
  OAI22_X1   g04189(.A1(new_n607_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n610_), .ZN(new_n4459_));
  OAI21_X1   g04190(.A1(new_n2102_), .A2(new_n684_), .B(new_n4459_), .ZN(new_n4460_));
  AOI21_X1   g04191(.A1(new_n4460_), .A2(new_n612_), .B(new_n607_), .ZN(new_n4461_));
  XNOR2_X1   g04192(.A1(new_n2443_), .A2(new_n4461_), .ZN(new_n4462_));
  AOI21_X1   g04193(.A1(new_n4458_), .A2(new_n4454_), .B(new_n4462_), .ZN(new_n4463_));
  NOR3_X1    g04194(.A1(new_n4457_), .A2(new_n4028_), .A3(new_n4205_), .ZN(new_n4464_));
  AOI21_X1   g04195(.A1(new_n4293_), .A2(new_n4453_), .B(new_n4292_), .ZN(new_n4465_));
  INV_X1     g04196(.I(new_n4462_), .ZN(new_n4466_));
  NOR3_X1    g04197(.A1(new_n4465_), .A2(new_n4464_), .A3(new_n4466_), .ZN(new_n4467_));
  OR2_X2     g04198(.A1(new_n4467_), .A2(new_n4463_), .Z(new_n4468_));
  OAI22_X1   g04199(.A1(new_n448_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n450_), .ZN(new_n4469_));
  OAI21_X1   g04200(.A1(new_n2643_), .A2(new_n496_), .B(new_n4469_), .ZN(new_n4470_));
  AOI21_X1   g04201(.A1(new_n4470_), .A2(new_n452_), .B(new_n448_), .ZN(new_n4471_));
  XNOR2_X1   g04202(.A1(new_n3022_), .A2(new_n4471_), .ZN(new_n4472_));
  NOR2_X1    g04203(.A1(new_n4468_), .A2(new_n4472_), .ZN(new_n4473_));
  NOR2_X1    g04204(.A1(new_n4467_), .A2(new_n4463_), .ZN(new_n4474_));
  INV_X1     g04205(.I(new_n4472_), .ZN(new_n4475_));
  NOR2_X1    g04206(.A1(new_n4474_), .A2(new_n4475_), .ZN(new_n4476_));
  NOR2_X1    g04207(.A1(new_n4473_), .A2(new_n4476_), .ZN(new_n4477_));
  NOR2_X1    g04208(.A1(new_n4477_), .A2(new_n4287_), .ZN(new_n4478_));
  NAND2_X1   g04209(.A1(new_n4023_), .A2(new_n4214_), .ZN(new_n4479_));
  NAND2_X1   g04210(.A1(new_n4479_), .A2(new_n4212_), .ZN(new_n4480_));
  XOR2_X1    g04211(.A1(new_n4474_), .A2(new_n4472_), .Z(new_n4481_));
  NOR2_X1    g04212(.A1(new_n4480_), .A2(new_n4481_), .ZN(new_n4482_));
  NOR2_X1    g04213(.A1(new_n4482_), .A2(new_n4478_), .ZN(new_n4483_));
  XOR2_X1    g04214(.A1(new_n4218_), .A2(new_n4223_), .Z(new_n4484_));
  NOR3_X1    g04215(.A1(new_n4484_), .A2(new_n4224_), .A3(new_n4483_), .ZN(new_n4485_));
  NOR2_X1    g04216(.A1(new_n4219_), .A2(new_n4223_), .ZN(new_n4486_));
  OR2_X2     g04217(.A1(new_n4485_), .A2(new_n4486_), .Z(new_n4487_));
  XOR2_X1    g04218(.A1(new_n4487_), .A2(new_n4231_), .Z(new_n4488_));
  INV_X1     g04219(.I(new_n4488_), .ZN(new_n4489_));
  OAI22_X1   g04220(.A1(new_n3709_), .A2(new_n341_), .B1(new_n404_), .B2(new_n3717_), .ZN(new_n4490_));
  OAI21_X1   g04221(.A1(new_n3260_), .A2(new_n366_), .B(new_n4490_), .ZN(new_n4491_));
  AOI21_X1   g04222(.A1(new_n4491_), .A2(new_n334_), .B(new_n341_), .ZN(new_n4492_));
  XOR2_X1    g04223(.A1(new_n3722_), .A2(new_n4492_), .Z(new_n4493_));
  NOR2_X1    g04224(.A1(new_n4489_), .A2(new_n4493_), .ZN(new_n4494_));
  XOR2_X1    g04225(.A1(new_n4494_), .A2(new_n4239_), .Z(new_n4495_));
  XNOR2_X1   g04226(.A1(new_n4495_), .A2(new_n4285_), .ZN(new_n4496_));
  XNOR2_X1   g04227(.A1(\b[33] ), .A2(\b[35] ), .ZN(new_n4497_));
  NOR2_X1    g04228(.A1(new_n4497_), .A2(new_n4252_), .ZN(new_n4498_));
  XOR2_X1    g04229(.A1(new_n4251_), .A2(new_n4498_), .Z(new_n4499_));
  INV_X1     g04230(.I(\b[35] ), .ZN(new_n4500_));
  OAI22_X1   g04231(.A1(new_n330_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n263_), .ZN(new_n4501_));
  OAI21_X1   g04232(.A1(new_n3989_), .A2(new_n289_), .B(new_n4501_), .ZN(new_n4502_));
  AOI21_X1   g04233(.A1(new_n4502_), .A2(new_n260_), .B(new_n426_), .ZN(new_n4503_));
  XOR2_X1    g04234(.A1(new_n4499_), .A2(new_n4503_), .Z(new_n4504_));
  XOR2_X1    g04235(.A1(new_n4496_), .A2(new_n4504_), .Z(new_n4505_));
  XOR2_X1    g04236(.A1(new_n4496_), .A2(new_n4504_), .Z(new_n4506_));
  NAND2_X1   g04237(.A1(new_n4269_), .A2(new_n4506_), .ZN(new_n4507_));
  OAI21_X1   g04238(.A1(new_n4269_), .A2(new_n4505_), .B(new_n4507_), .ZN(\f[35] ));
  INV_X1     g04239(.I(new_n4504_), .ZN(new_n4509_));
  NAND2_X1   g04240(.A1(new_n4496_), .A2(new_n4509_), .ZN(new_n4510_));
  NAND3_X1   g04241(.A1(new_n4284_), .A2(new_n4282_), .A3(new_n4488_), .ZN(new_n4511_));
  AOI21_X1   g04242(.A1(new_n4284_), .A2(new_n4282_), .B(new_n4488_), .ZN(new_n4512_));
  OR2_X2     g04243(.A1(new_n4238_), .A2(new_n4493_), .Z(new_n4513_));
  OAI21_X1   g04244(.A1(new_n4512_), .A2(new_n4513_), .B(new_n4511_), .ZN(new_n4514_));
  OAI21_X1   g04245(.A1(new_n4483_), .A2(new_n4223_), .B(new_n4219_), .ZN(new_n4515_));
  NAND2_X1   g04246(.A1(new_n4483_), .A2(new_n4223_), .ZN(new_n4516_));
  NAND3_X1   g04247(.A1(new_n4515_), .A2(new_n4231_), .A3(new_n4516_), .ZN(new_n4517_));
  XOR2_X1    g04248(.A1(new_n4287_), .A2(new_n4474_), .Z(new_n4518_));
  NOR2_X1    g04249(.A1(new_n4518_), .A2(new_n4475_), .ZN(new_n4519_));
  INV_X1     g04250(.I(new_n4519_), .ZN(new_n4520_));
  NAND2_X1   g04251(.A1(new_n4517_), .A2(new_n4520_), .ZN(new_n4521_));
  AOI21_X1   g04252(.A1(new_n4458_), .A2(new_n4454_), .B(new_n4466_), .ZN(new_n4522_));
  OAI21_X1   g04253(.A1(new_n4474_), .A2(new_n4206_), .B(new_n4210_), .ZN(new_n4523_));
  NAND2_X1   g04254(.A1(new_n4474_), .A2(new_n4206_), .ZN(new_n4524_));
  AND3_X2    g04255(.A1(new_n4023_), .A2(new_n4523_), .A3(new_n4524_), .Z(new_n4525_));
  NAND2_X1   g04256(.A1(new_n4435_), .A2(new_n4430_), .ZN(new_n4526_));
  NAND3_X1   g04257(.A1(new_n4442_), .A2(new_n4429_), .A3(new_n4434_), .ZN(new_n4527_));
  AOI21_X1   g04258(.A1(new_n4526_), .A2(new_n4527_), .B(new_n4449_), .ZN(new_n4528_));
  INV_X1     g04259(.I(new_n4528_), .ZN(new_n4529_));
  NAND3_X1   g04260(.A1(new_n4526_), .A2(new_n4527_), .A3(new_n4449_), .ZN(new_n4530_));
  NAND2_X1   g04261(.A1(new_n4529_), .A2(new_n4530_), .ZN(new_n4531_));
  NAND2_X1   g04262(.A1(new_n4531_), .A2(new_n4440_), .ZN(new_n4532_));
  OAI21_X1   g04263(.A1(new_n4456_), .A2(new_n4455_), .B(new_n4295_), .ZN(new_n4533_));
  AOI21_X1   g04264(.A1(new_n4533_), .A2(new_n4205_), .B(new_n4292_), .ZN(new_n4534_));
  OAI21_X1   g04265(.A1(new_n4428_), .A2(new_n4415_), .B(new_n4300_), .ZN(new_n4535_));
  OAI21_X1   g04266(.A1(new_n4428_), .A2(new_n4415_), .B(new_n4449_), .ZN(new_n4536_));
  OAI21_X1   g04267(.A1(new_n4427_), .A2(new_n4413_), .B(new_n4186_), .ZN(new_n4537_));
  NAND3_X1   g04268(.A1(new_n4410_), .A2(new_n4175_), .A3(new_n4414_), .ZN(new_n4538_));
  NAND3_X1   g04269(.A1(new_n4537_), .A2(new_n4538_), .A3(new_n4300_), .ZN(new_n4539_));
  AOI21_X1   g04270(.A1(new_n4536_), .A2(new_n4539_), .B(new_n4434_), .ZN(new_n4540_));
  OAI21_X1   g04271(.A1(new_n4540_), .A2(new_n4431_), .B(new_n4201_), .ZN(new_n4541_));
  NAND2_X1   g04272(.A1(new_n4301_), .A2(new_n4411_), .ZN(new_n4542_));
  NAND2_X1   g04273(.A1(new_n4412_), .A2(new_n4402_), .ZN(new_n4543_));
  AOI21_X1   g04274(.A1(new_n4543_), .A2(new_n4542_), .B(new_n4399_), .ZN(new_n4544_));
  INV_X1     g04275(.I(new_n4544_), .ZN(new_n4545_));
  AOI21_X1   g04276(.A1(new_n4406_), .A2(new_n4160_), .B(new_n4155_), .ZN(new_n4546_));
  NAND3_X1   g04277(.A1(new_n4405_), .A2(new_n4401_), .A3(new_n4159_), .ZN(new_n4547_));
  NAND2_X1   g04278(.A1(new_n4175_), .A2(new_n4547_), .ZN(new_n4548_));
  NOR2_X1    g04279(.A1(new_n4548_), .A2(new_n4546_), .ZN(new_n4549_));
  NOR3_X1    g04280(.A1(new_n4382_), .A2(new_n4377_), .A3(new_n4390_), .ZN(new_n4550_));
  NAND2_X1   g04281(.A1(new_n4134_), .A2(new_n4129_), .ZN(new_n4551_));
  AOI21_X1   g04282(.A1(new_n4411_), .A2(new_n4551_), .B(new_n4139_), .ZN(new_n4552_));
  OAI21_X1   g04283(.A1(new_n4411_), .A2(new_n4551_), .B(new_n4039_), .ZN(new_n4553_));
  AOI21_X1   g04284(.A1(new_n4372_), .A2(new_n4126_), .B(new_n4127_), .ZN(new_n4554_));
  NAND3_X1   g04285(.A1(new_n4371_), .A2(new_n4368_), .A3(new_n4117_), .ZN(new_n4555_));
  NAND2_X1   g04286(.A1(new_n4305_), .A2(new_n4555_), .ZN(new_n4556_));
  NOR2_X1    g04287(.A1(new_n4556_), .A2(new_n4554_), .ZN(new_n4557_));
  NAND2_X1   g04288(.A1(new_n4338_), .A2(new_n4337_), .ZN(new_n4558_));
  XOR2_X1    g04289(.A1(new_n4558_), .A2(new_n4342_), .Z(new_n4559_));
  NAND2_X1   g04290(.A1(new_n4559_), .A2(new_n4335_), .ZN(new_n4560_));
  XOR2_X1    g04291(.A1(new_n4558_), .A2(new_n4325_), .Z(new_n4561_));
  NAND2_X1   g04292(.A1(new_n4561_), .A2(new_n4339_), .ZN(new_n4562_));
  AOI21_X1   g04293(.A1(new_n4560_), .A2(new_n4562_), .B(new_n4311_), .ZN(new_n4563_));
  AOI21_X1   g04294(.A1(new_n4354_), .A2(new_n4103_), .B(new_n4104_), .ZN(new_n4564_));
  OAI21_X1   g04295(.A1(new_n4103_), .A2(new_n4354_), .B(new_n4358_), .ZN(new_n4565_));
  XOR2_X1    g04296(.A1(\a[35] ), .A2(\a[36] ), .Z(new_n4566_));
  NAND2_X1   g04297(.A1(new_n4566_), .A2(\b[0] ), .ZN(new_n4567_));
  NOR2_X1    g04298(.A1(new_n4318_), .A2(new_n269_), .ZN(new_n4568_));
  OAI22_X1   g04299(.A1(new_n280_), .A2(new_n4072_), .B1(new_n4067_), .B2(new_n298_), .ZN(new_n4569_));
  NOR2_X1    g04300(.A1(new_n4569_), .A2(new_n4568_), .ZN(new_n4570_));
  NOR3_X1    g04301(.A1(new_n4570_), .A2(new_n403_), .A3(new_n4072_), .ZN(new_n4571_));
  XOR2_X1    g04302(.A1(new_n4571_), .A2(\a[35] ), .Z(new_n4572_));
  INV_X1     g04303(.I(new_n4323_), .ZN(new_n4573_));
  NAND2_X1   g04304(.A1(new_n4573_), .A2(new_n4321_), .ZN(new_n4574_));
  AOI22_X1   g04305(.A1(new_n3346_), .A2(\b[5] ), .B1(\b[6] ), .B2(new_n3351_), .ZN(new_n4575_));
  NOR2_X1    g04306(.A1(new_n3569_), .A2(new_n325_), .ZN(new_n4576_));
  NOR2_X1    g04307(.A1(new_n4575_), .A2(new_n4576_), .ZN(new_n4577_));
  OAI21_X1   g04308(.A1(new_n4577_), .A2(\a[32] ), .B(new_n3346_), .ZN(new_n4578_));
  NOR3_X1    g04309(.A1(new_n424_), .A2(new_n417_), .A3(new_n4578_), .ZN(new_n4579_));
  INV_X1     g04310(.I(new_n4578_), .ZN(new_n4580_));
  AOI21_X1   g04311(.A1(new_n554_), .A2(new_n555_), .B(new_n4580_), .ZN(new_n4581_));
  OAI22_X1   g04312(.A1(new_n4581_), .A2(new_n4579_), .B1(new_n4313_), .B2(new_n4574_), .ZN(new_n4582_));
  NOR2_X1    g04313(.A1(new_n4574_), .A2(new_n4313_), .ZN(new_n4583_));
  NAND3_X1   g04314(.A1(new_n4580_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n4584_));
  OAI21_X1   g04315(.A1(new_n424_), .A2(new_n417_), .B(new_n4578_), .ZN(new_n4585_));
  NAND3_X1   g04316(.A1(new_n4583_), .A2(new_n4584_), .A3(new_n4585_), .ZN(new_n4586_));
  AOI21_X1   g04317(.A1(new_n4586_), .A2(new_n4582_), .B(new_n4572_), .ZN(new_n4587_));
  XOR2_X1    g04318(.A1(new_n4571_), .A2(new_n4069_), .Z(new_n4588_));
  NOR3_X1    g04319(.A1(new_n4077_), .A2(new_n4075_), .A3(new_n4078_), .ZN(new_n4589_));
  AOI22_X1   g04320(.A1(new_n4584_), .A2(new_n4585_), .B1(new_n4589_), .B2(new_n4324_), .ZN(new_n4590_));
  NAND2_X1   g04321(.A1(new_n4324_), .A2(new_n4589_), .ZN(new_n4591_));
  NOR3_X1    g04322(.A1(new_n4591_), .A2(new_n4579_), .A3(new_n4581_), .ZN(new_n4592_));
  NOR3_X1    g04323(.A1(new_n4592_), .A2(new_n4590_), .A3(new_n4588_), .ZN(new_n4593_));
  OAI21_X1   g04324(.A1(new_n4593_), .A2(new_n4587_), .B(new_n4567_), .ZN(new_n4594_));
  INV_X1     g04325(.I(new_n4567_), .ZN(new_n4595_));
  OAI21_X1   g04326(.A1(new_n4592_), .A2(new_n4590_), .B(new_n4588_), .ZN(new_n4596_));
  NAND3_X1   g04327(.A1(new_n4586_), .A2(new_n4582_), .A3(new_n4572_), .ZN(new_n4597_));
  NAND3_X1   g04328(.A1(new_n4596_), .A2(new_n4597_), .A3(new_n4595_), .ZN(new_n4598_));
  NAND2_X1   g04329(.A1(new_n4594_), .A2(new_n4598_), .ZN(new_n4599_));
  INV_X1     g04330(.I(new_n4599_), .ZN(new_n4600_));
  NOR2_X1    g04331(.A1(new_n4325_), .A2(new_n4339_), .ZN(new_n4601_));
  NOR2_X1    g04332(.A1(new_n4589_), .A2(new_n4334_), .ZN(new_n4602_));
  INV_X1     g04333(.I(new_n4334_), .ZN(new_n4603_));
  NOR2_X1    g04334(.A1(new_n4313_), .A2(new_n4603_), .ZN(new_n4604_));
  OAI21_X1   g04335(.A1(new_n4602_), .A2(new_n4604_), .B(new_n4324_), .ZN(new_n4605_));
  NAND2_X1   g04336(.A1(new_n4313_), .A2(new_n4603_), .ZN(new_n4606_));
  NAND2_X1   g04337(.A1(new_n4589_), .A2(new_n4334_), .ZN(new_n4607_));
  NAND3_X1   g04338(.A1(new_n4607_), .A2(new_n4606_), .A3(new_n4574_), .ZN(new_n4608_));
  AOI21_X1   g04339(.A1(new_n4605_), .A2(new_n4608_), .B(\a[32] ), .ZN(new_n4609_));
  AOI21_X1   g04340(.A1(new_n4607_), .A2(new_n4606_), .B(new_n4574_), .ZN(new_n4610_));
  NOR3_X1    g04341(.A1(new_n4602_), .A2(new_n4604_), .A3(new_n4324_), .ZN(new_n4611_));
  NOR3_X1    g04342(.A1(new_n4610_), .A2(new_n4611_), .A3(new_n3354_), .ZN(new_n4612_));
  OAI21_X1   g04343(.A1(new_n4612_), .A2(new_n4609_), .B(new_n4083_), .ZN(new_n4613_));
  OAI21_X1   g04344(.A1(new_n4610_), .A2(new_n4611_), .B(new_n3354_), .ZN(new_n4614_));
  NAND3_X1   g04345(.A1(new_n4605_), .A2(new_n4608_), .A3(\a[32] ), .ZN(new_n4615_));
  NAND3_X1   g04346(.A1(new_n4614_), .A2(new_n4615_), .A3(new_n4086_), .ZN(new_n4616_));
  NAND2_X1   g04347(.A1(new_n4616_), .A2(new_n4100_), .ZN(new_n4617_));
  AOI21_X1   g04348(.A1(new_n4085_), .A2(new_n4613_), .B(new_n4617_), .ZN(new_n4618_));
  OAI21_X1   g04349(.A1(new_n4618_), .A2(new_n4601_), .B(new_n4600_), .ZN(new_n4619_));
  INV_X1     g04350(.I(new_n4601_), .ZN(new_n4620_));
  NAND2_X1   g04351(.A1(new_n4613_), .A2(new_n4085_), .ZN(new_n4621_));
  NAND3_X1   g04352(.A1(new_n4621_), .A2(new_n4100_), .A3(new_n4616_), .ZN(new_n4622_));
  NAND3_X1   g04353(.A1(new_n4622_), .A2(new_n4599_), .A3(new_n4620_), .ZN(new_n4623_));
  OAI22_X1   g04354(.A1(new_n515_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n565_), .ZN(new_n4624_));
  OAI21_X1   g04355(.A1(new_n472_), .A2(new_n2884_), .B(new_n4624_), .ZN(new_n4625_));
  AOI21_X1   g04356(.A1(new_n4625_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n4626_));
  XOR2_X1    g04357(.A1(new_n759_), .A2(new_n4626_), .Z(new_n4627_));
  AOI21_X1   g04358(.A1(new_n4619_), .A2(new_n4623_), .B(new_n4627_), .ZN(new_n4628_));
  OAI21_X1   g04359(.A1(new_n4565_), .A2(new_n4564_), .B(new_n4628_), .ZN(new_n4629_));
  INV_X1     g04360(.I(new_n4564_), .ZN(new_n4630_));
  NOR2_X1    g04361(.A1(new_n4354_), .A2(new_n4103_), .ZN(new_n4631_));
  NOR2_X1    g04362(.A1(new_n4307_), .A2(new_n4631_), .ZN(new_n4632_));
  INV_X1     g04363(.I(new_n4628_), .ZN(new_n4633_));
  NAND3_X1   g04364(.A1(new_n4633_), .A2(new_n4632_), .A3(new_n4630_), .ZN(new_n4634_));
  AOI21_X1   g04365(.A1(new_n4629_), .A2(new_n4634_), .B(new_n4563_), .ZN(new_n4635_));
  NAND3_X1   g04366(.A1(new_n4629_), .A2(new_n4634_), .A3(new_n4563_), .ZN(new_n4636_));
  INV_X1     g04367(.I(new_n4636_), .ZN(new_n4637_));
  OAI22_X1   g04368(.A1(new_n2171_), .A2(new_n706_), .B1(new_n780_), .B2(new_n2166_), .ZN(new_n4638_));
  OAI21_X1   g04369(.A1(new_n656_), .A2(new_n2322_), .B(new_n4638_), .ZN(new_n4639_));
  AOI21_X1   g04370(.A1(new_n4639_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n4640_));
  XOR2_X1    g04371(.A1(new_n785_), .A2(new_n4640_), .Z(new_n4641_));
  INV_X1     g04372(.I(new_n4641_), .ZN(new_n4642_));
  OAI21_X1   g04373(.A1(new_n4637_), .A2(new_n4635_), .B(new_n4642_), .ZN(new_n4643_));
  NOR2_X1    g04374(.A1(new_n4557_), .A2(new_n4643_), .ZN(new_n4644_));
  OAI21_X1   g04375(.A1(new_n4378_), .A2(new_n4379_), .B(new_n4126_), .ZN(new_n4645_));
  NAND2_X1   g04376(.A1(new_n4645_), .A2(new_n4121_), .ZN(new_n4646_));
  NAND3_X1   g04377(.A1(new_n4646_), .A2(new_n4305_), .A3(new_n4555_), .ZN(new_n4647_));
  NOR2_X1    g04378(.A1(new_n4561_), .A2(new_n4339_), .ZN(new_n4648_));
  NOR2_X1    g04379(.A1(new_n4559_), .A2(new_n4335_), .ZN(new_n4649_));
  OAI21_X1   g04380(.A1(new_n4648_), .A2(new_n4649_), .B(new_n4312_), .ZN(new_n4650_));
  AOI21_X1   g04381(.A1(new_n4630_), .A2(new_n4632_), .B(new_n4633_), .ZN(new_n4651_));
  INV_X1     g04382(.I(new_n4634_), .ZN(new_n4652_));
  OAI21_X1   g04383(.A1(new_n4652_), .A2(new_n4651_), .B(new_n4650_), .ZN(new_n4653_));
  AOI21_X1   g04384(.A1(new_n4653_), .A2(new_n4636_), .B(new_n4641_), .ZN(new_n4654_));
  NOR2_X1    g04385(.A1(new_n4647_), .A2(new_n4654_), .ZN(new_n4655_));
  OAI21_X1   g04386(.A1(new_n4644_), .A2(new_n4655_), .B(new_n4371_), .ZN(new_n4656_));
  NAND2_X1   g04387(.A1(new_n4647_), .A2(new_n4654_), .ZN(new_n4657_));
  NAND2_X1   g04388(.A1(new_n4557_), .A2(new_n4643_), .ZN(new_n4658_));
  NAND3_X1   g04389(.A1(new_n4658_), .A2(new_n4657_), .A3(new_n4379_), .ZN(new_n4659_));
  OAI22_X1   g04390(.A1(new_n1712_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n1707_), .ZN(new_n4660_));
  OAI21_X1   g04391(.A1(new_n861_), .A2(new_n1850_), .B(new_n4660_), .ZN(new_n4661_));
  AOI21_X1   g04392(.A1(new_n4661_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n4662_));
  XOR2_X1    g04393(.A1(new_n1024_), .A2(new_n4662_), .Z(new_n4663_));
  AOI21_X1   g04394(.A1(new_n4656_), .A2(new_n4659_), .B(new_n4663_), .ZN(new_n4664_));
  OAI21_X1   g04395(.A1(new_n4552_), .A2(new_n4553_), .B(new_n4664_), .ZN(new_n4665_));
  OAI21_X1   g04396(.A1(new_n4387_), .A2(new_n4391_), .B(new_n4551_), .ZN(new_n4666_));
  NAND2_X1   g04397(.A1(new_n4666_), .A2(new_n4138_), .ZN(new_n4667_));
  NOR3_X1    g04398(.A1(new_n4387_), .A2(new_n4391_), .A3(new_n4551_), .ZN(new_n4668_));
  NOR2_X1    g04399(.A1(new_n4668_), .A2(new_n4147_), .ZN(new_n4669_));
  AOI21_X1   g04400(.A1(new_n4658_), .A2(new_n4657_), .B(new_n4379_), .ZN(new_n4670_));
  NOR3_X1    g04401(.A1(new_n4644_), .A2(new_n4655_), .A3(new_n4371_), .ZN(new_n4671_));
  INV_X1     g04402(.I(new_n4663_), .ZN(new_n4672_));
  OAI21_X1   g04403(.A1(new_n4671_), .A2(new_n4670_), .B(new_n4672_), .ZN(new_n4673_));
  NAND3_X1   g04404(.A1(new_n4667_), .A2(new_n4669_), .A3(new_n4673_), .ZN(new_n4674_));
  AOI21_X1   g04405(.A1(new_n4674_), .A2(new_n4665_), .B(new_n4550_), .ZN(new_n4675_));
  INV_X1     g04406(.I(new_n4550_), .ZN(new_n4676_));
  AOI21_X1   g04407(.A1(new_n4669_), .A2(new_n4667_), .B(new_n4673_), .ZN(new_n4677_));
  NOR3_X1    g04408(.A1(new_n4552_), .A2(new_n4553_), .A3(new_n4664_), .ZN(new_n4678_));
  NOR3_X1    g04409(.A1(new_n4677_), .A2(new_n4678_), .A3(new_n4676_), .ZN(new_n4679_));
  OAI22_X1   g04410(.A1(new_n1347_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n1344_), .ZN(new_n4680_));
  OAI21_X1   g04411(.A1(new_n1109_), .A2(new_n1457_), .B(new_n4680_), .ZN(new_n4681_));
  AOI21_X1   g04412(.A1(new_n4681_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n4682_));
  XOR2_X1    g04413(.A1(new_n1299_), .A2(new_n4682_), .Z(new_n4683_));
  INV_X1     g04414(.I(new_n4683_), .ZN(new_n4684_));
  OAI21_X1   g04415(.A1(new_n4675_), .A2(new_n4679_), .B(new_n4684_), .ZN(new_n4685_));
  NOR2_X1    g04416(.A1(new_n4549_), .A2(new_n4685_), .ZN(new_n4686_));
  OAI21_X1   g04417(.A1(new_n4419_), .A2(new_n4422_), .B(new_n4160_), .ZN(new_n4687_));
  NAND2_X1   g04418(.A1(new_n4687_), .A2(new_n4167_), .ZN(new_n4688_));
  NAND3_X1   g04419(.A1(new_n4688_), .A2(new_n4175_), .A3(new_n4547_), .ZN(new_n4689_));
  OAI21_X1   g04420(.A1(new_n4677_), .A2(new_n4678_), .B(new_n4676_), .ZN(new_n4690_));
  NAND3_X1   g04421(.A1(new_n4674_), .A2(new_n4665_), .A3(new_n4550_), .ZN(new_n4691_));
  AOI21_X1   g04422(.A1(new_n4690_), .A2(new_n4691_), .B(new_n4683_), .ZN(new_n4692_));
  NOR2_X1    g04423(.A1(new_n4692_), .A2(new_n4689_), .ZN(new_n4693_));
  OAI21_X1   g04424(.A1(new_n4686_), .A2(new_n4693_), .B(new_n4545_), .ZN(new_n4694_));
  NAND2_X1   g04425(.A1(new_n4692_), .A2(new_n4689_), .ZN(new_n4695_));
  NAND2_X1   g04426(.A1(new_n4549_), .A2(new_n4685_), .ZN(new_n4696_));
  NAND3_X1   g04427(.A1(new_n4696_), .A2(new_n4695_), .A3(new_n4544_), .ZN(new_n4697_));
  NAND2_X1   g04428(.A1(new_n4694_), .A2(new_n4697_), .ZN(new_n4698_));
  OAI22_X1   g04429(.A1(new_n1055_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n1061_), .ZN(new_n4699_));
  OAI21_X1   g04430(.A1(new_n1518_), .A2(new_n1332_), .B(new_n4699_), .ZN(new_n4700_));
  AOI21_X1   g04431(.A1(new_n4700_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n4701_));
  XNOR2_X1   g04432(.A1(new_n1638_), .A2(new_n4701_), .ZN(new_n4702_));
  INV_X1     g04433(.I(new_n4702_), .ZN(new_n4703_));
  NAND3_X1   g04434(.A1(new_n4541_), .A2(new_n4698_), .A3(new_n4703_), .ZN(new_n4704_));
  NAND2_X1   g04435(.A1(new_n4170_), .A2(new_n4175_), .ZN(new_n4705_));
  NAND2_X1   g04436(.A1(new_n4186_), .A2(new_n4169_), .ZN(new_n4706_));
  AOI21_X1   g04437(.A1(new_n4705_), .A2(new_n4706_), .B(new_n4180_), .ZN(new_n4707_));
  AOI21_X1   g04438(.A1(new_n4537_), .A2(new_n4538_), .B(new_n4300_), .ZN(new_n4708_));
  NOR3_X1    g04439(.A1(new_n4428_), .A2(new_n4415_), .A3(new_n4449_), .ZN(new_n4709_));
  OAI21_X1   g04440(.A1(new_n4709_), .A2(new_n4708_), .B(new_n4707_), .ZN(new_n4710_));
  AOI21_X1   g04441(.A1(new_n4710_), .A2(new_n4192_), .B(new_n4034_), .ZN(new_n4711_));
  AOI21_X1   g04442(.A1(new_n4696_), .A2(new_n4695_), .B(new_n4544_), .ZN(new_n4712_));
  NOR3_X1    g04443(.A1(new_n4686_), .A2(new_n4693_), .A3(new_n4545_), .ZN(new_n4713_));
  OAI21_X1   g04444(.A1(new_n4713_), .A2(new_n4712_), .B(new_n4703_), .ZN(new_n4714_));
  NAND2_X1   g04445(.A1(new_n4711_), .A2(new_n4714_), .ZN(new_n4715_));
  NAND2_X1   g04446(.A1(new_n4704_), .A2(new_n4715_), .ZN(new_n4716_));
  NAND2_X1   g04447(.A1(new_n4716_), .A2(new_n4535_), .ZN(new_n4717_));
  INV_X1     g04448(.I(new_n4535_), .ZN(new_n4718_));
  NAND3_X1   g04449(.A1(new_n4704_), .A2(new_n4715_), .A3(new_n4718_), .ZN(new_n4719_));
  NAND2_X1   g04450(.A1(new_n4717_), .A2(new_n4719_), .ZN(new_n4720_));
  OAI22_X1   g04451(.A1(new_n970_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n820_), .ZN(new_n4721_));
  OAI21_X1   g04452(.A1(new_n1803_), .A2(new_n894_), .B(new_n4721_), .ZN(new_n4722_));
  AOI21_X1   g04453(.A1(new_n4722_), .A2(new_n827_), .B(new_n970_), .ZN(new_n4723_));
  XOR2_X1    g04454(.A1(new_n2106_), .A2(new_n4723_), .Z(new_n4724_));
  INV_X1     g04455(.I(new_n4724_), .ZN(new_n4725_));
  NAND2_X1   g04456(.A1(new_n4720_), .A2(new_n4725_), .ZN(new_n4726_));
  NOR2_X1    g04457(.A1(new_n4534_), .A2(new_n4726_), .ZN(new_n4727_));
  AOI21_X1   g04458(.A1(new_n4448_), .A2(new_n4452_), .B(new_n4296_), .ZN(new_n4728_));
  OAI21_X1   g04459(.A1(new_n4728_), .A2(new_n4293_), .B(new_n4028_), .ZN(new_n4729_));
  INV_X1     g04460(.I(new_n4726_), .ZN(new_n4730_));
  NOR2_X1    g04461(.A1(new_n4730_), .A2(new_n4729_), .ZN(new_n4731_));
  OAI21_X1   g04462(.A1(new_n4727_), .A2(new_n4731_), .B(new_n4532_), .ZN(new_n4732_));
  INV_X1     g04463(.I(new_n4732_), .ZN(new_n4733_));
  NOR3_X1    g04464(.A1(new_n4727_), .A2(new_n4731_), .A3(new_n4532_), .ZN(new_n4734_));
  NOR2_X1    g04465(.A1(new_n4733_), .A2(new_n4734_), .ZN(new_n4735_));
  OAI22_X1   g04466(.A1(new_n607_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n610_), .ZN(new_n4736_));
  OAI21_X1   g04467(.A1(new_n2281_), .A2(new_n684_), .B(new_n4736_), .ZN(new_n4737_));
  AOI21_X1   g04468(.A1(new_n4737_), .A2(new_n612_), .B(new_n607_), .ZN(new_n4738_));
  XNOR2_X1   g04469(.A1(new_n2647_), .A2(new_n4738_), .ZN(new_n4739_));
  NOR3_X1    g04470(.A1(new_n4525_), .A2(new_n4735_), .A3(new_n4739_), .ZN(new_n4740_));
  NAND3_X1   g04471(.A1(new_n4023_), .A2(new_n4523_), .A3(new_n4524_), .ZN(new_n4741_));
  INV_X1     g04472(.I(new_n4734_), .ZN(new_n4742_));
  NAND2_X1   g04473(.A1(new_n4742_), .A2(new_n4732_), .ZN(new_n4743_));
  INV_X1     g04474(.I(new_n4739_), .ZN(new_n4744_));
  AOI21_X1   g04475(.A1(new_n4743_), .A2(new_n4744_), .B(new_n4741_), .ZN(new_n4745_));
  NOR2_X1    g04476(.A1(new_n4740_), .A2(new_n4745_), .ZN(new_n4746_));
  NOR2_X1    g04477(.A1(new_n4746_), .A2(new_n4522_), .ZN(new_n4747_));
  INV_X1     g04478(.I(new_n4522_), .ZN(new_n4748_));
  NOR3_X1    g04479(.A1(new_n4740_), .A2(new_n4748_), .A3(new_n4745_), .ZN(new_n4749_));
  NOR2_X1    g04480(.A1(new_n4747_), .A2(new_n4749_), .ZN(new_n4750_));
  OAI22_X1   g04481(.A1(new_n448_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n450_), .ZN(new_n4751_));
  OAI21_X1   g04482(.A1(new_n2842_), .A2(new_n496_), .B(new_n4751_), .ZN(new_n4752_));
  AOI21_X1   g04483(.A1(new_n4752_), .A2(new_n452_), .B(new_n448_), .ZN(new_n4753_));
  XNOR2_X1   g04484(.A1(new_n3264_), .A2(new_n4753_), .ZN(new_n4754_));
  XOR2_X1    g04485(.A1(new_n4750_), .A2(new_n4754_), .Z(new_n4755_));
  OAI22_X1   g04486(.A1(new_n3717_), .A2(new_n341_), .B1(new_n404_), .B2(new_n3989_), .ZN(new_n4756_));
  OAI21_X1   g04487(.A1(new_n3709_), .A2(new_n366_), .B(new_n4756_), .ZN(new_n4757_));
  AOI21_X1   g04488(.A1(new_n4757_), .A2(new_n334_), .B(new_n341_), .ZN(new_n4758_));
  XNOR2_X1   g04489(.A1(new_n3993_), .A2(new_n4758_), .ZN(new_n4759_));
  INV_X1     g04490(.I(new_n4759_), .ZN(new_n4760_));
  XOR2_X1    g04491(.A1(new_n4755_), .A2(new_n4760_), .Z(new_n4761_));
  NOR2_X1    g04492(.A1(new_n4761_), .A2(new_n4521_), .ZN(new_n4762_));
  INV_X1     g04493(.I(new_n4521_), .ZN(new_n4763_));
  XOR2_X1    g04494(.A1(new_n4755_), .A2(new_n4759_), .Z(new_n4764_));
  NOR2_X1    g04495(.A1(new_n4764_), .A2(new_n4763_), .ZN(new_n4765_));
  NOR2_X1    g04496(.A1(new_n4762_), .A2(new_n4765_), .ZN(new_n4766_));
  NOR2_X1    g04497(.A1(\b[34] ), .A2(\b[35] ), .ZN(new_n4767_));
  AOI21_X1   g04498(.A1(new_n4251_), .A2(new_n4767_), .B(new_n3989_), .ZN(new_n4768_));
  NOR2_X1    g04499(.A1(new_n4253_), .A2(new_n4500_), .ZN(new_n4769_));
  INV_X1     g04500(.I(new_n4769_), .ZN(new_n4770_));
  NOR2_X1    g04501(.A1(new_n4251_), .A2(new_n4770_), .ZN(new_n4771_));
  NOR2_X1    g04502(.A1(new_n4768_), .A2(new_n4771_), .ZN(new_n4772_));
  XNOR2_X1   g04503(.A1(\b[35] ), .A2(\b[36] ), .ZN(new_n4773_));
  INV_X1     g04504(.I(\b[36] ), .ZN(new_n4774_));
  NOR2_X1    g04505(.A1(new_n4500_), .A2(new_n4774_), .ZN(new_n4775_));
  NOR2_X1    g04506(.A1(\b[35] ), .A2(\b[36] ), .ZN(new_n4776_));
  OAI21_X1   g04507(.A1(new_n4775_), .A2(new_n4776_), .B(new_n4772_), .ZN(new_n4777_));
  OAI21_X1   g04508(.A1(new_n4772_), .A2(new_n4773_), .B(new_n4777_), .ZN(new_n4778_));
  OAI22_X1   g04509(.A1(new_n330_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n263_), .ZN(new_n4779_));
  OAI21_X1   g04510(.A1(new_n4253_), .A2(new_n289_), .B(new_n4779_), .ZN(new_n4780_));
  AOI21_X1   g04511(.A1(new_n4780_), .A2(new_n260_), .B(new_n426_), .ZN(new_n4781_));
  XNOR2_X1   g04512(.A1(new_n4778_), .A2(new_n4781_), .ZN(new_n4782_));
  XOR2_X1    g04513(.A1(new_n4766_), .A2(new_n4782_), .Z(new_n4783_));
  NAND2_X1   g04514(.A1(new_n4783_), .A2(new_n4514_), .ZN(new_n4784_));
  INV_X1     g04515(.I(new_n4514_), .ZN(new_n4785_));
  INV_X1     g04516(.I(new_n4782_), .ZN(new_n4786_));
  XOR2_X1    g04517(.A1(new_n4766_), .A2(new_n4786_), .Z(new_n4787_));
  NAND2_X1   g04518(.A1(new_n4787_), .A2(new_n4785_), .ZN(new_n4788_));
  AOI21_X1   g04519(.A1(new_n4784_), .A2(new_n4788_), .B(new_n4505_), .ZN(new_n4789_));
  XOR2_X1    g04520(.A1(new_n4789_), .A2(new_n4510_), .Z(new_n4790_));
  XOR2_X1    g04521(.A1(new_n4790_), .A2(new_n4269_), .Z(\f[36] ));
  NAND2_X1   g04522(.A1(new_n4788_), .A2(new_n4784_), .ZN(new_n4792_));
  AOI21_X1   g04523(.A1(new_n4792_), .A2(new_n4509_), .B(new_n4496_), .ZN(new_n4793_));
  OAI22_X1   g04524(.A1(new_n4268_), .A2(new_n4265_), .B1(new_n4509_), .B2(new_n4792_), .ZN(new_n4794_));
  NOR2_X1    g04525(.A1(new_n4794_), .A2(new_n4793_), .ZN(new_n4795_));
  XOR2_X1    g04526(.A1(new_n4514_), .A2(new_n4766_), .Z(new_n4796_));
  NAND2_X1   g04527(.A1(new_n4796_), .A2(new_n4782_), .ZN(new_n4797_));
  XOR2_X1    g04528(.A1(new_n4755_), .A2(new_n4763_), .Z(new_n4798_));
  NOR2_X1    g04529(.A1(new_n4798_), .A2(new_n4759_), .ZN(new_n4799_));
  OAI21_X1   g04530(.A1(new_n4747_), .A2(new_n4749_), .B(new_n4519_), .ZN(new_n4800_));
  NOR3_X1    g04531(.A1(new_n4747_), .A2(new_n4519_), .A3(new_n4749_), .ZN(new_n4801_));
  INV_X1     g04532(.I(new_n4754_), .ZN(new_n4802_));
  NAND4_X1   g04533(.A1(new_n4515_), .A2(new_n4231_), .A3(new_n4516_), .A4(new_n4802_), .ZN(new_n4803_));
  OAI21_X1   g04534(.A1(new_n4803_), .A2(new_n4801_), .B(new_n4800_), .ZN(new_n4804_));
  INV_X1     g04535(.I(new_n4804_), .ZN(new_n4805_));
  AOI21_X1   g04536(.A1(new_n4735_), .A2(new_n4748_), .B(new_n4739_), .ZN(new_n4806_));
  AOI22_X1   g04537(.A1(new_n4525_), .A2(new_n4806_), .B1(new_n4522_), .B2(new_n4743_), .ZN(new_n4807_));
  AOI21_X1   g04538(.A1(new_n4529_), .A2(new_n4530_), .B(new_n4439_), .ZN(new_n4808_));
  NAND2_X1   g04539(.A1(new_n4720_), .A2(new_n4808_), .ZN(new_n4809_));
  OAI21_X1   g04540(.A1(new_n4720_), .A2(new_n4808_), .B(new_n4725_), .ZN(new_n4810_));
  OAI21_X1   g04541(.A1(new_n4729_), .A2(new_n4810_), .B(new_n4809_), .ZN(new_n4811_));
  AOI21_X1   g04542(.A1(new_n4694_), .A2(new_n4697_), .B(new_n4535_), .ZN(new_n4812_));
  NOR3_X1    g04543(.A1(new_n4713_), .A2(new_n4712_), .A3(new_n4718_), .ZN(new_n4813_));
  NOR3_X1    g04544(.A1(new_n4541_), .A2(new_n4813_), .A3(new_n4702_), .ZN(new_n4814_));
  NOR2_X1    g04545(.A1(new_n4814_), .A2(new_n4812_), .ZN(new_n4815_));
  AOI21_X1   g04546(.A1(new_n4690_), .A2(new_n4691_), .B(new_n4545_), .ZN(new_n4816_));
  INV_X1     g04547(.I(new_n4816_), .ZN(new_n4817_));
  NAND3_X1   g04548(.A1(new_n4690_), .A2(new_n4691_), .A3(new_n4545_), .ZN(new_n4818_));
  NAND3_X1   g04549(.A1(new_n4549_), .A2(new_n4818_), .A3(new_n4684_), .ZN(new_n4819_));
  NAND2_X1   g04550(.A1(new_n4819_), .A2(new_n4817_), .ZN(new_n4820_));
  NAND2_X1   g04551(.A1(new_n4669_), .A2(new_n4667_), .ZN(new_n4821_));
  NOR2_X1    g04552(.A1(new_n4671_), .A2(new_n4670_), .ZN(new_n4822_));
  NAND3_X1   g04553(.A1(new_n4656_), .A2(new_n4659_), .A3(new_n4676_), .ZN(new_n4823_));
  NAND2_X1   g04554(.A1(new_n4823_), .A2(new_n4672_), .ZN(new_n4824_));
  OAI22_X1   g04555(.A1(new_n4821_), .A2(new_n4824_), .B1(new_n4676_), .B2(new_n4822_), .ZN(new_n4825_));
  OAI21_X1   g04556(.A1(new_n4637_), .A2(new_n4635_), .B(new_n4379_), .ZN(new_n4826_));
  NAND3_X1   g04557(.A1(new_n4653_), .A2(new_n4371_), .A3(new_n4636_), .ZN(new_n4827_));
  NAND2_X1   g04558(.A1(new_n4827_), .A2(new_n4642_), .ZN(new_n4828_));
  OAI21_X1   g04559(.A1(new_n4828_), .A2(new_n4647_), .B(new_n4826_), .ZN(new_n4829_));
  NAND2_X1   g04560(.A1(new_n4619_), .A2(new_n4623_), .ZN(new_n4830_));
  NAND2_X1   g04561(.A1(new_n4830_), .A2(new_n4563_), .ZN(new_n4831_));
  INV_X1     g04562(.I(new_n4831_), .ZN(new_n4832_));
  INV_X1     g04563(.I(new_n4627_), .ZN(new_n4833_));
  NAND3_X1   g04564(.A1(new_n4650_), .A2(new_n4619_), .A3(new_n4623_), .ZN(new_n4834_));
  NAND2_X1   g04565(.A1(new_n4834_), .A2(new_n4833_), .ZN(new_n4835_));
  NOR3_X1    g04566(.A1(new_n4835_), .A2(new_n4565_), .A3(new_n4564_), .ZN(new_n4836_));
  AOI21_X1   g04567(.A1(new_n4596_), .A2(new_n4597_), .B(new_n4595_), .ZN(new_n4837_));
  NOR3_X1    g04568(.A1(new_n4593_), .A2(new_n4587_), .A3(new_n4567_), .ZN(new_n4838_));
  NOR2_X1    g04569(.A1(new_n4583_), .A2(new_n4588_), .ZN(new_n4839_));
  NOR2_X1    g04570(.A1(new_n4591_), .A2(new_n4572_), .ZN(new_n4840_));
  OAI21_X1   g04571(.A1(new_n4840_), .A2(new_n4839_), .B(new_n4567_), .ZN(new_n4841_));
  NAND2_X1   g04572(.A1(new_n4591_), .A2(new_n4572_), .ZN(new_n4842_));
  NAND2_X1   g04573(.A1(new_n4583_), .A2(new_n4588_), .ZN(new_n4843_));
  NAND3_X1   g04574(.A1(new_n4842_), .A2(new_n4843_), .A3(new_n4595_), .ZN(new_n4844_));
  AOI22_X1   g04575(.A1(new_n4841_), .A2(new_n4844_), .B1(new_n4584_), .B2(new_n4585_), .ZN(new_n4845_));
  OAI21_X1   g04576(.A1(new_n4837_), .A2(new_n4838_), .B(new_n4845_), .ZN(new_n4846_));
  NAND2_X1   g04577(.A1(new_n4846_), .A2(new_n4620_), .ZN(new_n4847_));
  NOR2_X1    g04578(.A1(new_n4588_), .A2(new_n4324_), .ZN(new_n4848_));
  NAND2_X1   g04579(.A1(new_n4588_), .A2(new_n4324_), .ZN(new_n4849_));
  NOR2_X1    g04580(.A1(new_n4313_), .A2(new_n4567_), .ZN(new_n4850_));
  AOI21_X1   g04581(.A1(new_n4849_), .A2(new_n4850_), .B(new_n4848_), .ZN(new_n4851_));
  OAI22_X1   g04582(.A1(new_n298_), .A2(new_n4072_), .B1(new_n4067_), .B2(new_n325_), .ZN(new_n4852_));
  OAI21_X1   g04583(.A1(new_n280_), .A2(new_n4318_), .B(new_n4852_), .ZN(new_n4853_));
  AOI21_X1   g04584(.A1(new_n4853_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n4854_));
  XOR2_X1    g04585(.A1(new_n4854_), .A2(new_n807_), .Z(new_n4855_));
  INV_X1     g04586(.I(new_n4855_), .ZN(new_n4856_));
  XNOR2_X1   g04587(.A1(\a[36] ), .A2(\a[38] ), .ZN(new_n4857_));
  XNOR2_X1   g04588(.A1(\a[35] ), .A2(\a[37] ), .ZN(new_n4858_));
  NOR2_X1    g04589(.A1(new_n4858_), .A2(new_n4857_), .ZN(new_n4859_));
  INV_X1     g04590(.I(\a[38] ), .ZN(new_n4860_));
  INV_X1     g04591(.I(\a[37] ), .ZN(new_n4861_));
  NOR3_X1    g04592(.A1(new_n4861_), .A2(\a[35] ), .A3(\a[36] ), .ZN(new_n4862_));
  INV_X1     g04593(.I(new_n4862_), .ZN(new_n4863_));
  NAND3_X1   g04594(.A1(new_n4861_), .A2(\a[35] ), .A3(\a[36] ), .ZN(new_n4864_));
  NAND2_X1   g04595(.A1(new_n4863_), .A2(new_n4864_), .ZN(new_n4865_));
  NAND2_X1   g04596(.A1(new_n4865_), .A2(\b[1] ), .ZN(new_n4866_));
  NAND2_X1   g04597(.A1(new_n4859_), .A2(\b[0] ), .ZN(new_n4867_));
  NAND3_X1   g04598(.A1(new_n4867_), .A2(new_n4866_), .A3(new_n4860_), .ZN(new_n4868_));
  NAND3_X1   g04599(.A1(new_n4868_), .A2(new_n444_), .A3(new_n4859_), .ZN(new_n4869_));
  AOI21_X1   g04600(.A1(new_n4868_), .A2(new_n4859_), .B(new_n444_), .ZN(new_n4870_));
  INV_X1     g04601(.I(new_n4870_), .ZN(new_n4871_));
  NAND2_X1   g04602(.A1(new_n4871_), .A2(new_n4869_), .ZN(new_n4872_));
  NOR2_X1    g04603(.A1(new_n4595_), .A2(new_n4860_), .ZN(new_n4873_));
  INV_X1     g04604(.I(new_n4873_), .ZN(new_n4874_));
  XOR2_X1    g04605(.A1(new_n4872_), .A2(new_n4874_), .Z(new_n4875_));
  NAND2_X1   g04606(.A1(new_n4875_), .A2(new_n4856_), .ZN(new_n4876_));
  XOR2_X1    g04607(.A1(new_n4872_), .A2(new_n4873_), .Z(new_n4877_));
  NAND2_X1   g04608(.A1(new_n4877_), .A2(new_n4855_), .ZN(new_n4878_));
  AOI21_X1   g04609(.A1(new_n4876_), .A2(new_n4878_), .B(new_n4851_), .ZN(new_n4879_));
  NAND2_X1   g04610(.A1(new_n4572_), .A2(new_n4574_), .ZN(new_n4880_));
  NOR2_X1    g04611(.A1(new_n4572_), .A2(new_n4574_), .ZN(new_n4881_));
  INV_X1     g04612(.I(new_n4850_), .ZN(new_n4882_));
  OAI21_X1   g04613(.A1(new_n4881_), .A2(new_n4882_), .B(new_n4880_), .ZN(new_n4883_));
  NAND2_X1   g04614(.A1(new_n4875_), .A2(new_n4855_), .ZN(new_n4884_));
  NAND2_X1   g04615(.A1(new_n4877_), .A2(new_n4856_), .ZN(new_n4885_));
  AOI21_X1   g04616(.A1(new_n4884_), .A2(new_n4885_), .B(new_n4883_), .ZN(new_n4886_));
  AOI22_X1   g04617(.A1(new_n3346_), .A2(\b[6] ), .B1(\b[7] ), .B2(new_n3351_), .ZN(new_n4887_));
  AOI21_X1   g04618(.A1(\b[5] ), .A2(new_n4331_), .B(new_n4887_), .ZN(new_n4888_));
  OAI21_X1   g04619(.A1(new_n4888_), .A2(\a[32] ), .B(new_n3346_), .ZN(new_n4889_));
  XNOR2_X1   g04620(.A1(new_n471_), .A2(new_n4889_), .ZN(new_n4890_));
  INV_X1     g04621(.I(new_n4890_), .ZN(new_n4891_));
  OAI21_X1   g04622(.A1(new_n4879_), .A2(new_n4886_), .B(new_n4891_), .ZN(new_n4892_));
  NOR2_X1    g04623(.A1(new_n4877_), .A2(new_n4855_), .ZN(new_n4893_));
  NOR2_X1    g04624(.A1(new_n4875_), .A2(new_n4856_), .ZN(new_n4894_));
  OAI21_X1   g04625(.A1(new_n4893_), .A2(new_n4894_), .B(new_n4883_), .ZN(new_n4895_));
  NOR2_X1    g04626(.A1(new_n4877_), .A2(new_n4856_), .ZN(new_n4896_));
  NOR2_X1    g04627(.A1(new_n4875_), .A2(new_n4855_), .ZN(new_n4897_));
  OAI21_X1   g04628(.A1(new_n4896_), .A2(new_n4897_), .B(new_n4851_), .ZN(new_n4898_));
  NAND3_X1   g04629(.A1(new_n4898_), .A2(new_n4895_), .A3(new_n4890_), .ZN(new_n4899_));
  NAND2_X1   g04630(.A1(new_n4892_), .A2(new_n4899_), .ZN(new_n4900_));
  NAND3_X1   g04631(.A1(new_n4847_), .A2(new_n4618_), .A3(new_n4900_), .ZN(new_n4901_));
  AOI21_X1   g04632(.A1(new_n4599_), .A2(new_n4845_), .B(new_n4601_), .ZN(new_n4902_));
  NAND3_X1   g04633(.A1(new_n4898_), .A2(new_n4895_), .A3(new_n4891_), .ZN(new_n4903_));
  OAI21_X1   g04634(.A1(new_n4879_), .A2(new_n4886_), .B(new_n4890_), .ZN(new_n4904_));
  NAND2_X1   g04635(.A1(new_n4904_), .A2(new_n4903_), .ZN(new_n4905_));
  OAI21_X1   g04636(.A1(new_n4622_), .A2(new_n4902_), .B(new_n4905_), .ZN(new_n4906_));
  NAND2_X1   g04637(.A1(new_n4906_), .A2(new_n4901_), .ZN(new_n4907_));
  OAI22_X1   g04638(.A1(new_n565_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n656_), .ZN(new_n4908_));
  OAI21_X1   g04639(.A1(new_n515_), .A2(new_n2884_), .B(new_n4908_), .ZN(new_n4909_));
  AOI21_X1   g04640(.A1(new_n4909_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n4910_));
  XNOR2_X1   g04641(.A1(new_n660_), .A2(new_n4910_), .ZN(new_n4911_));
  INV_X1     g04642(.I(new_n4911_), .ZN(new_n4912_));
  NAND2_X1   g04643(.A1(new_n4907_), .A2(new_n4912_), .ZN(new_n4913_));
  AOI21_X1   g04644(.A1(new_n4898_), .A2(new_n4895_), .B(new_n4890_), .ZN(new_n4914_));
  NOR3_X1    g04645(.A1(new_n4879_), .A2(new_n4886_), .A3(new_n4891_), .ZN(new_n4915_));
  NOR2_X1    g04646(.A1(new_n4914_), .A2(new_n4915_), .ZN(new_n4916_));
  NOR3_X1    g04647(.A1(new_n4916_), .A2(new_n4622_), .A3(new_n4902_), .ZN(new_n4917_));
  NOR3_X1    g04648(.A1(new_n4879_), .A2(new_n4886_), .A3(new_n4890_), .ZN(new_n4918_));
  AOI21_X1   g04649(.A1(new_n4898_), .A2(new_n4895_), .B(new_n4891_), .ZN(new_n4919_));
  NOR2_X1    g04650(.A1(new_n4919_), .A2(new_n4918_), .ZN(new_n4920_));
  AOI21_X1   g04651(.A1(new_n4847_), .A2(new_n4618_), .B(new_n4920_), .ZN(new_n4921_));
  NOR2_X1    g04652(.A1(new_n4921_), .A2(new_n4917_), .ZN(new_n4922_));
  NAND2_X1   g04653(.A1(new_n4922_), .A2(new_n4911_), .ZN(new_n4923_));
  NAND2_X1   g04654(.A1(new_n4913_), .A2(new_n4923_), .ZN(new_n4924_));
  OAI21_X1   g04655(.A1(new_n4836_), .A2(new_n4832_), .B(new_n4924_), .ZN(new_n4925_));
  NAND4_X1   g04656(.A1(new_n4632_), .A2(new_n4630_), .A3(new_n4834_), .A4(new_n4833_), .ZN(new_n4926_));
  NAND3_X1   g04657(.A1(new_n4906_), .A2(new_n4901_), .A3(new_n4912_), .ZN(new_n4927_));
  OAI21_X1   g04658(.A1(new_n4921_), .A2(new_n4917_), .B(new_n4911_), .ZN(new_n4928_));
  NAND2_X1   g04659(.A1(new_n4928_), .A2(new_n4927_), .ZN(new_n4929_));
  NAND3_X1   g04660(.A1(new_n4926_), .A2(new_n4831_), .A3(new_n4929_), .ZN(new_n4930_));
  OAI22_X1   g04661(.A1(new_n2171_), .A2(new_n780_), .B1(new_n861_), .B2(new_n2166_), .ZN(new_n4931_));
  OAI21_X1   g04662(.A1(new_n706_), .A2(new_n2322_), .B(new_n4931_), .ZN(new_n4932_));
  AOI21_X1   g04663(.A1(new_n4932_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n4933_));
  XNOR2_X1   g04664(.A1(new_n860_), .A2(new_n4933_), .ZN(new_n4934_));
  AOI21_X1   g04665(.A1(new_n4925_), .A2(new_n4930_), .B(new_n4934_), .ZN(new_n4935_));
  INV_X1     g04666(.I(new_n4935_), .ZN(new_n4936_));
  NAND3_X1   g04667(.A1(new_n4925_), .A2(new_n4930_), .A3(new_n4934_), .ZN(new_n4937_));
  NAND2_X1   g04668(.A1(new_n4936_), .A2(new_n4937_), .ZN(new_n4938_));
  OAI22_X1   g04669(.A1(new_n1712_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n1707_), .ZN(new_n4939_));
  OAI21_X1   g04670(.A1(new_n930_), .A2(new_n1850_), .B(new_n4939_), .ZN(new_n4940_));
  AOI21_X1   g04671(.A1(new_n4940_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n4941_));
  XOR2_X1    g04672(.A1(new_n1114_), .A2(new_n4941_), .Z(new_n4942_));
  NOR2_X1    g04673(.A1(new_n4938_), .A2(new_n4942_), .ZN(new_n4943_));
  INV_X1     g04674(.I(new_n4937_), .ZN(new_n4944_));
  NOR2_X1    g04675(.A1(new_n4944_), .A2(new_n4935_), .ZN(new_n4945_));
  INV_X1     g04676(.I(new_n4942_), .ZN(new_n4946_));
  NOR2_X1    g04677(.A1(new_n4945_), .A2(new_n4946_), .ZN(new_n4947_));
  OAI21_X1   g04678(.A1(new_n4947_), .A2(new_n4943_), .B(new_n4829_), .ZN(new_n4948_));
  NAND2_X1   g04679(.A1(new_n4938_), .A2(new_n4946_), .ZN(new_n4949_));
  NAND2_X1   g04680(.A1(new_n4945_), .A2(new_n4942_), .ZN(new_n4950_));
  AOI21_X1   g04681(.A1(new_n4949_), .A2(new_n4950_), .B(new_n4829_), .ZN(new_n4951_));
  INV_X1     g04682(.I(new_n4951_), .ZN(new_n4952_));
  NAND2_X1   g04683(.A1(new_n4952_), .A2(new_n4948_), .ZN(new_n4953_));
  OAI22_X1   g04684(.A1(new_n1347_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n1344_), .ZN(new_n4954_));
  OAI21_X1   g04685(.A1(new_n1189_), .A2(new_n1457_), .B(new_n4954_), .ZN(new_n4955_));
  AOI21_X1   g04686(.A1(new_n4955_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n4956_));
  XNOR2_X1   g04687(.A1(new_n1421_), .A2(new_n4956_), .ZN(new_n4957_));
  INV_X1     g04688(.I(new_n4957_), .ZN(new_n4958_));
  NAND2_X1   g04689(.A1(new_n4953_), .A2(new_n4958_), .ZN(new_n4959_));
  INV_X1     g04690(.I(new_n4948_), .ZN(new_n4960_));
  NOR2_X1    g04691(.A1(new_n4960_), .A2(new_n4951_), .ZN(new_n4961_));
  NAND2_X1   g04692(.A1(new_n4961_), .A2(new_n4957_), .ZN(new_n4962_));
  NAND2_X1   g04693(.A1(new_n4962_), .A2(new_n4959_), .ZN(new_n4963_));
  NAND2_X1   g04694(.A1(new_n4963_), .A2(new_n4825_), .ZN(new_n4964_));
  NOR2_X1    g04695(.A1(new_n4552_), .A2(new_n4553_), .ZN(new_n4965_));
  INV_X1     g04696(.I(new_n4822_), .ZN(new_n4966_));
  AOI21_X1   g04697(.A1(new_n4822_), .A2(new_n4676_), .B(new_n4663_), .ZN(new_n4967_));
  AOI22_X1   g04698(.A1(new_n4965_), .A2(new_n4967_), .B1(new_n4550_), .B2(new_n4966_), .ZN(new_n4968_));
  NOR3_X1    g04699(.A1(new_n4960_), .A2(new_n4951_), .A3(new_n4957_), .ZN(new_n4969_));
  AOI21_X1   g04700(.A1(new_n4952_), .A2(new_n4948_), .B(new_n4958_), .ZN(new_n4970_));
  OAI21_X1   g04701(.A1(new_n4969_), .A2(new_n4970_), .B(new_n4968_), .ZN(new_n4971_));
  OAI22_X1   g04702(.A1(new_n1055_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n1061_), .ZN(new_n4972_));
  OAI21_X1   g04703(.A1(new_n1525_), .A2(new_n1332_), .B(new_n4972_), .ZN(new_n4973_));
  AOI21_X1   g04704(.A1(new_n4973_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n4974_));
  XOR2_X1    g04705(.A1(new_n1808_), .A2(new_n4974_), .Z(new_n4975_));
  AOI21_X1   g04706(.A1(new_n4964_), .A2(new_n4971_), .B(new_n4975_), .ZN(new_n4976_));
  AOI21_X1   g04707(.A1(new_n4959_), .A2(new_n4962_), .B(new_n4968_), .ZN(new_n4977_));
  NOR2_X1    g04708(.A1(new_n4969_), .A2(new_n4970_), .ZN(new_n4978_));
  NOR2_X1    g04709(.A1(new_n4978_), .A2(new_n4825_), .ZN(new_n4979_));
  INV_X1     g04710(.I(new_n4975_), .ZN(new_n4980_));
  NOR3_X1    g04711(.A1(new_n4977_), .A2(new_n4979_), .A3(new_n4980_), .ZN(new_n4981_));
  OAI21_X1   g04712(.A1(new_n4976_), .A2(new_n4981_), .B(new_n4820_), .ZN(new_n4982_));
  NOR2_X1    g04713(.A1(new_n4689_), .A2(new_n4683_), .ZN(new_n4983_));
  AOI21_X1   g04714(.A1(new_n4983_), .A2(new_n4818_), .B(new_n4816_), .ZN(new_n4984_));
  NOR3_X1    g04715(.A1(new_n4977_), .A2(new_n4979_), .A3(new_n4975_), .ZN(new_n4985_));
  AOI21_X1   g04716(.A1(new_n4964_), .A2(new_n4971_), .B(new_n4980_), .ZN(new_n4986_));
  OAI21_X1   g04717(.A1(new_n4985_), .A2(new_n4986_), .B(new_n4984_), .ZN(new_n4987_));
  NAND2_X1   g04718(.A1(new_n4982_), .A2(new_n4987_), .ZN(new_n4988_));
  NAND2_X1   g04719(.A1(new_n4815_), .A2(new_n4988_), .ZN(new_n4989_));
  INV_X1     g04720(.I(new_n4812_), .ZN(new_n4990_));
  NAND3_X1   g04721(.A1(new_n4694_), .A2(new_n4697_), .A3(new_n4535_), .ZN(new_n4991_));
  NAND3_X1   g04722(.A1(new_n4711_), .A2(new_n4991_), .A3(new_n4703_), .ZN(new_n4992_));
  NAND2_X1   g04723(.A1(new_n4992_), .A2(new_n4990_), .ZN(new_n4993_));
  NOR2_X1    g04724(.A1(new_n4976_), .A2(new_n4981_), .ZN(new_n4994_));
  NOR2_X1    g04725(.A1(new_n4994_), .A2(new_n4984_), .ZN(new_n4995_));
  NOR2_X1    g04726(.A1(new_n4986_), .A2(new_n4985_), .ZN(new_n4996_));
  NOR2_X1    g04727(.A1(new_n4996_), .A2(new_n4820_), .ZN(new_n4997_));
  NOR2_X1    g04728(.A1(new_n4995_), .A2(new_n4997_), .ZN(new_n4998_));
  NAND2_X1   g04729(.A1(new_n4993_), .A2(new_n4998_), .ZN(new_n4999_));
  OAI22_X1   g04730(.A1(new_n970_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n820_), .ZN(new_n5000_));
  OAI21_X1   g04731(.A1(new_n1936_), .A2(new_n894_), .B(new_n5000_), .ZN(new_n5001_));
  AOI21_X1   g04732(.A1(new_n5001_), .A2(new_n827_), .B(new_n970_), .ZN(new_n5002_));
  XNOR2_X1   g04733(.A1(new_n2280_), .A2(new_n5002_), .ZN(new_n5003_));
  INV_X1     g04734(.I(new_n5003_), .ZN(new_n5004_));
  NAND3_X1   g04735(.A1(new_n4989_), .A2(new_n4999_), .A3(new_n5004_), .ZN(new_n5005_));
  NOR2_X1    g04736(.A1(new_n4993_), .A2(new_n4998_), .ZN(new_n5006_));
  INV_X1     g04737(.I(new_n4999_), .ZN(new_n5007_));
  OAI21_X1   g04738(.A1(new_n5007_), .A2(new_n5006_), .B(new_n5003_), .ZN(new_n5008_));
  NAND2_X1   g04739(.A1(new_n5008_), .A2(new_n5005_), .ZN(new_n5009_));
  NAND2_X1   g04740(.A1(new_n4811_), .A2(new_n5009_), .ZN(new_n5010_));
  INV_X1     g04741(.I(new_n4809_), .ZN(new_n5011_));
  INV_X1     g04742(.I(new_n4810_), .ZN(new_n5012_));
  AOI21_X1   g04743(.A1(new_n5012_), .A2(new_n4534_), .B(new_n5011_), .ZN(new_n5013_));
  NAND2_X1   g04744(.A1(new_n4989_), .A2(new_n4999_), .ZN(new_n5014_));
  NAND2_X1   g04745(.A1(new_n5014_), .A2(new_n5004_), .ZN(new_n5015_));
  NOR2_X1    g04746(.A1(new_n5007_), .A2(new_n5006_), .ZN(new_n5016_));
  NAND2_X1   g04747(.A1(new_n5016_), .A2(new_n5003_), .ZN(new_n5017_));
  NAND2_X1   g04748(.A1(new_n5017_), .A2(new_n5015_), .ZN(new_n5018_));
  NAND2_X1   g04749(.A1(new_n5013_), .A2(new_n5018_), .ZN(new_n5019_));
  OAI22_X1   g04750(.A1(new_n607_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n610_), .ZN(new_n5020_));
  OAI21_X1   g04751(.A1(new_n2439_), .A2(new_n684_), .B(new_n5020_), .ZN(new_n5021_));
  AOI21_X1   g04752(.A1(new_n5021_), .A2(new_n612_), .B(new_n607_), .ZN(new_n5022_));
  XNOR2_X1   g04753(.A1(new_n2846_), .A2(new_n5022_), .ZN(new_n5023_));
  INV_X1     g04754(.I(new_n5023_), .ZN(new_n5024_));
  NAND3_X1   g04755(.A1(new_n5019_), .A2(new_n5010_), .A3(new_n5024_), .ZN(new_n5025_));
  INV_X1     g04756(.I(new_n5010_), .ZN(new_n5026_));
  AOI21_X1   g04757(.A1(new_n5015_), .A2(new_n5017_), .B(new_n4811_), .ZN(new_n5027_));
  OAI21_X1   g04758(.A1(new_n5026_), .A2(new_n5027_), .B(new_n5023_), .ZN(new_n5028_));
  NAND2_X1   g04759(.A1(new_n5028_), .A2(new_n5025_), .ZN(new_n5029_));
  INV_X1     g04760(.I(new_n5029_), .ZN(new_n5030_));
  NOR2_X1    g04761(.A1(new_n4807_), .A2(new_n5030_), .ZN(new_n5031_));
  OAI21_X1   g04762(.A1(new_n4743_), .A2(new_n4522_), .B(new_n4744_), .ZN(new_n5032_));
  OAI22_X1   g04763(.A1(new_n5032_), .A2(new_n4741_), .B1(new_n4748_), .B2(new_n4735_), .ZN(new_n5033_));
  NAND2_X1   g04764(.A1(new_n5019_), .A2(new_n5010_), .ZN(new_n5034_));
  NAND2_X1   g04765(.A1(new_n5034_), .A2(new_n5024_), .ZN(new_n5035_));
  INV_X1     g04766(.I(new_n5035_), .ZN(new_n5036_));
  NOR2_X1    g04767(.A1(new_n5034_), .A2(new_n5024_), .ZN(new_n5037_));
  NOR2_X1    g04768(.A1(new_n5036_), .A2(new_n5037_), .ZN(new_n5038_));
  NOR2_X1    g04769(.A1(new_n5033_), .A2(new_n5038_), .ZN(new_n5039_));
  NOR2_X1    g04770(.A1(new_n5031_), .A2(new_n5039_), .ZN(new_n5040_));
  OAI22_X1   g04771(.A1(new_n448_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n450_), .ZN(new_n5041_));
  OAI21_X1   g04772(.A1(new_n3018_), .A2(new_n496_), .B(new_n5041_), .ZN(new_n5042_));
  AOI21_X1   g04773(.A1(new_n5042_), .A2(new_n452_), .B(new_n448_), .ZN(new_n5043_));
  XNOR2_X1   g04774(.A1(new_n3514_), .A2(new_n5043_), .ZN(new_n5044_));
  XOR2_X1    g04775(.A1(new_n5040_), .A2(new_n5044_), .Z(new_n5045_));
  OAI22_X1   g04776(.A1(new_n3989_), .A2(new_n341_), .B1(new_n404_), .B2(new_n4253_), .ZN(new_n5046_));
  OAI21_X1   g04777(.A1(new_n3717_), .A2(new_n366_), .B(new_n5046_), .ZN(new_n5047_));
  AOI21_X1   g04778(.A1(new_n5047_), .A2(new_n334_), .B(new_n341_), .ZN(new_n5048_));
  XNOR2_X1   g04779(.A1(new_n4257_), .A2(new_n5048_), .ZN(new_n5049_));
  INV_X1     g04780(.I(new_n5049_), .ZN(new_n5050_));
  NAND2_X1   g04781(.A1(new_n5045_), .A2(new_n5050_), .ZN(new_n5051_));
  INV_X1     g04782(.I(new_n5045_), .ZN(new_n5052_));
  NAND2_X1   g04783(.A1(new_n5052_), .A2(new_n5049_), .ZN(new_n5053_));
  AOI21_X1   g04784(.A1(new_n5053_), .A2(new_n5051_), .B(new_n4805_), .ZN(new_n5054_));
  NAND2_X1   g04785(.A1(new_n5052_), .A2(new_n5050_), .ZN(new_n5055_));
  NAND2_X1   g04786(.A1(new_n5045_), .A2(new_n5049_), .ZN(new_n5056_));
  AOI21_X1   g04787(.A1(new_n5055_), .A2(new_n5056_), .B(new_n4804_), .ZN(new_n5057_));
  XOR2_X1    g04788(.A1(new_n4798_), .A2(new_n4759_), .Z(new_n5058_));
  OAI21_X1   g04789(.A1(new_n5054_), .A2(new_n5057_), .B(new_n5058_), .ZN(new_n5059_));
  NOR2_X1    g04790(.A1(new_n5059_), .A2(new_n4799_), .ZN(new_n5060_));
  NOR2_X1    g04791(.A1(new_n5054_), .A2(new_n5057_), .ZN(new_n5061_));
  NOR2_X1    g04792(.A1(new_n4798_), .A2(new_n4759_), .ZN(new_n5062_));
  NOR2_X1    g04793(.A1(new_n5060_), .A2(new_n5062_), .ZN(new_n5063_));
  XOR2_X1    g04794(.A1(new_n5063_), .A2(new_n4514_), .Z(new_n5064_));
  XNOR2_X1   g04795(.A1(\b[35] ), .A2(\b[37] ), .ZN(new_n5065_));
  NOR2_X1    g04796(.A1(new_n5065_), .A2(new_n4773_), .ZN(new_n5066_));
  XOR2_X1    g04797(.A1(new_n4772_), .A2(new_n5066_), .Z(new_n5067_));
  INV_X1     g04798(.I(\b[37] ), .ZN(new_n5068_));
  OAI22_X1   g04799(.A1(new_n330_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n263_), .ZN(new_n5069_));
  OAI21_X1   g04800(.A1(new_n4500_), .A2(new_n289_), .B(new_n5069_), .ZN(new_n5070_));
  AOI21_X1   g04801(.A1(new_n5070_), .A2(new_n260_), .B(new_n426_), .ZN(new_n5071_));
  XOR2_X1    g04802(.A1(new_n5067_), .A2(new_n5071_), .Z(new_n5072_));
  NOR2_X1    g04803(.A1(new_n5064_), .A2(new_n5072_), .ZN(new_n5073_));
  XOR2_X1    g04804(.A1(new_n5073_), .A2(new_n4797_), .Z(new_n5074_));
  XNOR2_X1   g04805(.A1(new_n5074_), .A2(new_n4795_), .ZN(\f[37] ));
  NOR2_X1    g04806(.A1(new_n4792_), .A2(new_n4509_), .ZN(new_n5076_));
  NOR4_X1    g04807(.A1(new_n4269_), .A2(new_n4793_), .A3(new_n5076_), .A4(new_n5064_), .ZN(new_n5077_));
  OAI21_X1   g04808(.A1(new_n4794_), .A2(new_n4793_), .B(new_n5064_), .ZN(new_n5078_));
  NOR2_X1    g04809(.A1(new_n4797_), .A2(new_n5072_), .ZN(new_n5079_));
  AOI21_X1   g04810(.A1(new_n5078_), .A2(new_n5079_), .B(new_n5077_), .ZN(new_n5080_));
  INV_X1     g04811(.I(new_n5080_), .ZN(new_n5081_));
  XNOR2_X1   g04812(.A1(new_n5045_), .A2(new_n4804_), .ZN(new_n5082_));
  NAND2_X1   g04813(.A1(new_n5061_), .A2(new_n4798_), .ZN(new_n5083_));
  OAI21_X1   g04814(.A1(new_n5061_), .A2(new_n4798_), .B(new_n4759_), .ZN(new_n5084_));
  NAND3_X1   g04815(.A1(new_n4514_), .A2(new_n5083_), .A3(new_n5084_), .ZN(new_n5085_));
  INV_X1     g04816(.I(new_n5040_), .ZN(new_n5086_));
  INV_X1     g04817(.I(new_n5044_), .ZN(new_n5087_));
  NAND2_X1   g04818(.A1(new_n5086_), .A2(new_n5087_), .ZN(new_n5088_));
  OAI22_X1   g04819(.A1(new_n1055_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n1061_), .ZN(new_n5089_));
  OAI21_X1   g04820(.A1(new_n1634_), .A2(new_n1332_), .B(new_n5089_), .ZN(new_n5090_));
  AOI21_X1   g04821(.A1(new_n5090_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n5091_));
  XNOR2_X1   g04822(.A1(new_n1940_), .A2(new_n5091_), .ZN(new_n5092_));
  NOR2_X1    g04823(.A1(new_n4977_), .A2(new_n4979_), .ZN(new_n5093_));
  INV_X1     g04824(.I(new_n5093_), .ZN(new_n5094_));
  NOR2_X1    g04825(.A1(new_n4825_), .A2(new_n4961_), .ZN(new_n5095_));
  NOR2_X1    g04826(.A1(new_n4968_), .A2(new_n4953_), .ZN(new_n5096_));
  OAI21_X1   g04827(.A1(new_n5096_), .A2(new_n5095_), .B(new_n4957_), .ZN(new_n5097_));
  NAND2_X1   g04828(.A1(new_n4829_), .A2(new_n4938_), .ZN(new_n5098_));
  INV_X1     g04829(.I(new_n5098_), .ZN(new_n5099_));
  NOR2_X1    g04830(.A1(new_n4829_), .A2(new_n4938_), .ZN(new_n5100_));
  OAI21_X1   g04831(.A1(new_n5099_), .A2(new_n5100_), .B(new_n4942_), .ZN(new_n5101_));
  INV_X1     g04832(.I(new_n4829_), .ZN(new_n5102_));
  NAND2_X1   g04833(.A1(new_n4926_), .A2(new_n4831_), .ZN(new_n5103_));
  NAND2_X1   g04834(.A1(new_n4847_), .A2(new_n4618_), .ZN(new_n5104_));
  AOI21_X1   g04835(.A1(new_n4883_), .A2(new_n4884_), .B(new_n4897_), .ZN(new_n5105_));
  INV_X1     g04836(.I(new_n4864_), .ZN(new_n5106_));
  NOR2_X1    g04837(.A1(new_n5106_), .A2(new_n4862_), .ZN(new_n5107_));
  OAI21_X1   g04838(.A1(\b[1] ), .A2(new_n282_), .B(new_n4859_), .ZN(new_n5108_));
  OAI21_X1   g04839(.A1(new_n280_), .A2(new_n5107_), .B(new_n5108_), .ZN(new_n5109_));
  XOR2_X1    g04840(.A1(\a[35] ), .A2(\a[37] ), .Z(new_n5110_));
  XOR2_X1    g04841(.A1(\a[35] ), .A2(\a[38] ), .Z(new_n5111_));
  NAND3_X1   g04842(.A1(new_n5110_), .A2(new_n4566_), .A3(new_n5111_), .ZN(new_n5112_));
  NOR2_X1    g04843(.A1(new_n5112_), .A2(new_n258_), .ZN(new_n5113_));
  AOI21_X1   g04844(.A1(new_n5109_), .A2(new_n5113_), .B(new_n4860_), .ZN(new_n5114_));
  INV_X1     g04845(.I(new_n5114_), .ZN(new_n5115_));
  NAND3_X1   g04846(.A1(new_n5109_), .A2(new_n4860_), .A3(new_n5113_), .ZN(new_n5116_));
  NAND2_X1   g04847(.A1(new_n5115_), .A2(new_n5116_), .ZN(new_n5117_));
  NAND3_X1   g04848(.A1(new_n4871_), .A2(new_n4869_), .A3(new_n4873_), .ZN(new_n5118_));
  NAND2_X1   g04849(.A1(new_n378_), .A2(new_n4062_), .ZN(new_n5119_));
  OAI22_X1   g04850(.A1(new_n4072_), .A2(new_n325_), .B1(new_n419_), .B2(new_n4067_), .ZN(new_n5120_));
  NAND2_X1   g04851(.A1(new_n4319_), .A2(\b[3] ), .ZN(new_n5121_));
  AND3_X2    g04852(.A1(new_n5119_), .A2(new_n5120_), .A3(new_n5121_), .Z(new_n5122_));
  NAND2_X1   g04853(.A1(new_n5118_), .A2(new_n5122_), .ZN(new_n5123_));
  NAND3_X1   g04854(.A1(new_n5119_), .A2(new_n5120_), .A3(new_n5121_), .ZN(new_n5124_));
  NAND4_X1   g04855(.A1(new_n4871_), .A2(new_n5124_), .A3(new_n4869_), .A4(new_n4873_), .ZN(new_n5125_));
  AOI21_X1   g04856(.A1(new_n5123_), .A2(new_n5125_), .B(new_n5117_), .ZN(new_n5126_));
  INV_X1     g04857(.I(new_n5116_), .ZN(new_n5127_));
  NOR2_X1    g04858(.A1(new_n5127_), .A2(new_n5114_), .ZN(new_n5128_));
  INV_X1     g04859(.I(new_n4869_), .ZN(new_n5129_));
  NOR2_X1    g04860(.A1(new_n5129_), .A2(new_n4870_), .ZN(new_n5130_));
  AOI21_X1   g04861(.A1(new_n5130_), .A2(new_n4873_), .B(new_n5124_), .ZN(new_n5131_));
  NOR4_X1    g04862(.A1(new_n5122_), .A2(new_n5129_), .A3(new_n4870_), .A4(new_n4874_), .ZN(new_n5132_));
  NOR3_X1    g04863(.A1(new_n5131_), .A2(new_n5132_), .A3(new_n5128_), .ZN(new_n5133_));
  OAI21_X1   g04864(.A1(new_n5133_), .A2(new_n5126_), .B(new_n4069_), .ZN(new_n5134_));
  OAI21_X1   g04865(.A1(new_n5131_), .A2(new_n5132_), .B(new_n5128_), .ZN(new_n5135_));
  NAND3_X1   g04866(.A1(new_n5123_), .A2(new_n5117_), .A3(new_n5125_), .ZN(new_n5136_));
  NAND3_X1   g04867(.A1(new_n5135_), .A2(new_n5136_), .A3(\a[35] ), .ZN(new_n5137_));
  OAI22_X1   g04868(.A1(new_n472_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n515_), .ZN(new_n5138_));
  OAI21_X1   g04869(.A1(new_n420_), .A2(new_n3569_), .B(new_n5138_), .ZN(new_n5139_));
  AOI21_X1   g04870(.A1(new_n5139_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n5140_));
  INV_X1     g04871(.I(new_n5140_), .ZN(new_n5141_));
  NOR3_X1    g04872(.A1(new_n699_), .A2(new_n520_), .A3(new_n5141_), .ZN(new_n5142_));
  AOI21_X1   g04873(.A1(new_n521_), .A2(new_n514_), .B(new_n5140_), .ZN(new_n5143_));
  OR2_X2     g04874(.A1(new_n5143_), .A2(new_n5142_), .Z(new_n5144_));
  NAND3_X1   g04875(.A1(new_n5134_), .A2(new_n5144_), .A3(new_n5137_), .ZN(new_n5145_));
  AOI21_X1   g04876(.A1(new_n5135_), .A2(new_n5136_), .B(\a[35] ), .ZN(new_n5146_));
  NOR3_X1    g04877(.A1(new_n5133_), .A2(new_n5126_), .A3(new_n4069_), .ZN(new_n5147_));
  NOR2_X1    g04878(.A1(new_n5143_), .A2(new_n5142_), .ZN(new_n5148_));
  OAI21_X1   g04879(.A1(new_n5146_), .A2(new_n5147_), .B(new_n5148_), .ZN(new_n5149_));
  AOI21_X1   g04880(.A1(new_n5145_), .A2(new_n5149_), .B(new_n5105_), .ZN(new_n5150_));
  OAI21_X1   g04881(.A1(new_n4851_), .A2(new_n4896_), .B(new_n4885_), .ZN(new_n5151_));
  OAI21_X1   g04882(.A1(new_n5146_), .A2(new_n5147_), .B(new_n5144_), .ZN(new_n5152_));
  NAND3_X1   g04883(.A1(new_n5134_), .A2(new_n5137_), .A3(new_n5148_), .ZN(new_n5153_));
  AOI21_X1   g04884(.A1(new_n5152_), .A2(new_n5153_), .B(new_n5151_), .ZN(new_n5154_));
  NOR2_X1    g04885(.A1(new_n5150_), .A2(new_n5154_), .ZN(new_n5155_));
  NOR3_X1    g04886(.A1(new_n5155_), .A2(new_n4920_), .A3(new_n4914_), .ZN(new_n5156_));
  NOR2_X1    g04887(.A1(new_n4879_), .A2(new_n4886_), .ZN(new_n5157_));
  NAND2_X1   g04888(.A1(new_n5134_), .A2(new_n5137_), .ZN(new_n5158_));
  INV_X1     g04889(.I(new_n5158_), .ZN(new_n5159_));
  NOR2_X1    g04890(.A1(new_n5157_), .A2(new_n4890_), .ZN(new_n5160_));
  OAI21_X1   g04891(.A1(new_n5156_), .A2(new_n5160_), .B(new_n5104_), .ZN(new_n5161_));
  NOR2_X1    g04892(.A1(new_n4622_), .A2(new_n4902_), .ZN(new_n5162_));
  NOR3_X1    g04893(.A1(new_n5146_), .A2(new_n5147_), .A3(new_n5148_), .ZN(new_n5163_));
  AOI21_X1   g04894(.A1(new_n5134_), .A2(new_n5137_), .B(new_n5144_), .ZN(new_n5164_));
  OAI21_X1   g04895(.A1(new_n5164_), .A2(new_n5163_), .B(new_n5151_), .ZN(new_n5165_));
  AOI21_X1   g04896(.A1(new_n5134_), .A2(new_n5137_), .B(new_n5148_), .ZN(new_n5166_));
  NOR3_X1    g04897(.A1(new_n5146_), .A2(new_n5147_), .A3(new_n5144_), .ZN(new_n5167_));
  OAI21_X1   g04898(.A1(new_n5167_), .A2(new_n5166_), .B(new_n5105_), .ZN(new_n5168_));
  NAND2_X1   g04899(.A1(new_n5168_), .A2(new_n5165_), .ZN(new_n5169_));
  NAND3_X1   g04900(.A1(new_n5169_), .A2(new_n4905_), .A3(new_n4892_), .ZN(new_n5170_));
  INV_X1     g04901(.I(new_n5160_), .ZN(new_n5171_));
  NAND3_X1   g04902(.A1(new_n5170_), .A2(new_n5162_), .A3(new_n5171_), .ZN(new_n5172_));
  OAI22_X1   g04903(.A1(new_n656_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n706_), .ZN(new_n5173_));
  OAI21_X1   g04904(.A1(new_n565_), .A2(new_n2884_), .B(new_n5173_), .ZN(new_n5174_));
  AOI21_X1   g04905(.A1(new_n5174_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n5175_));
  XNOR2_X1   g04906(.A1(new_n710_), .A2(new_n5175_), .ZN(new_n5176_));
  INV_X1     g04907(.I(new_n5176_), .ZN(new_n5177_));
  NAND3_X1   g04908(.A1(new_n5161_), .A2(new_n5172_), .A3(new_n5177_), .ZN(new_n5178_));
  AOI21_X1   g04909(.A1(new_n5170_), .A2(new_n5171_), .B(new_n5162_), .ZN(new_n5179_));
  NOR3_X1    g04910(.A1(new_n5156_), .A2(new_n5104_), .A3(new_n5160_), .ZN(new_n5180_));
  OAI21_X1   g04911(.A1(new_n5180_), .A2(new_n5179_), .B(new_n5176_), .ZN(new_n5181_));
  NAND2_X1   g04912(.A1(new_n5181_), .A2(new_n5178_), .ZN(new_n5182_));
  NAND3_X1   g04913(.A1(new_n5182_), .A2(new_n4913_), .A3(new_n4929_), .ZN(new_n5183_));
  INV_X1     g04914(.I(new_n5182_), .ZN(new_n5184_));
  NOR2_X1    g04915(.A1(new_n4922_), .A2(new_n4911_), .ZN(new_n5185_));
  INV_X1     g04916(.I(new_n5185_), .ZN(new_n5186_));
  AOI21_X1   g04917(.A1(new_n5183_), .A2(new_n5186_), .B(new_n5103_), .ZN(new_n5187_));
  NOR2_X1    g04918(.A1(new_n4836_), .A2(new_n4832_), .ZN(new_n5188_));
  INV_X1     g04919(.I(new_n4913_), .ZN(new_n5189_));
  NOR3_X1    g04920(.A1(new_n5180_), .A2(new_n5179_), .A3(new_n5176_), .ZN(new_n5190_));
  AOI21_X1   g04921(.A1(new_n5161_), .A2(new_n5172_), .B(new_n5177_), .ZN(new_n5191_));
  OAI21_X1   g04922(.A1(new_n5190_), .A2(new_n5191_), .B(new_n4929_), .ZN(new_n5192_));
  NOR2_X1    g04923(.A1(new_n5192_), .A2(new_n5189_), .ZN(new_n5193_));
  NOR3_X1    g04924(.A1(new_n5193_), .A2(new_n5188_), .A3(new_n5185_), .ZN(new_n5194_));
  OAI22_X1   g04925(.A1(new_n2171_), .A2(new_n861_), .B1(new_n930_), .B2(new_n2166_), .ZN(new_n5195_));
  OAI21_X1   g04926(.A1(new_n780_), .A2(new_n2322_), .B(new_n5195_), .ZN(new_n5196_));
  AOI21_X1   g04927(.A1(new_n5196_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n5197_));
  XNOR2_X1   g04928(.A1(new_n937_), .A2(new_n5197_), .ZN(new_n5198_));
  NOR3_X1    g04929(.A1(new_n5194_), .A2(new_n5187_), .A3(new_n5198_), .ZN(new_n5199_));
  OAI21_X1   g04930(.A1(new_n5193_), .A2(new_n5185_), .B(new_n5188_), .ZN(new_n5200_));
  NAND3_X1   g04931(.A1(new_n5183_), .A2(new_n5103_), .A3(new_n5186_), .ZN(new_n5201_));
  INV_X1     g04932(.I(new_n5198_), .ZN(new_n5202_));
  AOI21_X1   g04933(.A1(new_n5200_), .A2(new_n5201_), .B(new_n5202_), .ZN(new_n5203_));
  AOI22_X1   g04934(.A1(new_n4926_), .A2(new_n4831_), .B1(new_n4913_), .B2(new_n4923_), .ZN(new_n5204_));
  INV_X1     g04935(.I(new_n4930_), .ZN(new_n5205_));
  OAI21_X1   g04936(.A1(new_n5205_), .A2(new_n5204_), .B(new_n4934_), .ZN(new_n5206_));
  INV_X1     g04937(.I(new_n4934_), .ZN(new_n5207_));
  NAND3_X1   g04938(.A1(new_n4925_), .A2(new_n4930_), .A3(new_n5207_), .ZN(new_n5208_));
  NAND2_X1   g04939(.A1(new_n5206_), .A2(new_n5208_), .ZN(new_n5209_));
  OAI21_X1   g04940(.A1(new_n5199_), .A2(new_n5203_), .B(new_n5209_), .ZN(new_n5210_));
  NOR2_X1    g04941(.A1(new_n5210_), .A2(new_n4935_), .ZN(new_n5211_));
  NAND3_X1   g04942(.A1(new_n5200_), .A2(new_n5201_), .A3(new_n5202_), .ZN(new_n5212_));
  OAI21_X1   g04943(.A1(new_n5194_), .A2(new_n5187_), .B(new_n5198_), .ZN(new_n5213_));
  NAND2_X1   g04944(.A1(new_n5213_), .A2(new_n5212_), .ZN(new_n5214_));
  AOI21_X1   g04945(.A1(new_n4925_), .A2(new_n4930_), .B(new_n4934_), .ZN(new_n5216_));
  OAI21_X1   g04946(.A1(new_n5211_), .A2(new_n5216_), .B(new_n5102_), .ZN(new_n5217_));
  NAND3_X1   g04947(.A1(new_n5214_), .A2(new_n4936_), .A3(new_n5209_), .ZN(new_n5218_));
  INV_X1     g04948(.I(new_n5216_), .ZN(new_n5219_));
  NAND3_X1   g04949(.A1(new_n5218_), .A2(new_n4829_), .A3(new_n5219_), .ZN(new_n5220_));
  OAI22_X1   g04950(.A1(new_n1712_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n1707_), .ZN(new_n5221_));
  OAI21_X1   g04951(.A1(new_n1017_), .A2(new_n1850_), .B(new_n5221_), .ZN(new_n5222_));
  AOI21_X1   g04952(.A1(new_n5222_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n5223_));
  XNOR2_X1   g04953(.A1(new_n1196_), .A2(new_n5223_), .ZN(new_n5224_));
  INV_X1     g04954(.I(new_n5224_), .ZN(new_n5225_));
  NAND3_X1   g04955(.A1(new_n5217_), .A2(new_n5220_), .A3(new_n5225_), .ZN(new_n5226_));
  AOI21_X1   g04956(.A1(new_n5218_), .A2(new_n5219_), .B(new_n4829_), .ZN(new_n5227_));
  NOR3_X1    g04957(.A1(new_n5211_), .A2(new_n5102_), .A3(new_n5216_), .ZN(new_n5228_));
  OAI21_X1   g04958(.A1(new_n5228_), .A2(new_n5227_), .B(new_n5224_), .ZN(new_n5229_));
  NAND3_X1   g04959(.A1(new_n5229_), .A2(new_n5226_), .A3(new_n5101_), .ZN(new_n5230_));
  NAND3_X1   g04960(.A1(new_n5230_), .A2(new_n4968_), .A3(new_n4953_), .ZN(new_n5231_));
  INV_X1     g04961(.I(new_n5101_), .ZN(new_n5232_));
  NOR3_X1    g04962(.A1(new_n5228_), .A2(new_n5227_), .A3(new_n5224_), .ZN(new_n5233_));
  AOI21_X1   g04963(.A1(new_n5217_), .A2(new_n5220_), .B(new_n5225_), .ZN(new_n5234_));
  NOR3_X1    g04964(.A1(new_n5233_), .A2(new_n5234_), .A3(new_n5232_), .ZN(new_n5235_));
  OAI21_X1   g04965(.A1(new_n5235_), .A2(new_n4961_), .B(new_n4825_), .ZN(new_n5236_));
  OAI22_X1   g04966(.A1(new_n1347_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n1344_), .ZN(new_n5237_));
  OAI21_X1   g04967(.A1(new_n1294_), .A2(new_n1457_), .B(new_n5237_), .ZN(new_n5238_));
  AOI21_X1   g04968(.A1(new_n5238_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n5239_));
  XOR2_X1    g04969(.A1(new_n1530_), .A2(new_n5239_), .Z(new_n5240_));
  INV_X1     g04970(.I(new_n5240_), .ZN(new_n5241_));
  NAND3_X1   g04971(.A1(new_n5236_), .A2(new_n5231_), .A3(new_n5241_), .ZN(new_n5242_));
  NOR3_X1    g04972(.A1(new_n5235_), .A2(new_n4825_), .A3(new_n4961_), .ZN(new_n5243_));
  AOI21_X1   g04973(.A1(new_n5230_), .A2(new_n4953_), .B(new_n4968_), .ZN(new_n5244_));
  OAI21_X1   g04974(.A1(new_n5243_), .A2(new_n5244_), .B(new_n5240_), .ZN(new_n5245_));
  NAND3_X1   g04975(.A1(new_n5245_), .A2(new_n5242_), .A3(new_n5097_), .ZN(new_n5246_));
  NAND3_X1   g04976(.A1(new_n5246_), .A2(new_n4984_), .A3(new_n5094_), .ZN(new_n5247_));
  NAND2_X1   g04977(.A1(new_n4968_), .A2(new_n4953_), .ZN(new_n5248_));
  NAND2_X1   g04978(.A1(new_n4825_), .A2(new_n4961_), .ZN(new_n5249_));
  AOI21_X1   g04979(.A1(new_n5248_), .A2(new_n5249_), .B(new_n4958_), .ZN(new_n5250_));
  NOR3_X1    g04980(.A1(new_n5243_), .A2(new_n5244_), .A3(new_n5240_), .ZN(new_n5251_));
  AOI21_X1   g04981(.A1(new_n5236_), .A2(new_n5231_), .B(new_n5241_), .ZN(new_n5252_));
  NOR3_X1    g04982(.A1(new_n5251_), .A2(new_n5252_), .A3(new_n5250_), .ZN(new_n5253_));
  OAI21_X1   g04983(.A1(new_n5253_), .A2(new_n5093_), .B(new_n4820_), .ZN(new_n5254_));
  NAND2_X1   g04984(.A1(new_n5254_), .A2(new_n5247_), .ZN(new_n5255_));
  NAND2_X1   g04985(.A1(new_n4984_), .A2(new_n5094_), .ZN(new_n5256_));
  NAND2_X1   g04986(.A1(new_n4820_), .A2(new_n5093_), .ZN(new_n5257_));
  AOI21_X1   g04987(.A1(new_n5257_), .A2(new_n5256_), .B(new_n4980_), .ZN(new_n5258_));
  NOR3_X1    g04988(.A1(new_n4814_), .A2(new_n4812_), .A3(new_n4988_), .ZN(new_n5259_));
  OAI22_X1   g04989(.A1(new_n970_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n820_), .ZN(new_n5260_));
  OAI21_X1   g04990(.A1(new_n2102_), .A2(new_n894_), .B(new_n5260_), .ZN(new_n5261_));
  AOI21_X1   g04991(.A1(new_n5261_), .A2(new_n827_), .B(new_n970_), .ZN(new_n5262_));
  XNOR2_X1   g04992(.A1(new_n2443_), .A2(new_n5262_), .ZN(new_n5263_));
  INV_X1     g04993(.I(new_n5263_), .ZN(new_n5264_));
  OAI21_X1   g04994(.A1(new_n5259_), .A2(new_n5258_), .B(new_n5264_), .ZN(new_n5265_));
  INV_X1     g04995(.I(new_n5258_), .ZN(new_n5266_));
  NAND3_X1   g04996(.A1(new_n4992_), .A2(new_n4998_), .A3(new_n4990_), .ZN(new_n5267_));
  NAND3_X1   g04997(.A1(new_n5267_), .A2(new_n5266_), .A3(new_n5263_), .ZN(new_n5268_));
  AOI21_X1   g04998(.A1(new_n5265_), .A2(new_n5268_), .B(new_n5255_), .ZN(new_n5269_));
  NOR3_X1    g04999(.A1(new_n5253_), .A2(new_n4820_), .A3(new_n5093_), .ZN(new_n5270_));
  AOI21_X1   g05000(.A1(new_n5246_), .A2(new_n5094_), .B(new_n4984_), .ZN(new_n5271_));
  NOR2_X1    g05001(.A1(new_n5270_), .A2(new_n5271_), .ZN(new_n5272_));
  AOI21_X1   g05002(.A1(new_n5267_), .A2(new_n5266_), .B(new_n5263_), .ZN(new_n5273_));
  NOR3_X1    g05003(.A1(new_n5259_), .A2(new_n5258_), .A3(new_n5264_), .ZN(new_n5274_));
  NOR3_X1    g05004(.A1(new_n5274_), .A2(new_n5273_), .A3(new_n5272_), .ZN(new_n5275_));
  OAI21_X1   g05005(.A1(new_n5275_), .A2(new_n5269_), .B(new_n5092_), .ZN(new_n5276_));
  INV_X1     g05006(.I(new_n5092_), .ZN(new_n5277_));
  OAI21_X1   g05007(.A1(new_n5274_), .A2(new_n5273_), .B(new_n5272_), .ZN(new_n5278_));
  NAND3_X1   g05008(.A1(new_n5265_), .A2(new_n5268_), .A3(new_n5255_), .ZN(new_n5279_));
  NAND3_X1   g05009(.A1(new_n5278_), .A2(new_n5279_), .A3(new_n5277_), .ZN(new_n5280_));
  NAND2_X1   g05010(.A1(new_n5276_), .A2(new_n5280_), .ZN(new_n5281_));
  NAND3_X1   g05011(.A1(new_n5281_), .A2(new_n5009_), .A3(new_n5015_), .ZN(new_n5282_));
  NOR2_X1    g05012(.A1(new_n5016_), .A2(new_n5003_), .ZN(new_n5284_));
  INV_X1     g05013(.I(new_n5284_), .ZN(new_n5285_));
  AOI21_X1   g05014(.A1(new_n5282_), .A2(new_n5285_), .B(new_n4811_), .ZN(new_n5286_));
  INV_X1     g05015(.I(new_n5015_), .ZN(new_n5287_));
  AOI21_X1   g05016(.A1(new_n5278_), .A2(new_n5279_), .B(new_n5277_), .ZN(new_n5288_));
  NOR3_X1    g05017(.A1(new_n5275_), .A2(new_n5269_), .A3(new_n5092_), .ZN(new_n5289_));
  OAI21_X1   g05018(.A1(new_n5289_), .A2(new_n5288_), .B(new_n5009_), .ZN(new_n5290_));
  NOR2_X1    g05019(.A1(new_n5290_), .A2(new_n5287_), .ZN(new_n5291_));
  NOR3_X1    g05020(.A1(new_n5291_), .A2(new_n5013_), .A3(new_n5284_), .ZN(new_n5292_));
  OAI22_X1   g05021(.A1(new_n607_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n610_), .ZN(new_n5293_));
  OAI21_X1   g05022(.A1(new_n2643_), .A2(new_n684_), .B(new_n5293_), .ZN(new_n5294_));
  AOI21_X1   g05023(.A1(new_n5294_), .A2(new_n612_), .B(new_n607_), .ZN(new_n5295_));
  XNOR2_X1   g05024(.A1(new_n3022_), .A2(new_n5295_), .ZN(new_n5296_));
  INV_X1     g05025(.I(new_n5296_), .ZN(new_n5297_));
  OAI21_X1   g05026(.A1(new_n5292_), .A2(new_n5286_), .B(new_n5297_), .ZN(new_n5298_));
  OAI21_X1   g05027(.A1(new_n5291_), .A2(new_n5284_), .B(new_n5013_), .ZN(new_n5299_));
  NAND3_X1   g05028(.A1(new_n5282_), .A2(new_n4811_), .A3(new_n5285_), .ZN(new_n5300_));
  NAND3_X1   g05029(.A1(new_n5299_), .A2(new_n5300_), .A3(new_n5296_), .ZN(new_n5301_));
  NAND2_X1   g05030(.A1(new_n5298_), .A2(new_n5301_), .ZN(new_n5302_));
  NAND3_X1   g05031(.A1(new_n5302_), .A2(new_n5029_), .A3(new_n5035_), .ZN(new_n5303_));
  NOR2_X1    g05032(.A1(new_n5026_), .A2(new_n5027_), .ZN(new_n5304_));
  NOR2_X1    g05033(.A1(new_n5304_), .A2(new_n5023_), .ZN(new_n5306_));
  INV_X1     g05034(.I(new_n5306_), .ZN(new_n5307_));
  AOI21_X1   g05035(.A1(new_n5303_), .A2(new_n5307_), .B(new_n5033_), .ZN(new_n5308_));
  AOI21_X1   g05036(.A1(new_n5299_), .A2(new_n5300_), .B(new_n5296_), .ZN(new_n5309_));
  NOR3_X1    g05037(.A1(new_n5292_), .A2(new_n5286_), .A3(new_n5297_), .ZN(new_n5310_));
  OAI21_X1   g05038(.A1(new_n5310_), .A2(new_n5309_), .B(new_n5029_), .ZN(new_n5311_));
  NOR2_X1    g05039(.A1(new_n5311_), .A2(new_n5036_), .ZN(new_n5312_));
  NOR3_X1    g05040(.A1(new_n5312_), .A2(new_n4807_), .A3(new_n5306_), .ZN(new_n5313_));
  OAI22_X1   g05041(.A1(new_n448_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n450_), .ZN(new_n5314_));
  OAI21_X1   g05042(.A1(new_n3260_), .A2(new_n496_), .B(new_n5314_), .ZN(new_n5315_));
  AOI21_X1   g05043(.A1(new_n5315_), .A2(new_n452_), .B(new_n448_), .ZN(new_n5316_));
  XOR2_X1    g05044(.A1(new_n3722_), .A2(new_n5316_), .Z(new_n5317_));
  INV_X1     g05045(.I(new_n5317_), .ZN(new_n5318_));
  OAI21_X1   g05046(.A1(new_n5313_), .A2(new_n5308_), .B(new_n5318_), .ZN(new_n5319_));
  OAI21_X1   g05047(.A1(new_n5312_), .A2(new_n5306_), .B(new_n4807_), .ZN(new_n5320_));
  NAND3_X1   g05048(.A1(new_n5303_), .A2(new_n5033_), .A3(new_n5307_), .ZN(new_n5321_));
  NAND3_X1   g05049(.A1(new_n5320_), .A2(new_n5321_), .A3(new_n5317_), .ZN(new_n5322_));
  NAND2_X1   g05050(.A1(new_n5319_), .A2(new_n5322_), .ZN(new_n5323_));
  XOR2_X1    g05051(.A1(new_n5040_), .A2(new_n5044_), .Z(new_n5324_));
  NAND3_X1   g05052(.A1(new_n5324_), .A2(new_n5088_), .A3(new_n5323_), .ZN(new_n5325_));
  AOI21_X1   g05053(.A1(new_n5320_), .A2(new_n5321_), .B(new_n5317_), .ZN(new_n5326_));
  NOR3_X1    g05054(.A1(new_n5313_), .A2(new_n5308_), .A3(new_n5318_), .ZN(new_n5327_));
  NAND2_X1   g05055(.A1(new_n5086_), .A2(new_n5087_), .ZN(new_n5328_));
  AOI21_X1   g05056(.A1(new_n5325_), .A2(new_n5328_), .B(new_n4804_), .ZN(new_n5329_));
  AND3_X2    g05057(.A1(new_n5325_), .A2(new_n4804_), .A3(new_n5328_), .Z(new_n5330_));
  OR2_X2     g05058(.A1(new_n5330_), .A2(new_n5329_), .Z(new_n5331_));
  OAI22_X1   g05059(.A1(new_n4253_), .A2(new_n341_), .B1(new_n404_), .B2(new_n4500_), .ZN(new_n5332_));
  OAI21_X1   g05060(.A1(new_n3989_), .A2(new_n366_), .B(new_n5332_), .ZN(new_n5333_));
  AOI21_X1   g05061(.A1(new_n5333_), .A2(new_n334_), .B(new_n341_), .ZN(new_n5334_));
  XOR2_X1    g05062(.A1(new_n4499_), .A2(new_n5334_), .Z(new_n5335_));
  INV_X1     g05063(.I(new_n5335_), .ZN(new_n5336_));
  NAND2_X1   g05064(.A1(new_n5331_), .A2(new_n5336_), .ZN(new_n5337_));
  INV_X1     g05065(.I(new_n5337_), .ZN(new_n5338_));
  AND2_X2    g05066(.A1(new_n5085_), .A2(new_n5338_), .Z(new_n5339_));
  NOR2_X1    g05067(.A1(new_n5085_), .A2(new_n5338_), .ZN(new_n5340_));
  OAI22_X1   g05068(.A1(new_n5339_), .A2(new_n5340_), .B1(new_n5050_), .B2(new_n5082_), .ZN(new_n5341_));
  NOR2_X1    g05069(.A1(new_n5082_), .A2(new_n5050_), .ZN(new_n5342_));
  NOR2_X1    g05070(.A1(new_n5339_), .A2(new_n5340_), .ZN(new_n5343_));
  NAND2_X1   g05071(.A1(new_n5343_), .A2(new_n5342_), .ZN(new_n5344_));
  NAND2_X1   g05072(.A1(new_n5344_), .A2(new_n5341_), .ZN(new_n5345_));
  NOR2_X1    g05073(.A1(\b[36] ), .A2(\b[37] ), .ZN(new_n5346_));
  AOI21_X1   g05074(.A1(new_n4772_), .A2(new_n5346_), .B(new_n4500_), .ZN(new_n5347_));
  NOR2_X1    g05075(.A1(new_n4774_), .A2(new_n5068_), .ZN(new_n5348_));
  INV_X1     g05076(.I(new_n5348_), .ZN(new_n5349_));
  NOR2_X1    g05077(.A1(new_n4772_), .A2(new_n5349_), .ZN(new_n5350_));
  NOR2_X1    g05078(.A1(new_n5347_), .A2(new_n5350_), .ZN(new_n5351_));
  XNOR2_X1   g05079(.A1(\b[37] ), .A2(\b[38] ), .ZN(new_n5352_));
  INV_X1     g05080(.I(\b[38] ), .ZN(new_n5353_));
  NOR2_X1    g05081(.A1(new_n5068_), .A2(new_n5353_), .ZN(new_n5354_));
  NOR2_X1    g05082(.A1(\b[37] ), .A2(\b[38] ), .ZN(new_n5355_));
  OAI21_X1   g05083(.A1(new_n5354_), .A2(new_n5355_), .B(new_n5351_), .ZN(new_n5356_));
  OAI21_X1   g05084(.A1(new_n5351_), .A2(new_n5352_), .B(new_n5356_), .ZN(new_n5357_));
  OAI22_X1   g05085(.A1(new_n330_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n263_), .ZN(new_n5358_));
  OAI21_X1   g05086(.A1(new_n4774_), .A2(new_n289_), .B(new_n5358_), .ZN(new_n5359_));
  AOI21_X1   g05087(.A1(new_n5359_), .A2(new_n260_), .B(new_n426_), .ZN(new_n5360_));
  XNOR2_X1   g05088(.A1(new_n5357_), .A2(new_n5360_), .ZN(new_n5361_));
  XOR2_X1    g05089(.A1(new_n5345_), .A2(new_n5361_), .Z(new_n5362_));
  NAND2_X1   g05090(.A1(new_n5081_), .A2(new_n5362_), .ZN(new_n5363_));
  XOR2_X1    g05091(.A1(new_n5345_), .A2(new_n5361_), .Z(new_n5364_));
  OAI21_X1   g05092(.A1(new_n5081_), .A2(new_n5364_), .B(new_n5363_), .ZN(\f[38] ));
  INV_X1     g05093(.I(new_n5345_), .ZN(new_n5366_));
  NOR2_X1    g05094(.A1(new_n5366_), .A2(new_n5361_), .ZN(new_n5367_));
  NAND2_X1   g05095(.A1(new_n5331_), .A2(new_n5342_), .ZN(new_n5368_));
  NOR2_X1    g05096(.A1(new_n5331_), .A2(new_n5342_), .ZN(new_n5369_));
  NAND4_X1   g05097(.A1(new_n4514_), .A2(new_n5083_), .A3(new_n5084_), .A4(new_n5336_), .ZN(new_n5370_));
  OAI21_X1   g05098(.A1(new_n5370_), .A2(new_n5369_), .B(new_n5368_), .ZN(new_n5371_));
  INV_X1     g05099(.I(new_n5371_), .ZN(new_n5372_));
  AOI21_X1   g05100(.A1(new_n5320_), .A2(new_n5321_), .B(new_n5318_), .ZN(new_n5373_));
  INV_X1     g05101(.I(new_n5373_), .ZN(new_n5374_));
  AOI21_X1   g05102(.A1(new_n5323_), .A2(new_n5086_), .B(new_n5087_), .ZN(new_n5375_));
  NAND3_X1   g05103(.A1(new_n5319_), .A2(new_n5322_), .A3(new_n5040_), .ZN(new_n5376_));
  NAND2_X1   g05104(.A1(new_n4804_), .A2(new_n5376_), .ZN(new_n5377_));
  NOR2_X1    g05105(.A1(new_n5377_), .A2(new_n5375_), .ZN(new_n5378_));
  OAI21_X1   g05106(.A1(new_n5259_), .A2(new_n5258_), .B(new_n5255_), .ZN(new_n5379_));
  NAND3_X1   g05107(.A1(new_n5267_), .A2(new_n5272_), .A3(new_n5266_), .ZN(new_n5380_));
  AOI21_X1   g05108(.A1(new_n5379_), .A2(new_n5380_), .B(new_n5277_), .ZN(new_n5381_));
  NAND3_X1   g05109(.A1(new_n5379_), .A2(new_n5380_), .A3(new_n5277_), .ZN(new_n5382_));
  INV_X1     g05110(.I(new_n5382_), .ZN(new_n5383_));
  OAI21_X1   g05111(.A1(new_n5383_), .A2(new_n5381_), .B(new_n5264_), .ZN(new_n5384_));
  AOI21_X1   g05112(.A1(new_n5281_), .A2(new_n5014_), .B(new_n5004_), .ZN(new_n5385_));
  NAND3_X1   g05113(.A1(new_n5276_), .A2(new_n5280_), .A3(new_n5016_), .ZN(new_n5386_));
  NAND2_X1   g05114(.A1(new_n5386_), .A2(new_n4811_), .ZN(new_n5387_));
  NAND2_X1   g05115(.A1(new_n5255_), .A2(new_n5092_), .ZN(new_n5388_));
  NOR2_X1    g05116(.A1(new_n5272_), .A2(new_n5092_), .ZN(new_n5389_));
  NAND3_X1   g05117(.A1(new_n5254_), .A2(new_n5247_), .A3(new_n5092_), .ZN(new_n5390_));
  INV_X1     g05118(.I(new_n5390_), .ZN(new_n5391_));
  OAI21_X1   g05119(.A1(new_n5389_), .A2(new_n5391_), .B(new_n5258_), .ZN(new_n5392_));
  AOI21_X1   g05120(.A1(new_n5392_), .A2(new_n4998_), .B(new_n4815_), .ZN(new_n5393_));
  AOI21_X1   g05121(.A1(new_n5245_), .A2(new_n5242_), .B(new_n5097_), .ZN(new_n5394_));
  OAI21_X1   g05122(.A1(new_n5394_), .A2(new_n5094_), .B(new_n4820_), .ZN(new_n5395_));
  OAI21_X1   g05123(.A1(new_n5233_), .A2(new_n5234_), .B(new_n5232_), .ZN(new_n5396_));
  AOI21_X1   g05124(.A1(new_n5396_), .A2(new_n4961_), .B(new_n4968_), .ZN(new_n5397_));
  NOR3_X1    g05125(.A1(new_n5194_), .A2(new_n5187_), .A3(new_n5202_), .ZN(new_n5398_));
  NAND2_X1   g05126(.A1(new_n4925_), .A2(new_n4930_), .ZN(new_n5399_));
  AOI21_X1   g05127(.A1(new_n5214_), .A2(new_n5399_), .B(new_n5207_), .ZN(new_n5400_));
  OAI21_X1   g05128(.A1(new_n5214_), .A2(new_n5399_), .B(new_n4829_), .ZN(new_n5401_));
  AOI21_X1   g05129(.A1(new_n5182_), .A2(new_n4907_), .B(new_n4912_), .ZN(new_n5402_));
  INV_X1     g05130(.I(new_n5402_), .ZN(new_n5403_));
  AOI21_X1   g05131(.A1(new_n4922_), .A2(new_n5184_), .B(new_n5188_), .ZN(new_n5404_));
  NAND2_X1   g05132(.A1(new_n5105_), .A2(new_n5158_), .ZN(new_n5405_));
  NAND2_X1   g05133(.A1(new_n5159_), .A2(new_n5151_), .ZN(new_n5406_));
  AOI21_X1   g05134(.A1(new_n5406_), .A2(new_n5405_), .B(new_n5144_), .ZN(new_n5407_));
  OAI21_X1   g05135(.A1(new_n5155_), .A2(new_n5157_), .B(new_n4890_), .ZN(new_n5408_));
  NAND3_X1   g05136(.A1(new_n5168_), .A2(new_n5165_), .A3(new_n5157_), .ZN(new_n5409_));
  NAND3_X1   g05137(.A1(new_n5408_), .A2(new_n5162_), .A3(new_n5409_), .ZN(new_n5410_));
  XOR2_X1    g05138(.A1(new_n5124_), .A2(\a[35] ), .Z(new_n5411_));
  NAND2_X1   g05139(.A1(new_n5117_), .A2(new_n5118_), .ZN(new_n5412_));
  INV_X1     g05140(.I(new_n5118_), .ZN(new_n5413_));
  NAND2_X1   g05141(.A1(new_n5413_), .A2(new_n5128_), .ZN(new_n5414_));
  AOI21_X1   g05142(.A1(new_n5414_), .A2(new_n5412_), .B(new_n5411_), .ZN(new_n5415_));
  INV_X1     g05143(.I(new_n5415_), .ZN(new_n5416_));
  AOI21_X1   g05144(.A1(new_n5158_), .A2(new_n4875_), .B(new_n4856_), .ZN(new_n5417_));
  OAI21_X1   g05145(.A1(new_n5158_), .A2(new_n4875_), .B(new_n4883_), .ZN(new_n5418_));
  XOR2_X1    g05146(.A1(\a[36] ), .A2(\a[38] ), .Z(new_n5419_));
  NAND2_X1   g05147(.A1(new_n5110_), .A2(new_n5419_), .ZN(new_n5420_));
  NOR2_X1    g05148(.A1(new_n5112_), .A2(new_n269_), .ZN(new_n5421_));
  OAI22_X1   g05149(.A1(new_n280_), .A2(new_n5420_), .B1(new_n5107_), .B2(new_n298_), .ZN(new_n5422_));
  NOR2_X1    g05150(.A1(new_n5422_), .A2(new_n5421_), .ZN(new_n5423_));
  NOR3_X1    g05151(.A1(new_n5423_), .A2(new_n403_), .A3(new_n5420_), .ZN(new_n5424_));
  NOR2_X1    g05152(.A1(new_n5424_), .A2(new_n4860_), .ZN(new_n5425_));
  NOR4_X1    g05153(.A1(new_n5423_), .A2(\a[38] ), .A3(new_n403_), .A4(new_n5420_), .ZN(new_n5426_));
  XOR2_X1    g05154(.A1(\a[38] ), .A2(\a[39] ), .Z(new_n5427_));
  NAND2_X1   g05155(.A1(new_n5427_), .A2(\b[0] ), .ZN(new_n5428_));
  INV_X1     g05156(.I(new_n5428_), .ZN(new_n5429_));
  OAI21_X1   g05157(.A1(new_n5425_), .A2(new_n5426_), .B(new_n5429_), .ZN(new_n5430_));
  NOR2_X1    g05158(.A1(new_n5117_), .A2(new_n5430_), .ZN(new_n5431_));
  NAND2_X1   g05159(.A1(new_n5117_), .A2(new_n5430_), .ZN(new_n5432_));
  INV_X1     g05160(.I(new_n5432_), .ZN(new_n5433_));
  OAI21_X1   g05161(.A1(new_n5433_), .A2(new_n5431_), .B(new_n5118_), .ZN(new_n5434_));
  NOR2_X1    g05162(.A1(new_n5433_), .A2(new_n5431_), .ZN(new_n5435_));
  NAND2_X1   g05163(.A1(new_n5435_), .A2(new_n5413_), .ZN(new_n5436_));
  INV_X1     g05164(.I(new_n4064_), .ZN(new_n5437_));
  NAND2_X1   g05165(.A1(new_n5437_), .A2(new_n4065_), .ZN(new_n5438_));
  AOI22_X1   g05166(.A1(new_n4062_), .A2(\b[5] ), .B1(new_n5438_), .B2(\b[6] ), .ZN(new_n5439_));
  AOI21_X1   g05167(.A1(\b[4] ), .A2(new_n4319_), .B(new_n5439_), .ZN(new_n5440_));
  OAI21_X1   g05168(.A1(new_n5440_), .A2(\a[35] ), .B(new_n4062_), .ZN(new_n5441_));
  XOR2_X1    g05169(.A1(new_n556_), .A2(new_n5441_), .Z(new_n5442_));
  AOI21_X1   g05170(.A1(new_n5436_), .A2(new_n5434_), .B(new_n5442_), .ZN(new_n5443_));
  OAI21_X1   g05171(.A1(new_n5417_), .A2(new_n5418_), .B(new_n5443_), .ZN(new_n5444_));
  INV_X1     g05172(.I(new_n5444_), .ZN(new_n5445_));
  NOR3_X1    g05173(.A1(new_n5417_), .A2(new_n5418_), .A3(new_n5443_), .ZN(new_n5446_));
  OAI21_X1   g05174(.A1(new_n5445_), .A2(new_n5446_), .B(new_n5416_), .ZN(new_n5447_));
  INV_X1     g05175(.I(new_n5446_), .ZN(new_n5448_));
  NAND3_X1   g05176(.A1(new_n5448_), .A2(new_n5415_), .A3(new_n5444_), .ZN(new_n5449_));
  OAI22_X1   g05177(.A1(new_n515_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n565_), .ZN(new_n5450_));
  OAI21_X1   g05178(.A1(new_n472_), .A2(new_n3569_), .B(new_n5450_), .ZN(new_n5451_));
  AOI21_X1   g05179(.A1(new_n5451_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n5452_));
  XOR2_X1    g05180(.A1(new_n759_), .A2(new_n5452_), .Z(new_n5453_));
  AOI21_X1   g05181(.A1(new_n5447_), .A2(new_n5449_), .B(new_n5453_), .ZN(new_n5454_));
  NAND2_X1   g05182(.A1(new_n5454_), .A2(new_n5410_), .ZN(new_n5455_));
  AND3_X2    g05183(.A1(new_n5408_), .A2(new_n5162_), .A3(new_n5409_), .Z(new_n5456_));
  AOI21_X1   g05184(.A1(new_n5448_), .A2(new_n5444_), .B(new_n5415_), .ZN(new_n5457_));
  NOR3_X1    g05185(.A1(new_n5445_), .A2(new_n5416_), .A3(new_n5446_), .ZN(new_n5458_));
  INV_X1     g05186(.I(new_n5453_), .ZN(new_n5459_));
  OAI21_X1   g05187(.A1(new_n5458_), .A2(new_n5457_), .B(new_n5459_), .ZN(new_n5460_));
  NAND2_X1   g05188(.A1(new_n5460_), .A2(new_n5456_), .ZN(new_n5461_));
  AOI21_X1   g05189(.A1(new_n5461_), .A2(new_n5455_), .B(new_n5407_), .ZN(new_n5462_));
  INV_X1     g05190(.I(new_n5407_), .ZN(new_n5463_));
  NOR2_X1    g05191(.A1(new_n5460_), .A2(new_n5456_), .ZN(new_n5464_));
  NOR2_X1    g05192(.A1(new_n5454_), .A2(new_n5410_), .ZN(new_n5465_));
  NOR3_X1    g05193(.A1(new_n5464_), .A2(new_n5465_), .A3(new_n5463_), .ZN(new_n5466_));
  OAI22_X1   g05194(.A1(new_n706_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n780_), .ZN(new_n5467_));
  OAI21_X1   g05195(.A1(new_n656_), .A2(new_n2884_), .B(new_n5467_), .ZN(new_n5468_));
  AOI21_X1   g05196(.A1(new_n5468_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n5469_));
  XOR2_X1    g05197(.A1(new_n785_), .A2(new_n5469_), .Z(new_n5470_));
  INV_X1     g05198(.I(new_n5470_), .ZN(new_n5471_));
  OAI21_X1   g05199(.A1(new_n5466_), .A2(new_n5462_), .B(new_n5471_), .ZN(new_n5472_));
  AOI21_X1   g05200(.A1(new_n5404_), .A2(new_n5403_), .B(new_n5472_), .ZN(new_n5473_));
  OAI21_X1   g05201(.A1(new_n4907_), .A2(new_n5182_), .B(new_n5103_), .ZN(new_n5474_));
  OAI21_X1   g05202(.A1(new_n5464_), .A2(new_n5465_), .B(new_n5463_), .ZN(new_n5475_));
  NAND3_X1   g05203(.A1(new_n5461_), .A2(new_n5455_), .A3(new_n5407_), .ZN(new_n5476_));
  AOI21_X1   g05204(.A1(new_n5475_), .A2(new_n5476_), .B(new_n5470_), .ZN(new_n5477_));
  NOR3_X1    g05205(.A1(new_n5477_), .A2(new_n5474_), .A3(new_n5402_), .ZN(new_n5478_));
  OAI21_X1   g05206(.A1(new_n5473_), .A2(new_n5478_), .B(new_n5181_), .ZN(new_n5479_));
  OAI21_X1   g05207(.A1(new_n5402_), .A2(new_n5474_), .B(new_n5477_), .ZN(new_n5480_));
  NAND3_X1   g05208(.A1(new_n5404_), .A2(new_n5472_), .A3(new_n5403_), .ZN(new_n5481_));
  NAND3_X1   g05209(.A1(new_n5481_), .A2(new_n5191_), .A3(new_n5480_), .ZN(new_n5482_));
  OAI22_X1   g05210(.A1(new_n2171_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n2166_), .ZN(new_n5483_));
  OAI21_X1   g05211(.A1(new_n861_), .A2(new_n2322_), .B(new_n5483_), .ZN(new_n5484_));
  AOI21_X1   g05212(.A1(new_n5484_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n5485_));
  XOR2_X1    g05213(.A1(new_n1024_), .A2(new_n5485_), .Z(new_n5486_));
  AOI21_X1   g05214(.A1(new_n5479_), .A2(new_n5482_), .B(new_n5486_), .ZN(new_n5487_));
  OAI21_X1   g05215(.A1(new_n5401_), .A2(new_n5400_), .B(new_n5487_), .ZN(new_n5488_));
  INV_X1     g05216(.I(new_n5400_), .ZN(new_n5489_));
  INV_X1     g05217(.I(new_n5401_), .ZN(new_n5490_));
  AOI21_X1   g05218(.A1(new_n5481_), .A2(new_n5480_), .B(new_n5191_), .ZN(new_n5491_));
  NOR3_X1    g05219(.A1(new_n5473_), .A2(new_n5478_), .A3(new_n5181_), .ZN(new_n5492_));
  INV_X1     g05220(.I(new_n5486_), .ZN(new_n5493_));
  OAI21_X1   g05221(.A1(new_n5492_), .A2(new_n5491_), .B(new_n5493_), .ZN(new_n5494_));
  NAND3_X1   g05222(.A1(new_n5490_), .A2(new_n5489_), .A3(new_n5494_), .ZN(new_n5495_));
  AOI21_X1   g05223(.A1(new_n5495_), .A2(new_n5488_), .B(new_n5398_), .ZN(new_n5496_));
  INV_X1     g05224(.I(new_n5398_), .ZN(new_n5497_));
  NOR2_X1    g05225(.A1(new_n5401_), .A2(new_n5400_), .ZN(new_n5498_));
  NOR2_X1    g05226(.A1(new_n5498_), .A2(new_n5494_), .ZN(new_n5499_));
  NOR3_X1    g05227(.A1(new_n5487_), .A2(new_n5401_), .A3(new_n5400_), .ZN(new_n5500_));
  NOR3_X1    g05228(.A1(new_n5499_), .A2(new_n5497_), .A3(new_n5500_), .ZN(new_n5501_));
  OAI22_X1   g05229(.A1(new_n1712_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n1707_), .ZN(new_n5502_));
  OAI21_X1   g05230(.A1(new_n1109_), .A2(new_n1850_), .B(new_n5502_), .ZN(new_n5503_));
  AOI21_X1   g05231(.A1(new_n5503_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n5504_));
  XOR2_X1    g05232(.A1(new_n1299_), .A2(new_n5504_), .Z(new_n5505_));
  INV_X1     g05233(.I(new_n5505_), .ZN(new_n5506_));
  OAI21_X1   g05234(.A1(new_n5501_), .A2(new_n5496_), .B(new_n5506_), .ZN(new_n5507_));
  NOR2_X1    g05235(.A1(new_n5397_), .A2(new_n5507_), .ZN(new_n5508_));
  AOI21_X1   g05236(.A1(new_n5229_), .A2(new_n5226_), .B(new_n5101_), .ZN(new_n5509_));
  OAI21_X1   g05237(.A1(new_n5509_), .A2(new_n4953_), .B(new_n4825_), .ZN(new_n5510_));
  OAI21_X1   g05238(.A1(new_n5499_), .A2(new_n5500_), .B(new_n5497_), .ZN(new_n5511_));
  NAND3_X1   g05239(.A1(new_n5495_), .A2(new_n5398_), .A3(new_n5488_), .ZN(new_n5512_));
  AOI21_X1   g05240(.A1(new_n5511_), .A2(new_n5512_), .B(new_n5505_), .ZN(new_n5513_));
  NOR2_X1    g05241(.A1(new_n5510_), .A2(new_n5513_), .ZN(new_n5514_));
  OAI21_X1   g05242(.A1(new_n5508_), .A2(new_n5514_), .B(new_n5229_), .ZN(new_n5515_));
  NAND2_X1   g05243(.A1(new_n5510_), .A2(new_n5513_), .ZN(new_n5516_));
  NAND2_X1   g05244(.A1(new_n5397_), .A2(new_n5507_), .ZN(new_n5517_));
  NAND3_X1   g05245(.A1(new_n5517_), .A2(new_n5516_), .A3(new_n5234_), .ZN(new_n5518_));
  OAI22_X1   g05246(.A1(new_n1347_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n1344_), .ZN(new_n5519_));
  OAI21_X1   g05247(.A1(new_n1518_), .A2(new_n1457_), .B(new_n5519_), .ZN(new_n5520_));
  AOI21_X1   g05248(.A1(new_n5520_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n5521_));
  XNOR2_X1   g05249(.A1(new_n1638_), .A2(new_n5521_), .ZN(new_n5522_));
  AOI21_X1   g05250(.A1(new_n5515_), .A2(new_n5518_), .B(new_n5522_), .ZN(new_n5523_));
  NAND2_X1   g05251(.A1(new_n5395_), .A2(new_n5523_), .ZN(new_n5524_));
  OR2_X2     g05252(.A1(new_n5395_), .A2(new_n5523_), .Z(new_n5525_));
  AOI21_X1   g05253(.A1(new_n5525_), .A2(new_n5524_), .B(new_n5252_), .ZN(new_n5526_));
  INV_X1     g05254(.I(new_n5524_), .ZN(new_n5527_));
  NOR2_X1    g05255(.A1(new_n5395_), .A2(new_n5523_), .ZN(new_n5528_));
  NOR3_X1    g05256(.A1(new_n5527_), .A2(new_n5245_), .A3(new_n5528_), .ZN(new_n5529_));
  OAI22_X1   g05257(.A1(new_n1055_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n1061_), .ZN(new_n5530_));
  OAI21_X1   g05258(.A1(new_n1803_), .A2(new_n1332_), .B(new_n5530_), .ZN(new_n5531_));
  AOI21_X1   g05259(.A1(new_n5531_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n5532_));
  XOR2_X1    g05260(.A1(new_n2106_), .A2(new_n5532_), .Z(new_n5533_));
  INV_X1     g05261(.I(new_n5533_), .ZN(new_n5534_));
  OAI21_X1   g05262(.A1(new_n5529_), .A2(new_n5526_), .B(new_n5534_), .ZN(new_n5535_));
  NOR2_X1    g05263(.A1(new_n5393_), .A2(new_n5535_), .ZN(new_n5536_));
  NAND2_X1   g05264(.A1(new_n5255_), .A2(new_n5277_), .ZN(new_n5537_));
  AOI21_X1   g05265(.A1(new_n5537_), .A2(new_n5390_), .B(new_n5266_), .ZN(new_n5538_));
  OAI21_X1   g05266(.A1(new_n5538_), .A2(new_n4988_), .B(new_n4993_), .ZN(new_n5539_));
  OAI21_X1   g05267(.A1(new_n5527_), .A2(new_n5528_), .B(new_n5245_), .ZN(new_n5540_));
  NAND3_X1   g05268(.A1(new_n5525_), .A2(new_n5252_), .A3(new_n5524_), .ZN(new_n5541_));
  AOI21_X1   g05269(.A1(new_n5540_), .A2(new_n5541_), .B(new_n5533_), .ZN(new_n5542_));
  NOR2_X1    g05270(.A1(new_n5539_), .A2(new_n5542_), .ZN(new_n5543_));
  OAI21_X1   g05271(.A1(new_n5536_), .A2(new_n5543_), .B(new_n5388_), .ZN(new_n5544_));
  INV_X1     g05272(.I(new_n5388_), .ZN(new_n5545_));
  NAND2_X1   g05273(.A1(new_n5539_), .A2(new_n5542_), .ZN(new_n5546_));
  NAND2_X1   g05274(.A1(new_n5393_), .A2(new_n5535_), .ZN(new_n5547_));
  NAND3_X1   g05275(.A1(new_n5547_), .A2(new_n5546_), .A3(new_n5545_), .ZN(new_n5548_));
  OAI22_X1   g05276(.A1(new_n970_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n820_), .ZN(new_n5549_));
  OAI21_X1   g05277(.A1(new_n2281_), .A2(new_n894_), .B(new_n5549_), .ZN(new_n5550_));
  AOI21_X1   g05278(.A1(new_n5550_), .A2(new_n827_), .B(new_n970_), .ZN(new_n5551_));
  XNOR2_X1   g05279(.A1(new_n2647_), .A2(new_n5551_), .ZN(new_n5552_));
  AOI21_X1   g05280(.A1(new_n5544_), .A2(new_n5548_), .B(new_n5552_), .ZN(new_n5553_));
  OAI21_X1   g05281(.A1(new_n5385_), .A2(new_n5387_), .B(new_n5553_), .ZN(new_n5554_));
  INV_X1     g05282(.I(new_n5554_), .ZN(new_n5555_));
  NOR3_X1    g05283(.A1(new_n5385_), .A2(new_n5387_), .A3(new_n5553_), .ZN(new_n5556_));
  OAI21_X1   g05284(.A1(new_n5555_), .A2(new_n5556_), .B(new_n5384_), .ZN(new_n5557_));
  AOI21_X1   g05285(.A1(new_n5267_), .A2(new_n5266_), .B(new_n5272_), .ZN(new_n5558_));
  INV_X1     g05286(.I(new_n5380_), .ZN(new_n5559_));
  OAI21_X1   g05287(.A1(new_n5559_), .A2(new_n5558_), .B(new_n5092_), .ZN(new_n5560_));
  AOI21_X1   g05288(.A1(new_n5560_), .A2(new_n5382_), .B(new_n5263_), .ZN(new_n5561_));
  INV_X1     g05289(.I(new_n5556_), .ZN(new_n5562_));
  NAND3_X1   g05290(.A1(new_n5562_), .A2(new_n5561_), .A3(new_n5554_), .ZN(new_n5563_));
  OAI22_X1   g05291(.A1(new_n607_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n610_), .ZN(new_n5564_));
  OAI21_X1   g05292(.A1(new_n2842_), .A2(new_n684_), .B(new_n5564_), .ZN(new_n5565_));
  AOI21_X1   g05293(.A1(new_n5565_), .A2(new_n612_), .B(new_n607_), .ZN(new_n5566_));
  XNOR2_X1   g05294(.A1(new_n3264_), .A2(new_n5566_), .ZN(new_n5567_));
  INV_X1     g05295(.I(new_n5567_), .ZN(new_n5568_));
  NAND3_X1   g05296(.A1(new_n5557_), .A2(new_n5563_), .A3(new_n5568_), .ZN(new_n5569_));
  INV_X1     g05297(.I(new_n5569_), .ZN(new_n5570_));
  AOI21_X1   g05298(.A1(new_n5557_), .A2(new_n5563_), .B(new_n5568_), .ZN(new_n5571_));
  NOR2_X1    g05299(.A1(new_n5570_), .A2(new_n5571_), .ZN(new_n5572_));
  OAI21_X1   g05300(.A1(new_n5310_), .A2(new_n5309_), .B(new_n5024_), .ZN(new_n5573_));
  NAND2_X1   g05301(.A1(new_n5573_), .A2(new_n5304_), .ZN(new_n5574_));
  NAND3_X1   g05302(.A1(new_n5298_), .A2(new_n5301_), .A3(new_n5023_), .ZN(new_n5575_));
  NAND3_X1   g05303(.A1(new_n5574_), .A2(new_n5033_), .A3(new_n5575_), .ZN(new_n5576_));
  AOI21_X1   g05304(.A1(new_n5299_), .A2(new_n5300_), .B(new_n5297_), .ZN(new_n5577_));
  INV_X1     g05305(.I(new_n5577_), .ZN(new_n5578_));
  NAND2_X1   g05306(.A1(new_n5576_), .A2(new_n5578_), .ZN(new_n5579_));
  INV_X1     g05307(.I(new_n5571_), .ZN(new_n5580_));
  AOI21_X1   g05308(.A1(new_n5580_), .A2(new_n5569_), .B(new_n5577_), .ZN(new_n5581_));
  AOI22_X1   g05309(.A1(new_n5579_), .A2(new_n5572_), .B1(new_n5576_), .B2(new_n5581_), .ZN(new_n5582_));
  OAI22_X1   g05310(.A1(new_n448_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n450_), .ZN(new_n5583_));
  OAI21_X1   g05311(.A1(new_n3709_), .A2(new_n496_), .B(new_n5583_), .ZN(new_n5584_));
  AOI21_X1   g05312(.A1(new_n5584_), .A2(new_n452_), .B(new_n448_), .ZN(new_n5585_));
  XNOR2_X1   g05313(.A1(new_n3993_), .A2(new_n5585_), .ZN(new_n5586_));
  OR2_X2     g05314(.A1(new_n5582_), .A2(new_n5586_), .Z(new_n5587_));
  NOR2_X1    g05315(.A1(new_n5378_), .A2(new_n5587_), .ZN(new_n5588_));
  AND2_X2    g05316(.A1(new_n5378_), .A2(new_n5587_), .Z(new_n5589_));
  OAI21_X1   g05317(.A1(new_n5589_), .A2(new_n5588_), .B(new_n5374_), .ZN(new_n5590_));
  OR3_X2     g05318(.A1(new_n5589_), .A2(new_n5374_), .A3(new_n5588_), .Z(new_n5591_));
  NAND2_X1   g05319(.A1(new_n5591_), .A2(new_n5590_), .ZN(new_n5592_));
  OAI22_X1   g05320(.A1(new_n4500_), .A2(new_n341_), .B1(new_n404_), .B2(new_n4774_), .ZN(new_n5593_));
  OAI21_X1   g05321(.A1(new_n4253_), .A2(new_n366_), .B(new_n5593_), .ZN(new_n5594_));
  AOI21_X1   g05322(.A1(new_n5594_), .A2(new_n334_), .B(new_n341_), .ZN(new_n5595_));
  XNOR2_X1   g05323(.A1(new_n4778_), .A2(new_n5595_), .ZN(new_n5596_));
  XOR2_X1    g05324(.A1(new_n5592_), .A2(new_n5596_), .Z(new_n5597_));
  XNOR2_X1   g05325(.A1(\b[37] ), .A2(\b[39] ), .ZN(new_n5598_));
  NOR2_X1    g05326(.A1(new_n5598_), .A2(new_n5352_), .ZN(new_n5599_));
  XNOR2_X1   g05327(.A1(new_n5351_), .A2(new_n5599_), .ZN(new_n5600_));
  NAND2_X1   g05328(.A1(new_n286_), .A2(\b[38] ), .ZN(new_n5601_));
  AOI22_X1   g05329(.A1(new_n304_), .A2(\b[37] ), .B1(new_n262_), .B2(\b[39] ), .ZN(new_n5602_));
  AOI21_X1   g05330(.A1(new_n5601_), .A2(new_n5602_), .B(new_n426_), .ZN(new_n5603_));
  NAND2_X1   g05331(.A1(new_n5600_), .A2(new_n5603_), .ZN(new_n5604_));
  XOR2_X1    g05332(.A1(new_n5604_), .A2(\a[2] ), .Z(new_n5605_));
  XNOR2_X1   g05333(.A1(new_n5597_), .A2(new_n5605_), .ZN(new_n5606_));
  NOR2_X1    g05334(.A1(new_n5606_), .A2(new_n5372_), .ZN(new_n5607_));
  XOR2_X1    g05335(.A1(new_n5597_), .A2(new_n5605_), .Z(new_n5608_));
  NOR2_X1    g05336(.A1(new_n5608_), .A2(new_n5371_), .ZN(new_n5609_));
  NOR2_X1    g05337(.A1(new_n5607_), .A2(new_n5609_), .ZN(new_n5610_));
  NOR2_X1    g05338(.A1(new_n5364_), .A2(new_n5610_), .ZN(new_n5611_));
  XOR2_X1    g05339(.A1(new_n5611_), .A2(new_n5367_), .Z(new_n5612_));
  XOR2_X1    g05340(.A1(new_n5612_), .A2(new_n5081_), .Z(\f[39] ));
  INV_X1     g05341(.I(new_n5592_), .ZN(new_n5614_));
  INV_X1     g05342(.I(new_n5596_), .ZN(new_n5615_));
  OAI21_X1   g05343(.A1(new_n5592_), .A2(new_n5615_), .B(new_n5371_), .ZN(new_n5616_));
  OAI21_X1   g05344(.A1(new_n5614_), .A2(new_n5596_), .B(new_n5616_), .ZN(new_n5617_));
  NOR2_X1    g05345(.A1(new_n5582_), .A2(new_n5374_), .ZN(new_n5618_));
  AOI21_X1   g05346(.A1(new_n5582_), .A2(new_n5374_), .B(new_n5586_), .ZN(new_n5619_));
  AOI21_X1   g05347(.A1(new_n5378_), .A2(new_n5619_), .B(new_n5618_), .ZN(new_n5620_));
  AOI21_X1   g05348(.A1(new_n5557_), .A2(new_n5563_), .B(new_n5578_), .ZN(new_n5621_));
  INV_X1     g05349(.I(new_n5621_), .ZN(new_n5622_));
  NAND2_X1   g05350(.A1(new_n5557_), .A2(new_n5563_), .ZN(new_n5623_));
  OAI21_X1   g05351(.A1(new_n5623_), .A2(new_n5577_), .B(new_n5568_), .ZN(new_n5624_));
  OAI21_X1   g05352(.A1(new_n5576_), .A2(new_n5624_), .B(new_n5622_), .ZN(new_n5625_));
  AOI21_X1   g05353(.A1(new_n5544_), .A2(new_n5548_), .B(new_n5384_), .ZN(new_n5626_));
  AOI21_X1   g05354(.A1(new_n5547_), .A2(new_n5546_), .B(new_n5545_), .ZN(new_n5627_));
  NOR3_X1    g05355(.A1(new_n5536_), .A2(new_n5543_), .A3(new_n5388_), .ZN(new_n5628_));
  NOR3_X1    g05356(.A1(new_n5628_), .A2(new_n5627_), .A3(new_n5561_), .ZN(new_n5629_));
  NOR4_X1    g05357(.A1(new_n5385_), .A2(new_n5387_), .A3(new_n5629_), .A4(new_n5552_), .ZN(new_n5630_));
  NOR2_X1    g05358(.A1(new_n5529_), .A2(new_n5526_), .ZN(new_n5631_));
  NAND3_X1   g05359(.A1(new_n5540_), .A2(new_n5541_), .A3(new_n5388_), .ZN(new_n5632_));
  NAND2_X1   g05360(.A1(new_n5632_), .A2(new_n5534_), .ZN(new_n5633_));
  OAI22_X1   g05361(.A1(new_n5633_), .A2(new_n5539_), .B1(new_n5388_), .B2(new_n5631_), .ZN(new_n5634_));
  AOI21_X1   g05362(.A1(new_n5515_), .A2(new_n5518_), .B(new_n5245_), .ZN(new_n5635_));
  INV_X1     g05363(.I(new_n5635_), .ZN(new_n5636_));
  OAI21_X1   g05364(.A1(new_n5251_), .A2(new_n5252_), .B(new_n5250_), .ZN(new_n5637_));
  NAND2_X1   g05365(.A1(new_n5637_), .A2(new_n5093_), .ZN(new_n5638_));
  INV_X1     g05366(.I(new_n5522_), .ZN(new_n5639_));
  NAND3_X1   g05367(.A1(new_n5515_), .A2(new_n5518_), .A3(new_n5245_), .ZN(new_n5640_));
  NAND4_X1   g05368(.A1(new_n5638_), .A2(new_n5640_), .A3(new_n4820_), .A4(new_n5639_), .ZN(new_n5641_));
  NAND2_X1   g05369(.A1(new_n5641_), .A2(new_n5636_), .ZN(new_n5642_));
  NAND2_X1   g05370(.A1(new_n5511_), .A2(new_n5512_), .ZN(new_n5643_));
  NAND2_X1   g05371(.A1(new_n5643_), .A2(new_n5234_), .ZN(new_n5644_));
  OAI21_X1   g05372(.A1(new_n5643_), .A2(new_n5234_), .B(new_n5506_), .ZN(new_n5645_));
  OAI21_X1   g05373(.A1(new_n5645_), .A2(new_n5510_), .B(new_n5644_), .ZN(new_n5646_));
  NOR2_X1    g05374(.A1(new_n5474_), .A2(new_n5402_), .ZN(new_n5647_));
  NAND2_X1   g05375(.A1(new_n5475_), .A2(new_n5476_), .ZN(new_n5648_));
  NOR3_X1    g05376(.A1(new_n5466_), .A2(new_n5462_), .A3(new_n5191_), .ZN(new_n5649_));
  NOR2_X1    g05377(.A1(new_n5649_), .A2(new_n5470_), .ZN(new_n5650_));
  AOI22_X1   g05378(.A1(new_n5650_), .A2(new_n5647_), .B1(new_n5191_), .B2(new_n5648_), .ZN(new_n5651_));
  AOI21_X1   g05379(.A1(new_n5447_), .A2(new_n5449_), .B(new_n5463_), .ZN(new_n5652_));
  NOR3_X1    g05380(.A1(new_n5458_), .A2(new_n5457_), .A3(new_n5407_), .ZN(new_n5653_));
  NOR3_X1    g05381(.A1(new_n5653_), .A2(new_n5410_), .A3(new_n5453_), .ZN(new_n5654_));
  AOI21_X1   g05382(.A1(new_n5436_), .A2(new_n5434_), .B(new_n5416_), .ZN(new_n5655_));
  INV_X1     g05383(.I(new_n5655_), .ZN(new_n5656_));
  OAI21_X1   g05384(.A1(new_n5146_), .A2(new_n5147_), .B(new_n4875_), .ZN(new_n5657_));
  NAND2_X1   g05385(.A1(new_n5657_), .A2(new_n4855_), .ZN(new_n5658_));
  NOR3_X1    g05386(.A1(new_n5146_), .A2(new_n5147_), .A3(new_n4875_), .ZN(new_n5659_));
  NOR2_X1    g05387(.A1(new_n5659_), .A2(new_n4851_), .ZN(new_n5660_));
  INV_X1     g05388(.I(new_n5442_), .ZN(new_n5661_));
  NAND3_X1   g05389(.A1(new_n5436_), .A2(new_n5434_), .A3(new_n5416_), .ZN(new_n5662_));
  NAND4_X1   g05390(.A1(new_n5660_), .A2(new_n5658_), .A3(new_n5662_), .A4(new_n5661_), .ZN(new_n5663_));
  NAND2_X1   g05391(.A1(new_n5663_), .A2(new_n5656_), .ZN(new_n5664_));
  NOR2_X1    g05392(.A1(new_n5425_), .A2(new_n5426_), .ZN(new_n5665_));
  NOR2_X1    g05393(.A1(new_n5128_), .A2(new_n5665_), .ZN(new_n5666_));
  INV_X1     g05394(.I(new_n5666_), .ZN(new_n5667_));
  NAND2_X1   g05395(.A1(new_n5128_), .A2(new_n5665_), .ZN(new_n5668_));
  NOR2_X1    g05396(.A1(new_n5118_), .A2(new_n5428_), .ZN(new_n5669_));
  NAND2_X1   g05397(.A1(new_n5668_), .A2(new_n5669_), .ZN(new_n5670_));
  AOI22_X1   g05398(.A1(new_n4859_), .A2(\b[3] ), .B1(new_n4865_), .B2(\b[4] ), .ZN(new_n5671_));
  NOR2_X1    g05399(.A1(new_n5112_), .A2(new_n280_), .ZN(new_n5672_));
  OAI21_X1   g05400(.A1(new_n5671_), .A2(new_n5672_), .B(new_n4860_), .ZN(new_n5673_));
  NAND3_X1   g05401(.A1(new_n5673_), .A2(new_n807_), .A3(new_n4859_), .ZN(new_n5674_));
  INV_X1     g05402(.I(new_n5674_), .ZN(new_n5675_));
  AOI21_X1   g05403(.A1(new_n5673_), .A2(new_n4859_), .B(new_n807_), .ZN(new_n5676_));
  NOR2_X1    g05404(.A1(new_n5675_), .A2(new_n5676_), .ZN(new_n5677_));
  XNOR2_X1   g05405(.A1(\a[39] ), .A2(\a[41] ), .ZN(new_n5678_));
  XNOR2_X1   g05406(.A1(\a[38] ), .A2(\a[40] ), .ZN(new_n5679_));
  NOR2_X1    g05407(.A1(new_n5679_), .A2(new_n5678_), .ZN(new_n5680_));
  INV_X1     g05408(.I(\a[41] ), .ZN(new_n5681_));
  INV_X1     g05409(.I(\a[39] ), .ZN(new_n5682_));
  NAND3_X1   g05410(.A1(new_n4860_), .A2(new_n5682_), .A3(\a[40] ), .ZN(new_n5683_));
  INV_X1     g05411(.I(\a[40] ), .ZN(new_n5684_));
  NAND3_X1   g05412(.A1(new_n5684_), .A2(\a[38] ), .A3(\a[39] ), .ZN(new_n5685_));
  NAND2_X1   g05413(.A1(new_n5683_), .A2(new_n5685_), .ZN(new_n5686_));
  NAND2_X1   g05414(.A1(new_n5686_), .A2(\b[1] ), .ZN(new_n5687_));
  XOR2_X1    g05415(.A1(\a[39] ), .A2(\a[41] ), .Z(new_n5688_));
  XOR2_X1    g05416(.A1(\a[38] ), .A2(\a[40] ), .Z(new_n5689_));
  NAND3_X1   g05417(.A1(new_n5689_), .A2(new_n5688_), .A3(\b[0] ), .ZN(new_n5690_));
  NAND3_X1   g05418(.A1(new_n5687_), .A2(new_n5690_), .A3(new_n5681_), .ZN(new_n5691_));
  NAND3_X1   g05419(.A1(new_n5691_), .A2(new_n444_), .A3(new_n5680_), .ZN(new_n5692_));
  AOI21_X1   g05420(.A1(new_n5691_), .A2(new_n5680_), .B(new_n444_), .ZN(new_n5693_));
  INV_X1     g05421(.I(new_n5693_), .ZN(new_n5694_));
  NOR2_X1    g05422(.A1(new_n5429_), .A2(new_n5681_), .ZN(new_n5695_));
  INV_X1     g05423(.I(new_n5695_), .ZN(new_n5696_));
  NAND3_X1   g05424(.A1(new_n5694_), .A2(new_n5692_), .A3(new_n5696_), .ZN(new_n5697_));
  INV_X1     g05425(.I(new_n5692_), .ZN(new_n5698_));
  OAI21_X1   g05426(.A1(new_n5698_), .A2(new_n5693_), .B(new_n5695_), .ZN(new_n5699_));
  NAND2_X1   g05427(.A1(new_n5697_), .A2(new_n5699_), .ZN(new_n5700_));
  INV_X1     g05428(.I(new_n5700_), .ZN(new_n5701_));
  NOR2_X1    g05429(.A1(new_n5701_), .A2(new_n5677_), .ZN(new_n5702_));
  INV_X1     g05430(.I(new_n5702_), .ZN(new_n5703_));
  NAND2_X1   g05431(.A1(new_n5701_), .A2(new_n5677_), .ZN(new_n5704_));
  AOI22_X1   g05432(.A1(new_n5703_), .A2(new_n5704_), .B1(new_n5670_), .B2(new_n5667_), .ZN(new_n5705_));
  NAND2_X1   g05433(.A1(new_n5670_), .A2(new_n5667_), .ZN(new_n5706_));
  NAND2_X1   g05434(.A1(new_n5677_), .A2(new_n5700_), .ZN(new_n5707_));
  INV_X1     g05435(.I(new_n5676_), .ZN(new_n5708_));
  NAND2_X1   g05436(.A1(new_n5708_), .A2(new_n5674_), .ZN(new_n5709_));
  NAND3_X1   g05437(.A1(new_n5709_), .A2(new_n5697_), .A3(new_n5699_), .ZN(new_n5710_));
  AOI21_X1   g05438(.A1(new_n5707_), .A2(new_n5710_), .B(new_n5706_), .ZN(new_n5711_));
  AOI22_X1   g05439(.A1(new_n4062_), .A2(\b[6] ), .B1(new_n5438_), .B2(\b[7] ), .ZN(new_n5712_));
  AOI21_X1   g05440(.A1(\b[5] ), .A2(new_n4319_), .B(new_n5712_), .ZN(new_n5713_));
  OAI21_X1   g05441(.A1(new_n5713_), .A2(\a[35] ), .B(new_n4062_), .ZN(new_n5714_));
  XNOR2_X1   g05442(.A1(new_n471_), .A2(new_n5714_), .ZN(new_n5715_));
  INV_X1     g05443(.I(new_n5715_), .ZN(new_n5716_));
  OAI21_X1   g05444(.A1(new_n5711_), .A2(new_n5705_), .B(new_n5716_), .ZN(new_n5717_));
  INV_X1     g05445(.I(new_n5705_), .ZN(new_n5718_));
  INV_X1     g05446(.I(new_n5706_), .ZN(new_n5719_));
  NAND2_X1   g05447(.A1(new_n5710_), .A2(new_n5707_), .ZN(new_n5720_));
  NAND2_X1   g05448(.A1(new_n5719_), .A2(new_n5720_), .ZN(new_n5721_));
  NAND3_X1   g05449(.A1(new_n5721_), .A2(new_n5718_), .A3(new_n5715_), .ZN(new_n5722_));
  NAND2_X1   g05450(.A1(new_n5722_), .A2(new_n5717_), .ZN(new_n5723_));
  NAND2_X1   g05451(.A1(new_n5664_), .A2(new_n5723_), .ZN(new_n5724_));
  NAND3_X1   g05452(.A1(new_n5721_), .A2(new_n5718_), .A3(new_n5716_), .ZN(new_n5725_));
  OAI21_X1   g05453(.A1(new_n5711_), .A2(new_n5705_), .B(new_n5715_), .ZN(new_n5726_));
  NAND2_X1   g05454(.A1(new_n5725_), .A2(new_n5726_), .ZN(new_n5727_));
  NAND3_X1   g05455(.A1(new_n5727_), .A2(new_n5663_), .A3(new_n5656_), .ZN(new_n5728_));
  NAND2_X1   g05456(.A1(new_n5724_), .A2(new_n5728_), .ZN(new_n5729_));
  OAI22_X1   g05457(.A1(new_n565_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n656_), .ZN(new_n5730_));
  OAI21_X1   g05458(.A1(new_n515_), .A2(new_n3569_), .B(new_n5730_), .ZN(new_n5731_));
  AOI21_X1   g05459(.A1(new_n5731_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n5732_));
  XNOR2_X1   g05460(.A1(new_n660_), .A2(new_n5732_), .ZN(new_n5733_));
  NOR2_X1    g05461(.A1(new_n5729_), .A2(new_n5733_), .ZN(new_n5734_));
  INV_X1     g05462(.I(new_n5733_), .ZN(new_n5735_));
  AOI21_X1   g05463(.A1(new_n5724_), .A2(new_n5728_), .B(new_n5735_), .ZN(new_n5736_));
  OAI22_X1   g05464(.A1(new_n5654_), .A2(new_n5652_), .B1(new_n5734_), .B2(new_n5736_), .ZN(new_n5737_));
  NAND3_X1   g05465(.A1(new_n5447_), .A2(new_n5449_), .A3(new_n5463_), .ZN(new_n5738_));
  NOR2_X1    g05466(.A1(new_n5410_), .A2(new_n5453_), .ZN(new_n5739_));
  AOI21_X1   g05467(.A1(new_n5739_), .A2(new_n5738_), .B(new_n5652_), .ZN(new_n5740_));
  AOI22_X1   g05468(.A1(new_n5663_), .A2(new_n5656_), .B1(new_n5717_), .B2(new_n5722_), .ZN(new_n5741_));
  INV_X1     g05469(.I(new_n5728_), .ZN(new_n5742_));
  OAI21_X1   g05470(.A1(new_n5742_), .A2(new_n5741_), .B(new_n5735_), .ZN(new_n5743_));
  NAND3_X1   g05471(.A1(new_n5724_), .A2(new_n5728_), .A3(new_n5733_), .ZN(new_n5744_));
  NAND2_X1   g05472(.A1(new_n5743_), .A2(new_n5744_), .ZN(new_n5745_));
  NAND2_X1   g05473(.A1(new_n5740_), .A2(new_n5745_), .ZN(new_n5746_));
  OAI22_X1   g05474(.A1(new_n780_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n861_), .ZN(new_n5747_));
  OAI21_X1   g05475(.A1(new_n706_), .A2(new_n2884_), .B(new_n5747_), .ZN(new_n5748_));
  AOI21_X1   g05476(.A1(new_n5748_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n5749_));
  XNOR2_X1   g05477(.A1(new_n860_), .A2(new_n5749_), .ZN(new_n5750_));
  INV_X1     g05478(.I(new_n5750_), .ZN(new_n5751_));
  NAND3_X1   g05479(.A1(new_n5737_), .A2(new_n5746_), .A3(new_n5751_), .ZN(new_n5752_));
  NOR2_X1    g05480(.A1(new_n5734_), .A2(new_n5736_), .ZN(new_n5753_));
  NOR2_X1    g05481(.A1(new_n5753_), .A2(new_n5740_), .ZN(new_n5754_));
  AOI21_X1   g05482(.A1(new_n5724_), .A2(new_n5728_), .B(new_n5733_), .ZN(new_n5755_));
  NOR3_X1    g05483(.A1(new_n5742_), .A2(new_n5741_), .A3(new_n5735_), .ZN(new_n5756_));
  NOR2_X1    g05484(.A1(new_n5756_), .A2(new_n5755_), .ZN(new_n5757_));
  NOR3_X1    g05485(.A1(new_n5654_), .A2(new_n5757_), .A3(new_n5652_), .ZN(new_n5758_));
  OAI21_X1   g05486(.A1(new_n5754_), .A2(new_n5758_), .B(new_n5750_), .ZN(new_n5759_));
  AOI21_X1   g05487(.A1(new_n5752_), .A2(new_n5759_), .B(new_n5651_), .ZN(new_n5760_));
  NOR2_X1    g05488(.A1(new_n5754_), .A2(new_n5758_), .ZN(new_n5761_));
  NOR2_X1    g05489(.A1(new_n5761_), .A2(new_n5750_), .ZN(new_n5762_));
  INV_X1     g05490(.I(new_n5762_), .ZN(new_n5763_));
  NAND2_X1   g05491(.A1(new_n5761_), .A2(new_n5750_), .ZN(new_n5764_));
  NAND2_X1   g05492(.A1(new_n5763_), .A2(new_n5764_), .ZN(new_n5765_));
  NAND2_X1   g05493(.A1(new_n5765_), .A2(new_n5651_), .ZN(new_n5766_));
  INV_X1     g05494(.I(new_n5766_), .ZN(new_n5767_));
  OAI22_X1   g05495(.A1(new_n2171_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n2166_), .ZN(new_n5768_));
  OAI21_X1   g05496(.A1(new_n930_), .A2(new_n2322_), .B(new_n5768_), .ZN(new_n5769_));
  AOI21_X1   g05497(.A1(new_n5769_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n5770_));
  XOR2_X1    g05498(.A1(new_n1114_), .A2(new_n5770_), .Z(new_n5771_));
  NOR3_X1    g05499(.A1(new_n5767_), .A2(new_n5760_), .A3(new_n5771_), .ZN(new_n5772_));
  INV_X1     g05500(.I(new_n5760_), .ZN(new_n5773_));
  INV_X1     g05501(.I(new_n5771_), .ZN(new_n5774_));
  AOI21_X1   g05502(.A1(new_n5773_), .A2(new_n5766_), .B(new_n5774_), .ZN(new_n5775_));
  NOR2_X1    g05503(.A1(new_n5775_), .A2(new_n5772_), .ZN(new_n5776_));
  INV_X1     g05504(.I(new_n5498_), .ZN(new_n5777_));
  AOI21_X1   g05505(.A1(new_n5479_), .A2(new_n5482_), .B(new_n5497_), .ZN(new_n5778_));
  INV_X1     g05506(.I(new_n5778_), .ZN(new_n5779_));
  NAND3_X1   g05507(.A1(new_n5479_), .A2(new_n5482_), .A3(new_n5497_), .ZN(new_n5780_));
  NAND2_X1   g05508(.A1(new_n5780_), .A2(new_n5493_), .ZN(new_n5781_));
  OAI21_X1   g05509(.A1(new_n5777_), .A2(new_n5781_), .B(new_n5779_), .ZN(new_n5782_));
  OAI22_X1   g05510(.A1(new_n1712_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n1707_), .ZN(new_n5783_));
  OAI21_X1   g05511(.A1(new_n1189_), .A2(new_n1850_), .B(new_n5783_), .ZN(new_n5784_));
  AOI21_X1   g05512(.A1(new_n5784_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n5785_));
  XNOR2_X1   g05513(.A1(new_n1421_), .A2(new_n5785_), .ZN(new_n5786_));
  INV_X1     g05514(.I(new_n5786_), .ZN(new_n5787_));
  NAND2_X1   g05515(.A1(new_n5782_), .A2(new_n5787_), .ZN(new_n5788_));
  NOR3_X1    g05516(.A1(new_n5492_), .A2(new_n5491_), .A3(new_n5398_), .ZN(new_n5789_));
  NOR4_X1    g05517(.A1(new_n5789_), .A2(new_n5401_), .A3(new_n5400_), .A4(new_n5486_), .ZN(new_n5790_));
  NOR3_X1    g05518(.A1(new_n5790_), .A2(new_n5778_), .A3(new_n5787_), .ZN(new_n5791_));
  INV_X1     g05519(.I(new_n5791_), .ZN(new_n5792_));
  AOI21_X1   g05520(.A1(new_n5788_), .A2(new_n5792_), .B(new_n5776_), .ZN(new_n5793_));
  NAND3_X1   g05521(.A1(new_n5773_), .A2(new_n5766_), .A3(new_n5774_), .ZN(new_n5794_));
  OAI21_X1   g05522(.A1(new_n5767_), .A2(new_n5760_), .B(new_n5771_), .ZN(new_n5795_));
  NAND2_X1   g05523(.A1(new_n5794_), .A2(new_n5795_), .ZN(new_n5796_));
  NOR3_X1    g05524(.A1(new_n5790_), .A2(new_n5778_), .A3(new_n5786_), .ZN(new_n5797_));
  INV_X1     g05525(.I(new_n5797_), .ZN(new_n5798_));
  OAI21_X1   g05526(.A1(new_n5790_), .A2(new_n5778_), .B(new_n5786_), .ZN(new_n5799_));
  AOI21_X1   g05527(.A1(new_n5798_), .A2(new_n5799_), .B(new_n5796_), .ZN(new_n5800_));
  OAI22_X1   g05528(.A1(new_n1347_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n1344_), .ZN(new_n5801_));
  OAI21_X1   g05529(.A1(new_n1525_), .A2(new_n1457_), .B(new_n5801_), .ZN(new_n5802_));
  AOI21_X1   g05530(.A1(new_n5802_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n5803_));
  XOR2_X1    g05531(.A1(new_n1808_), .A2(new_n5803_), .Z(new_n5804_));
  INV_X1     g05532(.I(new_n5804_), .ZN(new_n5805_));
  OAI21_X1   g05533(.A1(new_n5793_), .A2(new_n5800_), .B(new_n5805_), .ZN(new_n5806_));
  NOR2_X1    g05534(.A1(new_n5790_), .A2(new_n5778_), .ZN(new_n5807_));
  NOR2_X1    g05535(.A1(new_n5807_), .A2(new_n5786_), .ZN(new_n5808_));
  OAI21_X1   g05536(.A1(new_n5808_), .A2(new_n5791_), .B(new_n5796_), .ZN(new_n5809_));
  INV_X1     g05537(.I(new_n5799_), .ZN(new_n5810_));
  OAI21_X1   g05538(.A1(new_n5810_), .A2(new_n5797_), .B(new_n5776_), .ZN(new_n5811_));
  NAND3_X1   g05539(.A1(new_n5809_), .A2(new_n5811_), .A3(new_n5804_), .ZN(new_n5812_));
  NAND2_X1   g05540(.A1(new_n5806_), .A2(new_n5812_), .ZN(new_n5813_));
  NAND2_X1   g05541(.A1(new_n5813_), .A2(new_n5646_), .ZN(new_n5814_));
  NOR3_X1    g05542(.A1(new_n5501_), .A2(new_n5496_), .A3(new_n5234_), .ZN(new_n5815_));
  NOR2_X1    g05543(.A1(new_n5815_), .A2(new_n5505_), .ZN(new_n5816_));
  AOI22_X1   g05544(.A1(new_n5816_), .A2(new_n5397_), .B1(new_n5234_), .B2(new_n5643_), .ZN(new_n5817_));
  NAND2_X1   g05545(.A1(new_n5809_), .A2(new_n5811_), .ZN(new_n5818_));
  NOR2_X1    g05546(.A1(new_n5818_), .A2(new_n5804_), .ZN(new_n5819_));
  NOR2_X1    g05547(.A1(new_n5793_), .A2(new_n5800_), .ZN(new_n5820_));
  NOR2_X1    g05548(.A1(new_n5820_), .A2(new_n5805_), .ZN(new_n5821_));
  OAI21_X1   g05549(.A1(new_n5821_), .A2(new_n5819_), .B(new_n5817_), .ZN(new_n5822_));
  NAND2_X1   g05550(.A1(new_n5822_), .A2(new_n5814_), .ZN(new_n5823_));
  OAI22_X1   g05551(.A1(new_n1055_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n1061_), .ZN(new_n5824_));
  OAI21_X1   g05552(.A1(new_n1936_), .A2(new_n1332_), .B(new_n5824_), .ZN(new_n5825_));
  AOI21_X1   g05553(.A1(new_n5825_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n5826_));
  XNOR2_X1   g05554(.A1(new_n2280_), .A2(new_n5826_), .ZN(new_n5827_));
  XOR2_X1    g05555(.A1(new_n5823_), .A2(new_n5827_), .Z(new_n5828_));
  NAND2_X1   g05556(.A1(new_n5828_), .A2(new_n5642_), .ZN(new_n5829_));
  AOI21_X1   g05557(.A1(new_n5517_), .A2(new_n5516_), .B(new_n5234_), .ZN(new_n5830_));
  NOR3_X1    g05558(.A1(new_n5508_), .A2(new_n5514_), .A3(new_n5229_), .ZN(new_n5831_));
  NOR3_X1    g05559(.A1(new_n5830_), .A2(new_n5831_), .A3(new_n5252_), .ZN(new_n5832_));
  NOR3_X1    g05560(.A1(new_n5395_), .A2(new_n5832_), .A3(new_n5522_), .ZN(new_n5833_));
  NOR2_X1    g05561(.A1(new_n5833_), .A2(new_n5635_), .ZN(new_n5834_));
  INV_X1     g05562(.I(new_n5827_), .ZN(new_n5835_));
  XOR2_X1    g05563(.A1(new_n5823_), .A2(new_n5835_), .Z(new_n5836_));
  NAND2_X1   g05564(.A1(new_n5836_), .A2(new_n5834_), .ZN(new_n5837_));
  NAND2_X1   g05565(.A1(new_n5829_), .A2(new_n5837_), .ZN(new_n5838_));
  INV_X1     g05566(.I(new_n5838_), .ZN(new_n5839_));
  OAI22_X1   g05567(.A1(new_n970_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n820_), .ZN(new_n5840_));
  OAI21_X1   g05568(.A1(new_n2439_), .A2(new_n894_), .B(new_n5840_), .ZN(new_n5841_));
  AOI21_X1   g05569(.A1(new_n5841_), .A2(new_n827_), .B(new_n970_), .ZN(new_n5842_));
  XNOR2_X1   g05570(.A1(new_n2846_), .A2(new_n5842_), .ZN(new_n5843_));
  NOR2_X1    g05571(.A1(new_n5839_), .A2(new_n5843_), .ZN(new_n5844_));
  INV_X1     g05572(.I(new_n5843_), .ZN(new_n5845_));
  NOR2_X1    g05573(.A1(new_n5838_), .A2(new_n5845_), .ZN(new_n5846_));
  OAI21_X1   g05574(.A1(new_n5844_), .A2(new_n5846_), .B(new_n5634_), .ZN(new_n5847_));
  NOR2_X1    g05575(.A1(new_n5631_), .A2(new_n5388_), .ZN(new_n5848_));
  AOI21_X1   g05576(.A1(new_n5631_), .A2(new_n5388_), .B(new_n5533_), .ZN(new_n5849_));
  AOI21_X1   g05577(.A1(new_n5849_), .A2(new_n5393_), .B(new_n5848_), .ZN(new_n5850_));
  NOR2_X1    g05578(.A1(new_n5838_), .A2(new_n5843_), .ZN(new_n5851_));
  NOR2_X1    g05579(.A1(new_n5839_), .A2(new_n5845_), .ZN(new_n5852_));
  OAI21_X1   g05580(.A1(new_n5852_), .A2(new_n5851_), .B(new_n5850_), .ZN(new_n5853_));
  NAND2_X1   g05581(.A1(new_n5847_), .A2(new_n5853_), .ZN(new_n5854_));
  OAI21_X1   g05582(.A1(new_n5630_), .A2(new_n5626_), .B(new_n5854_), .ZN(new_n5855_));
  INV_X1     g05583(.I(new_n5626_), .ZN(new_n5856_));
  OAI21_X1   g05584(.A1(new_n5289_), .A2(new_n5288_), .B(new_n5014_), .ZN(new_n5857_));
  NAND2_X1   g05585(.A1(new_n5857_), .A2(new_n5003_), .ZN(new_n5858_));
  NOR3_X1    g05586(.A1(new_n5289_), .A2(new_n5288_), .A3(new_n5014_), .ZN(new_n5859_));
  NOR2_X1    g05587(.A1(new_n5859_), .A2(new_n5013_), .ZN(new_n5860_));
  INV_X1     g05588(.I(new_n5552_), .ZN(new_n5861_));
  NAND3_X1   g05589(.A1(new_n5384_), .A2(new_n5544_), .A3(new_n5548_), .ZN(new_n5862_));
  NAND4_X1   g05590(.A1(new_n5860_), .A2(new_n5858_), .A3(new_n5861_), .A4(new_n5862_), .ZN(new_n5863_));
  XOR2_X1    g05591(.A1(new_n5838_), .A2(new_n5845_), .Z(new_n5864_));
  XOR2_X1    g05592(.A1(new_n5838_), .A2(new_n5843_), .Z(new_n5865_));
  MUX2_X1    g05593(.I0(new_n5865_), .I1(new_n5864_), .S(new_n5634_), .Z(new_n5866_));
  NAND3_X1   g05594(.A1(new_n5863_), .A2(new_n5866_), .A3(new_n5856_), .ZN(new_n5867_));
  OAI22_X1   g05595(.A1(new_n607_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n610_), .ZN(new_n5868_));
  OAI21_X1   g05596(.A1(new_n3018_), .A2(new_n684_), .B(new_n5868_), .ZN(new_n5869_));
  AOI21_X1   g05597(.A1(new_n5869_), .A2(new_n612_), .B(new_n607_), .ZN(new_n5870_));
  XNOR2_X1   g05598(.A1(new_n3514_), .A2(new_n5870_), .ZN(new_n5871_));
  INV_X1     g05599(.I(new_n5871_), .ZN(new_n5872_));
  NAND3_X1   g05600(.A1(new_n5867_), .A2(new_n5855_), .A3(new_n5872_), .ZN(new_n5873_));
  AOI21_X1   g05601(.A1(new_n5863_), .A2(new_n5856_), .B(new_n5866_), .ZN(new_n5874_));
  NOR3_X1    g05602(.A1(new_n5630_), .A2(new_n5626_), .A3(new_n5854_), .ZN(new_n5875_));
  OAI21_X1   g05603(.A1(new_n5874_), .A2(new_n5875_), .B(new_n5871_), .ZN(new_n5876_));
  NAND2_X1   g05604(.A1(new_n5876_), .A2(new_n5873_), .ZN(new_n5877_));
  NAND2_X1   g05605(.A1(new_n5625_), .A2(new_n5877_), .ZN(new_n5878_));
  NOR2_X1    g05606(.A1(new_n5874_), .A2(new_n5875_), .ZN(new_n5879_));
  NOR2_X1    g05607(.A1(new_n5879_), .A2(new_n5871_), .ZN(new_n5880_));
  INV_X1     g05608(.I(new_n5879_), .ZN(new_n5881_));
  NOR2_X1    g05609(.A1(new_n5881_), .A2(new_n5872_), .ZN(new_n5882_));
  NOR2_X1    g05610(.A1(new_n5882_), .A2(new_n5880_), .ZN(new_n5883_));
  OAI21_X1   g05611(.A1(new_n5625_), .A2(new_n5883_), .B(new_n5878_), .ZN(new_n5884_));
  OAI22_X1   g05612(.A1(new_n448_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n450_), .ZN(new_n5885_));
  OAI21_X1   g05613(.A1(new_n3717_), .A2(new_n496_), .B(new_n5885_), .ZN(new_n5886_));
  AOI21_X1   g05614(.A1(new_n5886_), .A2(new_n452_), .B(new_n448_), .ZN(new_n5887_));
  XNOR2_X1   g05615(.A1(new_n4257_), .A2(new_n5887_), .ZN(new_n5888_));
  INV_X1     g05616(.I(new_n5888_), .ZN(new_n5889_));
  XOR2_X1    g05617(.A1(new_n5884_), .A2(new_n5889_), .Z(new_n5890_));
  OAI22_X1   g05618(.A1(new_n4774_), .A2(new_n341_), .B1(new_n404_), .B2(new_n5068_), .ZN(new_n5891_));
  OAI21_X1   g05619(.A1(new_n4500_), .A2(new_n366_), .B(new_n5891_), .ZN(new_n5892_));
  AOI21_X1   g05620(.A1(new_n5892_), .A2(new_n334_), .B(new_n341_), .ZN(new_n5893_));
  XOR2_X1    g05621(.A1(new_n5067_), .A2(new_n5893_), .Z(new_n5894_));
  INV_X1     g05622(.I(new_n5894_), .ZN(new_n5895_));
  NAND2_X1   g05623(.A1(new_n5890_), .A2(new_n5895_), .ZN(new_n5896_));
  INV_X1     g05624(.I(new_n5890_), .ZN(new_n5897_));
  NAND2_X1   g05625(.A1(new_n5897_), .A2(new_n5894_), .ZN(new_n5898_));
  AOI21_X1   g05626(.A1(new_n5898_), .A2(new_n5896_), .B(new_n5620_), .ZN(new_n5899_));
  INV_X1     g05627(.I(new_n5899_), .ZN(new_n5900_));
  INV_X1     g05628(.I(new_n5618_), .ZN(new_n5901_));
  OAI21_X1   g05629(.A1(new_n5326_), .A2(new_n5327_), .B(new_n5086_), .ZN(new_n5902_));
  NAND2_X1   g05630(.A1(new_n5902_), .A2(new_n5044_), .ZN(new_n5903_));
  NAND4_X1   g05631(.A1(new_n5903_), .A2(new_n5619_), .A3(new_n4804_), .A4(new_n5376_), .ZN(new_n5904_));
  NAND2_X1   g05632(.A1(new_n5904_), .A2(new_n5901_), .ZN(new_n5905_));
  NAND2_X1   g05633(.A1(new_n5897_), .A2(new_n5895_), .ZN(new_n5906_));
  NAND2_X1   g05634(.A1(new_n5890_), .A2(new_n5894_), .ZN(new_n5907_));
  AOI21_X1   g05635(.A1(new_n5906_), .A2(new_n5907_), .B(new_n5905_), .ZN(new_n5908_));
  INV_X1     g05636(.I(new_n5908_), .ZN(new_n5909_));
  NAND2_X1   g05637(.A1(new_n5900_), .A2(new_n5909_), .ZN(new_n5910_));
  NOR2_X1    g05638(.A1(\b[38] ), .A2(\b[39] ), .ZN(new_n5911_));
  AOI21_X1   g05639(.A1(new_n5351_), .A2(new_n5911_), .B(new_n5068_), .ZN(new_n5912_));
  INV_X1     g05640(.I(\b[39] ), .ZN(new_n5913_));
  NOR2_X1    g05641(.A1(new_n5353_), .A2(new_n5913_), .ZN(new_n5914_));
  INV_X1     g05642(.I(new_n5914_), .ZN(new_n5915_));
  NOR2_X1    g05643(.A1(new_n5351_), .A2(new_n5915_), .ZN(new_n5916_));
  NOR2_X1    g05644(.A1(new_n5912_), .A2(new_n5916_), .ZN(new_n5917_));
  INV_X1     g05645(.I(new_n5917_), .ZN(new_n5918_));
  XNOR2_X1   g05646(.A1(\b[39] ), .A2(\b[40] ), .ZN(new_n5919_));
  INV_X1     g05647(.I(new_n5919_), .ZN(new_n5920_));
  INV_X1     g05648(.I(\b[40] ), .ZN(new_n5921_));
  NOR2_X1    g05649(.A1(new_n5913_), .A2(new_n5921_), .ZN(new_n5922_));
  INV_X1     g05650(.I(new_n5922_), .ZN(new_n5923_));
  NAND2_X1   g05651(.A1(new_n5913_), .A2(new_n5921_), .ZN(new_n5924_));
  AOI21_X1   g05652(.A1(new_n5923_), .A2(new_n5924_), .B(new_n5918_), .ZN(new_n5925_));
  AOI21_X1   g05653(.A1(new_n5918_), .A2(new_n5920_), .B(new_n5925_), .ZN(new_n5926_));
  OAI22_X1   g05654(.A1(new_n330_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n263_), .ZN(new_n5927_));
  OAI21_X1   g05655(.A1(new_n5353_), .A2(new_n289_), .B(new_n5927_), .ZN(new_n5928_));
  AOI21_X1   g05656(.A1(new_n5928_), .A2(new_n260_), .B(new_n426_), .ZN(new_n5929_));
  XOR2_X1    g05657(.A1(new_n5926_), .A2(new_n5929_), .Z(new_n5930_));
  INV_X1     g05658(.I(new_n5930_), .ZN(new_n5931_));
  XOR2_X1    g05659(.A1(new_n5910_), .A2(new_n5931_), .Z(new_n5932_));
  AND2_X2    g05660(.A1(new_n5617_), .A2(new_n5932_), .Z(new_n5933_));
  XOR2_X1    g05661(.A1(new_n5910_), .A2(new_n5931_), .Z(new_n5934_));
  NOR2_X1    g05662(.A1(new_n5617_), .A2(new_n5934_), .ZN(new_n5935_));
  OR2_X2     g05663(.A1(new_n5933_), .A2(new_n5935_), .Z(new_n5936_));
  XOR2_X1    g05664(.A1(new_n5597_), .A2(new_n5371_), .Z(new_n5937_));
  OAI21_X1   g05665(.A1(new_n5610_), .A2(new_n5366_), .B(new_n5361_), .ZN(new_n5938_));
  NOR3_X1    g05666(.A1(new_n5607_), .A2(new_n5609_), .A3(new_n5345_), .ZN(new_n5939_));
  NOR2_X1    g05667(.A1(new_n5080_), .A2(new_n5939_), .ZN(new_n5940_));
  AOI22_X1   g05668(.A1(new_n5940_), .A2(new_n5938_), .B1(new_n5605_), .B2(new_n5937_), .ZN(new_n5941_));
  NAND2_X1   g05669(.A1(new_n5937_), .A2(new_n5605_), .ZN(new_n5942_));
  NAND2_X1   g05670(.A1(new_n5940_), .A2(new_n5938_), .ZN(new_n5943_));
  NAND3_X1   g05671(.A1(new_n5943_), .A2(new_n5936_), .A3(new_n5942_), .ZN(new_n5944_));
  OAI21_X1   g05672(.A1(new_n5941_), .A2(new_n5936_), .B(new_n5944_), .ZN(\f[40] ));
  XNOR2_X1   g05673(.A1(new_n5617_), .A2(new_n5910_), .ZN(new_n5946_));
  NAND2_X1   g05674(.A1(new_n5936_), .A2(new_n5930_), .ZN(new_n5947_));
  OAI21_X1   g05675(.A1(new_n5947_), .A2(new_n5946_), .B(new_n5942_), .ZN(new_n5948_));
  NAND3_X1   g05676(.A1(new_n5940_), .A2(new_n5948_), .A3(new_n5938_), .ZN(new_n5949_));
  INV_X1     g05677(.I(new_n5884_), .ZN(new_n5950_));
  NAND2_X1   g05678(.A1(new_n5950_), .A2(new_n5889_), .ZN(new_n5951_));
  OAI21_X1   g05679(.A1(new_n5950_), .A2(new_n5889_), .B(new_n5905_), .ZN(new_n5952_));
  NAND2_X1   g05680(.A1(new_n5952_), .A2(new_n5951_), .ZN(new_n5953_));
  AOI21_X1   g05681(.A1(new_n5302_), .A2(new_n5024_), .B(new_n5034_), .ZN(new_n5954_));
  INV_X1     g05682(.I(new_n5575_), .ZN(new_n5955_));
  NOR3_X1    g05683(.A1(new_n5954_), .A2(new_n4807_), .A3(new_n5955_), .ZN(new_n5956_));
  AOI21_X1   g05684(.A1(new_n5562_), .A2(new_n5554_), .B(new_n5561_), .ZN(new_n5957_));
  NOR3_X1    g05685(.A1(new_n5555_), .A2(new_n5384_), .A3(new_n5556_), .ZN(new_n5958_));
  NOR3_X1    g05686(.A1(new_n5958_), .A2(new_n5957_), .A3(new_n5577_), .ZN(new_n5959_));
  NOR2_X1    g05687(.A1(new_n5959_), .A2(new_n5567_), .ZN(new_n5960_));
  AOI21_X1   g05688(.A1(new_n5956_), .A2(new_n5960_), .B(new_n5621_), .ZN(new_n5961_));
  NOR2_X1    g05689(.A1(new_n5385_), .A2(new_n5387_), .ZN(new_n5962_));
  NOR2_X1    g05690(.A1(new_n5629_), .A2(new_n5552_), .ZN(new_n5963_));
  AOI21_X1   g05691(.A1(new_n5962_), .A2(new_n5963_), .B(new_n5626_), .ZN(new_n5964_));
  NAND2_X1   g05692(.A1(new_n5850_), .A2(new_n5838_), .ZN(new_n5965_));
  NAND2_X1   g05693(.A1(new_n5634_), .A2(new_n5839_), .ZN(new_n5966_));
  AOI21_X1   g05694(.A1(new_n5965_), .A2(new_n5966_), .B(new_n5845_), .ZN(new_n5967_));
  INV_X1     g05695(.I(new_n5967_), .ZN(new_n5968_));
  AOI21_X1   g05696(.A1(new_n5806_), .A2(new_n5812_), .B(new_n5817_), .ZN(new_n5969_));
  NAND2_X1   g05697(.A1(new_n5820_), .A2(new_n5805_), .ZN(new_n5970_));
  NAND2_X1   g05698(.A1(new_n5818_), .A2(new_n5804_), .ZN(new_n5971_));
  AOI21_X1   g05699(.A1(new_n5970_), .A2(new_n5971_), .B(new_n5646_), .ZN(new_n5972_));
  NOR2_X1    g05700(.A1(new_n5969_), .A2(new_n5972_), .ZN(new_n5973_));
  XOR2_X1    g05701(.A1(new_n5642_), .A2(new_n5973_), .Z(new_n5974_));
  NOR2_X1    g05702(.A1(new_n5974_), .A2(new_n5835_), .ZN(new_n5975_));
  OAI22_X1   g05703(.A1(new_n1347_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n1344_), .ZN(new_n5976_));
  OAI21_X1   g05704(.A1(new_n1634_), .A2(new_n1457_), .B(new_n5976_), .ZN(new_n5977_));
  AOI21_X1   g05705(.A1(new_n5977_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n5978_));
  XNOR2_X1   g05706(.A1(new_n1940_), .A2(new_n5978_), .ZN(new_n5979_));
  INV_X1     g05707(.I(new_n5979_), .ZN(new_n5980_));
  NOR2_X1    g05708(.A1(new_n5796_), .A2(new_n5807_), .ZN(new_n5981_));
  INV_X1     g05709(.I(new_n5981_), .ZN(new_n5982_));
  NAND2_X1   g05710(.A1(new_n5796_), .A2(new_n5807_), .ZN(new_n5983_));
  AOI21_X1   g05711(.A1(new_n5982_), .A2(new_n5983_), .B(new_n5787_), .ZN(new_n5984_));
  NAND2_X1   g05712(.A1(new_n5759_), .A2(new_n5752_), .ZN(new_n5985_));
  INV_X1     g05713(.I(new_n5652_), .ZN(new_n5986_));
  NAND2_X1   g05714(.A1(new_n5739_), .A2(new_n5738_), .ZN(new_n5987_));
  NAND2_X1   g05715(.A1(new_n5987_), .A2(new_n5986_), .ZN(new_n5988_));
  INV_X1     g05716(.I(new_n5736_), .ZN(new_n5989_));
  AOI21_X1   g05717(.A1(new_n5988_), .A2(new_n5989_), .B(new_n5734_), .ZN(new_n5990_));
  INV_X1     g05718(.I(new_n5686_), .ZN(new_n5991_));
  NOR2_X1    g05719(.A1(new_n5991_), .A2(new_n280_), .ZN(new_n5992_));
  NAND2_X1   g05720(.A1(new_n5689_), .A2(new_n5688_), .ZN(new_n5993_));
  AOI21_X1   g05721(.A1(new_n269_), .A2(new_n490_), .B(new_n5993_), .ZN(new_n5994_));
  NOR2_X1    g05722(.A1(new_n5994_), .A2(new_n5992_), .ZN(new_n5995_));
  XOR2_X1    g05723(.A1(\a[38] ), .A2(\a[41] ), .Z(new_n5996_));
  NAND3_X1   g05724(.A1(new_n5689_), .A2(new_n5427_), .A3(new_n5996_), .ZN(new_n5997_));
  NOR2_X1    g05725(.A1(new_n5997_), .A2(new_n258_), .ZN(new_n5998_));
  INV_X1     g05726(.I(new_n5998_), .ZN(new_n5999_));
  OAI21_X1   g05727(.A1(new_n5995_), .A2(new_n5999_), .B(\a[41] ), .ZN(new_n6000_));
  INV_X1     g05728(.I(new_n6000_), .ZN(new_n6001_));
  NOR3_X1    g05729(.A1(new_n5995_), .A2(\a[41] ), .A3(new_n5999_), .ZN(new_n6002_));
  NOR2_X1    g05730(.A1(new_n6001_), .A2(new_n6002_), .ZN(new_n6003_));
  NOR2_X1    g05731(.A1(new_n5698_), .A2(new_n5693_), .ZN(new_n6004_));
  AND3_X2    g05732(.A1(new_n5110_), .A2(new_n4566_), .A3(new_n5111_), .Z(new_n6005_));
  NAND2_X1   g05733(.A1(new_n4859_), .A2(\b[4] ), .ZN(new_n6006_));
  NAND2_X1   g05734(.A1(new_n4865_), .A2(\b[5] ), .ZN(new_n6007_));
  AOI22_X1   g05735(.A1(new_n6006_), .A2(new_n6007_), .B1(new_n6005_), .B2(\b[3] ), .ZN(new_n6008_));
  OAI21_X1   g05736(.A1(new_n2333_), .A2(new_n5420_), .B(new_n6008_), .ZN(new_n6009_));
  AOI21_X1   g05737(.A1(new_n6004_), .A2(new_n5695_), .B(new_n6009_), .ZN(new_n6010_));
  NAND3_X1   g05738(.A1(new_n5694_), .A2(new_n5692_), .A3(new_n5695_), .ZN(new_n6011_));
  NOR2_X1    g05739(.A1(new_n5420_), .A2(new_n325_), .ZN(new_n6012_));
  NOR2_X1    g05740(.A1(new_n5107_), .A2(new_n419_), .ZN(new_n6013_));
  OAI22_X1   g05741(.A1(new_n6012_), .A2(new_n6013_), .B1(new_n298_), .B2(new_n5112_), .ZN(new_n6014_));
  AOI21_X1   g05742(.A1(new_n378_), .A2(new_n4859_), .B(new_n6014_), .ZN(new_n6015_));
  NOR2_X1    g05743(.A1(new_n6011_), .A2(new_n6015_), .ZN(new_n6016_));
  OAI21_X1   g05744(.A1(new_n6010_), .A2(new_n6016_), .B(new_n6003_), .ZN(new_n6017_));
  INV_X1     g05745(.I(new_n6002_), .ZN(new_n6018_));
  NAND2_X1   g05746(.A1(new_n6018_), .A2(new_n6000_), .ZN(new_n6019_));
  NAND2_X1   g05747(.A1(new_n6011_), .A2(new_n6015_), .ZN(new_n6020_));
  NAND4_X1   g05748(.A1(new_n6009_), .A2(new_n5692_), .A3(new_n5694_), .A4(new_n5695_), .ZN(new_n6021_));
  NAND3_X1   g05749(.A1(new_n6020_), .A2(new_n6019_), .A3(new_n6021_), .ZN(new_n6022_));
  AOI21_X1   g05750(.A1(new_n6017_), .A2(new_n6022_), .B(\a[38] ), .ZN(new_n6023_));
  AOI21_X1   g05751(.A1(new_n6020_), .A2(new_n6021_), .B(new_n6019_), .ZN(new_n6024_));
  NOR3_X1    g05752(.A1(new_n6010_), .A2(new_n6016_), .A3(new_n6003_), .ZN(new_n6025_));
  NOR3_X1    g05753(.A1(new_n6025_), .A2(new_n6024_), .A3(new_n4860_), .ZN(new_n6026_));
  OAI21_X1   g05754(.A1(new_n6026_), .A2(new_n6023_), .B(new_n5720_), .ZN(new_n6027_));
  NOR2_X1    g05755(.A1(new_n6027_), .A2(new_n5702_), .ZN(new_n6028_));
  OAI21_X1   g05756(.A1(new_n6025_), .A2(new_n6024_), .B(new_n4860_), .ZN(new_n6029_));
  NAND3_X1   g05757(.A1(new_n6017_), .A2(new_n6022_), .A3(\a[38] ), .ZN(new_n6030_));
  NAND2_X1   g05758(.A1(new_n6029_), .A2(new_n6030_), .ZN(new_n6031_));
  NAND2_X1   g05759(.A1(new_n5709_), .A2(new_n5700_), .ZN(new_n6033_));
  INV_X1     g05760(.I(new_n6033_), .ZN(new_n6034_));
  OAI21_X1   g05761(.A1(new_n6028_), .A2(new_n6034_), .B(new_n5719_), .ZN(new_n6035_));
  NAND3_X1   g05762(.A1(new_n6031_), .A2(new_n5703_), .A3(new_n5720_), .ZN(new_n6036_));
  NAND3_X1   g05763(.A1(new_n6036_), .A2(new_n5706_), .A3(new_n6033_), .ZN(new_n6037_));
  OAI22_X1   g05764(.A1(new_n4072_), .A2(new_n472_), .B1(new_n515_), .B2(new_n4067_), .ZN(new_n6038_));
  OAI21_X1   g05765(.A1(new_n420_), .A2(new_n4318_), .B(new_n6038_), .ZN(new_n6039_));
  AOI21_X1   g05766(.A1(new_n6039_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n6040_));
  XOR2_X1    g05767(.A1(new_n700_), .A2(new_n6040_), .Z(new_n6041_));
  INV_X1     g05768(.I(new_n6041_), .ZN(new_n6042_));
  NAND3_X1   g05769(.A1(new_n6035_), .A2(new_n6037_), .A3(new_n6042_), .ZN(new_n6043_));
  AOI21_X1   g05770(.A1(new_n6036_), .A2(new_n6033_), .B(new_n5706_), .ZN(new_n6044_));
  NOR3_X1    g05771(.A1(new_n6028_), .A2(new_n5719_), .A3(new_n6034_), .ZN(new_n6045_));
  OAI21_X1   g05772(.A1(new_n6045_), .A2(new_n6044_), .B(new_n6041_), .ZN(new_n6046_));
  NAND2_X1   g05773(.A1(new_n6046_), .A2(new_n6043_), .ZN(new_n6047_));
  NAND3_X1   g05774(.A1(new_n6047_), .A2(new_n5717_), .A3(new_n5727_), .ZN(new_n6048_));
  NOR2_X1    g05775(.A1(new_n5711_), .A2(new_n5705_), .ZN(new_n6049_));
  NOR2_X1    g05776(.A1(new_n6049_), .A2(new_n5715_), .ZN(new_n6051_));
  INV_X1     g05777(.I(new_n6051_), .ZN(new_n6052_));
  AOI21_X1   g05778(.A1(new_n6048_), .A2(new_n6052_), .B(new_n5664_), .ZN(new_n6053_));
  INV_X1     g05779(.I(new_n5664_), .ZN(new_n6054_));
  INV_X1     g05780(.I(new_n5717_), .ZN(new_n6055_));
  NOR3_X1    g05781(.A1(new_n6045_), .A2(new_n6044_), .A3(new_n6041_), .ZN(new_n6056_));
  AOI21_X1   g05782(.A1(new_n6035_), .A2(new_n6037_), .B(new_n6042_), .ZN(new_n6057_));
  OAI21_X1   g05783(.A1(new_n6056_), .A2(new_n6057_), .B(new_n5727_), .ZN(new_n6058_));
  NOR2_X1    g05784(.A1(new_n6058_), .A2(new_n6055_), .ZN(new_n6059_));
  NOR3_X1    g05785(.A1(new_n6059_), .A2(new_n6054_), .A3(new_n6051_), .ZN(new_n6060_));
  OAI22_X1   g05786(.A1(new_n656_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n706_), .ZN(new_n6061_));
  OAI21_X1   g05787(.A1(new_n565_), .A2(new_n3569_), .B(new_n6061_), .ZN(new_n6062_));
  AOI21_X1   g05788(.A1(new_n6062_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n6063_));
  XNOR2_X1   g05789(.A1(new_n710_), .A2(new_n6063_), .ZN(new_n6064_));
  NOR3_X1    g05790(.A1(new_n6060_), .A2(new_n6053_), .A3(new_n6064_), .ZN(new_n6065_));
  OAI21_X1   g05791(.A1(new_n6059_), .A2(new_n6051_), .B(new_n6054_), .ZN(new_n6066_));
  NAND3_X1   g05792(.A1(new_n6048_), .A2(new_n5664_), .A3(new_n6052_), .ZN(new_n6067_));
  INV_X1     g05793(.I(new_n6064_), .ZN(new_n6068_));
  AOI21_X1   g05794(.A1(new_n6066_), .A2(new_n6067_), .B(new_n6068_), .ZN(new_n6069_));
  OAI22_X1   g05795(.A1(new_n861_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n930_), .ZN(new_n6070_));
  OAI21_X1   g05796(.A1(new_n780_), .A2(new_n2884_), .B(new_n6070_), .ZN(new_n6071_));
  AOI21_X1   g05797(.A1(new_n6071_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n6072_));
  XNOR2_X1   g05798(.A1(new_n937_), .A2(new_n6072_), .ZN(new_n6073_));
  INV_X1     g05799(.I(new_n6073_), .ZN(new_n6074_));
  OAI21_X1   g05800(.A1(new_n6065_), .A2(new_n6069_), .B(new_n6074_), .ZN(new_n6075_));
  NAND3_X1   g05801(.A1(new_n6066_), .A2(new_n6067_), .A3(new_n6068_), .ZN(new_n6076_));
  OAI21_X1   g05802(.A1(new_n6060_), .A2(new_n6053_), .B(new_n6064_), .ZN(new_n6077_));
  NAND3_X1   g05803(.A1(new_n6077_), .A2(new_n6076_), .A3(new_n6073_), .ZN(new_n6078_));
  AOI21_X1   g05804(.A1(new_n6075_), .A2(new_n6078_), .B(new_n5990_), .ZN(new_n6079_));
  INV_X1     g05805(.I(new_n5734_), .ZN(new_n6080_));
  OAI21_X1   g05806(.A1(new_n5740_), .A2(new_n5736_), .B(new_n6080_), .ZN(new_n6081_));
  NAND3_X1   g05807(.A1(new_n6077_), .A2(new_n6076_), .A3(new_n6074_), .ZN(new_n6082_));
  OAI21_X1   g05808(.A1(new_n6065_), .A2(new_n6069_), .B(new_n6073_), .ZN(new_n6083_));
  AOI21_X1   g05809(.A1(new_n6083_), .A2(new_n6082_), .B(new_n6081_), .ZN(new_n6084_));
  OAI21_X1   g05810(.A1(new_n6079_), .A2(new_n6084_), .B(new_n5985_), .ZN(new_n6085_));
  NOR2_X1    g05811(.A1(new_n6085_), .A2(new_n5762_), .ZN(new_n6086_));
  AOI21_X1   g05812(.A1(new_n6077_), .A2(new_n6076_), .B(new_n6073_), .ZN(new_n6087_));
  NOR3_X1    g05813(.A1(new_n6065_), .A2(new_n6069_), .A3(new_n6074_), .ZN(new_n6088_));
  OAI21_X1   g05814(.A1(new_n6088_), .A2(new_n6087_), .B(new_n6081_), .ZN(new_n6089_));
  NOR3_X1    g05815(.A1(new_n6065_), .A2(new_n6069_), .A3(new_n6073_), .ZN(new_n6090_));
  AOI21_X1   g05816(.A1(new_n6077_), .A2(new_n6076_), .B(new_n6074_), .ZN(new_n6091_));
  OAI21_X1   g05817(.A1(new_n6090_), .A2(new_n6091_), .B(new_n5990_), .ZN(new_n6092_));
  NAND2_X1   g05818(.A1(new_n6092_), .A2(new_n6089_), .ZN(new_n6093_));
  NOR2_X1    g05819(.A1(new_n5761_), .A2(new_n5750_), .ZN(new_n6095_));
  OAI21_X1   g05820(.A1(new_n6086_), .A2(new_n6095_), .B(new_n5651_), .ZN(new_n6096_));
  NAND2_X1   g05821(.A1(new_n5648_), .A2(new_n5191_), .ZN(new_n6097_));
  NAND2_X1   g05822(.A1(new_n5650_), .A2(new_n5647_), .ZN(new_n6098_));
  NAND2_X1   g05823(.A1(new_n6098_), .A2(new_n6097_), .ZN(new_n6099_));
  NAND3_X1   g05824(.A1(new_n6093_), .A2(new_n5763_), .A3(new_n5985_), .ZN(new_n6100_));
  INV_X1     g05825(.I(new_n6095_), .ZN(new_n6101_));
  NAND3_X1   g05826(.A1(new_n6100_), .A2(new_n6099_), .A3(new_n6101_), .ZN(new_n6102_));
  OAI22_X1   g05827(.A1(new_n2171_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n2166_), .ZN(new_n6103_));
  OAI21_X1   g05828(.A1(new_n1017_), .A2(new_n2322_), .B(new_n6103_), .ZN(new_n6104_));
  AOI21_X1   g05829(.A1(new_n6104_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n6105_));
  XNOR2_X1   g05830(.A1(new_n1196_), .A2(new_n6105_), .ZN(new_n6106_));
  AOI21_X1   g05831(.A1(new_n6096_), .A2(new_n6102_), .B(new_n6106_), .ZN(new_n6107_));
  AOI21_X1   g05832(.A1(new_n6100_), .A2(new_n6101_), .B(new_n6099_), .ZN(new_n6108_));
  NOR3_X1    g05833(.A1(new_n6086_), .A2(new_n5651_), .A3(new_n6095_), .ZN(new_n6109_));
  INV_X1     g05834(.I(new_n6106_), .ZN(new_n6110_));
  NOR3_X1    g05835(.A1(new_n6109_), .A2(new_n6108_), .A3(new_n6110_), .ZN(new_n6111_));
  NOR3_X1    g05836(.A1(new_n6111_), .A2(new_n6107_), .A3(new_n5775_), .ZN(new_n6112_));
  NOR3_X1    g05837(.A1(new_n6112_), .A2(new_n5807_), .A3(new_n5796_), .ZN(new_n6113_));
  OAI21_X1   g05838(.A1(new_n6109_), .A2(new_n6108_), .B(new_n6110_), .ZN(new_n6114_));
  NAND3_X1   g05839(.A1(new_n6096_), .A2(new_n6102_), .A3(new_n6106_), .ZN(new_n6115_));
  NAND3_X1   g05840(.A1(new_n6114_), .A2(new_n6115_), .A3(new_n5795_), .ZN(new_n6116_));
  AOI21_X1   g05841(.A1(new_n6116_), .A2(new_n5782_), .B(new_n5776_), .ZN(new_n6117_));
  OAI22_X1   g05842(.A1(new_n1712_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n1707_), .ZN(new_n6118_));
  OAI21_X1   g05843(.A1(new_n1294_), .A2(new_n1850_), .B(new_n6118_), .ZN(new_n6119_));
  AOI21_X1   g05844(.A1(new_n6119_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n6120_));
  XOR2_X1    g05845(.A1(new_n1530_), .A2(new_n6120_), .Z(new_n6121_));
  NOR3_X1    g05846(.A1(new_n6113_), .A2(new_n6117_), .A3(new_n6121_), .ZN(new_n6122_));
  NAND3_X1   g05847(.A1(new_n6116_), .A2(new_n5782_), .A3(new_n5776_), .ZN(new_n6123_));
  OAI21_X1   g05848(.A1(new_n6112_), .A2(new_n5807_), .B(new_n5796_), .ZN(new_n6124_));
  INV_X1     g05849(.I(new_n6121_), .ZN(new_n6125_));
  AOI21_X1   g05850(.A1(new_n6124_), .A2(new_n6123_), .B(new_n6125_), .ZN(new_n6126_));
  NOR3_X1    g05851(.A1(new_n5984_), .A2(new_n6122_), .A3(new_n6126_), .ZN(new_n6127_));
  NOR3_X1    g05852(.A1(new_n6127_), .A2(new_n5646_), .A3(new_n5820_), .ZN(new_n6128_));
  INV_X1     g05853(.I(new_n5983_), .ZN(new_n6129_));
  OAI21_X1   g05854(.A1(new_n6129_), .A2(new_n5981_), .B(new_n5786_), .ZN(new_n6130_));
  NAND3_X1   g05855(.A1(new_n6124_), .A2(new_n6123_), .A3(new_n6125_), .ZN(new_n6131_));
  OAI21_X1   g05856(.A1(new_n6113_), .A2(new_n6117_), .B(new_n6121_), .ZN(new_n6132_));
  NAND3_X1   g05857(.A1(new_n6130_), .A2(new_n6132_), .A3(new_n6131_), .ZN(new_n6133_));
  AOI21_X1   g05858(.A1(new_n6133_), .A2(new_n5818_), .B(new_n5817_), .ZN(new_n6134_));
  NOR2_X1    g05859(.A1(new_n6134_), .A2(new_n6128_), .ZN(new_n6135_));
  NOR2_X1    g05860(.A1(new_n5646_), .A2(new_n5820_), .ZN(new_n6136_));
  NOR2_X1    g05861(.A1(new_n5817_), .A2(new_n5818_), .ZN(new_n6137_));
  OAI21_X1   g05862(.A1(new_n6137_), .A2(new_n6136_), .B(new_n5804_), .ZN(new_n6138_));
  NAND3_X1   g05863(.A1(new_n5641_), .A2(new_n5636_), .A3(new_n5973_), .ZN(new_n6139_));
  OAI22_X1   g05864(.A1(new_n1055_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n1061_), .ZN(new_n6140_));
  OAI21_X1   g05865(.A1(new_n2102_), .A2(new_n1332_), .B(new_n6140_), .ZN(new_n6141_));
  AOI21_X1   g05866(.A1(new_n6141_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n6142_));
  XNOR2_X1   g05867(.A1(new_n2443_), .A2(new_n6142_), .ZN(new_n6143_));
  AOI21_X1   g05868(.A1(new_n6139_), .A2(new_n6138_), .B(new_n6143_), .ZN(new_n6144_));
  INV_X1     g05869(.I(new_n6138_), .ZN(new_n6145_));
  NOR3_X1    g05870(.A1(new_n5833_), .A2(new_n5635_), .A3(new_n5823_), .ZN(new_n6146_));
  INV_X1     g05871(.I(new_n6143_), .ZN(new_n6147_));
  NOR3_X1    g05872(.A1(new_n6146_), .A2(new_n6145_), .A3(new_n6147_), .ZN(new_n6148_));
  OAI21_X1   g05873(.A1(new_n6148_), .A2(new_n6144_), .B(new_n6135_), .ZN(new_n6149_));
  INV_X1     g05874(.I(new_n6135_), .ZN(new_n6150_));
  OAI21_X1   g05875(.A1(new_n6146_), .A2(new_n6145_), .B(new_n6147_), .ZN(new_n6151_));
  NAND3_X1   g05876(.A1(new_n6139_), .A2(new_n6138_), .A3(new_n6143_), .ZN(new_n6152_));
  NAND3_X1   g05877(.A1(new_n6151_), .A2(new_n6152_), .A3(new_n6150_), .ZN(new_n6153_));
  AOI21_X1   g05878(.A1(new_n6149_), .A2(new_n6153_), .B(new_n5980_), .ZN(new_n6154_));
  AOI21_X1   g05879(.A1(new_n6151_), .A2(new_n6152_), .B(new_n6150_), .ZN(new_n6155_));
  NOR3_X1    g05880(.A1(new_n6148_), .A2(new_n6144_), .A3(new_n6135_), .ZN(new_n6156_));
  NOR3_X1    g05881(.A1(new_n6156_), .A2(new_n6155_), .A3(new_n5979_), .ZN(new_n6157_));
  NOR3_X1    g05882(.A1(new_n6157_), .A2(new_n6154_), .A3(new_n5975_), .ZN(new_n6158_));
  NOR3_X1    g05883(.A1(new_n6158_), .A2(new_n5634_), .A3(new_n5839_), .ZN(new_n6159_));
  XOR2_X1    g05884(.A1(new_n5642_), .A2(new_n5823_), .Z(new_n6160_));
  NAND2_X1   g05885(.A1(new_n6160_), .A2(new_n5827_), .ZN(new_n6161_));
  OAI21_X1   g05886(.A1(new_n6156_), .A2(new_n6155_), .B(new_n5979_), .ZN(new_n6162_));
  NAND3_X1   g05887(.A1(new_n6149_), .A2(new_n6153_), .A3(new_n5980_), .ZN(new_n6163_));
  NAND3_X1   g05888(.A1(new_n6162_), .A2(new_n6163_), .A3(new_n6161_), .ZN(new_n6164_));
  AOI21_X1   g05889(.A1(new_n6164_), .A2(new_n5838_), .B(new_n5850_), .ZN(new_n6165_));
  OAI22_X1   g05890(.A1(new_n970_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n820_), .ZN(new_n6166_));
  OAI21_X1   g05891(.A1(new_n2643_), .A2(new_n894_), .B(new_n6166_), .ZN(new_n6167_));
  AOI21_X1   g05892(.A1(new_n6167_), .A2(new_n827_), .B(new_n970_), .ZN(new_n6168_));
  XNOR2_X1   g05893(.A1(new_n3022_), .A2(new_n6168_), .ZN(new_n6169_));
  INV_X1     g05894(.I(new_n6169_), .ZN(new_n6170_));
  OAI21_X1   g05895(.A1(new_n6159_), .A2(new_n6165_), .B(new_n6170_), .ZN(new_n6171_));
  NAND3_X1   g05896(.A1(new_n6164_), .A2(new_n5850_), .A3(new_n5838_), .ZN(new_n6172_));
  OAI21_X1   g05897(.A1(new_n6158_), .A2(new_n5839_), .B(new_n5634_), .ZN(new_n6173_));
  NAND3_X1   g05898(.A1(new_n6173_), .A2(new_n6172_), .A3(new_n6169_), .ZN(new_n6174_));
  NAND3_X1   g05899(.A1(new_n6171_), .A2(new_n6174_), .A3(new_n5968_), .ZN(new_n6175_));
  NAND3_X1   g05900(.A1(new_n6175_), .A2(new_n5964_), .A3(new_n5854_), .ZN(new_n6176_));
  NAND2_X1   g05901(.A1(new_n5863_), .A2(new_n5856_), .ZN(new_n6177_));
  AOI21_X1   g05902(.A1(new_n6173_), .A2(new_n6172_), .B(new_n6169_), .ZN(new_n6178_));
  NOR3_X1    g05903(.A1(new_n6159_), .A2(new_n6165_), .A3(new_n6170_), .ZN(new_n6179_));
  NOR3_X1    g05904(.A1(new_n6179_), .A2(new_n6178_), .A3(new_n5967_), .ZN(new_n6180_));
  OAI21_X1   g05905(.A1(new_n6180_), .A2(new_n5866_), .B(new_n6177_), .ZN(new_n6181_));
  OAI22_X1   g05906(.A1(new_n607_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n610_), .ZN(new_n6182_));
  OAI21_X1   g05907(.A1(new_n3260_), .A2(new_n684_), .B(new_n6182_), .ZN(new_n6183_));
  AOI21_X1   g05908(.A1(new_n6183_), .A2(new_n612_), .B(new_n607_), .ZN(new_n6184_));
  XOR2_X1    g05909(.A1(new_n3722_), .A2(new_n6184_), .Z(new_n6185_));
  AOI21_X1   g05910(.A1(new_n6181_), .A2(new_n6176_), .B(new_n6185_), .ZN(new_n6186_));
  NOR3_X1    g05911(.A1(new_n6180_), .A2(new_n6177_), .A3(new_n5866_), .ZN(new_n6187_));
  AOI21_X1   g05912(.A1(new_n6175_), .A2(new_n5854_), .B(new_n5964_), .ZN(new_n6188_));
  INV_X1     g05913(.I(new_n6185_), .ZN(new_n6189_));
  NOR3_X1    g05914(.A1(new_n6187_), .A2(new_n6188_), .A3(new_n6189_), .ZN(new_n6190_));
  OAI21_X1   g05915(.A1(new_n6190_), .A2(new_n6186_), .B(new_n5877_), .ZN(new_n6191_));
  NOR2_X1    g05916(.A1(new_n6191_), .A2(new_n5880_), .ZN(new_n6192_));
  OAI21_X1   g05917(.A1(new_n6187_), .A2(new_n6188_), .B(new_n6189_), .ZN(new_n6193_));
  NAND3_X1   g05918(.A1(new_n6181_), .A2(new_n6176_), .A3(new_n6185_), .ZN(new_n6194_));
  NAND2_X1   g05919(.A1(new_n6193_), .A2(new_n6194_), .ZN(new_n6195_));
  NOR2_X1    g05920(.A1(new_n5879_), .A2(new_n5871_), .ZN(new_n6197_));
  OAI21_X1   g05921(.A1(new_n6192_), .A2(new_n6197_), .B(new_n5961_), .ZN(new_n6198_));
  INV_X1     g05922(.I(new_n5880_), .ZN(new_n6199_));
  NAND3_X1   g05923(.A1(new_n6195_), .A2(new_n5877_), .A3(new_n6199_), .ZN(new_n6200_));
  INV_X1     g05924(.I(new_n6197_), .ZN(new_n6201_));
  NAND3_X1   g05925(.A1(new_n6200_), .A2(new_n5625_), .A3(new_n6201_), .ZN(new_n6202_));
  OAI22_X1   g05926(.A1(new_n448_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n450_), .ZN(new_n6203_));
  OAI21_X1   g05927(.A1(new_n3989_), .A2(new_n496_), .B(new_n6203_), .ZN(new_n6204_));
  AOI21_X1   g05928(.A1(new_n6204_), .A2(new_n452_), .B(new_n448_), .ZN(new_n6205_));
  XOR2_X1    g05929(.A1(new_n4499_), .A2(new_n6205_), .Z(new_n6206_));
  INV_X1     g05930(.I(new_n6206_), .ZN(new_n6207_));
  NAND3_X1   g05931(.A1(new_n6198_), .A2(new_n6202_), .A3(new_n6207_), .ZN(new_n6208_));
  AOI21_X1   g05932(.A1(new_n6200_), .A2(new_n6201_), .B(new_n5625_), .ZN(new_n6209_));
  NOR3_X1    g05933(.A1(new_n6192_), .A2(new_n5961_), .A3(new_n6197_), .ZN(new_n6210_));
  OAI21_X1   g05934(.A1(new_n6210_), .A2(new_n6209_), .B(new_n6206_), .ZN(new_n6211_));
  NAND2_X1   g05935(.A1(new_n6211_), .A2(new_n6208_), .ZN(new_n6212_));
  OAI22_X1   g05936(.A1(new_n5068_), .A2(new_n341_), .B1(new_n404_), .B2(new_n5353_), .ZN(new_n6213_));
  OAI21_X1   g05937(.A1(new_n4774_), .A2(new_n366_), .B(new_n6213_), .ZN(new_n6214_));
  AOI21_X1   g05938(.A1(new_n6214_), .A2(new_n334_), .B(new_n341_), .ZN(new_n6215_));
  XNOR2_X1   g05939(.A1(new_n5357_), .A2(new_n6215_), .ZN(new_n6216_));
  INV_X1     g05940(.I(new_n6216_), .ZN(new_n6217_));
  XOR2_X1    g05941(.A1(new_n6212_), .A2(new_n6217_), .Z(new_n6218_));
  NAND2_X1   g05942(.A1(new_n5953_), .A2(new_n6218_), .ZN(new_n6219_));
  XOR2_X1    g05943(.A1(new_n6212_), .A2(new_n6217_), .Z(new_n6220_));
  OAI21_X1   g05944(.A1(new_n5953_), .A2(new_n6220_), .B(new_n6219_), .ZN(new_n6221_));
  OAI21_X1   g05945(.A1(new_n5899_), .A2(new_n5908_), .B(new_n5615_), .ZN(new_n6222_));
  NAND2_X1   g05946(.A1(new_n6222_), .A2(new_n5614_), .ZN(new_n6223_));
  NAND3_X1   g05947(.A1(new_n5900_), .A2(new_n5909_), .A3(new_n5596_), .ZN(new_n6224_));
  NAND3_X1   g05948(.A1(new_n5371_), .A2(new_n6223_), .A3(new_n6224_), .ZN(new_n6225_));
  XOR2_X1    g05949(.A1(new_n5620_), .A2(new_n5890_), .Z(new_n6226_));
  OAI21_X1   g05950(.A1(new_n5895_), .A2(new_n6226_), .B(new_n6225_), .ZN(new_n6227_));
  XOR2_X1    g05951(.A1(new_n6227_), .A2(new_n6221_), .Z(new_n6228_));
  INV_X1     g05952(.I(\b[41] ), .ZN(new_n6229_));
  NOR2_X1    g05953(.A1(new_n6229_), .A2(\b[39] ), .ZN(new_n6230_));
  NOR2_X1    g05954(.A1(new_n5913_), .A2(\b[41] ), .ZN(new_n6231_));
  OAI21_X1   g05955(.A1(new_n6230_), .A2(new_n6231_), .B(new_n5920_), .ZN(new_n6232_));
  XNOR2_X1   g05956(.A1(new_n5917_), .A2(new_n6232_), .ZN(new_n6233_));
  OAI22_X1   g05957(.A1(new_n330_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n263_), .ZN(new_n6234_));
  OAI21_X1   g05958(.A1(new_n5913_), .A2(new_n289_), .B(new_n6234_), .ZN(new_n6235_));
  AOI21_X1   g05959(.A1(new_n6235_), .A2(new_n260_), .B(new_n426_), .ZN(new_n6236_));
  XOR2_X1    g05960(.A1(new_n6233_), .A2(new_n6236_), .Z(new_n6237_));
  INV_X1     g05961(.I(new_n6237_), .ZN(new_n6238_));
  XOR2_X1    g05962(.A1(new_n6228_), .A2(new_n6238_), .Z(new_n6239_));
  XOR2_X1    g05963(.A1(new_n6228_), .A2(new_n6238_), .Z(new_n6240_));
  NAND2_X1   g05964(.A1(new_n5949_), .A2(new_n6240_), .ZN(new_n6241_));
  OAI21_X1   g05965(.A1(new_n5949_), .A2(new_n6239_), .B(new_n6241_), .ZN(\f[41] ));
  NAND2_X1   g05966(.A1(new_n6228_), .A2(new_n6238_), .ZN(new_n6243_));
  OAI22_X1   g05967(.A1(new_n5353_), .A2(new_n341_), .B1(new_n404_), .B2(new_n5913_), .ZN(new_n6244_));
  OAI21_X1   g05968(.A1(new_n5068_), .A2(new_n366_), .B(new_n6244_), .ZN(new_n6245_));
  AOI21_X1   g05969(.A1(new_n6245_), .A2(new_n334_), .B(new_n341_), .ZN(new_n6246_));
  XNOR2_X1   g05970(.A1(new_n5600_), .A2(new_n6246_), .ZN(new_n6247_));
  INV_X1     g05971(.I(new_n6247_), .ZN(new_n6248_));
  AOI21_X1   g05972(.A1(new_n6198_), .A2(new_n6202_), .B(new_n6207_), .ZN(new_n6249_));
  NOR3_X1    g05973(.A1(new_n6210_), .A2(new_n6209_), .A3(new_n6206_), .ZN(new_n6250_));
  OAI21_X1   g05974(.A1(new_n6250_), .A2(new_n6249_), .B(new_n5884_), .ZN(new_n6251_));
  NAND2_X1   g05975(.A1(new_n6251_), .A2(new_n5888_), .ZN(new_n6252_));
  NAND3_X1   g05976(.A1(new_n5950_), .A2(new_n6208_), .A3(new_n6211_), .ZN(new_n6253_));
  NAND3_X1   g05977(.A1(new_n6252_), .A2(new_n5905_), .A3(new_n6253_), .ZN(new_n6254_));
  AOI21_X1   g05978(.A1(new_n6181_), .A2(new_n6176_), .B(new_n6189_), .ZN(new_n6255_));
  INV_X1     g05979(.I(new_n6255_), .ZN(new_n6256_));
  AOI21_X1   g05980(.A1(new_n6195_), .A2(new_n5872_), .B(new_n5881_), .ZN(new_n6257_));
  NOR2_X1    g05981(.A1(new_n6195_), .A2(new_n5872_), .ZN(new_n6258_));
  NOR3_X1    g05982(.A1(new_n6257_), .A2(new_n6258_), .A3(new_n5961_), .ZN(new_n6259_));
  AOI21_X1   g05983(.A1(new_n6173_), .A2(new_n6172_), .B(new_n6170_), .ZN(new_n6260_));
  OAI21_X1   g05984(.A1(new_n6179_), .A2(new_n6178_), .B(new_n5967_), .ZN(new_n6261_));
  AOI21_X1   g05985(.A1(new_n6261_), .A2(new_n5866_), .B(new_n5964_), .ZN(new_n6262_));
  NOR2_X1    g05986(.A1(new_n6146_), .A2(new_n6145_), .ZN(new_n6263_));
  NOR2_X1    g05987(.A1(new_n6263_), .A2(new_n6135_), .ZN(new_n6264_));
  NAND2_X1   g05988(.A1(new_n6139_), .A2(new_n6138_), .ZN(new_n6265_));
  NOR2_X1    g05989(.A1(new_n6265_), .A2(new_n6150_), .ZN(new_n6266_));
  OAI21_X1   g05990(.A1(new_n6264_), .A2(new_n6266_), .B(new_n5979_), .ZN(new_n6267_));
  NAND2_X1   g05991(.A1(new_n6265_), .A2(new_n6150_), .ZN(new_n6268_));
  NAND2_X1   g05992(.A1(new_n6263_), .A2(new_n6135_), .ZN(new_n6269_));
  NAND3_X1   g05993(.A1(new_n6269_), .A2(new_n6268_), .A3(new_n5980_), .ZN(new_n6270_));
  AOI21_X1   g05994(.A1(new_n6267_), .A2(new_n6270_), .B(new_n6143_), .ZN(new_n6271_));
  AOI21_X1   g05995(.A1(new_n6162_), .A2(new_n6163_), .B(new_n6161_), .ZN(new_n6272_));
  OAI21_X1   g05996(.A1(new_n6272_), .A2(new_n5838_), .B(new_n5634_), .ZN(new_n6273_));
  NOR2_X1    g05997(.A1(new_n6135_), .A2(new_n5980_), .ZN(new_n6274_));
  OAI21_X1   g05998(.A1(new_n6134_), .A2(new_n6128_), .B(new_n5980_), .ZN(new_n6275_));
  NAND3_X1   g05999(.A1(new_n6133_), .A2(new_n5817_), .A3(new_n5818_), .ZN(new_n6276_));
  OAI21_X1   g06000(.A1(new_n6127_), .A2(new_n5820_), .B(new_n5646_), .ZN(new_n6277_));
  NAND3_X1   g06001(.A1(new_n6277_), .A2(new_n6276_), .A3(new_n5979_), .ZN(new_n6278_));
  AOI21_X1   g06002(.A1(new_n6275_), .A2(new_n6278_), .B(new_n6138_), .ZN(new_n6279_));
  OAI21_X1   g06003(.A1(new_n6279_), .A2(new_n5823_), .B(new_n5642_), .ZN(new_n6280_));
  OAI21_X1   g06004(.A1(new_n6122_), .A2(new_n6126_), .B(new_n5984_), .ZN(new_n6281_));
  AOI21_X1   g06005(.A1(new_n6281_), .A2(new_n5820_), .B(new_n5817_), .ZN(new_n6282_));
  OAI21_X1   g06006(.A1(new_n6109_), .A2(new_n6108_), .B(new_n6106_), .ZN(new_n6283_));
  OAI21_X1   g06007(.A1(new_n6111_), .A2(new_n6107_), .B(new_n5775_), .ZN(new_n6284_));
  AOI21_X1   g06008(.A1(new_n6284_), .A2(new_n5807_), .B(new_n5776_), .ZN(new_n6285_));
  NAND2_X1   g06009(.A1(new_n6077_), .A2(new_n6076_), .ZN(new_n6286_));
  NAND2_X1   g06010(.A1(new_n6081_), .A2(new_n6286_), .ZN(new_n6287_));
  NAND3_X1   g06011(.A1(new_n5990_), .A2(new_n6076_), .A3(new_n6077_), .ZN(new_n6288_));
  AOI21_X1   g06012(.A1(new_n6288_), .A2(new_n6287_), .B(new_n6074_), .ZN(new_n6289_));
  OAI21_X1   g06013(.A1(new_n6079_), .A2(new_n6084_), .B(new_n5751_), .ZN(new_n6290_));
  NAND2_X1   g06014(.A1(new_n6290_), .A2(new_n5761_), .ZN(new_n6291_));
  NAND3_X1   g06015(.A1(new_n6092_), .A2(new_n6089_), .A3(new_n5750_), .ZN(new_n6292_));
  NAND3_X1   g06016(.A1(new_n6291_), .A2(new_n6099_), .A3(new_n6292_), .ZN(new_n6293_));
  NOR3_X1    g06017(.A1(new_n6060_), .A2(new_n6053_), .A3(new_n6068_), .ZN(new_n6294_));
  INV_X1     g06018(.I(new_n6294_), .ZN(new_n6295_));
  OAI21_X1   g06019(.A1(new_n6065_), .A2(new_n6069_), .B(new_n5729_), .ZN(new_n6296_));
  NAND2_X1   g06020(.A1(new_n6296_), .A2(new_n5733_), .ZN(new_n6297_));
  NOR3_X1    g06021(.A1(new_n6065_), .A2(new_n6069_), .A3(new_n5729_), .ZN(new_n6298_));
  NOR2_X1    g06022(.A1(new_n6298_), .A2(new_n5740_), .ZN(new_n6299_));
  INV_X1     g06023(.I(new_n6049_), .ZN(new_n6300_));
  OAI21_X1   g06024(.A1(new_n6056_), .A2(new_n6057_), .B(new_n6300_), .ZN(new_n6301_));
  NAND2_X1   g06025(.A1(new_n6301_), .A2(new_n5715_), .ZN(new_n6302_));
  NAND3_X1   g06026(.A1(new_n6046_), .A2(new_n6043_), .A3(new_n6049_), .ZN(new_n6303_));
  NAND3_X1   g06027(.A1(new_n6302_), .A2(new_n5664_), .A3(new_n6303_), .ZN(new_n6304_));
  XOR2_X1    g06028(.A1(new_n6015_), .A2(new_n4860_), .Z(new_n6305_));
  NAND2_X1   g06029(.A1(new_n6019_), .A2(new_n6011_), .ZN(new_n6306_));
  INV_X1     g06030(.I(new_n6011_), .ZN(new_n6307_));
  NAND2_X1   g06031(.A1(new_n6003_), .A2(new_n6307_), .ZN(new_n6308_));
  AOI21_X1   g06032(.A1(new_n6308_), .A2(new_n6306_), .B(new_n6305_), .ZN(new_n6309_));
  INV_X1     g06033(.I(new_n6309_), .ZN(new_n6310_));
  AOI21_X1   g06034(.A1(new_n6031_), .A2(new_n5700_), .B(new_n5709_), .ZN(new_n6311_));
  OAI21_X1   g06035(.A1(new_n6031_), .A2(new_n5700_), .B(new_n5706_), .ZN(new_n6312_));
  NOR2_X1    g06036(.A1(new_n6311_), .A2(new_n6312_), .ZN(new_n6313_));
  NOR2_X1    g06037(.A1(new_n5997_), .A2(new_n269_), .ZN(new_n6314_));
  OAI22_X1   g06038(.A1(new_n298_), .A2(new_n5991_), .B1(new_n5993_), .B2(new_n280_), .ZN(new_n6315_));
  NOR2_X1    g06039(.A1(new_n403_), .A2(new_n5993_), .ZN(new_n6316_));
  OAI21_X1   g06040(.A1(new_n6314_), .A2(new_n6315_), .B(new_n6316_), .ZN(new_n6317_));
  NAND2_X1   g06041(.A1(new_n6317_), .A2(\a[41] ), .ZN(new_n6318_));
  NOR2_X1    g06042(.A1(new_n6315_), .A2(new_n6314_), .ZN(new_n6319_));
  NOR3_X1    g06043(.A1(new_n6319_), .A2(new_n403_), .A3(new_n5993_), .ZN(new_n6320_));
  NAND2_X1   g06044(.A1(new_n6320_), .A2(new_n5681_), .ZN(new_n6321_));
  XNOR2_X1   g06045(.A1(\a[41] ), .A2(\a[42] ), .ZN(new_n6322_));
  NOR2_X1    g06046(.A1(new_n6322_), .A2(new_n258_), .ZN(new_n6323_));
  INV_X1     g06047(.I(new_n6323_), .ZN(new_n6324_));
  AOI21_X1   g06048(.A1(new_n6318_), .A2(new_n6321_), .B(new_n6324_), .ZN(new_n6325_));
  NAND2_X1   g06049(.A1(new_n6325_), .A2(new_n6003_), .ZN(new_n6326_));
  NOR2_X1    g06050(.A1(new_n6320_), .A2(new_n5681_), .ZN(new_n6327_));
  NOR2_X1    g06051(.A1(new_n6317_), .A2(\a[41] ), .ZN(new_n6328_));
  OAI21_X1   g06052(.A1(new_n6328_), .A2(new_n6327_), .B(new_n6323_), .ZN(new_n6329_));
  NAND2_X1   g06053(.A1(new_n6329_), .A2(new_n6019_), .ZN(new_n6330_));
  AOI21_X1   g06054(.A1(new_n6330_), .A2(new_n6326_), .B(new_n6307_), .ZN(new_n6331_));
  NOR2_X1    g06055(.A1(new_n6329_), .A2(new_n6019_), .ZN(new_n6332_));
  NOR2_X1    g06056(.A1(new_n6325_), .A2(new_n6003_), .ZN(new_n6333_));
  NOR3_X1    g06057(.A1(new_n6332_), .A2(new_n6333_), .A3(new_n6011_), .ZN(new_n6334_));
  AOI22_X1   g06058(.A1(new_n4859_), .A2(\b[5] ), .B1(new_n4865_), .B2(\b[6] ), .ZN(new_n6335_));
  AOI21_X1   g06059(.A1(\b[4] ), .A2(new_n6005_), .B(new_n6335_), .ZN(new_n6336_));
  OAI21_X1   g06060(.A1(new_n6336_), .A2(\a[38] ), .B(new_n4859_), .ZN(new_n6337_));
  XOR2_X1    g06061(.A1(new_n556_), .A2(new_n6337_), .Z(new_n6338_));
  INV_X1     g06062(.I(new_n6338_), .ZN(new_n6339_));
  OAI21_X1   g06063(.A1(new_n6331_), .A2(new_n6334_), .B(new_n6339_), .ZN(new_n6340_));
  NOR2_X1    g06064(.A1(new_n6313_), .A2(new_n6340_), .ZN(new_n6341_));
  INV_X1     g06065(.I(new_n6340_), .ZN(new_n6342_));
  NOR3_X1    g06066(.A1(new_n6342_), .A2(new_n6311_), .A3(new_n6312_), .ZN(new_n6343_));
  OAI21_X1   g06067(.A1(new_n6341_), .A2(new_n6343_), .B(new_n6310_), .ZN(new_n6344_));
  OAI21_X1   g06068(.A1(new_n6312_), .A2(new_n6311_), .B(new_n6342_), .ZN(new_n6345_));
  NAND2_X1   g06069(.A1(new_n6313_), .A2(new_n6340_), .ZN(new_n6346_));
  NAND3_X1   g06070(.A1(new_n6346_), .A2(new_n6345_), .A3(new_n6309_), .ZN(new_n6347_));
  OAI22_X1   g06071(.A1(new_n4072_), .A2(new_n515_), .B1(new_n565_), .B2(new_n4067_), .ZN(new_n6348_));
  OAI21_X1   g06072(.A1(new_n472_), .A2(new_n4318_), .B(new_n6348_), .ZN(new_n6349_));
  AOI21_X1   g06073(.A1(new_n6349_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n6350_));
  XOR2_X1    g06074(.A1(new_n759_), .A2(new_n6350_), .Z(new_n6351_));
  AOI21_X1   g06075(.A1(new_n6344_), .A2(new_n6347_), .B(new_n6351_), .ZN(new_n6352_));
  NAND2_X1   g06076(.A1(new_n6304_), .A2(new_n6352_), .ZN(new_n6353_));
  AOI21_X1   g06077(.A1(new_n6047_), .A2(new_n6300_), .B(new_n5716_), .ZN(new_n6354_));
  NAND2_X1   g06078(.A1(new_n6303_), .A2(new_n5664_), .ZN(new_n6355_));
  NOR2_X1    g06079(.A1(new_n6354_), .A2(new_n6355_), .ZN(new_n6356_));
  INV_X1     g06080(.I(new_n6352_), .ZN(new_n6357_));
  NAND2_X1   g06081(.A1(new_n6356_), .A2(new_n6357_), .ZN(new_n6358_));
  AOI21_X1   g06082(.A1(new_n6353_), .A2(new_n6358_), .B(new_n6057_), .ZN(new_n6359_));
  NOR2_X1    g06083(.A1(new_n6356_), .A2(new_n6357_), .ZN(new_n6360_));
  NOR2_X1    g06084(.A1(new_n6304_), .A2(new_n6352_), .ZN(new_n6361_));
  NOR3_X1    g06085(.A1(new_n6361_), .A2(new_n6360_), .A3(new_n6046_), .ZN(new_n6362_));
  OAI22_X1   g06086(.A1(new_n706_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n780_), .ZN(new_n6363_));
  OAI21_X1   g06087(.A1(new_n656_), .A2(new_n3569_), .B(new_n6363_), .ZN(new_n6364_));
  AOI21_X1   g06088(.A1(new_n6364_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n6365_));
  XOR2_X1    g06089(.A1(new_n785_), .A2(new_n6365_), .Z(new_n6366_));
  INV_X1     g06090(.I(new_n6366_), .ZN(new_n6367_));
  OAI21_X1   g06091(.A1(new_n6359_), .A2(new_n6362_), .B(new_n6367_), .ZN(new_n6368_));
  AOI21_X1   g06092(.A1(new_n6297_), .A2(new_n6299_), .B(new_n6368_), .ZN(new_n6369_));
  AOI21_X1   g06093(.A1(new_n6286_), .A2(new_n5729_), .B(new_n5735_), .ZN(new_n6370_));
  OAI21_X1   g06094(.A1(new_n6286_), .A2(new_n5729_), .B(new_n5988_), .ZN(new_n6371_));
  OAI21_X1   g06095(.A1(new_n6361_), .A2(new_n6360_), .B(new_n6046_), .ZN(new_n6372_));
  NAND3_X1   g06096(.A1(new_n6353_), .A2(new_n6358_), .A3(new_n6057_), .ZN(new_n6373_));
  AOI21_X1   g06097(.A1(new_n6372_), .A2(new_n6373_), .B(new_n6366_), .ZN(new_n6374_));
  NOR3_X1    g06098(.A1(new_n6370_), .A2(new_n6371_), .A3(new_n6374_), .ZN(new_n6375_));
  OAI21_X1   g06099(.A1(new_n6369_), .A2(new_n6375_), .B(new_n6295_), .ZN(new_n6376_));
  OAI21_X1   g06100(.A1(new_n6370_), .A2(new_n6371_), .B(new_n6374_), .ZN(new_n6377_));
  NAND3_X1   g06101(.A1(new_n6297_), .A2(new_n6299_), .A3(new_n6368_), .ZN(new_n6378_));
  NAND3_X1   g06102(.A1(new_n6378_), .A2(new_n6377_), .A3(new_n6294_), .ZN(new_n6379_));
  OAI22_X1   g06103(.A1(new_n930_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1017_), .ZN(new_n6380_));
  OAI21_X1   g06104(.A1(new_n861_), .A2(new_n2884_), .B(new_n6380_), .ZN(new_n6381_));
  AOI21_X1   g06105(.A1(new_n6381_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n6382_));
  XOR2_X1    g06106(.A1(new_n1024_), .A2(new_n6382_), .Z(new_n6383_));
  AOI21_X1   g06107(.A1(new_n6376_), .A2(new_n6379_), .B(new_n6383_), .ZN(new_n6384_));
  NAND2_X1   g06108(.A1(new_n6384_), .A2(new_n6293_), .ZN(new_n6385_));
  INV_X1     g06109(.I(new_n5761_), .ZN(new_n6386_));
  AOI21_X1   g06110(.A1(new_n6093_), .A2(new_n5751_), .B(new_n6386_), .ZN(new_n6387_));
  INV_X1     g06111(.I(new_n6292_), .ZN(new_n6388_));
  NOR3_X1    g06112(.A1(new_n6387_), .A2(new_n6388_), .A3(new_n5651_), .ZN(new_n6389_));
  AOI21_X1   g06113(.A1(new_n6378_), .A2(new_n6377_), .B(new_n6294_), .ZN(new_n6390_));
  NOR3_X1    g06114(.A1(new_n6369_), .A2(new_n6375_), .A3(new_n6295_), .ZN(new_n6391_));
  INV_X1     g06115(.I(new_n6383_), .ZN(new_n6392_));
  OAI21_X1   g06116(.A1(new_n6390_), .A2(new_n6391_), .B(new_n6392_), .ZN(new_n6393_));
  NAND2_X1   g06117(.A1(new_n6393_), .A2(new_n6389_), .ZN(new_n6394_));
  AOI21_X1   g06118(.A1(new_n6394_), .A2(new_n6385_), .B(new_n6289_), .ZN(new_n6395_));
  INV_X1     g06119(.I(new_n6289_), .ZN(new_n6396_));
  NOR2_X1    g06120(.A1(new_n6393_), .A2(new_n6389_), .ZN(new_n6397_));
  NOR2_X1    g06121(.A1(new_n6384_), .A2(new_n6293_), .ZN(new_n6398_));
  NOR3_X1    g06122(.A1(new_n6397_), .A2(new_n6398_), .A3(new_n6396_), .ZN(new_n6399_));
  OAI22_X1   g06123(.A1(new_n2171_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n2166_), .ZN(new_n6400_));
  OAI21_X1   g06124(.A1(new_n1109_), .A2(new_n2322_), .B(new_n6400_), .ZN(new_n6401_));
  AOI21_X1   g06125(.A1(new_n6401_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n6402_));
  XOR2_X1    g06126(.A1(new_n1299_), .A2(new_n6402_), .Z(new_n6403_));
  INV_X1     g06127(.I(new_n6403_), .ZN(new_n6404_));
  OAI21_X1   g06128(.A1(new_n6395_), .A2(new_n6399_), .B(new_n6404_), .ZN(new_n6405_));
  NOR2_X1    g06129(.A1(new_n6285_), .A2(new_n6405_), .ZN(new_n6406_));
  AOI21_X1   g06130(.A1(new_n6114_), .A2(new_n6115_), .B(new_n5795_), .ZN(new_n6407_));
  OAI21_X1   g06131(.A1(new_n6407_), .A2(new_n5782_), .B(new_n5796_), .ZN(new_n6408_));
  OAI21_X1   g06132(.A1(new_n6397_), .A2(new_n6398_), .B(new_n6396_), .ZN(new_n6409_));
  NAND3_X1   g06133(.A1(new_n6394_), .A2(new_n6385_), .A3(new_n6289_), .ZN(new_n6410_));
  AOI21_X1   g06134(.A1(new_n6409_), .A2(new_n6410_), .B(new_n6403_), .ZN(new_n6411_));
  NOR2_X1    g06135(.A1(new_n6408_), .A2(new_n6411_), .ZN(new_n6412_));
  OAI21_X1   g06136(.A1(new_n6406_), .A2(new_n6412_), .B(new_n6283_), .ZN(new_n6413_));
  AOI21_X1   g06137(.A1(new_n6096_), .A2(new_n6102_), .B(new_n6110_), .ZN(new_n6414_));
  NAND2_X1   g06138(.A1(new_n6408_), .A2(new_n6411_), .ZN(new_n6415_));
  NAND2_X1   g06139(.A1(new_n6285_), .A2(new_n6405_), .ZN(new_n6416_));
  NAND3_X1   g06140(.A1(new_n6416_), .A2(new_n6415_), .A3(new_n6414_), .ZN(new_n6417_));
  NAND2_X1   g06141(.A1(new_n6413_), .A2(new_n6417_), .ZN(new_n6418_));
  OAI22_X1   g06142(.A1(new_n1712_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n1707_), .ZN(new_n6419_));
  OAI21_X1   g06143(.A1(new_n1518_), .A2(new_n1850_), .B(new_n6419_), .ZN(new_n6420_));
  AOI21_X1   g06144(.A1(new_n6420_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n6421_));
  XNOR2_X1   g06145(.A1(new_n1638_), .A2(new_n6421_), .ZN(new_n6422_));
  INV_X1     g06146(.I(new_n6422_), .ZN(new_n6423_));
  NAND2_X1   g06147(.A1(new_n6418_), .A2(new_n6423_), .ZN(new_n6424_));
  NOR2_X1    g06148(.A1(new_n6424_), .A2(new_n6282_), .ZN(new_n6425_));
  AOI21_X1   g06149(.A1(new_n6132_), .A2(new_n6131_), .B(new_n6130_), .ZN(new_n6426_));
  OAI21_X1   g06150(.A1(new_n6426_), .A2(new_n5818_), .B(new_n5646_), .ZN(new_n6427_));
  AOI21_X1   g06151(.A1(new_n6418_), .A2(new_n6423_), .B(new_n6427_), .ZN(new_n6428_));
  OAI21_X1   g06152(.A1(new_n6428_), .A2(new_n6425_), .B(new_n6132_), .ZN(new_n6429_));
  NAND3_X1   g06153(.A1(new_n6427_), .A2(new_n6418_), .A3(new_n6423_), .ZN(new_n6430_));
  NAND2_X1   g06154(.A1(new_n6424_), .A2(new_n6282_), .ZN(new_n6431_));
  NAND3_X1   g06155(.A1(new_n6431_), .A2(new_n6430_), .A3(new_n6126_), .ZN(new_n6432_));
  OAI22_X1   g06156(.A1(new_n1347_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n1344_), .ZN(new_n6433_));
  OAI21_X1   g06157(.A1(new_n1803_), .A2(new_n1457_), .B(new_n6433_), .ZN(new_n6434_));
  AOI21_X1   g06158(.A1(new_n6434_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n6435_));
  XOR2_X1    g06159(.A1(new_n2106_), .A2(new_n6435_), .Z(new_n6436_));
  AOI21_X1   g06160(.A1(new_n6429_), .A2(new_n6432_), .B(new_n6436_), .ZN(new_n6437_));
  NAND2_X1   g06161(.A1(new_n6437_), .A2(new_n6280_), .ZN(new_n6438_));
  AOI21_X1   g06162(.A1(new_n6277_), .A2(new_n6276_), .B(new_n5979_), .ZN(new_n6439_));
  NOR3_X1    g06163(.A1(new_n6134_), .A2(new_n6128_), .A3(new_n5980_), .ZN(new_n6440_));
  OAI21_X1   g06164(.A1(new_n6439_), .A2(new_n6440_), .B(new_n6145_), .ZN(new_n6441_));
  AOI21_X1   g06165(.A1(new_n6441_), .A2(new_n5973_), .B(new_n5834_), .ZN(new_n6442_));
  AOI21_X1   g06166(.A1(new_n6431_), .A2(new_n6430_), .B(new_n6126_), .ZN(new_n6443_));
  NOR3_X1    g06167(.A1(new_n6428_), .A2(new_n6425_), .A3(new_n6132_), .ZN(new_n6444_));
  INV_X1     g06168(.I(new_n6436_), .ZN(new_n6445_));
  OAI21_X1   g06169(.A1(new_n6444_), .A2(new_n6443_), .B(new_n6445_), .ZN(new_n6446_));
  NAND2_X1   g06170(.A1(new_n6442_), .A2(new_n6446_), .ZN(new_n6447_));
  AOI21_X1   g06171(.A1(new_n6447_), .A2(new_n6438_), .B(new_n6274_), .ZN(new_n6448_));
  INV_X1     g06172(.I(new_n6274_), .ZN(new_n6449_));
  NOR2_X1    g06173(.A1(new_n6442_), .A2(new_n6446_), .ZN(new_n6450_));
  NOR2_X1    g06174(.A1(new_n6437_), .A2(new_n6280_), .ZN(new_n6451_));
  NOR3_X1    g06175(.A1(new_n6450_), .A2(new_n6451_), .A3(new_n6449_), .ZN(new_n6452_));
  NOR2_X1    g06176(.A1(new_n6448_), .A2(new_n6452_), .ZN(new_n6453_));
  OAI22_X1   g06177(.A1(new_n1055_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n1061_), .ZN(new_n6454_));
  OAI21_X1   g06178(.A1(new_n2281_), .A2(new_n1332_), .B(new_n6454_), .ZN(new_n6455_));
  AOI21_X1   g06179(.A1(new_n6455_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n6456_));
  XNOR2_X1   g06180(.A1(new_n2647_), .A2(new_n6456_), .ZN(new_n6457_));
  NOR2_X1    g06181(.A1(new_n6453_), .A2(new_n6457_), .ZN(new_n6458_));
  NAND2_X1   g06182(.A1(new_n6273_), .A2(new_n6458_), .ZN(new_n6459_));
  OAI21_X1   g06183(.A1(new_n6157_), .A2(new_n6154_), .B(new_n5975_), .ZN(new_n6460_));
  AOI21_X1   g06184(.A1(new_n6460_), .A2(new_n5839_), .B(new_n5850_), .ZN(new_n6461_));
  OAI21_X1   g06185(.A1(new_n6450_), .A2(new_n6451_), .B(new_n6449_), .ZN(new_n6462_));
  NAND3_X1   g06186(.A1(new_n6447_), .A2(new_n6438_), .A3(new_n6274_), .ZN(new_n6463_));
  NAND2_X1   g06187(.A1(new_n6462_), .A2(new_n6463_), .ZN(new_n6464_));
  INV_X1     g06188(.I(new_n6457_), .ZN(new_n6465_));
  NAND2_X1   g06189(.A1(new_n6464_), .A2(new_n6465_), .ZN(new_n6466_));
  NAND2_X1   g06190(.A1(new_n6461_), .A2(new_n6466_), .ZN(new_n6467_));
  AOI21_X1   g06191(.A1(new_n6467_), .A2(new_n6459_), .B(new_n6271_), .ZN(new_n6468_));
  AOI21_X1   g06192(.A1(new_n6269_), .A2(new_n6268_), .B(new_n5980_), .ZN(new_n6469_));
  NOR3_X1    g06193(.A1(new_n6264_), .A2(new_n6266_), .A3(new_n5979_), .ZN(new_n6470_));
  OAI21_X1   g06194(.A1(new_n6469_), .A2(new_n6470_), .B(new_n6147_), .ZN(new_n6471_));
  NOR2_X1    g06195(.A1(new_n6461_), .A2(new_n6466_), .ZN(new_n6472_));
  NOR2_X1    g06196(.A1(new_n6273_), .A2(new_n6458_), .ZN(new_n6473_));
  NOR3_X1    g06197(.A1(new_n6472_), .A2(new_n6473_), .A3(new_n6471_), .ZN(new_n6474_));
  OAI22_X1   g06198(.A1(new_n970_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n820_), .ZN(new_n6475_));
  OAI21_X1   g06199(.A1(new_n2842_), .A2(new_n894_), .B(new_n6475_), .ZN(new_n6476_));
  AOI21_X1   g06200(.A1(new_n6476_), .A2(new_n827_), .B(new_n970_), .ZN(new_n6477_));
  XNOR2_X1   g06201(.A1(new_n3264_), .A2(new_n6477_), .ZN(new_n6478_));
  INV_X1     g06202(.I(new_n6478_), .ZN(new_n6479_));
  OAI21_X1   g06203(.A1(new_n6468_), .A2(new_n6474_), .B(new_n6479_), .ZN(new_n6480_));
  OR2_X2     g06204(.A1(new_n6262_), .A2(new_n6480_), .Z(new_n6481_));
  NAND2_X1   g06205(.A1(new_n6262_), .A2(new_n6480_), .ZN(new_n6482_));
  AOI21_X1   g06206(.A1(new_n6481_), .A2(new_n6482_), .B(new_n6260_), .ZN(new_n6483_));
  INV_X1     g06207(.I(new_n6260_), .ZN(new_n6484_));
  NOR2_X1    g06208(.A1(new_n6262_), .A2(new_n6480_), .ZN(new_n6485_));
  INV_X1     g06209(.I(new_n6482_), .ZN(new_n6486_));
  NOR3_X1    g06210(.A1(new_n6486_), .A2(new_n6484_), .A3(new_n6485_), .ZN(new_n6487_));
  OAI22_X1   g06211(.A1(new_n607_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n610_), .ZN(new_n6488_));
  OAI21_X1   g06212(.A1(new_n3709_), .A2(new_n684_), .B(new_n6488_), .ZN(new_n6489_));
  AOI21_X1   g06213(.A1(new_n6489_), .A2(new_n612_), .B(new_n607_), .ZN(new_n6490_));
  XNOR2_X1   g06214(.A1(new_n3993_), .A2(new_n6490_), .ZN(new_n6491_));
  INV_X1     g06215(.I(new_n6491_), .ZN(new_n6492_));
  OAI21_X1   g06216(.A1(new_n6487_), .A2(new_n6483_), .B(new_n6492_), .ZN(new_n6493_));
  NOR2_X1    g06217(.A1(new_n6259_), .A2(new_n6493_), .ZN(new_n6494_));
  NOR2_X1    g06218(.A1(new_n5576_), .A2(new_n5624_), .ZN(new_n6495_));
  OAI22_X1   g06219(.A1(new_n6495_), .A2(new_n5621_), .B1(new_n5872_), .B2(new_n6195_), .ZN(new_n6496_));
  OAI21_X1   g06220(.A1(new_n6486_), .A2(new_n6485_), .B(new_n6484_), .ZN(new_n6497_));
  NAND3_X1   g06221(.A1(new_n6481_), .A2(new_n6260_), .A3(new_n6482_), .ZN(new_n6498_));
  AOI21_X1   g06222(.A1(new_n6497_), .A2(new_n6498_), .B(new_n6491_), .ZN(new_n6499_));
  NOR3_X1    g06223(.A1(new_n6496_), .A2(new_n6499_), .A3(new_n6257_), .ZN(new_n6500_));
  OAI21_X1   g06224(.A1(new_n6494_), .A2(new_n6500_), .B(new_n6256_), .ZN(new_n6501_));
  OAI21_X1   g06225(.A1(new_n6496_), .A2(new_n6257_), .B(new_n6499_), .ZN(new_n6502_));
  NAND2_X1   g06226(.A1(new_n6259_), .A2(new_n6493_), .ZN(new_n6503_));
  NAND3_X1   g06227(.A1(new_n6502_), .A2(new_n6503_), .A3(new_n6255_), .ZN(new_n6504_));
  NAND2_X1   g06228(.A1(new_n6504_), .A2(new_n6501_), .ZN(new_n6505_));
  OAI22_X1   g06229(.A1(new_n448_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n450_), .ZN(new_n6506_));
  OAI21_X1   g06230(.A1(new_n4253_), .A2(new_n496_), .B(new_n6506_), .ZN(new_n6507_));
  AOI21_X1   g06231(.A1(new_n6507_), .A2(new_n452_), .B(new_n448_), .ZN(new_n6508_));
  XNOR2_X1   g06232(.A1(new_n4778_), .A2(new_n6508_), .ZN(new_n6509_));
  INV_X1     g06233(.I(new_n6509_), .ZN(new_n6510_));
  NAND3_X1   g06234(.A1(new_n6254_), .A2(new_n6505_), .A3(new_n6510_), .ZN(new_n6511_));
  AOI21_X1   g06235(.A1(new_n6212_), .A2(new_n5884_), .B(new_n5889_), .ZN(new_n6512_));
  NOR2_X1    g06236(.A1(new_n6212_), .A2(new_n5884_), .ZN(new_n6513_));
  NOR3_X1    g06237(.A1(new_n6512_), .A2(new_n5620_), .A3(new_n6513_), .ZN(new_n6514_));
  AOI21_X1   g06238(.A1(new_n6502_), .A2(new_n6503_), .B(new_n6255_), .ZN(new_n6515_));
  NOR3_X1    g06239(.A1(new_n6494_), .A2(new_n6500_), .A3(new_n6256_), .ZN(new_n6516_));
  NOR2_X1    g06240(.A1(new_n6515_), .A2(new_n6516_), .ZN(new_n6517_));
  OAI21_X1   g06241(.A1(new_n6517_), .A2(new_n6509_), .B(new_n6514_), .ZN(new_n6518_));
  AOI21_X1   g06242(.A1(new_n6518_), .A2(new_n6511_), .B(new_n6249_), .ZN(new_n6519_));
  AND3_X2    g06243(.A1(new_n6518_), .A2(new_n6511_), .A3(new_n6249_), .Z(new_n6520_));
  NOR2_X1    g06244(.A1(new_n6520_), .A2(new_n6519_), .ZN(new_n6521_));
  INV_X1     g06245(.I(new_n6521_), .ZN(new_n6522_));
  INV_X1     g06246(.I(new_n6226_), .ZN(new_n6523_));
  NAND3_X1   g06247(.A1(new_n5952_), .A2(new_n5951_), .A3(new_n6212_), .ZN(new_n6524_));
  NAND3_X1   g06248(.A1(new_n5953_), .A2(new_n6208_), .A3(new_n6211_), .ZN(new_n6525_));
  AOI21_X1   g06249(.A1(new_n6525_), .A2(new_n6524_), .B(new_n6217_), .ZN(new_n6526_));
  AOI22_X1   g06250(.A1(new_n6221_), .A2(new_n6526_), .B1(new_n5894_), .B2(new_n6523_), .ZN(new_n6527_));
  NOR2_X1    g06251(.A1(new_n6225_), .A2(new_n6527_), .ZN(new_n6528_));
  NOR2_X1    g06252(.A1(\b[40] ), .A2(\b[41] ), .ZN(new_n6529_));
  AOI21_X1   g06253(.A1(new_n5917_), .A2(new_n6529_), .B(new_n5913_), .ZN(new_n6530_));
  NOR2_X1    g06254(.A1(new_n5921_), .A2(new_n6229_), .ZN(new_n6531_));
  INV_X1     g06255(.I(new_n6531_), .ZN(new_n6532_));
  NOR2_X1    g06256(.A1(new_n5917_), .A2(new_n6532_), .ZN(new_n6533_));
  NOR2_X1    g06257(.A1(new_n6530_), .A2(new_n6533_), .ZN(new_n6534_));
  INV_X1     g06258(.I(new_n6534_), .ZN(new_n6535_));
  XNOR2_X1   g06259(.A1(\b[41] ), .A2(\b[42] ), .ZN(new_n6536_));
  INV_X1     g06260(.I(new_n6536_), .ZN(new_n6537_));
  INV_X1     g06261(.I(\b[42] ), .ZN(new_n6538_));
  NOR2_X1    g06262(.A1(new_n6229_), .A2(new_n6538_), .ZN(new_n6539_));
  INV_X1     g06263(.I(new_n6539_), .ZN(new_n6540_));
  NAND2_X1   g06264(.A1(new_n6229_), .A2(new_n6538_), .ZN(new_n6541_));
  AOI21_X1   g06265(.A1(new_n6540_), .A2(new_n6541_), .B(new_n6535_), .ZN(new_n6542_));
  AOI21_X1   g06266(.A1(new_n6535_), .A2(new_n6537_), .B(new_n6542_), .ZN(new_n6543_));
  OAI22_X1   g06267(.A1(new_n330_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n263_), .ZN(new_n6544_));
  OAI21_X1   g06268(.A1(new_n5921_), .A2(new_n289_), .B(new_n6544_), .ZN(new_n6545_));
  AOI21_X1   g06269(.A1(new_n6545_), .A2(new_n260_), .B(new_n426_), .ZN(new_n6546_));
  XOR2_X1    g06270(.A1(new_n6543_), .A2(new_n6546_), .Z(new_n6547_));
  NOR2_X1    g06271(.A1(new_n6528_), .A2(new_n6547_), .ZN(new_n6548_));
  AND2_X2    g06272(.A1(new_n6528_), .A2(new_n6547_), .Z(new_n6549_));
  NOR2_X1    g06273(.A1(new_n6549_), .A2(new_n6548_), .ZN(new_n6550_));
  NOR2_X1    g06274(.A1(new_n6550_), .A2(new_n6522_), .ZN(new_n6551_));
  NOR3_X1    g06275(.A1(new_n6549_), .A2(new_n6521_), .A3(new_n6548_), .ZN(new_n6552_));
  NOR2_X1    g06276(.A1(new_n6551_), .A2(new_n6552_), .ZN(new_n6553_));
  NOR2_X1    g06277(.A1(new_n6553_), .A2(new_n6248_), .ZN(new_n6554_));
  NOR3_X1    g06278(.A1(new_n6551_), .A2(new_n6247_), .A3(new_n6552_), .ZN(new_n6555_));
  OAI21_X1   g06279(.A1(new_n6554_), .A2(new_n6555_), .B(new_n6240_), .ZN(new_n6556_));
  XNOR2_X1   g06280(.A1(new_n6556_), .A2(new_n6243_), .ZN(new_n6557_));
  XOR2_X1    g06281(.A1(new_n6557_), .A2(new_n5949_), .Z(\f[42] ));
  NOR2_X1    g06282(.A1(new_n6521_), .A2(new_n6247_), .ZN(new_n6559_));
  XOR2_X1    g06283(.A1(new_n6521_), .A2(new_n6248_), .Z(new_n6560_));
  OAI22_X1   g06284(.A1(new_n448_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n450_), .ZN(new_n6561_));
  OAI21_X1   g06285(.A1(new_n4500_), .A2(new_n496_), .B(new_n6561_), .ZN(new_n6562_));
  AOI21_X1   g06286(.A1(new_n6562_), .A2(new_n452_), .B(new_n448_), .ZN(new_n6563_));
  XOR2_X1    g06287(.A1(new_n5067_), .A2(new_n6563_), .Z(new_n6564_));
  NAND2_X1   g06288(.A1(new_n6497_), .A2(new_n6498_), .ZN(new_n6565_));
  NOR2_X1    g06289(.A1(new_n6487_), .A2(new_n6483_), .ZN(new_n6566_));
  AOI21_X1   g06290(.A1(new_n6566_), .A2(new_n6256_), .B(new_n6491_), .ZN(new_n6567_));
  AOI22_X1   g06291(.A1(new_n6567_), .A2(new_n6259_), .B1(new_n6565_), .B2(new_n6255_), .ZN(new_n6568_));
  OAI21_X1   g06292(.A1(new_n6472_), .A2(new_n6473_), .B(new_n6471_), .ZN(new_n6569_));
  NAND3_X1   g06293(.A1(new_n6467_), .A2(new_n6459_), .A3(new_n6271_), .ZN(new_n6570_));
  NAND2_X1   g06294(.A1(new_n6569_), .A2(new_n6570_), .ZN(new_n6571_));
  NAND2_X1   g06295(.A1(new_n6571_), .A2(new_n6260_), .ZN(new_n6572_));
  NAND3_X1   g06296(.A1(new_n6569_), .A2(new_n6570_), .A3(new_n6484_), .ZN(new_n6573_));
  NAND3_X1   g06297(.A1(new_n6262_), .A2(new_n6573_), .A3(new_n6479_), .ZN(new_n6574_));
  NAND2_X1   g06298(.A1(new_n6574_), .A2(new_n6572_), .ZN(new_n6575_));
  INV_X1     g06299(.I(new_n6575_), .ZN(new_n6576_));
  NAND2_X1   g06300(.A1(new_n6464_), .A2(new_n6271_), .ZN(new_n6577_));
  OAI21_X1   g06301(.A1(new_n6464_), .A2(new_n6271_), .B(new_n6465_), .ZN(new_n6578_));
  OAI21_X1   g06302(.A1(new_n6273_), .A2(new_n6578_), .B(new_n6577_), .ZN(new_n6579_));
  NAND2_X1   g06303(.A1(new_n6429_), .A2(new_n6432_), .ZN(new_n6580_));
  INV_X1     g06304(.I(new_n6580_), .ZN(new_n6581_));
  OAI21_X1   g06305(.A1(new_n6580_), .A2(new_n6274_), .B(new_n6445_), .ZN(new_n6582_));
  OAI22_X1   g06306(.A1(new_n6582_), .A2(new_n6280_), .B1(new_n6449_), .B2(new_n6581_), .ZN(new_n6583_));
  INV_X1     g06307(.I(new_n6583_), .ZN(new_n6584_));
  AOI21_X1   g06308(.A1(new_n6413_), .A2(new_n6417_), .B(new_n6132_), .ZN(new_n6585_));
  INV_X1     g06309(.I(new_n6585_), .ZN(new_n6586_));
  NAND3_X1   g06310(.A1(new_n6413_), .A2(new_n6417_), .A3(new_n6132_), .ZN(new_n6587_));
  NAND3_X1   g06311(.A1(new_n6282_), .A2(new_n6423_), .A3(new_n6587_), .ZN(new_n6588_));
  NAND2_X1   g06312(.A1(new_n6588_), .A2(new_n6586_), .ZN(new_n6589_));
  OAI21_X1   g06313(.A1(new_n6395_), .A2(new_n6399_), .B(new_n6414_), .ZN(new_n6590_));
  NAND3_X1   g06314(.A1(new_n6409_), .A2(new_n6410_), .A3(new_n6283_), .ZN(new_n6591_));
  NAND2_X1   g06315(.A1(new_n6591_), .A2(new_n6404_), .ZN(new_n6592_));
  OAI21_X1   g06316(.A1(new_n6592_), .A2(new_n6408_), .B(new_n6590_), .ZN(new_n6593_));
  AOI21_X1   g06317(.A1(new_n6376_), .A2(new_n6379_), .B(new_n6396_), .ZN(new_n6594_));
  INV_X1     g06318(.I(new_n6594_), .ZN(new_n6595_));
  NAND3_X1   g06319(.A1(new_n6376_), .A2(new_n6379_), .A3(new_n6396_), .ZN(new_n6596_));
  NOR4_X1    g06320(.A1(new_n6387_), .A2(new_n6388_), .A3(new_n5651_), .A4(new_n6383_), .ZN(new_n6597_));
  NAND2_X1   g06321(.A1(new_n6597_), .A2(new_n6596_), .ZN(new_n6598_));
  NAND2_X1   g06322(.A1(new_n6598_), .A2(new_n6595_), .ZN(new_n6599_));
  NOR2_X1    g06323(.A1(new_n6370_), .A2(new_n6371_), .ZN(new_n6600_));
  AOI21_X1   g06324(.A1(new_n6372_), .A2(new_n6373_), .B(new_n6295_), .ZN(new_n6601_));
  NOR3_X1    g06325(.A1(new_n6359_), .A2(new_n6362_), .A3(new_n6294_), .ZN(new_n6602_));
  NOR2_X1    g06326(.A1(new_n6602_), .A2(new_n6366_), .ZN(new_n6603_));
  AOI21_X1   g06327(.A1(new_n6600_), .A2(new_n6603_), .B(new_n6601_), .ZN(new_n6604_));
  AOI21_X1   g06328(.A1(new_n6344_), .A2(new_n6347_), .B(new_n6046_), .ZN(new_n6605_));
  AOI21_X1   g06329(.A1(new_n6346_), .A2(new_n6345_), .B(new_n6309_), .ZN(new_n6606_));
  NOR3_X1    g06330(.A1(new_n6341_), .A2(new_n6310_), .A3(new_n6343_), .ZN(new_n6607_));
  NOR3_X1    g06331(.A1(new_n6607_), .A2(new_n6606_), .A3(new_n6057_), .ZN(new_n6608_));
  NOR2_X1    g06332(.A1(new_n6608_), .A2(new_n6351_), .ZN(new_n6609_));
  AOI21_X1   g06333(.A1(new_n6356_), .A2(new_n6609_), .B(new_n6605_), .ZN(new_n6610_));
  OAI21_X1   g06334(.A1(new_n6331_), .A2(new_n6334_), .B(new_n6309_), .ZN(new_n6611_));
  OR3_X2     g06335(.A1(new_n6331_), .A2(new_n6334_), .A3(new_n6309_), .Z(new_n6612_));
  NAND3_X1   g06336(.A1(new_n6313_), .A2(new_n6339_), .A3(new_n6612_), .ZN(new_n6613_));
  NAND2_X1   g06337(.A1(new_n6318_), .A2(new_n6321_), .ZN(new_n6614_));
  NAND2_X1   g06338(.A1(new_n6614_), .A2(new_n6019_), .ZN(new_n6615_));
  NOR2_X1    g06339(.A1(new_n6614_), .A2(new_n6019_), .ZN(new_n6616_));
  NOR2_X1    g06340(.A1(new_n6011_), .A2(new_n6324_), .ZN(new_n6617_));
  INV_X1     g06341(.I(new_n6617_), .ZN(new_n6618_));
  OAI21_X1   g06342(.A1(new_n6616_), .A2(new_n6618_), .B(new_n6615_), .ZN(new_n6619_));
  AOI22_X1   g06343(.A1(new_n5680_), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n5686_), .ZN(new_n6620_));
  NOR2_X1    g06344(.A1(new_n5997_), .A2(new_n280_), .ZN(new_n6621_));
  OAI21_X1   g06345(.A1(new_n6620_), .A2(new_n6621_), .B(new_n5681_), .ZN(new_n6622_));
  NAND3_X1   g06346(.A1(new_n6622_), .A2(new_n807_), .A3(new_n5680_), .ZN(new_n6623_));
  OAI22_X1   g06347(.A1(new_n325_), .A2(new_n5991_), .B1(new_n5993_), .B2(new_n298_), .ZN(new_n6624_));
  INV_X1     g06348(.I(new_n6621_), .ZN(new_n6625_));
  AOI21_X1   g06349(.A1(new_n6625_), .A2(new_n6624_), .B(\a[41] ), .ZN(new_n6626_));
  OAI21_X1   g06350(.A1(new_n6626_), .A2(new_n5993_), .B(new_n329_), .ZN(new_n6627_));
  NAND2_X1   g06351(.A1(new_n6627_), .A2(new_n6623_), .ZN(new_n6628_));
  XNOR2_X1   g06352(.A1(\a[42] ), .A2(\a[44] ), .ZN(new_n6629_));
  XNOR2_X1   g06353(.A1(\a[41] ), .A2(\a[43] ), .ZN(new_n6630_));
  NOR2_X1    g06354(.A1(new_n6630_), .A2(new_n6629_), .ZN(new_n6631_));
  INV_X1     g06355(.I(\a[44] ), .ZN(new_n6632_));
  INV_X1     g06356(.I(\a[42] ), .ZN(new_n6633_));
  NAND3_X1   g06357(.A1(new_n5681_), .A2(new_n6633_), .A3(\a[43] ), .ZN(new_n6634_));
  INV_X1     g06358(.I(\a[43] ), .ZN(new_n6635_));
  NAND3_X1   g06359(.A1(new_n6635_), .A2(\a[41] ), .A3(\a[42] ), .ZN(new_n6636_));
  NAND2_X1   g06360(.A1(new_n6634_), .A2(new_n6636_), .ZN(new_n6637_));
  NAND2_X1   g06361(.A1(new_n6637_), .A2(\b[1] ), .ZN(new_n6638_));
  XOR2_X1    g06362(.A1(\a[42] ), .A2(\a[44] ), .Z(new_n6639_));
  XOR2_X1    g06363(.A1(\a[41] ), .A2(\a[43] ), .Z(new_n6640_));
  NAND3_X1   g06364(.A1(new_n6640_), .A2(new_n6639_), .A3(\b[0] ), .ZN(new_n6641_));
  NAND3_X1   g06365(.A1(new_n6638_), .A2(new_n6641_), .A3(new_n6632_), .ZN(new_n6642_));
  NAND3_X1   g06366(.A1(new_n6642_), .A2(new_n444_), .A3(new_n6631_), .ZN(new_n6643_));
  NAND2_X1   g06367(.A1(new_n6640_), .A2(new_n6639_), .ZN(new_n6644_));
  NOR3_X1    g06368(.A1(new_n6635_), .A2(\a[41] ), .A3(\a[42] ), .ZN(new_n6645_));
  NOR3_X1    g06369(.A1(new_n5681_), .A2(new_n6633_), .A3(\a[43] ), .ZN(new_n6646_));
  NOR2_X1    g06370(.A1(new_n6646_), .A2(new_n6645_), .ZN(new_n6647_));
  NOR2_X1    g06371(.A1(new_n6647_), .A2(new_n269_), .ZN(new_n6648_));
  NOR3_X1    g06372(.A1(new_n6630_), .A2(new_n6629_), .A3(new_n258_), .ZN(new_n6649_));
  NOR3_X1    g06373(.A1(new_n6648_), .A2(new_n6649_), .A3(\a[44] ), .ZN(new_n6650_));
  OAI21_X1   g06374(.A1(new_n6650_), .A2(new_n6644_), .B(new_n271_), .ZN(new_n6651_));
  NOR2_X1    g06375(.A1(new_n6323_), .A2(new_n6632_), .ZN(new_n6652_));
  INV_X1     g06376(.I(new_n6652_), .ZN(new_n6653_));
  NAND3_X1   g06377(.A1(new_n6651_), .A2(new_n6643_), .A3(new_n6653_), .ZN(new_n6654_));
  NOR3_X1    g06378(.A1(new_n6650_), .A2(new_n271_), .A3(new_n6644_), .ZN(new_n6655_));
  AOI21_X1   g06379(.A1(new_n6642_), .A2(new_n6631_), .B(new_n444_), .ZN(new_n6656_));
  OAI21_X1   g06380(.A1(new_n6655_), .A2(new_n6656_), .B(new_n6652_), .ZN(new_n6657_));
  NAND2_X1   g06381(.A1(new_n6657_), .A2(new_n6654_), .ZN(new_n6658_));
  NAND2_X1   g06382(.A1(new_n6628_), .A2(new_n6658_), .ZN(new_n6659_));
  NOR3_X1    g06383(.A1(new_n6626_), .A2(new_n329_), .A3(new_n5993_), .ZN(new_n6660_));
  AOI21_X1   g06384(.A1(new_n6622_), .A2(new_n5680_), .B(new_n807_), .ZN(new_n6661_));
  NOR2_X1    g06385(.A1(new_n6660_), .A2(new_n6661_), .ZN(new_n6662_));
  AND2_X2    g06386(.A1(new_n6657_), .A2(new_n6654_), .Z(new_n6663_));
  NAND2_X1   g06387(.A1(new_n6663_), .A2(new_n6662_), .ZN(new_n6664_));
  NAND2_X1   g06388(.A1(new_n6664_), .A2(new_n6659_), .ZN(new_n6665_));
  NAND2_X1   g06389(.A1(new_n6619_), .A2(new_n6665_), .ZN(new_n6666_));
  NOR2_X1    g06390(.A1(new_n6328_), .A2(new_n6327_), .ZN(new_n6667_));
  NOR2_X1    g06391(.A1(new_n6667_), .A2(new_n6003_), .ZN(new_n6668_));
  NAND2_X1   g06392(.A1(new_n6667_), .A2(new_n6003_), .ZN(new_n6669_));
  AOI21_X1   g06393(.A1(new_n6669_), .A2(new_n6617_), .B(new_n6668_), .ZN(new_n6670_));
  NAND2_X1   g06394(.A1(new_n6662_), .A2(new_n6658_), .ZN(new_n6671_));
  NAND2_X1   g06395(.A1(new_n6663_), .A2(new_n6628_), .ZN(new_n6672_));
  NAND2_X1   g06396(.A1(new_n6672_), .A2(new_n6671_), .ZN(new_n6673_));
  NAND2_X1   g06397(.A1(new_n6670_), .A2(new_n6673_), .ZN(new_n6674_));
  NAND2_X1   g06398(.A1(new_n6674_), .A2(new_n6666_), .ZN(new_n6675_));
  AOI22_X1   g06399(.A1(new_n4859_), .A2(\b[6] ), .B1(new_n4865_), .B2(\b[7] ), .ZN(new_n6676_));
  AOI21_X1   g06400(.A1(\b[5] ), .A2(new_n6005_), .B(new_n6676_), .ZN(new_n6677_));
  OAI21_X1   g06401(.A1(new_n6677_), .A2(\a[38] ), .B(new_n4859_), .ZN(new_n6678_));
  XNOR2_X1   g06402(.A1(new_n471_), .A2(new_n6678_), .ZN(new_n6679_));
  INV_X1     g06403(.I(new_n6679_), .ZN(new_n6680_));
  NAND2_X1   g06404(.A1(new_n6675_), .A2(new_n6680_), .ZN(new_n6681_));
  INV_X1     g06405(.I(new_n6675_), .ZN(new_n6682_));
  NAND2_X1   g06406(.A1(new_n6682_), .A2(new_n6679_), .ZN(new_n6683_));
  AOI22_X1   g06407(.A1(new_n6613_), .A2(new_n6611_), .B1(new_n6683_), .B2(new_n6681_), .ZN(new_n6684_));
  INV_X1     g06408(.I(new_n6684_), .ZN(new_n6685_));
  NAND3_X1   g06409(.A1(new_n6674_), .A2(new_n6666_), .A3(new_n6680_), .ZN(new_n6686_));
  NAND2_X1   g06410(.A1(new_n6675_), .A2(new_n6679_), .ZN(new_n6687_));
  NAND2_X1   g06411(.A1(new_n6687_), .A2(new_n6686_), .ZN(new_n6688_));
  NAND3_X1   g06412(.A1(new_n6613_), .A2(new_n6688_), .A3(new_n6611_), .ZN(new_n6689_));
  OAI22_X1   g06413(.A1(new_n4072_), .A2(new_n565_), .B1(new_n656_), .B2(new_n4067_), .ZN(new_n6690_));
  OAI21_X1   g06414(.A1(new_n515_), .A2(new_n4318_), .B(new_n6690_), .ZN(new_n6691_));
  AOI21_X1   g06415(.A1(new_n6691_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n6692_));
  XNOR2_X1   g06416(.A1(new_n660_), .A2(new_n6692_), .ZN(new_n6693_));
  INV_X1     g06417(.I(new_n6693_), .ZN(new_n6694_));
  NAND3_X1   g06418(.A1(new_n6685_), .A2(new_n6689_), .A3(new_n6694_), .ZN(new_n6695_));
  INV_X1     g06419(.I(new_n6689_), .ZN(new_n6696_));
  OAI21_X1   g06420(.A1(new_n6696_), .A2(new_n6684_), .B(new_n6693_), .ZN(new_n6697_));
  AOI21_X1   g06421(.A1(new_n6695_), .A2(new_n6697_), .B(new_n6610_), .ZN(new_n6698_));
  INV_X1     g06422(.I(new_n6605_), .ZN(new_n6699_));
  INV_X1     g06423(.I(new_n6351_), .ZN(new_n6700_));
  NAND3_X1   g06424(.A1(new_n6344_), .A2(new_n6347_), .A3(new_n6046_), .ZN(new_n6701_));
  NAND2_X1   g06425(.A1(new_n6701_), .A2(new_n6700_), .ZN(new_n6702_));
  OAI21_X1   g06426(.A1(new_n6304_), .A2(new_n6702_), .B(new_n6699_), .ZN(new_n6703_));
  AOI21_X1   g06427(.A1(new_n6685_), .A2(new_n6689_), .B(new_n6693_), .ZN(new_n6704_));
  NAND3_X1   g06428(.A1(new_n6685_), .A2(new_n6689_), .A3(new_n6693_), .ZN(new_n6705_));
  INV_X1     g06429(.I(new_n6705_), .ZN(new_n6706_));
  NOR2_X1    g06430(.A1(new_n6706_), .A2(new_n6704_), .ZN(new_n6707_));
  NOR2_X1    g06431(.A1(new_n6707_), .A2(new_n6703_), .ZN(new_n6708_));
  OAI22_X1   g06432(.A1(new_n780_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n861_), .ZN(new_n6709_));
  OAI21_X1   g06433(.A1(new_n706_), .A2(new_n3569_), .B(new_n6709_), .ZN(new_n6710_));
  AOI21_X1   g06434(.A1(new_n6710_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n6711_));
  XNOR2_X1   g06435(.A1(new_n860_), .A2(new_n6711_), .ZN(new_n6712_));
  NOR3_X1    g06436(.A1(new_n6698_), .A2(new_n6708_), .A3(new_n6712_), .ZN(new_n6713_));
  NAND2_X1   g06437(.A1(new_n6695_), .A2(new_n6697_), .ZN(new_n6714_));
  NAND2_X1   g06438(.A1(new_n6703_), .A2(new_n6714_), .ZN(new_n6715_));
  OAI21_X1   g06439(.A1(new_n6704_), .A2(new_n6706_), .B(new_n6610_), .ZN(new_n6716_));
  INV_X1     g06440(.I(new_n6712_), .ZN(new_n6717_));
  AOI21_X1   g06441(.A1(new_n6716_), .A2(new_n6715_), .B(new_n6717_), .ZN(new_n6718_));
  NOR2_X1    g06442(.A1(new_n6713_), .A2(new_n6718_), .ZN(new_n6719_));
  OAI22_X1   g06443(.A1(new_n1017_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1109_), .ZN(new_n6720_));
  OAI21_X1   g06444(.A1(new_n930_), .A2(new_n2884_), .B(new_n6720_), .ZN(new_n6721_));
  AOI21_X1   g06445(.A1(new_n6721_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n6722_));
  XOR2_X1    g06446(.A1(new_n1114_), .A2(new_n6722_), .Z(new_n6723_));
  INV_X1     g06447(.I(new_n6723_), .ZN(new_n6724_));
  NAND2_X1   g06448(.A1(new_n6719_), .A2(new_n6724_), .ZN(new_n6725_));
  NAND3_X1   g06449(.A1(new_n6716_), .A2(new_n6715_), .A3(new_n6717_), .ZN(new_n6726_));
  OAI21_X1   g06450(.A1(new_n6698_), .A2(new_n6708_), .B(new_n6712_), .ZN(new_n6727_));
  NAND2_X1   g06451(.A1(new_n6727_), .A2(new_n6726_), .ZN(new_n6728_));
  NAND2_X1   g06452(.A1(new_n6728_), .A2(new_n6723_), .ZN(new_n6729_));
  AOI21_X1   g06453(.A1(new_n6725_), .A2(new_n6729_), .B(new_n6604_), .ZN(new_n6730_));
  NAND2_X1   g06454(.A1(new_n6299_), .A2(new_n6297_), .ZN(new_n6731_));
  INV_X1     g06455(.I(new_n6601_), .ZN(new_n6732_));
  NAND3_X1   g06456(.A1(new_n6372_), .A2(new_n6373_), .A3(new_n6295_), .ZN(new_n6733_));
  NAND2_X1   g06457(.A1(new_n6733_), .A2(new_n6367_), .ZN(new_n6734_));
  OAI21_X1   g06458(.A1(new_n6731_), .A2(new_n6734_), .B(new_n6732_), .ZN(new_n6735_));
  NAND2_X1   g06459(.A1(new_n6728_), .A2(new_n6724_), .ZN(new_n6736_));
  NAND2_X1   g06460(.A1(new_n6719_), .A2(new_n6723_), .ZN(new_n6737_));
  AOI21_X1   g06461(.A1(new_n6736_), .A2(new_n6737_), .B(new_n6735_), .ZN(new_n6738_));
  NOR2_X1    g06462(.A1(new_n6738_), .A2(new_n6730_), .ZN(new_n6739_));
  OAI22_X1   g06463(.A1(new_n2171_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n2166_), .ZN(new_n6740_));
  OAI21_X1   g06464(.A1(new_n1189_), .A2(new_n2322_), .B(new_n6740_), .ZN(new_n6741_));
  AOI21_X1   g06465(.A1(new_n6741_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n6742_));
  XNOR2_X1   g06466(.A1(new_n1421_), .A2(new_n6742_), .ZN(new_n6743_));
  NOR2_X1    g06467(.A1(new_n6739_), .A2(new_n6743_), .ZN(new_n6744_));
  OR2_X2     g06468(.A1(new_n6738_), .A2(new_n6730_), .Z(new_n6745_));
  INV_X1     g06469(.I(new_n6743_), .ZN(new_n6746_));
  NOR2_X1    g06470(.A1(new_n6745_), .A2(new_n6746_), .ZN(new_n6747_));
  OAI21_X1   g06471(.A1(new_n6747_), .A2(new_n6744_), .B(new_n6599_), .ZN(new_n6748_));
  AOI21_X1   g06472(.A1(new_n6597_), .A2(new_n6596_), .B(new_n6594_), .ZN(new_n6749_));
  NOR2_X1    g06473(.A1(new_n6745_), .A2(new_n6743_), .ZN(new_n6750_));
  NOR2_X1    g06474(.A1(new_n6739_), .A2(new_n6746_), .ZN(new_n6751_));
  OAI21_X1   g06475(.A1(new_n6750_), .A2(new_n6751_), .B(new_n6749_), .ZN(new_n6752_));
  NAND2_X1   g06476(.A1(new_n6748_), .A2(new_n6752_), .ZN(new_n6753_));
  OAI22_X1   g06477(.A1(new_n1712_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n1707_), .ZN(new_n6754_));
  OAI21_X1   g06478(.A1(new_n1525_), .A2(new_n1850_), .B(new_n6754_), .ZN(new_n6755_));
  AOI21_X1   g06479(.A1(new_n6755_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n6756_));
  XOR2_X1    g06480(.A1(new_n1808_), .A2(new_n6756_), .Z(new_n6757_));
  INV_X1     g06481(.I(new_n6757_), .ZN(new_n6758_));
  NAND2_X1   g06482(.A1(new_n6753_), .A2(new_n6758_), .ZN(new_n6759_));
  NAND3_X1   g06483(.A1(new_n6748_), .A2(new_n6752_), .A3(new_n6757_), .ZN(new_n6760_));
  NAND2_X1   g06484(.A1(new_n6759_), .A2(new_n6760_), .ZN(new_n6761_));
  NAND3_X1   g06485(.A1(new_n6748_), .A2(new_n6752_), .A3(new_n6758_), .ZN(new_n6762_));
  NAND2_X1   g06486(.A1(new_n6753_), .A2(new_n6757_), .ZN(new_n6763_));
  AOI21_X1   g06487(.A1(new_n6762_), .A2(new_n6763_), .B(new_n6593_), .ZN(new_n6764_));
  AOI21_X1   g06488(.A1(new_n6593_), .A2(new_n6761_), .B(new_n6764_), .ZN(new_n6765_));
  OAI22_X1   g06489(.A1(new_n1347_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n1344_), .ZN(new_n6766_));
  OAI21_X1   g06490(.A1(new_n1936_), .A2(new_n1457_), .B(new_n6766_), .ZN(new_n6767_));
  AOI21_X1   g06491(.A1(new_n6767_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n6768_));
  XNOR2_X1   g06492(.A1(new_n2280_), .A2(new_n6768_), .ZN(new_n6769_));
  INV_X1     g06493(.I(new_n6769_), .ZN(new_n6770_));
  XOR2_X1    g06494(.A1(new_n6765_), .A2(new_n6770_), .Z(new_n6771_));
  NAND2_X1   g06495(.A1(new_n6771_), .A2(new_n6589_), .ZN(new_n6772_));
  XOR2_X1    g06496(.A1(new_n6765_), .A2(new_n6770_), .Z(new_n6773_));
  OAI21_X1   g06497(.A1(new_n6589_), .A2(new_n6773_), .B(new_n6772_), .ZN(new_n6774_));
  OAI22_X1   g06498(.A1(new_n1055_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n1061_), .ZN(new_n6775_));
  OAI21_X1   g06499(.A1(new_n2439_), .A2(new_n1332_), .B(new_n6775_), .ZN(new_n6776_));
  AOI21_X1   g06500(.A1(new_n6776_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n6777_));
  XNOR2_X1   g06501(.A1(new_n2846_), .A2(new_n6777_), .ZN(new_n6778_));
  INV_X1     g06502(.I(new_n6778_), .ZN(new_n6779_));
  NAND2_X1   g06503(.A1(new_n6774_), .A2(new_n6779_), .ZN(new_n6780_));
  NOR2_X1    g06504(.A1(new_n6773_), .A2(new_n6589_), .ZN(new_n6781_));
  AOI21_X1   g06505(.A1(new_n6589_), .A2(new_n6771_), .B(new_n6781_), .ZN(new_n6782_));
  NAND2_X1   g06506(.A1(new_n6782_), .A2(new_n6778_), .ZN(new_n6783_));
  AND2_X2    g06507(.A1(new_n6783_), .A2(new_n6780_), .Z(new_n6784_));
  NOR2_X1    g06508(.A1(new_n6774_), .A2(new_n6778_), .ZN(new_n6785_));
  NOR2_X1    g06509(.A1(new_n6782_), .A2(new_n6779_), .ZN(new_n6786_));
  OAI21_X1   g06510(.A1(new_n6786_), .A2(new_n6785_), .B(new_n6584_), .ZN(new_n6787_));
  OAI21_X1   g06511(.A1(new_n6784_), .A2(new_n6584_), .B(new_n6787_), .ZN(new_n6788_));
  NAND2_X1   g06512(.A1(new_n6579_), .A2(new_n6788_), .ZN(new_n6789_));
  AOI21_X1   g06513(.A1(new_n6453_), .A2(new_n6471_), .B(new_n6457_), .ZN(new_n6790_));
  AOI22_X1   g06514(.A1(new_n6461_), .A2(new_n6790_), .B1(new_n6271_), .B2(new_n6464_), .ZN(new_n6791_));
  AOI21_X1   g06515(.A1(new_n6780_), .A2(new_n6783_), .B(new_n6584_), .ZN(new_n6792_));
  OR2_X2     g06516(.A1(new_n6786_), .A2(new_n6785_), .Z(new_n6793_));
  AOI21_X1   g06517(.A1(new_n6793_), .A2(new_n6584_), .B(new_n6792_), .ZN(new_n6794_));
  NAND2_X1   g06518(.A1(new_n6791_), .A2(new_n6794_), .ZN(new_n6795_));
  OAI22_X1   g06519(.A1(new_n970_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n820_), .ZN(new_n6796_));
  OAI21_X1   g06520(.A1(new_n3018_), .A2(new_n894_), .B(new_n6796_), .ZN(new_n6797_));
  AOI21_X1   g06521(.A1(new_n6797_), .A2(new_n827_), .B(new_n970_), .ZN(new_n6798_));
  XNOR2_X1   g06522(.A1(new_n3514_), .A2(new_n6798_), .ZN(new_n6799_));
  INV_X1     g06523(.I(new_n6799_), .ZN(new_n6800_));
  NAND3_X1   g06524(.A1(new_n6795_), .A2(new_n6789_), .A3(new_n6800_), .ZN(new_n6801_));
  NOR2_X1    g06525(.A1(new_n6791_), .A2(new_n6794_), .ZN(new_n6802_));
  NOR2_X1    g06526(.A1(new_n6579_), .A2(new_n6788_), .ZN(new_n6803_));
  OAI21_X1   g06527(.A1(new_n6802_), .A2(new_n6803_), .B(new_n6799_), .ZN(new_n6804_));
  NAND2_X1   g06528(.A1(new_n6804_), .A2(new_n6801_), .ZN(new_n6805_));
  OAI22_X1   g06529(.A1(new_n607_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n610_), .ZN(new_n6806_));
  OAI21_X1   g06530(.A1(new_n3717_), .A2(new_n684_), .B(new_n6806_), .ZN(new_n6807_));
  AOI21_X1   g06531(.A1(new_n6807_), .A2(new_n612_), .B(new_n607_), .ZN(new_n6808_));
  XNOR2_X1   g06532(.A1(new_n4257_), .A2(new_n6808_), .ZN(new_n6809_));
  XOR2_X1    g06533(.A1(new_n6805_), .A2(new_n6809_), .Z(new_n6810_));
  NOR2_X1    g06534(.A1(new_n6810_), .A2(new_n6576_), .ZN(new_n6811_));
  INV_X1     g06535(.I(new_n6809_), .ZN(new_n6812_));
  XOR2_X1    g06536(.A1(new_n6805_), .A2(new_n6812_), .Z(new_n6813_));
  NOR2_X1    g06537(.A1(new_n6813_), .A2(new_n6575_), .ZN(new_n6814_));
  NOR2_X1    g06538(.A1(new_n6811_), .A2(new_n6814_), .ZN(new_n6815_));
  XOR2_X1    g06539(.A1(new_n6568_), .A2(new_n6815_), .Z(new_n6816_));
  NOR2_X1    g06540(.A1(new_n6517_), .A2(new_n6211_), .ZN(new_n6817_));
  AOI21_X1   g06541(.A1(new_n6517_), .A2(new_n6211_), .B(new_n6509_), .ZN(new_n6818_));
  AOI21_X1   g06542(.A1(new_n6514_), .A2(new_n6818_), .B(new_n6817_), .ZN(new_n6819_));
  OAI22_X1   g06543(.A1(new_n5913_), .A2(new_n341_), .B1(new_n404_), .B2(new_n5921_), .ZN(new_n6820_));
  OAI21_X1   g06544(.A1(new_n5353_), .A2(new_n366_), .B(new_n6820_), .ZN(new_n6821_));
  AOI21_X1   g06545(.A1(new_n6821_), .A2(new_n334_), .B(new_n341_), .ZN(new_n6822_));
  XOR2_X1    g06546(.A1(new_n5926_), .A2(new_n6822_), .Z(new_n6823_));
  INV_X1     g06547(.I(new_n6823_), .ZN(new_n6824_));
  NAND2_X1   g06548(.A1(new_n6819_), .A2(new_n6824_), .ZN(new_n6825_));
  NAND2_X1   g06549(.A1(new_n6505_), .A2(new_n6249_), .ZN(new_n6826_));
  NAND3_X1   g06550(.A1(new_n6504_), .A2(new_n6501_), .A3(new_n6211_), .ZN(new_n6827_));
  NAND2_X1   g06551(.A1(new_n6827_), .A2(new_n6510_), .ZN(new_n6828_));
  OAI21_X1   g06552(.A1(new_n6254_), .A2(new_n6828_), .B(new_n6826_), .ZN(new_n6829_));
  NAND2_X1   g06553(.A1(new_n6829_), .A2(new_n6823_), .ZN(new_n6830_));
  AOI21_X1   g06554(.A1(new_n6825_), .A2(new_n6830_), .B(new_n6816_), .ZN(new_n6831_));
  INV_X1     g06555(.I(new_n6815_), .ZN(new_n6832_));
  XOR2_X1    g06556(.A1(new_n6568_), .A2(new_n6832_), .Z(new_n6833_));
  NOR2_X1    g06557(.A1(new_n6829_), .A2(new_n6823_), .ZN(new_n6834_));
  NOR2_X1    g06558(.A1(new_n6819_), .A2(new_n6824_), .ZN(new_n6835_));
  NOR3_X1    g06559(.A1(new_n6835_), .A2(new_n6834_), .A3(new_n6833_), .ZN(new_n6836_));
  OAI21_X1   g06560(.A1(new_n6831_), .A2(new_n6836_), .B(new_n6564_), .ZN(new_n6837_));
  INV_X1     g06561(.I(new_n6564_), .ZN(new_n6838_));
  OAI21_X1   g06562(.A1(new_n6835_), .A2(new_n6834_), .B(new_n6833_), .ZN(new_n6839_));
  NAND3_X1   g06563(.A1(new_n6825_), .A2(new_n6830_), .A3(new_n6816_), .ZN(new_n6840_));
  NAND3_X1   g06564(.A1(new_n6839_), .A2(new_n6840_), .A3(new_n6838_), .ZN(new_n6841_));
  NAND2_X1   g06565(.A1(new_n6837_), .A2(new_n6841_), .ZN(new_n6842_));
  INV_X1     g06566(.I(new_n6842_), .ZN(new_n6843_));
  NOR2_X1    g06567(.A1(new_n6560_), .A2(new_n6843_), .ZN(new_n6844_));
  XOR2_X1    g06568(.A1(new_n6844_), .A2(new_n6559_), .Z(new_n6845_));
  XOR2_X1    g06569(.A1(new_n6845_), .A2(new_n6528_), .Z(new_n6846_));
  INV_X1     g06570(.I(\b[43] ), .ZN(new_n6847_));
  NOR2_X1    g06571(.A1(new_n6847_), .A2(\b[41] ), .ZN(new_n6848_));
  NOR2_X1    g06572(.A1(new_n6229_), .A2(\b[43] ), .ZN(new_n6849_));
  OAI21_X1   g06573(.A1(new_n6848_), .A2(new_n6849_), .B(new_n6537_), .ZN(new_n6850_));
  XNOR2_X1   g06574(.A1(new_n6534_), .A2(new_n6850_), .ZN(new_n6851_));
  OAI22_X1   g06575(.A1(new_n330_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n263_), .ZN(new_n6852_));
  OAI21_X1   g06576(.A1(new_n6229_), .A2(new_n289_), .B(new_n6852_), .ZN(new_n6853_));
  AOI21_X1   g06577(.A1(new_n6853_), .A2(new_n260_), .B(new_n426_), .ZN(new_n6854_));
  XOR2_X1    g06578(.A1(new_n6851_), .A2(new_n6854_), .Z(new_n6855_));
  XOR2_X1    g06579(.A1(new_n6846_), .A2(new_n6855_), .Z(new_n6856_));
  INV_X1     g06580(.I(new_n6528_), .ZN(new_n6857_));
  NOR2_X1    g06581(.A1(new_n6522_), .A2(new_n6248_), .ZN(new_n6858_));
  OAI21_X1   g06582(.A1(new_n6559_), .A2(new_n6858_), .B(new_n6857_), .ZN(new_n6859_));
  INV_X1     g06583(.I(new_n6560_), .ZN(new_n6860_));
  NAND2_X1   g06584(.A1(new_n6860_), .A2(new_n6528_), .ZN(new_n6861_));
  NAND3_X1   g06585(.A1(new_n6861_), .A2(new_n6859_), .A3(new_n6547_), .ZN(new_n6862_));
  OAI21_X1   g06586(.A1(new_n6554_), .A2(new_n6555_), .B(new_n6228_), .ZN(new_n6863_));
  NAND2_X1   g06587(.A1(new_n6863_), .A2(new_n6237_), .ZN(new_n6864_));
  NOR3_X1    g06588(.A1(new_n6554_), .A2(new_n6228_), .A3(new_n6555_), .ZN(new_n6865_));
  NOR2_X1    g06589(.A1(new_n5949_), .A2(new_n6865_), .ZN(new_n6866_));
  NAND2_X1   g06590(.A1(new_n6866_), .A2(new_n6864_), .ZN(new_n6867_));
  NAND2_X1   g06591(.A1(new_n6867_), .A2(new_n6862_), .ZN(new_n6868_));
  XOR2_X1    g06592(.A1(new_n6868_), .A2(new_n6856_), .Z(\f[43] ));
  NAND3_X1   g06593(.A1(new_n6866_), .A2(new_n6864_), .A3(new_n6846_), .ZN(new_n6870_));
  AOI21_X1   g06594(.A1(new_n6866_), .A2(new_n6864_), .B(new_n6846_), .ZN(new_n6871_));
  NOR2_X1    g06595(.A1(new_n6862_), .A2(new_n6855_), .ZN(new_n6872_));
  INV_X1     g06596(.I(new_n6872_), .ZN(new_n6873_));
  OAI21_X1   g06597(.A1(new_n6871_), .A2(new_n6873_), .B(new_n6870_), .ZN(new_n6874_));
  INV_X1     g06598(.I(new_n6874_), .ZN(new_n6875_));
  NAND2_X1   g06599(.A1(new_n6833_), .A2(new_n6838_), .ZN(new_n6876_));
  OAI21_X1   g06600(.A1(new_n6838_), .A2(new_n6833_), .B(new_n6829_), .ZN(new_n6877_));
  NAND2_X1   g06601(.A1(new_n6877_), .A2(new_n6876_), .ZN(new_n6878_));
  NAND2_X1   g06602(.A1(new_n6575_), .A2(new_n6805_), .ZN(new_n6879_));
  INV_X1     g06603(.I(new_n6879_), .ZN(new_n6880_));
  NOR2_X1    g06604(.A1(new_n6575_), .A2(new_n6805_), .ZN(new_n6881_));
  OAI21_X1   g06605(.A1(new_n6880_), .A2(new_n6881_), .B(new_n6809_), .ZN(new_n6882_));
  NOR2_X1    g06606(.A1(new_n6802_), .A2(new_n6803_), .ZN(new_n6883_));
  NOR2_X1    g06607(.A1(new_n6883_), .A2(new_n6799_), .ZN(new_n6884_));
  NAND2_X1   g06608(.A1(new_n6584_), .A2(new_n6774_), .ZN(new_n6885_));
  NAND2_X1   g06609(.A1(new_n6583_), .A2(new_n6782_), .ZN(new_n6886_));
  AOI21_X1   g06610(.A1(new_n6885_), .A2(new_n6886_), .B(new_n6779_), .ZN(new_n6887_));
  INV_X1     g06611(.I(new_n6887_), .ZN(new_n6888_));
  XOR2_X1    g06612(.A1(new_n6589_), .A2(new_n6765_), .Z(new_n6889_));
  NOR2_X1    g06613(.A1(new_n6889_), .A2(new_n6770_), .ZN(new_n6890_));
  OAI22_X1   g06614(.A1(new_n1712_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n1707_), .ZN(new_n6891_));
  OAI21_X1   g06615(.A1(new_n1634_), .A2(new_n1850_), .B(new_n6891_), .ZN(new_n6892_));
  AOI21_X1   g06616(.A1(new_n6892_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n6893_));
  XNOR2_X1   g06617(.A1(new_n1940_), .A2(new_n6893_), .ZN(new_n6894_));
  INV_X1     g06618(.I(new_n6894_), .ZN(new_n6895_));
  INV_X1     g06619(.I(new_n6753_), .ZN(new_n6896_));
  NAND2_X1   g06620(.A1(new_n6745_), .A2(new_n6749_), .ZN(new_n6897_));
  NOR2_X1    g06621(.A1(new_n6745_), .A2(new_n6749_), .ZN(new_n6898_));
  INV_X1     g06622(.I(new_n6898_), .ZN(new_n6899_));
  AOI21_X1   g06623(.A1(new_n6899_), .A2(new_n6897_), .B(new_n6746_), .ZN(new_n6900_));
  NAND2_X1   g06624(.A1(new_n6735_), .A2(new_n6728_), .ZN(new_n6901_));
  NAND2_X1   g06625(.A1(new_n6604_), .A2(new_n6719_), .ZN(new_n6902_));
  AOI21_X1   g06626(.A1(new_n6901_), .A2(new_n6902_), .B(new_n6724_), .ZN(new_n6903_));
  NOR2_X1    g06627(.A1(new_n6698_), .A2(new_n6708_), .ZN(new_n6904_));
  NOR2_X1    g06628(.A1(new_n6904_), .A2(new_n6712_), .ZN(new_n6905_));
  INV_X1     g06629(.I(new_n6695_), .ZN(new_n6906_));
  AOI21_X1   g06630(.A1(new_n6703_), .A2(new_n6697_), .B(new_n6906_), .ZN(new_n6907_));
  NAND2_X1   g06631(.A1(new_n6613_), .A2(new_n6611_), .ZN(new_n6908_));
  INV_X1     g06632(.I(new_n6659_), .ZN(new_n6909_));
  NOR2_X1    g06633(.A1(new_n6647_), .A2(new_n280_), .ZN(new_n6910_));
  INV_X1     g06634(.I(new_n6910_), .ZN(new_n6911_));
  OAI21_X1   g06635(.A1(\b[1] ), .A2(new_n282_), .B(new_n6631_), .ZN(new_n6912_));
  XNOR2_X1   g06636(.A1(\a[41] ), .A2(\a[44] ), .ZN(new_n6913_));
  NOR3_X1    g06637(.A1(new_n6630_), .A2(new_n6322_), .A3(new_n6913_), .ZN(new_n6914_));
  NAND2_X1   g06638(.A1(new_n6914_), .A2(\b[0] ), .ZN(new_n6915_));
  AOI21_X1   g06639(.A1(new_n6912_), .A2(new_n6911_), .B(new_n6915_), .ZN(new_n6916_));
  NOR2_X1    g06640(.A1(new_n6916_), .A2(new_n6632_), .ZN(new_n6917_));
  AOI21_X1   g06641(.A1(new_n269_), .A2(new_n490_), .B(new_n6644_), .ZN(new_n6918_));
  NOR2_X1    g06642(.A1(new_n6918_), .A2(new_n6910_), .ZN(new_n6919_));
  NOR3_X1    g06643(.A1(new_n6919_), .A2(\a[44] ), .A3(new_n6915_), .ZN(new_n6920_));
  NOR2_X1    g06644(.A1(new_n6917_), .A2(new_n6920_), .ZN(new_n6921_));
  NOR3_X1    g06645(.A1(new_n6655_), .A2(new_n6656_), .A3(new_n6653_), .ZN(new_n6922_));
  INV_X1     g06646(.I(new_n5997_), .ZN(new_n6923_));
  NAND3_X1   g06647(.A1(new_n5689_), .A2(new_n5688_), .A3(\b[4] ), .ZN(new_n6924_));
  NAND2_X1   g06648(.A1(new_n5686_), .A2(\b[5] ), .ZN(new_n6925_));
  AOI22_X1   g06649(.A1(new_n6923_), .A2(\b[3] ), .B1(new_n6924_), .B2(new_n6925_), .ZN(new_n6926_));
  OAI21_X1   g06650(.A1(new_n2333_), .A2(new_n5993_), .B(new_n6926_), .ZN(new_n6927_));
  NOR2_X1    g06651(.A1(new_n6922_), .A2(new_n6927_), .ZN(new_n6928_));
  NAND3_X1   g06652(.A1(new_n6651_), .A2(new_n6643_), .A3(new_n6652_), .ZN(new_n6929_));
  INV_X1     g06653(.I(new_n6924_), .ZN(new_n6930_));
  INV_X1     g06654(.I(new_n6925_), .ZN(new_n6931_));
  OAI22_X1   g06655(.A1(new_n6931_), .A2(new_n6930_), .B1(new_n298_), .B2(new_n5997_), .ZN(new_n6932_));
  AOI21_X1   g06656(.A1(new_n378_), .A2(new_n5680_), .B(new_n6932_), .ZN(new_n6933_));
  NOR2_X1    g06657(.A1(new_n6929_), .A2(new_n6933_), .ZN(new_n6934_));
  OAI21_X1   g06658(.A1(new_n6934_), .A2(new_n6928_), .B(new_n6921_), .ZN(new_n6935_));
  OAI21_X1   g06659(.A1(new_n6919_), .A2(new_n6915_), .B(\a[44] ), .ZN(new_n6936_));
  NAND2_X1   g06660(.A1(new_n6916_), .A2(new_n6632_), .ZN(new_n6937_));
  NAND2_X1   g06661(.A1(new_n6937_), .A2(new_n6936_), .ZN(new_n6938_));
  NAND2_X1   g06662(.A1(new_n6929_), .A2(new_n6933_), .ZN(new_n6939_));
  NAND2_X1   g06663(.A1(new_n6922_), .A2(new_n6927_), .ZN(new_n6940_));
  NAND3_X1   g06664(.A1(new_n6939_), .A2(new_n6940_), .A3(new_n6938_), .ZN(new_n6941_));
  AOI21_X1   g06665(.A1(new_n6935_), .A2(new_n6941_), .B(\a[41] ), .ZN(new_n6942_));
  AOI21_X1   g06666(.A1(new_n6939_), .A2(new_n6940_), .B(new_n6938_), .ZN(new_n6943_));
  NOR3_X1    g06667(.A1(new_n6934_), .A2(new_n6928_), .A3(new_n6921_), .ZN(new_n6944_));
  NOR3_X1    g06668(.A1(new_n6943_), .A2(new_n6944_), .A3(new_n5681_), .ZN(new_n6945_));
  OAI21_X1   g06669(.A1(new_n6945_), .A2(new_n6942_), .B(new_n6673_), .ZN(new_n6946_));
  NOR2_X1    g06670(.A1(new_n6946_), .A2(new_n6909_), .ZN(new_n6947_));
  OAI21_X1   g06671(.A1(new_n6943_), .A2(new_n6944_), .B(new_n5681_), .ZN(new_n6948_));
  NAND3_X1   g06672(.A1(new_n6935_), .A2(new_n6941_), .A3(\a[41] ), .ZN(new_n6949_));
  NAND2_X1   g06673(.A1(new_n6948_), .A2(new_n6949_), .ZN(new_n6950_));
  NAND2_X1   g06674(.A1(new_n6628_), .A2(new_n6658_), .ZN(new_n6952_));
  INV_X1     g06675(.I(new_n6952_), .ZN(new_n6953_));
  OAI21_X1   g06676(.A1(new_n6947_), .A2(new_n6953_), .B(new_n6670_), .ZN(new_n6954_));
  NAND3_X1   g06677(.A1(new_n6950_), .A2(new_n6659_), .A3(new_n6673_), .ZN(new_n6955_));
  NAND3_X1   g06678(.A1(new_n6955_), .A2(new_n6619_), .A3(new_n6952_), .ZN(new_n6956_));
  OAI22_X1   g06679(.A1(new_n5420_), .A2(new_n472_), .B1(new_n515_), .B2(new_n5107_), .ZN(new_n6957_));
  OAI21_X1   g06680(.A1(new_n420_), .A2(new_n5112_), .B(new_n6957_), .ZN(new_n6958_));
  AOI21_X1   g06681(.A1(new_n6958_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n6959_));
  XOR2_X1    g06682(.A1(new_n700_), .A2(new_n6959_), .Z(new_n6960_));
  INV_X1     g06683(.I(new_n6960_), .ZN(new_n6961_));
  NAND3_X1   g06684(.A1(new_n6954_), .A2(new_n6956_), .A3(new_n6961_), .ZN(new_n6962_));
  AOI21_X1   g06685(.A1(new_n6955_), .A2(new_n6952_), .B(new_n6619_), .ZN(new_n6963_));
  NOR3_X1    g06686(.A1(new_n6947_), .A2(new_n6670_), .A3(new_n6953_), .ZN(new_n6964_));
  OAI21_X1   g06687(.A1(new_n6964_), .A2(new_n6963_), .B(new_n6960_), .ZN(new_n6965_));
  NAND2_X1   g06688(.A1(new_n6965_), .A2(new_n6962_), .ZN(new_n6966_));
  NAND3_X1   g06689(.A1(new_n6966_), .A2(new_n6681_), .A3(new_n6688_), .ZN(new_n6967_));
  NAND2_X1   g06690(.A1(new_n6675_), .A2(new_n6680_), .ZN(new_n6969_));
  AOI21_X1   g06691(.A1(new_n6967_), .A2(new_n6969_), .B(new_n6908_), .ZN(new_n6970_));
  INV_X1     g06692(.I(new_n6908_), .ZN(new_n6971_));
  INV_X1     g06693(.I(new_n6681_), .ZN(new_n6972_));
  NOR3_X1    g06694(.A1(new_n6964_), .A2(new_n6963_), .A3(new_n6960_), .ZN(new_n6973_));
  AOI21_X1   g06695(.A1(new_n6954_), .A2(new_n6956_), .B(new_n6961_), .ZN(new_n6974_));
  OAI21_X1   g06696(.A1(new_n6973_), .A2(new_n6974_), .B(new_n6688_), .ZN(new_n6975_));
  NOR2_X1    g06697(.A1(new_n6975_), .A2(new_n6972_), .ZN(new_n6976_));
  INV_X1     g06698(.I(new_n6969_), .ZN(new_n6977_));
  NOR3_X1    g06699(.A1(new_n6976_), .A2(new_n6971_), .A3(new_n6977_), .ZN(new_n6978_));
  OAI22_X1   g06700(.A1(new_n4072_), .A2(new_n656_), .B1(new_n706_), .B2(new_n4067_), .ZN(new_n6979_));
  OAI21_X1   g06701(.A1(new_n565_), .A2(new_n4318_), .B(new_n6979_), .ZN(new_n6980_));
  AOI21_X1   g06702(.A1(new_n6980_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n6981_));
  XNOR2_X1   g06703(.A1(new_n710_), .A2(new_n6981_), .ZN(new_n6982_));
  NOR3_X1    g06704(.A1(new_n6978_), .A2(new_n6970_), .A3(new_n6982_), .ZN(new_n6983_));
  OAI21_X1   g06705(.A1(new_n6976_), .A2(new_n6977_), .B(new_n6971_), .ZN(new_n6984_));
  NAND3_X1   g06706(.A1(new_n6967_), .A2(new_n6908_), .A3(new_n6969_), .ZN(new_n6985_));
  INV_X1     g06707(.I(new_n6982_), .ZN(new_n6986_));
  AOI21_X1   g06708(.A1(new_n6984_), .A2(new_n6985_), .B(new_n6986_), .ZN(new_n6987_));
  OAI22_X1   g06709(.A1(new_n861_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n930_), .ZN(new_n6988_));
  OAI21_X1   g06710(.A1(new_n780_), .A2(new_n3569_), .B(new_n6988_), .ZN(new_n6989_));
  AOI21_X1   g06711(.A1(new_n6989_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n6990_));
  XNOR2_X1   g06712(.A1(new_n937_), .A2(new_n6990_), .ZN(new_n6991_));
  INV_X1     g06713(.I(new_n6991_), .ZN(new_n6992_));
  OAI21_X1   g06714(.A1(new_n6983_), .A2(new_n6987_), .B(new_n6992_), .ZN(new_n6993_));
  NAND3_X1   g06715(.A1(new_n6984_), .A2(new_n6985_), .A3(new_n6986_), .ZN(new_n6994_));
  OAI21_X1   g06716(.A1(new_n6978_), .A2(new_n6970_), .B(new_n6982_), .ZN(new_n6995_));
  NAND3_X1   g06717(.A1(new_n6995_), .A2(new_n6994_), .A3(new_n6991_), .ZN(new_n6996_));
  AOI21_X1   g06718(.A1(new_n6993_), .A2(new_n6996_), .B(new_n6907_), .ZN(new_n6997_));
  INV_X1     g06719(.I(new_n6697_), .ZN(new_n6998_));
  OAI21_X1   g06720(.A1(new_n6610_), .A2(new_n6998_), .B(new_n6695_), .ZN(new_n6999_));
  NAND3_X1   g06721(.A1(new_n6995_), .A2(new_n6994_), .A3(new_n6992_), .ZN(new_n7000_));
  OAI21_X1   g06722(.A1(new_n6983_), .A2(new_n6987_), .B(new_n6991_), .ZN(new_n7001_));
  AOI21_X1   g06723(.A1(new_n7001_), .A2(new_n7000_), .B(new_n6999_), .ZN(new_n7002_));
  NOR2_X1    g06724(.A1(new_n6997_), .A2(new_n7002_), .ZN(new_n7003_));
  NOR3_X1    g06725(.A1(new_n7003_), .A2(new_n6719_), .A3(new_n6905_), .ZN(new_n7004_));
  NAND2_X1   g06726(.A1(new_n6995_), .A2(new_n6994_), .ZN(new_n7005_));
  INV_X1     g06727(.I(new_n7005_), .ZN(new_n7006_));
  NOR2_X1    g06728(.A1(new_n6904_), .A2(new_n6712_), .ZN(new_n7007_));
  OAI21_X1   g06729(.A1(new_n7004_), .A2(new_n7007_), .B(new_n6604_), .ZN(new_n7008_));
  NAND2_X1   g06730(.A1(new_n6716_), .A2(new_n6715_), .ZN(new_n7009_));
  NAND2_X1   g06731(.A1(new_n7009_), .A2(new_n6717_), .ZN(new_n7010_));
  AOI21_X1   g06732(.A1(new_n6995_), .A2(new_n6994_), .B(new_n6991_), .ZN(new_n7011_));
  NOR3_X1    g06733(.A1(new_n6983_), .A2(new_n6987_), .A3(new_n6992_), .ZN(new_n7012_));
  OAI21_X1   g06734(.A1(new_n7012_), .A2(new_n7011_), .B(new_n6999_), .ZN(new_n7013_));
  NOR3_X1    g06735(.A1(new_n6983_), .A2(new_n6987_), .A3(new_n6991_), .ZN(new_n7014_));
  AOI21_X1   g06736(.A1(new_n6995_), .A2(new_n6994_), .B(new_n6992_), .ZN(new_n7015_));
  OAI21_X1   g06737(.A1(new_n7014_), .A2(new_n7015_), .B(new_n6907_), .ZN(new_n7016_));
  NAND2_X1   g06738(.A1(new_n7016_), .A2(new_n7013_), .ZN(new_n7017_));
  NAND3_X1   g06739(.A1(new_n7017_), .A2(new_n6728_), .A3(new_n7010_), .ZN(new_n7018_));
  INV_X1     g06740(.I(new_n7007_), .ZN(new_n7019_));
  NAND3_X1   g06741(.A1(new_n7018_), .A2(new_n6735_), .A3(new_n7019_), .ZN(new_n7020_));
  OAI22_X1   g06742(.A1(new_n1109_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1189_), .ZN(new_n7021_));
  OAI21_X1   g06743(.A1(new_n1017_), .A2(new_n2884_), .B(new_n7021_), .ZN(new_n7022_));
  AOI21_X1   g06744(.A1(new_n7022_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n7023_));
  XNOR2_X1   g06745(.A1(new_n1196_), .A2(new_n7023_), .ZN(new_n7024_));
  AOI21_X1   g06746(.A1(new_n7008_), .A2(new_n7020_), .B(new_n7024_), .ZN(new_n7025_));
  AOI21_X1   g06747(.A1(new_n7018_), .A2(new_n7019_), .B(new_n6735_), .ZN(new_n7026_));
  NOR3_X1    g06748(.A1(new_n7004_), .A2(new_n6604_), .A3(new_n7007_), .ZN(new_n7027_));
  INV_X1     g06749(.I(new_n7024_), .ZN(new_n7028_));
  NOR3_X1    g06750(.A1(new_n7027_), .A2(new_n7026_), .A3(new_n7028_), .ZN(new_n7029_));
  NOR3_X1    g06751(.A1(new_n7029_), .A2(new_n7025_), .A3(new_n6903_), .ZN(new_n7030_));
  NOR3_X1    g06752(.A1(new_n7030_), .A2(new_n6599_), .A3(new_n6739_), .ZN(new_n7031_));
  NOR2_X1    g06753(.A1(new_n6604_), .A2(new_n6719_), .ZN(new_n7032_));
  NOR2_X1    g06754(.A1(new_n6735_), .A2(new_n6728_), .ZN(new_n7033_));
  OAI21_X1   g06755(.A1(new_n7033_), .A2(new_n7032_), .B(new_n6723_), .ZN(new_n7034_));
  OAI21_X1   g06756(.A1(new_n7027_), .A2(new_n7026_), .B(new_n7028_), .ZN(new_n7035_));
  NAND3_X1   g06757(.A1(new_n7008_), .A2(new_n7020_), .A3(new_n7024_), .ZN(new_n7036_));
  NAND3_X1   g06758(.A1(new_n7035_), .A2(new_n7036_), .A3(new_n7034_), .ZN(new_n7037_));
  AOI21_X1   g06759(.A1(new_n7037_), .A2(new_n6745_), .B(new_n6749_), .ZN(new_n7038_));
  OAI22_X1   g06760(.A1(new_n2171_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n2166_), .ZN(new_n7039_));
  OAI21_X1   g06761(.A1(new_n1294_), .A2(new_n2322_), .B(new_n7039_), .ZN(new_n7040_));
  AOI21_X1   g06762(.A1(new_n7040_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n7041_));
  XOR2_X1    g06763(.A1(new_n1530_), .A2(new_n7041_), .Z(new_n7042_));
  NOR3_X1    g06764(.A1(new_n7031_), .A2(new_n7038_), .A3(new_n7042_), .ZN(new_n7043_));
  NAND3_X1   g06765(.A1(new_n7037_), .A2(new_n6749_), .A3(new_n6745_), .ZN(new_n7044_));
  OAI21_X1   g06766(.A1(new_n7030_), .A2(new_n6739_), .B(new_n6599_), .ZN(new_n7045_));
  INV_X1     g06767(.I(new_n7042_), .ZN(new_n7046_));
  AOI21_X1   g06768(.A1(new_n7045_), .A2(new_n7044_), .B(new_n7046_), .ZN(new_n7047_));
  NOR3_X1    g06769(.A1(new_n7043_), .A2(new_n7047_), .A3(new_n6900_), .ZN(new_n7048_));
  NOR3_X1    g06770(.A1(new_n7048_), .A2(new_n6593_), .A3(new_n6896_), .ZN(new_n7049_));
  AOI21_X1   g06771(.A1(new_n6409_), .A2(new_n6410_), .B(new_n6283_), .ZN(new_n7050_));
  NOR3_X1    g06772(.A1(new_n6395_), .A2(new_n6399_), .A3(new_n6414_), .ZN(new_n7051_));
  NOR2_X1    g06773(.A1(new_n7051_), .A2(new_n6403_), .ZN(new_n7052_));
  AOI21_X1   g06774(.A1(new_n7052_), .A2(new_n6285_), .B(new_n7050_), .ZN(new_n7053_));
  INV_X1     g06775(.I(new_n6897_), .ZN(new_n7054_));
  OAI21_X1   g06776(.A1(new_n7054_), .A2(new_n6898_), .B(new_n6743_), .ZN(new_n7055_));
  NAND3_X1   g06777(.A1(new_n7045_), .A2(new_n7044_), .A3(new_n7046_), .ZN(new_n7056_));
  OAI21_X1   g06778(.A1(new_n7031_), .A2(new_n7038_), .B(new_n7042_), .ZN(new_n7057_));
  NAND3_X1   g06779(.A1(new_n7057_), .A2(new_n7056_), .A3(new_n7055_), .ZN(new_n7058_));
  AOI21_X1   g06780(.A1(new_n7058_), .A2(new_n6753_), .B(new_n7053_), .ZN(new_n7059_));
  NOR2_X1    g06781(.A1(new_n7059_), .A2(new_n7049_), .ZN(new_n7060_));
  NOR2_X1    g06782(.A1(new_n6593_), .A2(new_n6896_), .ZN(new_n7061_));
  NOR2_X1    g06783(.A1(new_n7053_), .A2(new_n6753_), .ZN(new_n7062_));
  OAI21_X1   g06784(.A1(new_n7062_), .A2(new_n7061_), .B(new_n6757_), .ZN(new_n7063_));
  NAND3_X1   g06785(.A1(new_n6588_), .A2(new_n6765_), .A3(new_n6586_), .ZN(new_n7064_));
  OAI22_X1   g06786(.A1(new_n1347_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n1344_), .ZN(new_n7065_));
  OAI21_X1   g06787(.A1(new_n2102_), .A2(new_n1457_), .B(new_n7065_), .ZN(new_n7066_));
  AOI21_X1   g06788(.A1(new_n7066_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n7067_));
  XNOR2_X1   g06789(.A1(new_n2443_), .A2(new_n7067_), .ZN(new_n7068_));
  AOI21_X1   g06790(.A1(new_n7064_), .A2(new_n7063_), .B(new_n7068_), .ZN(new_n7069_));
  INV_X1     g06791(.I(new_n7063_), .ZN(new_n7070_));
  AOI21_X1   g06792(.A1(new_n6416_), .A2(new_n6415_), .B(new_n6414_), .ZN(new_n7071_));
  NOR3_X1    g06793(.A1(new_n6406_), .A2(new_n6412_), .A3(new_n6283_), .ZN(new_n7072_));
  NOR3_X1    g06794(.A1(new_n7071_), .A2(new_n7072_), .A3(new_n6126_), .ZN(new_n7073_));
  NOR3_X1    g06795(.A1(new_n6427_), .A2(new_n7073_), .A3(new_n6422_), .ZN(new_n7074_));
  NAND2_X1   g06796(.A1(new_n6761_), .A2(new_n6593_), .ZN(new_n7075_));
  NAND2_X1   g06797(.A1(new_n6763_), .A2(new_n6762_), .ZN(new_n7076_));
  NAND2_X1   g06798(.A1(new_n7076_), .A2(new_n7053_), .ZN(new_n7077_));
  NAND2_X1   g06799(.A1(new_n7075_), .A2(new_n7077_), .ZN(new_n7078_));
  NOR3_X1    g06800(.A1(new_n7074_), .A2(new_n6585_), .A3(new_n7078_), .ZN(new_n7079_));
  INV_X1     g06801(.I(new_n7068_), .ZN(new_n7080_));
  NOR3_X1    g06802(.A1(new_n7079_), .A2(new_n7070_), .A3(new_n7080_), .ZN(new_n7081_));
  OAI21_X1   g06803(.A1(new_n7081_), .A2(new_n7069_), .B(new_n7060_), .ZN(new_n7082_));
  NAND3_X1   g06804(.A1(new_n7058_), .A2(new_n7053_), .A3(new_n6753_), .ZN(new_n7083_));
  OAI21_X1   g06805(.A1(new_n7048_), .A2(new_n6896_), .B(new_n6593_), .ZN(new_n7084_));
  NAND2_X1   g06806(.A1(new_n7084_), .A2(new_n7083_), .ZN(new_n7085_));
  OAI21_X1   g06807(.A1(new_n7079_), .A2(new_n7070_), .B(new_n7080_), .ZN(new_n7086_));
  NAND3_X1   g06808(.A1(new_n7064_), .A2(new_n7063_), .A3(new_n7068_), .ZN(new_n7087_));
  NAND3_X1   g06809(.A1(new_n7086_), .A2(new_n7087_), .A3(new_n7085_), .ZN(new_n7088_));
  AOI21_X1   g06810(.A1(new_n7082_), .A2(new_n7088_), .B(new_n6895_), .ZN(new_n7089_));
  AOI21_X1   g06811(.A1(new_n7086_), .A2(new_n7087_), .B(new_n7085_), .ZN(new_n7090_));
  NOR3_X1    g06812(.A1(new_n7081_), .A2(new_n7069_), .A3(new_n7060_), .ZN(new_n7091_));
  NOR3_X1    g06813(.A1(new_n7091_), .A2(new_n7090_), .A3(new_n6894_), .ZN(new_n7092_));
  NOR3_X1    g06814(.A1(new_n7092_), .A2(new_n7089_), .A3(new_n6890_), .ZN(new_n7093_));
  NOR3_X1    g06815(.A1(new_n7093_), .A2(new_n6583_), .A3(new_n6782_), .ZN(new_n7094_));
  XOR2_X1    g06816(.A1(new_n6589_), .A2(new_n7078_), .Z(new_n7095_));
  NAND2_X1   g06817(.A1(new_n7095_), .A2(new_n6769_), .ZN(new_n7096_));
  OAI21_X1   g06818(.A1(new_n7091_), .A2(new_n7090_), .B(new_n6894_), .ZN(new_n7097_));
  NAND3_X1   g06819(.A1(new_n7082_), .A2(new_n7088_), .A3(new_n6895_), .ZN(new_n7098_));
  NAND3_X1   g06820(.A1(new_n7097_), .A2(new_n7098_), .A3(new_n7096_), .ZN(new_n7099_));
  AOI21_X1   g06821(.A1(new_n7099_), .A2(new_n6774_), .B(new_n6584_), .ZN(new_n7100_));
  OAI22_X1   g06822(.A1(new_n1055_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n1061_), .ZN(new_n7101_));
  OAI21_X1   g06823(.A1(new_n2643_), .A2(new_n1332_), .B(new_n7101_), .ZN(new_n7102_));
  AOI21_X1   g06824(.A1(new_n7102_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n7103_));
  XNOR2_X1   g06825(.A1(new_n3022_), .A2(new_n7103_), .ZN(new_n7104_));
  INV_X1     g06826(.I(new_n7104_), .ZN(new_n7105_));
  OAI21_X1   g06827(.A1(new_n7094_), .A2(new_n7100_), .B(new_n7105_), .ZN(new_n7106_));
  NAND3_X1   g06828(.A1(new_n7099_), .A2(new_n6584_), .A3(new_n6774_), .ZN(new_n7107_));
  OAI21_X1   g06829(.A1(new_n7093_), .A2(new_n6782_), .B(new_n6583_), .ZN(new_n7108_));
  NAND3_X1   g06830(.A1(new_n7108_), .A2(new_n7107_), .A3(new_n7104_), .ZN(new_n7109_));
  NAND3_X1   g06831(.A1(new_n6888_), .A2(new_n7106_), .A3(new_n7109_), .ZN(new_n7110_));
  NAND3_X1   g06832(.A1(new_n7110_), .A2(new_n6791_), .A3(new_n6788_), .ZN(new_n7111_));
  AOI21_X1   g06833(.A1(new_n7108_), .A2(new_n7107_), .B(new_n7104_), .ZN(new_n7112_));
  NOR3_X1    g06834(.A1(new_n7094_), .A2(new_n7100_), .A3(new_n7105_), .ZN(new_n7113_));
  NOR3_X1    g06835(.A1(new_n7113_), .A2(new_n7112_), .A3(new_n6887_), .ZN(new_n7114_));
  OAI21_X1   g06836(.A1(new_n7114_), .A2(new_n6794_), .B(new_n6579_), .ZN(new_n7115_));
  OAI22_X1   g06837(.A1(new_n970_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n820_), .ZN(new_n7116_));
  OAI21_X1   g06838(.A1(new_n3260_), .A2(new_n894_), .B(new_n7116_), .ZN(new_n7117_));
  AOI21_X1   g06839(.A1(new_n7117_), .A2(new_n827_), .B(new_n970_), .ZN(new_n7118_));
  XOR2_X1    g06840(.A1(new_n3722_), .A2(new_n7118_), .Z(new_n7119_));
  AOI21_X1   g06841(.A1(new_n7111_), .A2(new_n7115_), .B(new_n7119_), .ZN(new_n7120_));
  NOR3_X1    g06842(.A1(new_n7114_), .A2(new_n6579_), .A3(new_n6794_), .ZN(new_n7121_));
  AOI21_X1   g06843(.A1(new_n7110_), .A2(new_n6788_), .B(new_n6791_), .ZN(new_n7122_));
  INV_X1     g06844(.I(new_n7119_), .ZN(new_n7123_));
  NOR3_X1    g06845(.A1(new_n7122_), .A2(new_n7121_), .A3(new_n7123_), .ZN(new_n7124_));
  OAI21_X1   g06846(.A1(new_n7120_), .A2(new_n7124_), .B(new_n6805_), .ZN(new_n7125_));
  NOR2_X1    g06847(.A1(new_n7125_), .A2(new_n6884_), .ZN(new_n7126_));
  OAI21_X1   g06848(.A1(new_n7122_), .A2(new_n7121_), .B(new_n7123_), .ZN(new_n7127_));
  NAND3_X1   g06849(.A1(new_n7111_), .A2(new_n7115_), .A3(new_n7119_), .ZN(new_n7128_));
  NAND2_X1   g06850(.A1(new_n7127_), .A2(new_n7128_), .ZN(new_n7129_));
  NOR2_X1    g06851(.A1(new_n6883_), .A2(new_n6799_), .ZN(new_n7131_));
  OAI21_X1   g06852(.A1(new_n7126_), .A2(new_n7131_), .B(new_n6576_), .ZN(new_n7132_));
  INV_X1     g06853(.I(new_n6884_), .ZN(new_n7133_));
  NAND3_X1   g06854(.A1(new_n7129_), .A2(new_n6805_), .A3(new_n7133_), .ZN(new_n7134_));
  INV_X1     g06855(.I(new_n7131_), .ZN(new_n7135_));
  NAND3_X1   g06856(.A1(new_n7134_), .A2(new_n6575_), .A3(new_n7135_), .ZN(new_n7136_));
  OAI22_X1   g06857(.A1(new_n607_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n610_), .ZN(new_n7137_));
  OAI21_X1   g06858(.A1(new_n3989_), .A2(new_n684_), .B(new_n7137_), .ZN(new_n7138_));
  AOI21_X1   g06859(.A1(new_n7138_), .A2(new_n612_), .B(new_n607_), .ZN(new_n7139_));
  XOR2_X1    g06860(.A1(new_n4499_), .A2(new_n7139_), .Z(new_n7140_));
  INV_X1     g06861(.I(new_n7140_), .ZN(new_n7141_));
  NAND3_X1   g06862(.A1(new_n7132_), .A2(new_n7136_), .A3(new_n7141_), .ZN(new_n7142_));
  AOI21_X1   g06863(.A1(new_n7134_), .A2(new_n7135_), .B(new_n6575_), .ZN(new_n7143_));
  NOR3_X1    g06864(.A1(new_n7126_), .A2(new_n6576_), .A3(new_n7131_), .ZN(new_n7144_));
  OAI21_X1   g06865(.A1(new_n7144_), .A2(new_n7143_), .B(new_n7140_), .ZN(new_n7145_));
  NAND3_X1   g06866(.A1(new_n7145_), .A2(new_n7142_), .A3(new_n6882_), .ZN(new_n7146_));
  NAND3_X1   g06867(.A1(new_n7146_), .A2(new_n6568_), .A3(new_n6832_), .ZN(new_n7147_));
  OR3_X2     g06868(.A1(new_n6257_), .A2(new_n5961_), .A3(new_n6258_), .Z(new_n7148_));
  OAI21_X1   g06869(.A1(new_n6565_), .A2(new_n6255_), .B(new_n6492_), .ZN(new_n7149_));
  OAI22_X1   g06870(.A1(new_n7148_), .A2(new_n7149_), .B1(new_n6256_), .B2(new_n6566_), .ZN(new_n7150_));
  INV_X1     g06871(.I(new_n6881_), .ZN(new_n7151_));
  AOI21_X1   g06872(.A1(new_n7151_), .A2(new_n6879_), .B(new_n6812_), .ZN(new_n7152_));
  NOR3_X1    g06873(.A1(new_n7144_), .A2(new_n7143_), .A3(new_n7140_), .ZN(new_n7153_));
  AOI21_X1   g06874(.A1(new_n7132_), .A2(new_n7136_), .B(new_n7141_), .ZN(new_n7154_));
  NOR3_X1    g06875(.A1(new_n7153_), .A2(new_n7154_), .A3(new_n7152_), .ZN(new_n7155_));
  OAI21_X1   g06876(.A1(new_n7155_), .A2(new_n6815_), .B(new_n7150_), .ZN(new_n7156_));
  OAI22_X1   g06877(.A1(new_n448_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n450_), .ZN(new_n7157_));
  OAI21_X1   g06878(.A1(new_n4774_), .A2(new_n496_), .B(new_n7157_), .ZN(new_n7158_));
  AOI21_X1   g06879(.A1(new_n7158_), .A2(new_n452_), .B(new_n448_), .ZN(new_n7159_));
  XNOR2_X1   g06880(.A1(new_n5357_), .A2(new_n7159_), .ZN(new_n7160_));
  INV_X1     g06881(.I(new_n7160_), .ZN(new_n7161_));
  NAND3_X1   g06882(.A1(new_n7156_), .A2(new_n7147_), .A3(new_n7161_), .ZN(new_n7162_));
  NOR3_X1    g06883(.A1(new_n7155_), .A2(new_n7150_), .A3(new_n6815_), .ZN(new_n7163_));
  AOI21_X1   g06884(.A1(new_n7146_), .A2(new_n6832_), .B(new_n6568_), .ZN(new_n7164_));
  OAI21_X1   g06885(.A1(new_n7163_), .A2(new_n7164_), .B(new_n7160_), .ZN(new_n7165_));
  NAND2_X1   g06886(.A1(new_n7165_), .A2(new_n7162_), .ZN(new_n7166_));
  OAI22_X1   g06887(.A1(new_n5921_), .A2(new_n341_), .B1(new_n404_), .B2(new_n6229_), .ZN(new_n7167_));
  OAI21_X1   g06888(.A1(new_n5913_), .A2(new_n366_), .B(new_n7167_), .ZN(new_n7168_));
  AOI21_X1   g06889(.A1(new_n7168_), .A2(new_n334_), .B(new_n341_), .ZN(new_n7169_));
  XOR2_X1    g06890(.A1(new_n6233_), .A2(new_n7169_), .Z(new_n7170_));
  XOR2_X1    g06891(.A1(new_n7166_), .A2(new_n7170_), .Z(new_n7171_));
  NAND2_X1   g06892(.A1(new_n7171_), .A2(new_n6878_), .ZN(new_n7172_));
  XOR2_X1    g06893(.A1(new_n7166_), .A2(new_n7170_), .Z(new_n7173_));
  OAI21_X1   g06894(.A1(new_n6878_), .A2(new_n7173_), .B(new_n7172_), .ZN(new_n7174_));
  INV_X1     g06895(.I(new_n7174_), .ZN(new_n7175_));
  AOI21_X1   g06896(.A1(new_n6842_), .A2(new_n6522_), .B(new_n6248_), .ZN(new_n7176_));
  NAND3_X1   g06897(.A1(new_n6837_), .A2(new_n6841_), .A3(new_n6521_), .ZN(new_n7177_));
  NAND2_X1   g06898(.A1(new_n6528_), .A2(new_n7177_), .ZN(new_n7178_));
  OR2_X2     g06899(.A1(new_n7178_), .A2(new_n7176_), .Z(new_n7179_));
  NAND2_X1   g06900(.A1(new_n6819_), .A2(new_n6816_), .ZN(new_n7180_));
  NAND2_X1   g06901(.A1(new_n6829_), .A2(new_n6833_), .ZN(new_n7181_));
  NAND2_X1   g06902(.A1(new_n7180_), .A2(new_n7181_), .ZN(new_n7182_));
  NAND2_X1   g06903(.A1(new_n7182_), .A2(new_n6564_), .ZN(new_n7183_));
  NAND3_X1   g06904(.A1(new_n7180_), .A2(new_n7181_), .A3(new_n6838_), .ZN(new_n7184_));
  AOI21_X1   g06905(.A1(new_n7183_), .A2(new_n7184_), .B(new_n6823_), .ZN(new_n7185_));
  INV_X1     g06906(.I(new_n7185_), .ZN(new_n7186_));
  NAND2_X1   g06907(.A1(new_n7179_), .A2(new_n7186_), .ZN(new_n7187_));
  NAND2_X1   g06908(.A1(new_n7187_), .A2(new_n7175_), .ZN(new_n7188_));
  NAND3_X1   g06909(.A1(new_n7179_), .A2(new_n7174_), .A3(new_n7186_), .ZN(new_n7189_));
  NAND2_X1   g06910(.A1(new_n7188_), .A2(new_n7189_), .ZN(new_n7190_));
  NOR2_X1    g06911(.A1(\b[42] ), .A2(\b[43] ), .ZN(new_n7191_));
  AOI21_X1   g06912(.A1(new_n6534_), .A2(new_n7191_), .B(new_n6229_), .ZN(new_n7192_));
  NOR2_X1    g06913(.A1(new_n6538_), .A2(new_n6847_), .ZN(new_n7193_));
  INV_X1     g06914(.I(new_n7193_), .ZN(new_n7194_));
  NOR2_X1    g06915(.A1(new_n6534_), .A2(new_n7194_), .ZN(new_n7195_));
  NOR2_X1    g06916(.A1(new_n7192_), .A2(new_n7195_), .ZN(new_n7196_));
  XNOR2_X1   g06917(.A1(\b[43] ), .A2(\b[44] ), .ZN(new_n7197_));
  INV_X1     g06918(.I(\b[44] ), .ZN(new_n7198_));
  NOR2_X1    g06919(.A1(new_n6847_), .A2(new_n7198_), .ZN(new_n7199_));
  NOR2_X1    g06920(.A1(\b[43] ), .A2(\b[44] ), .ZN(new_n7200_));
  OAI21_X1   g06921(.A1(new_n7199_), .A2(new_n7200_), .B(new_n7196_), .ZN(new_n7201_));
  OAI21_X1   g06922(.A1(new_n7196_), .A2(new_n7197_), .B(new_n7201_), .ZN(new_n7202_));
  OAI22_X1   g06923(.A1(new_n330_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n263_), .ZN(new_n7203_));
  OAI21_X1   g06924(.A1(new_n6538_), .A2(new_n289_), .B(new_n7203_), .ZN(new_n7204_));
  AOI21_X1   g06925(.A1(new_n7204_), .A2(new_n260_), .B(new_n426_), .ZN(new_n7205_));
  XNOR2_X1   g06926(.A1(new_n7202_), .A2(new_n7205_), .ZN(new_n7206_));
  XOR2_X1    g06927(.A1(new_n7190_), .A2(new_n7206_), .Z(new_n7207_));
  XOR2_X1    g06928(.A1(new_n7190_), .A2(new_n7206_), .Z(new_n7208_));
  NAND2_X1   g06929(.A1(new_n6875_), .A2(new_n7208_), .ZN(new_n7209_));
  OAI21_X1   g06930(.A1(new_n6875_), .A2(new_n7207_), .B(new_n7209_), .ZN(\f[44] ));
  INV_X1     g06931(.I(new_n7206_), .ZN(new_n7211_));
  NAND2_X1   g06932(.A1(new_n7190_), .A2(new_n7211_), .ZN(new_n7212_));
  INV_X1     g06933(.I(new_n7170_), .ZN(new_n7213_));
  NAND3_X1   g06934(.A1(new_n6877_), .A2(new_n6876_), .A3(new_n7166_), .ZN(new_n7214_));
  NOR3_X1    g06935(.A1(new_n7163_), .A2(new_n7164_), .A3(new_n7160_), .ZN(new_n7215_));
  AOI21_X1   g06936(.A1(new_n7156_), .A2(new_n7147_), .B(new_n7161_), .ZN(new_n7216_));
  NOR2_X1    g06937(.A1(new_n7215_), .A2(new_n7216_), .ZN(new_n7217_));
  NAND2_X1   g06938(.A1(new_n6878_), .A2(new_n7217_), .ZN(new_n7218_));
  AOI21_X1   g06939(.A1(new_n7218_), .A2(new_n7214_), .B(new_n7213_), .ZN(new_n7219_));
  AOI21_X1   g06940(.A1(new_n7174_), .A2(new_n7219_), .B(new_n7185_), .ZN(new_n7220_));
  OR3_X2     g06941(.A1(new_n7220_), .A2(new_n7178_), .A3(new_n7176_), .Z(new_n7221_));
  OAI21_X1   g06942(.A1(new_n7217_), .A2(new_n6833_), .B(new_n6564_), .ZN(new_n7222_));
  NOR3_X1    g06943(.A1(new_n7215_), .A2(new_n7216_), .A3(new_n6816_), .ZN(new_n7223_));
  NOR2_X1    g06944(.A1(new_n7223_), .A2(new_n6819_), .ZN(new_n7224_));
  NAND2_X1   g06945(.A1(new_n7224_), .A2(new_n7222_), .ZN(new_n7225_));
  OAI21_X1   g06946(.A1(new_n7153_), .A2(new_n7154_), .B(new_n7152_), .ZN(new_n7226_));
  AOI21_X1   g06947(.A1(new_n7226_), .A2(new_n6815_), .B(new_n6568_), .ZN(new_n7227_));
  OAI21_X1   g06948(.A1(new_n7122_), .A2(new_n7121_), .B(new_n7119_), .ZN(new_n7228_));
  INV_X1     g06949(.I(new_n7228_), .ZN(new_n7229_));
  INV_X1     g06950(.I(new_n6883_), .ZN(new_n7230_));
  AOI21_X1   g06951(.A1(new_n7129_), .A2(new_n6800_), .B(new_n7230_), .ZN(new_n7231_));
  OAI21_X1   g06952(.A1(new_n6800_), .A2(new_n7129_), .B(new_n6575_), .ZN(new_n7232_));
  AOI21_X1   g06953(.A1(new_n7108_), .A2(new_n7107_), .B(new_n7105_), .ZN(new_n7233_));
  INV_X1     g06954(.I(new_n7233_), .ZN(new_n7234_));
  OAI21_X1   g06955(.A1(new_n7113_), .A2(new_n7112_), .B(new_n6887_), .ZN(new_n7235_));
  AOI21_X1   g06956(.A1(new_n7235_), .A2(new_n6794_), .B(new_n6791_), .ZN(new_n7236_));
  NOR2_X1    g06957(.A1(new_n7079_), .A2(new_n7070_), .ZN(new_n7237_));
  NOR2_X1    g06958(.A1(new_n7237_), .A2(new_n7060_), .ZN(new_n7238_));
  NAND2_X1   g06959(.A1(new_n7064_), .A2(new_n7063_), .ZN(new_n7239_));
  NOR2_X1    g06960(.A1(new_n7239_), .A2(new_n7085_), .ZN(new_n7240_));
  OAI21_X1   g06961(.A1(new_n7238_), .A2(new_n7240_), .B(new_n6894_), .ZN(new_n7241_));
  NAND2_X1   g06962(.A1(new_n7239_), .A2(new_n7085_), .ZN(new_n7242_));
  NAND2_X1   g06963(.A1(new_n7237_), .A2(new_n7060_), .ZN(new_n7243_));
  NAND3_X1   g06964(.A1(new_n7243_), .A2(new_n7242_), .A3(new_n6895_), .ZN(new_n7244_));
  AOI21_X1   g06965(.A1(new_n7241_), .A2(new_n7244_), .B(new_n7068_), .ZN(new_n7245_));
  AOI21_X1   g06966(.A1(new_n7097_), .A2(new_n7098_), .B(new_n7096_), .ZN(new_n7246_));
  OAI21_X1   g06967(.A1(new_n7246_), .A2(new_n6774_), .B(new_n6583_), .ZN(new_n7247_));
  NOR2_X1    g06968(.A1(new_n7060_), .A2(new_n6895_), .ZN(new_n7248_));
  INV_X1     g06969(.I(new_n7248_), .ZN(new_n7249_));
  NOR2_X1    g06970(.A1(new_n7060_), .A2(new_n6894_), .ZN(new_n7250_));
  NOR2_X1    g06971(.A1(new_n7085_), .A2(new_n6895_), .ZN(new_n7251_));
  OAI21_X1   g06972(.A1(new_n7250_), .A2(new_n7251_), .B(new_n7070_), .ZN(new_n7252_));
  AOI22_X1   g06973(.A1(new_n7252_), .A2(new_n6765_), .B1(new_n6586_), .B2(new_n6588_), .ZN(new_n7253_));
  AOI21_X1   g06974(.A1(new_n7057_), .A2(new_n7056_), .B(new_n7055_), .ZN(new_n7254_));
  OAI21_X1   g06975(.A1(new_n7254_), .A2(new_n6753_), .B(new_n6593_), .ZN(new_n7255_));
  AOI21_X1   g06976(.A1(new_n7008_), .A2(new_n7020_), .B(new_n7028_), .ZN(new_n7256_));
  INV_X1     g06977(.I(new_n7256_), .ZN(new_n7257_));
  OAI21_X1   g06978(.A1(new_n7029_), .A2(new_n7025_), .B(new_n6903_), .ZN(new_n7258_));
  AOI21_X1   g06979(.A1(new_n7258_), .A2(new_n6739_), .B(new_n6749_), .ZN(new_n7259_));
  NAND2_X1   g06980(.A1(new_n6999_), .A2(new_n7005_), .ZN(new_n7260_));
  NAND2_X1   g06981(.A1(new_n7006_), .A2(new_n6907_), .ZN(new_n7261_));
  AOI21_X1   g06982(.A1(new_n7261_), .A2(new_n7260_), .B(new_n6992_), .ZN(new_n7262_));
  OAI21_X1   g06983(.A1(new_n7003_), .A2(new_n6712_), .B(new_n6904_), .ZN(new_n7263_));
  NAND3_X1   g06984(.A1(new_n7016_), .A2(new_n7013_), .A3(new_n6712_), .ZN(new_n7264_));
  NAND3_X1   g06985(.A1(new_n7263_), .A2(new_n6735_), .A3(new_n7264_), .ZN(new_n7265_));
  NOR3_X1    g06986(.A1(new_n6978_), .A2(new_n6970_), .A3(new_n6986_), .ZN(new_n7266_));
  INV_X1     g06987(.I(new_n7266_), .ZN(new_n7267_));
  NAND2_X1   g06988(.A1(new_n6685_), .A2(new_n6689_), .ZN(new_n7268_));
  OAI21_X1   g06989(.A1(new_n6983_), .A2(new_n6987_), .B(new_n7268_), .ZN(new_n7269_));
  NAND2_X1   g06990(.A1(new_n7269_), .A2(new_n6693_), .ZN(new_n7270_));
  NOR3_X1    g06991(.A1(new_n6983_), .A2(new_n6987_), .A3(new_n7268_), .ZN(new_n7271_));
  NOR2_X1    g06992(.A1(new_n7271_), .A2(new_n6610_), .ZN(new_n7272_));
  OAI21_X1   g06993(.A1(new_n6973_), .A2(new_n6974_), .B(new_n6675_), .ZN(new_n7273_));
  NAND2_X1   g06994(.A1(new_n7273_), .A2(new_n6679_), .ZN(new_n7274_));
  NAND3_X1   g06995(.A1(new_n6965_), .A2(new_n6962_), .A3(new_n6682_), .ZN(new_n7275_));
  NAND3_X1   g06996(.A1(new_n7274_), .A2(new_n6908_), .A3(new_n7275_), .ZN(new_n7276_));
  XOR2_X1    g06997(.A1(new_n6927_), .A2(new_n5681_), .Z(new_n7277_));
  XOR2_X1    g06998(.A1(new_n6938_), .A2(new_n6922_), .Z(new_n7278_));
  NAND2_X1   g06999(.A1(new_n7278_), .A2(new_n7277_), .ZN(new_n7279_));
  AOI21_X1   g07000(.A1(new_n6950_), .A2(new_n6658_), .B(new_n6628_), .ZN(new_n7280_));
  OAI21_X1   g07001(.A1(new_n6950_), .A2(new_n6658_), .B(new_n6619_), .ZN(new_n7281_));
  XOR2_X1    g07002(.A1(\a[41] ), .A2(\a[42] ), .Z(new_n7282_));
  XOR2_X1    g07003(.A1(\a[41] ), .A2(\a[44] ), .Z(new_n7283_));
  NAND3_X1   g07004(.A1(new_n6640_), .A2(new_n7282_), .A3(new_n7283_), .ZN(new_n7284_));
  NOR2_X1    g07005(.A1(new_n7284_), .A2(new_n269_), .ZN(new_n7285_));
  OAI22_X1   g07006(.A1(new_n6644_), .A2(new_n280_), .B1(new_n298_), .B2(new_n6647_), .ZN(new_n7286_));
  NOR2_X1    g07007(.A1(new_n7286_), .A2(new_n7285_), .ZN(new_n7287_));
  NAND2_X1   g07008(.A1(new_n301_), .A2(new_n6631_), .ZN(new_n7288_));
  OAI21_X1   g07009(.A1(new_n7287_), .A2(new_n7288_), .B(\a[44] ), .ZN(new_n7289_));
  INV_X1     g07010(.I(new_n7289_), .ZN(new_n7290_));
  NOR3_X1    g07011(.A1(new_n7287_), .A2(\a[44] ), .A3(new_n7288_), .ZN(new_n7291_));
  XNOR2_X1   g07012(.A1(\a[44] ), .A2(\a[45] ), .ZN(new_n7292_));
  NOR2_X1    g07013(.A1(new_n7292_), .A2(new_n258_), .ZN(new_n7293_));
  OAI21_X1   g07014(.A1(new_n7290_), .A2(new_n7291_), .B(new_n7293_), .ZN(new_n7294_));
  NOR2_X1    g07015(.A1(new_n7294_), .A2(new_n6938_), .ZN(new_n7295_));
  OR3_X2     g07016(.A1(new_n7287_), .A2(\a[44] ), .A3(new_n7288_), .Z(new_n7296_));
  INV_X1     g07017(.I(new_n7293_), .ZN(new_n7297_));
  AOI21_X1   g07018(.A1(new_n7296_), .A2(new_n7289_), .B(new_n7297_), .ZN(new_n7298_));
  NOR2_X1    g07019(.A1(new_n7298_), .A2(new_n6921_), .ZN(new_n7299_));
  OAI21_X1   g07020(.A1(new_n7295_), .A2(new_n7299_), .B(new_n6929_), .ZN(new_n7300_));
  NOR2_X1    g07021(.A1(new_n7295_), .A2(new_n7299_), .ZN(new_n7301_));
  NAND2_X1   g07022(.A1(new_n7301_), .A2(new_n6922_), .ZN(new_n7302_));
  AOI22_X1   g07023(.A1(new_n5680_), .A2(\b[5] ), .B1(\b[6] ), .B2(new_n5686_), .ZN(new_n7303_));
  AOI21_X1   g07024(.A1(\b[4] ), .A2(new_n6923_), .B(new_n7303_), .ZN(new_n7304_));
  OAI21_X1   g07025(.A1(new_n7304_), .A2(\a[41] ), .B(new_n5680_), .ZN(new_n7305_));
  XOR2_X1    g07026(.A1(new_n556_), .A2(new_n7305_), .Z(new_n7306_));
  AOI21_X1   g07027(.A1(new_n7302_), .A2(new_n7300_), .B(new_n7306_), .ZN(new_n7307_));
  OAI21_X1   g07028(.A1(new_n7280_), .A2(new_n7281_), .B(new_n7307_), .ZN(new_n7308_));
  INV_X1     g07029(.I(new_n7308_), .ZN(new_n7309_));
  NOR3_X1    g07030(.A1(new_n7280_), .A2(new_n7281_), .A3(new_n7307_), .ZN(new_n7310_));
  OAI21_X1   g07031(.A1(new_n7309_), .A2(new_n7310_), .B(new_n7279_), .ZN(new_n7311_));
  INV_X1     g07032(.I(new_n7279_), .ZN(new_n7312_));
  INV_X1     g07033(.I(new_n7310_), .ZN(new_n7313_));
  NAND3_X1   g07034(.A1(new_n7313_), .A2(new_n7312_), .A3(new_n7308_), .ZN(new_n7314_));
  OAI22_X1   g07035(.A1(new_n5420_), .A2(new_n515_), .B1(new_n565_), .B2(new_n5107_), .ZN(new_n7315_));
  OAI21_X1   g07036(.A1(new_n472_), .A2(new_n5112_), .B(new_n7315_), .ZN(new_n7316_));
  AOI21_X1   g07037(.A1(new_n7316_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n7317_));
  XOR2_X1    g07038(.A1(new_n759_), .A2(new_n7317_), .Z(new_n7318_));
  AOI21_X1   g07039(.A1(new_n7311_), .A2(new_n7314_), .B(new_n7318_), .ZN(new_n7319_));
  NAND2_X1   g07040(.A1(new_n7276_), .A2(new_n7319_), .ZN(new_n7320_));
  AOI21_X1   g07041(.A1(new_n6966_), .A2(new_n6675_), .B(new_n6680_), .ZN(new_n7321_));
  NAND2_X1   g07042(.A1(new_n7275_), .A2(new_n6908_), .ZN(new_n7322_));
  NOR2_X1    g07043(.A1(new_n7322_), .A2(new_n7321_), .ZN(new_n7323_));
  INV_X1     g07044(.I(new_n7319_), .ZN(new_n7324_));
  NAND2_X1   g07045(.A1(new_n7323_), .A2(new_n7324_), .ZN(new_n7325_));
  AOI21_X1   g07046(.A1(new_n7325_), .A2(new_n7320_), .B(new_n6974_), .ZN(new_n7326_));
  NOR2_X1    g07047(.A1(new_n7323_), .A2(new_n7324_), .ZN(new_n7327_));
  NOR2_X1    g07048(.A1(new_n7276_), .A2(new_n7319_), .ZN(new_n7328_));
  NOR3_X1    g07049(.A1(new_n7327_), .A2(new_n7328_), .A3(new_n6965_), .ZN(new_n7329_));
  OAI22_X1   g07050(.A1(new_n4072_), .A2(new_n706_), .B1(new_n780_), .B2(new_n4067_), .ZN(new_n7330_));
  OAI21_X1   g07051(.A1(new_n656_), .A2(new_n4318_), .B(new_n7330_), .ZN(new_n7331_));
  AOI21_X1   g07052(.A1(new_n7331_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n7332_));
  XOR2_X1    g07053(.A1(new_n785_), .A2(new_n7332_), .Z(new_n7333_));
  INV_X1     g07054(.I(new_n7333_), .ZN(new_n7334_));
  OAI21_X1   g07055(.A1(new_n7326_), .A2(new_n7329_), .B(new_n7334_), .ZN(new_n7335_));
  AOI21_X1   g07056(.A1(new_n7272_), .A2(new_n7270_), .B(new_n7335_), .ZN(new_n7336_));
  AOI21_X1   g07057(.A1(new_n7005_), .A2(new_n7268_), .B(new_n6694_), .ZN(new_n7337_));
  OAI21_X1   g07058(.A1(new_n7005_), .A2(new_n7268_), .B(new_n6703_), .ZN(new_n7338_));
  OAI21_X1   g07059(.A1(new_n7327_), .A2(new_n7328_), .B(new_n6965_), .ZN(new_n7339_));
  NAND3_X1   g07060(.A1(new_n7325_), .A2(new_n7320_), .A3(new_n6974_), .ZN(new_n7340_));
  AOI21_X1   g07061(.A1(new_n7339_), .A2(new_n7340_), .B(new_n7333_), .ZN(new_n7341_));
  NOR3_X1    g07062(.A1(new_n7337_), .A2(new_n7338_), .A3(new_n7341_), .ZN(new_n7342_));
  OAI21_X1   g07063(.A1(new_n7336_), .A2(new_n7342_), .B(new_n7267_), .ZN(new_n7343_));
  OAI21_X1   g07064(.A1(new_n7337_), .A2(new_n7338_), .B(new_n7341_), .ZN(new_n7344_));
  NAND3_X1   g07065(.A1(new_n7270_), .A2(new_n7272_), .A3(new_n7335_), .ZN(new_n7345_));
  NAND3_X1   g07066(.A1(new_n7345_), .A2(new_n7344_), .A3(new_n7266_), .ZN(new_n7346_));
  OAI22_X1   g07067(.A1(new_n930_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1017_), .ZN(new_n7347_));
  OAI21_X1   g07068(.A1(new_n861_), .A2(new_n3569_), .B(new_n7347_), .ZN(new_n7348_));
  AOI21_X1   g07069(.A1(new_n7348_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n7349_));
  XOR2_X1    g07070(.A1(new_n1024_), .A2(new_n7349_), .Z(new_n7350_));
  AOI21_X1   g07071(.A1(new_n7343_), .A2(new_n7346_), .B(new_n7350_), .ZN(new_n7351_));
  NAND2_X1   g07072(.A1(new_n7351_), .A2(new_n7265_), .ZN(new_n7352_));
  AOI21_X1   g07073(.A1(new_n7017_), .A2(new_n6717_), .B(new_n7009_), .ZN(new_n7353_));
  INV_X1     g07074(.I(new_n7264_), .ZN(new_n7354_));
  NOR3_X1    g07075(.A1(new_n7353_), .A2(new_n6604_), .A3(new_n7354_), .ZN(new_n7355_));
  AOI21_X1   g07076(.A1(new_n7345_), .A2(new_n7344_), .B(new_n7266_), .ZN(new_n7356_));
  NOR3_X1    g07077(.A1(new_n7336_), .A2(new_n7342_), .A3(new_n7267_), .ZN(new_n7357_));
  INV_X1     g07078(.I(new_n7350_), .ZN(new_n7358_));
  OAI21_X1   g07079(.A1(new_n7356_), .A2(new_n7357_), .B(new_n7358_), .ZN(new_n7359_));
  NAND2_X1   g07080(.A1(new_n7359_), .A2(new_n7355_), .ZN(new_n7360_));
  AOI21_X1   g07081(.A1(new_n7360_), .A2(new_n7352_), .B(new_n7262_), .ZN(new_n7361_));
  INV_X1     g07082(.I(new_n7262_), .ZN(new_n7362_));
  NOR2_X1    g07083(.A1(new_n7359_), .A2(new_n7355_), .ZN(new_n7363_));
  NOR2_X1    g07084(.A1(new_n7351_), .A2(new_n7265_), .ZN(new_n7364_));
  NOR3_X1    g07085(.A1(new_n7363_), .A2(new_n7364_), .A3(new_n7362_), .ZN(new_n7365_));
  OAI22_X1   g07086(.A1(new_n1189_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1294_), .ZN(new_n7366_));
  OAI21_X1   g07087(.A1(new_n1109_), .A2(new_n2884_), .B(new_n7366_), .ZN(new_n7367_));
  AOI21_X1   g07088(.A1(new_n7367_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n7368_));
  XOR2_X1    g07089(.A1(new_n1299_), .A2(new_n7368_), .Z(new_n7369_));
  INV_X1     g07090(.I(new_n7369_), .ZN(new_n7370_));
  OAI21_X1   g07091(.A1(new_n7361_), .A2(new_n7365_), .B(new_n7370_), .ZN(new_n7371_));
  NOR2_X1    g07092(.A1(new_n7259_), .A2(new_n7371_), .ZN(new_n7372_));
  AOI21_X1   g07093(.A1(new_n7035_), .A2(new_n7036_), .B(new_n7034_), .ZN(new_n7373_));
  OAI21_X1   g07094(.A1(new_n7373_), .A2(new_n6745_), .B(new_n6599_), .ZN(new_n7374_));
  OAI21_X1   g07095(.A1(new_n7363_), .A2(new_n7364_), .B(new_n7362_), .ZN(new_n7375_));
  NAND3_X1   g07096(.A1(new_n7360_), .A2(new_n7352_), .A3(new_n7262_), .ZN(new_n7376_));
  AOI21_X1   g07097(.A1(new_n7375_), .A2(new_n7376_), .B(new_n7369_), .ZN(new_n7377_));
  NOR2_X1    g07098(.A1(new_n7374_), .A2(new_n7377_), .ZN(new_n7378_));
  OAI21_X1   g07099(.A1(new_n7372_), .A2(new_n7378_), .B(new_n7257_), .ZN(new_n7379_));
  NAND2_X1   g07100(.A1(new_n7374_), .A2(new_n7377_), .ZN(new_n7380_));
  NAND2_X1   g07101(.A1(new_n7259_), .A2(new_n7371_), .ZN(new_n7381_));
  NAND3_X1   g07102(.A1(new_n7381_), .A2(new_n7380_), .A3(new_n7256_), .ZN(new_n7382_));
  NAND2_X1   g07103(.A1(new_n7379_), .A2(new_n7382_), .ZN(new_n7383_));
  OAI22_X1   g07104(.A1(new_n2171_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n2166_), .ZN(new_n7384_));
  OAI21_X1   g07105(.A1(new_n1518_), .A2(new_n2322_), .B(new_n7384_), .ZN(new_n7385_));
  AOI21_X1   g07106(.A1(new_n7385_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n7386_));
  XNOR2_X1   g07107(.A1(new_n1638_), .A2(new_n7386_), .ZN(new_n7387_));
  INV_X1     g07108(.I(new_n7387_), .ZN(new_n7388_));
  NAND3_X1   g07109(.A1(new_n7255_), .A2(new_n7383_), .A3(new_n7388_), .ZN(new_n7389_));
  OAI21_X1   g07110(.A1(new_n7043_), .A2(new_n7047_), .B(new_n6900_), .ZN(new_n7390_));
  AOI21_X1   g07111(.A1(new_n7390_), .A2(new_n6896_), .B(new_n7053_), .ZN(new_n7391_));
  NAND2_X1   g07112(.A1(new_n7383_), .A2(new_n7388_), .ZN(new_n7392_));
  NAND2_X1   g07113(.A1(new_n7392_), .A2(new_n7391_), .ZN(new_n7393_));
  AOI21_X1   g07114(.A1(new_n7393_), .A2(new_n7389_), .B(new_n7047_), .ZN(new_n7394_));
  NAND3_X1   g07115(.A1(new_n7393_), .A2(new_n7047_), .A3(new_n7389_), .ZN(new_n7395_));
  INV_X1     g07116(.I(new_n7395_), .ZN(new_n7396_));
  OAI22_X1   g07117(.A1(new_n1712_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n1707_), .ZN(new_n7397_));
  OAI21_X1   g07118(.A1(new_n1803_), .A2(new_n1850_), .B(new_n7397_), .ZN(new_n7398_));
  AOI21_X1   g07119(.A1(new_n7398_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n7399_));
  XOR2_X1    g07120(.A1(new_n2106_), .A2(new_n7399_), .Z(new_n7400_));
  INV_X1     g07121(.I(new_n7400_), .ZN(new_n7401_));
  OAI21_X1   g07122(.A1(new_n7396_), .A2(new_n7394_), .B(new_n7401_), .ZN(new_n7402_));
  NOR2_X1    g07123(.A1(new_n7253_), .A2(new_n7402_), .ZN(new_n7403_));
  NAND2_X1   g07124(.A1(new_n7085_), .A2(new_n6895_), .ZN(new_n7404_));
  NAND2_X1   g07125(.A1(new_n7060_), .A2(new_n6894_), .ZN(new_n7405_));
  AOI21_X1   g07126(.A1(new_n7405_), .A2(new_n7404_), .B(new_n7063_), .ZN(new_n7406_));
  OAI21_X1   g07127(.A1(new_n7406_), .A2(new_n7078_), .B(new_n6589_), .ZN(new_n7407_));
  INV_X1     g07128(.I(new_n7389_), .ZN(new_n7408_));
  AOI21_X1   g07129(.A1(new_n7383_), .A2(new_n7388_), .B(new_n7255_), .ZN(new_n7409_));
  OAI21_X1   g07130(.A1(new_n7408_), .A2(new_n7409_), .B(new_n7057_), .ZN(new_n7410_));
  NAND2_X1   g07131(.A1(new_n7410_), .A2(new_n7395_), .ZN(new_n7411_));
  AOI21_X1   g07132(.A1(new_n7411_), .A2(new_n7401_), .B(new_n7407_), .ZN(new_n7412_));
  OAI21_X1   g07133(.A1(new_n7412_), .A2(new_n7403_), .B(new_n7249_), .ZN(new_n7413_));
  NAND3_X1   g07134(.A1(new_n7407_), .A2(new_n7411_), .A3(new_n7401_), .ZN(new_n7414_));
  NAND2_X1   g07135(.A1(new_n7253_), .A2(new_n7402_), .ZN(new_n7415_));
  NAND3_X1   g07136(.A1(new_n7415_), .A2(new_n7414_), .A3(new_n7248_), .ZN(new_n7416_));
  OAI22_X1   g07137(.A1(new_n1347_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n1344_), .ZN(new_n7417_));
  OAI21_X1   g07138(.A1(new_n2281_), .A2(new_n1457_), .B(new_n7417_), .ZN(new_n7418_));
  AOI21_X1   g07139(.A1(new_n7418_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n7419_));
  XNOR2_X1   g07140(.A1(new_n2647_), .A2(new_n7419_), .ZN(new_n7420_));
  AOI21_X1   g07141(.A1(new_n7413_), .A2(new_n7416_), .B(new_n7420_), .ZN(new_n7421_));
  NAND2_X1   g07142(.A1(new_n7247_), .A2(new_n7421_), .ZN(new_n7422_));
  OAI21_X1   g07143(.A1(new_n7092_), .A2(new_n7089_), .B(new_n6890_), .ZN(new_n7423_));
  AOI21_X1   g07144(.A1(new_n7423_), .A2(new_n6782_), .B(new_n6584_), .ZN(new_n7424_));
  NAND2_X1   g07145(.A1(new_n7413_), .A2(new_n7416_), .ZN(new_n7425_));
  INV_X1     g07146(.I(new_n7420_), .ZN(new_n7426_));
  NAND2_X1   g07147(.A1(new_n7425_), .A2(new_n7426_), .ZN(new_n7427_));
  NAND2_X1   g07148(.A1(new_n7424_), .A2(new_n7427_), .ZN(new_n7428_));
  AOI21_X1   g07149(.A1(new_n7428_), .A2(new_n7422_), .B(new_n7245_), .ZN(new_n7429_));
  AOI21_X1   g07150(.A1(new_n7243_), .A2(new_n7242_), .B(new_n6895_), .ZN(new_n7430_));
  NOR3_X1    g07151(.A1(new_n7238_), .A2(new_n7240_), .A3(new_n6894_), .ZN(new_n7431_));
  OAI21_X1   g07152(.A1(new_n7430_), .A2(new_n7431_), .B(new_n7080_), .ZN(new_n7432_));
  NOR2_X1    g07153(.A1(new_n7424_), .A2(new_n7427_), .ZN(new_n7433_));
  NOR2_X1    g07154(.A1(new_n7247_), .A2(new_n7421_), .ZN(new_n7434_));
  NOR3_X1    g07155(.A1(new_n7433_), .A2(new_n7434_), .A3(new_n7432_), .ZN(new_n7435_));
  OAI22_X1   g07156(.A1(new_n1055_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n1061_), .ZN(new_n7436_));
  OAI21_X1   g07157(.A1(new_n2842_), .A2(new_n1332_), .B(new_n7436_), .ZN(new_n7437_));
  AOI21_X1   g07158(.A1(new_n7437_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n7438_));
  XNOR2_X1   g07159(.A1(new_n3264_), .A2(new_n7438_), .ZN(new_n7439_));
  INV_X1     g07160(.I(new_n7439_), .ZN(new_n7440_));
  OAI21_X1   g07161(.A1(new_n7429_), .A2(new_n7435_), .B(new_n7440_), .ZN(new_n7441_));
  NOR2_X1    g07162(.A1(new_n7236_), .A2(new_n7441_), .ZN(new_n7442_));
  AOI21_X1   g07163(.A1(new_n7106_), .A2(new_n7109_), .B(new_n6888_), .ZN(new_n7443_));
  OAI21_X1   g07164(.A1(new_n7443_), .A2(new_n6788_), .B(new_n6579_), .ZN(new_n7444_));
  OAI21_X1   g07165(.A1(new_n7433_), .A2(new_n7434_), .B(new_n7432_), .ZN(new_n7445_));
  NAND3_X1   g07166(.A1(new_n7428_), .A2(new_n7422_), .A3(new_n7245_), .ZN(new_n7446_));
  AOI21_X1   g07167(.A1(new_n7445_), .A2(new_n7446_), .B(new_n7439_), .ZN(new_n7447_));
  NOR2_X1    g07168(.A1(new_n7444_), .A2(new_n7447_), .ZN(new_n7448_));
  OAI21_X1   g07169(.A1(new_n7448_), .A2(new_n7442_), .B(new_n7234_), .ZN(new_n7449_));
  NAND2_X1   g07170(.A1(new_n7444_), .A2(new_n7447_), .ZN(new_n7450_));
  NAND2_X1   g07171(.A1(new_n7236_), .A2(new_n7441_), .ZN(new_n7451_));
  NAND3_X1   g07172(.A1(new_n7450_), .A2(new_n7451_), .A3(new_n7233_), .ZN(new_n7452_));
  OAI22_X1   g07173(.A1(new_n970_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n820_), .ZN(new_n7453_));
  OAI21_X1   g07174(.A1(new_n3709_), .A2(new_n894_), .B(new_n7453_), .ZN(new_n7454_));
  AOI21_X1   g07175(.A1(new_n7454_), .A2(new_n827_), .B(new_n970_), .ZN(new_n7455_));
  XNOR2_X1   g07176(.A1(new_n3993_), .A2(new_n7455_), .ZN(new_n7456_));
  AOI21_X1   g07177(.A1(new_n7449_), .A2(new_n7452_), .B(new_n7456_), .ZN(new_n7457_));
  OAI21_X1   g07178(.A1(new_n7232_), .A2(new_n7231_), .B(new_n7457_), .ZN(new_n7458_));
  OAI21_X1   g07179(.A1(new_n7120_), .A2(new_n7124_), .B(new_n6800_), .ZN(new_n7459_));
  NAND2_X1   g07180(.A1(new_n7459_), .A2(new_n6883_), .ZN(new_n7460_));
  NOR3_X1    g07181(.A1(new_n7120_), .A2(new_n7124_), .A3(new_n6800_), .ZN(new_n7461_));
  NOR2_X1    g07182(.A1(new_n6576_), .A2(new_n7461_), .ZN(new_n7462_));
  AOI21_X1   g07183(.A1(new_n7450_), .A2(new_n7451_), .B(new_n7233_), .ZN(new_n7463_));
  NOR3_X1    g07184(.A1(new_n7448_), .A2(new_n7442_), .A3(new_n7234_), .ZN(new_n7464_));
  INV_X1     g07185(.I(new_n7456_), .ZN(new_n7465_));
  OAI21_X1   g07186(.A1(new_n7464_), .A2(new_n7463_), .B(new_n7465_), .ZN(new_n7466_));
  NAND3_X1   g07187(.A1(new_n7462_), .A2(new_n7466_), .A3(new_n7460_), .ZN(new_n7467_));
  AOI21_X1   g07188(.A1(new_n7467_), .A2(new_n7458_), .B(new_n7229_), .ZN(new_n7468_));
  NAND3_X1   g07189(.A1(new_n7467_), .A2(new_n7458_), .A3(new_n7229_), .ZN(new_n7469_));
  INV_X1     g07190(.I(new_n7469_), .ZN(new_n7470_));
  OAI22_X1   g07191(.A1(new_n607_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n610_), .ZN(new_n7471_));
  OAI21_X1   g07192(.A1(new_n4253_), .A2(new_n684_), .B(new_n7471_), .ZN(new_n7472_));
  AOI21_X1   g07193(.A1(new_n7472_), .A2(new_n612_), .B(new_n607_), .ZN(new_n7473_));
  XNOR2_X1   g07194(.A1(new_n4778_), .A2(new_n7473_), .ZN(new_n7474_));
  INV_X1     g07195(.I(new_n7474_), .ZN(new_n7475_));
  OAI21_X1   g07196(.A1(new_n7470_), .A2(new_n7468_), .B(new_n7475_), .ZN(new_n7476_));
  NOR2_X1    g07197(.A1(new_n7227_), .A2(new_n7476_), .ZN(new_n7477_));
  AOI21_X1   g07198(.A1(new_n7145_), .A2(new_n7142_), .B(new_n6882_), .ZN(new_n7478_));
  OAI21_X1   g07199(.A1(new_n7478_), .A2(new_n6832_), .B(new_n7150_), .ZN(new_n7479_));
  AOI21_X1   g07200(.A1(new_n7462_), .A2(new_n7460_), .B(new_n7466_), .ZN(new_n7480_));
  NOR3_X1    g07201(.A1(new_n7232_), .A2(new_n7457_), .A3(new_n7231_), .ZN(new_n7481_));
  OAI21_X1   g07202(.A1(new_n7480_), .A2(new_n7481_), .B(new_n7228_), .ZN(new_n7482_));
  AOI21_X1   g07203(.A1(new_n7482_), .A2(new_n7469_), .B(new_n7474_), .ZN(new_n7483_));
  NOR2_X1    g07204(.A1(new_n7479_), .A2(new_n7483_), .ZN(new_n7484_));
  OAI21_X1   g07205(.A1(new_n7477_), .A2(new_n7484_), .B(new_n7145_), .ZN(new_n7485_));
  NAND2_X1   g07206(.A1(new_n7479_), .A2(new_n7483_), .ZN(new_n7486_));
  NAND2_X1   g07207(.A1(new_n7227_), .A2(new_n7476_), .ZN(new_n7487_));
  NAND3_X1   g07208(.A1(new_n7487_), .A2(new_n7486_), .A3(new_n7154_), .ZN(new_n7488_));
  OAI22_X1   g07209(.A1(new_n448_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n450_), .ZN(new_n7489_));
  OAI21_X1   g07210(.A1(new_n5068_), .A2(new_n496_), .B(new_n7489_), .ZN(new_n7490_));
  AOI21_X1   g07211(.A1(new_n7490_), .A2(new_n452_), .B(new_n448_), .ZN(new_n7491_));
  XNOR2_X1   g07212(.A1(new_n5600_), .A2(new_n7491_), .ZN(new_n7492_));
  AOI21_X1   g07213(.A1(new_n7485_), .A2(new_n7488_), .B(new_n7492_), .ZN(new_n7493_));
  NAND2_X1   g07214(.A1(new_n7225_), .A2(new_n7493_), .ZN(new_n7494_));
  AOI21_X1   g07215(.A1(new_n7166_), .A2(new_n6816_), .B(new_n6838_), .ZN(new_n7495_));
  NAND3_X1   g07216(.A1(new_n7165_), .A2(new_n7162_), .A3(new_n6833_), .ZN(new_n7496_));
  NAND2_X1   g07217(.A1(new_n7496_), .A2(new_n6829_), .ZN(new_n7497_));
  NOR2_X1    g07218(.A1(new_n7497_), .A2(new_n7495_), .ZN(new_n7498_));
  INV_X1     g07219(.I(new_n7493_), .ZN(new_n7499_));
  NAND2_X1   g07220(.A1(new_n7498_), .A2(new_n7499_), .ZN(new_n7500_));
  AOI21_X1   g07221(.A1(new_n7494_), .A2(new_n7500_), .B(new_n7216_), .ZN(new_n7501_));
  NOR2_X1    g07222(.A1(new_n7498_), .A2(new_n7499_), .ZN(new_n7502_));
  NOR2_X1    g07223(.A1(new_n7225_), .A2(new_n7493_), .ZN(new_n7503_));
  NOR3_X1    g07224(.A1(new_n7503_), .A2(new_n7502_), .A3(new_n7165_), .ZN(new_n7504_));
  NOR2_X1    g07225(.A1(new_n7501_), .A2(new_n7504_), .ZN(new_n7505_));
  OAI22_X1   g07226(.A1(new_n6229_), .A2(new_n341_), .B1(new_n404_), .B2(new_n6538_), .ZN(new_n7506_));
  OAI21_X1   g07227(.A1(new_n5921_), .A2(new_n366_), .B(new_n7506_), .ZN(new_n7507_));
  AOI21_X1   g07228(.A1(new_n7507_), .A2(new_n334_), .B(new_n341_), .ZN(new_n7508_));
  XOR2_X1    g07229(.A1(new_n6543_), .A2(new_n7508_), .Z(new_n7509_));
  XOR2_X1    g07230(.A1(new_n7505_), .A2(new_n7509_), .Z(new_n7510_));
  INV_X1     g07231(.I(new_n7510_), .ZN(new_n7511_));
  XNOR2_X1   g07232(.A1(\b[43] ), .A2(\b[45] ), .ZN(new_n7512_));
  NOR4_X1    g07233(.A1(new_n7192_), .A2(new_n7195_), .A3(new_n7197_), .A4(new_n7512_), .ZN(new_n7513_));
  NOR2_X1    g07234(.A1(new_n7512_), .A2(new_n7197_), .ZN(new_n7514_));
  NOR2_X1    g07235(.A1(new_n7196_), .A2(new_n7514_), .ZN(new_n7515_));
  NOR2_X1    g07236(.A1(new_n7515_), .A2(new_n7513_), .ZN(new_n7516_));
  INV_X1     g07237(.I(new_n7516_), .ZN(new_n7517_));
  NAND2_X1   g07238(.A1(new_n286_), .A2(\b[44] ), .ZN(new_n7518_));
  AOI22_X1   g07239(.A1(new_n304_), .A2(\b[43] ), .B1(new_n262_), .B2(\b[45] ), .ZN(new_n7519_));
  AOI21_X1   g07240(.A1(new_n7518_), .A2(new_n7519_), .B(new_n426_), .ZN(new_n7520_));
  AND3_X2    g07241(.A1(new_n7511_), .A2(new_n7517_), .A3(new_n7520_), .Z(new_n7521_));
  AOI21_X1   g07242(.A1(new_n7517_), .A2(new_n7520_), .B(new_n7511_), .ZN(new_n7522_));
  OAI21_X1   g07243(.A1(new_n7521_), .A2(new_n7522_), .B(new_n7221_), .ZN(new_n7523_));
  NOR3_X1    g07244(.A1(new_n7521_), .A2(new_n7221_), .A3(new_n7522_), .ZN(new_n7524_));
  INV_X1     g07245(.I(new_n7524_), .ZN(new_n7525_));
  NAND2_X1   g07246(.A1(new_n7525_), .A2(new_n7523_), .ZN(new_n7526_));
  NAND2_X1   g07247(.A1(new_n7526_), .A2(new_n260_), .ZN(new_n7527_));
  NAND3_X1   g07248(.A1(new_n7525_), .A2(\a[2] ), .A3(new_n7523_), .ZN(new_n7528_));
  AOI21_X1   g07249(.A1(new_n7527_), .A2(new_n7528_), .B(new_n7207_), .ZN(new_n7529_));
  XOR2_X1    g07250(.A1(new_n7529_), .A2(new_n7212_), .Z(new_n7530_));
  XOR2_X1    g07251(.A1(new_n7530_), .A2(new_n6875_), .Z(\f[45] ));
  NOR3_X1    g07252(.A1(new_n7220_), .A2(new_n7178_), .A3(new_n7176_), .ZN(new_n7532_));
  OAI22_X1   g07253(.A1(new_n448_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n450_), .ZN(new_n7533_));
  OAI21_X1   g07254(.A1(new_n5353_), .A2(new_n496_), .B(new_n7533_), .ZN(new_n7534_));
  AOI21_X1   g07255(.A1(new_n7534_), .A2(new_n452_), .B(new_n448_), .ZN(new_n7535_));
  XOR2_X1    g07256(.A1(new_n5926_), .A2(new_n7535_), .Z(new_n7536_));
  NOR2_X1    g07257(.A1(new_n7470_), .A2(new_n7468_), .ZN(new_n7537_));
  NAND3_X1   g07258(.A1(new_n7482_), .A2(new_n7469_), .A3(new_n7145_), .ZN(new_n7538_));
  NAND2_X1   g07259(.A1(new_n7538_), .A2(new_n7475_), .ZN(new_n7539_));
  OAI22_X1   g07260(.A1(new_n7539_), .A2(new_n7479_), .B1(new_n7145_), .B2(new_n7537_), .ZN(new_n7540_));
  NOR2_X1    g07261(.A1(new_n7232_), .A2(new_n7231_), .ZN(new_n7541_));
  NAND2_X1   g07262(.A1(new_n7449_), .A2(new_n7452_), .ZN(new_n7542_));
  NAND3_X1   g07263(.A1(new_n7449_), .A2(new_n7452_), .A3(new_n7228_), .ZN(new_n7543_));
  AND2_X2    g07264(.A1(new_n7543_), .A2(new_n7465_), .Z(new_n7544_));
  AOI22_X1   g07265(.A1(new_n7544_), .A2(new_n7541_), .B1(new_n7542_), .B2(new_n7229_), .ZN(new_n7545_));
  OAI21_X1   g07266(.A1(new_n7429_), .A2(new_n7435_), .B(new_n7233_), .ZN(new_n7546_));
  NAND3_X1   g07267(.A1(new_n7445_), .A2(new_n7446_), .A3(new_n7234_), .ZN(new_n7547_));
  NAND2_X1   g07268(.A1(new_n7547_), .A2(new_n7440_), .ZN(new_n7548_));
  OAI21_X1   g07269(.A1(new_n7548_), .A2(new_n7444_), .B(new_n7546_), .ZN(new_n7549_));
  AOI21_X1   g07270(.A1(new_n7415_), .A2(new_n7414_), .B(new_n7248_), .ZN(new_n7550_));
  NOR3_X1    g07271(.A1(new_n7412_), .A2(new_n7403_), .A3(new_n7249_), .ZN(new_n7551_));
  NOR2_X1    g07272(.A1(new_n7551_), .A2(new_n7550_), .ZN(new_n7552_));
  OAI21_X1   g07273(.A1(new_n7425_), .A2(new_n7245_), .B(new_n7426_), .ZN(new_n7553_));
  OAI22_X1   g07274(.A1(new_n7553_), .A2(new_n7247_), .B1(new_n7432_), .B2(new_n7552_), .ZN(new_n7554_));
  INV_X1     g07275(.I(new_n7411_), .ZN(new_n7555_));
  NOR2_X1    g07276(.A1(new_n7555_), .A2(new_n7249_), .ZN(new_n7556_));
  OAI21_X1   g07277(.A1(new_n7411_), .A2(new_n7248_), .B(new_n7401_), .ZN(new_n7557_));
  NOR2_X1    g07278(.A1(new_n7557_), .A2(new_n7407_), .ZN(new_n7558_));
  NOR2_X1    g07279(.A1(new_n7558_), .A2(new_n7556_), .ZN(new_n7559_));
  AOI21_X1   g07280(.A1(new_n7379_), .A2(new_n7382_), .B(new_n7057_), .ZN(new_n7560_));
  INV_X1     g07281(.I(new_n7560_), .ZN(new_n7561_));
  NAND3_X1   g07282(.A1(new_n7379_), .A2(new_n7382_), .A3(new_n7057_), .ZN(new_n7562_));
  NAND3_X1   g07283(.A1(new_n7391_), .A2(new_n7562_), .A3(new_n7388_), .ZN(new_n7563_));
  NAND2_X1   g07284(.A1(new_n7563_), .A2(new_n7561_), .ZN(new_n7564_));
  OAI21_X1   g07285(.A1(new_n7361_), .A2(new_n7365_), .B(new_n7256_), .ZN(new_n7565_));
  NAND3_X1   g07286(.A1(new_n7375_), .A2(new_n7376_), .A3(new_n7257_), .ZN(new_n7566_));
  NAND2_X1   g07287(.A1(new_n7566_), .A2(new_n7370_), .ZN(new_n7567_));
  OAI21_X1   g07288(.A1(new_n7567_), .A2(new_n7374_), .B(new_n7565_), .ZN(new_n7568_));
  AOI21_X1   g07289(.A1(new_n7343_), .A2(new_n7346_), .B(new_n7362_), .ZN(new_n7569_));
  NAND3_X1   g07290(.A1(new_n7343_), .A2(new_n7346_), .A3(new_n7362_), .ZN(new_n7570_));
  NOR2_X1    g07291(.A1(new_n7265_), .A2(new_n7350_), .ZN(new_n7571_));
  AOI21_X1   g07292(.A1(new_n7571_), .A2(new_n7570_), .B(new_n7569_), .ZN(new_n7572_));
  NOR2_X1    g07293(.A1(new_n7337_), .A2(new_n7338_), .ZN(new_n7573_));
  AOI21_X1   g07294(.A1(new_n7339_), .A2(new_n7340_), .B(new_n7267_), .ZN(new_n7574_));
  NOR3_X1    g07295(.A1(new_n7326_), .A2(new_n7329_), .A3(new_n7266_), .ZN(new_n7575_));
  NOR2_X1    g07296(.A1(new_n7575_), .A2(new_n7333_), .ZN(new_n7576_));
  AOI21_X1   g07297(.A1(new_n7573_), .A2(new_n7576_), .B(new_n7574_), .ZN(new_n7577_));
  AOI21_X1   g07298(.A1(new_n7311_), .A2(new_n7314_), .B(new_n6965_), .ZN(new_n7578_));
  AOI21_X1   g07299(.A1(new_n7313_), .A2(new_n7308_), .B(new_n7312_), .ZN(new_n7579_));
  NOR3_X1    g07300(.A1(new_n7309_), .A2(new_n7279_), .A3(new_n7310_), .ZN(new_n7580_));
  NOR3_X1    g07301(.A1(new_n7580_), .A2(new_n7579_), .A3(new_n6974_), .ZN(new_n7581_));
  NOR2_X1    g07302(.A1(new_n7581_), .A2(new_n7318_), .ZN(new_n7582_));
  AOI21_X1   g07303(.A1(new_n7323_), .A2(new_n7582_), .B(new_n7578_), .ZN(new_n7583_));
  NAND2_X1   g07304(.A1(new_n7302_), .A2(new_n7300_), .ZN(new_n7584_));
  NAND2_X1   g07305(.A1(new_n7584_), .A2(new_n7312_), .ZN(new_n7585_));
  INV_X1     g07306(.I(new_n7585_), .ZN(new_n7586_));
  INV_X1     g07307(.I(new_n7306_), .ZN(new_n7587_));
  OAI21_X1   g07308(.A1(new_n7584_), .A2(new_n7312_), .B(new_n7587_), .ZN(new_n7588_));
  NOR3_X1    g07309(.A1(new_n7588_), .A2(new_n7280_), .A3(new_n7281_), .ZN(new_n7589_));
  NOR2_X1    g07310(.A1(new_n7589_), .A2(new_n7586_), .ZN(new_n7590_));
  OAI21_X1   g07311(.A1(new_n7290_), .A2(new_n7291_), .B(new_n6938_), .ZN(new_n7591_));
  NAND3_X1   g07312(.A1(new_n6921_), .A2(new_n7289_), .A3(new_n7296_), .ZN(new_n7592_));
  NOR2_X1    g07313(.A1(new_n6929_), .A2(new_n7297_), .ZN(new_n7593_));
  NAND2_X1   g07314(.A1(new_n7592_), .A2(new_n7593_), .ZN(new_n7594_));
  NAND2_X1   g07315(.A1(new_n7594_), .A2(new_n7591_), .ZN(new_n7595_));
  AOI22_X1   g07316(.A1(new_n6631_), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n6637_), .ZN(new_n7596_));
  NOR2_X1    g07317(.A1(new_n7284_), .A2(new_n280_), .ZN(new_n7597_));
  OAI21_X1   g07318(.A1(new_n7596_), .A2(new_n7597_), .B(new_n6632_), .ZN(new_n7598_));
  NAND3_X1   g07319(.A1(new_n7598_), .A2(new_n807_), .A3(new_n6631_), .ZN(new_n7599_));
  OAI22_X1   g07320(.A1(new_n6644_), .A2(new_n298_), .B1(new_n325_), .B2(new_n6647_), .ZN(new_n7600_));
  NAND2_X1   g07321(.A1(new_n6914_), .A2(\b[2] ), .ZN(new_n7601_));
  AOI21_X1   g07322(.A1(new_n7600_), .A2(new_n7601_), .B(\a[44] ), .ZN(new_n7602_));
  OAI21_X1   g07323(.A1(new_n7602_), .A2(new_n6644_), .B(new_n329_), .ZN(new_n7603_));
  NAND2_X1   g07324(.A1(new_n7603_), .A2(new_n7599_), .ZN(new_n7604_));
  XNOR2_X1   g07325(.A1(\a[45] ), .A2(\a[47] ), .ZN(new_n7605_));
  XNOR2_X1   g07326(.A1(\a[44] ), .A2(\a[46] ), .ZN(new_n7606_));
  NOR2_X1    g07327(.A1(new_n7605_), .A2(new_n7606_), .ZN(new_n7607_));
  INV_X1     g07328(.I(\a[47] ), .ZN(new_n7608_));
  INV_X1     g07329(.I(\a[46] ), .ZN(new_n7609_));
  NOR3_X1    g07330(.A1(new_n7609_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n7610_));
  INV_X1     g07331(.I(\a[45] ), .ZN(new_n7611_));
  NOR3_X1    g07332(.A1(new_n6632_), .A2(new_n7611_), .A3(\a[46] ), .ZN(new_n7612_));
  OAI21_X1   g07333(.A1(new_n7612_), .A2(new_n7610_), .B(\b[1] ), .ZN(new_n7613_));
  XOR2_X1    g07334(.A1(\a[45] ), .A2(\a[47] ), .Z(new_n7614_));
  XOR2_X1    g07335(.A1(\a[44] ), .A2(\a[46] ), .Z(new_n7615_));
  NAND3_X1   g07336(.A1(new_n7614_), .A2(new_n7615_), .A3(\b[0] ), .ZN(new_n7616_));
  NAND3_X1   g07337(.A1(new_n7616_), .A2(new_n7608_), .A3(new_n7613_), .ZN(new_n7617_));
  NAND3_X1   g07338(.A1(new_n7617_), .A2(new_n444_), .A3(new_n7607_), .ZN(new_n7618_));
  NAND2_X1   g07339(.A1(new_n7614_), .A2(new_n7615_), .ZN(new_n7619_));
  NAND3_X1   g07340(.A1(new_n6632_), .A2(new_n7611_), .A3(\a[46] ), .ZN(new_n7620_));
  NAND3_X1   g07341(.A1(new_n7609_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n7621_));
  AOI21_X1   g07342(.A1(new_n7620_), .A2(new_n7621_), .B(new_n269_), .ZN(new_n7622_));
  NOR3_X1    g07343(.A1(new_n7605_), .A2(new_n7606_), .A3(new_n258_), .ZN(new_n7623_));
  NOR3_X1    g07344(.A1(new_n7623_), .A2(\a[47] ), .A3(new_n7622_), .ZN(new_n7624_));
  OAI21_X1   g07345(.A1(new_n7624_), .A2(new_n7619_), .B(new_n271_), .ZN(new_n7625_));
  NOR2_X1    g07346(.A1(new_n7293_), .A2(new_n7608_), .ZN(new_n7626_));
  INV_X1     g07347(.I(new_n7626_), .ZN(new_n7627_));
  NAND3_X1   g07348(.A1(new_n7625_), .A2(new_n7618_), .A3(new_n7627_), .ZN(new_n7628_));
  NOR3_X1    g07349(.A1(new_n7624_), .A2(new_n271_), .A3(new_n7619_), .ZN(new_n7629_));
  AOI21_X1   g07350(.A1(new_n7617_), .A2(new_n7607_), .B(new_n444_), .ZN(new_n7630_));
  OAI21_X1   g07351(.A1(new_n7629_), .A2(new_n7630_), .B(new_n7626_), .ZN(new_n7631_));
  NAND2_X1   g07352(.A1(new_n7631_), .A2(new_n7628_), .ZN(new_n7632_));
  NAND2_X1   g07353(.A1(new_n7604_), .A2(new_n7632_), .ZN(new_n7633_));
  NOR3_X1    g07354(.A1(new_n7602_), .A2(new_n329_), .A3(new_n6644_), .ZN(new_n7634_));
  AOI21_X1   g07355(.A1(new_n7598_), .A2(new_n6631_), .B(new_n807_), .ZN(new_n7635_));
  NOR2_X1    g07356(.A1(new_n7634_), .A2(new_n7635_), .ZN(new_n7636_));
  INV_X1     g07357(.I(new_n7632_), .ZN(new_n7637_));
  NAND2_X1   g07358(.A1(new_n7637_), .A2(new_n7636_), .ZN(new_n7638_));
  NAND2_X1   g07359(.A1(new_n7638_), .A2(new_n7633_), .ZN(new_n7639_));
  NAND2_X1   g07360(.A1(new_n7595_), .A2(new_n7639_), .ZN(new_n7640_));
  AOI21_X1   g07361(.A1(new_n7289_), .A2(new_n7296_), .B(new_n6921_), .ZN(new_n7641_));
  AOI21_X1   g07362(.A1(new_n7592_), .A2(new_n7593_), .B(new_n7641_), .ZN(new_n7642_));
  NAND2_X1   g07363(.A1(new_n7636_), .A2(new_n7632_), .ZN(new_n7643_));
  NAND3_X1   g07364(.A1(new_n7604_), .A2(new_n7628_), .A3(new_n7631_), .ZN(new_n7644_));
  NAND2_X1   g07365(.A1(new_n7644_), .A2(new_n7643_), .ZN(new_n7645_));
  NAND2_X1   g07366(.A1(new_n7642_), .A2(new_n7645_), .ZN(new_n7646_));
  NAND2_X1   g07367(.A1(new_n7640_), .A2(new_n7646_), .ZN(new_n7647_));
  AOI22_X1   g07368(.A1(new_n5680_), .A2(\b[6] ), .B1(\b[7] ), .B2(new_n5686_), .ZN(new_n7648_));
  NOR2_X1    g07369(.A1(new_n5997_), .A2(new_n419_), .ZN(new_n7649_));
  OAI21_X1   g07370(.A1(new_n7648_), .A2(new_n7649_), .B(new_n5681_), .ZN(new_n7650_));
  NAND2_X1   g07371(.A1(new_n7650_), .A2(new_n5680_), .ZN(new_n7651_));
  XNOR2_X1   g07372(.A1(new_n471_), .A2(new_n7651_), .ZN(new_n7652_));
  INV_X1     g07373(.I(new_n7652_), .ZN(new_n7653_));
  NAND2_X1   g07374(.A1(new_n7647_), .A2(new_n7653_), .ZN(new_n7654_));
  INV_X1     g07375(.I(new_n7654_), .ZN(new_n7655_));
  NOR2_X1    g07376(.A1(new_n7647_), .A2(new_n7653_), .ZN(new_n7656_));
  NOR2_X1    g07377(.A1(new_n7655_), .A2(new_n7656_), .ZN(new_n7657_));
  NOR2_X1    g07378(.A1(new_n7590_), .A2(new_n7657_), .ZN(new_n7658_));
  NOR2_X1    g07379(.A1(new_n7280_), .A2(new_n7281_), .ZN(new_n7659_));
  INV_X1     g07380(.I(new_n7659_), .ZN(new_n7660_));
  OAI21_X1   g07381(.A1(new_n7660_), .A2(new_n7588_), .B(new_n7585_), .ZN(new_n7661_));
  NAND3_X1   g07382(.A1(new_n7640_), .A2(new_n7646_), .A3(new_n7653_), .ZN(new_n7662_));
  NAND2_X1   g07383(.A1(new_n7647_), .A2(new_n7652_), .ZN(new_n7663_));
  NAND2_X1   g07384(.A1(new_n7663_), .A2(new_n7662_), .ZN(new_n7664_));
  INV_X1     g07385(.I(new_n7664_), .ZN(new_n7665_));
  NOR2_X1    g07386(.A1(new_n7661_), .A2(new_n7665_), .ZN(new_n7666_));
  NOR2_X1    g07387(.A1(new_n7666_), .A2(new_n7658_), .ZN(new_n7667_));
  OAI22_X1   g07388(.A1(new_n5420_), .A2(new_n565_), .B1(new_n656_), .B2(new_n5107_), .ZN(new_n7668_));
  OAI21_X1   g07389(.A1(new_n515_), .A2(new_n5112_), .B(new_n7668_), .ZN(new_n7669_));
  AOI21_X1   g07390(.A1(new_n7669_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n7670_));
  XNOR2_X1   g07391(.A1(new_n660_), .A2(new_n7670_), .ZN(new_n7671_));
  INV_X1     g07392(.I(new_n7671_), .ZN(new_n7672_));
  NAND2_X1   g07393(.A1(new_n7667_), .A2(new_n7672_), .ZN(new_n7673_));
  NOR2_X1    g07394(.A1(new_n7667_), .A2(new_n7672_), .ZN(new_n7674_));
  INV_X1     g07395(.I(new_n7674_), .ZN(new_n7675_));
  AOI21_X1   g07396(.A1(new_n7673_), .A2(new_n7675_), .B(new_n7583_), .ZN(new_n7676_));
  INV_X1     g07397(.I(new_n7578_), .ZN(new_n7677_));
  INV_X1     g07398(.I(new_n7318_), .ZN(new_n7678_));
  NAND3_X1   g07399(.A1(new_n7311_), .A2(new_n7314_), .A3(new_n6965_), .ZN(new_n7679_));
  NAND2_X1   g07400(.A1(new_n7679_), .A2(new_n7678_), .ZN(new_n7680_));
  OAI21_X1   g07401(.A1(new_n7276_), .A2(new_n7680_), .B(new_n7677_), .ZN(new_n7681_));
  NOR2_X1    g07402(.A1(new_n7667_), .A2(new_n7671_), .ZN(new_n7682_));
  NOR3_X1    g07403(.A1(new_n7666_), .A2(new_n7658_), .A3(new_n7672_), .ZN(new_n7683_));
  NOR2_X1    g07404(.A1(new_n7682_), .A2(new_n7683_), .ZN(new_n7684_));
  NOR2_X1    g07405(.A1(new_n7684_), .A2(new_n7681_), .ZN(new_n7685_));
  OAI22_X1   g07406(.A1(new_n4072_), .A2(new_n780_), .B1(new_n861_), .B2(new_n4067_), .ZN(new_n7686_));
  OAI21_X1   g07407(.A1(new_n706_), .A2(new_n4318_), .B(new_n7686_), .ZN(new_n7687_));
  AOI21_X1   g07408(.A1(new_n7687_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n7688_));
  XNOR2_X1   g07409(.A1(new_n860_), .A2(new_n7688_), .ZN(new_n7689_));
  NOR3_X1    g07410(.A1(new_n7676_), .A2(new_n7685_), .A3(new_n7689_), .ZN(new_n7690_));
  OR2_X2     g07411(.A1(new_n7666_), .A2(new_n7658_), .Z(new_n7691_));
  NOR2_X1    g07412(.A1(new_n7691_), .A2(new_n7671_), .ZN(new_n7692_));
  OAI21_X1   g07413(.A1(new_n7692_), .A2(new_n7674_), .B(new_n7681_), .ZN(new_n7693_));
  OAI21_X1   g07414(.A1(new_n7682_), .A2(new_n7683_), .B(new_n7583_), .ZN(new_n7694_));
  INV_X1     g07415(.I(new_n7689_), .ZN(new_n7695_));
  AOI21_X1   g07416(.A1(new_n7694_), .A2(new_n7693_), .B(new_n7695_), .ZN(new_n7696_));
  NOR2_X1    g07417(.A1(new_n7696_), .A2(new_n7690_), .ZN(new_n7697_));
  OAI22_X1   g07418(.A1(new_n1017_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1109_), .ZN(new_n7698_));
  OAI21_X1   g07419(.A1(new_n930_), .A2(new_n3569_), .B(new_n7698_), .ZN(new_n7699_));
  AOI21_X1   g07420(.A1(new_n7699_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n7700_));
  XOR2_X1    g07421(.A1(new_n1114_), .A2(new_n7700_), .Z(new_n7701_));
  INV_X1     g07422(.I(new_n7701_), .ZN(new_n7702_));
  NAND2_X1   g07423(.A1(new_n7697_), .A2(new_n7702_), .ZN(new_n7703_));
  NAND3_X1   g07424(.A1(new_n7694_), .A2(new_n7693_), .A3(new_n7695_), .ZN(new_n7704_));
  OAI21_X1   g07425(.A1(new_n7676_), .A2(new_n7685_), .B(new_n7689_), .ZN(new_n7705_));
  NAND2_X1   g07426(.A1(new_n7704_), .A2(new_n7705_), .ZN(new_n7706_));
  NAND2_X1   g07427(.A1(new_n7706_), .A2(new_n7701_), .ZN(new_n7707_));
  AOI21_X1   g07428(.A1(new_n7703_), .A2(new_n7707_), .B(new_n7577_), .ZN(new_n7708_));
  NAND2_X1   g07429(.A1(new_n7272_), .A2(new_n7270_), .ZN(new_n7709_));
  INV_X1     g07430(.I(new_n7574_), .ZN(new_n7710_));
  NAND2_X1   g07431(.A1(new_n7339_), .A2(new_n7340_), .ZN(new_n7711_));
  OAI21_X1   g07432(.A1(new_n7711_), .A2(new_n7266_), .B(new_n7334_), .ZN(new_n7712_));
  OAI21_X1   g07433(.A1(new_n7709_), .A2(new_n7712_), .B(new_n7710_), .ZN(new_n7713_));
  NAND2_X1   g07434(.A1(new_n7706_), .A2(new_n7702_), .ZN(new_n7714_));
  NAND2_X1   g07435(.A1(new_n7697_), .A2(new_n7701_), .ZN(new_n7715_));
  AOI21_X1   g07436(.A1(new_n7714_), .A2(new_n7715_), .B(new_n7713_), .ZN(new_n7716_));
  OAI22_X1   g07437(.A1(new_n1294_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1518_), .ZN(new_n7717_));
  OAI21_X1   g07438(.A1(new_n1189_), .A2(new_n2884_), .B(new_n7717_), .ZN(new_n7718_));
  AOI21_X1   g07439(.A1(new_n7718_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n7719_));
  XNOR2_X1   g07440(.A1(new_n1421_), .A2(new_n7719_), .ZN(new_n7720_));
  INV_X1     g07441(.I(new_n7720_), .ZN(new_n7721_));
  OAI21_X1   g07442(.A1(new_n7716_), .A2(new_n7708_), .B(new_n7721_), .ZN(new_n7722_));
  NOR2_X1    g07443(.A1(new_n7716_), .A2(new_n7708_), .ZN(new_n7723_));
  NAND2_X1   g07444(.A1(new_n7723_), .A2(new_n7720_), .ZN(new_n7724_));
  AOI21_X1   g07445(.A1(new_n7722_), .A2(new_n7724_), .B(new_n7572_), .ZN(new_n7725_));
  INV_X1     g07446(.I(new_n7569_), .ZN(new_n7726_));
  NAND3_X1   g07447(.A1(new_n7570_), .A2(new_n7355_), .A3(new_n7358_), .ZN(new_n7727_));
  NAND2_X1   g07448(.A1(new_n7727_), .A2(new_n7726_), .ZN(new_n7728_));
  NAND2_X1   g07449(.A1(new_n7723_), .A2(new_n7721_), .ZN(new_n7729_));
  NOR2_X1    g07450(.A1(new_n7723_), .A2(new_n7721_), .ZN(new_n7730_));
  INV_X1     g07451(.I(new_n7730_), .ZN(new_n7731_));
  AOI21_X1   g07452(.A1(new_n7731_), .A2(new_n7729_), .B(new_n7728_), .ZN(new_n7732_));
  OAI22_X1   g07453(.A1(new_n2171_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n2166_), .ZN(new_n7733_));
  OAI21_X1   g07454(.A1(new_n1525_), .A2(new_n2322_), .B(new_n7733_), .ZN(new_n7734_));
  AOI21_X1   g07455(.A1(new_n7734_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n7735_));
  XOR2_X1    g07456(.A1(new_n1808_), .A2(new_n7735_), .Z(new_n7736_));
  INV_X1     g07457(.I(new_n7736_), .ZN(new_n7737_));
  OAI21_X1   g07458(.A1(new_n7732_), .A2(new_n7725_), .B(new_n7737_), .ZN(new_n7738_));
  NAND2_X1   g07459(.A1(new_n7724_), .A2(new_n7722_), .ZN(new_n7739_));
  NAND2_X1   g07460(.A1(new_n7739_), .A2(new_n7728_), .ZN(new_n7740_));
  OR2_X2     g07461(.A1(new_n7716_), .A2(new_n7708_), .Z(new_n7741_));
  NOR2_X1    g07462(.A1(new_n7741_), .A2(new_n7720_), .ZN(new_n7742_));
  OAI21_X1   g07463(.A1(new_n7742_), .A2(new_n7730_), .B(new_n7572_), .ZN(new_n7743_));
  NAND3_X1   g07464(.A1(new_n7740_), .A2(new_n7743_), .A3(new_n7736_), .ZN(new_n7744_));
  NAND2_X1   g07465(.A1(new_n7738_), .A2(new_n7744_), .ZN(new_n7745_));
  NAND2_X1   g07466(.A1(new_n7745_), .A2(new_n7568_), .ZN(new_n7746_));
  AOI21_X1   g07467(.A1(new_n7375_), .A2(new_n7376_), .B(new_n7257_), .ZN(new_n7747_));
  NOR3_X1    g07468(.A1(new_n7361_), .A2(new_n7365_), .A3(new_n7256_), .ZN(new_n7748_));
  NOR2_X1    g07469(.A1(new_n7748_), .A2(new_n7369_), .ZN(new_n7749_));
  AOI21_X1   g07470(.A1(new_n7749_), .A2(new_n7259_), .B(new_n7747_), .ZN(new_n7750_));
  NAND2_X1   g07471(.A1(new_n7740_), .A2(new_n7743_), .ZN(new_n7751_));
  NOR2_X1    g07472(.A1(new_n7751_), .A2(new_n7736_), .ZN(new_n7752_));
  NOR2_X1    g07473(.A1(new_n7732_), .A2(new_n7725_), .ZN(new_n7753_));
  NOR2_X1    g07474(.A1(new_n7753_), .A2(new_n7737_), .ZN(new_n7754_));
  OAI21_X1   g07475(.A1(new_n7752_), .A2(new_n7754_), .B(new_n7750_), .ZN(new_n7755_));
  NAND2_X1   g07476(.A1(new_n7755_), .A2(new_n7746_), .ZN(new_n7756_));
  OAI22_X1   g07477(.A1(new_n1712_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n1707_), .ZN(new_n7757_));
  OAI21_X1   g07478(.A1(new_n1936_), .A2(new_n1850_), .B(new_n7757_), .ZN(new_n7758_));
  AOI21_X1   g07479(.A1(new_n7758_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n7759_));
  XNOR2_X1   g07480(.A1(new_n2280_), .A2(new_n7759_), .ZN(new_n7760_));
  XOR2_X1    g07481(.A1(new_n7756_), .A2(new_n7760_), .Z(new_n7761_));
  NAND2_X1   g07482(.A1(new_n7761_), .A2(new_n7564_), .ZN(new_n7762_));
  AOI21_X1   g07483(.A1(new_n7381_), .A2(new_n7380_), .B(new_n7256_), .ZN(new_n7763_));
  NOR3_X1    g07484(.A1(new_n7372_), .A2(new_n7378_), .A3(new_n7257_), .ZN(new_n7764_));
  NOR3_X1    g07485(.A1(new_n7763_), .A2(new_n7764_), .A3(new_n7047_), .ZN(new_n7765_));
  NOR3_X1    g07486(.A1(new_n7765_), .A2(new_n7255_), .A3(new_n7387_), .ZN(new_n7766_));
  NOR2_X1    g07487(.A1(new_n7766_), .A2(new_n7560_), .ZN(new_n7767_));
  INV_X1     g07488(.I(new_n7760_), .ZN(new_n7768_));
  XOR2_X1    g07489(.A1(new_n7756_), .A2(new_n7768_), .Z(new_n7769_));
  NAND2_X1   g07490(.A1(new_n7769_), .A2(new_n7767_), .ZN(new_n7770_));
  NAND2_X1   g07491(.A1(new_n7762_), .A2(new_n7770_), .ZN(new_n7771_));
  OAI22_X1   g07492(.A1(new_n1347_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n1344_), .ZN(new_n7772_));
  OAI21_X1   g07493(.A1(new_n2439_), .A2(new_n1457_), .B(new_n7772_), .ZN(new_n7773_));
  AOI21_X1   g07494(.A1(new_n7773_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n7774_));
  XNOR2_X1   g07495(.A1(new_n2846_), .A2(new_n7774_), .ZN(new_n7775_));
  INV_X1     g07496(.I(new_n7775_), .ZN(new_n7776_));
  XOR2_X1    g07497(.A1(new_n7771_), .A2(new_n7776_), .Z(new_n7777_));
  XOR2_X1    g07498(.A1(new_n7771_), .A2(new_n7776_), .Z(new_n7778_));
  NAND2_X1   g07499(.A1(new_n7778_), .A2(new_n7559_), .ZN(new_n7779_));
  OAI21_X1   g07500(.A1(new_n7559_), .A2(new_n7777_), .B(new_n7779_), .ZN(new_n7780_));
  NAND2_X1   g07501(.A1(new_n7554_), .A2(new_n7780_), .ZN(new_n7781_));
  AOI21_X1   g07502(.A1(new_n7552_), .A2(new_n7432_), .B(new_n7420_), .ZN(new_n7782_));
  AOI22_X1   g07503(.A1(new_n7782_), .A2(new_n7424_), .B1(new_n7245_), .B2(new_n7425_), .ZN(new_n7783_));
  NOR2_X1    g07504(.A1(new_n7777_), .A2(new_n7559_), .ZN(new_n7784_));
  AOI21_X1   g07505(.A1(new_n7559_), .A2(new_n7778_), .B(new_n7784_), .ZN(new_n7785_));
  NAND2_X1   g07506(.A1(new_n7783_), .A2(new_n7785_), .ZN(new_n7786_));
  OAI22_X1   g07507(.A1(new_n1055_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n1061_), .ZN(new_n7787_));
  OAI21_X1   g07508(.A1(new_n3018_), .A2(new_n1332_), .B(new_n7787_), .ZN(new_n7788_));
  AOI21_X1   g07509(.A1(new_n7788_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n7789_));
  XNOR2_X1   g07510(.A1(new_n3514_), .A2(new_n7789_), .ZN(new_n7790_));
  INV_X1     g07511(.I(new_n7790_), .ZN(new_n7791_));
  NAND3_X1   g07512(.A1(new_n7786_), .A2(new_n7781_), .A3(new_n7791_), .ZN(new_n7792_));
  NOR2_X1    g07513(.A1(new_n7783_), .A2(new_n7785_), .ZN(new_n7793_));
  NOR2_X1    g07514(.A1(new_n7554_), .A2(new_n7780_), .ZN(new_n7794_));
  OAI21_X1   g07515(.A1(new_n7793_), .A2(new_n7794_), .B(new_n7790_), .ZN(new_n7795_));
  NAND2_X1   g07516(.A1(new_n7795_), .A2(new_n7792_), .ZN(new_n7796_));
  OAI22_X1   g07517(.A1(new_n970_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n820_), .ZN(new_n7797_));
  OAI21_X1   g07518(.A1(new_n3717_), .A2(new_n894_), .B(new_n7797_), .ZN(new_n7798_));
  AOI21_X1   g07519(.A1(new_n7798_), .A2(new_n827_), .B(new_n970_), .ZN(new_n7799_));
  XNOR2_X1   g07520(.A1(new_n4257_), .A2(new_n7799_), .ZN(new_n7800_));
  NOR2_X1    g07521(.A1(new_n7796_), .A2(new_n7800_), .ZN(new_n7801_));
  INV_X1     g07522(.I(new_n7796_), .ZN(new_n7802_));
  INV_X1     g07523(.I(new_n7800_), .ZN(new_n7803_));
  NOR2_X1    g07524(.A1(new_n7802_), .A2(new_n7803_), .ZN(new_n7804_));
  OAI21_X1   g07525(.A1(new_n7804_), .A2(new_n7801_), .B(new_n7549_), .ZN(new_n7805_));
  INV_X1     g07526(.I(new_n7549_), .ZN(new_n7806_));
  XOR2_X1    g07527(.A1(new_n7796_), .A2(new_n7800_), .Z(new_n7807_));
  NAND2_X1   g07528(.A1(new_n7807_), .A2(new_n7806_), .ZN(new_n7808_));
  NAND2_X1   g07529(.A1(new_n7808_), .A2(new_n7805_), .ZN(new_n7809_));
  OAI22_X1   g07530(.A1(new_n607_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n610_), .ZN(new_n7810_));
  OAI21_X1   g07531(.A1(new_n4500_), .A2(new_n684_), .B(new_n7810_), .ZN(new_n7811_));
  AOI21_X1   g07532(.A1(new_n7811_), .A2(new_n612_), .B(new_n607_), .ZN(new_n7812_));
  XOR2_X1    g07533(.A1(new_n5067_), .A2(new_n7812_), .Z(new_n7813_));
  INV_X1     g07534(.I(new_n7813_), .ZN(new_n7814_));
  NAND2_X1   g07535(.A1(new_n7809_), .A2(new_n7814_), .ZN(new_n7815_));
  INV_X1     g07536(.I(new_n7809_), .ZN(new_n7816_));
  NAND2_X1   g07537(.A1(new_n7816_), .A2(new_n7813_), .ZN(new_n7817_));
  AOI21_X1   g07538(.A1(new_n7817_), .A2(new_n7815_), .B(new_n7545_), .ZN(new_n7818_));
  NAND2_X1   g07539(.A1(new_n7542_), .A2(new_n7229_), .ZN(new_n7819_));
  NAND3_X1   g07540(.A1(new_n7541_), .A2(new_n7465_), .A3(new_n7543_), .ZN(new_n7820_));
  NAND2_X1   g07541(.A1(new_n7820_), .A2(new_n7819_), .ZN(new_n7821_));
  XOR2_X1    g07542(.A1(new_n7809_), .A2(new_n7813_), .Z(new_n7822_));
  NOR2_X1    g07543(.A1(new_n7822_), .A2(new_n7821_), .ZN(new_n7823_));
  NOR2_X1    g07544(.A1(new_n7823_), .A2(new_n7818_), .ZN(new_n7824_));
  XOR2_X1    g07545(.A1(new_n7540_), .A2(new_n7824_), .Z(new_n7825_));
  INV_X1     g07546(.I(new_n7825_), .ZN(new_n7826_));
  AOI21_X1   g07547(.A1(new_n7485_), .A2(new_n7488_), .B(new_n7165_), .ZN(new_n7827_));
  INV_X1     g07548(.I(new_n7827_), .ZN(new_n7828_));
  INV_X1     g07549(.I(new_n7492_), .ZN(new_n7829_));
  NAND3_X1   g07550(.A1(new_n7485_), .A2(new_n7488_), .A3(new_n7165_), .ZN(new_n7830_));
  NAND4_X1   g07551(.A1(new_n7222_), .A2(new_n7224_), .A3(new_n7830_), .A4(new_n7829_), .ZN(new_n7831_));
  OAI22_X1   g07552(.A1(new_n6538_), .A2(new_n341_), .B1(new_n404_), .B2(new_n6847_), .ZN(new_n7832_));
  OAI21_X1   g07553(.A1(new_n6229_), .A2(new_n366_), .B(new_n7832_), .ZN(new_n7833_));
  AOI21_X1   g07554(.A1(new_n7833_), .A2(new_n334_), .B(new_n341_), .ZN(new_n7834_));
  XOR2_X1    g07555(.A1(new_n6851_), .A2(new_n7834_), .Z(new_n7835_));
  INV_X1     g07556(.I(new_n7835_), .ZN(new_n7836_));
  NAND3_X1   g07557(.A1(new_n7831_), .A2(new_n7828_), .A3(new_n7836_), .ZN(new_n7837_));
  AOI21_X1   g07558(.A1(new_n7487_), .A2(new_n7486_), .B(new_n7154_), .ZN(new_n7838_));
  NOR3_X1    g07559(.A1(new_n7477_), .A2(new_n7484_), .A3(new_n7145_), .ZN(new_n7839_));
  NOR3_X1    g07560(.A1(new_n7838_), .A2(new_n7839_), .A3(new_n7216_), .ZN(new_n7840_));
  NOR4_X1    g07561(.A1(new_n7840_), .A2(new_n7497_), .A3(new_n7495_), .A4(new_n7492_), .ZN(new_n7841_));
  OAI21_X1   g07562(.A1(new_n7841_), .A2(new_n7827_), .B(new_n7835_), .ZN(new_n7842_));
  AOI21_X1   g07563(.A1(new_n7842_), .A2(new_n7837_), .B(new_n7826_), .ZN(new_n7843_));
  NOR3_X1    g07564(.A1(new_n7841_), .A2(new_n7827_), .A3(new_n7835_), .ZN(new_n7844_));
  AOI21_X1   g07565(.A1(new_n7831_), .A2(new_n7828_), .B(new_n7836_), .ZN(new_n7845_));
  NOR3_X1    g07566(.A1(new_n7844_), .A2(new_n7845_), .A3(new_n7825_), .ZN(new_n7846_));
  OAI21_X1   g07567(.A1(new_n7846_), .A2(new_n7843_), .B(new_n7536_), .ZN(new_n7847_));
  INV_X1     g07568(.I(new_n7536_), .ZN(new_n7848_));
  OAI21_X1   g07569(.A1(new_n7844_), .A2(new_n7845_), .B(new_n7825_), .ZN(new_n7849_));
  NAND3_X1   g07570(.A1(new_n7842_), .A2(new_n7837_), .A3(new_n7826_), .ZN(new_n7850_));
  NAND3_X1   g07571(.A1(new_n7849_), .A2(new_n7850_), .A3(new_n7848_), .ZN(new_n7851_));
  NAND2_X1   g07572(.A1(new_n7847_), .A2(new_n7851_), .ZN(new_n7852_));
  INV_X1     g07573(.I(new_n7852_), .ZN(new_n7853_));
  NOR2_X1    g07574(.A1(new_n7511_), .A2(new_n7853_), .ZN(new_n7854_));
  OAI21_X1   g07575(.A1(new_n7505_), .A2(new_n7509_), .B(new_n7854_), .ZN(new_n7855_));
  INV_X1     g07576(.I(new_n7855_), .ZN(new_n7856_));
  NOR2_X1    g07577(.A1(new_n7505_), .A2(new_n7509_), .ZN(new_n7857_));
  NOR2_X1    g07578(.A1(new_n7856_), .A2(new_n7857_), .ZN(new_n7858_));
  NOR2_X1    g07579(.A1(new_n7858_), .A2(new_n7532_), .ZN(new_n7859_));
  NOR3_X1    g07580(.A1(new_n7856_), .A2(new_n7221_), .A3(new_n7857_), .ZN(new_n7860_));
  NOR2_X1    g07581(.A1(new_n7859_), .A2(new_n7860_), .ZN(new_n7861_));
  NOR2_X1    g07582(.A1(\b[44] ), .A2(\b[45] ), .ZN(new_n7862_));
  AOI21_X1   g07583(.A1(new_n7196_), .A2(new_n7862_), .B(new_n6847_), .ZN(new_n7863_));
  INV_X1     g07584(.I(\b[45] ), .ZN(new_n7864_));
  NOR2_X1    g07585(.A1(new_n7198_), .A2(new_n7864_), .ZN(new_n7865_));
  INV_X1     g07586(.I(new_n7865_), .ZN(new_n7866_));
  NOR2_X1    g07587(.A1(new_n7196_), .A2(new_n7866_), .ZN(new_n7867_));
  NOR2_X1    g07588(.A1(new_n7863_), .A2(new_n7867_), .ZN(new_n7868_));
  XNOR2_X1   g07589(.A1(\b[45] ), .A2(\b[46] ), .ZN(new_n7869_));
  INV_X1     g07590(.I(\b[46] ), .ZN(new_n7870_));
  NOR2_X1    g07591(.A1(new_n7864_), .A2(new_n7870_), .ZN(new_n7871_));
  NOR2_X1    g07592(.A1(\b[45] ), .A2(\b[46] ), .ZN(new_n7872_));
  OAI21_X1   g07593(.A1(new_n7871_), .A2(new_n7872_), .B(new_n7868_), .ZN(new_n7873_));
  OAI21_X1   g07594(.A1(new_n7868_), .A2(new_n7869_), .B(new_n7873_), .ZN(new_n7874_));
  OAI22_X1   g07595(.A1(new_n330_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n263_), .ZN(new_n7875_));
  OAI21_X1   g07596(.A1(new_n7198_), .A2(new_n289_), .B(new_n7875_), .ZN(new_n7876_));
  AOI21_X1   g07597(.A1(new_n7876_), .A2(new_n260_), .B(new_n426_), .ZN(new_n7877_));
  XNOR2_X1   g07598(.A1(new_n7874_), .A2(new_n7877_), .ZN(new_n7878_));
  XOR2_X1    g07599(.A1(new_n7861_), .A2(new_n7878_), .Z(new_n7879_));
  NAND2_X1   g07600(.A1(new_n7527_), .A2(new_n7528_), .ZN(new_n7880_));
  AOI21_X1   g07601(.A1(new_n7880_), .A2(new_n7211_), .B(new_n7190_), .ZN(new_n7881_));
  NAND3_X1   g07602(.A1(new_n7527_), .A2(new_n7528_), .A3(new_n7206_), .ZN(new_n7882_));
  NAND2_X1   g07603(.A1(new_n6874_), .A2(new_n7882_), .ZN(new_n7883_));
  NOR2_X1    g07604(.A1(new_n7883_), .A2(new_n7881_), .ZN(new_n7884_));
  NOR2_X1    g07605(.A1(new_n7521_), .A2(new_n7522_), .ZN(new_n7885_));
  XOR2_X1    g07606(.A1(new_n7532_), .A2(new_n260_), .Z(new_n7886_));
  NOR2_X1    g07607(.A1(new_n7885_), .A2(new_n7886_), .ZN(new_n7887_));
  NOR2_X1    g07608(.A1(new_n7884_), .A2(new_n7887_), .ZN(new_n7888_));
  XOR2_X1    g07609(.A1(new_n7888_), .A2(new_n7879_), .Z(\f[46] ));
  OR2_X2     g07610(.A1(new_n7501_), .A2(new_n7504_), .Z(new_n7890_));
  INV_X1     g07611(.I(new_n7509_), .ZN(new_n7891_));
  AOI21_X1   g07612(.A1(new_n7852_), .A2(new_n7890_), .B(new_n7891_), .ZN(new_n7892_));
  NAND3_X1   g07613(.A1(new_n7847_), .A2(new_n7851_), .A3(new_n7505_), .ZN(new_n7893_));
  NAND2_X1   g07614(.A1(new_n7893_), .A2(new_n7532_), .ZN(new_n7894_));
  NAND2_X1   g07615(.A1(new_n7831_), .A2(new_n7828_), .ZN(new_n7895_));
  XOR2_X1    g07616(.A1(new_n7895_), .A2(new_n7825_), .Z(new_n7896_));
  NOR2_X1    g07617(.A1(new_n7896_), .A2(new_n7848_), .ZN(new_n7897_));
  XOR2_X1    g07618(.A1(new_n7895_), .A2(new_n7826_), .Z(new_n7898_));
  NOR2_X1    g07619(.A1(new_n7898_), .A2(new_n7536_), .ZN(new_n7899_));
  OAI21_X1   g07620(.A1(new_n7897_), .A2(new_n7899_), .B(new_n7836_), .ZN(new_n7900_));
  OAI21_X1   g07621(.A1(new_n7892_), .A2(new_n7894_), .B(new_n7900_), .ZN(new_n7901_));
  NOR2_X1    g07622(.A1(new_n7841_), .A2(new_n7827_), .ZN(new_n7902_));
  NAND2_X1   g07623(.A1(new_n7825_), .A2(new_n7848_), .ZN(new_n7903_));
  NOR2_X1    g07624(.A1(new_n7825_), .A2(new_n7848_), .ZN(new_n7904_));
  OAI21_X1   g07625(.A1(new_n7902_), .A2(new_n7904_), .B(new_n7903_), .ZN(new_n7905_));
  NOR2_X1    g07626(.A1(new_n7537_), .A2(new_n7145_), .ZN(new_n7906_));
  NOR2_X1    g07627(.A1(new_n7539_), .A2(new_n7479_), .ZN(new_n7907_));
  NOR2_X1    g07628(.A1(new_n7907_), .A2(new_n7906_), .ZN(new_n7908_));
  INV_X1     g07629(.I(new_n7824_), .ZN(new_n7909_));
  NOR2_X1    g07630(.A1(new_n7821_), .A2(new_n7816_), .ZN(new_n7910_));
  NOR2_X1    g07631(.A1(new_n7545_), .A2(new_n7809_), .ZN(new_n7911_));
  OAI21_X1   g07632(.A1(new_n7910_), .A2(new_n7911_), .B(new_n7813_), .ZN(new_n7912_));
  NOR2_X1    g07633(.A1(new_n7806_), .A2(new_n7802_), .ZN(new_n7913_));
  NOR2_X1    g07634(.A1(new_n7549_), .A2(new_n7796_), .ZN(new_n7914_));
  OAI21_X1   g07635(.A1(new_n7913_), .A2(new_n7914_), .B(new_n7800_), .ZN(new_n7915_));
  NAND2_X1   g07636(.A1(new_n7786_), .A2(new_n7781_), .ZN(new_n7916_));
  NAND2_X1   g07637(.A1(new_n7916_), .A2(new_n7791_), .ZN(new_n7917_));
  OAI22_X1   g07638(.A1(new_n7557_), .A2(new_n7407_), .B1(new_n7249_), .B2(new_n7555_), .ZN(new_n7918_));
  INV_X1     g07639(.I(new_n7771_), .ZN(new_n7919_));
  NOR2_X1    g07640(.A1(new_n7918_), .A2(new_n7919_), .ZN(new_n7920_));
  INV_X1     g07641(.I(new_n7920_), .ZN(new_n7921_));
  NAND2_X1   g07642(.A1(new_n7918_), .A2(new_n7919_), .ZN(new_n7922_));
  AOI21_X1   g07643(.A1(new_n7921_), .A2(new_n7922_), .B(new_n7776_), .ZN(new_n7923_));
  XOR2_X1    g07644(.A1(new_n7564_), .A2(new_n7756_), .Z(new_n7924_));
  NAND2_X1   g07645(.A1(new_n7924_), .A2(new_n7760_), .ZN(new_n7925_));
  OAI22_X1   g07646(.A1(new_n2171_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n2166_), .ZN(new_n7926_));
  OAI21_X1   g07647(.A1(new_n1634_), .A2(new_n2322_), .B(new_n7926_), .ZN(new_n7927_));
  AOI21_X1   g07648(.A1(new_n7927_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n7928_));
  XNOR2_X1   g07649(.A1(new_n1940_), .A2(new_n7928_), .ZN(new_n7929_));
  NOR2_X1    g07650(.A1(new_n7728_), .A2(new_n7723_), .ZN(new_n7930_));
  NOR2_X1    g07651(.A1(new_n7572_), .A2(new_n7741_), .ZN(new_n7931_));
  OAI21_X1   g07652(.A1(new_n7930_), .A2(new_n7931_), .B(new_n7720_), .ZN(new_n7932_));
  NAND2_X1   g07653(.A1(new_n7713_), .A2(new_n7706_), .ZN(new_n7933_));
  NAND2_X1   g07654(.A1(new_n7577_), .A2(new_n7697_), .ZN(new_n7934_));
  AOI21_X1   g07655(.A1(new_n7933_), .A2(new_n7934_), .B(new_n7702_), .ZN(new_n7935_));
  NAND2_X1   g07656(.A1(new_n7694_), .A2(new_n7693_), .ZN(new_n7936_));
  NAND2_X1   g07657(.A1(new_n7936_), .A2(new_n7695_), .ZN(new_n7937_));
  OAI21_X1   g07658(.A1(new_n7583_), .A2(new_n7674_), .B(new_n7673_), .ZN(new_n7938_));
  INV_X1     g07659(.I(new_n7633_), .ZN(new_n7939_));
  NAND2_X1   g07660(.A1(new_n7620_), .A2(new_n7621_), .ZN(new_n7940_));
  NAND2_X1   g07661(.A1(new_n7940_), .A2(\b[2] ), .ZN(new_n7941_));
  NAND2_X1   g07662(.A1(new_n7607_), .A2(new_n282_), .ZN(new_n7942_));
  NAND3_X1   g07663(.A1(new_n7614_), .A2(new_n7615_), .A3(\b[1] ), .ZN(new_n7943_));
  NAND3_X1   g07664(.A1(new_n7942_), .A2(new_n7941_), .A3(new_n7943_), .ZN(new_n7944_));
  XOR2_X1    g07665(.A1(\a[44] ), .A2(\a[45] ), .Z(new_n7945_));
  XOR2_X1    g07666(.A1(\a[44] ), .A2(\a[47] ), .Z(new_n7946_));
  NAND3_X1   g07667(.A1(new_n7945_), .A2(new_n7615_), .A3(new_n7946_), .ZN(new_n7947_));
  NOR2_X1    g07668(.A1(new_n7947_), .A2(new_n258_), .ZN(new_n7948_));
  AOI21_X1   g07669(.A1(new_n7944_), .A2(new_n7948_), .B(new_n7608_), .ZN(new_n7949_));
  INV_X1     g07670(.I(new_n7941_), .ZN(new_n7950_));
  NOR2_X1    g07671(.A1(new_n7619_), .A2(new_n490_), .ZN(new_n7951_));
  INV_X1     g07672(.I(new_n7943_), .ZN(new_n7952_));
  NOR3_X1    g07673(.A1(new_n7951_), .A2(new_n7950_), .A3(new_n7952_), .ZN(new_n7953_));
  INV_X1     g07674(.I(new_n7948_), .ZN(new_n7954_));
  NOR3_X1    g07675(.A1(new_n7953_), .A2(\a[47] ), .A3(new_n7954_), .ZN(new_n7955_));
  NOR2_X1    g07676(.A1(new_n7955_), .A2(new_n7949_), .ZN(new_n7956_));
  NOR3_X1    g07677(.A1(new_n7629_), .A2(new_n7630_), .A3(new_n7627_), .ZN(new_n7957_));
  OAI21_X1   g07678(.A1(new_n2332_), .A2(new_n2331_), .B(new_n6631_), .ZN(new_n7958_));
  OAI22_X1   g07679(.A1(new_n6644_), .A2(new_n325_), .B1(new_n419_), .B2(new_n6647_), .ZN(new_n7959_));
  NAND4_X1   g07680(.A1(new_n6640_), .A2(new_n7282_), .A3(new_n7283_), .A4(\b[3] ), .ZN(new_n7960_));
  NAND3_X1   g07681(.A1(new_n7958_), .A2(new_n7959_), .A3(new_n7960_), .ZN(new_n7961_));
  NOR2_X1    g07682(.A1(new_n7957_), .A2(new_n7961_), .ZN(new_n7962_));
  NAND3_X1   g07683(.A1(new_n7625_), .A2(new_n7618_), .A3(new_n7626_), .ZN(new_n7963_));
  AOI21_X1   g07684(.A1(new_n374_), .A2(new_n377_), .B(new_n6644_), .ZN(new_n7964_));
  NAND2_X1   g07685(.A1(new_n7959_), .A2(new_n7960_), .ZN(new_n7965_));
  NOR2_X1    g07686(.A1(new_n7965_), .A2(new_n7964_), .ZN(new_n7966_));
  NOR2_X1    g07687(.A1(new_n7963_), .A2(new_n7966_), .ZN(new_n7967_));
  OAI21_X1   g07688(.A1(new_n7962_), .A2(new_n7967_), .B(new_n7956_), .ZN(new_n7968_));
  OAI21_X1   g07689(.A1(new_n7953_), .A2(new_n7954_), .B(\a[47] ), .ZN(new_n7969_));
  NAND3_X1   g07690(.A1(new_n7944_), .A2(new_n7608_), .A3(new_n7948_), .ZN(new_n7970_));
  NAND2_X1   g07691(.A1(new_n7969_), .A2(new_n7970_), .ZN(new_n7971_));
  NAND2_X1   g07692(.A1(new_n7963_), .A2(new_n7966_), .ZN(new_n7972_));
  NAND4_X1   g07693(.A1(new_n7961_), .A2(new_n7618_), .A3(new_n7625_), .A4(new_n7626_), .ZN(new_n7973_));
  NAND3_X1   g07694(.A1(new_n7972_), .A2(new_n7973_), .A3(new_n7971_), .ZN(new_n7974_));
  AOI21_X1   g07695(.A1(new_n7968_), .A2(new_n7974_), .B(\a[44] ), .ZN(new_n7975_));
  AOI21_X1   g07696(.A1(new_n7972_), .A2(new_n7973_), .B(new_n7971_), .ZN(new_n7976_));
  NOR3_X1    g07697(.A1(new_n7962_), .A2(new_n7967_), .A3(new_n7956_), .ZN(new_n7977_));
  NOR3_X1    g07698(.A1(new_n7977_), .A2(new_n7976_), .A3(new_n6632_), .ZN(new_n7978_));
  OAI21_X1   g07699(.A1(new_n7978_), .A2(new_n7975_), .B(new_n7645_), .ZN(new_n7979_));
  NOR2_X1    g07700(.A1(new_n7979_), .A2(new_n7939_), .ZN(new_n7980_));
  OAI21_X1   g07701(.A1(new_n7977_), .A2(new_n7976_), .B(new_n6632_), .ZN(new_n7981_));
  NAND3_X1   g07702(.A1(new_n7968_), .A2(new_n7974_), .A3(\a[44] ), .ZN(new_n7982_));
  NAND2_X1   g07703(.A1(new_n7981_), .A2(new_n7982_), .ZN(new_n7983_));
  NAND2_X1   g07704(.A1(new_n7604_), .A2(new_n7632_), .ZN(new_n7985_));
  INV_X1     g07705(.I(new_n7985_), .ZN(new_n7986_));
  OAI21_X1   g07706(.A1(new_n7980_), .A2(new_n7986_), .B(new_n7642_), .ZN(new_n7987_));
  NAND3_X1   g07707(.A1(new_n7983_), .A2(new_n7633_), .A3(new_n7645_), .ZN(new_n7988_));
  NAND3_X1   g07708(.A1(new_n7988_), .A2(new_n7595_), .A3(new_n7985_), .ZN(new_n7989_));
  OAI22_X1   g07709(.A1(new_n5993_), .A2(new_n472_), .B1(new_n515_), .B2(new_n5991_), .ZN(new_n7990_));
  OAI21_X1   g07710(.A1(new_n420_), .A2(new_n5997_), .B(new_n7990_), .ZN(new_n7991_));
  AOI21_X1   g07711(.A1(new_n7991_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n7992_));
  XOR2_X1    g07712(.A1(new_n700_), .A2(new_n7992_), .Z(new_n7993_));
  INV_X1     g07713(.I(new_n7993_), .ZN(new_n7994_));
  NAND3_X1   g07714(.A1(new_n7987_), .A2(new_n7989_), .A3(new_n7994_), .ZN(new_n7995_));
  AOI21_X1   g07715(.A1(new_n7988_), .A2(new_n7985_), .B(new_n7595_), .ZN(new_n7996_));
  NOR3_X1    g07716(.A1(new_n7980_), .A2(new_n7642_), .A3(new_n7986_), .ZN(new_n7997_));
  OAI21_X1   g07717(.A1(new_n7997_), .A2(new_n7996_), .B(new_n7993_), .ZN(new_n7998_));
  NAND2_X1   g07718(.A1(new_n7998_), .A2(new_n7995_), .ZN(new_n7999_));
  NAND3_X1   g07719(.A1(new_n7999_), .A2(new_n7654_), .A3(new_n7664_), .ZN(new_n8000_));
  NAND2_X1   g07720(.A1(new_n7647_), .A2(new_n7653_), .ZN(new_n8002_));
  AOI21_X1   g07721(.A1(new_n8000_), .A2(new_n8002_), .B(new_n7661_), .ZN(new_n8003_));
  NOR3_X1    g07722(.A1(new_n7997_), .A2(new_n7996_), .A3(new_n7993_), .ZN(new_n8004_));
  AOI21_X1   g07723(.A1(new_n7987_), .A2(new_n7989_), .B(new_n7994_), .ZN(new_n8005_));
  OAI21_X1   g07724(.A1(new_n8004_), .A2(new_n8005_), .B(new_n7664_), .ZN(new_n8006_));
  NOR2_X1    g07725(.A1(new_n8006_), .A2(new_n7655_), .ZN(new_n8007_));
  INV_X1     g07726(.I(new_n8002_), .ZN(new_n8008_));
  NOR3_X1    g07727(.A1(new_n8007_), .A2(new_n7590_), .A3(new_n8008_), .ZN(new_n8009_));
  OAI22_X1   g07728(.A1(new_n5420_), .A2(new_n656_), .B1(new_n706_), .B2(new_n5107_), .ZN(new_n8010_));
  OAI21_X1   g07729(.A1(new_n565_), .A2(new_n5112_), .B(new_n8010_), .ZN(new_n8011_));
  AOI21_X1   g07730(.A1(new_n8011_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n8012_));
  XNOR2_X1   g07731(.A1(new_n710_), .A2(new_n8012_), .ZN(new_n8013_));
  NOR3_X1    g07732(.A1(new_n8009_), .A2(new_n8003_), .A3(new_n8013_), .ZN(new_n8014_));
  OAI21_X1   g07733(.A1(new_n8007_), .A2(new_n8008_), .B(new_n7590_), .ZN(new_n8015_));
  NAND3_X1   g07734(.A1(new_n8000_), .A2(new_n7661_), .A3(new_n8002_), .ZN(new_n8016_));
  INV_X1     g07735(.I(new_n8013_), .ZN(new_n8017_));
  AOI21_X1   g07736(.A1(new_n8015_), .A2(new_n8016_), .B(new_n8017_), .ZN(new_n8018_));
  OAI22_X1   g07737(.A1(new_n4072_), .A2(new_n861_), .B1(new_n930_), .B2(new_n4067_), .ZN(new_n8019_));
  OAI21_X1   g07738(.A1(new_n780_), .A2(new_n4318_), .B(new_n8019_), .ZN(new_n8020_));
  AOI21_X1   g07739(.A1(new_n8020_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n8021_));
  XNOR2_X1   g07740(.A1(new_n937_), .A2(new_n8021_), .ZN(new_n8022_));
  NOR3_X1    g07741(.A1(new_n8014_), .A2(new_n8018_), .A3(new_n8022_), .ZN(new_n8023_));
  NAND3_X1   g07742(.A1(new_n8015_), .A2(new_n8016_), .A3(new_n8017_), .ZN(new_n8024_));
  OAI21_X1   g07743(.A1(new_n8009_), .A2(new_n8003_), .B(new_n8013_), .ZN(new_n8025_));
  INV_X1     g07744(.I(new_n8022_), .ZN(new_n8026_));
  AOI21_X1   g07745(.A1(new_n8025_), .A2(new_n8024_), .B(new_n8026_), .ZN(new_n8027_));
  OAI21_X1   g07746(.A1(new_n8023_), .A2(new_n8027_), .B(new_n7938_), .ZN(new_n8028_));
  AOI21_X1   g07747(.A1(new_n7681_), .A2(new_n7675_), .B(new_n7692_), .ZN(new_n8029_));
  AOI21_X1   g07748(.A1(new_n8025_), .A2(new_n8024_), .B(new_n8022_), .ZN(new_n8030_));
  NOR3_X1    g07749(.A1(new_n8014_), .A2(new_n8018_), .A3(new_n8026_), .ZN(new_n8031_));
  OAI21_X1   g07750(.A1(new_n8030_), .A2(new_n8031_), .B(new_n8029_), .ZN(new_n8032_));
  NAND2_X1   g07751(.A1(new_n8032_), .A2(new_n8028_), .ZN(new_n8033_));
  NAND3_X1   g07752(.A1(new_n7706_), .A2(new_n8033_), .A3(new_n7937_), .ZN(new_n8034_));
  NOR2_X1    g07753(.A1(new_n7676_), .A2(new_n7685_), .ZN(new_n8035_));
  NAND2_X1   g07754(.A1(new_n8025_), .A2(new_n8024_), .ZN(new_n8036_));
  INV_X1     g07755(.I(new_n8036_), .ZN(new_n8037_));
  NOR2_X1    g07756(.A1(new_n8035_), .A2(new_n7689_), .ZN(new_n8038_));
  INV_X1     g07757(.I(new_n8038_), .ZN(new_n8039_));
  AOI21_X1   g07758(.A1(new_n8034_), .A2(new_n8039_), .B(new_n7713_), .ZN(new_n8040_));
  NOR2_X1    g07759(.A1(new_n8035_), .A2(new_n7689_), .ZN(new_n8041_));
  NAND3_X1   g07760(.A1(new_n8025_), .A2(new_n8024_), .A3(new_n8026_), .ZN(new_n8042_));
  OAI21_X1   g07761(.A1(new_n8014_), .A2(new_n8018_), .B(new_n8022_), .ZN(new_n8043_));
  AOI21_X1   g07762(.A1(new_n8042_), .A2(new_n8043_), .B(new_n8029_), .ZN(new_n8044_));
  OAI21_X1   g07763(.A1(new_n8014_), .A2(new_n8018_), .B(new_n8026_), .ZN(new_n8045_));
  NAND3_X1   g07764(.A1(new_n8025_), .A2(new_n8024_), .A3(new_n8022_), .ZN(new_n8046_));
  AOI21_X1   g07765(.A1(new_n8045_), .A2(new_n8046_), .B(new_n7938_), .ZN(new_n8047_));
  NOR2_X1    g07766(.A1(new_n8044_), .A2(new_n8047_), .ZN(new_n8048_));
  NOR3_X1    g07767(.A1(new_n7697_), .A2(new_n8048_), .A3(new_n8041_), .ZN(new_n8049_));
  NOR3_X1    g07768(.A1(new_n8049_), .A2(new_n7577_), .A3(new_n8038_), .ZN(new_n8050_));
  OAI22_X1   g07769(.A1(new_n1109_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1189_), .ZN(new_n8051_));
  OAI21_X1   g07770(.A1(new_n1017_), .A2(new_n3569_), .B(new_n8051_), .ZN(new_n8052_));
  AOI21_X1   g07771(.A1(new_n8052_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n8053_));
  XNOR2_X1   g07772(.A1(new_n1196_), .A2(new_n8053_), .ZN(new_n8054_));
  NOR3_X1    g07773(.A1(new_n8040_), .A2(new_n8050_), .A3(new_n8054_), .ZN(new_n8055_));
  OAI21_X1   g07774(.A1(new_n8049_), .A2(new_n8038_), .B(new_n7577_), .ZN(new_n8056_));
  NAND3_X1   g07775(.A1(new_n8034_), .A2(new_n7713_), .A3(new_n8039_), .ZN(new_n8057_));
  INV_X1     g07776(.I(new_n8054_), .ZN(new_n8058_));
  AOI21_X1   g07777(.A1(new_n8056_), .A2(new_n8057_), .B(new_n8058_), .ZN(new_n8059_));
  NOR3_X1    g07778(.A1(new_n8055_), .A2(new_n8059_), .A3(new_n7935_), .ZN(new_n8060_));
  NOR3_X1    g07779(.A1(new_n8060_), .A2(new_n7728_), .A3(new_n7723_), .ZN(new_n8061_));
  NOR2_X1    g07780(.A1(new_n7577_), .A2(new_n7697_), .ZN(new_n8062_));
  NOR2_X1    g07781(.A1(new_n7713_), .A2(new_n7706_), .ZN(new_n8063_));
  OAI21_X1   g07782(.A1(new_n8063_), .A2(new_n8062_), .B(new_n7701_), .ZN(new_n8064_));
  NAND3_X1   g07783(.A1(new_n8056_), .A2(new_n8057_), .A3(new_n8058_), .ZN(new_n8065_));
  OAI21_X1   g07784(.A1(new_n8040_), .A2(new_n8050_), .B(new_n8054_), .ZN(new_n8066_));
  NAND3_X1   g07785(.A1(new_n8066_), .A2(new_n8065_), .A3(new_n8064_), .ZN(new_n8067_));
  AOI21_X1   g07786(.A1(new_n8067_), .A2(new_n7741_), .B(new_n7572_), .ZN(new_n8068_));
  OAI22_X1   g07787(.A1(new_n1518_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1525_), .ZN(new_n8069_));
  OAI21_X1   g07788(.A1(new_n1294_), .A2(new_n2884_), .B(new_n8069_), .ZN(new_n8070_));
  AOI21_X1   g07789(.A1(new_n8070_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n8071_));
  XOR2_X1    g07790(.A1(new_n1530_), .A2(new_n8071_), .Z(new_n8072_));
  INV_X1     g07791(.I(new_n8072_), .ZN(new_n8073_));
  OAI21_X1   g07792(.A1(new_n8061_), .A2(new_n8068_), .B(new_n8073_), .ZN(new_n8074_));
  NAND3_X1   g07793(.A1(new_n8067_), .A2(new_n7572_), .A3(new_n7741_), .ZN(new_n8075_));
  OAI21_X1   g07794(.A1(new_n8060_), .A2(new_n7723_), .B(new_n7728_), .ZN(new_n8076_));
  NAND3_X1   g07795(.A1(new_n8076_), .A2(new_n8075_), .A3(new_n8072_), .ZN(new_n8077_));
  NAND3_X1   g07796(.A1(new_n8074_), .A2(new_n8077_), .A3(new_n7932_), .ZN(new_n8078_));
  NAND3_X1   g07797(.A1(new_n8078_), .A2(new_n7750_), .A3(new_n7751_), .ZN(new_n8079_));
  NAND2_X1   g07798(.A1(new_n7572_), .A2(new_n7741_), .ZN(new_n8080_));
  NAND2_X1   g07799(.A1(new_n7728_), .A2(new_n7723_), .ZN(new_n8081_));
  AOI21_X1   g07800(.A1(new_n8081_), .A2(new_n8080_), .B(new_n7721_), .ZN(new_n8082_));
  AOI21_X1   g07801(.A1(new_n8076_), .A2(new_n8075_), .B(new_n8072_), .ZN(new_n8083_));
  NOR3_X1    g07802(.A1(new_n8061_), .A2(new_n8068_), .A3(new_n8073_), .ZN(new_n8084_));
  NOR3_X1    g07803(.A1(new_n8084_), .A2(new_n8083_), .A3(new_n8082_), .ZN(new_n8085_));
  OAI21_X1   g07804(.A1(new_n8085_), .A2(new_n7753_), .B(new_n7568_), .ZN(new_n8086_));
  NAND2_X1   g07805(.A1(new_n8086_), .A2(new_n8079_), .ZN(new_n8087_));
  XOR2_X1    g07806(.A1(new_n7568_), .A2(new_n7753_), .Z(new_n8088_));
  NOR2_X1    g07807(.A1(new_n8088_), .A2(new_n7737_), .ZN(new_n8089_));
  NOR3_X1    g07808(.A1(new_n7766_), .A2(new_n7560_), .A3(new_n7756_), .ZN(new_n8090_));
  OAI22_X1   g07809(.A1(new_n1712_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n1707_), .ZN(new_n8091_));
  OAI21_X1   g07810(.A1(new_n2102_), .A2(new_n1850_), .B(new_n8091_), .ZN(new_n8092_));
  AOI21_X1   g07811(.A1(new_n8092_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n8093_));
  XNOR2_X1   g07812(.A1(new_n2443_), .A2(new_n8093_), .ZN(new_n8094_));
  INV_X1     g07813(.I(new_n8094_), .ZN(new_n8095_));
  OAI21_X1   g07814(.A1(new_n8090_), .A2(new_n8089_), .B(new_n8095_), .ZN(new_n8096_));
  XOR2_X1    g07815(.A1(new_n7568_), .A2(new_n7751_), .Z(new_n8097_));
  NAND2_X1   g07816(.A1(new_n8097_), .A2(new_n7736_), .ZN(new_n8098_));
  AOI21_X1   g07817(.A1(new_n7738_), .A2(new_n7744_), .B(new_n7750_), .ZN(new_n8099_));
  NAND2_X1   g07818(.A1(new_n7753_), .A2(new_n7737_), .ZN(new_n8100_));
  NAND2_X1   g07819(.A1(new_n7751_), .A2(new_n7736_), .ZN(new_n8101_));
  AOI21_X1   g07820(.A1(new_n8100_), .A2(new_n8101_), .B(new_n7568_), .ZN(new_n8102_));
  NOR2_X1    g07821(.A1(new_n8099_), .A2(new_n8102_), .ZN(new_n8103_));
  NAND3_X1   g07822(.A1(new_n7563_), .A2(new_n7561_), .A3(new_n8103_), .ZN(new_n8104_));
  NAND3_X1   g07823(.A1(new_n8104_), .A2(new_n8098_), .A3(new_n8094_), .ZN(new_n8105_));
  AOI21_X1   g07824(.A1(new_n8096_), .A2(new_n8105_), .B(new_n8087_), .ZN(new_n8106_));
  NOR3_X1    g07825(.A1(new_n8085_), .A2(new_n7568_), .A3(new_n7753_), .ZN(new_n8107_));
  AOI21_X1   g07826(.A1(new_n8078_), .A2(new_n7751_), .B(new_n7750_), .ZN(new_n8108_));
  NOR2_X1    g07827(.A1(new_n8108_), .A2(new_n8107_), .ZN(new_n8109_));
  AOI21_X1   g07828(.A1(new_n8104_), .A2(new_n8098_), .B(new_n8094_), .ZN(new_n8110_));
  NOR3_X1    g07829(.A1(new_n8090_), .A2(new_n8089_), .A3(new_n8095_), .ZN(new_n8111_));
  NOR3_X1    g07830(.A1(new_n8111_), .A2(new_n8110_), .A3(new_n8109_), .ZN(new_n8112_));
  OAI21_X1   g07831(.A1(new_n8112_), .A2(new_n8106_), .B(new_n7929_), .ZN(new_n8113_));
  INV_X1     g07832(.I(new_n7929_), .ZN(new_n8114_));
  OAI21_X1   g07833(.A1(new_n8111_), .A2(new_n8110_), .B(new_n8109_), .ZN(new_n8115_));
  NAND3_X1   g07834(.A1(new_n8096_), .A2(new_n8105_), .A3(new_n8087_), .ZN(new_n8116_));
  NAND3_X1   g07835(.A1(new_n8115_), .A2(new_n8116_), .A3(new_n8114_), .ZN(new_n8117_));
  NAND3_X1   g07836(.A1(new_n8113_), .A2(new_n8117_), .A3(new_n7925_), .ZN(new_n8118_));
  NAND3_X1   g07837(.A1(new_n8118_), .A2(new_n7559_), .A3(new_n7771_), .ZN(new_n8119_));
  XOR2_X1    g07838(.A1(new_n7564_), .A2(new_n8103_), .Z(new_n8120_));
  NOR2_X1    g07839(.A1(new_n8120_), .A2(new_n7768_), .ZN(new_n8121_));
  AOI21_X1   g07840(.A1(new_n8115_), .A2(new_n8116_), .B(new_n8114_), .ZN(new_n8122_));
  NOR3_X1    g07841(.A1(new_n8112_), .A2(new_n8106_), .A3(new_n7929_), .ZN(new_n8123_));
  NOR3_X1    g07842(.A1(new_n8123_), .A2(new_n8122_), .A3(new_n8121_), .ZN(new_n8124_));
  OAI21_X1   g07843(.A1(new_n8124_), .A2(new_n7919_), .B(new_n7918_), .ZN(new_n8125_));
  OAI22_X1   g07844(.A1(new_n1347_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n1344_), .ZN(new_n8126_));
  OAI21_X1   g07845(.A1(new_n2643_), .A2(new_n1457_), .B(new_n8126_), .ZN(new_n8127_));
  AOI21_X1   g07846(.A1(new_n8127_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n8128_));
  XNOR2_X1   g07847(.A1(new_n3022_), .A2(new_n8128_), .ZN(new_n8129_));
  AOI21_X1   g07848(.A1(new_n8125_), .A2(new_n8119_), .B(new_n8129_), .ZN(new_n8130_));
  NOR3_X1    g07849(.A1(new_n8124_), .A2(new_n7918_), .A3(new_n7919_), .ZN(new_n8131_));
  AOI21_X1   g07850(.A1(new_n8118_), .A2(new_n7771_), .B(new_n7559_), .ZN(new_n8132_));
  INV_X1     g07851(.I(new_n8129_), .ZN(new_n8133_));
  NOR3_X1    g07852(.A1(new_n8131_), .A2(new_n8132_), .A3(new_n8133_), .ZN(new_n8134_));
  NOR3_X1    g07853(.A1(new_n8134_), .A2(new_n8130_), .A3(new_n7923_), .ZN(new_n8135_));
  NOR3_X1    g07854(.A1(new_n8135_), .A2(new_n7554_), .A3(new_n7785_), .ZN(new_n8136_));
  INV_X1     g07855(.I(new_n7922_), .ZN(new_n8137_));
  OAI21_X1   g07856(.A1(new_n8137_), .A2(new_n7920_), .B(new_n7775_), .ZN(new_n8138_));
  OAI21_X1   g07857(.A1(new_n8131_), .A2(new_n8132_), .B(new_n8133_), .ZN(new_n8139_));
  NAND3_X1   g07858(.A1(new_n8125_), .A2(new_n8119_), .A3(new_n8129_), .ZN(new_n8140_));
  NAND3_X1   g07859(.A1(new_n8139_), .A2(new_n8140_), .A3(new_n8138_), .ZN(new_n8141_));
  AOI21_X1   g07860(.A1(new_n8141_), .A2(new_n7780_), .B(new_n7783_), .ZN(new_n8142_));
  OAI22_X1   g07861(.A1(new_n1055_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n1061_), .ZN(new_n8143_));
  OAI21_X1   g07862(.A1(new_n3260_), .A2(new_n1332_), .B(new_n8143_), .ZN(new_n8144_));
  AOI21_X1   g07863(.A1(new_n8144_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n8145_));
  XOR2_X1    g07864(.A1(new_n3722_), .A2(new_n8145_), .Z(new_n8146_));
  INV_X1     g07865(.I(new_n8146_), .ZN(new_n8147_));
  OAI21_X1   g07866(.A1(new_n8136_), .A2(new_n8142_), .B(new_n8147_), .ZN(new_n8148_));
  NAND3_X1   g07867(.A1(new_n8141_), .A2(new_n7783_), .A3(new_n7780_), .ZN(new_n8149_));
  OAI21_X1   g07868(.A1(new_n8135_), .A2(new_n7785_), .B(new_n7554_), .ZN(new_n8150_));
  NAND3_X1   g07869(.A1(new_n8150_), .A2(new_n8149_), .A3(new_n8146_), .ZN(new_n8151_));
  NAND2_X1   g07870(.A1(new_n8148_), .A2(new_n8151_), .ZN(new_n8152_));
  NAND3_X1   g07871(.A1(new_n8152_), .A2(new_n7796_), .A3(new_n7917_), .ZN(new_n8153_));
  AOI21_X1   g07872(.A1(new_n8150_), .A2(new_n8149_), .B(new_n8146_), .ZN(new_n8154_));
  NOR3_X1    g07873(.A1(new_n8136_), .A2(new_n8142_), .A3(new_n8147_), .ZN(new_n8155_));
  NAND2_X1   g07874(.A1(new_n7916_), .A2(new_n7791_), .ZN(new_n8156_));
  AOI21_X1   g07875(.A1(new_n8153_), .A2(new_n8156_), .B(new_n7549_), .ZN(new_n8157_));
  INV_X1     g07876(.I(new_n8157_), .ZN(new_n8158_));
  NAND3_X1   g07877(.A1(new_n8153_), .A2(new_n7549_), .A3(new_n8156_), .ZN(new_n8159_));
  OAI22_X1   g07878(.A1(new_n970_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n820_), .ZN(new_n8160_));
  OAI21_X1   g07879(.A1(new_n3989_), .A2(new_n894_), .B(new_n8160_), .ZN(new_n8161_));
  AOI21_X1   g07880(.A1(new_n8161_), .A2(new_n827_), .B(new_n970_), .ZN(new_n8162_));
  XOR2_X1    g07881(.A1(new_n4499_), .A2(new_n8162_), .Z(new_n8163_));
  INV_X1     g07882(.I(new_n8163_), .ZN(new_n8164_));
  NAND3_X1   g07883(.A1(new_n8158_), .A2(new_n8159_), .A3(new_n8164_), .ZN(new_n8165_));
  INV_X1     g07884(.I(new_n8159_), .ZN(new_n8166_));
  OAI21_X1   g07885(.A1(new_n8166_), .A2(new_n8157_), .B(new_n8163_), .ZN(new_n8167_));
  NAND3_X1   g07886(.A1(new_n8165_), .A2(new_n8167_), .A3(new_n7915_), .ZN(new_n8168_));
  NAND3_X1   g07887(.A1(new_n8168_), .A2(new_n7545_), .A3(new_n7809_), .ZN(new_n8169_));
  INV_X1     g07888(.I(new_n7915_), .ZN(new_n8170_));
  NOR3_X1    g07889(.A1(new_n8166_), .A2(new_n8157_), .A3(new_n8163_), .ZN(new_n8171_));
  AOI21_X1   g07890(.A1(new_n8158_), .A2(new_n8159_), .B(new_n8164_), .ZN(new_n8172_));
  NOR3_X1    g07891(.A1(new_n8172_), .A2(new_n8171_), .A3(new_n8170_), .ZN(new_n8173_));
  OAI21_X1   g07892(.A1(new_n8173_), .A2(new_n7816_), .B(new_n7821_), .ZN(new_n8174_));
  OAI22_X1   g07893(.A1(new_n607_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n610_), .ZN(new_n8175_));
  OAI21_X1   g07894(.A1(new_n4774_), .A2(new_n684_), .B(new_n8175_), .ZN(new_n8176_));
  AOI21_X1   g07895(.A1(new_n8176_), .A2(new_n612_), .B(new_n607_), .ZN(new_n8177_));
  XNOR2_X1   g07896(.A1(new_n5357_), .A2(new_n8177_), .ZN(new_n8178_));
  INV_X1     g07897(.I(new_n8178_), .ZN(new_n8179_));
  NAND3_X1   g07898(.A1(new_n8174_), .A2(new_n8169_), .A3(new_n8179_), .ZN(new_n8180_));
  NOR3_X1    g07899(.A1(new_n8173_), .A2(new_n7821_), .A3(new_n7816_), .ZN(new_n8181_));
  AOI21_X1   g07900(.A1(new_n8168_), .A2(new_n7809_), .B(new_n7545_), .ZN(new_n8182_));
  OAI21_X1   g07901(.A1(new_n8181_), .A2(new_n8182_), .B(new_n8178_), .ZN(new_n8183_));
  NAND3_X1   g07902(.A1(new_n8183_), .A2(new_n8180_), .A3(new_n7912_), .ZN(new_n8184_));
  NAND3_X1   g07903(.A1(new_n8184_), .A2(new_n7909_), .A3(new_n7908_), .ZN(new_n8185_));
  NAND2_X1   g07904(.A1(new_n7545_), .A2(new_n7809_), .ZN(new_n8186_));
  INV_X1     g07905(.I(new_n7911_), .ZN(new_n8187_));
  AOI21_X1   g07906(.A1(new_n8187_), .A2(new_n8186_), .B(new_n7814_), .ZN(new_n8188_));
  NOR3_X1    g07907(.A1(new_n8181_), .A2(new_n8182_), .A3(new_n8178_), .ZN(new_n8189_));
  AOI21_X1   g07908(.A1(new_n8174_), .A2(new_n8169_), .B(new_n8179_), .ZN(new_n8190_));
  NOR3_X1    g07909(.A1(new_n8188_), .A2(new_n8189_), .A3(new_n8190_), .ZN(new_n8191_));
  OAI21_X1   g07910(.A1(new_n8191_), .A2(new_n7824_), .B(new_n7540_), .ZN(new_n8192_));
  OAI22_X1   g07911(.A1(new_n448_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n450_), .ZN(new_n8193_));
  OAI21_X1   g07912(.A1(new_n5913_), .A2(new_n496_), .B(new_n8193_), .ZN(new_n8194_));
  AOI21_X1   g07913(.A1(new_n8194_), .A2(new_n452_), .B(new_n448_), .ZN(new_n8195_));
  XOR2_X1    g07914(.A1(new_n6233_), .A2(new_n8195_), .Z(new_n8196_));
  INV_X1     g07915(.I(new_n8196_), .ZN(new_n8197_));
  NAND3_X1   g07916(.A1(new_n8192_), .A2(new_n8185_), .A3(new_n8197_), .ZN(new_n8198_));
  AOI21_X1   g07917(.A1(new_n8192_), .A2(new_n8185_), .B(new_n8197_), .ZN(new_n8199_));
  INV_X1     g07918(.I(new_n8199_), .ZN(new_n8200_));
  NAND2_X1   g07919(.A1(new_n8200_), .A2(new_n8198_), .ZN(new_n8201_));
  AND2_X2    g07920(.A1(new_n7905_), .A2(new_n8201_), .Z(new_n8202_));
  AOI21_X1   g07921(.A1(new_n8192_), .A2(new_n8185_), .B(new_n8196_), .ZN(new_n8203_));
  NOR3_X1    g07922(.A1(new_n8191_), .A2(new_n7540_), .A3(new_n7824_), .ZN(new_n8204_));
  AOI21_X1   g07923(.A1(new_n8184_), .A2(new_n7909_), .B(new_n7908_), .ZN(new_n8205_));
  NOR3_X1    g07924(.A1(new_n8204_), .A2(new_n8205_), .A3(new_n8197_), .ZN(new_n8206_));
  NOR2_X1    g07925(.A1(new_n8206_), .A2(new_n8203_), .ZN(new_n8207_));
  NOR2_X1    g07926(.A1(new_n7905_), .A2(new_n8207_), .ZN(new_n8208_));
  NOR2_X1    g07927(.A1(new_n8202_), .A2(new_n8208_), .ZN(new_n8209_));
  OAI22_X1   g07928(.A1(new_n6847_), .A2(new_n341_), .B1(new_n404_), .B2(new_n7198_), .ZN(new_n8210_));
  OAI21_X1   g07929(.A1(new_n6538_), .A2(new_n366_), .B(new_n8210_), .ZN(new_n8211_));
  AOI21_X1   g07930(.A1(new_n8211_), .A2(new_n334_), .B(new_n341_), .ZN(new_n8212_));
  XNOR2_X1   g07931(.A1(new_n7202_), .A2(new_n8212_), .ZN(new_n8213_));
  XNOR2_X1   g07932(.A1(new_n8209_), .A2(new_n8213_), .ZN(new_n8214_));
  XNOR2_X1   g07933(.A1(\b[45] ), .A2(\b[47] ), .ZN(new_n8215_));
  NOR2_X1    g07934(.A1(new_n8215_), .A2(new_n7869_), .ZN(new_n8216_));
  XOR2_X1    g07935(.A1(new_n7868_), .A2(new_n8216_), .Z(new_n8217_));
  INV_X1     g07936(.I(\b[47] ), .ZN(new_n8218_));
  OAI22_X1   g07937(.A1(new_n330_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n263_), .ZN(new_n8219_));
  OAI21_X1   g07938(.A1(new_n7864_), .A2(new_n289_), .B(new_n8219_), .ZN(new_n8220_));
  AOI21_X1   g07939(.A1(new_n8220_), .A2(new_n260_), .B(new_n426_), .ZN(new_n8221_));
  XOR2_X1    g07940(.A1(new_n8217_), .A2(new_n8221_), .Z(new_n8222_));
  INV_X1     g07941(.I(new_n8222_), .ZN(new_n8223_));
  XOR2_X1    g07942(.A1(new_n8214_), .A2(new_n8223_), .Z(new_n8224_));
  XOR2_X1    g07943(.A1(new_n8214_), .A2(new_n8222_), .Z(new_n8225_));
  MUX2_X1    g07944(.I0(new_n8224_), .I1(new_n8225_), .S(new_n7901_), .Z(new_n8226_));
  NOR3_X1    g07945(.A1(new_n7861_), .A2(new_n7885_), .A3(new_n7886_), .ZN(new_n8227_));
  INV_X1     g07946(.I(new_n7887_), .ZN(new_n8228_));
  AOI21_X1   g07947(.A1(new_n7861_), .A2(new_n8228_), .B(new_n7878_), .ZN(new_n8229_));
  AOI21_X1   g07948(.A1(new_n7884_), .A2(new_n8229_), .B(new_n8227_), .ZN(new_n8230_));
  XOR2_X1    g07949(.A1(new_n8230_), .A2(new_n8226_), .Z(\f[47] ));
  XOR2_X1    g07950(.A1(new_n8214_), .A2(new_n7901_), .Z(new_n8232_));
  NOR2_X1    g07951(.A1(new_n8232_), .A2(new_n8223_), .ZN(new_n8233_));
  AOI21_X1   g07952(.A1(new_n7849_), .A2(new_n7850_), .B(new_n7848_), .ZN(new_n8234_));
  NOR3_X1    g07953(.A1(new_n7846_), .A2(new_n7843_), .A3(new_n7536_), .ZN(new_n8235_));
  OAI21_X1   g07954(.A1(new_n8235_), .A2(new_n8234_), .B(new_n7890_), .ZN(new_n8236_));
  NAND2_X1   g07955(.A1(new_n8236_), .A2(new_n7509_), .ZN(new_n8237_));
  NOR3_X1    g07956(.A1(new_n8235_), .A2(new_n8234_), .A3(new_n7890_), .ZN(new_n8238_));
  NOR2_X1    g07957(.A1(new_n7221_), .A2(new_n8238_), .ZN(new_n8239_));
  INV_X1     g07958(.I(new_n8209_), .ZN(new_n8240_));
  NAND3_X1   g07959(.A1(new_n8239_), .A2(new_n8237_), .A3(new_n8240_), .ZN(new_n8241_));
  AOI21_X1   g07960(.A1(new_n8239_), .A2(new_n8237_), .B(new_n8240_), .ZN(new_n8242_));
  NOR2_X1    g07961(.A1(new_n7900_), .A2(new_n8213_), .ZN(new_n8243_));
  INV_X1     g07962(.I(new_n8243_), .ZN(new_n8244_));
  OAI21_X1   g07963(.A1(new_n8242_), .A2(new_n8244_), .B(new_n8241_), .ZN(new_n8245_));
  OAI21_X1   g07964(.A1(new_n8204_), .A2(new_n8205_), .B(new_n8197_), .ZN(new_n8246_));
  NAND3_X1   g07965(.A1(new_n8192_), .A2(new_n8185_), .A3(new_n8196_), .ZN(new_n8247_));
  NAND2_X1   g07966(.A1(new_n8246_), .A2(new_n8247_), .ZN(new_n8248_));
  AOI21_X1   g07967(.A1(new_n8248_), .A2(new_n7826_), .B(new_n7848_), .ZN(new_n8249_));
  OAI21_X1   g07968(.A1(new_n7826_), .A2(new_n8248_), .B(new_n7895_), .ZN(new_n8250_));
  NOR2_X1    g07969(.A1(new_n8250_), .A2(new_n8249_), .ZN(new_n8251_));
  OAI21_X1   g07970(.A1(new_n8189_), .A2(new_n8190_), .B(new_n8188_), .ZN(new_n8252_));
  AOI21_X1   g07971(.A1(new_n8252_), .A2(new_n7824_), .B(new_n7908_), .ZN(new_n8253_));
  AOI21_X1   g07972(.A1(new_n8165_), .A2(new_n8167_), .B(new_n7915_), .ZN(new_n8254_));
  OAI21_X1   g07973(.A1(new_n8254_), .A2(new_n7809_), .B(new_n7821_), .ZN(new_n8255_));
  AOI21_X1   g07974(.A1(new_n8150_), .A2(new_n8149_), .B(new_n8147_), .ZN(new_n8256_));
  AOI21_X1   g07975(.A1(new_n8152_), .A2(new_n7791_), .B(new_n7916_), .ZN(new_n8257_));
  NAND3_X1   g07976(.A1(new_n8148_), .A2(new_n8151_), .A3(new_n7790_), .ZN(new_n8258_));
  NAND2_X1   g07977(.A1(new_n7549_), .A2(new_n8258_), .ZN(new_n8259_));
  AOI21_X1   g07978(.A1(new_n8125_), .A2(new_n8119_), .B(new_n8133_), .ZN(new_n8260_));
  INV_X1     g07979(.I(new_n8260_), .ZN(new_n8261_));
  OAI21_X1   g07980(.A1(new_n8134_), .A2(new_n8130_), .B(new_n7923_), .ZN(new_n8262_));
  AOI21_X1   g07981(.A1(new_n8262_), .A2(new_n7785_), .B(new_n7783_), .ZN(new_n8263_));
  OAI21_X1   g07982(.A1(new_n8090_), .A2(new_n8089_), .B(new_n8087_), .ZN(new_n8264_));
  NAND3_X1   g07983(.A1(new_n8104_), .A2(new_n8109_), .A3(new_n8098_), .ZN(new_n8265_));
  AOI21_X1   g07984(.A1(new_n8264_), .A2(new_n8265_), .B(new_n8114_), .ZN(new_n8266_));
  INV_X1     g07985(.I(new_n8266_), .ZN(new_n8267_));
  NAND3_X1   g07986(.A1(new_n8264_), .A2(new_n8265_), .A3(new_n8114_), .ZN(new_n8268_));
  AOI21_X1   g07987(.A1(new_n8267_), .A2(new_n8268_), .B(new_n8094_), .ZN(new_n8269_));
  AOI21_X1   g07988(.A1(new_n8113_), .A2(new_n8117_), .B(new_n7925_), .ZN(new_n8270_));
  OAI21_X1   g07989(.A1(new_n8270_), .A2(new_n7771_), .B(new_n7918_), .ZN(new_n8271_));
  NAND2_X1   g07990(.A1(new_n8087_), .A2(new_n7929_), .ZN(new_n8272_));
  NOR2_X1    g07991(.A1(new_n8109_), .A2(new_n7929_), .ZN(new_n8273_));
  NAND3_X1   g07992(.A1(new_n8086_), .A2(new_n8079_), .A3(new_n7929_), .ZN(new_n8274_));
  INV_X1     g07993(.I(new_n8274_), .ZN(new_n8275_));
  OAI21_X1   g07994(.A1(new_n8273_), .A2(new_n8275_), .B(new_n8089_), .ZN(new_n8276_));
  AOI21_X1   g07995(.A1(new_n8276_), .A2(new_n8103_), .B(new_n7767_), .ZN(new_n8277_));
  OAI21_X1   g07996(.A1(new_n8084_), .A2(new_n8083_), .B(new_n8082_), .ZN(new_n8278_));
  AOI21_X1   g07997(.A1(new_n8278_), .A2(new_n7753_), .B(new_n7750_), .ZN(new_n8279_));
  OAI21_X1   g07998(.A1(new_n8055_), .A2(new_n8059_), .B(new_n7935_), .ZN(new_n8280_));
  AOI21_X1   g07999(.A1(new_n8280_), .A2(new_n7723_), .B(new_n7572_), .ZN(new_n8281_));
  NAND2_X1   g08000(.A1(new_n7938_), .A2(new_n8036_), .ZN(new_n8282_));
  NAND2_X1   g08001(.A1(new_n8037_), .A2(new_n8029_), .ZN(new_n8283_));
  AOI21_X1   g08002(.A1(new_n8283_), .A2(new_n8282_), .B(new_n8026_), .ZN(new_n8284_));
  OAI21_X1   g08003(.A1(new_n8048_), .A2(new_n7689_), .B(new_n8035_), .ZN(new_n8285_));
  NAND2_X1   g08004(.A1(new_n8048_), .A2(new_n7689_), .ZN(new_n8286_));
  NAND3_X1   g08005(.A1(new_n8285_), .A2(new_n7713_), .A3(new_n8286_), .ZN(new_n8287_));
  NAND3_X1   g08006(.A1(new_n8015_), .A2(new_n8016_), .A3(new_n8013_), .ZN(new_n8288_));
  OAI21_X1   g08007(.A1(new_n8014_), .A2(new_n8018_), .B(new_n7691_), .ZN(new_n8289_));
  NAND2_X1   g08008(.A1(new_n8289_), .A2(new_n7671_), .ZN(new_n8290_));
  NOR3_X1    g08009(.A1(new_n8014_), .A2(new_n8018_), .A3(new_n7691_), .ZN(new_n8291_));
  NOR2_X1    g08010(.A1(new_n8291_), .A2(new_n7583_), .ZN(new_n8292_));
  OAI21_X1   g08011(.A1(new_n8004_), .A2(new_n8005_), .B(new_n7647_), .ZN(new_n8293_));
  NAND2_X1   g08012(.A1(new_n8293_), .A2(new_n7652_), .ZN(new_n8294_));
  NOR3_X1    g08013(.A1(new_n8004_), .A2(new_n8005_), .A3(new_n7647_), .ZN(new_n8295_));
  NOR2_X1    g08014(.A1(new_n8295_), .A2(new_n7590_), .ZN(new_n8296_));
  XOR2_X1    g08015(.A1(new_n7961_), .A2(new_n6632_), .Z(new_n8297_));
  XOR2_X1    g08016(.A1(new_n7971_), .A2(new_n7957_), .Z(new_n8298_));
  NAND2_X1   g08017(.A1(new_n8298_), .A2(new_n8297_), .ZN(new_n8299_));
  INV_X1     g08018(.I(new_n8299_), .ZN(new_n8300_));
  AOI21_X1   g08019(.A1(new_n7983_), .A2(new_n7632_), .B(new_n7604_), .ZN(new_n8301_));
  OAI21_X1   g08020(.A1(new_n7983_), .A2(new_n7632_), .B(new_n7595_), .ZN(new_n8302_));
  AOI22_X1   g08021(.A1(new_n7607_), .A2(\b[2] ), .B1(\b[3] ), .B2(new_n7940_), .ZN(new_n8303_));
  OAI21_X1   g08022(.A1(new_n269_), .A2(new_n7947_), .B(new_n8303_), .ZN(new_n8304_));
  NOR2_X1    g08023(.A1(new_n403_), .A2(new_n7619_), .ZN(new_n8305_));
  AOI21_X1   g08024(.A1(new_n8304_), .A2(new_n8305_), .B(new_n7608_), .ZN(new_n8306_));
  XNOR2_X1   g08025(.A1(\a[44] ), .A2(\a[47] ), .ZN(new_n8307_));
  NOR3_X1    g08026(.A1(new_n7292_), .A2(new_n7606_), .A3(new_n8307_), .ZN(new_n8308_));
  NOR2_X1    g08027(.A1(new_n7612_), .A2(new_n7610_), .ZN(new_n8309_));
  OAI22_X1   g08028(.A1(new_n7619_), .A2(new_n280_), .B1(new_n298_), .B2(new_n8309_), .ZN(new_n8310_));
  AOI21_X1   g08029(.A1(\b[1] ), .A2(new_n8308_), .B(new_n8310_), .ZN(new_n8311_));
  NOR4_X1    g08030(.A1(new_n8311_), .A2(\a[47] ), .A3(new_n403_), .A4(new_n7619_), .ZN(new_n8312_));
  XNOR2_X1   g08031(.A1(\a[47] ), .A2(\a[48] ), .ZN(new_n8313_));
  NOR2_X1    g08032(.A1(new_n8313_), .A2(new_n258_), .ZN(new_n8314_));
  OAI21_X1   g08033(.A1(new_n8312_), .A2(new_n8306_), .B(new_n8314_), .ZN(new_n8315_));
  NOR2_X1    g08034(.A1(new_n8315_), .A2(new_n7971_), .ZN(new_n8316_));
  INV_X1     g08035(.I(new_n8306_), .ZN(new_n8317_));
  NAND3_X1   g08036(.A1(new_n8304_), .A2(new_n8305_), .A3(new_n7608_), .ZN(new_n8318_));
  INV_X1     g08037(.I(new_n8314_), .ZN(new_n8319_));
  AOI21_X1   g08038(.A1(new_n8317_), .A2(new_n8318_), .B(new_n8319_), .ZN(new_n8320_));
  NOR2_X1    g08039(.A1(new_n8320_), .A2(new_n7956_), .ZN(new_n8321_));
  OAI21_X1   g08040(.A1(new_n8321_), .A2(new_n8316_), .B(new_n7963_), .ZN(new_n8322_));
  NAND2_X1   g08041(.A1(new_n8320_), .A2(new_n7956_), .ZN(new_n8323_));
  NAND2_X1   g08042(.A1(new_n8315_), .A2(new_n7971_), .ZN(new_n8324_));
  NAND3_X1   g08043(.A1(new_n8323_), .A2(new_n7957_), .A3(new_n8324_), .ZN(new_n8325_));
  OAI22_X1   g08044(.A1(new_n6644_), .A2(new_n419_), .B1(new_n420_), .B2(new_n6647_), .ZN(new_n8326_));
  OAI21_X1   g08045(.A1(new_n325_), .A2(new_n7284_), .B(new_n8326_), .ZN(new_n8327_));
  AOI21_X1   g08046(.A1(new_n8327_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n8328_));
  XOR2_X1    g08047(.A1(new_n425_), .A2(new_n8328_), .Z(new_n8329_));
  AOI21_X1   g08048(.A1(new_n8322_), .A2(new_n8325_), .B(new_n8329_), .ZN(new_n8330_));
  OAI21_X1   g08049(.A1(new_n8301_), .A2(new_n8302_), .B(new_n8330_), .ZN(new_n8331_));
  NOR2_X1    g08050(.A1(new_n8301_), .A2(new_n8302_), .ZN(new_n8332_));
  INV_X1     g08051(.I(new_n8330_), .ZN(new_n8333_));
  NAND2_X1   g08052(.A1(new_n8332_), .A2(new_n8333_), .ZN(new_n8334_));
  AOI21_X1   g08053(.A1(new_n8334_), .A2(new_n8331_), .B(new_n8300_), .ZN(new_n8335_));
  INV_X1     g08054(.I(new_n8331_), .ZN(new_n8336_));
  NOR3_X1    g08055(.A1(new_n8301_), .A2(new_n8302_), .A3(new_n8330_), .ZN(new_n8337_));
  NOR3_X1    g08056(.A1(new_n8336_), .A2(new_n8299_), .A3(new_n8337_), .ZN(new_n8338_));
  OAI22_X1   g08057(.A1(new_n5993_), .A2(new_n515_), .B1(new_n565_), .B2(new_n5991_), .ZN(new_n8339_));
  OAI21_X1   g08058(.A1(new_n472_), .A2(new_n5997_), .B(new_n8339_), .ZN(new_n8340_));
  AOI21_X1   g08059(.A1(new_n8340_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n8341_));
  XOR2_X1    g08060(.A1(new_n759_), .A2(new_n8341_), .Z(new_n8342_));
  INV_X1     g08061(.I(new_n8342_), .ZN(new_n8343_));
  OAI21_X1   g08062(.A1(new_n8338_), .A2(new_n8335_), .B(new_n8343_), .ZN(new_n8344_));
  AOI21_X1   g08063(.A1(new_n8296_), .A2(new_n8294_), .B(new_n8344_), .ZN(new_n8345_));
  AOI21_X1   g08064(.A1(new_n7999_), .A2(new_n7647_), .B(new_n7653_), .ZN(new_n8346_));
  AOI21_X1   g08065(.A1(new_n7633_), .A2(new_n7638_), .B(new_n7642_), .ZN(new_n8347_));
  INV_X1     g08066(.I(new_n7645_), .ZN(new_n8348_));
  NOR2_X1    g08067(.A1(new_n8348_), .A2(new_n7595_), .ZN(new_n8349_));
  NOR2_X1    g08068(.A1(new_n8347_), .A2(new_n8349_), .ZN(new_n8350_));
  NAND3_X1   g08069(.A1(new_n7998_), .A2(new_n7995_), .A3(new_n8350_), .ZN(new_n8351_));
  NAND2_X1   g08070(.A1(new_n8351_), .A2(new_n7661_), .ZN(new_n8352_));
  OAI21_X1   g08071(.A1(new_n8336_), .A2(new_n8337_), .B(new_n8299_), .ZN(new_n8353_));
  NAND3_X1   g08072(.A1(new_n8334_), .A2(new_n8300_), .A3(new_n8331_), .ZN(new_n8354_));
  AOI21_X1   g08073(.A1(new_n8353_), .A2(new_n8354_), .B(new_n8342_), .ZN(new_n8355_));
  NOR3_X1    g08074(.A1(new_n8346_), .A2(new_n8352_), .A3(new_n8355_), .ZN(new_n8356_));
  OAI21_X1   g08075(.A1(new_n8345_), .A2(new_n8356_), .B(new_n7998_), .ZN(new_n8357_));
  OAI21_X1   g08076(.A1(new_n8346_), .A2(new_n8352_), .B(new_n8355_), .ZN(new_n8358_));
  NAND3_X1   g08077(.A1(new_n8294_), .A2(new_n8296_), .A3(new_n8344_), .ZN(new_n8359_));
  NAND3_X1   g08078(.A1(new_n8359_), .A2(new_n8358_), .A3(new_n8005_), .ZN(new_n8360_));
  OAI22_X1   g08079(.A1(new_n5420_), .A2(new_n706_), .B1(new_n780_), .B2(new_n5107_), .ZN(new_n8361_));
  OAI21_X1   g08080(.A1(new_n656_), .A2(new_n5112_), .B(new_n8361_), .ZN(new_n8362_));
  AOI21_X1   g08081(.A1(new_n8362_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n8363_));
  XOR2_X1    g08082(.A1(new_n785_), .A2(new_n8363_), .Z(new_n8364_));
  AOI21_X1   g08083(.A1(new_n8357_), .A2(new_n8360_), .B(new_n8364_), .ZN(new_n8365_));
  INV_X1     g08084(.I(new_n8365_), .ZN(new_n8366_));
  AOI21_X1   g08085(.A1(new_n8292_), .A2(new_n8290_), .B(new_n8366_), .ZN(new_n8367_));
  AOI21_X1   g08086(.A1(new_n8036_), .A2(new_n7691_), .B(new_n7672_), .ZN(new_n8368_));
  NAND3_X1   g08087(.A1(new_n8025_), .A2(new_n8024_), .A3(new_n7667_), .ZN(new_n8369_));
  NAND2_X1   g08088(.A1(new_n8369_), .A2(new_n7681_), .ZN(new_n8370_));
  NOR3_X1    g08089(.A1(new_n8368_), .A2(new_n8370_), .A3(new_n8365_), .ZN(new_n8371_));
  OAI21_X1   g08090(.A1(new_n8367_), .A2(new_n8371_), .B(new_n8288_), .ZN(new_n8372_));
  INV_X1     g08091(.I(new_n8288_), .ZN(new_n8373_));
  OAI21_X1   g08092(.A1(new_n8368_), .A2(new_n8370_), .B(new_n8365_), .ZN(new_n8374_));
  NAND3_X1   g08093(.A1(new_n8292_), .A2(new_n8290_), .A3(new_n8366_), .ZN(new_n8375_));
  NAND3_X1   g08094(.A1(new_n8375_), .A2(new_n8374_), .A3(new_n8373_), .ZN(new_n8376_));
  OAI22_X1   g08095(.A1(new_n4072_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n4067_), .ZN(new_n8377_));
  OAI21_X1   g08096(.A1(new_n861_), .A2(new_n4318_), .B(new_n8377_), .ZN(new_n8378_));
  AOI21_X1   g08097(.A1(new_n8378_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n8379_));
  XOR2_X1    g08098(.A1(new_n1024_), .A2(new_n8379_), .Z(new_n8380_));
  AOI21_X1   g08099(.A1(new_n8372_), .A2(new_n8376_), .B(new_n8380_), .ZN(new_n8381_));
  NAND2_X1   g08100(.A1(new_n8287_), .A2(new_n8381_), .ZN(new_n8382_));
  AOI21_X1   g08101(.A1(new_n8033_), .A2(new_n7695_), .B(new_n7936_), .ZN(new_n8383_));
  NOR2_X1    g08102(.A1(new_n8033_), .A2(new_n7695_), .ZN(new_n8384_));
  NOR3_X1    g08103(.A1(new_n8383_), .A2(new_n7577_), .A3(new_n8384_), .ZN(new_n8385_));
  AOI21_X1   g08104(.A1(new_n8375_), .A2(new_n8374_), .B(new_n8373_), .ZN(new_n8386_));
  NOR3_X1    g08105(.A1(new_n8367_), .A2(new_n8371_), .A3(new_n8288_), .ZN(new_n8387_));
  INV_X1     g08106(.I(new_n8380_), .ZN(new_n8388_));
  OAI21_X1   g08107(.A1(new_n8387_), .A2(new_n8386_), .B(new_n8388_), .ZN(new_n8389_));
  NAND2_X1   g08108(.A1(new_n8385_), .A2(new_n8389_), .ZN(new_n8390_));
  AOI21_X1   g08109(.A1(new_n8390_), .A2(new_n8382_), .B(new_n8284_), .ZN(new_n8391_));
  INV_X1     g08110(.I(new_n8284_), .ZN(new_n8392_));
  NOR2_X1    g08111(.A1(new_n8385_), .A2(new_n8389_), .ZN(new_n8393_));
  NOR2_X1    g08112(.A1(new_n8287_), .A2(new_n8381_), .ZN(new_n8394_));
  NOR3_X1    g08113(.A1(new_n8393_), .A2(new_n8394_), .A3(new_n8392_), .ZN(new_n8395_));
  OAI22_X1   g08114(.A1(new_n1189_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1294_), .ZN(new_n8396_));
  OAI21_X1   g08115(.A1(new_n1109_), .A2(new_n3569_), .B(new_n8396_), .ZN(new_n8397_));
  AOI21_X1   g08116(.A1(new_n8397_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n8398_));
  XOR2_X1    g08117(.A1(new_n1299_), .A2(new_n8398_), .Z(new_n8399_));
  INV_X1     g08118(.I(new_n8399_), .ZN(new_n8400_));
  OAI21_X1   g08119(.A1(new_n8391_), .A2(new_n8395_), .B(new_n8400_), .ZN(new_n8401_));
  NOR2_X1    g08120(.A1(new_n8281_), .A2(new_n8401_), .ZN(new_n8402_));
  AOI21_X1   g08121(.A1(new_n8066_), .A2(new_n8065_), .B(new_n8064_), .ZN(new_n8403_));
  OAI21_X1   g08122(.A1(new_n8403_), .A2(new_n7741_), .B(new_n7728_), .ZN(new_n8404_));
  OAI21_X1   g08123(.A1(new_n8393_), .A2(new_n8394_), .B(new_n8392_), .ZN(new_n8405_));
  NAND3_X1   g08124(.A1(new_n8390_), .A2(new_n8382_), .A3(new_n8284_), .ZN(new_n8406_));
  AOI21_X1   g08125(.A1(new_n8405_), .A2(new_n8406_), .B(new_n8399_), .ZN(new_n8407_));
  NOR2_X1    g08126(.A1(new_n8404_), .A2(new_n8407_), .ZN(new_n8408_));
  OAI21_X1   g08127(.A1(new_n8408_), .A2(new_n8402_), .B(new_n8066_), .ZN(new_n8409_));
  NAND2_X1   g08128(.A1(new_n8404_), .A2(new_n8407_), .ZN(new_n8410_));
  NAND2_X1   g08129(.A1(new_n8281_), .A2(new_n8401_), .ZN(new_n8411_));
  NAND3_X1   g08130(.A1(new_n8410_), .A2(new_n8411_), .A3(new_n8059_), .ZN(new_n8412_));
  NAND2_X1   g08131(.A1(new_n8409_), .A2(new_n8412_), .ZN(new_n8413_));
  OAI22_X1   g08132(.A1(new_n1525_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1634_), .ZN(new_n8414_));
  OAI21_X1   g08133(.A1(new_n1518_), .A2(new_n2884_), .B(new_n8414_), .ZN(new_n8415_));
  AOI21_X1   g08134(.A1(new_n8415_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n8416_));
  XNOR2_X1   g08135(.A1(new_n1638_), .A2(new_n8416_), .ZN(new_n8417_));
  INV_X1     g08136(.I(new_n8417_), .ZN(new_n8418_));
  NAND2_X1   g08137(.A1(new_n8413_), .A2(new_n8418_), .ZN(new_n8419_));
  NOR2_X1    g08138(.A1(new_n8419_), .A2(new_n8279_), .ZN(new_n8420_));
  AOI21_X1   g08139(.A1(new_n8074_), .A2(new_n8077_), .B(new_n7932_), .ZN(new_n8421_));
  OAI21_X1   g08140(.A1(new_n8421_), .A2(new_n7751_), .B(new_n7568_), .ZN(new_n8422_));
  AOI21_X1   g08141(.A1(new_n8413_), .A2(new_n8418_), .B(new_n8422_), .ZN(new_n8423_));
  OAI21_X1   g08142(.A1(new_n8420_), .A2(new_n8423_), .B(new_n8077_), .ZN(new_n8424_));
  NAND3_X1   g08143(.A1(new_n8422_), .A2(new_n8413_), .A3(new_n8418_), .ZN(new_n8425_));
  NAND2_X1   g08144(.A1(new_n8419_), .A2(new_n8279_), .ZN(new_n8426_));
  NAND3_X1   g08145(.A1(new_n8426_), .A2(new_n8084_), .A3(new_n8425_), .ZN(new_n8427_));
  OAI22_X1   g08146(.A1(new_n2171_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n2166_), .ZN(new_n8428_));
  OAI21_X1   g08147(.A1(new_n1803_), .A2(new_n2322_), .B(new_n8428_), .ZN(new_n8429_));
  AOI21_X1   g08148(.A1(new_n8429_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n8430_));
  XOR2_X1    g08149(.A1(new_n2106_), .A2(new_n8430_), .Z(new_n8431_));
  AOI21_X1   g08150(.A1(new_n8424_), .A2(new_n8427_), .B(new_n8431_), .ZN(new_n8432_));
  INV_X1     g08151(.I(new_n8432_), .ZN(new_n8433_));
  NOR2_X1    g08152(.A1(new_n8433_), .A2(new_n8277_), .ZN(new_n8434_));
  NAND2_X1   g08153(.A1(new_n8087_), .A2(new_n8114_), .ZN(new_n8435_));
  AOI21_X1   g08154(.A1(new_n8435_), .A2(new_n8274_), .B(new_n8098_), .ZN(new_n8436_));
  OAI21_X1   g08155(.A1(new_n8436_), .A2(new_n7756_), .B(new_n7564_), .ZN(new_n8437_));
  NOR2_X1    g08156(.A1(new_n8437_), .A2(new_n8432_), .ZN(new_n8438_));
  OAI21_X1   g08157(.A1(new_n8434_), .A2(new_n8438_), .B(new_n8272_), .ZN(new_n8439_));
  INV_X1     g08158(.I(new_n8272_), .ZN(new_n8440_));
  NAND2_X1   g08159(.A1(new_n8437_), .A2(new_n8432_), .ZN(new_n8441_));
  NAND2_X1   g08160(.A1(new_n8433_), .A2(new_n8277_), .ZN(new_n8442_));
  NAND3_X1   g08161(.A1(new_n8442_), .A2(new_n8441_), .A3(new_n8440_), .ZN(new_n8443_));
  OAI22_X1   g08162(.A1(new_n1712_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n1707_), .ZN(new_n8444_));
  OAI21_X1   g08163(.A1(new_n2281_), .A2(new_n1850_), .B(new_n8444_), .ZN(new_n8445_));
  AOI21_X1   g08164(.A1(new_n8445_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n8446_));
  XNOR2_X1   g08165(.A1(new_n2647_), .A2(new_n8446_), .ZN(new_n8447_));
  AOI21_X1   g08166(.A1(new_n8439_), .A2(new_n8443_), .B(new_n8447_), .ZN(new_n8448_));
  NAND2_X1   g08167(.A1(new_n8271_), .A2(new_n8448_), .ZN(new_n8449_));
  OAI21_X1   g08168(.A1(new_n8123_), .A2(new_n8122_), .B(new_n8121_), .ZN(new_n8450_));
  AOI21_X1   g08169(.A1(new_n8450_), .A2(new_n7919_), .B(new_n7559_), .ZN(new_n8451_));
  AOI21_X1   g08170(.A1(new_n8442_), .A2(new_n8441_), .B(new_n8440_), .ZN(new_n8452_));
  NOR3_X1    g08171(.A1(new_n8434_), .A2(new_n8438_), .A3(new_n8272_), .ZN(new_n8453_));
  INV_X1     g08172(.I(new_n8447_), .ZN(new_n8454_));
  OAI21_X1   g08173(.A1(new_n8453_), .A2(new_n8452_), .B(new_n8454_), .ZN(new_n8455_));
  NAND2_X1   g08174(.A1(new_n8451_), .A2(new_n8455_), .ZN(new_n8456_));
  AOI21_X1   g08175(.A1(new_n8456_), .A2(new_n8449_), .B(new_n8269_), .ZN(new_n8457_));
  INV_X1     g08176(.I(new_n8269_), .ZN(new_n8458_));
  NOR2_X1    g08177(.A1(new_n8451_), .A2(new_n8455_), .ZN(new_n8459_));
  NOR2_X1    g08178(.A1(new_n8271_), .A2(new_n8448_), .ZN(new_n8460_));
  NOR3_X1    g08179(.A1(new_n8459_), .A2(new_n8460_), .A3(new_n8458_), .ZN(new_n8461_));
  OAI22_X1   g08180(.A1(new_n1347_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n1344_), .ZN(new_n8462_));
  OAI21_X1   g08181(.A1(new_n2842_), .A2(new_n1457_), .B(new_n8462_), .ZN(new_n8463_));
  AOI21_X1   g08182(.A1(new_n8463_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n8464_));
  XNOR2_X1   g08183(.A1(new_n3264_), .A2(new_n8464_), .ZN(new_n8465_));
  INV_X1     g08184(.I(new_n8465_), .ZN(new_n8466_));
  OAI21_X1   g08185(.A1(new_n8457_), .A2(new_n8461_), .B(new_n8466_), .ZN(new_n8467_));
  NOR2_X1    g08186(.A1(new_n8263_), .A2(new_n8467_), .ZN(new_n8468_));
  AOI21_X1   g08187(.A1(new_n8139_), .A2(new_n8140_), .B(new_n8138_), .ZN(new_n8469_));
  OAI21_X1   g08188(.A1(new_n8469_), .A2(new_n7780_), .B(new_n7554_), .ZN(new_n8470_));
  OAI21_X1   g08189(.A1(new_n8459_), .A2(new_n8460_), .B(new_n8458_), .ZN(new_n8471_));
  NAND3_X1   g08190(.A1(new_n8456_), .A2(new_n8449_), .A3(new_n8269_), .ZN(new_n8472_));
  AOI21_X1   g08191(.A1(new_n8471_), .A2(new_n8472_), .B(new_n8465_), .ZN(new_n8473_));
  NOR2_X1    g08192(.A1(new_n8470_), .A2(new_n8473_), .ZN(new_n8474_));
  OAI21_X1   g08193(.A1(new_n8468_), .A2(new_n8474_), .B(new_n8261_), .ZN(new_n8475_));
  NAND2_X1   g08194(.A1(new_n8470_), .A2(new_n8473_), .ZN(new_n8476_));
  NAND2_X1   g08195(.A1(new_n8263_), .A2(new_n8467_), .ZN(new_n8477_));
  NAND3_X1   g08196(.A1(new_n8477_), .A2(new_n8476_), .A3(new_n8260_), .ZN(new_n8478_));
  OAI22_X1   g08197(.A1(new_n1055_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n1061_), .ZN(new_n8479_));
  OAI21_X1   g08198(.A1(new_n3709_), .A2(new_n1332_), .B(new_n8479_), .ZN(new_n8480_));
  AOI21_X1   g08199(.A1(new_n8480_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n8481_));
  XNOR2_X1   g08200(.A1(new_n3993_), .A2(new_n8481_), .ZN(new_n8482_));
  AOI21_X1   g08201(.A1(new_n8475_), .A2(new_n8478_), .B(new_n8482_), .ZN(new_n8483_));
  OAI21_X1   g08202(.A1(new_n8257_), .A2(new_n8259_), .B(new_n8483_), .ZN(new_n8484_));
  INV_X1     g08203(.I(new_n7916_), .ZN(new_n8485_));
  OAI21_X1   g08204(.A1(new_n8155_), .A2(new_n8154_), .B(new_n7791_), .ZN(new_n8486_));
  NAND2_X1   g08205(.A1(new_n8486_), .A2(new_n8485_), .ZN(new_n8487_));
  AOI21_X1   g08206(.A1(new_n8477_), .A2(new_n8476_), .B(new_n8260_), .ZN(new_n8488_));
  NOR3_X1    g08207(.A1(new_n8468_), .A2(new_n8474_), .A3(new_n8261_), .ZN(new_n8489_));
  INV_X1     g08208(.I(new_n8482_), .ZN(new_n8490_));
  OAI21_X1   g08209(.A1(new_n8488_), .A2(new_n8489_), .B(new_n8490_), .ZN(new_n8491_));
  NAND4_X1   g08210(.A1(new_n8491_), .A2(new_n8487_), .A3(new_n7549_), .A4(new_n8258_), .ZN(new_n8492_));
  AOI21_X1   g08211(.A1(new_n8484_), .A2(new_n8492_), .B(new_n8256_), .ZN(new_n8493_));
  INV_X1     g08212(.I(new_n8256_), .ZN(new_n8494_));
  NOR2_X1    g08213(.A1(new_n8259_), .A2(new_n8257_), .ZN(new_n8495_));
  NOR2_X1    g08214(.A1(new_n8495_), .A2(new_n8491_), .ZN(new_n8496_));
  NOR3_X1    g08215(.A1(new_n8483_), .A2(new_n8259_), .A3(new_n8257_), .ZN(new_n8497_));
  NOR3_X1    g08216(.A1(new_n8496_), .A2(new_n8494_), .A3(new_n8497_), .ZN(new_n8498_));
  OAI22_X1   g08217(.A1(new_n970_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n820_), .ZN(new_n8499_));
  OAI21_X1   g08218(.A1(new_n4253_), .A2(new_n894_), .B(new_n8499_), .ZN(new_n8500_));
  AOI21_X1   g08219(.A1(new_n8500_), .A2(new_n827_), .B(new_n970_), .ZN(new_n8501_));
  XNOR2_X1   g08220(.A1(new_n4778_), .A2(new_n8501_), .ZN(new_n8502_));
  INV_X1     g08221(.I(new_n8502_), .ZN(new_n8503_));
  OAI21_X1   g08222(.A1(new_n8498_), .A2(new_n8493_), .B(new_n8503_), .ZN(new_n8504_));
  INV_X1     g08223(.I(new_n8504_), .ZN(new_n8505_));
  NAND2_X1   g08224(.A1(new_n8255_), .A2(new_n8505_), .ZN(new_n8506_));
  OAI21_X1   g08225(.A1(new_n8172_), .A2(new_n8171_), .B(new_n8170_), .ZN(new_n8507_));
  AOI21_X1   g08226(.A1(new_n8507_), .A2(new_n7816_), .B(new_n7545_), .ZN(new_n8508_));
  NAND2_X1   g08227(.A1(new_n8508_), .A2(new_n8504_), .ZN(new_n8509_));
  AOI21_X1   g08228(.A1(new_n8509_), .A2(new_n8506_), .B(new_n8172_), .ZN(new_n8510_));
  NOR2_X1    g08229(.A1(new_n8508_), .A2(new_n8504_), .ZN(new_n8511_));
  NOR2_X1    g08230(.A1(new_n8255_), .A2(new_n8505_), .ZN(new_n8512_));
  NOR3_X1    g08231(.A1(new_n8511_), .A2(new_n8512_), .A3(new_n8167_), .ZN(new_n8513_));
  OAI22_X1   g08232(.A1(new_n607_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n610_), .ZN(new_n8514_));
  OAI21_X1   g08233(.A1(new_n5068_), .A2(new_n684_), .B(new_n8514_), .ZN(new_n8515_));
  AOI21_X1   g08234(.A1(new_n8515_), .A2(new_n612_), .B(new_n607_), .ZN(new_n8516_));
  XNOR2_X1   g08235(.A1(new_n5600_), .A2(new_n8516_), .ZN(new_n8517_));
  INV_X1     g08236(.I(new_n8517_), .ZN(new_n8518_));
  OAI21_X1   g08237(.A1(new_n8510_), .A2(new_n8513_), .B(new_n8518_), .ZN(new_n8519_));
  NOR2_X1    g08238(.A1(new_n8253_), .A2(new_n8519_), .ZN(new_n8520_));
  AOI21_X1   g08239(.A1(new_n8183_), .A2(new_n8180_), .B(new_n7912_), .ZN(new_n8521_));
  OAI21_X1   g08240(.A1(new_n8521_), .A2(new_n7909_), .B(new_n7540_), .ZN(new_n8522_));
  OAI21_X1   g08241(.A1(new_n8511_), .A2(new_n8512_), .B(new_n8167_), .ZN(new_n8523_));
  NAND3_X1   g08242(.A1(new_n8509_), .A2(new_n8506_), .A3(new_n8172_), .ZN(new_n8524_));
  AOI21_X1   g08243(.A1(new_n8523_), .A2(new_n8524_), .B(new_n8517_), .ZN(new_n8525_));
  NOR2_X1    g08244(.A1(new_n8522_), .A2(new_n8525_), .ZN(new_n8526_));
  OAI21_X1   g08245(.A1(new_n8520_), .A2(new_n8526_), .B(new_n8183_), .ZN(new_n8527_));
  NAND2_X1   g08246(.A1(new_n8522_), .A2(new_n8525_), .ZN(new_n8528_));
  NAND2_X1   g08247(.A1(new_n8253_), .A2(new_n8519_), .ZN(new_n8529_));
  NAND3_X1   g08248(.A1(new_n8529_), .A2(new_n8528_), .A3(new_n8190_), .ZN(new_n8530_));
  NAND2_X1   g08249(.A1(new_n8527_), .A2(new_n8530_), .ZN(new_n8531_));
  OAI22_X1   g08250(.A1(new_n448_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n450_), .ZN(new_n8532_));
  OAI21_X1   g08251(.A1(new_n5921_), .A2(new_n496_), .B(new_n8532_), .ZN(new_n8533_));
  AOI21_X1   g08252(.A1(new_n8533_), .A2(new_n452_), .B(new_n448_), .ZN(new_n8534_));
  XOR2_X1    g08253(.A1(new_n6543_), .A2(new_n8534_), .Z(new_n8535_));
  INV_X1     g08254(.I(new_n8535_), .ZN(new_n8536_));
  NAND2_X1   g08255(.A1(new_n8531_), .A2(new_n8536_), .ZN(new_n8537_));
  NOR2_X1    g08256(.A1(new_n8251_), .A2(new_n8537_), .ZN(new_n8538_));
  OAI21_X1   g08257(.A1(new_n8207_), .A2(new_n7825_), .B(new_n7536_), .ZN(new_n8539_));
  AOI21_X1   g08258(.A1(new_n7825_), .A2(new_n8207_), .B(new_n7902_), .ZN(new_n8540_));
  NAND2_X1   g08259(.A1(new_n8540_), .A2(new_n8539_), .ZN(new_n8541_));
  AOI21_X1   g08260(.A1(new_n8531_), .A2(new_n8536_), .B(new_n8541_), .ZN(new_n8542_));
  OAI21_X1   g08261(.A1(new_n8542_), .A2(new_n8538_), .B(new_n8200_), .ZN(new_n8543_));
  NAND3_X1   g08262(.A1(new_n8541_), .A2(new_n8531_), .A3(new_n8536_), .ZN(new_n8544_));
  NAND2_X1   g08263(.A1(new_n8251_), .A2(new_n8537_), .ZN(new_n8545_));
  NAND3_X1   g08264(.A1(new_n8544_), .A2(new_n8545_), .A3(new_n8199_), .ZN(new_n8546_));
  NAND2_X1   g08265(.A1(new_n8543_), .A2(new_n8546_), .ZN(new_n8547_));
  OAI22_X1   g08266(.A1(new_n7198_), .A2(new_n341_), .B1(new_n404_), .B2(new_n7864_), .ZN(new_n8548_));
  OAI21_X1   g08267(.A1(new_n6847_), .A2(new_n366_), .B(new_n8548_), .ZN(new_n8549_));
  AOI21_X1   g08268(.A1(new_n8549_), .A2(new_n334_), .B(new_n341_), .ZN(new_n8550_));
  XOR2_X1    g08269(.A1(new_n7516_), .A2(new_n8550_), .Z(new_n8551_));
  INV_X1     g08270(.I(new_n8551_), .ZN(new_n8552_));
  XOR2_X1    g08271(.A1(new_n8547_), .A2(new_n8552_), .Z(new_n8553_));
  NOR2_X1    g08272(.A1(\b[46] ), .A2(\b[47] ), .ZN(new_n8554_));
  AOI21_X1   g08273(.A1(new_n7868_), .A2(new_n8554_), .B(new_n7864_), .ZN(new_n8555_));
  NOR2_X1    g08274(.A1(new_n7870_), .A2(new_n8218_), .ZN(new_n8556_));
  INV_X1     g08275(.I(new_n8556_), .ZN(new_n8557_));
  NOR2_X1    g08276(.A1(new_n7868_), .A2(new_n8557_), .ZN(new_n8558_));
  NOR2_X1    g08277(.A1(new_n8555_), .A2(new_n8558_), .ZN(new_n8559_));
  INV_X1     g08278(.I(new_n8559_), .ZN(new_n8560_));
  XNOR2_X1   g08279(.A1(\b[47] ), .A2(\b[48] ), .ZN(new_n8561_));
  INV_X1     g08280(.I(new_n8561_), .ZN(new_n8562_));
  INV_X1     g08281(.I(\b[48] ), .ZN(new_n8563_));
  NOR2_X1    g08282(.A1(new_n8218_), .A2(new_n8563_), .ZN(new_n8564_));
  INV_X1     g08283(.I(new_n8564_), .ZN(new_n8565_));
  NAND2_X1   g08284(.A1(new_n8218_), .A2(new_n8563_), .ZN(new_n8566_));
  AOI21_X1   g08285(.A1(new_n8565_), .A2(new_n8566_), .B(new_n8560_), .ZN(new_n8567_));
  AOI21_X1   g08286(.A1(new_n8560_), .A2(new_n8562_), .B(new_n8567_), .ZN(new_n8568_));
  OAI22_X1   g08287(.A1(new_n330_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n263_), .ZN(new_n8569_));
  OAI21_X1   g08288(.A1(new_n7870_), .A2(new_n289_), .B(new_n8569_), .ZN(new_n8570_));
  AOI21_X1   g08289(.A1(new_n8570_), .A2(new_n260_), .B(new_n426_), .ZN(new_n8571_));
  XOR2_X1    g08290(.A1(new_n8568_), .A2(new_n8571_), .Z(new_n8572_));
  XOR2_X1    g08291(.A1(new_n8553_), .A2(new_n8572_), .Z(new_n8573_));
  NAND2_X1   g08292(.A1(new_n8573_), .A2(new_n8245_), .ZN(new_n8574_));
  XOR2_X1    g08293(.A1(new_n8553_), .A2(new_n8572_), .Z(new_n8575_));
  OAI21_X1   g08294(.A1(new_n8245_), .A2(new_n8575_), .B(new_n8574_), .ZN(new_n8576_));
  NOR2_X1    g08295(.A1(new_n8576_), .A2(new_n8233_), .ZN(new_n8577_));
  NOR2_X1    g08296(.A1(new_n8230_), .A2(new_n8577_), .ZN(new_n8578_));
  XNOR2_X1   g08297(.A1(new_n8578_), .A2(new_n8226_), .ZN(\f[48] ));
  OAI22_X1   g08298(.A1(new_n7864_), .A2(new_n341_), .B1(new_n404_), .B2(new_n7870_), .ZN(new_n8580_));
  OAI21_X1   g08299(.A1(new_n7198_), .A2(new_n366_), .B(new_n8580_), .ZN(new_n8581_));
  AOI21_X1   g08300(.A1(new_n8581_), .A2(new_n334_), .B(new_n341_), .ZN(new_n8582_));
  XNOR2_X1   g08301(.A1(new_n7874_), .A2(new_n8582_), .ZN(new_n8583_));
  INV_X1     g08302(.I(new_n8583_), .ZN(new_n8584_));
  NOR2_X1    g08303(.A1(new_n8453_), .A2(new_n8452_), .ZN(new_n8585_));
  NAND2_X1   g08304(.A1(new_n8439_), .A2(new_n8443_), .ZN(new_n8586_));
  OAI21_X1   g08305(.A1(new_n8586_), .A2(new_n8269_), .B(new_n8454_), .ZN(new_n8587_));
  OAI22_X1   g08306(.A1(new_n8587_), .A2(new_n8271_), .B1(new_n8458_), .B2(new_n8585_), .ZN(new_n8588_));
  AOI21_X1   g08307(.A1(new_n8357_), .A2(new_n8360_), .B(new_n8288_), .ZN(new_n8589_));
  INV_X1     g08308(.I(new_n8364_), .ZN(new_n8590_));
  NAND3_X1   g08309(.A1(new_n8357_), .A2(new_n8360_), .A3(new_n8288_), .ZN(new_n8591_));
  NAND2_X1   g08310(.A1(new_n8591_), .A2(new_n8590_), .ZN(new_n8592_));
  NOR3_X1    g08311(.A1(new_n8592_), .A2(new_n8368_), .A3(new_n8370_), .ZN(new_n8593_));
  NAND2_X1   g08312(.A1(new_n8296_), .A2(new_n8294_), .ZN(new_n8594_));
  AOI21_X1   g08313(.A1(new_n8353_), .A2(new_n8354_), .B(new_n7998_), .ZN(new_n8595_));
  INV_X1     g08314(.I(new_n8595_), .ZN(new_n8596_));
  NAND3_X1   g08315(.A1(new_n8353_), .A2(new_n8354_), .A3(new_n7998_), .ZN(new_n8597_));
  NAND2_X1   g08316(.A1(new_n8597_), .A2(new_n8343_), .ZN(new_n8598_));
  OAI21_X1   g08317(.A1(new_n8594_), .A2(new_n8598_), .B(new_n8596_), .ZN(new_n8599_));
  INV_X1     g08318(.I(new_n8332_), .ZN(new_n8600_));
  NAND2_X1   g08319(.A1(new_n8322_), .A2(new_n8325_), .ZN(new_n8601_));
  NAND2_X1   g08320(.A1(new_n8601_), .A2(new_n8300_), .ZN(new_n8602_));
  INV_X1     g08321(.I(new_n8329_), .ZN(new_n8603_));
  NAND3_X1   g08322(.A1(new_n8322_), .A2(new_n8325_), .A3(new_n8299_), .ZN(new_n8604_));
  NAND2_X1   g08323(.A1(new_n8604_), .A2(new_n8603_), .ZN(new_n8605_));
  OAI21_X1   g08324(.A1(new_n8600_), .A2(new_n8605_), .B(new_n8602_), .ZN(new_n8606_));
  NOR2_X1    g08325(.A1(new_n8312_), .A2(new_n8306_), .ZN(new_n8607_));
  NOR2_X1    g08326(.A1(new_n8607_), .A2(new_n7956_), .ZN(new_n8608_));
  INV_X1     g08327(.I(new_n8608_), .ZN(new_n8609_));
  NAND2_X1   g08328(.A1(new_n8607_), .A2(new_n7956_), .ZN(new_n8610_));
  NOR2_X1    g08329(.A1(new_n7963_), .A2(new_n8319_), .ZN(new_n8611_));
  NAND2_X1   g08330(.A1(new_n8610_), .A2(new_n8611_), .ZN(new_n8612_));
  NAND2_X1   g08331(.A1(new_n8612_), .A2(new_n8609_), .ZN(new_n8613_));
  AOI21_X1   g08332(.A1(new_n7620_), .A2(new_n7621_), .B(new_n325_), .ZN(new_n8614_));
  AOI21_X1   g08333(.A1(new_n7607_), .A2(\b[3] ), .B(new_n8614_), .ZN(new_n8615_));
  NAND4_X1   g08334(.A1(new_n7945_), .A2(new_n7615_), .A3(new_n7946_), .A4(\b[2] ), .ZN(new_n8616_));
  INV_X1     g08335(.I(new_n8616_), .ZN(new_n8617_));
  OAI21_X1   g08336(.A1(new_n8615_), .A2(new_n8617_), .B(new_n7608_), .ZN(new_n8618_));
  NAND3_X1   g08337(.A1(new_n8618_), .A2(new_n807_), .A3(new_n7607_), .ZN(new_n8619_));
  OAI22_X1   g08338(.A1(new_n7619_), .A2(new_n298_), .B1(new_n325_), .B2(new_n8309_), .ZN(new_n8620_));
  AOI21_X1   g08339(.A1(new_n8620_), .A2(new_n8616_), .B(\a[47] ), .ZN(new_n8621_));
  OAI21_X1   g08340(.A1(new_n8621_), .A2(new_n7619_), .B(new_n329_), .ZN(new_n8622_));
  NAND2_X1   g08341(.A1(new_n8622_), .A2(new_n8619_), .ZN(new_n8623_));
  INV_X1     g08342(.I(\a[50] ), .ZN(new_n8624_));
  NAND2_X1   g08343(.A1(new_n8624_), .A2(\a[48] ), .ZN(new_n8625_));
  INV_X1     g08344(.I(\a[48] ), .ZN(new_n8626_));
  NAND2_X1   g08345(.A1(new_n8626_), .A2(\a[50] ), .ZN(new_n8627_));
  NAND2_X1   g08346(.A1(new_n7608_), .A2(\a[49] ), .ZN(new_n8628_));
  INV_X1     g08347(.I(\a[49] ), .ZN(new_n8629_));
  NAND2_X1   g08348(.A1(new_n8629_), .A2(\a[47] ), .ZN(new_n8630_));
  AOI22_X1   g08349(.A1(new_n8625_), .A2(new_n8627_), .B1(new_n8628_), .B2(new_n8630_), .ZN(new_n8631_));
  NOR3_X1    g08350(.A1(new_n8629_), .A2(\a[47] ), .A3(\a[48] ), .ZN(new_n8632_));
  NOR3_X1    g08351(.A1(new_n7608_), .A2(new_n8626_), .A3(\a[49] ), .ZN(new_n8633_));
  OAI21_X1   g08352(.A1(new_n8633_), .A2(new_n8632_), .B(\b[1] ), .ZN(new_n8634_));
  XOR2_X1    g08353(.A1(\a[48] ), .A2(\a[50] ), .Z(new_n8635_));
  XOR2_X1    g08354(.A1(\a[47] ), .A2(\a[49] ), .Z(new_n8636_));
  NAND3_X1   g08355(.A1(new_n8635_), .A2(new_n8636_), .A3(\b[0] ), .ZN(new_n8637_));
  NAND3_X1   g08356(.A1(new_n8637_), .A2(new_n8624_), .A3(new_n8634_), .ZN(new_n8638_));
  NAND3_X1   g08357(.A1(new_n8638_), .A2(new_n444_), .A3(new_n8631_), .ZN(new_n8639_));
  NOR2_X1    g08358(.A1(new_n8626_), .A2(\a[50] ), .ZN(new_n8640_));
  NOR2_X1    g08359(.A1(new_n8624_), .A2(\a[48] ), .ZN(new_n8641_));
  NOR2_X1    g08360(.A1(new_n8629_), .A2(\a[47] ), .ZN(new_n8642_));
  NOR2_X1    g08361(.A1(new_n7608_), .A2(\a[49] ), .ZN(new_n8643_));
  OAI22_X1   g08362(.A1(new_n8640_), .A2(new_n8641_), .B1(new_n8642_), .B2(new_n8643_), .ZN(new_n8644_));
  NAND3_X1   g08363(.A1(new_n7608_), .A2(new_n8626_), .A3(\a[49] ), .ZN(new_n8645_));
  NAND3_X1   g08364(.A1(new_n8629_), .A2(\a[47] ), .A3(\a[48] ), .ZN(new_n8646_));
  AOI21_X1   g08365(.A1(new_n8645_), .A2(new_n8646_), .B(new_n269_), .ZN(new_n8647_));
  XNOR2_X1   g08366(.A1(\a[48] ), .A2(\a[50] ), .ZN(new_n8648_));
  XNOR2_X1   g08367(.A1(\a[47] ), .A2(\a[49] ), .ZN(new_n8649_));
  NOR3_X1    g08368(.A1(new_n8648_), .A2(new_n8649_), .A3(new_n258_), .ZN(new_n8650_));
  NOR3_X1    g08369(.A1(new_n8650_), .A2(\a[50] ), .A3(new_n8647_), .ZN(new_n8651_));
  OAI21_X1   g08370(.A1(new_n8651_), .A2(new_n8644_), .B(new_n271_), .ZN(new_n8652_));
  NOR2_X1    g08371(.A1(new_n8314_), .A2(new_n8624_), .ZN(new_n8653_));
  INV_X1     g08372(.I(new_n8653_), .ZN(new_n8654_));
  NAND3_X1   g08373(.A1(new_n8652_), .A2(new_n8639_), .A3(new_n8654_), .ZN(new_n8655_));
  NOR3_X1    g08374(.A1(new_n8651_), .A2(new_n271_), .A3(new_n8644_), .ZN(new_n8656_));
  AOI21_X1   g08375(.A1(new_n8638_), .A2(new_n8631_), .B(new_n444_), .ZN(new_n8657_));
  OAI21_X1   g08376(.A1(new_n8656_), .A2(new_n8657_), .B(new_n8653_), .ZN(new_n8658_));
  NAND2_X1   g08377(.A1(new_n8658_), .A2(new_n8655_), .ZN(new_n8659_));
  NAND2_X1   g08378(.A1(new_n8659_), .A2(new_n8623_), .ZN(new_n8660_));
  NOR3_X1    g08379(.A1(new_n8621_), .A2(new_n329_), .A3(new_n7619_), .ZN(new_n8661_));
  AOI21_X1   g08380(.A1(new_n8618_), .A2(new_n7607_), .B(new_n807_), .ZN(new_n8662_));
  NOR2_X1    g08381(.A1(new_n8661_), .A2(new_n8662_), .ZN(new_n8663_));
  NAND3_X1   g08382(.A1(new_n8663_), .A2(new_n8655_), .A3(new_n8658_), .ZN(new_n8664_));
  NAND2_X1   g08383(.A1(new_n8664_), .A2(new_n8660_), .ZN(new_n8665_));
  NAND2_X1   g08384(.A1(new_n8613_), .A2(new_n8665_), .ZN(new_n8666_));
  AOI21_X1   g08385(.A1(new_n8610_), .A2(new_n8611_), .B(new_n8608_), .ZN(new_n8667_));
  NAND2_X1   g08386(.A1(new_n8659_), .A2(new_n8663_), .ZN(new_n8668_));
  NAND3_X1   g08387(.A1(new_n8623_), .A2(new_n8655_), .A3(new_n8658_), .ZN(new_n8669_));
  NAND2_X1   g08388(.A1(new_n8668_), .A2(new_n8669_), .ZN(new_n8670_));
  NAND2_X1   g08389(.A1(new_n8667_), .A2(new_n8670_), .ZN(new_n8671_));
  NAND2_X1   g08390(.A1(new_n8666_), .A2(new_n8671_), .ZN(new_n8672_));
  OAI22_X1   g08391(.A1(new_n6644_), .A2(new_n420_), .B1(new_n472_), .B2(new_n6647_), .ZN(new_n8673_));
  OAI21_X1   g08392(.A1(new_n419_), .A2(new_n7284_), .B(new_n8673_), .ZN(new_n8674_));
  AOI21_X1   g08393(.A1(new_n8674_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n8675_));
  XOR2_X1    g08394(.A1(new_n471_), .A2(new_n8675_), .Z(new_n8676_));
  INV_X1     g08395(.I(new_n8676_), .ZN(new_n8677_));
  NAND2_X1   g08396(.A1(new_n8672_), .A2(new_n8677_), .ZN(new_n8678_));
  INV_X1     g08397(.I(new_n8672_), .ZN(new_n8679_));
  NAND2_X1   g08398(.A1(new_n8679_), .A2(new_n8676_), .ZN(new_n8680_));
  NAND2_X1   g08399(.A1(new_n8680_), .A2(new_n8678_), .ZN(new_n8681_));
  NAND2_X1   g08400(.A1(new_n8681_), .A2(new_n8606_), .ZN(new_n8682_));
  NOR3_X1    g08401(.A1(new_n8605_), .A2(new_n8301_), .A3(new_n8302_), .ZN(new_n8683_));
  AOI21_X1   g08402(.A1(new_n8300_), .A2(new_n8601_), .B(new_n8683_), .ZN(new_n8684_));
  NAND3_X1   g08403(.A1(new_n8666_), .A2(new_n8671_), .A3(new_n8677_), .ZN(new_n8685_));
  AOI21_X1   g08404(.A1(new_n8660_), .A2(new_n8664_), .B(new_n8667_), .ZN(new_n8686_));
  INV_X1     g08405(.I(new_n8671_), .ZN(new_n8687_));
  OAI21_X1   g08406(.A1(new_n8687_), .A2(new_n8686_), .B(new_n8676_), .ZN(new_n8688_));
  NAND2_X1   g08407(.A1(new_n8688_), .A2(new_n8685_), .ZN(new_n8689_));
  NAND2_X1   g08408(.A1(new_n8684_), .A2(new_n8689_), .ZN(new_n8690_));
  OAI22_X1   g08409(.A1(new_n5993_), .A2(new_n565_), .B1(new_n656_), .B2(new_n5991_), .ZN(new_n8691_));
  OAI21_X1   g08410(.A1(new_n515_), .A2(new_n5997_), .B(new_n8691_), .ZN(new_n8692_));
  AOI21_X1   g08411(.A1(new_n8692_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n8693_));
  XNOR2_X1   g08412(.A1(new_n660_), .A2(new_n8693_), .ZN(new_n8694_));
  INV_X1     g08413(.I(new_n8694_), .ZN(new_n8695_));
  NAND3_X1   g08414(.A1(new_n8690_), .A2(new_n8682_), .A3(new_n8695_), .ZN(new_n8696_));
  AOI21_X1   g08415(.A1(new_n8678_), .A2(new_n8680_), .B(new_n8684_), .ZN(new_n8697_));
  AOI21_X1   g08416(.A1(new_n8685_), .A2(new_n8688_), .B(new_n8606_), .ZN(new_n8698_));
  OAI21_X1   g08417(.A1(new_n8697_), .A2(new_n8698_), .B(new_n8694_), .ZN(new_n8699_));
  NAND2_X1   g08418(.A1(new_n8699_), .A2(new_n8696_), .ZN(new_n8700_));
  NAND2_X1   g08419(.A1(new_n8599_), .A2(new_n8700_), .ZN(new_n8701_));
  NOR2_X1    g08420(.A1(new_n8346_), .A2(new_n8352_), .ZN(new_n8702_));
  NOR3_X1    g08421(.A1(new_n8338_), .A2(new_n8335_), .A3(new_n8005_), .ZN(new_n8703_));
  NOR2_X1    g08422(.A1(new_n8703_), .A2(new_n8342_), .ZN(new_n8704_));
  AOI21_X1   g08423(.A1(new_n8702_), .A2(new_n8704_), .B(new_n8595_), .ZN(new_n8705_));
  AOI21_X1   g08424(.A1(new_n8690_), .A2(new_n8682_), .B(new_n8694_), .ZN(new_n8706_));
  NOR3_X1    g08425(.A1(new_n8697_), .A2(new_n8698_), .A3(new_n8695_), .ZN(new_n8707_));
  OAI21_X1   g08426(.A1(new_n8706_), .A2(new_n8707_), .B(new_n8705_), .ZN(new_n8708_));
  OAI22_X1   g08427(.A1(new_n5420_), .A2(new_n780_), .B1(new_n861_), .B2(new_n5107_), .ZN(new_n8709_));
  OAI21_X1   g08428(.A1(new_n706_), .A2(new_n5112_), .B(new_n8709_), .ZN(new_n8710_));
  AOI21_X1   g08429(.A1(new_n8710_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n8711_));
  XNOR2_X1   g08430(.A1(new_n860_), .A2(new_n8711_), .ZN(new_n8712_));
  INV_X1     g08431(.I(new_n8712_), .ZN(new_n8713_));
  NAND3_X1   g08432(.A1(new_n8708_), .A2(new_n8701_), .A3(new_n8713_), .ZN(new_n8714_));
  AOI21_X1   g08433(.A1(new_n8696_), .A2(new_n8699_), .B(new_n8705_), .ZN(new_n8715_));
  NOR2_X1    g08434(.A1(new_n8707_), .A2(new_n8706_), .ZN(new_n8716_));
  NOR2_X1    g08435(.A1(new_n8716_), .A2(new_n8599_), .ZN(new_n8717_));
  OAI21_X1   g08436(.A1(new_n8715_), .A2(new_n8717_), .B(new_n8712_), .ZN(new_n8718_));
  NAND2_X1   g08437(.A1(new_n8718_), .A2(new_n8714_), .ZN(new_n8719_));
  OAI21_X1   g08438(.A1(new_n8593_), .A2(new_n8589_), .B(new_n8719_), .ZN(new_n8720_));
  INV_X1     g08439(.I(new_n8589_), .ZN(new_n8721_));
  NAND4_X1   g08440(.A1(new_n8292_), .A2(new_n8290_), .A3(new_n8590_), .A4(new_n8591_), .ZN(new_n8722_));
  AOI21_X1   g08441(.A1(new_n8708_), .A2(new_n8701_), .B(new_n8712_), .ZN(new_n8723_));
  INV_X1     g08442(.I(new_n8723_), .ZN(new_n8724_));
  NAND3_X1   g08443(.A1(new_n8708_), .A2(new_n8701_), .A3(new_n8712_), .ZN(new_n8725_));
  NAND2_X1   g08444(.A1(new_n8724_), .A2(new_n8725_), .ZN(new_n8726_));
  NAND3_X1   g08445(.A1(new_n8726_), .A2(new_n8721_), .A3(new_n8722_), .ZN(new_n8727_));
  OAI22_X1   g08446(.A1(new_n4072_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n4067_), .ZN(new_n8728_));
  OAI21_X1   g08447(.A1(new_n930_), .A2(new_n4318_), .B(new_n8728_), .ZN(new_n8729_));
  AOI21_X1   g08448(.A1(new_n8729_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n8730_));
  XOR2_X1    g08449(.A1(new_n1114_), .A2(new_n8730_), .Z(new_n8731_));
  INV_X1     g08450(.I(new_n8731_), .ZN(new_n8732_));
  NAND3_X1   g08451(.A1(new_n8727_), .A2(new_n8720_), .A3(new_n8732_), .ZN(new_n8733_));
  NOR2_X1    g08452(.A1(new_n8593_), .A2(new_n8589_), .ZN(new_n8734_));
  NOR3_X1    g08453(.A1(new_n8715_), .A2(new_n8717_), .A3(new_n8712_), .ZN(new_n8735_));
  AOI21_X1   g08454(.A1(new_n8708_), .A2(new_n8701_), .B(new_n8713_), .ZN(new_n8736_));
  NOR2_X1    g08455(.A1(new_n8735_), .A2(new_n8736_), .ZN(new_n8737_));
  NOR2_X1    g08456(.A1(new_n8734_), .A2(new_n8737_), .ZN(new_n8738_));
  INV_X1     g08457(.I(new_n8725_), .ZN(new_n8739_));
  NOR2_X1    g08458(.A1(new_n8739_), .A2(new_n8723_), .ZN(new_n8740_));
  NOR3_X1    g08459(.A1(new_n8740_), .A2(new_n8589_), .A3(new_n8593_), .ZN(new_n8741_));
  OAI21_X1   g08460(.A1(new_n8738_), .A2(new_n8741_), .B(new_n8731_), .ZN(new_n8742_));
  NAND2_X1   g08461(.A1(new_n8742_), .A2(new_n8733_), .ZN(new_n8743_));
  AOI21_X1   g08462(.A1(new_n8372_), .A2(new_n8376_), .B(new_n8392_), .ZN(new_n8744_));
  NAND3_X1   g08463(.A1(new_n8372_), .A2(new_n8376_), .A3(new_n8392_), .ZN(new_n8745_));
  NOR4_X1    g08464(.A1(new_n8383_), .A2(new_n7577_), .A3(new_n8384_), .A4(new_n8380_), .ZN(new_n8746_));
  AOI21_X1   g08465(.A1(new_n8746_), .A2(new_n8745_), .B(new_n8744_), .ZN(new_n8747_));
  NOR2_X1    g08466(.A1(new_n8747_), .A2(new_n8743_), .ZN(new_n8748_));
  NOR3_X1    g08467(.A1(new_n8738_), .A2(new_n8741_), .A3(new_n8731_), .ZN(new_n8749_));
  AOI21_X1   g08468(.A1(new_n8727_), .A2(new_n8720_), .B(new_n8732_), .ZN(new_n8750_));
  NOR2_X1    g08469(.A1(new_n8749_), .A2(new_n8750_), .ZN(new_n8751_));
  OAI21_X1   g08470(.A1(new_n8387_), .A2(new_n8386_), .B(new_n8284_), .ZN(new_n8752_));
  NOR3_X1    g08471(.A1(new_n8387_), .A2(new_n8386_), .A3(new_n8284_), .ZN(new_n8753_));
  NAND4_X1   g08472(.A1(new_n8285_), .A2(new_n7713_), .A3(new_n8286_), .A4(new_n8388_), .ZN(new_n8754_));
  OAI21_X1   g08473(.A1(new_n8754_), .A2(new_n8753_), .B(new_n8752_), .ZN(new_n8755_));
  NOR2_X1    g08474(.A1(new_n8755_), .A2(new_n8751_), .ZN(new_n8756_));
  OAI22_X1   g08475(.A1(new_n1294_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1518_), .ZN(new_n8757_));
  OAI21_X1   g08476(.A1(new_n1189_), .A2(new_n3569_), .B(new_n8757_), .ZN(new_n8758_));
  AOI21_X1   g08477(.A1(new_n8758_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n8759_));
  XNOR2_X1   g08478(.A1(new_n1421_), .A2(new_n8759_), .ZN(new_n8760_));
  NOR3_X1    g08479(.A1(new_n8756_), .A2(new_n8748_), .A3(new_n8760_), .ZN(new_n8761_));
  NAND2_X1   g08480(.A1(new_n8755_), .A2(new_n8751_), .ZN(new_n8762_));
  NAND2_X1   g08481(.A1(new_n8747_), .A2(new_n8743_), .ZN(new_n8763_));
  INV_X1     g08482(.I(new_n8760_), .ZN(new_n8764_));
  AOI21_X1   g08483(.A1(new_n8762_), .A2(new_n8763_), .B(new_n8764_), .ZN(new_n8765_));
  NOR2_X1    g08484(.A1(new_n8765_), .A2(new_n8761_), .ZN(new_n8766_));
  AOI21_X1   g08485(.A1(new_n8405_), .A2(new_n8406_), .B(new_n8066_), .ZN(new_n8767_));
  NOR3_X1    g08486(.A1(new_n8391_), .A2(new_n8395_), .A3(new_n8059_), .ZN(new_n8768_));
  NOR3_X1    g08487(.A1(new_n8404_), .A2(new_n8768_), .A3(new_n8399_), .ZN(new_n8769_));
  OAI21_X1   g08488(.A1(new_n8769_), .A2(new_n8767_), .B(new_n8766_), .ZN(new_n8770_));
  NAND3_X1   g08489(.A1(new_n8762_), .A2(new_n8763_), .A3(new_n8764_), .ZN(new_n8771_));
  OAI21_X1   g08490(.A1(new_n8756_), .A2(new_n8748_), .B(new_n8760_), .ZN(new_n8772_));
  NAND2_X1   g08491(.A1(new_n8772_), .A2(new_n8771_), .ZN(new_n8773_));
  INV_X1     g08492(.I(new_n8767_), .ZN(new_n8774_));
  NAND3_X1   g08493(.A1(new_n8405_), .A2(new_n8406_), .A3(new_n8066_), .ZN(new_n8775_));
  NAND3_X1   g08494(.A1(new_n8281_), .A2(new_n8400_), .A3(new_n8775_), .ZN(new_n8776_));
  NAND3_X1   g08495(.A1(new_n8776_), .A2(new_n8773_), .A3(new_n8774_), .ZN(new_n8777_));
  OAI22_X1   g08496(.A1(new_n1634_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1803_), .ZN(new_n8778_));
  OAI21_X1   g08497(.A1(new_n1525_), .A2(new_n2884_), .B(new_n8778_), .ZN(new_n8779_));
  AOI21_X1   g08498(.A1(new_n8779_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n8780_));
  XOR2_X1    g08499(.A1(new_n1808_), .A2(new_n8780_), .Z(new_n8781_));
  INV_X1     g08500(.I(new_n8781_), .ZN(new_n8782_));
  NAND3_X1   g08501(.A1(new_n8770_), .A2(new_n8777_), .A3(new_n8782_), .ZN(new_n8783_));
  AOI21_X1   g08502(.A1(new_n8776_), .A2(new_n8774_), .B(new_n8773_), .ZN(new_n8784_));
  NOR3_X1    g08503(.A1(new_n8769_), .A2(new_n8766_), .A3(new_n8767_), .ZN(new_n8785_));
  OAI21_X1   g08504(.A1(new_n8784_), .A2(new_n8785_), .B(new_n8781_), .ZN(new_n8786_));
  NAND2_X1   g08505(.A1(new_n8786_), .A2(new_n8783_), .ZN(new_n8787_));
  AOI21_X1   g08506(.A1(new_n8409_), .A2(new_n8412_), .B(new_n8077_), .ZN(new_n8788_));
  INV_X1     g08507(.I(new_n8788_), .ZN(new_n8789_));
  NAND3_X1   g08508(.A1(new_n8409_), .A2(new_n8412_), .A3(new_n8077_), .ZN(new_n8790_));
  NAND3_X1   g08509(.A1(new_n8279_), .A2(new_n8790_), .A3(new_n8418_), .ZN(new_n8791_));
  NAND2_X1   g08510(.A1(new_n8791_), .A2(new_n8789_), .ZN(new_n8792_));
  XOR2_X1    g08511(.A1(new_n8792_), .A2(new_n8787_), .Z(new_n8793_));
  OAI22_X1   g08512(.A1(new_n2171_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n2166_), .ZN(new_n8794_));
  OAI21_X1   g08513(.A1(new_n1936_), .A2(new_n2322_), .B(new_n8794_), .ZN(new_n8795_));
  AOI21_X1   g08514(.A1(new_n8795_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n8796_));
  XNOR2_X1   g08515(.A1(new_n2280_), .A2(new_n8796_), .ZN(new_n8797_));
  NOR2_X1    g08516(.A1(new_n8793_), .A2(new_n8797_), .ZN(new_n8798_));
  NOR3_X1    g08517(.A1(new_n8784_), .A2(new_n8785_), .A3(new_n8781_), .ZN(new_n8799_));
  AOI21_X1   g08518(.A1(new_n8770_), .A2(new_n8777_), .B(new_n8782_), .ZN(new_n8800_));
  NOR2_X1    g08519(.A1(new_n8799_), .A2(new_n8800_), .ZN(new_n8801_));
  XOR2_X1    g08520(.A1(new_n8792_), .A2(new_n8801_), .Z(new_n8802_));
  INV_X1     g08521(.I(new_n8797_), .ZN(new_n8803_));
  NOR2_X1    g08522(.A1(new_n8802_), .A2(new_n8803_), .ZN(new_n8804_));
  NOR2_X1    g08523(.A1(new_n8804_), .A2(new_n8798_), .ZN(new_n8805_));
  NAND2_X1   g08524(.A1(new_n8424_), .A2(new_n8427_), .ZN(new_n8806_));
  NAND2_X1   g08525(.A1(new_n8806_), .A2(new_n8440_), .ZN(new_n8807_));
  INV_X1     g08526(.I(new_n8431_), .ZN(new_n8808_));
  NAND3_X1   g08527(.A1(new_n8424_), .A2(new_n8427_), .A3(new_n8272_), .ZN(new_n8809_));
  NAND2_X1   g08528(.A1(new_n8809_), .A2(new_n8808_), .ZN(new_n8810_));
  OAI21_X1   g08529(.A1(new_n8810_), .A2(new_n8437_), .B(new_n8807_), .ZN(new_n8811_));
  NAND2_X1   g08530(.A1(new_n8805_), .A2(new_n8811_), .ZN(new_n8812_));
  NAND2_X1   g08531(.A1(new_n8802_), .A2(new_n8803_), .ZN(new_n8813_));
  NAND2_X1   g08532(.A1(new_n8793_), .A2(new_n8797_), .ZN(new_n8814_));
  NAND2_X1   g08533(.A1(new_n8813_), .A2(new_n8814_), .ZN(new_n8815_));
  INV_X1     g08534(.I(new_n8811_), .ZN(new_n8816_));
  NAND2_X1   g08535(.A1(new_n8816_), .A2(new_n8815_), .ZN(new_n8817_));
  OAI22_X1   g08536(.A1(new_n1712_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n1707_), .ZN(new_n8818_));
  OAI21_X1   g08537(.A1(new_n2439_), .A2(new_n1850_), .B(new_n8818_), .ZN(new_n8819_));
  AOI21_X1   g08538(.A1(new_n8819_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n8820_));
  XNOR2_X1   g08539(.A1(new_n2846_), .A2(new_n8820_), .ZN(new_n8821_));
  INV_X1     g08540(.I(new_n8821_), .ZN(new_n8822_));
  NAND3_X1   g08541(.A1(new_n8817_), .A2(new_n8812_), .A3(new_n8822_), .ZN(new_n8823_));
  NOR2_X1    g08542(.A1(new_n8816_), .A2(new_n8815_), .ZN(new_n8824_));
  NOR2_X1    g08543(.A1(new_n8805_), .A2(new_n8811_), .ZN(new_n8825_));
  OAI21_X1   g08544(.A1(new_n8824_), .A2(new_n8825_), .B(new_n8821_), .ZN(new_n8826_));
  NAND2_X1   g08545(.A1(new_n8826_), .A2(new_n8823_), .ZN(new_n8827_));
  NAND2_X1   g08546(.A1(new_n8588_), .A2(new_n8827_), .ZN(new_n8828_));
  AOI21_X1   g08547(.A1(new_n8585_), .A2(new_n8458_), .B(new_n8447_), .ZN(new_n8829_));
  AOI22_X1   g08548(.A1(new_n8829_), .A2(new_n8451_), .B1(new_n8269_), .B2(new_n8586_), .ZN(new_n8830_));
  INV_X1     g08549(.I(new_n8827_), .ZN(new_n8831_));
  NAND2_X1   g08550(.A1(new_n8831_), .A2(new_n8830_), .ZN(new_n8832_));
  OAI22_X1   g08551(.A1(new_n1347_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n1344_), .ZN(new_n8833_));
  OAI21_X1   g08552(.A1(new_n3018_), .A2(new_n1457_), .B(new_n8833_), .ZN(new_n8834_));
  AOI21_X1   g08553(.A1(new_n8834_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n8835_));
  XNOR2_X1   g08554(.A1(new_n3514_), .A2(new_n8835_), .ZN(new_n8836_));
  AOI21_X1   g08555(.A1(new_n8832_), .A2(new_n8828_), .B(new_n8836_), .ZN(new_n8837_));
  NOR2_X1    g08556(.A1(new_n8831_), .A2(new_n8830_), .ZN(new_n8838_));
  NOR2_X1    g08557(.A1(new_n8588_), .A2(new_n8827_), .ZN(new_n8839_));
  INV_X1     g08558(.I(new_n8836_), .ZN(new_n8840_));
  NOR3_X1    g08559(.A1(new_n8838_), .A2(new_n8839_), .A3(new_n8840_), .ZN(new_n8841_));
  NOR2_X1    g08560(.A1(new_n8841_), .A2(new_n8837_), .ZN(new_n8842_));
  NOR2_X1    g08561(.A1(new_n8457_), .A2(new_n8461_), .ZN(new_n8843_));
  NAND3_X1   g08562(.A1(new_n8471_), .A2(new_n8472_), .A3(new_n8261_), .ZN(new_n8844_));
  NAND2_X1   g08563(.A1(new_n8844_), .A2(new_n8466_), .ZN(new_n8845_));
  OAI22_X1   g08564(.A1(new_n8845_), .A2(new_n8470_), .B1(new_n8261_), .B2(new_n8843_), .ZN(new_n8846_));
  NAND2_X1   g08565(.A1(new_n8846_), .A2(new_n8842_), .ZN(new_n8847_));
  OAI21_X1   g08566(.A1(new_n8838_), .A2(new_n8839_), .B(new_n8840_), .ZN(new_n8848_));
  NAND3_X1   g08567(.A1(new_n8832_), .A2(new_n8828_), .A3(new_n8836_), .ZN(new_n8849_));
  NAND2_X1   g08568(.A1(new_n8848_), .A2(new_n8849_), .ZN(new_n8850_));
  NOR2_X1    g08569(.A1(new_n8843_), .A2(new_n8261_), .ZN(new_n8851_));
  AOI21_X1   g08570(.A1(new_n8843_), .A2(new_n8261_), .B(new_n8465_), .ZN(new_n8852_));
  AOI21_X1   g08571(.A1(new_n8852_), .A2(new_n8263_), .B(new_n8851_), .ZN(new_n8853_));
  NAND2_X1   g08572(.A1(new_n8853_), .A2(new_n8850_), .ZN(new_n8854_));
  OAI22_X1   g08573(.A1(new_n1055_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n1061_), .ZN(new_n8855_));
  OAI21_X1   g08574(.A1(new_n3717_), .A2(new_n1332_), .B(new_n8855_), .ZN(new_n8856_));
  AOI21_X1   g08575(.A1(new_n8856_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n8857_));
  XNOR2_X1   g08576(.A1(new_n4257_), .A2(new_n8857_), .ZN(new_n8858_));
  INV_X1     g08577(.I(new_n8858_), .ZN(new_n8859_));
  NAND3_X1   g08578(.A1(new_n8854_), .A2(new_n8847_), .A3(new_n8859_), .ZN(new_n8860_));
  NOR2_X1    g08579(.A1(new_n8853_), .A2(new_n8850_), .ZN(new_n8861_));
  NOR2_X1    g08580(.A1(new_n8846_), .A2(new_n8842_), .ZN(new_n8862_));
  OAI21_X1   g08581(.A1(new_n8861_), .A2(new_n8862_), .B(new_n8858_), .ZN(new_n8863_));
  NAND2_X1   g08582(.A1(new_n8863_), .A2(new_n8860_), .ZN(new_n8864_));
  AOI21_X1   g08583(.A1(new_n8475_), .A2(new_n8478_), .B(new_n8494_), .ZN(new_n8865_));
  NOR3_X1    g08584(.A1(new_n8488_), .A2(new_n8489_), .A3(new_n8256_), .ZN(new_n8866_));
  NOR2_X1    g08585(.A1(new_n8866_), .A2(new_n8482_), .ZN(new_n8867_));
  AOI21_X1   g08586(.A1(new_n8867_), .A2(new_n8495_), .B(new_n8865_), .ZN(new_n8868_));
  NOR2_X1    g08587(.A1(new_n8868_), .A2(new_n8864_), .ZN(new_n8869_));
  NOR3_X1    g08588(.A1(new_n8861_), .A2(new_n8862_), .A3(new_n8858_), .ZN(new_n8870_));
  AOI21_X1   g08589(.A1(new_n8854_), .A2(new_n8847_), .B(new_n8859_), .ZN(new_n8871_));
  NOR2_X1    g08590(.A1(new_n8871_), .A2(new_n8870_), .ZN(new_n8872_));
  NAND3_X1   g08591(.A1(new_n8487_), .A2(new_n7549_), .A3(new_n8258_), .ZN(new_n8873_));
  INV_X1     g08592(.I(new_n8865_), .ZN(new_n8874_));
  NAND3_X1   g08593(.A1(new_n8475_), .A2(new_n8478_), .A3(new_n8494_), .ZN(new_n8875_));
  NAND2_X1   g08594(.A1(new_n8875_), .A2(new_n8490_), .ZN(new_n8876_));
  OAI21_X1   g08595(.A1(new_n8873_), .A2(new_n8876_), .B(new_n8874_), .ZN(new_n8877_));
  NOR2_X1    g08596(.A1(new_n8877_), .A2(new_n8872_), .ZN(new_n8878_));
  OAI22_X1   g08597(.A1(new_n970_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n820_), .ZN(new_n8879_));
  OAI21_X1   g08598(.A1(new_n4500_), .A2(new_n894_), .B(new_n8879_), .ZN(new_n8880_));
  AOI21_X1   g08599(.A1(new_n8880_), .A2(new_n827_), .B(new_n970_), .ZN(new_n8881_));
  XOR2_X1    g08600(.A1(new_n5067_), .A2(new_n8881_), .Z(new_n8882_));
  NOR3_X1    g08601(.A1(new_n8869_), .A2(new_n8878_), .A3(new_n8882_), .ZN(new_n8883_));
  NAND2_X1   g08602(.A1(new_n8877_), .A2(new_n8872_), .ZN(new_n8884_));
  NAND2_X1   g08603(.A1(new_n8868_), .A2(new_n8864_), .ZN(new_n8885_));
  INV_X1     g08604(.I(new_n8882_), .ZN(new_n8886_));
  AOI21_X1   g08605(.A1(new_n8885_), .A2(new_n8884_), .B(new_n8886_), .ZN(new_n8887_));
  NOR2_X1    g08606(.A1(new_n8887_), .A2(new_n8883_), .ZN(new_n8888_));
  NOR2_X1    g08607(.A1(new_n8498_), .A2(new_n8493_), .ZN(new_n8889_));
  OAI21_X1   g08608(.A1(new_n8496_), .A2(new_n8497_), .B(new_n8494_), .ZN(new_n8890_));
  NAND3_X1   g08609(.A1(new_n8484_), .A2(new_n8492_), .A3(new_n8256_), .ZN(new_n8891_));
  NAND3_X1   g08610(.A1(new_n8890_), .A2(new_n8167_), .A3(new_n8891_), .ZN(new_n8892_));
  NAND2_X1   g08611(.A1(new_n8892_), .A2(new_n8503_), .ZN(new_n8893_));
  OAI22_X1   g08612(.A1(new_n8255_), .A2(new_n8893_), .B1(new_n8167_), .B2(new_n8889_), .ZN(new_n8894_));
  NAND2_X1   g08613(.A1(new_n8894_), .A2(new_n8888_), .ZN(new_n8895_));
  INV_X1     g08614(.I(new_n8888_), .ZN(new_n8896_));
  NOR2_X1    g08615(.A1(new_n8889_), .A2(new_n8167_), .ZN(new_n8897_));
  AOI21_X1   g08616(.A1(new_n8889_), .A2(new_n8167_), .B(new_n8502_), .ZN(new_n8898_));
  AOI21_X1   g08617(.A1(new_n8508_), .A2(new_n8898_), .B(new_n8897_), .ZN(new_n8899_));
  NAND2_X1   g08618(.A1(new_n8899_), .A2(new_n8896_), .ZN(new_n8900_));
  OAI22_X1   g08619(.A1(new_n607_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n610_), .ZN(new_n8901_));
  OAI21_X1   g08620(.A1(new_n5353_), .A2(new_n684_), .B(new_n8901_), .ZN(new_n8902_));
  AOI21_X1   g08621(.A1(new_n8902_), .A2(new_n612_), .B(new_n607_), .ZN(new_n8903_));
  XOR2_X1    g08622(.A1(new_n5926_), .A2(new_n8903_), .Z(new_n8904_));
  INV_X1     g08623(.I(new_n8904_), .ZN(new_n8905_));
  NAND3_X1   g08624(.A1(new_n8895_), .A2(new_n8900_), .A3(new_n8905_), .ZN(new_n8906_));
  NOR2_X1    g08625(.A1(new_n8899_), .A2(new_n8896_), .ZN(new_n8907_));
  NOR2_X1    g08626(.A1(new_n8894_), .A2(new_n8888_), .ZN(new_n8908_));
  OAI21_X1   g08627(.A1(new_n8908_), .A2(new_n8907_), .B(new_n8904_), .ZN(new_n8909_));
  NAND2_X1   g08628(.A1(new_n8909_), .A2(new_n8906_), .ZN(new_n8910_));
  INV_X1     g08629(.I(new_n8910_), .ZN(new_n8911_));
  OAI21_X1   g08630(.A1(new_n8510_), .A2(new_n8513_), .B(new_n8190_), .ZN(new_n8912_));
  NAND3_X1   g08631(.A1(new_n8523_), .A2(new_n8524_), .A3(new_n8183_), .ZN(new_n8913_));
  NAND2_X1   g08632(.A1(new_n8913_), .A2(new_n8518_), .ZN(new_n8914_));
  OAI21_X1   g08633(.A1(new_n8914_), .A2(new_n8522_), .B(new_n8912_), .ZN(new_n8915_));
  NAND2_X1   g08634(.A1(new_n8915_), .A2(new_n8911_), .ZN(new_n8916_));
  AOI21_X1   g08635(.A1(new_n8523_), .A2(new_n8524_), .B(new_n8183_), .ZN(new_n8917_));
  NOR3_X1    g08636(.A1(new_n8510_), .A2(new_n8513_), .A3(new_n8190_), .ZN(new_n8918_));
  NOR2_X1    g08637(.A1(new_n8918_), .A2(new_n8517_), .ZN(new_n8919_));
  AOI21_X1   g08638(.A1(new_n8919_), .A2(new_n8253_), .B(new_n8917_), .ZN(new_n8920_));
  NAND2_X1   g08639(.A1(new_n8920_), .A2(new_n8910_), .ZN(new_n8921_));
  OAI22_X1   g08640(.A1(new_n448_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n450_), .ZN(new_n8922_));
  OAI21_X1   g08641(.A1(new_n6229_), .A2(new_n496_), .B(new_n8922_), .ZN(new_n8923_));
  AOI21_X1   g08642(.A1(new_n8923_), .A2(new_n452_), .B(new_n448_), .ZN(new_n8924_));
  XOR2_X1    g08643(.A1(new_n6851_), .A2(new_n8924_), .Z(new_n8925_));
  INV_X1     g08644(.I(new_n8925_), .ZN(new_n8926_));
  NAND3_X1   g08645(.A1(new_n8921_), .A2(new_n8916_), .A3(new_n8926_), .ZN(new_n8927_));
  NOR2_X1    g08646(.A1(new_n8920_), .A2(new_n8910_), .ZN(new_n8928_));
  NOR2_X1    g08647(.A1(new_n8915_), .A2(new_n8911_), .ZN(new_n8929_));
  OAI21_X1   g08648(.A1(new_n8928_), .A2(new_n8929_), .B(new_n8925_), .ZN(new_n8930_));
  NAND2_X1   g08649(.A1(new_n8930_), .A2(new_n8927_), .ZN(new_n8931_));
  INV_X1     g08650(.I(new_n8931_), .ZN(new_n8932_));
  NAND2_X1   g08651(.A1(new_n8531_), .A2(new_n8199_), .ZN(new_n8933_));
  NAND3_X1   g08652(.A1(new_n8527_), .A2(new_n8530_), .A3(new_n8200_), .ZN(new_n8934_));
  NAND2_X1   g08653(.A1(new_n8934_), .A2(new_n8536_), .ZN(new_n8935_));
  OAI21_X1   g08654(.A1(new_n8541_), .A2(new_n8935_), .B(new_n8933_), .ZN(new_n8936_));
  NAND2_X1   g08655(.A1(new_n8932_), .A2(new_n8936_), .ZN(new_n8937_));
  NOR2_X1    g08656(.A1(new_n8932_), .A2(new_n8936_), .ZN(new_n8938_));
  INV_X1     g08657(.I(new_n8938_), .ZN(new_n8939_));
  NAND2_X1   g08658(.A1(new_n8939_), .A2(new_n8937_), .ZN(new_n8940_));
  INV_X1     g08659(.I(new_n8940_), .ZN(new_n8941_));
  INV_X1     g08660(.I(new_n8547_), .ZN(new_n8942_));
  NOR2_X1    g08661(.A1(new_n8942_), .A2(new_n8551_), .ZN(new_n8943_));
  NOR3_X1    g08662(.A1(new_n7892_), .A2(new_n7894_), .A3(new_n8209_), .ZN(new_n8944_));
  OAI21_X1   g08663(.A1(new_n7892_), .A2(new_n7894_), .B(new_n8209_), .ZN(new_n8945_));
  AOI21_X1   g08664(.A1(new_n8945_), .A2(new_n8243_), .B(new_n8944_), .ZN(new_n8946_));
  AOI21_X1   g08665(.A1(new_n8942_), .A2(new_n8551_), .B(new_n8946_), .ZN(new_n8947_));
  INV_X1     g08666(.I(\b[49] ), .ZN(new_n8948_));
  NOR2_X1    g08667(.A1(new_n8948_), .A2(\b[47] ), .ZN(new_n8949_));
  NOR2_X1    g08668(.A1(new_n8218_), .A2(\b[49] ), .ZN(new_n8950_));
  OAI21_X1   g08669(.A1(new_n8949_), .A2(new_n8950_), .B(new_n8562_), .ZN(new_n8951_));
  XNOR2_X1   g08670(.A1(new_n8559_), .A2(new_n8951_), .ZN(new_n8952_));
  OAI22_X1   g08671(.A1(new_n330_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n263_), .ZN(new_n8953_));
  OAI21_X1   g08672(.A1(new_n8218_), .A2(new_n289_), .B(new_n8953_), .ZN(new_n8954_));
  AOI21_X1   g08673(.A1(new_n8954_), .A2(new_n260_), .B(new_n426_), .ZN(new_n8955_));
  XOR2_X1    g08674(.A1(new_n8952_), .A2(new_n8955_), .Z(new_n8956_));
  NOR3_X1    g08675(.A1(new_n8947_), .A2(new_n8943_), .A3(new_n8956_), .ZN(new_n8957_));
  OAI21_X1   g08676(.A1(new_n8947_), .A2(new_n8943_), .B(new_n8956_), .ZN(new_n8958_));
  INV_X1     g08677(.I(new_n8958_), .ZN(new_n8959_));
  OAI21_X1   g08678(.A1(new_n8959_), .A2(new_n8957_), .B(new_n8941_), .ZN(new_n8960_));
  INV_X1     g08679(.I(new_n8957_), .ZN(new_n8961_));
  NAND3_X1   g08680(.A1(new_n8961_), .A2(new_n8940_), .A3(new_n8958_), .ZN(new_n8962_));
  AOI21_X1   g08681(.A1(new_n8960_), .A2(new_n8962_), .B(new_n8584_), .ZN(new_n8963_));
  AND3_X2    g08682(.A1(new_n8960_), .A2(new_n8962_), .A3(new_n8584_), .Z(new_n8964_));
  NOR2_X1    g08683(.A1(new_n8964_), .A2(new_n8963_), .ZN(new_n8965_));
  XOR2_X1    g08684(.A1(new_n8553_), .A2(new_n8946_), .Z(new_n8966_));
  NAND2_X1   g08685(.A1(new_n8576_), .A2(new_n8233_), .ZN(new_n8967_));
  AOI21_X1   g08686(.A1(new_n8230_), .A2(new_n8967_), .B(new_n8226_), .ZN(new_n8968_));
  AOI21_X1   g08687(.A1(new_n8572_), .A2(new_n8966_), .B(new_n8968_), .ZN(new_n8969_));
  XOR2_X1    g08688(.A1(new_n8969_), .A2(new_n8965_), .Z(\f[49] ));
  NAND2_X1   g08689(.A1(new_n8966_), .A2(new_n8572_), .ZN(new_n8971_));
  INV_X1     g08690(.I(new_n8956_), .ZN(new_n8972_));
  OR3_X2     g08691(.A1(new_n8947_), .A2(new_n8941_), .A3(new_n8943_), .Z(new_n8973_));
  OAI21_X1   g08692(.A1(new_n8947_), .A2(new_n8943_), .B(new_n8941_), .ZN(new_n8974_));
  AOI21_X1   g08693(.A1(new_n8973_), .A2(new_n8974_), .B(new_n8584_), .ZN(new_n8975_));
  AND3_X2    g08694(.A1(new_n8973_), .A2(new_n8584_), .A3(new_n8974_), .Z(new_n8976_));
  OAI21_X1   g08695(.A1(new_n8976_), .A2(new_n8975_), .B(new_n8972_), .ZN(new_n8977_));
  OAI21_X1   g08696(.A1(new_n8965_), .A2(new_n8977_), .B(new_n8971_), .ZN(new_n8978_));
  NAND2_X1   g08697(.A1(new_n8968_), .A2(new_n8978_), .ZN(new_n8979_));
  NAND4_X1   g08698(.A1(new_n8540_), .A2(new_n8539_), .A3(new_n8934_), .A4(new_n8536_), .ZN(new_n8980_));
  AOI21_X1   g08699(.A1(new_n8980_), .A2(new_n8933_), .B(new_n8583_), .ZN(new_n8981_));
  INV_X1     g08700(.I(new_n8933_), .ZN(new_n8982_));
  AOI21_X1   g08701(.A1(new_n8529_), .A2(new_n8528_), .B(new_n8190_), .ZN(new_n8983_));
  NOR3_X1    g08702(.A1(new_n8520_), .A2(new_n8526_), .A3(new_n8183_), .ZN(new_n8984_));
  NOR3_X1    g08703(.A1(new_n8983_), .A2(new_n8984_), .A3(new_n8199_), .ZN(new_n8985_));
  NOR4_X1    g08704(.A1(new_n8250_), .A2(new_n8985_), .A3(new_n8249_), .A4(new_n8535_), .ZN(new_n8986_));
  NOR3_X1    g08705(.A1(new_n8986_), .A2(new_n8982_), .A3(new_n8584_), .ZN(new_n8987_));
  OAI21_X1   g08706(.A1(new_n8987_), .A2(new_n8981_), .B(new_n8931_), .ZN(new_n8988_));
  NOR3_X1    g08707(.A1(new_n8986_), .A2(new_n8982_), .A3(new_n8583_), .ZN(new_n8989_));
  AOI21_X1   g08708(.A1(new_n8980_), .A2(new_n8933_), .B(new_n8584_), .ZN(new_n8990_));
  OAI21_X1   g08709(.A1(new_n8989_), .A2(new_n8990_), .B(new_n8932_), .ZN(new_n8991_));
  NAND2_X1   g08710(.A1(new_n8988_), .A2(new_n8991_), .ZN(new_n8992_));
  AOI21_X1   g08711(.A1(new_n8992_), .A2(new_n8552_), .B(new_n8547_), .ZN(new_n8993_));
  NAND2_X1   g08712(.A1(new_n8936_), .A2(new_n8584_), .ZN(new_n8994_));
  NAND3_X1   g08713(.A1(new_n8980_), .A2(new_n8583_), .A3(new_n8933_), .ZN(new_n8995_));
  AOI21_X1   g08714(.A1(new_n8994_), .A2(new_n8995_), .B(new_n8932_), .ZN(new_n8996_));
  NAND3_X1   g08715(.A1(new_n8980_), .A2(new_n8584_), .A3(new_n8933_), .ZN(new_n8997_));
  OAI21_X1   g08716(.A1(new_n8986_), .A2(new_n8982_), .B(new_n8583_), .ZN(new_n8998_));
  AOI21_X1   g08717(.A1(new_n8998_), .A2(new_n8997_), .B(new_n8931_), .ZN(new_n8999_));
  NOR3_X1    g08718(.A1(new_n8996_), .A2(new_n8552_), .A3(new_n8999_), .ZN(new_n9000_));
  NOR3_X1    g08719(.A1(new_n8946_), .A2(new_n8993_), .A3(new_n9000_), .ZN(new_n9001_));
  NAND2_X1   g08720(.A1(new_n8940_), .A2(new_n8583_), .ZN(new_n9002_));
  OAI21_X1   g08721(.A1(new_n8936_), .A2(new_n8931_), .B(new_n8930_), .ZN(new_n9003_));
  AOI21_X1   g08722(.A1(new_n8895_), .A2(new_n8900_), .B(new_n8905_), .ZN(new_n9004_));
  OAI22_X1   g08723(.A1(new_n1803_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n1936_), .ZN(new_n9005_));
  OAI21_X1   g08724(.A1(new_n1634_), .A2(new_n2884_), .B(new_n9005_), .ZN(new_n9006_));
  AOI21_X1   g08725(.A1(new_n9006_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n9007_));
  XNOR2_X1   g08726(.A1(new_n1940_), .A2(new_n9007_), .ZN(new_n9008_));
  INV_X1     g08727(.I(new_n9008_), .ZN(new_n9009_));
  NOR2_X1    g08728(.A1(new_n8768_), .A2(new_n8399_), .ZN(new_n9010_));
  AOI21_X1   g08729(.A1(new_n9010_), .A2(new_n8281_), .B(new_n8767_), .ZN(new_n9011_));
  INV_X1     g08730(.I(new_n8696_), .ZN(new_n9012_));
  AOI21_X1   g08731(.A1(new_n8599_), .A2(new_n8699_), .B(new_n9012_), .ZN(new_n9013_));
  INV_X1     g08732(.I(new_n8678_), .ZN(new_n9014_));
  AOI21_X1   g08733(.A1(new_n8645_), .A2(new_n8646_), .B(new_n280_), .ZN(new_n9015_));
  AOI21_X1   g08734(.A1(new_n8631_), .A2(\b[1] ), .B(new_n9015_), .ZN(new_n9016_));
  XNOR2_X1   g08735(.A1(\a[47] ), .A2(\a[50] ), .ZN(new_n9017_));
  NOR4_X1    g08736(.A1(new_n8313_), .A2(new_n8649_), .A3(new_n9017_), .A4(new_n258_), .ZN(new_n9018_));
  OAI21_X1   g08737(.A1(new_n9016_), .A2(new_n9018_), .B(new_n8624_), .ZN(new_n9019_));
  NAND3_X1   g08738(.A1(new_n9019_), .A2(new_n490_), .A3(new_n8631_), .ZN(new_n9020_));
  OAI21_X1   g08739(.A1(new_n8633_), .A2(new_n8632_), .B(\b[2] ), .ZN(new_n9021_));
  OAI21_X1   g08740(.A1(new_n8644_), .A2(new_n269_), .B(new_n9021_), .ZN(new_n9022_));
  XOR2_X1    g08741(.A1(\a[47] ), .A2(\a[48] ), .Z(new_n9023_));
  XOR2_X1    g08742(.A1(\a[47] ), .A2(\a[50] ), .Z(new_n9024_));
  NAND4_X1   g08743(.A1(new_n9023_), .A2(new_n8636_), .A3(new_n9024_), .A4(\b[0] ), .ZN(new_n9025_));
  AOI21_X1   g08744(.A1(new_n9022_), .A2(new_n9025_), .B(\a[50] ), .ZN(new_n9026_));
  OAI21_X1   g08745(.A1(new_n9026_), .A2(new_n8644_), .B(new_n282_), .ZN(new_n9027_));
  NAND2_X1   g08746(.A1(new_n9027_), .A2(new_n9020_), .ZN(new_n9028_));
  NAND3_X1   g08747(.A1(new_n8652_), .A2(new_n8639_), .A3(new_n8653_), .ZN(new_n9029_));
  AOI21_X1   g08748(.A1(new_n374_), .A2(new_n377_), .B(new_n7619_), .ZN(new_n9030_));
  NOR3_X1    g08749(.A1(new_n7605_), .A2(new_n7606_), .A3(new_n325_), .ZN(new_n9031_));
  NOR2_X1    g08750(.A1(new_n8309_), .A2(new_n419_), .ZN(new_n9032_));
  OAI22_X1   g08751(.A1(new_n9031_), .A2(new_n9032_), .B1(new_n7947_), .B2(new_n298_), .ZN(new_n9033_));
  NOR2_X1    g08752(.A1(new_n9030_), .A2(new_n9033_), .ZN(new_n9034_));
  NAND2_X1   g08753(.A1(new_n9029_), .A2(new_n9034_), .ZN(new_n9035_));
  OAI21_X1   g08754(.A1(new_n2332_), .A2(new_n2331_), .B(new_n7607_), .ZN(new_n9036_));
  NAND3_X1   g08755(.A1(new_n7614_), .A2(new_n7615_), .A3(\b[4] ), .ZN(new_n9037_));
  NAND2_X1   g08756(.A1(new_n7940_), .A2(\b[5] ), .ZN(new_n9038_));
  AOI22_X1   g08757(.A1(new_n8308_), .A2(\b[3] ), .B1(new_n9038_), .B2(new_n9037_), .ZN(new_n9039_));
  NAND2_X1   g08758(.A1(new_n9036_), .A2(new_n9039_), .ZN(new_n9040_));
  NAND4_X1   g08759(.A1(new_n9040_), .A2(new_n8639_), .A3(new_n8652_), .A4(new_n8653_), .ZN(new_n9041_));
  AOI21_X1   g08760(.A1(new_n9035_), .A2(new_n9041_), .B(new_n9028_), .ZN(new_n9042_));
  NOR3_X1    g08761(.A1(new_n9026_), .A2(new_n282_), .A3(new_n8644_), .ZN(new_n9043_));
  AOI21_X1   g08762(.A1(new_n9019_), .A2(new_n8631_), .B(new_n490_), .ZN(new_n9044_));
  NOR2_X1    g08763(.A1(new_n9043_), .A2(new_n9044_), .ZN(new_n9045_));
  NOR3_X1    g08764(.A1(new_n8656_), .A2(new_n8657_), .A3(new_n8654_), .ZN(new_n9046_));
  NOR2_X1    g08765(.A1(new_n9046_), .A2(new_n9040_), .ZN(new_n9047_));
  NOR4_X1    g08766(.A1(new_n9034_), .A2(new_n8656_), .A3(new_n8657_), .A4(new_n8654_), .ZN(new_n9048_));
  NOR3_X1    g08767(.A1(new_n9047_), .A2(new_n9048_), .A3(new_n9045_), .ZN(new_n9049_));
  OAI21_X1   g08768(.A1(new_n9049_), .A2(new_n9042_), .B(new_n7608_), .ZN(new_n9050_));
  OAI21_X1   g08769(.A1(new_n9047_), .A2(new_n9048_), .B(new_n9045_), .ZN(new_n9051_));
  NAND3_X1   g08770(.A1(new_n9035_), .A2(new_n9041_), .A3(new_n9028_), .ZN(new_n9052_));
  NAND3_X1   g08771(.A1(new_n9051_), .A2(new_n9052_), .A3(\a[47] ), .ZN(new_n9053_));
  NAND2_X1   g08772(.A1(new_n9050_), .A2(new_n9053_), .ZN(new_n9054_));
  NAND3_X1   g08773(.A1(new_n9054_), .A2(new_n8660_), .A3(new_n8670_), .ZN(new_n9055_));
  NAND2_X1   g08774(.A1(new_n8659_), .A2(new_n8623_), .ZN(new_n9057_));
  AOI21_X1   g08775(.A1(new_n9055_), .A2(new_n9057_), .B(new_n8613_), .ZN(new_n9058_));
  INV_X1     g08776(.I(new_n8660_), .ZN(new_n9059_));
  AOI21_X1   g08777(.A1(new_n9051_), .A2(new_n9052_), .B(\a[47] ), .ZN(new_n9060_));
  NOR3_X1    g08778(.A1(new_n9049_), .A2(new_n9042_), .A3(new_n7608_), .ZN(new_n9061_));
  OAI21_X1   g08779(.A1(new_n9061_), .A2(new_n9060_), .B(new_n8670_), .ZN(new_n9062_));
  NOR2_X1    g08780(.A1(new_n9062_), .A2(new_n9059_), .ZN(new_n9063_));
  INV_X1     g08781(.I(new_n9057_), .ZN(new_n9064_));
  NOR3_X1    g08782(.A1(new_n9063_), .A2(new_n8667_), .A3(new_n9064_), .ZN(new_n9065_));
  OAI22_X1   g08783(.A1(new_n6644_), .A2(new_n472_), .B1(new_n515_), .B2(new_n6647_), .ZN(new_n9066_));
  OAI21_X1   g08784(.A1(new_n420_), .A2(new_n7284_), .B(new_n9066_), .ZN(new_n9067_));
  AOI21_X1   g08785(.A1(new_n9067_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n9068_));
  XOR2_X1    g08786(.A1(new_n700_), .A2(new_n9068_), .Z(new_n9069_));
  NOR3_X1    g08787(.A1(new_n9065_), .A2(new_n9058_), .A3(new_n9069_), .ZN(new_n9070_));
  OAI21_X1   g08788(.A1(new_n9063_), .A2(new_n9064_), .B(new_n8667_), .ZN(new_n9071_));
  NAND3_X1   g08789(.A1(new_n9055_), .A2(new_n8613_), .A3(new_n9057_), .ZN(new_n9072_));
  INV_X1     g08790(.I(new_n9069_), .ZN(new_n9073_));
  AOI21_X1   g08791(.A1(new_n9071_), .A2(new_n9072_), .B(new_n9073_), .ZN(new_n9074_));
  OAI21_X1   g08792(.A1(new_n9070_), .A2(new_n9074_), .B(new_n8689_), .ZN(new_n9075_));
  NOR2_X1    g08793(.A1(new_n9075_), .A2(new_n9014_), .ZN(new_n9076_));
  NAND3_X1   g08794(.A1(new_n9071_), .A2(new_n9072_), .A3(new_n9073_), .ZN(new_n9077_));
  OAI21_X1   g08795(.A1(new_n9065_), .A2(new_n9058_), .B(new_n9069_), .ZN(new_n9078_));
  NAND2_X1   g08796(.A1(new_n9078_), .A2(new_n9077_), .ZN(new_n9079_));
  NOR2_X1    g08797(.A1(new_n8679_), .A2(new_n8676_), .ZN(new_n9081_));
  OAI21_X1   g08798(.A1(new_n9076_), .A2(new_n9081_), .B(new_n8684_), .ZN(new_n9082_));
  NAND3_X1   g08799(.A1(new_n9079_), .A2(new_n8678_), .A3(new_n8689_), .ZN(new_n9083_));
  INV_X1     g08800(.I(new_n9081_), .ZN(new_n9084_));
  NAND3_X1   g08801(.A1(new_n9083_), .A2(new_n8606_), .A3(new_n9084_), .ZN(new_n9085_));
  OAI22_X1   g08802(.A1(new_n5993_), .A2(new_n656_), .B1(new_n706_), .B2(new_n5991_), .ZN(new_n9086_));
  OAI21_X1   g08803(.A1(new_n565_), .A2(new_n5997_), .B(new_n9086_), .ZN(new_n9087_));
  AOI21_X1   g08804(.A1(new_n9087_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n9088_));
  XOR2_X1    g08805(.A1(new_n710_), .A2(new_n9088_), .Z(new_n9089_));
  NAND3_X1   g08806(.A1(new_n9082_), .A2(new_n9085_), .A3(new_n9089_), .ZN(new_n9090_));
  AOI21_X1   g08807(.A1(new_n9083_), .A2(new_n9084_), .B(new_n8606_), .ZN(new_n9091_));
  NOR3_X1    g08808(.A1(new_n9076_), .A2(new_n8684_), .A3(new_n9081_), .ZN(new_n9092_));
  INV_X1     g08809(.I(new_n9089_), .ZN(new_n9093_));
  OAI21_X1   g08810(.A1(new_n9092_), .A2(new_n9091_), .B(new_n9093_), .ZN(new_n9094_));
  OAI22_X1   g08811(.A1(new_n5420_), .A2(new_n861_), .B1(new_n930_), .B2(new_n5107_), .ZN(new_n9095_));
  OAI21_X1   g08812(.A1(new_n780_), .A2(new_n5112_), .B(new_n9095_), .ZN(new_n9096_));
  AOI21_X1   g08813(.A1(new_n9096_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n9097_));
  XOR2_X1    g08814(.A1(new_n937_), .A2(new_n9097_), .Z(new_n9098_));
  NAND3_X1   g08815(.A1(new_n9094_), .A2(new_n9090_), .A3(new_n9098_), .ZN(new_n9099_));
  NOR3_X1    g08816(.A1(new_n9092_), .A2(new_n9091_), .A3(new_n9093_), .ZN(new_n9100_));
  AOI21_X1   g08817(.A1(new_n9082_), .A2(new_n9085_), .B(new_n9089_), .ZN(new_n9101_));
  XNOR2_X1   g08818(.A1(new_n937_), .A2(new_n9097_), .ZN(new_n9102_));
  OAI21_X1   g08819(.A1(new_n9100_), .A2(new_n9101_), .B(new_n9102_), .ZN(new_n9103_));
  AOI21_X1   g08820(.A1(new_n9103_), .A2(new_n9099_), .B(new_n9013_), .ZN(new_n9104_));
  AOI21_X1   g08821(.A1(new_n8690_), .A2(new_n8682_), .B(new_n8695_), .ZN(new_n9105_));
  OAI21_X1   g08822(.A1(new_n8705_), .A2(new_n9105_), .B(new_n8696_), .ZN(new_n9106_));
  OAI21_X1   g08823(.A1(new_n9100_), .A2(new_n9101_), .B(new_n9098_), .ZN(new_n9107_));
  NAND3_X1   g08824(.A1(new_n9094_), .A2(new_n9090_), .A3(new_n9102_), .ZN(new_n9108_));
  AOI21_X1   g08825(.A1(new_n9107_), .A2(new_n9108_), .B(new_n9106_), .ZN(new_n9109_));
  NOR2_X1    g08826(.A1(new_n9104_), .A2(new_n9109_), .ZN(new_n9110_));
  NOR3_X1    g08827(.A1(new_n9110_), .A2(new_n8737_), .A3(new_n8723_), .ZN(new_n9111_));
  NAND2_X1   g08828(.A1(new_n8708_), .A2(new_n8701_), .ZN(new_n9112_));
  NOR2_X1    g08829(.A1(new_n9100_), .A2(new_n9101_), .ZN(new_n9113_));
  NAND2_X1   g08830(.A1(new_n9112_), .A2(new_n8713_), .ZN(new_n9114_));
  INV_X1     g08831(.I(new_n9114_), .ZN(new_n9115_));
  OAI21_X1   g08832(.A1(new_n9111_), .A2(new_n9115_), .B(new_n8734_), .ZN(new_n9116_));
  NAND2_X1   g08833(.A1(new_n8292_), .A2(new_n8290_), .ZN(new_n9117_));
  OAI21_X1   g08834(.A1(new_n9117_), .A2(new_n8592_), .B(new_n8721_), .ZN(new_n9118_));
  NOR3_X1    g08835(.A1(new_n9100_), .A2(new_n9101_), .A3(new_n9102_), .ZN(new_n9119_));
  AOI21_X1   g08836(.A1(new_n9094_), .A2(new_n9090_), .B(new_n9098_), .ZN(new_n9120_));
  OAI21_X1   g08837(.A1(new_n9119_), .A2(new_n9120_), .B(new_n9106_), .ZN(new_n9121_));
  AOI21_X1   g08838(.A1(new_n9094_), .A2(new_n9090_), .B(new_n9102_), .ZN(new_n9122_));
  NOR3_X1    g08839(.A1(new_n9100_), .A2(new_n9101_), .A3(new_n9098_), .ZN(new_n9123_));
  OAI21_X1   g08840(.A1(new_n9123_), .A2(new_n9122_), .B(new_n9013_), .ZN(new_n9124_));
  NAND2_X1   g08841(.A1(new_n9121_), .A2(new_n9124_), .ZN(new_n9125_));
  NAND3_X1   g08842(.A1(new_n9125_), .A2(new_n8719_), .A3(new_n8724_), .ZN(new_n9126_));
  NAND3_X1   g08843(.A1(new_n9126_), .A2(new_n9118_), .A3(new_n9114_), .ZN(new_n9127_));
  OAI22_X1   g08844(.A1(new_n4072_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n4067_), .ZN(new_n9128_));
  OAI21_X1   g08845(.A1(new_n1017_), .A2(new_n4318_), .B(new_n9128_), .ZN(new_n9129_));
  AOI21_X1   g08846(.A1(new_n9129_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n9130_));
  XNOR2_X1   g08847(.A1(new_n1196_), .A2(new_n9130_), .ZN(new_n9131_));
  INV_X1     g08848(.I(new_n9131_), .ZN(new_n9132_));
  NAND3_X1   g08849(.A1(new_n9116_), .A2(new_n9127_), .A3(new_n9132_), .ZN(new_n9133_));
  AOI21_X1   g08850(.A1(new_n9126_), .A2(new_n9114_), .B(new_n9118_), .ZN(new_n9134_));
  NOR3_X1    g08851(.A1(new_n9111_), .A2(new_n8734_), .A3(new_n9115_), .ZN(new_n9135_));
  OAI21_X1   g08852(.A1(new_n9135_), .A2(new_n9134_), .B(new_n9131_), .ZN(new_n9136_));
  NAND3_X1   g08853(.A1(new_n9136_), .A2(new_n9133_), .A3(new_n8742_), .ZN(new_n9137_));
  NAND3_X1   g08854(.A1(new_n9137_), .A2(new_n8751_), .A3(new_n8755_), .ZN(new_n9138_));
  NOR3_X1    g08855(.A1(new_n9135_), .A2(new_n9134_), .A3(new_n9131_), .ZN(new_n9139_));
  AOI21_X1   g08856(.A1(new_n9116_), .A2(new_n9127_), .B(new_n9132_), .ZN(new_n9140_));
  NOR3_X1    g08857(.A1(new_n9139_), .A2(new_n9140_), .A3(new_n8750_), .ZN(new_n9141_));
  OAI21_X1   g08858(.A1(new_n9141_), .A2(new_n8747_), .B(new_n8743_), .ZN(new_n9142_));
  OAI22_X1   g08859(.A1(new_n1518_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1525_), .ZN(new_n9143_));
  OAI21_X1   g08860(.A1(new_n1294_), .A2(new_n3569_), .B(new_n9143_), .ZN(new_n9144_));
  AOI21_X1   g08861(.A1(new_n9144_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n9145_));
  XOR2_X1    g08862(.A1(new_n1530_), .A2(new_n9145_), .Z(new_n9146_));
  AOI21_X1   g08863(.A1(new_n9142_), .A2(new_n9138_), .B(new_n9146_), .ZN(new_n9147_));
  NOR3_X1    g08864(.A1(new_n9141_), .A2(new_n8743_), .A3(new_n8747_), .ZN(new_n9148_));
  AOI21_X1   g08865(.A1(new_n9137_), .A2(new_n8755_), .B(new_n8751_), .ZN(new_n9149_));
  INV_X1     g08866(.I(new_n9146_), .ZN(new_n9150_));
  NOR3_X1    g08867(.A1(new_n9148_), .A2(new_n9149_), .A3(new_n9150_), .ZN(new_n9151_));
  NOR3_X1    g08868(.A1(new_n9151_), .A2(new_n9147_), .A3(new_n8765_), .ZN(new_n9152_));
  NOR3_X1    g08869(.A1(new_n9152_), .A2(new_n9011_), .A3(new_n8773_), .ZN(new_n9153_));
  NAND2_X1   g08870(.A1(new_n8776_), .A2(new_n8774_), .ZN(new_n9154_));
  OAI21_X1   g08871(.A1(new_n9148_), .A2(new_n9149_), .B(new_n9150_), .ZN(new_n9155_));
  NAND3_X1   g08872(.A1(new_n9142_), .A2(new_n9138_), .A3(new_n9146_), .ZN(new_n9156_));
  NAND3_X1   g08873(.A1(new_n9155_), .A2(new_n9156_), .A3(new_n8772_), .ZN(new_n9157_));
  AOI21_X1   g08874(.A1(new_n9154_), .A2(new_n9157_), .B(new_n8766_), .ZN(new_n9158_));
  NOR2_X1    g08875(.A1(new_n9158_), .A2(new_n9153_), .ZN(new_n9159_));
  NAND3_X1   g08876(.A1(new_n8791_), .A2(new_n8801_), .A3(new_n8789_), .ZN(new_n9160_));
  OAI22_X1   g08877(.A1(new_n2171_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n2166_), .ZN(new_n9161_));
  OAI21_X1   g08878(.A1(new_n2102_), .A2(new_n2322_), .B(new_n9161_), .ZN(new_n9162_));
  AOI21_X1   g08879(.A1(new_n9162_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n9163_));
  XNOR2_X1   g08880(.A1(new_n2443_), .A2(new_n9163_), .ZN(new_n9164_));
  AOI21_X1   g08881(.A1(new_n9160_), .A2(new_n8786_), .B(new_n9164_), .ZN(new_n9165_));
  AOI21_X1   g08882(.A1(new_n8410_), .A2(new_n8411_), .B(new_n8059_), .ZN(new_n9166_));
  NOR3_X1    g08883(.A1(new_n8408_), .A2(new_n8402_), .A3(new_n8066_), .ZN(new_n9167_));
  NOR3_X1    g08884(.A1(new_n9166_), .A2(new_n9167_), .A3(new_n8084_), .ZN(new_n9168_));
  NOR3_X1    g08885(.A1(new_n8422_), .A2(new_n9168_), .A3(new_n8417_), .ZN(new_n9169_));
  NOR3_X1    g08886(.A1(new_n9169_), .A2(new_n8787_), .A3(new_n8788_), .ZN(new_n9170_));
  INV_X1     g08887(.I(new_n9164_), .ZN(new_n9171_));
  NOR3_X1    g08888(.A1(new_n9170_), .A2(new_n8800_), .A3(new_n9171_), .ZN(new_n9172_));
  OAI21_X1   g08889(.A1(new_n9172_), .A2(new_n9165_), .B(new_n9159_), .ZN(new_n9173_));
  INV_X1     g08890(.I(new_n9159_), .ZN(new_n9174_));
  OAI21_X1   g08891(.A1(new_n9170_), .A2(new_n8800_), .B(new_n9171_), .ZN(new_n9175_));
  NAND3_X1   g08892(.A1(new_n9160_), .A2(new_n8786_), .A3(new_n9164_), .ZN(new_n9176_));
  NAND3_X1   g08893(.A1(new_n9175_), .A2(new_n9176_), .A3(new_n9174_), .ZN(new_n9177_));
  AOI21_X1   g08894(.A1(new_n9173_), .A2(new_n9177_), .B(new_n9009_), .ZN(new_n9178_));
  AOI21_X1   g08895(.A1(new_n9175_), .A2(new_n9176_), .B(new_n9174_), .ZN(new_n9179_));
  NOR3_X1    g08896(.A1(new_n9172_), .A2(new_n9165_), .A3(new_n9159_), .ZN(new_n9180_));
  NOR3_X1    g08897(.A1(new_n9180_), .A2(new_n9179_), .A3(new_n9008_), .ZN(new_n9181_));
  NOR3_X1    g08898(.A1(new_n9181_), .A2(new_n9178_), .A3(new_n8804_), .ZN(new_n9182_));
  NOR3_X1    g08899(.A1(new_n9182_), .A2(new_n8816_), .A3(new_n8815_), .ZN(new_n9183_));
  OAI21_X1   g08900(.A1(new_n9180_), .A2(new_n9179_), .B(new_n9008_), .ZN(new_n9184_));
  NAND3_X1   g08901(.A1(new_n9173_), .A2(new_n9177_), .A3(new_n9009_), .ZN(new_n9185_));
  NAND3_X1   g08902(.A1(new_n9184_), .A2(new_n9185_), .A3(new_n8814_), .ZN(new_n9186_));
  AOI21_X1   g08903(.A1(new_n9186_), .A2(new_n8811_), .B(new_n8805_), .ZN(new_n9187_));
  OAI22_X1   g08904(.A1(new_n1712_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n1707_), .ZN(new_n9188_));
  OAI21_X1   g08905(.A1(new_n2643_), .A2(new_n1850_), .B(new_n9188_), .ZN(new_n9189_));
  AOI21_X1   g08906(.A1(new_n9189_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n9190_));
  XNOR2_X1   g08907(.A1(new_n3022_), .A2(new_n9190_), .ZN(new_n9191_));
  INV_X1     g08908(.I(new_n9191_), .ZN(new_n9192_));
  OAI21_X1   g08909(.A1(new_n9183_), .A2(new_n9187_), .B(new_n9192_), .ZN(new_n9193_));
  NAND3_X1   g08910(.A1(new_n9186_), .A2(new_n8805_), .A3(new_n8811_), .ZN(new_n9194_));
  OAI21_X1   g08911(.A1(new_n9182_), .A2(new_n8816_), .B(new_n8815_), .ZN(new_n9195_));
  NAND3_X1   g08912(.A1(new_n9195_), .A2(new_n9194_), .A3(new_n9191_), .ZN(new_n9196_));
  NAND3_X1   g08913(.A1(new_n9193_), .A2(new_n9196_), .A3(new_n8826_), .ZN(new_n9197_));
  NAND3_X1   g08914(.A1(new_n9197_), .A2(new_n8830_), .A3(new_n8827_), .ZN(new_n9198_));
  AOI21_X1   g08915(.A1(new_n8817_), .A2(new_n8812_), .B(new_n8822_), .ZN(new_n9199_));
  AOI21_X1   g08916(.A1(new_n9195_), .A2(new_n9194_), .B(new_n9191_), .ZN(new_n9200_));
  NOR3_X1    g08917(.A1(new_n9183_), .A2(new_n9187_), .A3(new_n9192_), .ZN(new_n9201_));
  NOR3_X1    g08918(.A1(new_n9201_), .A2(new_n9200_), .A3(new_n9199_), .ZN(new_n9202_));
  OAI21_X1   g08919(.A1(new_n9202_), .A2(new_n8831_), .B(new_n8588_), .ZN(new_n9203_));
  OAI22_X1   g08920(.A1(new_n1347_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n1344_), .ZN(new_n9204_));
  OAI21_X1   g08921(.A1(new_n3260_), .A2(new_n1457_), .B(new_n9204_), .ZN(new_n9205_));
  AOI21_X1   g08922(.A1(new_n9205_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n9206_));
  XOR2_X1    g08923(.A1(new_n3722_), .A2(new_n9206_), .Z(new_n9207_));
  AOI21_X1   g08924(.A1(new_n9203_), .A2(new_n9198_), .B(new_n9207_), .ZN(new_n9208_));
  NOR3_X1    g08925(.A1(new_n9202_), .A2(new_n8831_), .A3(new_n8588_), .ZN(new_n9209_));
  AOI21_X1   g08926(.A1(new_n9197_), .A2(new_n8827_), .B(new_n8830_), .ZN(new_n9210_));
  INV_X1     g08927(.I(new_n9207_), .ZN(new_n9211_));
  NOR3_X1    g08928(.A1(new_n9209_), .A2(new_n9210_), .A3(new_n9211_), .ZN(new_n9212_));
  NOR3_X1    g08929(.A1(new_n9212_), .A2(new_n9208_), .A3(new_n8841_), .ZN(new_n9213_));
  NOR3_X1    g08930(.A1(new_n9213_), .A2(new_n8853_), .A3(new_n8850_), .ZN(new_n9214_));
  OAI21_X1   g08931(.A1(new_n9209_), .A2(new_n9210_), .B(new_n9211_), .ZN(new_n9215_));
  NAND3_X1   g08932(.A1(new_n9203_), .A2(new_n9198_), .A3(new_n9207_), .ZN(new_n9216_));
  NAND3_X1   g08933(.A1(new_n9215_), .A2(new_n9216_), .A3(new_n8849_), .ZN(new_n9217_));
  AOI21_X1   g08934(.A1(new_n9217_), .A2(new_n8846_), .B(new_n8842_), .ZN(new_n9218_));
  OAI22_X1   g08935(.A1(new_n1055_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n1061_), .ZN(new_n9219_));
  OAI21_X1   g08936(.A1(new_n3989_), .A2(new_n1332_), .B(new_n9219_), .ZN(new_n9220_));
  AOI21_X1   g08937(.A1(new_n9220_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n9221_));
  XOR2_X1    g08938(.A1(new_n4499_), .A2(new_n9221_), .Z(new_n9222_));
  NOR3_X1    g08939(.A1(new_n9214_), .A2(new_n9218_), .A3(new_n9222_), .ZN(new_n9223_));
  NAND3_X1   g08940(.A1(new_n9217_), .A2(new_n8846_), .A3(new_n8842_), .ZN(new_n9224_));
  OAI21_X1   g08941(.A1(new_n9213_), .A2(new_n8853_), .B(new_n8850_), .ZN(new_n9225_));
  INV_X1     g08942(.I(new_n9222_), .ZN(new_n9226_));
  AOI21_X1   g08943(.A1(new_n9225_), .A2(new_n9224_), .B(new_n9226_), .ZN(new_n9227_));
  NOR3_X1    g08944(.A1(new_n9223_), .A2(new_n9227_), .A3(new_n8871_), .ZN(new_n9228_));
  NOR3_X1    g08945(.A1(new_n9228_), .A2(new_n8868_), .A3(new_n8864_), .ZN(new_n9229_));
  NAND3_X1   g08946(.A1(new_n9225_), .A2(new_n9224_), .A3(new_n9226_), .ZN(new_n9230_));
  OAI21_X1   g08947(.A1(new_n9214_), .A2(new_n9218_), .B(new_n9222_), .ZN(new_n9231_));
  NAND3_X1   g08948(.A1(new_n9231_), .A2(new_n9230_), .A3(new_n8863_), .ZN(new_n9232_));
  AOI21_X1   g08949(.A1(new_n9232_), .A2(new_n8877_), .B(new_n8872_), .ZN(new_n9233_));
  OAI22_X1   g08950(.A1(new_n970_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n820_), .ZN(new_n9234_));
  OAI21_X1   g08951(.A1(new_n4774_), .A2(new_n894_), .B(new_n9234_), .ZN(new_n9235_));
  AOI21_X1   g08952(.A1(new_n9235_), .A2(new_n827_), .B(new_n970_), .ZN(new_n9236_));
  XNOR2_X1   g08953(.A1(new_n5357_), .A2(new_n9236_), .ZN(new_n9237_));
  NOR3_X1    g08954(.A1(new_n9229_), .A2(new_n9233_), .A3(new_n9237_), .ZN(new_n9238_));
  NAND3_X1   g08955(.A1(new_n9232_), .A2(new_n8877_), .A3(new_n8872_), .ZN(new_n9239_));
  OAI21_X1   g08956(.A1(new_n9228_), .A2(new_n8868_), .B(new_n8864_), .ZN(new_n9240_));
  INV_X1     g08957(.I(new_n9237_), .ZN(new_n9241_));
  AOI21_X1   g08958(.A1(new_n9240_), .A2(new_n9239_), .B(new_n9241_), .ZN(new_n9242_));
  NOR3_X1    g08959(.A1(new_n9238_), .A2(new_n9242_), .A3(new_n8887_), .ZN(new_n9243_));
  NOR3_X1    g08960(.A1(new_n8899_), .A2(new_n8896_), .A3(new_n9243_), .ZN(new_n9244_));
  OAI21_X1   g08961(.A1(new_n8869_), .A2(new_n8878_), .B(new_n8882_), .ZN(new_n9245_));
  NAND3_X1   g08962(.A1(new_n9240_), .A2(new_n9239_), .A3(new_n9241_), .ZN(new_n9246_));
  OAI21_X1   g08963(.A1(new_n9229_), .A2(new_n9233_), .B(new_n9237_), .ZN(new_n9247_));
  NAND3_X1   g08964(.A1(new_n9247_), .A2(new_n9246_), .A3(new_n9245_), .ZN(new_n9248_));
  AOI21_X1   g08965(.A1(new_n8894_), .A2(new_n9248_), .B(new_n8888_), .ZN(new_n9249_));
  OAI22_X1   g08966(.A1(new_n607_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n610_), .ZN(new_n9250_));
  OAI21_X1   g08967(.A1(new_n5913_), .A2(new_n684_), .B(new_n9250_), .ZN(new_n9251_));
  AOI21_X1   g08968(.A1(new_n9251_), .A2(new_n612_), .B(new_n607_), .ZN(new_n9252_));
  XOR2_X1    g08969(.A1(new_n6233_), .A2(new_n9252_), .Z(new_n9253_));
  NOR3_X1    g08970(.A1(new_n9249_), .A2(new_n9244_), .A3(new_n9253_), .ZN(new_n9254_));
  NAND3_X1   g08971(.A1(new_n8894_), .A2(new_n8888_), .A3(new_n9248_), .ZN(new_n9255_));
  OAI21_X1   g08972(.A1(new_n8899_), .A2(new_n9243_), .B(new_n8896_), .ZN(new_n9256_));
  INV_X1     g08973(.I(new_n9253_), .ZN(new_n9257_));
  AOI21_X1   g08974(.A1(new_n9255_), .A2(new_n9256_), .B(new_n9257_), .ZN(new_n9258_));
  NOR3_X1    g08975(.A1(new_n9258_), .A2(new_n9254_), .A3(new_n9004_), .ZN(new_n9259_));
  NOR3_X1    g08976(.A1(new_n8920_), .A2(new_n8910_), .A3(new_n9259_), .ZN(new_n9260_));
  NAND3_X1   g08977(.A1(new_n9255_), .A2(new_n9256_), .A3(new_n9257_), .ZN(new_n9261_));
  OAI21_X1   g08978(.A1(new_n9249_), .A2(new_n9244_), .B(new_n9253_), .ZN(new_n9262_));
  NAND3_X1   g08979(.A1(new_n9262_), .A2(new_n9261_), .A3(new_n8909_), .ZN(new_n9263_));
  AOI21_X1   g08980(.A1(new_n8915_), .A2(new_n9263_), .B(new_n8911_), .ZN(new_n9264_));
  OAI22_X1   g08981(.A1(new_n448_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n450_), .ZN(new_n9265_));
  OAI21_X1   g08982(.A1(new_n6538_), .A2(new_n496_), .B(new_n9265_), .ZN(new_n9266_));
  AOI21_X1   g08983(.A1(new_n9266_), .A2(new_n452_), .B(new_n448_), .ZN(new_n9267_));
  XNOR2_X1   g08984(.A1(new_n7202_), .A2(new_n9267_), .ZN(new_n9268_));
  NOR3_X1    g08985(.A1(new_n9260_), .A2(new_n9264_), .A3(new_n9268_), .ZN(new_n9269_));
  NAND3_X1   g08986(.A1(new_n8915_), .A2(new_n8911_), .A3(new_n9263_), .ZN(new_n9270_));
  OAI21_X1   g08987(.A1(new_n8920_), .A2(new_n9259_), .B(new_n8910_), .ZN(new_n9271_));
  INV_X1     g08988(.I(new_n9268_), .ZN(new_n9272_));
  AOI21_X1   g08989(.A1(new_n9271_), .A2(new_n9270_), .B(new_n9272_), .ZN(new_n9273_));
  NOR2_X1    g08990(.A1(new_n9269_), .A2(new_n9273_), .ZN(new_n9274_));
  OAI21_X1   g08991(.A1(new_n9260_), .A2(new_n9264_), .B(new_n9272_), .ZN(new_n9275_));
  NAND3_X1   g08992(.A1(new_n9271_), .A2(new_n9270_), .A3(new_n9268_), .ZN(new_n9276_));
  NAND2_X1   g08993(.A1(new_n9275_), .A2(new_n9276_), .ZN(new_n9277_));
  NAND2_X1   g08994(.A1(new_n9003_), .A2(new_n9277_), .ZN(new_n9278_));
  OAI21_X1   g08995(.A1(new_n9003_), .A2(new_n9274_), .B(new_n9278_), .ZN(new_n9279_));
  OAI22_X1   g08996(.A1(new_n7870_), .A2(new_n341_), .B1(new_n404_), .B2(new_n8218_), .ZN(new_n9280_));
  OAI21_X1   g08997(.A1(new_n7864_), .A2(new_n366_), .B(new_n9280_), .ZN(new_n9281_));
  AOI21_X1   g08998(.A1(new_n9281_), .A2(new_n334_), .B(new_n341_), .ZN(new_n9282_));
  XOR2_X1    g08999(.A1(new_n8217_), .A2(new_n9282_), .Z(new_n9283_));
  INV_X1     g09000(.I(new_n9283_), .ZN(new_n9284_));
  NAND2_X1   g09001(.A1(new_n9279_), .A2(new_n9284_), .ZN(new_n9285_));
  XOR2_X1    g09002(.A1(new_n9285_), .A2(new_n9002_), .Z(new_n9286_));
  XOR2_X1    g09003(.A1(new_n9286_), .A2(new_n9001_), .Z(new_n9287_));
  NOR2_X1    g09004(.A1(\b[48] ), .A2(\b[49] ), .ZN(new_n9288_));
  AOI21_X1   g09005(.A1(new_n8559_), .A2(new_n9288_), .B(new_n8218_), .ZN(new_n9289_));
  NOR2_X1    g09006(.A1(new_n8563_), .A2(new_n8948_), .ZN(new_n9290_));
  INV_X1     g09007(.I(new_n9290_), .ZN(new_n9291_));
  NOR2_X1    g09008(.A1(new_n8559_), .A2(new_n9291_), .ZN(new_n9292_));
  NOR2_X1    g09009(.A1(new_n9289_), .A2(new_n9292_), .ZN(new_n9293_));
  XNOR2_X1   g09010(.A1(\b[49] ), .A2(\b[50] ), .ZN(new_n9294_));
  INV_X1     g09011(.I(\b[50] ), .ZN(new_n9295_));
  NOR2_X1    g09012(.A1(new_n8948_), .A2(new_n9295_), .ZN(new_n9296_));
  NOR2_X1    g09013(.A1(\b[49] ), .A2(\b[50] ), .ZN(new_n9297_));
  OAI21_X1   g09014(.A1(new_n9296_), .A2(new_n9297_), .B(new_n9293_), .ZN(new_n9298_));
  OAI21_X1   g09015(.A1(new_n9293_), .A2(new_n9294_), .B(new_n9298_), .ZN(new_n9299_));
  OAI22_X1   g09016(.A1(new_n330_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n263_), .ZN(new_n9300_));
  OAI21_X1   g09017(.A1(new_n8563_), .A2(new_n289_), .B(new_n9300_), .ZN(new_n9301_));
  AOI21_X1   g09018(.A1(new_n9301_), .A2(new_n260_), .B(new_n426_), .ZN(new_n9302_));
  XNOR2_X1   g09019(.A1(new_n9299_), .A2(new_n9302_), .ZN(new_n9303_));
  INV_X1     g09020(.I(new_n9303_), .ZN(new_n9304_));
  AND2_X2    g09021(.A1(new_n9287_), .A2(new_n9304_), .Z(new_n9305_));
  NOR2_X1    g09022(.A1(new_n9287_), .A2(new_n9304_), .ZN(new_n9306_));
  NOR2_X1    g09023(.A1(new_n9305_), .A2(new_n9306_), .ZN(new_n9307_));
  XOR2_X1    g09024(.A1(new_n9287_), .A2(new_n9304_), .Z(new_n9308_));
  NAND2_X1   g09025(.A1(new_n8979_), .A2(new_n9308_), .ZN(new_n9309_));
  OAI21_X1   g09026(.A1(new_n8979_), .A2(new_n9307_), .B(new_n9309_), .ZN(\f[50] ));
  OAI21_X1   g09027(.A1(new_n8996_), .A2(new_n8999_), .B(new_n8552_), .ZN(new_n9311_));
  NAND2_X1   g09028(.A1(new_n9311_), .A2(new_n8942_), .ZN(new_n9312_));
  INV_X1     g09029(.I(new_n9000_), .ZN(new_n9313_));
  NAND4_X1   g09030(.A1(new_n9312_), .A2(new_n8245_), .A3(new_n9313_), .A4(new_n9279_), .ZN(new_n9314_));
  NAND2_X1   g09031(.A1(new_n8945_), .A2(new_n8243_), .ZN(new_n9315_));
  AOI21_X1   g09032(.A1(new_n9315_), .A2(new_n8241_), .B(new_n9000_), .ZN(new_n9316_));
  AOI21_X1   g09033(.A1(new_n9316_), .A2(new_n9312_), .B(new_n9279_), .ZN(new_n9317_));
  NOR2_X1    g09034(.A1(new_n9002_), .A2(new_n9283_), .ZN(new_n9318_));
  INV_X1     g09035(.I(new_n9318_), .ZN(new_n9319_));
  OAI21_X1   g09036(.A1(new_n9317_), .A2(new_n9319_), .B(new_n9314_), .ZN(new_n9320_));
  INV_X1     g09037(.I(new_n9320_), .ZN(new_n9321_));
  INV_X1     g09038(.I(new_n9273_), .ZN(new_n9322_));
  AOI21_X1   g09039(.A1(new_n9275_), .A2(new_n9276_), .B(new_n8930_), .ZN(new_n9323_));
  OAI21_X1   g09040(.A1(new_n8936_), .A2(new_n9323_), .B(new_n8931_), .ZN(new_n9324_));
  NAND2_X1   g09041(.A1(new_n9324_), .A2(new_n9322_), .ZN(new_n9325_));
  INV_X1     g09042(.I(new_n9325_), .ZN(new_n9326_));
  NAND3_X1   g09043(.A1(new_n8253_), .A2(new_n8913_), .A3(new_n8518_), .ZN(new_n9327_));
  OAI21_X1   g09044(.A1(new_n9258_), .A2(new_n9254_), .B(new_n9004_), .ZN(new_n9328_));
  NAND3_X1   g09045(.A1(new_n9328_), .A2(new_n9327_), .A3(new_n8912_), .ZN(new_n9329_));
  AOI21_X1   g09046(.A1(new_n9247_), .A2(new_n9246_), .B(new_n9245_), .ZN(new_n9330_));
  OAI21_X1   g09047(.A1(new_n8894_), .A2(new_n9330_), .B(new_n8896_), .ZN(new_n9331_));
  OAI21_X1   g09048(.A1(new_n9223_), .A2(new_n9227_), .B(new_n8871_), .ZN(new_n9332_));
  AOI21_X1   g09049(.A1(new_n9332_), .A2(new_n8868_), .B(new_n8872_), .ZN(new_n9333_));
  AOI21_X1   g09050(.A1(new_n9203_), .A2(new_n9198_), .B(new_n9211_), .ZN(new_n9334_));
  AOI21_X1   g09051(.A1(new_n9215_), .A2(new_n9216_), .B(new_n8849_), .ZN(new_n9335_));
  OAI21_X1   g09052(.A1(new_n9335_), .A2(new_n8846_), .B(new_n8850_), .ZN(new_n9336_));
  AOI21_X1   g09053(.A1(new_n9195_), .A2(new_n9194_), .B(new_n9192_), .ZN(new_n9337_));
  INV_X1     g09054(.I(new_n9337_), .ZN(new_n9338_));
  AOI21_X1   g09055(.A1(new_n8823_), .A2(new_n8826_), .B(new_n8830_), .ZN(new_n9340_));
  OAI21_X1   g09056(.A1(new_n9170_), .A2(new_n8800_), .B(new_n9174_), .ZN(new_n9341_));
  NAND3_X1   g09057(.A1(new_n9160_), .A2(new_n8786_), .A3(new_n9159_), .ZN(new_n9342_));
  NAND2_X1   g09058(.A1(new_n9341_), .A2(new_n9342_), .ZN(new_n9343_));
  NAND2_X1   g09059(.A1(new_n9343_), .A2(new_n9008_), .ZN(new_n9344_));
  NAND3_X1   g09060(.A1(new_n9341_), .A2(new_n9342_), .A3(new_n9009_), .ZN(new_n9345_));
  AOI21_X1   g09061(.A1(new_n9344_), .A2(new_n9345_), .B(new_n9164_), .ZN(new_n9346_));
  AOI21_X1   g09062(.A1(new_n9184_), .A2(new_n9185_), .B(new_n8814_), .ZN(new_n9347_));
  OAI21_X1   g09063(.A1(new_n9347_), .A2(new_n8811_), .B(new_n8815_), .ZN(new_n9348_));
  NOR2_X1    g09064(.A1(new_n9159_), .A2(new_n9009_), .ZN(new_n9349_));
  INV_X1     g09065(.I(new_n9349_), .ZN(new_n9350_));
  NOR2_X1    g09066(.A1(new_n9169_), .A2(new_n8788_), .ZN(new_n9351_));
  NAND3_X1   g09067(.A1(new_n9154_), .A2(new_n9157_), .A3(new_n8766_), .ZN(new_n9352_));
  OAI21_X1   g09068(.A1(new_n9152_), .A2(new_n9011_), .B(new_n8773_), .ZN(new_n9353_));
  AOI21_X1   g09069(.A1(new_n9353_), .A2(new_n9352_), .B(new_n9008_), .ZN(new_n9354_));
  NOR3_X1    g09070(.A1(new_n9158_), .A2(new_n9153_), .A3(new_n9009_), .ZN(new_n9355_));
  OAI21_X1   g09071(.A1(new_n9355_), .A2(new_n9354_), .B(new_n8800_), .ZN(new_n9356_));
  AOI21_X1   g09072(.A1(new_n9351_), .A2(new_n9356_), .B(new_n8801_), .ZN(new_n9357_));
  AOI21_X1   g09073(.A1(new_n9155_), .A2(new_n9156_), .B(new_n8772_), .ZN(new_n9358_));
  OAI21_X1   g09074(.A1(new_n9154_), .A2(new_n9358_), .B(new_n8773_), .ZN(new_n9359_));
  OAI21_X1   g09075(.A1(new_n9139_), .A2(new_n9140_), .B(new_n8750_), .ZN(new_n9360_));
  AOI21_X1   g09076(.A1(new_n9360_), .A2(new_n8747_), .B(new_n8751_), .ZN(new_n9361_));
  NAND2_X1   g09077(.A1(new_n9094_), .A2(new_n9090_), .ZN(new_n9362_));
  XOR2_X1    g09078(.A1(new_n9013_), .A2(new_n9362_), .Z(new_n9363_));
  NAND2_X1   g09079(.A1(new_n9363_), .A2(new_n9102_), .ZN(new_n9364_));
  INV_X1     g09080(.I(new_n9364_), .ZN(new_n9365_));
  AOI21_X1   g09081(.A1(new_n9125_), .A2(new_n8713_), .B(new_n9112_), .ZN(new_n9366_));
  OAI22_X1   g09082(.A1(new_n8713_), .A2(new_n9125_), .B1(new_n8593_), .B2(new_n8589_), .ZN(new_n9367_));
  NAND3_X1   g09083(.A1(new_n9082_), .A2(new_n9085_), .A3(new_n9093_), .ZN(new_n9368_));
  AOI21_X1   g09084(.A1(new_n9079_), .A2(new_n8672_), .B(new_n8677_), .ZN(new_n9369_));
  NAND3_X1   g09085(.A1(new_n9078_), .A2(new_n9077_), .A3(new_n8679_), .ZN(new_n9370_));
  NAND2_X1   g09086(.A1(new_n9370_), .A2(new_n8606_), .ZN(new_n9371_));
  XOR2_X1    g09087(.A1(new_n9040_), .A2(\a[47] ), .Z(new_n9372_));
  NAND2_X1   g09088(.A1(new_n9028_), .A2(new_n9029_), .ZN(new_n9373_));
  NAND2_X1   g09089(.A1(new_n9045_), .A2(new_n9046_), .ZN(new_n9374_));
  AOI21_X1   g09090(.A1(new_n9373_), .A2(new_n9374_), .B(new_n9372_), .ZN(new_n9375_));
  INV_X1     g09091(.I(new_n9375_), .ZN(new_n9376_));
  OAI21_X1   g09092(.A1(new_n9061_), .A2(new_n9060_), .B(new_n8659_), .ZN(new_n9377_));
  NAND2_X1   g09093(.A1(new_n9377_), .A2(new_n8663_), .ZN(new_n9378_));
  NOR3_X1    g09094(.A1(new_n9061_), .A2(new_n9060_), .A3(new_n8659_), .ZN(new_n9379_));
  NOR2_X1    g09095(.A1(new_n9379_), .A2(new_n8667_), .ZN(new_n9380_));
  NAND4_X1   g09096(.A1(new_n9023_), .A2(new_n8636_), .A3(new_n9024_), .A4(\b[1] ), .ZN(new_n9381_));
  NAND2_X1   g09097(.A1(new_n8645_), .A2(new_n8646_), .ZN(new_n9382_));
  AOI22_X1   g09098(.A1(new_n8631_), .A2(\b[2] ), .B1(\b[3] ), .B2(new_n9382_), .ZN(new_n9383_));
  NAND2_X1   g09099(.A1(new_n9383_), .A2(new_n9381_), .ZN(new_n9384_));
  AOI21_X1   g09100(.A1(new_n296_), .A2(new_n300_), .B(new_n8644_), .ZN(new_n9385_));
  AOI21_X1   g09101(.A1(new_n9384_), .A2(new_n9385_), .B(new_n8624_), .ZN(new_n9386_));
  NOR4_X1    g09102(.A1(new_n8313_), .A2(new_n8649_), .A3(new_n9017_), .A4(new_n269_), .ZN(new_n9387_));
  NOR2_X1    g09103(.A1(new_n8633_), .A2(new_n8632_), .ZN(new_n9388_));
  OAI22_X1   g09104(.A1(new_n8644_), .A2(new_n280_), .B1(new_n298_), .B2(new_n9388_), .ZN(new_n9389_));
  NOR2_X1    g09105(.A1(new_n9389_), .A2(new_n9387_), .ZN(new_n9390_));
  INV_X1     g09106(.I(new_n9385_), .ZN(new_n9391_));
  NOR3_X1    g09107(.A1(new_n9390_), .A2(new_n9391_), .A3(\a[50] ), .ZN(new_n9392_));
  NOR2_X1    g09108(.A1(new_n9392_), .A2(new_n9386_), .ZN(new_n9393_));
  NAND2_X1   g09109(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n9394_));
  NOR2_X1    g09110(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n9395_));
  INV_X1     g09111(.I(new_n9395_), .ZN(new_n9396_));
  NAND2_X1   g09112(.A1(new_n9396_), .A2(new_n9394_), .ZN(new_n9397_));
  NOR2_X1    g09113(.A1(new_n9397_), .A2(new_n258_), .ZN(new_n9398_));
  INV_X1     g09114(.I(new_n9398_), .ZN(new_n9399_));
  NOR2_X1    g09115(.A1(new_n9393_), .A2(new_n9399_), .ZN(new_n9400_));
  NAND2_X1   g09116(.A1(new_n9400_), .A2(new_n9045_), .ZN(new_n9401_));
  OAI21_X1   g09117(.A1(new_n9393_), .A2(new_n9399_), .B(new_n9028_), .ZN(new_n9402_));
  AOI21_X1   g09118(.A1(new_n9401_), .A2(new_n9402_), .B(new_n9046_), .ZN(new_n9403_));
  NOR3_X1    g09119(.A1(new_n9393_), .A2(new_n9028_), .A3(new_n9399_), .ZN(new_n9404_));
  NOR2_X1    g09120(.A1(new_n9400_), .A2(new_n9045_), .ZN(new_n9405_));
  NOR3_X1    g09121(.A1(new_n9405_), .A2(new_n9404_), .A3(new_n9029_), .ZN(new_n9406_));
  OAI22_X1   g09122(.A1(new_n7619_), .A2(new_n419_), .B1(new_n420_), .B2(new_n8309_), .ZN(new_n9407_));
  OAI21_X1   g09123(.A1(new_n325_), .A2(new_n7947_), .B(new_n9407_), .ZN(new_n9408_));
  AOI21_X1   g09124(.A1(new_n9408_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n9409_));
  XOR2_X1    g09125(.A1(new_n556_), .A2(new_n9409_), .Z(new_n9410_));
  OAI21_X1   g09126(.A1(new_n9403_), .A2(new_n9406_), .B(new_n9410_), .ZN(new_n9411_));
  AOI21_X1   g09127(.A1(new_n9380_), .A2(new_n9378_), .B(new_n9411_), .ZN(new_n9412_));
  AOI21_X1   g09128(.A1(new_n9054_), .A2(new_n8659_), .B(new_n8623_), .ZN(new_n9413_));
  OAI21_X1   g09129(.A1(new_n9054_), .A2(new_n8659_), .B(new_n8613_), .ZN(new_n9414_));
  INV_X1     g09130(.I(new_n9403_), .ZN(new_n9415_));
  NAND3_X1   g09131(.A1(new_n9401_), .A2(new_n9046_), .A3(new_n9402_), .ZN(new_n9416_));
  XOR2_X1    g09132(.A1(new_n425_), .A2(new_n9409_), .Z(new_n9417_));
  AOI21_X1   g09133(.A1(new_n9415_), .A2(new_n9416_), .B(new_n9417_), .ZN(new_n9418_));
  NOR3_X1    g09134(.A1(new_n9414_), .A2(new_n9418_), .A3(new_n9413_), .ZN(new_n9419_));
  OAI21_X1   g09135(.A1(new_n9419_), .A2(new_n9412_), .B(new_n9376_), .ZN(new_n9420_));
  OAI21_X1   g09136(.A1(new_n9414_), .A2(new_n9413_), .B(new_n9418_), .ZN(new_n9421_));
  NAND3_X1   g09137(.A1(new_n9380_), .A2(new_n9378_), .A3(new_n9411_), .ZN(new_n9422_));
  NAND3_X1   g09138(.A1(new_n9421_), .A2(new_n9422_), .A3(new_n9375_), .ZN(new_n9423_));
  OAI22_X1   g09139(.A1(new_n6644_), .A2(new_n515_), .B1(new_n565_), .B2(new_n6647_), .ZN(new_n9424_));
  OAI21_X1   g09140(.A1(new_n472_), .A2(new_n7284_), .B(new_n9424_), .ZN(new_n9425_));
  AOI21_X1   g09141(.A1(new_n9425_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n9426_));
  XOR2_X1    g09142(.A1(new_n759_), .A2(new_n9426_), .Z(new_n9427_));
  AOI21_X1   g09143(.A1(new_n9420_), .A2(new_n9423_), .B(new_n9427_), .ZN(new_n9428_));
  OAI21_X1   g09144(.A1(new_n9369_), .A2(new_n9371_), .B(new_n9428_), .ZN(new_n9429_));
  OAI21_X1   g09145(.A1(new_n9070_), .A2(new_n9074_), .B(new_n8672_), .ZN(new_n9430_));
  NAND2_X1   g09146(.A1(new_n9430_), .A2(new_n8676_), .ZN(new_n9431_));
  NOR3_X1    g09147(.A1(new_n9070_), .A2(new_n9074_), .A3(new_n8672_), .ZN(new_n9432_));
  NOR2_X1    g09148(.A1(new_n9432_), .A2(new_n8684_), .ZN(new_n9433_));
  AOI21_X1   g09149(.A1(new_n9421_), .A2(new_n9422_), .B(new_n9375_), .ZN(new_n9434_));
  NOR3_X1    g09150(.A1(new_n9419_), .A2(new_n9412_), .A3(new_n9376_), .ZN(new_n9435_));
  INV_X1     g09151(.I(new_n9427_), .ZN(new_n9436_));
  OAI21_X1   g09152(.A1(new_n9435_), .A2(new_n9434_), .B(new_n9436_), .ZN(new_n9437_));
  NAND3_X1   g09153(.A1(new_n9433_), .A2(new_n9431_), .A3(new_n9437_), .ZN(new_n9438_));
  AOI21_X1   g09154(.A1(new_n9438_), .A2(new_n9429_), .B(new_n9074_), .ZN(new_n9439_));
  AOI21_X1   g09155(.A1(new_n9433_), .A2(new_n9431_), .B(new_n9437_), .ZN(new_n9440_));
  NOR3_X1    g09156(.A1(new_n9369_), .A2(new_n9371_), .A3(new_n9428_), .ZN(new_n9441_));
  NOR3_X1    g09157(.A1(new_n9440_), .A2(new_n9441_), .A3(new_n9078_), .ZN(new_n9442_));
  OAI22_X1   g09158(.A1(new_n5993_), .A2(new_n706_), .B1(new_n780_), .B2(new_n5991_), .ZN(new_n9443_));
  OAI21_X1   g09159(.A1(new_n656_), .A2(new_n5997_), .B(new_n9443_), .ZN(new_n9444_));
  AOI21_X1   g09160(.A1(new_n9444_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n9445_));
  XOR2_X1    g09161(.A1(new_n785_), .A2(new_n9445_), .Z(new_n9446_));
  INV_X1     g09162(.I(new_n9446_), .ZN(new_n9447_));
  OAI21_X1   g09163(.A1(new_n9439_), .A2(new_n9442_), .B(new_n9447_), .ZN(new_n9448_));
  AOI21_X1   g09164(.A1(new_n9013_), .A2(new_n9362_), .B(new_n9448_), .ZN(new_n9449_));
  OAI21_X1   g09165(.A1(new_n9440_), .A2(new_n9441_), .B(new_n9078_), .ZN(new_n9450_));
  NAND3_X1   g09166(.A1(new_n9438_), .A2(new_n9429_), .A3(new_n9074_), .ZN(new_n9451_));
  AOI21_X1   g09167(.A1(new_n9450_), .A2(new_n9451_), .B(new_n9446_), .ZN(new_n9452_));
  NOR3_X1    g09168(.A1(new_n9452_), .A2(new_n9113_), .A3(new_n9106_), .ZN(new_n9453_));
  OAI21_X1   g09169(.A1(new_n9449_), .A2(new_n9453_), .B(new_n9368_), .ZN(new_n9454_));
  INV_X1     g09170(.I(new_n9368_), .ZN(new_n9455_));
  OAI21_X1   g09171(.A1(new_n9106_), .A2(new_n9113_), .B(new_n9452_), .ZN(new_n9456_));
  NAND3_X1   g09172(.A1(new_n9448_), .A2(new_n9013_), .A3(new_n9362_), .ZN(new_n9457_));
  NAND3_X1   g09173(.A1(new_n9456_), .A2(new_n9457_), .A3(new_n9455_), .ZN(new_n9458_));
  OAI22_X1   g09174(.A1(new_n5420_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n5107_), .ZN(new_n9459_));
  OAI21_X1   g09175(.A1(new_n861_), .A2(new_n5112_), .B(new_n9459_), .ZN(new_n9460_));
  AOI21_X1   g09176(.A1(new_n9460_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n9461_));
  XOR2_X1    g09177(.A1(new_n1024_), .A2(new_n9461_), .Z(new_n9462_));
  AOI21_X1   g09178(.A1(new_n9454_), .A2(new_n9458_), .B(new_n9462_), .ZN(new_n9463_));
  OAI21_X1   g09179(.A1(new_n9366_), .A2(new_n9367_), .B(new_n9463_), .ZN(new_n9464_));
  INV_X1     g09180(.I(new_n9112_), .ZN(new_n9465_));
  OAI21_X1   g09181(.A1(new_n9110_), .A2(new_n8712_), .B(new_n9465_), .ZN(new_n9466_));
  NOR3_X1    g09182(.A1(new_n9104_), .A2(new_n9109_), .A3(new_n8713_), .ZN(new_n9467_));
  AOI21_X1   g09183(.A1(new_n8721_), .A2(new_n8722_), .B(new_n9467_), .ZN(new_n9468_));
  AOI21_X1   g09184(.A1(new_n9456_), .A2(new_n9457_), .B(new_n9455_), .ZN(new_n9469_));
  NOR3_X1    g09185(.A1(new_n9449_), .A2(new_n9368_), .A3(new_n9453_), .ZN(new_n9470_));
  INV_X1     g09186(.I(new_n9462_), .ZN(new_n9471_));
  OAI21_X1   g09187(.A1(new_n9470_), .A2(new_n9469_), .B(new_n9471_), .ZN(new_n9472_));
  NAND3_X1   g09188(.A1(new_n9472_), .A2(new_n9468_), .A3(new_n9466_), .ZN(new_n9473_));
  AOI21_X1   g09189(.A1(new_n9464_), .A2(new_n9473_), .B(new_n9365_), .ZN(new_n9474_));
  AOI21_X1   g09190(.A1(new_n9466_), .A2(new_n9468_), .B(new_n9472_), .ZN(new_n9475_));
  NOR3_X1    g09191(.A1(new_n9367_), .A2(new_n9463_), .A3(new_n9366_), .ZN(new_n9476_));
  NOR3_X1    g09192(.A1(new_n9475_), .A2(new_n9476_), .A3(new_n9364_), .ZN(new_n9477_));
  OAI22_X1   g09193(.A1(new_n4072_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n4067_), .ZN(new_n9478_));
  OAI21_X1   g09194(.A1(new_n1109_), .A2(new_n4318_), .B(new_n9478_), .ZN(new_n9479_));
  AOI21_X1   g09195(.A1(new_n9479_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n9480_));
  XOR2_X1    g09196(.A1(new_n1299_), .A2(new_n9480_), .Z(new_n9481_));
  INV_X1     g09197(.I(new_n9481_), .ZN(new_n9482_));
  OAI21_X1   g09198(.A1(new_n9477_), .A2(new_n9474_), .B(new_n9482_), .ZN(new_n9483_));
  NOR2_X1    g09199(.A1(new_n9361_), .A2(new_n9483_), .ZN(new_n9484_));
  AOI21_X1   g09200(.A1(new_n9136_), .A2(new_n9133_), .B(new_n8742_), .ZN(new_n9485_));
  OAI21_X1   g09201(.A1(new_n9485_), .A2(new_n8755_), .B(new_n8743_), .ZN(new_n9486_));
  OAI21_X1   g09202(.A1(new_n9475_), .A2(new_n9476_), .B(new_n9364_), .ZN(new_n9487_));
  NAND3_X1   g09203(.A1(new_n9464_), .A2(new_n9473_), .A3(new_n9365_), .ZN(new_n9488_));
  AOI21_X1   g09204(.A1(new_n9487_), .A2(new_n9488_), .B(new_n9481_), .ZN(new_n9489_));
  NOR2_X1    g09205(.A1(new_n9486_), .A2(new_n9489_), .ZN(new_n9490_));
  OAI21_X1   g09206(.A1(new_n9484_), .A2(new_n9490_), .B(new_n9136_), .ZN(new_n9491_));
  NAND2_X1   g09207(.A1(new_n9486_), .A2(new_n9489_), .ZN(new_n9492_));
  NAND2_X1   g09208(.A1(new_n9361_), .A2(new_n9483_), .ZN(new_n9493_));
  NAND3_X1   g09209(.A1(new_n9493_), .A2(new_n9492_), .A3(new_n9140_), .ZN(new_n9494_));
  OAI22_X1   g09210(.A1(new_n1525_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1634_), .ZN(new_n9495_));
  OAI21_X1   g09211(.A1(new_n1518_), .A2(new_n3569_), .B(new_n9495_), .ZN(new_n9496_));
  AOI21_X1   g09212(.A1(new_n9496_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n9497_));
  XNOR2_X1   g09213(.A1(new_n1638_), .A2(new_n9497_), .ZN(new_n9498_));
  AOI21_X1   g09214(.A1(new_n9491_), .A2(new_n9494_), .B(new_n9498_), .ZN(new_n9499_));
  NAND2_X1   g09215(.A1(new_n9359_), .A2(new_n9499_), .ZN(new_n9500_));
  OR2_X2     g09216(.A1(new_n9359_), .A2(new_n9499_), .Z(new_n9501_));
  AOI21_X1   g09217(.A1(new_n9501_), .A2(new_n9500_), .B(new_n9151_), .ZN(new_n9502_));
  INV_X1     g09218(.I(new_n9500_), .ZN(new_n9503_));
  NOR2_X1    g09219(.A1(new_n9359_), .A2(new_n9499_), .ZN(new_n9504_));
  NOR3_X1    g09220(.A1(new_n9503_), .A2(new_n9156_), .A3(new_n9504_), .ZN(new_n9505_));
  OAI22_X1   g09221(.A1(new_n1936_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n2102_), .ZN(new_n9506_));
  OAI21_X1   g09222(.A1(new_n1803_), .A2(new_n2884_), .B(new_n9506_), .ZN(new_n9507_));
  AOI21_X1   g09223(.A1(new_n9507_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n9508_));
  XOR2_X1    g09224(.A1(new_n2106_), .A2(new_n9508_), .Z(new_n9509_));
  INV_X1     g09225(.I(new_n9509_), .ZN(new_n9510_));
  OAI21_X1   g09226(.A1(new_n9505_), .A2(new_n9502_), .B(new_n9510_), .ZN(new_n9511_));
  NOR2_X1    g09227(.A1(new_n9511_), .A2(new_n9357_), .ZN(new_n9512_));
  OAI21_X1   g09228(.A1(new_n9158_), .A2(new_n9153_), .B(new_n9009_), .ZN(new_n9513_));
  NAND3_X1   g09229(.A1(new_n9353_), .A2(new_n9352_), .A3(new_n9008_), .ZN(new_n9514_));
  AOI21_X1   g09230(.A1(new_n9513_), .A2(new_n9514_), .B(new_n8786_), .ZN(new_n9515_));
  OAI21_X1   g09231(.A1(new_n8792_), .A2(new_n9515_), .B(new_n8787_), .ZN(new_n9516_));
  OAI21_X1   g09232(.A1(new_n9503_), .A2(new_n9504_), .B(new_n9156_), .ZN(new_n9517_));
  NAND3_X1   g09233(.A1(new_n9501_), .A2(new_n9151_), .A3(new_n9500_), .ZN(new_n9518_));
  AOI21_X1   g09234(.A1(new_n9517_), .A2(new_n9518_), .B(new_n9509_), .ZN(new_n9519_));
  NOR2_X1    g09235(.A1(new_n9519_), .A2(new_n9516_), .ZN(new_n9520_));
  OAI21_X1   g09236(.A1(new_n9512_), .A2(new_n9520_), .B(new_n9350_), .ZN(new_n9521_));
  NAND2_X1   g09237(.A1(new_n9519_), .A2(new_n9516_), .ZN(new_n9522_));
  NAND2_X1   g09238(.A1(new_n9511_), .A2(new_n9357_), .ZN(new_n9523_));
  NAND3_X1   g09239(.A1(new_n9523_), .A2(new_n9522_), .A3(new_n9349_), .ZN(new_n9524_));
  OAI22_X1   g09240(.A1(new_n2171_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n2166_), .ZN(new_n9525_));
  OAI21_X1   g09241(.A1(new_n2281_), .A2(new_n2322_), .B(new_n9525_), .ZN(new_n9526_));
  AOI21_X1   g09242(.A1(new_n9526_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n9527_));
  XNOR2_X1   g09243(.A1(new_n2647_), .A2(new_n9527_), .ZN(new_n9528_));
  AOI21_X1   g09244(.A1(new_n9521_), .A2(new_n9524_), .B(new_n9528_), .ZN(new_n9529_));
  NAND2_X1   g09245(.A1(new_n9348_), .A2(new_n9529_), .ZN(new_n9530_));
  OAI21_X1   g09246(.A1(new_n9181_), .A2(new_n9178_), .B(new_n8804_), .ZN(new_n9531_));
  AOI21_X1   g09247(.A1(new_n9531_), .A2(new_n8816_), .B(new_n8805_), .ZN(new_n9532_));
  INV_X1     g09248(.I(new_n9529_), .ZN(new_n9533_));
  NAND2_X1   g09249(.A1(new_n9532_), .A2(new_n9533_), .ZN(new_n9534_));
  AOI21_X1   g09250(.A1(new_n9534_), .A2(new_n9530_), .B(new_n9346_), .ZN(new_n9535_));
  INV_X1     g09251(.I(new_n9346_), .ZN(new_n9536_));
  NOR2_X1    g09252(.A1(new_n9532_), .A2(new_n9533_), .ZN(new_n9537_));
  NOR2_X1    g09253(.A1(new_n9348_), .A2(new_n9529_), .ZN(new_n9538_));
  NOR3_X1    g09254(.A1(new_n9537_), .A2(new_n9538_), .A3(new_n9536_), .ZN(new_n9539_));
  OAI22_X1   g09255(.A1(new_n1712_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n1707_), .ZN(new_n9540_));
  OAI21_X1   g09256(.A1(new_n2842_), .A2(new_n1850_), .B(new_n9540_), .ZN(new_n9541_));
  AOI21_X1   g09257(.A1(new_n9541_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n9542_));
  XNOR2_X1   g09258(.A1(new_n3264_), .A2(new_n9542_), .ZN(new_n9543_));
  INV_X1     g09259(.I(new_n9543_), .ZN(new_n9544_));
  OAI21_X1   g09260(.A1(new_n9535_), .A2(new_n9539_), .B(new_n9544_), .ZN(new_n9545_));
  NOR2_X1    g09261(.A1(new_n9545_), .A2(new_n9340_), .ZN(new_n9546_));
  NAND2_X1   g09262(.A1(new_n8826_), .A2(new_n8823_), .ZN(new_n9547_));
  NAND2_X1   g09263(.A1(new_n8588_), .A2(new_n9547_), .ZN(new_n9548_));
  OAI21_X1   g09264(.A1(new_n9537_), .A2(new_n9538_), .B(new_n9536_), .ZN(new_n9549_));
  NAND3_X1   g09265(.A1(new_n9534_), .A2(new_n9530_), .A3(new_n9346_), .ZN(new_n9550_));
  NAND2_X1   g09266(.A1(new_n9549_), .A2(new_n9550_), .ZN(new_n9551_));
  AOI21_X1   g09267(.A1(new_n9551_), .A2(new_n9544_), .B(new_n9548_), .ZN(new_n9552_));
  OAI21_X1   g09268(.A1(new_n9546_), .A2(new_n9552_), .B(new_n9338_), .ZN(new_n9553_));
  NAND3_X1   g09269(.A1(new_n9551_), .A2(new_n9548_), .A3(new_n9544_), .ZN(new_n9554_));
  NAND2_X1   g09270(.A1(new_n9545_), .A2(new_n9340_), .ZN(new_n9555_));
  NAND3_X1   g09271(.A1(new_n9555_), .A2(new_n9554_), .A3(new_n9337_), .ZN(new_n9556_));
  OAI22_X1   g09272(.A1(new_n1347_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n1344_), .ZN(new_n9557_));
  OAI21_X1   g09273(.A1(new_n3709_), .A2(new_n1457_), .B(new_n9557_), .ZN(new_n9558_));
  AOI21_X1   g09274(.A1(new_n9558_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n9559_));
  XNOR2_X1   g09275(.A1(new_n3993_), .A2(new_n9559_), .ZN(new_n9560_));
  AOI21_X1   g09276(.A1(new_n9553_), .A2(new_n9556_), .B(new_n9560_), .ZN(new_n9561_));
  NAND2_X1   g09277(.A1(new_n9336_), .A2(new_n9561_), .ZN(new_n9562_));
  OAI21_X1   g09278(.A1(new_n9212_), .A2(new_n9208_), .B(new_n8841_), .ZN(new_n9563_));
  AOI21_X1   g09279(.A1(new_n9563_), .A2(new_n8853_), .B(new_n8842_), .ZN(new_n9564_));
  AOI21_X1   g09280(.A1(new_n9555_), .A2(new_n9554_), .B(new_n9337_), .ZN(new_n9565_));
  NOR3_X1    g09281(.A1(new_n9546_), .A2(new_n9552_), .A3(new_n9338_), .ZN(new_n9566_));
  INV_X1     g09282(.I(new_n9560_), .ZN(new_n9567_));
  OAI21_X1   g09283(.A1(new_n9566_), .A2(new_n9565_), .B(new_n9567_), .ZN(new_n9568_));
  NAND2_X1   g09284(.A1(new_n9564_), .A2(new_n9568_), .ZN(new_n9569_));
  AOI21_X1   g09285(.A1(new_n9569_), .A2(new_n9562_), .B(new_n9334_), .ZN(new_n9570_));
  INV_X1     g09286(.I(new_n9334_), .ZN(new_n9571_));
  NOR2_X1    g09287(.A1(new_n9564_), .A2(new_n9568_), .ZN(new_n9572_));
  NOR2_X1    g09288(.A1(new_n9336_), .A2(new_n9561_), .ZN(new_n9573_));
  NOR3_X1    g09289(.A1(new_n9572_), .A2(new_n9573_), .A3(new_n9571_), .ZN(new_n9574_));
  OAI22_X1   g09290(.A1(new_n1055_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n1061_), .ZN(new_n9575_));
  OAI21_X1   g09291(.A1(new_n4253_), .A2(new_n1332_), .B(new_n9575_), .ZN(new_n9576_));
  AOI21_X1   g09292(.A1(new_n9576_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n9577_));
  XNOR2_X1   g09293(.A1(new_n4778_), .A2(new_n9577_), .ZN(new_n9578_));
  INV_X1     g09294(.I(new_n9578_), .ZN(new_n9579_));
  OAI21_X1   g09295(.A1(new_n9570_), .A2(new_n9574_), .B(new_n9579_), .ZN(new_n9580_));
  NOR2_X1    g09296(.A1(new_n9333_), .A2(new_n9580_), .ZN(new_n9581_));
  AOI21_X1   g09297(.A1(new_n9231_), .A2(new_n9230_), .B(new_n8863_), .ZN(new_n9582_));
  OAI21_X1   g09298(.A1(new_n9582_), .A2(new_n8877_), .B(new_n8864_), .ZN(new_n9583_));
  OAI21_X1   g09299(.A1(new_n9572_), .A2(new_n9573_), .B(new_n9571_), .ZN(new_n9584_));
  NAND3_X1   g09300(.A1(new_n9569_), .A2(new_n9562_), .A3(new_n9334_), .ZN(new_n9585_));
  AOI21_X1   g09301(.A1(new_n9584_), .A2(new_n9585_), .B(new_n9578_), .ZN(new_n9586_));
  NOR2_X1    g09302(.A1(new_n9583_), .A2(new_n9586_), .ZN(new_n9587_));
  OAI21_X1   g09303(.A1(new_n9581_), .A2(new_n9587_), .B(new_n9231_), .ZN(new_n9588_));
  NAND2_X1   g09304(.A1(new_n9583_), .A2(new_n9586_), .ZN(new_n9589_));
  NAND2_X1   g09305(.A1(new_n9333_), .A2(new_n9580_), .ZN(new_n9590_));
  NAND3_X1   g09306(.A1(new_n9590_), .A2(new_n9589_), .A3(new_n9227_), .ZN(new_n9591_));
  OAI22_X1   g09307(.A1(new_n970_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n820_), .ZN(new_n9592_));
  OAI21_X1   g09308(.A1(new_n5068_), .A2(new_n894_), .B(new_n9592_), .ZN(new_n9593_));
  AOI21_X1   g09309(.A1(new_n9593_), .A2(new_n827_), .B(new_n970_), .ZN(new_n9594_));
  XNOR2_X1   g09310(.A1(new_n5600_), .A2(new_n9594_), .ZN(new_n9595_));
  AOI21_X1   g09311(.A1(new_n9588_), .A2(new_n9591_), .B(new_n9595_), .ZN(new_n9596_));
  NAND2_X1   g09312(.A1(new_n9331_), .A2(new_n9596_), .ZN(new_n9597_));
  OAI21_X1   g09313(.A1(new_n9238_), .A2(new_n9242_), .B(new_n8887_), .ZN(new_n9598_));
  AOI21_X1   g09314(.A1(new_n8899_), .A2(new_n9598_), .B(new_n8888_), .ZN(new_n9599_));
  AOI21_X1   g09315(.A1(new_n9590_), .A2(new_n9589_), .B(new_n9227_), .ZN(new_n9600_));
  NOR3_X1    g09316(.A1(new_n9581_), .A2(new_n9587_), .A3(new_n9231_), .ZN(new_n9601_));
  INV_X1     g09317(.I(new_n9595_), .ZN(new_n9602_));
  OAI21_X1   g09318(.A1(new_n9600_), .A2(new_n9601_), .B(new_n9602_), .ZN(new_n9603_));
  NAND2_X1   g09319(.A1(new_n9599_), .A2(new_n9603_), .ZN(new_n9604_));
  AOI21_X1   g09320(.A1(new_n9597_), .A2(new_n9604_), .B(new_n9242_), .ZN(new_n9605_));
  NOR2_X1    g09321(.A1(new_n9599_), .A2(new_n9603_), .ZN(new_n9606_));
  NOR2_X1    g09322(.A1(new_n9331_), .A2(new_n9596_), .ZN(new_n9607_));
  NOR3_X1    g09323(.A1(new_n9607_), .A2(new_n9606_), .A3(new_n9247_), .ZN(new_n9608_));
  OAI22_X1   g09324(.A1(new_n607_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n610_), .ZN(new_n9609_));
  OAI21_X1   g09325(.A1(new_n5921_), .A2(new_n684_), .B(new_n9609_), .ZN(new_n9610_));
  AOI21_X1   g09326(.A1(new_n9610_), .A2(new_n612_), .B(new_n607_), .ZN(new_n9611_));
  XOR2_X1    g09327(.A1(new_n6543_), .A2(new_n9611_), .Z(new_n9612_));
  INV_X1     g09328(.I(new_n9612_), .ZN(new_n9613_));
  OAI21_X1   g09329(.A1(new_n9605_), .A2(new_n9608_), .B(new_n9613_), .ZN(new_n9614_));
  AOI21_X1   g09330(.A1(new_n9329_), .A2(new_n8910_), .B(new_n9614_), .ZN(new_n9615_));
  AOI21_X1   g09331(.A1(new_n9262_), .A2(new_n9261_), .B(new_n8909_), .ZN(new_n9616_));
  OAI21_X1   g09332(.A1(new_n8915_), .A2(new_n9616_), .B(new_n8910_), .ZN(new_n9617_));
  INV_X1     g09333(.I(new_n9614_), .ZN(new_n9618_));
  NOR2_X1    g09334(.A1(new_n9618_), .A2(new_n9617_), .ZN(new_n9619_));
  OAI21_X1   g09335(.A1(new_n9619_), .A2(new_n9615_), .B(new_n9262_), .ZN(new_n9620_));
  NAND2_X1   g09336(.A1(new_n9618_), .A2(new_n9617_), .ZN(new_n9621_));
  NAND3_X1   g09337(.A1(new_n9329_), .A2(new_n9614_), .A3(new_n8910_), .ZN(new_n9622_));
  NAND3_X1   g09338(.A1(new_n9621_), .A2(new_n9622_), .A3(new_n9258_), .ZN(new_n9623_));
  NAND2_X1   g09339(.A1(new_n9620_), .A2(new_n9623_), .ZN(new_n9624_));
  OAI22_X1   g09340(.A1(new_n448_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n450_), .ZN(new_n9625_));
  OAI21_X1   g09341(.A1(new_n6847_), .A2(new_n496_), .B(new_n9625_), .ZN(new_n9626_));
  AOI21_X1   g09342(.A1(new_n9626_), .A2(new_n452_), .B(new_n448_), .ZN(new_n9627_));
  XOR2_X1    g09343(.A1(new_n7516_), .A2(new_n9627_), .Z(new_n9628_));
  INV_X1     g09344(.I(new_n9628_), .ZN(new_n9629_));
  XOR2_X1    g09345(.A1(new_n9624_), .A2(new_n9629_), .Z(new_n9630_));
  OAI22_X1   g09346(.A1(new_n8218_), .A2(new_n341_), .B1(new_n404_), .B2(new_n8563_), .ZN(new_n9631_));
  OAI21_X1   g09347(.A1(new_n7870_), .A2(new_n366_), .B(new_n9631_), .ZN(new_n9632_));
  AOI21_X1   g09348(.A1(new_n9632_), .A2(new_n334_), .B(new_n341_), .ZN(new_n9633_));
  XOR2_X1    g09349(.A1(new_n8568_), .A2(new_n9633_), .Z(new_n9634_));
  INV_X1     g09350(.I(new_n9634_), .ZN(new_n9635_));
  XOR2_X1    g09351(.A1(new_n9630_), .A2(new_n9635_), .Z(new_n9636_));
  NAND2_X1   g09352(.A1(new_n9636_), .A2(new_n9326_), .ZN(new_n9637_));
  XOR2_X1    g09353(.A1(new_n9630_), .A2(new_n9635_), .Z(new_n9638_));
  OAI21_X1   g09354(.A1(new_n9326_), .A2(new_n9638_), .B(new_n9637_), .ZN(new_n9639_));
  XNOR2_X1   g09355(.A1(\b[49] ), .A2(\b[51] ), .ZN(new_n9640_));
  NOR2_X1    g09356(.A1(new_n9640_), .A2(new_n9294_), .ZN(new_n9641_));
  XNOR2_X1   g09357(.A1(new_n9293_), .A2(new_n9641_), .ZN(new_n9642_));
  NAND2_X1   g09358(.A1(new_n286_), .A2(\b[50] ), .ZN(new_n9643_));
  AOI22_X1   g09359(.A1(new_n304_), .A2(\b[49] ), .B1(new_n262_), .B2(\b[51] ), .ZN(new_n9644_));
  AOI21_X1   g09360(.A1(new_n9643_), .A2(new_n9644_), .B(new_n426_), .ZN(new_n9645_));
  NAND2_X1   g09361(.A1(new_n9642_), .A2(new_n9645_), .ZN(new_n9646_));
  XOR2_X1    g09362(.A1(new_n9646_), .A2(\a[2] ), .Z(new_n9647_));
  INV_X1     g09363(.I(new_n9647_), .ZN(new_n9648_));
  NAND2_X1   g09364(.A1(new_n9639_), .A2(new_n9648_), .ZN(new_n9649_));
  NOR2_X1    g09365(.A1(new_n9638_), .A2(new_n9326_), .ZN(new_n9650_));
  AOI21_X1   g09366(.A1(new_n9326_), .A2(new_n9636_), .B(new_n9650_), .ZN(new_n9651_));
  NAND2_X1   g09367(.A1(new_n9651_), .A2(new_n9647_), .ZN(new_n9652_));
  AOI21_X1   g09368(.A1(new_n9652_), .A2(new_n9649_), .B(new_n9321_), .ZN(new_n9653_));
  NAND2_X1   g09369(.A1(new_n9651_), .A2(new_n9648_), .ZN(new_n9654_));
  NAND2_X1   g09370(.A1(new_n9639_), .A2(new_n9647_), .ZN(new_n9655_));
  AOI21_X1   g09371(.A1(new_n9654_), .A2(new_n9655_), .B(new_n9320_), .ZN(new_n9656_));
  OAI21_X1   g09372(.A1(new_n9653_), .A2(new_n9656_), .B(new_n9308_), .ZN(new_n9657_));
  XOR2_X1    g09373(.A1(new_n9657_), .A2(new_n9305_), .Z(new_n9658_));
  XOR2_X1    g09374(.A1(new_n9658_), .A2(new_n8979_), .Z(\f[51] ));
  NOR2_X1    g09375(.A1(new_n9321_), .A2(new_n9634_), .ZN(new_n9660_));
  XOR2_X1    g09376(.A1(new_n9630_), .A2(new_n9325_), .Z(new_n9661_));
  AOI21_X1   g09377(.A1(new_n9321_), .A2(new_n9634_), .B(new_n9661_), .ZN(new_n9662_));
  OAI21_X1   g09378(.A1(new_n9607_), .A2(new_n9606_), .B(new_n9247_), .ZN(new_n9663_));
  NAND3_X1   g09379(.A1(new_n9597_), .A2(new_n9604_), .A3(new_n9242_), .ZN(new_n9664_));
  AOI21_X1   g09380(.A1(new_n9663_), .A2(new_n9664_), .B(new_n9262_), .ZN(new_n9665_));
  INV_X1     g09381(.I(new_n9665_), .ZN(new_n9666_));
  NAND3_X1   g09382(.A1(new_n9663_), .A2(new_n9664_), .A3(new_n9262_), .ZN(new_n9667_));
  NAND4_X1   g09383(.A1(new_n9329_), .A2(new_n9667_), .A3(new_n8910_), .A4(new_n9613_), .ZN(new_n9668_));
  NAND2_X1   g09384(.A1(new_n9668_), .A2(new_n9666_), .ZN(new_n9669_));
  AOI21_X1   g09385(.A1(new_n9588_), .A2(new_n9591_), .B(new_n9247_), .ZN(new_n9670_));
  NOR3_X1    g09386(.A1(new_n9600_), .A2(new_n9601_), .A3(new_n9242_), .ZN(new_n9671_));
  NOR2_X1    g09387(.A1(new_n9671_), .A2(new_n9595_), .ZN(new_n9672_));
  AOI21_X1   g09388(.A1(new_n9672_), .A2(new_n9599_), .B(new_n9670_), .ZN(new_n9673_));
  NOR2_X1    g09389(.A1(new_n9570_), .A2(new_n9574_), .ZN(new_n9674_));
  NAND3_X1   g09390(.A1(new_n9584_), .A2(new_n9585_), .A3(new_n9231_), .ZN(new_n9675_));
  NAND2_X1   g09391(.A1(new_n9675_), .A2(new_n9579_), .ZN(new_n9676_));
  OAI22_X1   g09392(.A1(new_n9676_), .A2(new_n9583_), .B1(new_n9231_), .B2(new_n9674_), .ZN(new_n9677_));
  NOR2_X1    g09393(.A1(new_n9566_), .A2(new_n9565_), .ZN(new_n9678_));
  NAND3_X1   g09394(.A1(new_n9553_), .A2(new_n9556_), .A3(new_n9571_), .ZN(new_n9679_));
  NAND2_X1   g09395(.A1(new_n9679_), .A2(new_n9567_), .ZN(new_n9680_));
  OAI22_X1   g09396(.A1(new_n9680_), .A2(new_n9336_), .B1(new_n9571_), .B2(new_n9678_), .ZN(new_n9681_));
  AOI21_X1   g09397(.A1(new_n9549_), .A2(new_n9550_), .B(new_n9338_), .ZN(new_n9682_));
  INV_X1     g09398(.I(new_n9682_), .ZN(new_n9683_));
  NAND3_X1   g09399(.A1(new_n9549_), .A2(new_n9550_), .A3(new_n9338_), .ZN(new_n9684_));
  NAND3_X1   g09400(.A1(new_n9340_), .A2(new_n9684_), .A3(new_n9544_), .ZN(new_n9685_));
  NAND2_X1   g09401(.A1(new_n9685_), .A2(new_n9683_), .ZN(new_n9686_));
  NAND2_X1   g09402(.A1(new_n9521_), .A2(new_n9524_), .ZN(new_n9687_));
  INV_X1     g09403(.I(new_n9687_), .ZN(new_n9688_));
  INV_X1     g09404(.I(new_n9528_), .ZN(new_n9689_));
  OAI21_X1   g09405(.A1(new_n9687_), .A2(new_n9346_), .B(new_n9689_), .ZN(new_n9690_));
  OAI22_X1   g09406(.A1(new_n9348_), .A2(new_n9690_), .B1(new_n9536_), .B2(new_n9688_), .ZN(new_n9691_));
  AOI21_X1   g09407(.A1(new_n9517_), .A2(new_n9518_), .B(new_n9350_), .ZN(new_n9692_));
  NOR3_X1    g09408(.A1(new_n9505_), .A2(new_n9502_), .A3(new_n9349_), .ZN(new_n9693_));
  NOR3_X1    g09409(.A1(new_n9693_), .A2(new_n9516_), .A3(new_n9509_), .ZN(new_n9694_));
  OAI21_X1   g09410(.A1(new_n9477_), .A2(new_n9474_), .B(new_n9140_), .ZN(new_n9695_));
  NAND3_X1   g09411(.A1(new_n9487_), .A2(new_n9488_), .A3(new_n9136_), .ZN(new_n9696_));
  NAND2_X1   g09412(.A1(new_n9696_), .A2(new_n9482_), .ZN(new_n9697_));
  OAI21_X1   g09413(.A1(new_n9697_), .A2(new_n9486_), .B(new_n9695_), .ZN(new_n9698_));
  AOI21_X1   g09414(.A1(new_n9450_), .A2(new_n9451_), .B(new_n9368_), .ZN(new_n9699_));
  NAND3_X1   g09415(.A1(new_n9450_), .A2(new_n9451_), .A3(new_n9368_), .ZN(new_n9700_));
  NOR3_X1    g09416(.A1(new_n9113_), .A2(new_n9106_), .A3(new_n9446_), .ZN(new_n9701_));
  AOI21_X1   g09417(.A1(new_n9701_), .A2(new_n9700_), .B(new_n9699_), .ZN(new_n9702_));
  NAND2_X1   g09418(.A1(new_n9420_), .A2(new_n9423_), .ZN(new_n9703_));
  NAND2_X1   g09419(.A1(new_n9703_), .A2(new_n9074_), .ZN(new_n9704_));
  NAND3_X1   g09420(.A1(new_n9420_), .A2(new_n9423_), .A3(new_n9078_), .ZN(new_n9705_));
  NAND4_X1   g09421(.A1(new_n9433_), .A2(new_n9431_), .A3(new_n9436_), .A4(new_n9705_), .ZN(new_n9706_));
  AOI21_X1   g09422(.A1(new_n9415_), .A2(new_n9416_), .B(new_n9376_), .ZN(new_n9707_));
  NOR3_X1    g09423(.A1(new_n9406_), .A2(new_n9403_), .A3(new_n9375_), .ZN(new_n9708_));
  NOR4_X1    g09424(.A1(new_n9414_), .A2(new_n9413_), .A3(new_n9417_), .A4(new_n9708_), .ZN(new_n9709_));
  NOR2_X1    g09425(.A1(new_n9709_), .A2(new_n9707_), .ZN(new_n9710_));
  XNOR2_X1   g09426(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n9711_));
  NOR2_X1    g09427(.A1(new_n9397_), .A2(new_n9711_), .ZN(new_n9712_));
  INV_X1     g09428(.I(new_n9712_), .ZN(new_n9713_));
  NAND2_X1   g09429(.A1(new_n9395_), .A2(\a[52] ), .ZN(new_n9714_));
  OAI21_X1   g09430(.A1(\a[52] ), .A2(new_n9394_), .B(new_n9714_), .ZN(new_n9715_));
  XOR2_X1    g09431(.A1(\a[52] ), .A2(\a[53] ), .Z(new_n9716_));
  NOR2_X1    g09432(.A1(new_n9397_), .A2(new_n9716_), .ZN(new_n9717_));
  INV_X1     g09433(.I(\a[53] ), .ZN(new_n9718_));
  NAND2_X1   g09434(.A1(new_n268_), .A2(new_n9718_), .ZN(new_n9719_));
  AOI21_X1   g09435(.A1(new_n9717_), .A2(new_n9715_), .B(new_n9719_), .ZN(new_n9720_));
  NOR3_X1    g09436(.A1(new_n9720_), .A2(new_n271_), .A3(new_n9713_), .ZN(new_n9721_));
  INV_X1     g09437(.I(new_n9721_), .ZN(new_n9722_));
  OAI21_X1   g09438(.A1(new_n9720_), .A2(new_n9713_), .B(new_n271_), .ZN(new_n9723_));
  NAND2_X1   g09439(.A1(new_n9722_), .A2(new_n9723_), .ZN(new_n9724_));
  NOR2_X1    g09440(.A1(new_n9398_), .A2(new_n9718_), .ZN(new_n9725_));
  XOR2_X1    g09441(.A1(new_n9724_), .A2(new_n9725_), .Z(new_n9726_));
  NOR2_X1    g09442(.A1(new_n9045_), .A2(new_n9393_), .ZN(new_n9727_));
  NAND4_X1   g09443(.A1(new_n8652_), .A2(new_n8639_), .A3(new_n8653_), .A4(new_n9398_), .ZN(new_n9728_));
  AOI21_X1   g09444(.A1(new_n9045_), .A2(new_n9393_), .B(new_n9728_), .ZN(new_n9729_));
  OAI22_X1   g09445(.A1(new_n8644_), .A2(new_n298_), .B1(new_n325_), .B2(new_n9388_), .ZN(new_n9730_));
  NOR3_X1    g09446(.A1(new_n8313_), .A2(new_n8649_), .A3(new_n9017_), .ZN(new_n9731_));
  NAND2_X1   g09447(.A1(new_n9731_), .A2(\b[2] ), .ZN(new_n9732_));
  NAND2_X1   g09448(.A1(new_n9732_), .A2(new_n9730_), .ZN(new_n9733_));
  AOI21_X1   g09449(.A1(new_n329_), .A2(new_n8631_), .B(new_n9733_), .ZN(new_n9734_));
  INV_X1     g09450(.I(new_n9734_), .ZN(new_n9735_));
  NOR3_X1    g09451(.A1(new_n9729_), .A2(new_n9727_), .A3(new_n9735_), .ZN(new_n9736_));
  OAI21_X1   g09452(.A1(new_n9390_), .A2(new_n9391_), .B(\a[50] ), .ZN(new_n9737_));
  NAND3_X1   g09453(.A1(new_n9384_), .A2(new_n8624_), .A3(new_n9385_), .ZN(new_n9738_));
  NAND2_X1   g09454(.A1(new_n9737_), .A2(new_n9738_), .ZN(new_n9739_));
  NAND2_X1   g09455(.A1(new_n9028_), .A2(new_n9739_), .ZN(new_n9740_));
  NOR4_X1    g09456(.A1(new_n8656_), .A2(new_n8657_), .A3(new_n8654_), .A4(new_n9399_), .ZN(new_n9741_));
  OAI21_X1   g09457(.A1(new_n9028_), .A2(new_n9739_), .B(new_n9741_), .ZN(new_n9742_));
  AOI21_X1   g09458(.A1(new_n9742_), .A2(new_n9740_), .B(new_n9734_), .ZN(new_n9743_));
  OAI21_X1   g09459(.A1(new_n9736_), .A2(new_n9743_), .B(new_n9726_), .ZN(new_n9744_));
  INV_X1     g09460(.I(new_n9725_), .ZN(new_n9745_));
  XOR2_X1    g09461(.A1(new_n9724_), .A2(new_n9745_), .Z(new_n9746_));
  NAND3_X1   g09462(.A1(new_n9742_), .A2(new_n9740_), .A3(new_n9734_), .ZN(new_n9747_));
  OAI21_X1   g09463(.A1(new_n9729_), .A2(new_n9727_), .B(new_n9735_), .ZN(new_n9748_));
  NAND3_X1   g09464(.A1(new_n9748_), .A2(new_n9747_), .A3(new_n9746_), .ZN(new_n9749_));
  AOI21_X1   g09465(.A1(new_n9744_), .A2(new_n9749_), .B(\a[50] ), .ZN(new_n9750_));
  AOI21_X1   g09466(.A1(new_n9748_), .A2(new_n9747_), .B(new_n9746_), .ZN(new_n9751_));
  NOR3_X1    g09467(.A1(new_n9736_), .A2(new_n9743_), .A3(new_n9726_), .ZN(new_n9752_));
  NOR3_X1    g09468(.A1(new_n9752_), .A2(new_n9751_), .A3(new_n8624_), .ZN(new_n9753_));
  OAI22_X1   g09469(.A1(new_n7619_), .A2(new_n420_), .B1(new_n472_), .B2(new_n8309_), .ZN(new_n9754_));
  OAI21_X1   g09470(.A1(new_n419_), .A2(new_n7947_), .B(new_n9754_), .ZN(new_n9755_));
  AOI21_X1   g09471(.A1(new_n9755_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n9756_));
  XOR2_X1    g09472(.A1(new_n471_), .A2(new_n9756_), .Z(new_n9757_));
  INV_X1     g09473(.I(new_n9757_), .ZN(new_n9758_));
  OAI21_X1   g09474(.A1(new_n9753_), .A2(new_n9750_), .B(new_n9758_), .ZN(new_n9759_));
  OAI21_X1   g09475(.A1(new_n9752_), .A2(new_n9751_), .B(new_n8624_), .ZN(new_n9760_));
  NAND3_X1   g09476(.A1(new_n9744_), .A2(new_n9749_), .A3(\a[50] ), .ZN(new_n9761_));
  NAND3_X1   g09477(.A1(new_n9760_), .A2(new_n9761_), .A3(new_n9757_), .ZN(new_n9762_));
  AOI21_X1   g09478(.A1(new_n9759_), .A2(new_n9762_), .B(new_n9710_), .ZN(new_n9763_));
  INV_X1     g09479(.I(new_n9707_), .ZN(new_n9764_));
  NOR2_X1    g09480(.A1(new_n9708_), .A2(new_n9417_), .ZN(new_n9765_));
  NAND3_X1   g09481(.A1(new_n9765_), .A2(new_n9378_), .A3(new_n9380_), .ZN(new_n9766_));
  NAND2_X1   g09482(.A1(new_n9766_), .A2(new_n9764_), .ZN(new_n9767_));
  NOR3_X1    g09483(.A1(new_n9753_), .A2(new_n9750_), .A3(new_n9757_), .ZN(new_n9768_));
  INV_X1     g09484(.I(new_n9768_), .ZN(new_n9769_));
  OAI21_X1   g09485(.A1(new_n9753_), .A2(new_n9750_), .B(new_n9757_), .ZN(new_n9770_));
  AOI21_X1   g09486(.A1(new_n9769_), .A2(new_n9770_), .B(new_n9767_), .ZN(new_n9771_));
  OAI22_X1   g09487(.A1(new_n6644_), .A2(new_n565_), .B1(new_n656_), .B2(new_n6647_), .ZN(new_n9772_));
  OAI21_X1   g09488(.A1(new_n515_), .A2(new_n7284_), .B(new_n9772_), .ZN(new_n9773_));
  AOI21_X1   g09489(.A1(new_n9773_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n9774_));
  XNOR2_X1   g09490(.A1(new_n660_), .A2(new_n9774_), .ZN(new_n9775_));
  NOR3_X1    g09491(.A1(new_n9763_), .A2(new_n9771_), .A3(new_n9775_), .ZN(new_n9776_));
  INV_X1     g09492(.I(new_n9776_), .ZN(new_n9777_));
  NAND2_X1   g09493(.A1(new_n9759_), .A2(new_n9762_), .ZN(new_n9778_));
  NAND2_X1   g09494(.A1(new_n9767_), .A2(new_n9778_), .ZN(new_n9779_));
  AOI21_X1   g09495(.A1(new_n9760_), .A2(new_n9761_), .B(new_n9758_), .ZN(new_n9780_));
  OAI21_X1   g09496(.A1(new_n9768_), .A2(new_n9780_), .B(new_n9710_), .ZN(new_n9781_));
  INV_X1     g09497(.I(new_n9775_), .ZN(new_n9782_));
  AOI21_X1   g09498(.A1(new_n9781_), .A2(new_n9779_), .B(new_n9782_), .ZN(new_n9783_));
  INV_X1     g09499(.I(new_n9783_), .ZN(new_n9784_));
  AOI22_X1   g09500(.A1(new_n9706_), .A2(new_n9704_), .B1(new_n9777_), .B2(new_n9784_), .ZN(new_n9785_));
  INV_X1     g09501(.I(new_n9704_), .ZN(new_n9786_));
  NAND2_X1   g09502(.A1(new_n9705_), .A2(new_n9436_), .ZN(new_n9787_));
  NOR3_X1    g09503(.A1(new_n9787_), .A2(new_n9369_), .A3(new_n9371_), .ZN(new_n9788_));
  AOI21_X1   g09504(.A1(new_n9781_), .A2(new_n9779_), .B(new_n9775_), .ZN(new_n9789_));
  NOR3_X1    g09505(.A1(new_n9763_), .A2(new_n9771_), .A3(new_n9782_), .ZN(new_n9790_));
  NOR2_X1    g09506(.A1(new_n9790_), .A2(new_n9789_), .ZN(new_n9791_));
  NOR3_X1    g09507(.A1(new_n9791_), .A2(new_n9788_), .A3(new_n9786_), .ZN(new_n9792_));
  OAI22_X1   g09508(.A1(new_n5993_), .A2(new_n780_), .B1(new_n861_), .B2(new_n5991_), .ZN(new_n9793_));
  OAI21_X1   g09509(.A1(new_n706_), .A2(new_n5997_), .B(new_n9793_), .ZN(new_n9794_));
  AOI21_X1   g09510(.A1(new_n9794_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n9795_));
  XNOR2_X1   g09511(.A1(new_n860_), .A2(new_n9795_), .ZN(new_n9796_));
  NOR3_X1    g09512(.A1(new_n9785_), .A2(new_n9792_), .A3(new_n9796_), .ZN(new_n9797_));
  OAI22_X1   g09513(.A1(new_n9788_), .A2(new_n9786_), .B1(new_n9776_), .B2(new_n9783_), .ZN(new_n9798_));
  INV_X1     g09514(.I(new_n9792_), .ZN(new_n9799_));
  INV_X1     g09515(.I(new_n9796_), .ZN(new_n9800_));
  AOI21_X1   g09516(.A1(new_n9799_), .A2(new_n9798_), .B(new_n9800_), .ZN(new_n9801_));
  NOR2_X1    g09517(.A1(new_n9801_), .A2(new_n9797_), .ZN(new_n9802_));
  OAI22_X1   g09518(.A1(new_n5420_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n5107_), .ZN(new_n9803_));
  OAI21_X1   g09519(.A1(new_n930_), .A2(new_n5112_), .B(new_n9803_), .ZN(new_n9804_));
  AOI21_X1   g09520(.A1(new_n9804_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n9805_));
  XOR2_X1    g09521(.A1(new_n1114_), .A2(new_n9805_), .Z(new_n9806_));
  INV_X1     g09522(.I(new_n9806_), .ZN(new_n9807_));
  NAND2_X1   g09523(.A1(new_n9802_), .A2(new_n9807_), .ZN(new_n9808_));
  NAND3_X1   g09524(.A1(new_n9799_), .A2(new_n9798_), .A3(new_n9800_), .ZN(new_n9809_));
  OAI21_X1   g09525(.A1(new_n9785_), .A2(new_n9792_), .B(new_n9796_), .ZN(new_n9810_));
  NAND2_X1   g09526(.A1(new_n9809_), .A2(new_n9810_), .ZN(new_n9811_));
  NAND2_X1   g09527(.A1(new_n9811_), .A2(new_n9806_), .ZN(new_n9812_));
  AND2_X2    g09528(.A1(new_n9808_), .A2(new_n9812_), .Z(new_n9813_));
  NOR2_X1    g09529(.A1(new_n9802_), .A2(new_n9806_), .ZN(new_n9814_));
  NOR2_X1    g09530(.A1(new_n9811_), .A2(new_n9807_), .ZN(new_n9815_));
  OAI21_X1   g09531(.A1(new_n9814_), .A2(new_n9815_), .B(new_n9702_), .ZN(new_n9816_));
  OAI21_X1   g09532(.A1(new_n9813_), .A2(new_n9702_), .B(new_n9816_), .ZN(new_n9817_));
  INV_X1     g09533(.I(new_n9467_), .ZN(new_n9818_));
  NAND3_X1   g09534(.A1(new_n9466_), .A2(new_n9118_), .A3(new_n9818_), .ZN(new_n9819_));
  NOR2_X1    g09535(.A1(new_n9470_), .A2(new_n9469_), .ZN(new_n9820_));
  NOR2_X1    g09536(.A1(new_n9819_), .A2(new_n9820_), .ZN(new_n9821_));
  NAND3_X1   g09537(.A1(new_n9363_), .A2(new_n9102_), .A3(new_n9471_), .ZN(new_n9822_));
  AOI21_X1   g09538(.A1(new_n9819_), .A2(new_n9820_), .B(new_n9822_), .ZN(new_n9823_));
  NOR2_X1    g09539(.A1(new_n9823_), .A2(new_n9821_), .ZN(new_n9824_));
  NOR2_X1    g09540(.A1(new_n9824_), .A2(new_n9817_), .ZN(new_n9825_));
  AOI21_X1   g09541(.A1(new_n9808_), .A2(new_n9812_), .B(new_n9702_), .ZN(new_n9826_));
  OR2_X2     g09542(.A1(new_n9814_), .A2(new_n9815_), .Z(new_n9827_));
  AOI21_X1   g09543(.A1(new_n9827_), .A2(new_n9702_), .B(new_n9826_), .ZN(new_n9828_));
  NAND2_X1   g09544(.A1(new_n9454_), .A2(new_n9458_), .ZN(new_n9829_));
  NAND3_X1   g09545(.A1(new_n9468_), .A2(new_n9829_), .A3(new_n9466_), .ZN(new_n9830_));
  NOR3_X1    g09546(.A1(new_n9366_), .A2(new_n8734_), .A3(new_n9467_), .ZN(new_n9831_));
  INV_X1     g09547(.I(new_n9822_), .ZN(new_n9832_));
  OAI21_X1   g09548(.A1(new_n9831_), .A2(new_n9829_), .B(new_n9832_), .ZN(new_n9833_));
  NAND2_X1   g09549(.A1(new_n9833_), .A2(new_n9830_), .ZN(new_n9834_));
  NOR2_X1    g09550(.A1(new_n9834_), .A2(new_n9828_), .ZN(new_n9835_));
  OAI22_X1   g09551(.A1(new_n4072_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n4067_), .ZN(new_n9836_));
  OAI21_X1   g09552(.A1(new_n1189_), .A2(new_n4318_), .B(new_n9836_), .ZN(new_n9837_));
  AOI21_X1   g09553(.A1(new_n9837_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n9838_));
  XNOR2_X1   g09554(.A1(new_n1421_), .A2(new_n9838_), .ZN(new_n9839_));
  NOR3_X1    g09555(.A1(new_n9835_), .A2(new_n9825_), .A3(new_n9839_), .ZN(new_n9840_));
  NAND2_X1   g09556(.A1(new_n9834_), .A2(new_n9828_), .ZN(new_n9841_));
  NAND2_X1   g09557(.A1(new_n9824_), .A2(new_n9817_), .ZN(new_n9842_));
  INV_X1     g09558(.I(new_n9839_), .ZN(new_n9843_));
  AOI21_X1   g09559(.A1(new_n9841_), .A2(new_n9842_), .B(new_n9843_), .ZN(new_n9844_));
  OAI21_X1   g09560(.A1(new_n9840_), .A2(new_n9844_), .B(new_n9698_), .ZN(new_n9845_));
  AOI21_X1   g09561(.A1(new_n9487_), .A2(new_n9488_), .B(new_n9136_), .ZN(new_n9846_));
  NOR3_X1    g09562(.A1(new_n9477_), .A2(new_n9474_), .A3(new_n9140_), .ZN(new_n9847_));
  NOR2_X1    g09563(.A1(new_n9847_), .A2(new_n9481_), .ZN(new_n9848_));
  AOI21_X1   g09564(.A1(new_n9848_), .A2(new_n9361_), .B(new_n9846_), .ZN(new_n9849_));
  OAI21_X1   g09565(.A1(new_n9835_), .A2(new_n9825_), .B(new_n9843_), .ZN(new_n9850_));
  NAND3_X1   g09566(.A1(new_n9841_), .A2(new_n9842_), .A3(new_n9839_), .ZN(new_n9851_));
  NAND2_X1   g09567(.A1(new_n9850_), .A2(new_n9851_), .ZN(new_n9852_));
  NAND2_X1   g09568(.A1(new_n9852_), .A2(new_n9849_), .ZN(new_n9853_));
  NAND2_X1   g09569(.A1(new_n9845_), .A2(new_n9853_), .ZN(new_n9854_));
  OAI22_X1   g09570(.A1(new_n1634_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1803_), .ZN(new_n9855_));
  OAI21_X1   g09571(.A1(new_n1525_), .A2(new_n3569_), .B(new_n9855_), .ZN(new_n9856_));
  AOI21_X1   g09572(.A1(new_n9856_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n9857_));
  XOR2_X1    g09573(.A1(new_n1808_), .A2(new_n9857_), .Z(new_n9858_));
  INV_X1     g09574(.I(new_n9858_), .ZN(new_n9859_));
  NAND2_X1   g09575(.A1(new_n9854_), .A2(new_n9859_), .ZN(new_n9860_));
  NAND3_X1   g09576(.A1(new_n9841_), .A2(new_n9842_), .A3(new_n9843_), .ZN(new_n9861_));
  OAI21_X1   g09577(.A1(new_n9835_), .A2(new_n9825_), .B(new_n9839_), .ZN(new_n9862_));
  AOI21_X1   g09578(.A1(new_n9861_), .A2(new_n9862_), .B(new_n9849_), .ZN(new_n9863_));
  AOI21_X1   g09579(.A1(new_n9850_), .A2(new_n9851_), .B(new_n9698_), .ZN(new_n9864_));
  NOR2_X1    g09580(.A1(new_n9863_), .A2(new_n9864_), .ZN(new_n9865_));
  NAND2_X1   g09581(.A1(new_n9865_), .A2(new_n9858_), .ZN(new_n9866_));
  NAND2_X1   g09582(.A1(new_n9866_), .A2(new_n9860_), .ZN(new_n9867_));
  AOI21_X1   g09583(.A1(new_n9493_), .A2(new_n9492_), .B(new_n9140_), .ZN(new_n9868_));
  NOR3_X1    g09584(.A1(new_n9484_), .A2(new_n9490_), .A3(new_n9136_), .ZN(new_n9869_));
  OAI21_X1   g09585(.A1(new_n9868_), .A2(new_n9869_), .B(new_n9151_), .ZN(new_n9870_));
  OAI21_X1   g09586(.A1(new_n9151_), .A2(new_n9147_), .B(new_n8765_), .ZN(new_n9871_));
  NAND2_X1   g09587(.A1(new_n9871_), .A2(new_n9011_), .ZN(new_n9872_));
  INV_X1     g09588(.I(new_n9498_), .ZN(new_n9873_));
  NAND3_X1   g09589(.A1(new_n9491_), .A2(new_n9494_), .A3(new_n9156_), .ZN(new_n9874_));
  NAND4_X1   g09590(.A1(new_n9872_), .A2(new_n9874_), .A3(new_n8773_), .A4(new_n9873_), .ZN(new_n9875_));
  OAI22_X1   g09591(.A1(new_n2102_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n2281_), .ZN(new_n9876_));
  OAI21_X1   g09592(.A1(new_n1936_), .A2(new_n2884_), .B(new_n9876_), .ZN(new_n9877_));
  AOI21_X1   g09593(.A1(new_n9877_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n9878_));
  XNOR2_X1   g09594(.A1(new_n2280_), .A2(new_n9878_), .ZN(new_n9879_));
  AOI21_X1   g09595(.A1(new_n9875_), .A2(new_n9870_), .B(new_n9879_), .ZN(new_n9880_));
  NAND3_X1   g09596(.A1(new_n9875_), .A2(new_n9870_), .A3(new_n9879_), .ZN(new_n9881_));
  INV_X1     g09597(.I(new_n9881_), .ZN(new_n9882_));
  OAI21_X1   g09598(.A1(new_n9882_), .A2(new_n9880_), .B(new_n9867_), .ZN(new_n9883_));
  NOR2_X1    g09599(.A1(new_n9865_), .A2(new_n9858_), .ZN(new_n9884_));
  NOR2_X1    g09600(.A1(new_n9854_), .A2(new_n9859_), .ZN(new_n9885_));
  NOR2_X1    g09601(.A1(new_n9884_), .A2(new_n9885_), .ZN(new_n9886_));
  NAND2_X1   g09602(.A1(new_n9874_), .A2(new_n9873_), .ZN(new_n9887_));
  OAI21_X1   g09603(.A1(new_n9887_), .A2(new_n9359_), .B(new_n9870_), .ZN(new_n9888_));
  NOR2_X1    g09604(.A1(new_n9888_), .A2(new_n9879_), .ZN(new_n9889_));
  INV_X1     g09605(.I(new_n9879_), .ZN(new_n9890_));
  AOI21_X1   g09606(.A1(new_n9875_), .A2(new_n9870_), .B(new_n9890_), .ZN(new_n9891_));
  OAI21_X1   g09607(.A1(new_n9889_), .A2(new_n9891_), .B(new_n9886_), .ZN(new_n9892_));
  NAND2_X1   g09608(.A1(new_n9883_), .A2(new_n9892_), .ZN(new_n9893_));
  OAI21_X1   g09609(.A1(new_n9694_), .A2(new_n9692_), .B(new_n9893_), .ZN(new_n9894_));
  INV_X1     g09610(.I(new_n9692_), .ZN(new_n9895_));
  NAND3_X1   g09611(.A1(new_n9517_), .A2(new_n9518_), .A3(new_n9350_), .ZN(new_n9896_));
  NAND3_X1   g09612(.A1(new_n9896_), .A2(new_n9357_), .A3(new_n9510_), .ZN(new_n9897_));
  INV_X1     g09613(.I(new_n9880_), .ZN(new_n9898_));
  AOI21_X1   g09614(.A1(new_n9898_), .A2(new_n9881_), .B(new_n9886_), .ZN(new_n9899_));
  NAND3_X1   g09615(.A1(new_n9875_), .A2(new_n9870_), .A3(new_n9890_), .ZN(new_n9900_));
  NAND2_X1   g09616(.A1(new_n9888_), .A2(new_n9879_), .ZN(new_n9901_));
  AOI21_X1   g09617(.A1(new_n9901_), .A2(new_n9900_), .B(new_n9867_), .ZN(new_n9902_));
  NOR2_X1    g09618(.A1(new_n9899_), .A2(new_n9902_), .ZN(new_n9903_));
  NAND3_X1   g09619(.A1(new_n9897_), .A2(new_n9903_), .A3(new_n9895_), .ZN(new_n9904_));
  OAI22_X1   g09620(.A1(new_n2171_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n2166_), .ZN(new_n9905_));
  OAI21_X1   g09621(.A1(new_n2439_), .A2(new_n2322_), .B(new_n9905_), .ZN(new_n9906_));
  AOI21_X1   g09622(.A1(new_n9906_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n9907_));
  XNOR2_X1   g09623(.A1(new_n2846_), .A2(new_n9907_), .ZN(new_n9908_));
  INV_X1     g09624(.I(new_n9908_), .ZN(new_n9909_));
  NAND3_X1   g09625(.A1(new_n9894_), .A2(new_n9904_), .A3(new_n9909_), .ZN(new_n9910_));
  AOI21_X1   g09626(.A1(new_n9897_), .A2(new_n9895_), .B(new_n9903_), .ZN(new_n9911_));
  NOR3_X1    g09627(.A1(new_n9694_), .A2(new_n9692_), .A3(new_n9893_), .ZN(new_n9912_));
  OAI21_X1   g09628(.A1(new_n9911_), .A2(new_n9912_), .B(new_n9908_), .ZN(new_n9913_));
  NAND2_X1   g09629(.A1(new_n9913_), .A2(new_n9910_), .ZN(new_n9914_));
  OAI22_X1   g09630(.A1(new_n1712_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n1707_), .ZN(new_n9915_));
  OAI21_X1   g09631(.A1(new_n3018_), .A2(new_n1850_), .B(new_n9915_), .ZN(new_n9916_));
  AOI21_X1   g09632(.A1(new_n9916_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n9917_));
  XNOR2_X1   g09633(.A1(new_n3514_), .A2(new_n9917_), .ZN(new_n9918_));
  INV_X1     g09634(.I(new_n9918_), .ZN(new_n9919_));
  XOR2_X1    g09635(.A1(new_n9914_), .A2(new_n9919_), .Z(new_n9920_));
  XOR2_X1    g09636(.A1(new_n9914_), .A2(new_n9919_), .Z(new_n9921_));
  NOR2_X1    g09637(.A1(new_n9921_), .A2(new_n9691_), .ZN(new_n9922_));
  AOI21_X1   g09638(.A1(new_n9691_), .A2(new_n9920_), .B(new_n9922_), .ZN(new_n9923_));
  OAI22_X1   g09639(.A1(new_n1347_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n1344_), .ZN(new_n9924_));
  OAI21_X1   g09640(.A1(new_n3717_), .A2(new_n1457_), .B(new_n9924_), .ZN(new_n9925_));
  AOI21_X1   g09641(.A1(new_n9925_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n9926_));
  XNOR2_X1   g09642(.A1(new_n4257_), .A2(new_n9926_), .ZN(new_n9927_));
  NOR2_X1    g09643(.A1(new_n9923_), .A2(new_n9927_), .ZN(new_n9928_));
  NAND2_X1   g09644(.A1(new_n9920_), .A2(new_n9691_), .ZN(new_n9929_));
  OAI21_X1   g09645(.A1(new_n9691_), .A2(new_n9921_), .B(new_n9929_), .ZN(new_n9930_));
  INV_X1     g09646(.I(new_n9927_), .ZN(new_n9931_));
  NOR2_X1    g09647(.A1(new_n9930_), .A2(new_n9931_), .ZN(new_n9932_));
  OAI21_X1   g09648(.A1(new_n9928_), .A2(new_n9932_), .B(new_n9686_), .ZN(new_n9933_));
  NOR3_X1    g09649(.A1(new_n9535_), .A2(new_n9539_), .A3(new_n9337_), .ZN(new_n9934_));
  NOR2_X1    g09650(.A1(new_n9934_), .A2(new_n9543_), .ZN(new_n9935_));
  AOI21_X1   g09651(.A1(new_n9935_), .A2(new_n9340_), .B(new_n9682_), .ZN(new_n9936_));
  NOR2_X1    g09652(.A1(new_n9930_), .A2(new_n9927_), .ZN(new_n9937_));
  NOR2_X1    g09653(.A1(new_n9923_), .A2(new_n9931_), .ZN(new_n9938_));
  OAI21_X1   g09654(.A1(new_n9938_), .A2(new_n9937_), .B(new_n9936_), .ZN(new_n9939_));
  NAND2_X1   g09655(.A1(new_n9939_), .A2(new_n9933_), .ZN(new_n9940_));
  OAI22_X1   g09656(.A1(new_n1055_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n1061_), .ZN(new_n9941_));
  OAI21_X1   g09657(.A1(new_n4500_), .A2(new_n1332_), .B(new_n9941_), .ZN(new_n9942_));
  AOI21_X1   g09658(.A1(new_n9942_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n9943_));
  XOR2_X1    g09659(.A1(new_n5067_), .A2(new_n9943_), .Z(new_n9944_));
  INV_X1     g09660(.I(new_n9944_), .ZN(new_n9945_));
  NAND2_X1   g09661(.A1(new_n9940_), .A2(new_n9945_), .ZN(new_n9946_));
  NAND3_X1   g09662(.A1(new_n9939_), .A2(new_n9933_), .A3(new_n9944_), .ZN(new_n9947_));
  NAND2_X1   g09663(.A1(new_n9946_), .A2(new_n9947_), .ZN(new_n9948_));
  NAND2_X1   g09664(.A1(new_n9948_), .A2(new_n9681_), .ZN(new_n9949_));
  XOR2_X1    g09665(.A1(new_n9940_), .A2(new_n9944_), .Z(new_n9950_));
  OAI21_X1   g09666(.A1(new_n9681_), .A2(new_n9950_), .B(new_n9949_), .ZN(new_n9951_));
  OAI22_X1   g09667(.A1(new_n970_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n820_), .ZN(new_n9952_));
  OAI21_X1   g09668(.A1(new_n5353_), .A2(new_n894_), .B(new_n9952_), .ZN(new_n9953_));
  AOI21_X1   g09669(.A1(new_n9953_), .A2(new_n827_), .B(new_n970_), .ZN(new_n9954_));
  XOR2_X1    g09670(.A1(new_n5926_), .A2(new_n9954_), .Z(new_n9955_));
  XOR2_X1    g09671(.A1(new_n9951_), .A2(new_n9955_), .Z(new_n9956_));
  NAND2_X1   g09672(.A1(new_n9956_), .A2(new_n9677_), .ZN(new_n9957_));
  AOI21_X1   g09673(.A1(new_n9584_), .A2(new_n9585_), .B(new_n9231_), .ZN(new_n9958_));
  AOI21_X1   g09674(.A1(new_n9674_), .A2(new_n9231_), .B(new_n9578_), .ZN(new_n9959_));
  AOI21_X1   g09675(.A1(new_n9959_), .A2(new_n9333_), .B(new_n9958_), .ZN(new_n9960_));
  INV_X1     g09676(.I(new_n9955_), .ZN(new_n9961_));
  XOR2_X1    g09677(.A1(new_n9951_), .A2(new_n9961_), .Z(new_n9962_));
  NAND2_X1   g09678(.A1(new_n9962_), .A2(new_n9960_), .ZN(new_n9963_));
  NAND2_X1   g09679(.A1(new_n9957_), .A2(new_n9963_), .ZN(new_n9964_));
  NAND2_X1   g09680(.A1(new_n9964_), .A2(new_n9673_), .ZN(new_n9965_));
  OAI21_X1   g09681(.A1(new_n9600_), .A2(new_n9601_), .B(new_n9242_), .ZN(new_n9966_));
  NAND3_X1   g09682(.A1(new_n9588_), .A2(new_n9591_), .A3(new_n9247_), .ZN(new_n9967_));
  NAND2_X1   g09683(.A1(new_n9967_), .A2(new_n9602_), .ZN(new_n9968_));
  OAI21_X1   g09684(.A1(new_n9968_), .A2(new_n9331_), .B(new_n9966_), .ZN(new_n9969_));
  XOR2_X1    g09685(.A1(new_n9951_), .A2(new_n9961_), .Z(new_n9970_));
  XOR2_X1    g09686(.A1(new_n9951_), .A2(new_n9955_), .Z(new_n9971_));
  MUX2_X1    g09687(.I0(new_n9971_), .I1(new_n9970_), .S(new_n9677_), .Z(new_n9972_));
  NAND2_X1   g09688(.A1(new_n9972_), .A2(new_n9969_), .ZN(new_n9973_));
  NAND2_X1   g09689(.A1(new_n9965_), .A2(new_n9973_), .ZN(new_n9974_));
  OAI22_X1   g09690(.A1(new_n607_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n610_), .ZN(new_n9975_));
  OAI21_X1   g09691(.A1(new_n6229_), .A2(new_n684_), .B(new_n9975_), .ZN(new_n9976_));
  AOI21_X1   g09692(.A1(new_n9976_), .A2(new_n612_), .B(new_n607_), .ZN(new_n9977_));
  XOR2_X1    g09693(.A1(new_n6851_), .A2(new_n9977_), .Z(new_n9978_));
  NOR2_X1    g09694(.A1(new_n9974_), .A2(new_n9978_), .ZN(new_n9979_));
  INV_X1     g09695(.I(new_n9978_), .ZN(new_n9980_));
  AOI21_X1   g09696(.A1(new_n9965_), .A2(new_n9973_), .B(new_n9980_), .ZN(new_n9981_));
  OAI21_X1   g09697(.A1(new_n9979_), .A2(new_n9981_), .B(new_n9669_), .ZN(new_n9982_));
  NAND2_X1   g09698(.A1(new_n9667_), .A2(new_n9613_), .ZN(new_n9983_));
  NOR2_X1    g09699(.A1(new_n9983_), .A2(new_n9617_), .ZN(new_n9984_));
  NOR2_X1    g09700(.A1(new_n9984_), .A2(new_n9665_), .ZN(new_n9985_));
  XOR2_X1    g09701(.A1(new_n9974_), .A2(new_n9978_), .Z(new_n9986_));
  NAND2_X1   g09702(.A1(new_n9985_), .A2(new_n9986_), .ZN(new_n9987_));
  OAI22_X1   g09703(.A1(new_n448_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n450_), .ZN(new_n9988_));
  OAI21_X1   g09704(.A1(new_n7198_), .A2(new_n496_), .B(new_n9988_), .ZN(new_n9989_));
  AOI21_X1   g09705(.A1(new_n9989_), .A2(new_n452_), .B(new_n448_), .ZN(new_n9990_));
  XNOR2_X1   g09706(.A1(new_n7874_), .A2(new_n9990_), .ZN(new_n9991_));
  AOI21_X1   g09707(.A1(new_n9982_), .A2(new_n9987_), .B(new_n9991_), .ZN(new_n9992_));
  NAND3_X1   g09708(.A1(new_n9982_), .A2(new_n9987_), .A3(new_n9991_), .ZN(new_n9993_));
  INV_X1     g09709(.I(new_n9993_), .ZN(new_n9994_));
  NOR2_X1    g09710(.A1(new_n9994_), .A2(new_n9992_), .ZN(new_n9995_));
  NAND2_X1   g09711(.A1(new_n9624_), .A2(new_n9273_), .ZN(new_n9996_));
  INV_X1     g09712(.I(new_n9996_), .ZN(new_n9997_));
  AOI21_X1   g09713(.A1(new_n9621_), .A2(new_n9622_), .B(new_n9258_), .ZN(new_n9998_));
  NOR3_X1    g09714(.A1(new_n9619_), .A2(new_n9615_), .A3(new_n9262_), .ZN(new_n9999_));
  NOR3_X1    g09715(.A1(new_n9999_), .A2(new_n9998_), .A3(new_n9273_), .ZN(new_n10000_));
  NOR3_X1    g09716(.A1(new_n9324_), .A2(new_n9628_), .A3(new_n10000_), .ZN(new_n10001_));
  OAI22_X1   g09717(.A1(new_n8563_), .A2(new_n341_), .B1(new_n404_), .B2(new_n8948_), .ZN(new_n10002_));
  OAI21_X1   g09718(.A1(new_n8218_), .A2(new_n366_), .B(new_n10002_), .ZN(new_n10003_));
  AOI21_X1   g09719(.A1(new_n10003_), .A2(new_n334_), .B(new_n341_), .ZN(new_n10004_));
  XOR2_X1    g09720(.A1(new_n8952_), .A2(new_n10004_), .Z(new_n10005_));
  INV_X1     g09721(.I(new_n10005_), .ZN(new_n10006_));
  OAI21_X1   g09722(.A1(new_n10001_), .A2(new_n9997_), .B(new_n10006_), .ZN(new_n10007_));
  AOI21_X1   g09723(.A1(new_n8921_), .A2(new_n8916_), .B(new_n8926_), .ZN(new_n10008_));
  AOI21_X1   g09724(.A1(new_n9271_), .A2(new_n9270_), .B(new_n9268_), .ZN(new_n10009_));
  NOR3_X1    g09725(.A1(new_n9260_), .A2(new_n9264_), .A3(new_n9272_), .ZN(new_n10010_));
  OAI21_X1   g09726(.A1(new_n10010_), .A2(new_n10009_), .B(new_n10008_), .ZN(new_n10011_));
  NAND3_X1   g09727(.A1(new_n10011_), .A2(new_n8933_), .A3(new_n8980_), .ZN(new_n10012_));
  NAND3_X1   g09728(.A1(new_n9620_), .A2(new_n9623_), .A3(new_n9322_), .ZN(new_n10013_));
  NAND4_X1   g09729(.A1(new_n10012_), .A2(new_n8931_), .A3(new_n10013_), .A4(new_n9629_), .ZN(new_n10014_));
  NAND3_X1   g09730(.A1(new_n10014_), .A2(new_n9996_), .A3(new_n10005_), .ZN(new_n10015_));
  AOI21_X1   g09731(.A1(new_n10007_), .A2(new_n10015_), .B(new_n9995_), .ZN(new_n10016_));
  INV_X1     g09732(.I(new_n9992_), .ZN(new_n10017_));
  NAND2_X1   g09733(.A1(new_n10017_), .A2(new_n9993_), .ZN(new_n10018_));
  NAND3_X1   g09734(.A1(new_n10014_), .A2(new_n9996_), .A3(new_n10006_), .ZN(new_n10019_));
  OAI21_X1   g09735(.A1(new_n10001_), .A2(new_n9997_), .B(new_n10005_), .ZN(new_n10020_));
  AOI21_X1   g09736(.A1(new_n10020_), .A2(new_n10019_), .B(new_n10018_), .ZN(new_n10021_));
  NOR2_X1    g09737(.A1(new_n10016_), .A2(new_n10021_), .ZN(new_n10022_));
  NOR2_X1    g09738(.A1(\b[50] ), .A2(\b[51] ), .ZN(new_n10023_));
  AOI21_X1   g09739(.A1(new_n9293_), .A2(new_n10023_), .B(new_n8948_), .ZN(new_n10024_));
  INV_X1     g09740(.I(\b[51] ), .ZN(new_n10025_));
  NOR2_X1    g09741(.A1(new_n9295_), .A2(new_n10025_), .ZN(new_n10026_));
  INV_X1     g09742(.I(new_n10026_), .ZN(new_n10027_));
  NOR2_X1    g09743(.A1(new_n9293_), .A2(new_n10027_), .ZN(new_n10028_));
  NOR2_X1    g09744(.A1(new_n10024_), .A2(new_n10028_), .ZN(new_n10029_));
  XNOR2_X1   g09745(.A1(\b[51] ), .A2(\b[52] ), .ZN(new_n10030_));
  INV_X1     g09746(.I(\b[52] ), .ZN(new_n10031_));
  NOR2_X1    g09747(.A1(new_n10025_), .A2(new_n10031_), .ZN(new_n10032_));
  NOR2_X1    g09748(.A1(\b[51] ), .A2(\b[52] ), .ZN(new_n10033_));
  OAI21_X1   g09749(.A1(new_n10032_), .A2(new_n10033_), .B(new_n10029_), .ZN(new_n10034_));
  OAI21_X1   g09750(.A1(new_n10029_), .A2(new_n10030_), .B(new_n10034_), .ZN(new_n10035_));
  OAI22_X1   g09751(.A1(new_n330_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n263_), .ZN(new_n10036_));
  OAI21_X1   g09752(.A1(new_n9295_), .A2(new_n289_), .B(new_n10036_), .ZN(new_n10037_));
  AOI21_X1   g09753(.A1(new_n10037_), .A2(new_n260_), .B(new_n426_), .ZN(new_n10038_));
  XNOR2_X1   g09754(.A1(new_n10035_), .A2(new_n10038_), .ZN(new_n10039_));
  XOR2_X1    g09755(.A1(new_n10022_), .A2(new_n10039_), .Z(new_n10040_));
  OAI21_X1   g09756(.A1(new_n9662_), .A2(new_n9660_), .B(new_n10040_), .ZN(new_n10041_));
  NOR2_X1    g09757(.A1(new_n9662_), .A2(new_n9660_), .ZN(new_n10042_));
  INV_X1     g09758(.I(new_n10039_), .ZN(new_n10043_));
  XOR2_X1    g09759(.A1(new_n10022_), .A2(new_n10043_), .Z(new_n10044_));
  NAND2_X1   g09760(.A1(new_n10042_), .A2(new_n10044_), .ZN(new_n10045_));
  NAND2_X1   g09761(.A1(new_n10045_), .A2(new_n10041_), .ZN(new_n10046_));
  NOR3_X1    g09762(.A1(new_n9653_), .A2(new_n9656_), .A3(new_n9287_), .ZN(new_n10047_));
  OAI21_X1   g09763(.A1(new_n9653_), .A2(new_n9656_), .B(new_n9287_), .ZN(new_n10048_));
  AOI21_X1   g09764(.A1(new_n10048_), .A2(new_n9303_), .B(new_n10047_), .ZN(new_n10049_));
  NAND3_X1   g09765(.A1(new_n8968_), .A2(new_n10049_), .A3(new_n8978_), .ZN(new_n10050_));
  INV_X1     g09766(.I(new_n10050_), .ZN(new_n10051_));
  XOR2_X1    g09767(.A1(new_n9639_), .A2(new_n9320_), .Z(new_n10052_));
  NOR2_X1    g09768(.A1(new_n10052_), .A2(new_n9648_), .ZN(new_n10053_));
  NOR2_X1    g09769(.A1(new_n10051_), .A2(new_n10053_), .ZN(new_n10054_));
  OAI21_X1   g09770(.A1(new_n9648_), .A2(new_n10052_), .B(new_n10046_), .ZN(new_n10055_));
  OAI22_X1   g09771(.A1(new_n10054_), .A2(new_n10046_), .B1(new_n10051_), .B2(new_n10055_), .ZN(\f[52] ));
  XOR2_X1    g09772(.A1(new_n10042_), .A2(new_n10022_), .Z(new_n10057_));
  AOI21_X1   g09773(.A1(new_n10045_), .A2(new_n10041_), .B(new_n10043_), .ZN(new_n10058_));
  AOI21_X1   g09774(.A1(new_n10057_), .A2(new_n10058_), .B(new_n10053_), .ZN(new_n10059_));
  NOR2_X1    g09775(.A1(new_n10050_), .A2(new_n10059_), .ZN(new_n10060_));
  INV_X1     g09776(.I(new_n10060_), .ZN(new_n10061_));
  NAND2_X1   g09777(.A1(new_n10014_), .A2(new_n9996_), .ZN(new_n10062_));
  NAND2_X1   g09778(.A1(new_n9995_), .A2(new_n10062_), .ZN(new_n10063_));
  NOR2_X1    g09779(.A1(new_n10001_), .A2(new_n9997_), .ZN(new_n10064_));
  NAND2_X1   g09780(.A1(new_n10064_), .A2(new_n10018_), .ZN(new_n10065_));
  AOI21_X1   g09781(.A1(new_n10065_), .A2(new_n10063_), .B(new_n10006_), .ZN(new_n10066_));
  OAI21_X1   g09782(.A1(new_n10016_), .A2(new_n10021_), .B(new_n9635_), .ZN(new_n10067_));
  XNOR2_X1   g09783(.A1(new_n9630_), .A2(new_n9325_), .ZN(new_n10068_));
  NAND2_X1   g09784(.A1(new_n10067_), .A2(new_n10068_), .ZN(new_n10069_));
  OAI21_X1   g09785(.A1(new_n9001_), .A2(new_n9279_), .B(new_n9318_), .ZN(new_n10070_));
  NOR3_X1    g09786(.A1(new_n10016_), .A2(new_n10021_), .A3(new_n9635_), .ZN(new_n10071_));
  AOI21_X1   g09787(.A1(new_n10070_), .A2(new_n9314_), .B(new_n10071_), .ZN(new_n10072_));
  NAND2_X1   g09788(.A1(new_n10072_), .A2(new_n10069_), .ZN(new_n10073_));
  OAI22_X1   g09789(.A1(new_n607_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n610_), .ZN(new_n10074_));
  OAI21_X1   g09790(.A1(new_n6538_), .A2(new_n684_), .B(new_n10074_), .ZN(new_n10075_));
  AOI21_X1   g09791(.A1(new_n10075_), .A2(new_n612_), .B(new_n607_), .ZN(new_n10076_));
  XNOR2_X1   g09792(.A1(new_n7202_), .A2(new_n10076_), .ZN(new_n10077_));
  INV_X1     g09793(.I(new_n10077_), .ZN(new_n10078_));
  NAND2_X1   g09794(.A1(new_n9960_), .A2(new_n9951_), .ZN(new_n10079_));
  INV_X1     g09795(.I(new_n9951_), .ZN(new_n10080_));
  NAND2_X1   g09796(.A1(new_n10080_), .A2(new_n9677_), .ZN(new_n10081_));
  AOI21_X1   g09797(.A1(new_n10081_), .A2(new_n10079_), .B(new_n9961_), .ZN(new_n10082_));
  NOR2_X1    g09798(.A1(new_n9678_), .A2(new_n9571_), .ZN(new_n10083_));
  AOI21_X1   g09799(.A1(new_n9678_), .A2(new_n9571_), .B(new_n9560_), .ZN(new_n10084_));
  AOI21_X1   g09800(.A1(new_n10084_), .A2(new_n9564_), .B(new_n10083_), .ZN(new_n10085_));
  NAND2_X1   g09801(.A1(new_n10085_), .A2(new_n9940_), .ZN(new_n10086_));
  AND2_X2    g09802(.A1(new_n9939_), .A2(new_n9933_), .Z(new_n10087_));
  NAND2_X1   g09803(.A1(new_n9681_), .A2(new_n10087_), .ZN(new_n10088_));
  AOI21_X1   g09804(.A1(new_n10088_), .A2(new_n10086_), .B(new_n9945_), .ZN(new_n10089_));
  NAND2_X1   g09805(.A1(new_n9936_), .A2(new_n9930_), .ZN(new_n10090_));
  NAND2_X1   g09806(.A1(new_n9686_), .A2(new_n9923_), .ZN(new_n10091_));
  AOI21_X1   g09807(.A1(new_n10090_), .A2(new_n10091_), .B(new_n9931_), .ZN(new_n10092_));
  NAND2_X1   g09808(.A1(new_n9691_), .A2(new_n9914_), .ZN(new_n10093_));
  NOR2_X1    g09809(.A1(new_n9691_), .A2(new_n9914_), .ZN(new_n10094_));
  INV_X1     g09810(.I(new_n10094_), .ZN(new_n10095_));
  AOI21_X1   g09811(.A1(new_n10095_), .A2(new_n10093_), .B(new_n9919_), .ZN(new_n10096_));
  INV_X1     g09812(.I(new_n9690_), .ZN(new_n10097_));
  AOI22_X1   g09813(.A1(new_n10097_), .A2(new_n9532_), .B1(new_n9346_), .B2(new_n9687_), .ZN(new_n10098_));
  NOR2_X1    g09814(.A1(new_n9911_), .A2(new_n9912_), .ZN(new_n10099_));
  NOR2_X1    g09815(.A1(new_n10099_), .A2(new_n9908_), .ZN(new_n10100_));
  NOR2_X1    g09816(.A1(new_n9694_), .A2(new_n9692_), .ZN(new_n10101_));
  INV_X1     g09817(.I(new_n9870_), .ZN(new_n10102_));
  NOR3_X1    g09818(.A1(new_n9868_), .A2(new_n9869_), .A3(new_n9151_), .ZN(new_n10103_));
  NOR3_X1    g09819(.A1(new_n9359_), .A2(new_n10103_), .A3(new_n9498_), .ZN(new_n10104_));
  NOR2_X1    g09820(.A1(new_n10104_), .A2(new_n10102_), .ZN(new_n10105_));
  NOR2_X1    g09821(.A1(new_n10105_), .A2(new_n9867_), .ZN(new_n10106_));
  NOR2_X1    g09822(.A1(new_n9886_), .A2(new_n9888_), .ZN(new_n10107_));
  OAI21_X1   g09823(.A1(new_n10106_), .A2(new_n10107_), .B(new_n9879_), .ZN(new_n10108_));
  NOR3_X1    g09824(.A1(new_n9486_), .A2(new_n9481_), .A3(new_n9847_), .ZN(new_n10109_));
  OAI21_X1   g09825(.A1(new_n10109_), .A2(new_n9846_), .B(new_n9862_), .ZN(new_n10110_));
  XOR2_X1    g09826(.A1(new_n9702_), .A2(new_n9802_), .Z(new_n10111_));
  NOR2_X1    g09827(.A1(new_n10111_), .A2(new_n9807_), .ZN(new_n10112_));
  INV_X1     g09828(.I(new_n10112_), .ZN(new_n10113_));
  NAND3_X1   g09829(.A1(new_n9833_), .A2(new_n9828_), .A3(new_n9830_), .ZN(new_n10114_));
  NOR2_X1    g09830(.A1(new_n9785_), .A2(new_n9792_), .ZN(new_n10115_));
  NOR2_X1    g09831(.A1(new_n10115_), .A2(new_n9796_), .ZN(new_n10116_));
  OAI21_X1   g09832(.A1(new_n9788_), .A2(new_n9786_), .B(new_n9784_), .ZN(new_n10117_));
  OAI21_X1   g09833(.A1(new_n9709_), .A2(new_n9707_), .B(new_n9770_), .ZN(new_n10118_));
  NAND2_X1   g09834(.A1(new_n9742_), .A2(new_n9740_), .ZN(new_n10119_));
  NAND2_X1   g09835(.A1(new_n10119_), .A2(new_n9746_), .ZN(new_n10120_));
  XOR2_X1    g09836(.A1(new_n9734_), .A2(\a[50] ), .Z(new_n10121_));
  OAI21_X1   g09837(.A1(new_n10119_), .A2(new_n9746_), .B(new_n10121_), .ZN(new_n10122_));
  NOR2_X1    g09838(.A1(new_n9394_), .A2(\a[52] ), .ZN(new_n10123_));
  AOI21_X1   g09839(.A1(\a[52] ), .A2(new_n9395_), .B(new_n10123_), .ZN(new_n10124_));
  XNOR2_X1   g09840(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n10125_));
  NAND3_X1   g09841(.A1(new_n10125_), .A2(new_n9394_), .A3(new_n9396_), .ZN(new_n10126_));
  INV_X1     g09842(.I(new_n9719_), .ZN(new_n10127_));
  OAI21_X1   g09843(.A1(new_n10126_), .A2(new_n10124_), .B(new_n10127_), .ZN(new_n10128_));
  AOI21_X1   g09844(.A1(new_n10128_), .A2(new_n9712_), .B(new_n444_), .ZN(new_n10129_));
  NOR3_X1    g09845(.A1(new_n9721_), .A2(new_n10129_), .A3(new_n9745_), .ZN(new_n10130_));
  NAND2_X1   g09846(.A1(\b[1] ), .A2(\b[2] ), .ZN(new_n10131_));
  INV_X1     g09847(.I(new_n10131_), .ZN(new_n10132_));
  AOI21_X1   g09848(.A1(new_n9717_), .A2(new_n9715_), .B(new_n10132_), .ZN(new_n10133_));
  XOR2_X1    g09849(.A1(\a[50] ), .A2(\a[52] ), .Z(new_n10134_));
  XOR2_X1    g09850(.A1(\a[50] ), .A2(\a[53] ), .Z(new_n10135_));
  XOR2_X1    g09851(.A1(\a[50] ), .A2(\a[51] ), .Z(new_n10136_));
  NAND3_X1   g09852(.A1(new_n10134_), .A2(new_n10135_), .A3(new_n10136_), .ZN(new_n10137_));
  NOR2_X1    g09853(.A1(new_n10137_), .A2(new_n258_), .ZN(new_n10138_));
  OAI21_X1   g09854(.A1(new_n10133_), .A2(new_n10138_), .B(new_n9718_), .ZN(new_n10139_));
  NAND3_X1   g09855(.A1(new_n10139_), .A2(new_n282_), .A3(new_n9713_), .ZN(new_n10140_));
  OAI21_X1   g09856(.A1(new_n10126_), .A2(new_n10124_), .B(new_n10131_), .ZN(new_n10141_));
  XNOR2_X1   g09857(.A1(\a[50] ), .A2(\a[52] ), .ZN(new_n10142_));
  XNOR2_X1   g09858(.A1(\a[50] ), .A2(\a[53] ), .ZN(new_n10143_));
  XNOR2_X1   g09859(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n10144_));
  NOR3_X1    g09860(.A1(new_n10142_), .A2(new_n10143_), .A3(new_n10144_), .ZN(new_n10145_));
  NAND2_X1   g09861(.A1(new_n10145_), .A2(\b[0] ), .ZN(new_n10146_));
  AOI21_X1   g09862(.A1(new_n10146_), .A2(new_n10141_), .B(\a[53] ), .ZN(new_n10147_));
  OAI21_X1   g09863(.A1(new_n10147_), .A2(new_n490_), .B(new_n9712_), .ZN(new_n10148_));
  NAND2_X1   g09864(.A1(new_n10148_), .A2(new_n10140_), .ZN(new_n10149_));
  NAND2_X1   g09865(.A1(new_n10149_), .A2(new_n10130_), .ZN(new_n10150_));
  NAND3_X1   g09866(.A1(new_n9722_), .A2(new_n9723_), .A3(new_n9725_), .ZN(new_n10151_));
  NAND3_X1   g09867(.A1(new_n10151_), .A2(new_n10140_), .A3(new_n10148_), .ZN(new_n10152_));
  AOI22_X1   g09868(.A1(new_n8631_), .A2(\b[4] ), .B1(\b[5] ), .B2(new_n9382_), .ZN(new_n10153_));
  NAND3_X1   g09869(.A1(new_n9023_), .A2(new_n8636_), .A3(new_n9024_), .ZN(new_n10154_));
  NOR2_X1    g09870(.A1(new_n10154_), .A2(new_n298_), .ZN(new_n10155_));
  OAI21_X1   g09871(.A1(new_n10155_), .A2(new_n10153_), .B(new_n8624_), .ZN(new_n10156_));
  NAND3_X1   g09872(.A1(new_n10156_), .A2(new_n2333_), .A3(new_n8631_), .ZN(new_n10157_));
  AOI21_X1   g09873(.A1(new_n10156_), .A2(new_n8631_), .B(new_n2333_), .ZN(new_n10158_));
  INV_X1     g09874(.I(new_n10158_), .ZN(new_n10159_));
  NAND2_X1   g09875(.A1(new_n10159_), .A2(new_n10157_), .ZN(new_n10160_));
  NAND3_X1   g09876(.A1(new_n10150_), .A2(new_n10152_), .A3(new_n10160_), .ZN(new_n10161_));
  AOI21_X1   g09877(.A1(new_n10140_), .A2(new_n10148_), .B(new_n10151_), .ZN(new_n10162_));
  NOR2_X1    g09878(.A1(new_n10149_), .A2(new_n10130_), .ZN(new_n10163_));
  INV_X1     g09879(.I(new_n10157_), .ZN(new_n10164_));
  NOR2_X1    g09880(.A1(new_n10164_), .A2(new_n10158_), .ZN(new_n10165_));
  OAI21_X1   g09881(.A1(new_n10163_), .A2(new_n10162_), .B(new_n10165_), .ZN(new_n10166_));
  AOI22_X1   g09882(.A1(new_n10122_), .A2(new_n10120_), .B1(new_n10161_), .B2(new_n10166_), .ZN(new_n10167_));
  NOR2_X1    g09883(.A1(new_n9729_), .A2(new_n9727_), .ZN(new_n10168_));
  NOR2_X1    g09884(.A1(new_n10168_), .A2(new_n9726_), .ZN(new_n10169_));
  XOR2_X1    g09885(.A1(new_n9734_), .A2(new_n8624_), .Z(new_n10170_));
  AOI21_X1   g09886(.A1(new_n10168_), .A2(new_n9726_), .B(new_n10170_), .ZN(new_n10171_));
  AOI21_X1   g09887(.A1(new_n10150_), .A2(new_n10152_), .B(new_n10165_), .ZN(new_n10172_));
  NOR3_X1    g09888(.A1(new_n10163_), .A2(new_n10162_), .A3(new_n10160_), .ZN(new_n10173_));
  NOR2_X1    g09889(.A1(new_n10173_), .A2(new_n10172_), .ZN(new_n10174_));
  NOR3_X1    g09890(.A1(new_n10174_), .A2(new_n10171_), .A3(new_n10169_), .ZN(new_n10175_));
  OAI22_X1   g09891(.A1(new_n7619_), .A2(new_n472_), .B1(new_n515_), .B2(new_n8309_), .ZN(new_n10176_));
  OAI21_X1   g09892(.A1(new_n420_), .A2(new_n7947_), .B(new_n10176_), .ZN(new_n10177_));
  AOI21_X1   g09893(.A1(new_n10177_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n10178_));
  XOR2_X1    g09894(.A1(new_n700_), .A2(new_n10178_), .Z(new_n10179_));
  NOR3_X1    g09895(.A1(new_n10167_), .A2(new_n10175_), .A3(new_n10179_), .ZN(new_n10180_));
  NAND2_X1   g09896(.A1(new_n10166_), .A2(new_n10161_), .ZN(new_n10181_));
  OAI21_X1   g09897(.A1(new_n10169_), .A2(new_n10171_), .B(new_n10181_), .ZN(new_n10182_));
  OAI21_X1   g09898(.A1(new_n10163_), .A2(new_n10162_), .B(new_n10160_), .ZN(new_n10183_));
  NAND3_X1   g09899(.A1(new_n10150_), .A2(new_n10152_), .A3(new_n10165_), .ZN(new_n10184_));
  NAND2_X1   g09900(.A1(new_n10183_), .A2(new_n10184_), .ZN(new_n10185_));
  NAND3_X1   g09901(.A1(new_n10185_), .A2(new_n10122_), .A3(new_n10120_), .ZN(new_n10186_));
  XOR2_X1    g09902(.A1(new_n522_), .A2(new_n10178_), .Z(new_n10187_));
  AOI21_X1   g09903(.A1(new_n10182_), .A2(new_n10186_), .B(new_n10187_), .ZN(new_n10188_));
  NOR2_X1    g09904(.A1(new_n10188_), .A2(new_n10180_), .ZN(new_n10189_));
  AOI21_X1   g09905(.A1(new_n10118_), .A2(new_n9769_), .B(new_n10189_), .ZN(new_n10190_));
  AOI21_X1   g09906(.A1(new_n9766_), .A2(new_n9764_), .B(new_n9780_), .ZN(new_n10191_));
  AOI21_X1   g09907(.A1(new_n10182_), .A2(new_n10186_), .B(new_n10179_), .ZN(new_n10192_));
  NOR3_X1    g09908(.A1(new_n10167_), .A2(new_n10175_), .A3(new_n10187_), .ZN(new_n10193_));
  NOR2_X1    g09909(.A1(new_n10192_), .A2(new_n10193_), .ZN(new_n10194_));
  NOR3_X1    g09910(.A1(new_n10191_), .A2(new_n9768_), .A3(new_n10194_), .ZN(new_n10195_));
  OAI22_X1   g09911(.A1(new_n6644_), .A2(new_n656_), .B1(new_n706_), .B2(new_n6647_), .ZN(new_n10196_));
  OAI21_X1   g09912(.A1(new_n565_), .A2(new_n7284_), .B(new_n10196_), .ZN(new_n10197_));
  AOI21_X1   g09913(.A1(new_n10197_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n10198_));
  XNOR2_X1   g09914(.A1(new_n710_), .A2(new_n10198_), .ZN(new_n10199_));
  INV_X1     g09915(.I(new_n10199_), .ZN(new_n10200_));
  OAI21_X1   g09916(.A1(new_n10190_), .A2(new_n10195_), .B(new_n10200_), .ZN(new_n10201_));
  NAND3_X1   g09917(.A1(new_n10182_), .A2(new_n10186_), .A3(new_n10187_), .ZN(new_n10202_));
  OAI21_X1   g09918(.A1(new_n10167_), .A2(new_n10175_), .B(new_n10179_), .ZN(new_n10203_));
  NAND2_X1   g09919(.A1(new_n10203_), .A2(new_n10202_), .ZN(new_n10204_));
  OAI21_X1   g09920(.A1(new_n10191_), .A2(new_n9768_), .B(new_n10204_), .ZN(new_n10205_));
  OAI21_X1   g09921(.A1(new_n10167_), .A2(new_n10175_), .B(new_n10187_), .ZN(new_n10206_));
  NAND3_X1   g09922(.A1(new_n10182_), .A2(new_n10186_), .A3(new_n10179_), .ZN(new_n10207_));
  NAND2_X1   g09923(.A1(new_n10206_), .A2(new_n10207_), .ZN(new_n10208_));
  NAND3_X1   g09924(.A1(new_n10118_), .A2(new_n9769_), .A3(new_n10208_), .ZN(new_n10209_));
  NAND3_X1   g09925(.A1(new_n10209_), .A2(new_n10205_), .A3(new_n10199_), .ZN(new_n10210_));
  OAI22_X1   g09926(.A1(new_n5993_), .A2(new_n861_), .B1(new_n930_), .B2(new_n5991_), .ZN(new_n10211_));
  OAI21_X1   g09927(.A1(new_n780_), .A2(new_n5997_), .B(new_n10211_), .ZN(new_n10212_));
  AOI21_X1   g09928(.A1(new_n10212_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n10213_));
  NAND3_X1   g09929(.A1(new_n936_), .A2(new_n925_), .A3(new_n10213_), .ZN(new_n10214_));
  NOR2_X1    g09930(.A1(new_n1015_), .A2(new_n934_), .ZN(new_n10215_));
  INV_X1     g09931(.I(new_n10213_), .ZN(new_n10216_));
  OAI21_X1   g09932(.A1(new_n10215_), .A2(new_n924_), .B(new_n10216_), .ZN(new_n10217_));
  NAND2_X1   g09933(.A1(new_n10214_), .A2(new_n10217_), .ZN(new_n10218_));
  NAND3_X1   g09934(.A1(new_n10201_), .A2(new_n10210_), .A3(new_n10218_), .ZN(new_n10219_));
  AOI21_X1   g09935(.A1(new_n10209_), .A2(new_n10205_), .B(new_n10199_), .ZN(new_n10220_));
  NOR3_X1    g09936(.A1(new_n10190_), .A2(new_n10195_), .A3(new_n10200_), .ZN(new_n10221_));
  NOR3_X1    g09937(.A1(new_n10215_), .A2(new_n924_), .A3(new_n10216_), .ZN(new_n10222_));
  AOI21_X1   g09938(.A1(new_n936_), .A2(new_n925_), .B(new_n10213_), .ZN(new_n10223_));
  NOR2_X1    g09939(.A1(new_n10223_), .A2(new_n10222_), .ZN(new_n10224_));
  OAI21_X1   g09940(.A1(new_n10220_), .A2(new_n10221_), .B(new_n10224_), .ZN(new_n10225_));
  AOI22_X1   g09941(.A1(new_n10117_), .A2(new_n9777_), .B1(new_n10219_), .B2(new_n10225_), .ZN(new_n10226_));
  AOI21_X1   g09942(.A1(new_n9706_), .A2(new_n9704_), .B(new_n9783_), .ZN(new_n10227_));
  AOI21_X1   g09943(.A1(new_n10201_), .A2(new_n10210_), .B(new_n10224_), .ZN(new_n10228_));
  NOR3_X1    g09944(.A1(new_n10220_), .A2(new_n10221_), .A3(new_n10218_), .ZN(new_n10229_));
  NOR2_X1    g09945(.A1(new_n10229_), .A2(new_n10228_), .ZN(new_n10230_));
  NOR3_X1    g09946(.A1(new_n10230_), .A2(new_n9776_), .A3(new_n10227_), .ZN(new_n10231_));
  NOR2_X1    g09947(.A1(new_n10231_), .A2(new_n10226_), .ZN(new_n10232_));
  NOR3_X1    g09948(.A1(new_n9802_), .A2(new_n10232_), .A3(new_n10116_), .ZN(new_n10233_));
  NOR2_X1    g09949(.A1(new_n10227_), .A2(new_n9776_), .ZN(new_n10234_));
  NOR2_X1    g09950(.A1(new_n10220_), .A2(new_n10221_), .ZN(new_n10235_));
  NOR2_X1    g09951(.A1(new_n10115_), .A2(new_n9796_), .ZN(new_n10236_));
  OAI21_X1   g09952(.A1(new_n10233_), .A2(new_n10236_), .B(new_n9702_), .ZN(new_n10237_));
  INV_X1     g09953(.I(new_n9699_), .ZN(new_n10238_));
  NAND4_X1   g09954(.A1(new_n9700_), .A2(new_n9013_), .A3(new_n9362_), .A4(new_n9447_), .ZN(new_n10239_));
  NAND2_X1   g09955(.A1(new_n10239_), .A2(new_n10238_), .ZN(new_n10240_));
  INV_X1     g09956(.I(new_n10116_), .ZN(new_n10241_));
  NAND2_X1   g09957(.A1(new_n10225_), .A2(new_n10219_), .ZN(new_n10242_));
  OAI21_X1   g09958(.A1(new_n9776_), .A2(new_n10227_), .B(new_n10242_), .ZN(new_n10243_));
  OAI21_X1   g09959(.A1(new_n10220_), .A2(new_n10221_), .B(new_n10218_), .ZN(new_n10244_));
  NAND3_X1   g09960(.A1(new_n10201_), .A2(new_n10210_), .A3(new_n10224_), .ZN(new_n10245_));
  NAND2_X1   g09961(.A1(new_n10244_), .A2(new_n10245_), .ZN(new_n10246_));
  NAND3_X1   g09962(.A1(new_n10246_), .A2(new_n10117_), .A3(new_n9777_), .ZN(new_n10247_));
  NAND2_X1   g09963(.A1(new_n10243_), .A2(new_n10247_), .ZN(new_n10248_));
  NAND3_X1   g09964(.A1(new_n10241_), .A2(new_n9811_), .A3(new_n10248_), .ZN(new_n10249_));
  INV_X1     g09965(.I(new_n10236_), .ZN(new_n10250_));
  NAND3_X1   g09966(.A1(new_n10249_), .A2(new_n10240_), .A3(new_n10250_), .ZN(new_n10251_));
  OAI22_X1   g09967(.A1(new_n5420_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n5107_), .ZN(new_n10252_));
  OAI21_X1   g09968(.A1(new_n1017_), .A2(new_n5112_), .B(new_n10252_), .ZN(new_n10253_));
  AOI21_X1   g09969(.A1(new_n10253_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n10254_));
  XNOR2_X1   g09970(.A1(new_n1196_), .A2(new_n10254_), .ZN(new_n10255_));
  INV_X1     g09971(.I(new_n10255_), .ZN(new_n10256_));
  NAND3_X1   g09972(.A1(new_n10237_), .A2(new_n10251_), .A3(new_n10256_), .ZN(new_n10257_));
  AOI21_X1   g09973(.A1(new_n10249_), .A2(new_n10250_), .B(new_n10240_), .ZN(new_n10258_));
  NOR3_X1    g09974(.A1(new_n10233_), .A2(new_n9702_), .A3(new_n10236_), .ZN(new_n10259_));
  OAI21_X1   g09975(.A1(new_n10258_), .A2(new_n10259_), .B(new_n10255_), .ZN(new_n10260_));
  NAND2_X1   g09976(.A1(new_n10260_), .A2(new_n10257_), .ZN(new_n10261_));
  NAND3_X1   g09977(.A1(new_n10114_), .A2(new_n10113_), .A3(new_n10261_), .ZN(new_n10262_));
  NOR3_X1    g09978(.A1(new_n9823_), .A2(new_n9817_), .A3(new_n9821_), .ZN(new_n10263_));
  OAI21_X1   g09979(.A1(new_n10258_), .A2(new_n10259_), .B(new_n10256_), .ZN(new_n10264_));
  NAND3_X1   g09980(.A1(new_n10237_), .A2(new_n10251_), .A3(new_n10255_), .ZN(new_n10265_));
  NAND2_X1   g09981(.A1(new_n10264_), .A2(new_n10265_), .ZN(new_n10266_));
  OAI21_X1   g09982(.A1(new_n10263_), .A2(new_n10112_), .B(new_n10266_), .ZN(new_n10267_));
  OAI22_X1   g09983(.A1(new_n4072_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n4067_), .ZN(new_n10268_));
  OAI21_X1   g09984(.A1(new_n1294_), .A2(new_n4318_), .B(new_n10268_), .ZN(new_n10269_));
  AOI21_X1   g09985(.A1(new_n10269_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n10270_));
  XOR2_X1    g09986(.A1(new_n1530_), .A2(new_n10270_), .Z(new_n10271_));
  AOI21_X1   g09987(.A1(new_n10267_), .A2(new_n10262_), .B(new_n10271_), .ZN(new_n10272_));
  NOR3_X1    g09988(.A1(new_n10258_), .A2(new_n10259_), .A3(new_n10255_), .ZN(new_n10273_));
  AOI21_X1   g09989(.A1(new_n10237_), .A2(new_n10251_), .B(new_n10256_), .ZN(new_n10274_));
  NOR2_X1    g09990(.A1(new_n10274_), .A2(new_n10273_), .ZN(new_n10275_));
  NOR3_X1    g09991(.A1(new_n10263_), .A2(new_n10112_), .A3(new_n10275_), .ZN(new_n10276_));
  AOI22_X1   g09992(.A1(new_n10114_), .A2(new_n10113_), .B1(new_n10264_), .B2(new_n10265_), .ZN(new_n10277_));
  INV_X1     g09993(.I(new_n10271_), .ZN(new_n10278_));
  NOR3_X1    g09994(.A1(new_n10277_), .A2(new_n10276_), .A3(new_n10278_), .ZN(new_n10279_));
  OAI22_X1   g09995(.A1(new_n1803_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n1936_), .ZN(new_n10280_));
  OAI21_X1   g09996(.A1(new_n1634_), .A2(new_n3569_), .B(new_n10280_), .ZN(new_n10281_));
  AOI21_X1   g09997(.A1(new_n10281_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n10282_));
  XNOR2_X1   g09998(.A1(new_n1940_), .A2(new_n10282_), .ZN(new_n10283_));
  INV_X1     g09999(.I(new_n10283_), .ZN(new_n10284_));
  OAI21_X1   g10000(.A1(new_n10279_), .A2(new_n10272_), .B(new_n10284_), .ZN(new_n10285_));
  OAI21_X1   g10001(.A1(new_n10277_), .A2(new_n10276_), .B(new_n10278_), .ZN(new_n10286_));
  NAND3_X1   g10002(.A1(new_n10267_), .A2(new_n10262_), .A3(new_n10271_), .ZN(new_n10287_));
  NAND3_X1   g10003(.A1(new_n10286_), .A2(new_n10287_), .A3(new_n10283_), .ZN(new_n10288_));
  AOI22_X1   g10004(.A1(new_n10285_), .A2(new_n10288_), .B1(new_n10110_), .B2(new_n9861_), .ZN(new_n10289_));
  OAI21_X1   g10005(.A1(new_n9849_), .A2(new_n9844_), .B(new_n9861_), .ZN(new_n10290_));
  NAND3_X1   g10006(.A1(new_n10286_), .A2(new_n10287_), .A3(new_n10284_), .ZN(new_n10291_));
  OAI21_X1   g10007(.A1(new_n10279_), .A2(new_n10272_), .B(new_n10283_), .ZN(new_n10292_));
  AOI21_X1   g10008(.A1(new_n10291_), .A2(new_n10292_), .B(new_n10290_), .ZN(new_n10293_));
  NOR2_X1    g10009(.A1(new_n10293_), .A2(new_n10289_), .ZN(new_n10294_));
  NOR3_X1    g10010(.A1(new_n9863_), .A2(new_n9864_), .A3(new_n9858_), .ZN(new_n10295_));
  AOI21_X1   g10011(.A1(new_n9845_), .A2(new_n9853_), .B(new_n9859_), .ZN(new_n10296_));
  NOR2_X1    g10012(.A1(new_n10295_), .A2(new_n10296_), .ZN(new_n10297_));
  NOR3_X1    g10013(.A1(new_n10297_), .A2(new_n10294_), .A3(new_n9884_), .ZN(new_n10298_));
  AOI21_X1   g10014(.A1(new_n9698_), .A2(new_n9862_), .B(new_n9840_), .ZN(new_n10299_));
  NOR2_X1    g10015(.A1(new_n10279_), .A2(new_n10272_), .ZN(new_n10300_));
  NOR2_X1    g10016(.A1(new_n9865_), .A2(new_n9858_), .ZN(new_n10301_));
  OAI21_X1   g10017(.A1(new_n10298_), .A2(new_n10301_), .B(new_n10105_), .ZN(new_n10302_));
  NAND3_X1   g10018(.A1(new_n9361_), .A2(new_n9482_), .A3(new_n9696_), .ZN(new_n10303_));
  AOI21_X1   g10019(.A1(new_n10303_), .A2(new_n9695_), .B(new_n9844_), .ZN(new_n10304_));
  AOI21_X1   g10020(.A1(new_n10286_), .A2(new_n10287_), .B(new_n10283_), .ZN(new_n10305_));
  NOR3_X1    g10021(.A1(new_n10279_), .A2(new_n10272_), .A3(new_n10284_), .ZN(new_n10306_));
  OAI22_X1   g10022(.A1(new_n10305_), .A2(new_n10306_), .B1(new_n10304_), .B2(new_n9840_), .ZN(new_n10307_));
  NOR3_X1    g10023(.A1(new_n10279_), .A2(new_n10272_), .A3(new_n10283_), .ZN(new_n10308_));
  AOI21_X1   g10024(.A1(new_n10286_), .A2(new_n10287_), .B(new_n10284_), .ZN(new_n10309_));
  OAI21_X1   g10025(.A1(new_n10308_), .A2(new_n10309_), .B(new_n10299_), .ZN(new_n10310_));
  NAND2_X1   g10026(.A1(new_n10310_), .A2(new_n10307_), .ZN(new_n10311_));
  NAND3_X1   g10027(.A1(new_n9845_), .A2(new_n9853_), .A3(new_n9859_), .ZN(new_n10312_));
  OAI21_X1   g10028(.A1(new_n9863_), .A2(new_n9864_), .B(new_n9858_), .ZN(new_n10313_));
  NAND2_X1   g10029(.A1(new_n10313_), .A2(new_n10312_), .ZN(new_n10314_));
  NAND3_X1   g10030(.A1(new_n10314_), .A2(new_n10311_), .A3(new_n9860_), .ZN(new_n10315_));
  INV_X1     g10031(.I(new_n10301_), .ZN(new_n10316_));
  NAND3_X1   g10032(.A1(new_n10315_), .A2(new_n9888_), .A3(new_n10316_), .ZN(new_n10317_));
  OAI22_X1   g10033(.A1(new_n2281_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n2439_), .ZN(new_n10318_));
  OAI21_X1   g10034(.A1(new_n2102_), .A2(new_n2884_), .B(new_n10318_), .ZN(new_n10319_));
  AOI21_X1   g10035(.A1(new_n10319_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n10320_));
  XNOR2_X1   g10036(.A1(new_n2443_), .A2(new_n10320_), .ZN(new_n10321_));
  INV_X1     g10037(.I(new_n10321_), .ZN(new_n10322_));
  NAND3_X1   g10038(.A1(new_n10302_), .A2(new_n10317_), .A3(new_n10322_), .ZN(new_n10323_));
  AOI21_X1   g10039(.A1(new_n10315_), .A2(new_n10316_), .B(new_n9888_), .ZN(new_n10324_));
  NOR3_X1    g10040(.A1(new_n10298_), .A2(new_n10105_), .A3(new_n10301_), .ZN(new_n10325_));
  OAI21_X1   g10041(.A1(new_n10325_), .A2(new_n10324_), .B(new_n10321_), .ZN(new_n10326_));
  NAND3_X1   g10042(.A1(new_n10326_), .A2(new_n10323_), .A3(new_n10108_), .ZN(new_n10327_));
  NAND3_X1   g10043(.A1(new_n10101_), .A2(new_n10327_), .A3(new_n9893_), .ZN(new_n10328_));
  NAND2_X1   g10044(.A1(new_n9897_), .A2(new_n9895_), .ZN(new_n10329_));
  NAND2_X1   g10045(.A1(new_n9886_), .A2(new_n9888_), .ZN(new_n10330_));
  INV_X1     g10046(.I(new_n10107_), .ZN(new_n10331_));
  AOI21_X1   g10047(.A1(new_n10331_), .A2(new_n10330_), .B(new_n9890_), .ZN(new_n10332_));
  NOR3_X1    g10048(.A1(new_n10325_), .A2(new_n10324_), .A3(new_n10321_), .ZN(new_n10333_));
  AOI21_X1   g10049(.A1(new_n10302_), .A2(new_n10317_), .B(new_n10322_), .ZN(new_n10334_));
  NOR3_X1    g10050(.A1(new_n10332_), .A2(new_n10333_), .A3(new_n10334_), .ZN(new_n10335_));
  OAI21_X1   g10051(.A1(new_n10335_), .A2(new_n9903_), .B(new_n10329_), .ZN(new_n10336_));
  OAI22_X1   g10052(.A1(new_n2171_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n2166_), .ZN(new_n10337_));
  OAI21_X1   g10053(.A1(new_n2643_), .A2(new_n2322_), .B(new_n10337_), .ZN(new_n10338_));
  AOI21_X1   g10054(.A1(new_n10338_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n10339_));
  XNOR2_X1   g10055(.A1(new_n3022_), .A2(new_n10339_), .ZN(new_n10340_));
  AOI21_X1   g10056(.A1(new_n10336_), .A2(new_n10328_), .B(new_n10340_), .ZN(new_n10341_));
  NOR3_X1    g10057(.A1(new_n10335_), .A2(new_n10329_), .A3(new_n9903_), .ZN(new_n10342_));
  AOI21_X1   g10058(.A1(new_n9893_), .A2(new_n10327_), .B(new_n10101_), .ZN(new_n10343_));
  INV_X1     g10059(.I(new_n10340_), .ZN(new_n10344_));
  NOR3_X1    g10060(.A1(new_n10343_), .A2(new_n10342_), .A3(new_n10344_), .ZN(new_n10345_));
  OAI21_X1   g10061(.A1(new_n10345_), .A2(new_n10341_), .B(new_n9914_), .ZN(new_n10346_));
  NOR2_X1    g10062(.A1(new_n10346_), .A2(new_n10100_), .ZN(new_n10347_));
  OAI21_X1   g10063(.A1(new_n10343_), .A2(new_n10342_), .B(new_n10344_), .ZN(new_n10348_));
  NAND3_X1   g10064(.A1(new_n10336_), .A2(new_n10328_), .A3(new_n10340_), .ZN(new_n10349_));
  NAND2_X1   g10065(.A1(new_n10348_), .A2(new_n10349_), .ZN(new_n10350_));
  NOR2_X1    g10066(.A1(new_n10099_), .A2(new_n9908_), .ZN(new_n10352_));
  OAI21_X1   g10067(.A1(new_n10347_), .A2(new_n10352_), .B(new_n10098_), .ZN(new_n10353_));
  INV_X1     g10068(.I(new_n10100_), .ZN(new_n10354_));
  NAND3_X1   g10069(.A1(new_n10350_), .A2(new_n9914_), .A3(new_n10354_), .ZN(new_n10355_));
  INV_X1     g10070(.I(new_n10352_), .ZN(new_n10356_));
  NAND3_X1   g10071(.A1(new_n10355_), .A2(new_n9691_), .A3(new_n10356_), .ZN(new_n10357_));
  OAI22_X1   g10072(.A1(new_n1712_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n1707_), .ZN(new_n10358_));
  OAI21_X1   g10073(.A1(new_n3260_), .A2(new_n1850_), .B(new_n10358_), .ZN(new_n10359_));
  AOI21_X1   g10074(.A1(new_n10359_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n10360_));
  XOR2_X1    g10075(.A1(new_n3722_), .A2(new_n10360_), .Z(new_n10361_));
  AOI21_X1   g10076(.A1(new_n10353_), .A2(new_n10357_), .B(new_n10361_), .ZN(new_n10362_));
  AOI21_X1   g10077(.A1(new_n10355_), .A2(new_n10356_), .B(new_n9691_), .ZN(new_n10363_));
  NOR3_X1    g10078(.A1(new_n10347_), .A2(new_n10098_), .A3(new_n10352_), .ZN(new_n10364_));
  INV_X1     g10079(.I(new_n10361_), .ZN(new_n10365_));
  NOR3_X1    g10080(.A1(new_n10364_), .A2(new_n10363_), .A3(new_n10365_), .ZN(new_n10366_));
  NOR3_X1    g10081(.A1(new_n10366_), .A2(new_n10362_), .A3(new_n10096_), .ZN(new_n10367_));
  NOR3_X1    g10082(.A1(new_n10367_), .A2(new_n9686_), .A3(new_n9923_), .ZN(new_n10368_));
  INV_X1     g10083(.I(new_n10093_), .ZN(new_n10369_));
  OAI21_X1   g10084(.A1(new_n10369_), .A2(new_n10094_), .B(new_n9918_), .ZN(new_n10370_));
  OAI21_X1   g10085(.A1(new_n10364_), .A2(new_n10363_), .B(new_n10365_), .ZN(new_n10371_));
  NAND3_X1   g10086(.A1(new_n10353_), .A2(new_n10357_), .A3(new_n10361_), .ZN(new_n10372_));
  NAND3_X1   g10087(.A1(new_n10371_), .A2(new_n10372_), .A3(new_n10370_), .ZN(new_n10373_));
  AOI21_X1   g10088(.A1(new_n10373_), .A2(new_n9930_), .B(new_n9936_), .ZN(new_n10374_));
  OAI22_X1   g10089(.A1(new_n1347_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n1344_), .ZN(new_n10375_));
  OAI21_X1   g10090(.A1(new_n3989_), .A2(new_n1457_), .B(new_n10375_), .ZN(new_n10376_));
  AOI21_X1   g10091(.A1(new_n10376_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n10377_));
  XOR2_X1    g10092(.A1(new_n4499_), .A2(new_n10377_), .Z(new_n10378_));
  NOR3_X1    g10093(.A1(new_n10374_), .A2(new_n10368_), .A3(new_n10378_), .ZN(new_n10379_));
  NAND3_X1   g10094(.A1(new_n10373_), .A2(new_n9936_), .A3(new_n9930_), .ZN(new_n10380_));
  OAI21_X1   g10095(.A1(new_n10367_), .A2(new_n9923_), .B(new_n9686_), .ZN(new_n10381_));
  INV_X1     g10096(.I(new_n10378_), .ZN(new_n10382_));
  AOI21_X1   g10097(.A1(new_n10381_), .A2(new_n10380_), .B(new_n10382_), .ZN(new_n10383_));
  NOR3_X1    g10098(.A1(new_n10379_), .A2(new_n10383_), .A3(new_n10092_), .ZN(new_n10384_));
  NOR3_X1    g10099(.A1(new_n10384_), .A2(new_n9681_), .A3(new_n10087_), .ZN(new_n10385_));
  NOR2_X1    g10100(.A1(new_n9686_), .A2(new_n9923_), .ZN(new_n10386_));
  NOR2_X1    g10101(.A1(new_n9936_), .A2(new_n9930_), .ZN(new_n10387_));
  OAI21_X1   g10102(.A1(new_n10387_), .A2(new_n10386_), .B(new_n9927_), .ZN(new_n10388_));
  NAND3_X1   g10103(.A1(new_n10381_), .A2(new_n10380_), .A3(new_n10382_), .ZN(new_n10389_));
  OAI21_X1   g10104(.A1(new_n10374_), .A2(new_n10368_), .B(new_n10378_), .ZN(new_n10390_));
  NAND3_X1   g10105(.A1(new_n10390_), .A2(new_n10389_), .A3(new_n10388_), .ZN(new_n10391_));
  AOI21_X1   g10106(.A1(new_n10391_), .A2(new_n9940_), .B(new_n10085_), .ZN(new_n10392_));
  OAI22_X1   g10107(.A1(new_n1055_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n1061_), .ZN(new_n10393_));
  OAI21_X1   g10108(.A1(new_n4774_), .A2(new_n1332_), .B(new_n10393_), .ZN(new_n10394_));
  AOI21_X1   g10109(.A1(new_n10394_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n10395_));
  XNOR2_X1   g10110(.A1(new_n5357_), .A2(new_n10395_), .ZN(new_n10396_));
  NOR3_X1    g10111(.A1(new_n10385_), .A2(new_n10392_), .A3(new_n10396_), .ZN(new_n10397_));
  NAND3_X1   g10112(.A1(new_n10391_), .A2(new_n10085_), .A3(new_n9940_), .ZN(new_n10398_));
  OAI21_X1   g10113(.A1(new_n10384_), .A2(new_n10087_), .B(new_n9681_), .ZN(new_n10399_));
  INV_X1     g10114(.I(new_n10396_), .ZN(new_n10400_));
  AOI21_X1   g10115(.A1(new_n10399_), .A2(new_n10398_), .B(new_n10400_), .ZN(new_n10401_));
  NOR3_X1    g10116(.A1(new_n10397_), .A2(new_n10401_), .A3(new_n10089_), .ZN(new_n10402_));
  NOR3_X1    g10117(.A1(new_n10402_), .A2(new_n10080_), .A3(new_n9677_), .ZN(new_n10403_));
  NOR2_X1    g10118(.A1(new_n9681_), .A2(new_n10087_), .ZN(new_n10404_));
  NOR2_X1    g10119(.A1(new_n10085_), .A2(new_n9940_), .ZN(new_n10405_));
  OAI21_X1   g10120(.A1(new_n10404_), .A2(new_n10405_), .B(new_n9944_), .ZN(new_n10406_));
  NAND3_X1   g10121(.A1(new_n10399_), .A2(new_n10398_), .A3(new_n10400_), .ZN(new_n10407_));
  OAI21_X1   g10122(.A1(new_n10385_), .A2(new_n10392_), .B(new_n10396_), .ZN(new_n10408_));
  NAND3_X1   g10123(.A1(new_n10408_), .A2(new_n10407_), .A3(new_n10406_), .ZN(new_n10409_));
  AOI21_X1   g10124(.A1(new_n10409_), .A2(new_n9951_), .B(new_n9960_), .ZN(new_n10410_));
  OAI22_X1   g10125(.A1(new_n970_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n820_), .ZN(new_n10411_));
  OAI21_X1   g10126(.A1(new_n5913_), .A2(new_n894_), .B(new_n10411_), .ZN(new_n10412_));
  AOI21_X1   g10127(.A1(new_n10412_), .A2(new_n827_), .B(new_n970_), .ZN(new_n10413_));
  XOR2_X1    g10128(.A1(new_n6233_), .A2(new_n10413_), .Z(new_n10414_));
  NOR3_X1    g10129(.A1(new_n10403_), .A2(new_n10410_), .A3(new_n10414_), .ZN(new_n10415_));
  NAND3_X1   g10130(.A1(new_n10409_), .A2(new_n9960_), .A3(new_n9951_), .ZN(new_n10416_));
  OAI21_X1   g10131(.A1(new_n10402_), .A2(new_n10080_), .B(new_n9677_), .ZN(new_n10417_));
  INV_X1     g10132(.I(new_n10414_), .ZN(new_n10418_));
  AOI21_X1   g10133(.A1(new_n10417_), .A2(new_n10416_), .B(new_n10418_), .ZN(new_n10419_));
  NOR3_X1    g10134(.A1(new_n10415_), .A2(new_n10419_), .A3(new_n10082_), .ZN(new_n10420_));
  NOR3_X1    g10135(.A1(new_n10420_), .A2(new_n9972_), .A3(new_n9969_), .ZN(new_n10421_));
  NOR2_X1    g10136(.A1(new_n10080_), .A2(new_n9677_), .ZN(new_n10422_));
  NOR2_X1    g10137(.A1(new_n9960_), .A2(new_n9951_), .ZN(new_n10423_));
  OAI21_X1   g10138(.A1(new_n10422_), .A2(new_n10423_), .B(new_n9955_), .ZN(new_n10424_));
  NAND3_X1   g10139(.A1(new_n10417_), .A2(new_n10416_), .A3(new_n10418_), .ZN(new_n10425_));
  OAI21_X1   g10140(.A1(new_n10403_), .A2(new_n10410_), .B(new_n10414_), .ZN(new_n10426_));
  NAND3_X1   g10141(.A1(new_n10426_), .A2(new_n10425_), .A3(new_n10424_), .ZN(new_n10427_));
  AOI21_X1   g10142(.A1(new_n10427_), .A2(new_n9964_), .B(new_n9673_), .ZN(new_n10428_));
  NOR2_X1    g10143(.A1(new_n10428_), .A2(new_n10421_), .ZN(new_n10429_));
  AOI21_X1   g10144(.A1(new_n9668_), .A2(new_n9666_), .B(new_n9981_), .ZN(new_n10430_));
  OAI22_X1   g10145(.A1(new_n448_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n450_), .ZN(new_n10431_));
  OAI21_X1   g10146(.A1(new_n7864_), .A2(new_n496_), .B(new_n10431_), .ZN(new_n10432_));
  AOI21_X1   g10147(.A1(new_n10432_), .A2(new_n452_), .B(new_n448_), .ZN(new_n10433_));
  XOR2_X1    g10148(.A1(new_n8217_), .A2(new_n10433_), .Z(new_n10434_));
  NOR3_X1    g10149(.A1(new_n10430_), .A2(new_n9979_), .A3(new_n10434_), .ZN(new_n10435_));
  INV_X1     g10150(.I(new_n9979_), .ZN(new_n10436_));
  INV_X1     g10151(.I(new_n9981_), .ZN(new_n10437_));
  OAI21_X1   g10152(.A1(new_n9984_), .A2(new_n9665_), .B(new_n10437_), .ZN(new_n10438_));
  INV_X1     g10153(.I(new_n10434_), .ZN(new_n10439_));
  AOI21_X1   g10154(.A1(new_n10438_), .A2(new_n10436_), .B(new_n10439_), .ZN(new_n10440_));
  OAI21_X1   g10155(.A1(new_n10440_), .A2(new_n10435_), .B(new_n10429_), .ZN(new_n10441_));
  INV_X1     g10156(.I(new_n10429_), .ZN(new_n10442_));
  NAND3_X1   g10157(.A1(new_n10438_), .A2(new_n10436_), .A3(new_n10439_), .ZN(new_n10443_));
  OAI21_X1   g10158(.A1(new_n10430_), .A2(new_n9979_), .B(new_n10434_), .ZN(new_n10444_));
  NAND3_X1   g10159(.A1(new_n10443_), .A2(new_n10444_), .A3(new_n10442_), .ZN(new_n10445_));
  AOI21_X1   g10160(.A1(new_n10441_), .A2(new_n10445_), .B(new_n10078_), .ZN(new_n10446_));
  AOI21_X1   g10161(.A1(new_n10443_), .A2(new_n10444_), .B(new_n10442_), .ZN(new_n10447_));
  NOR3_X1    g10162(.A1(new_n10440_), .A2(new_n10435_), .A3(new_n10429_), .ZN(new_n10448_));
  NOR3_X1    g10163(.A1(new_n10448_), .A2(new_n10447_), .A3(new_n10077_), .ZN(new_n10449_));
  INV_X1     g10164(.I(new_n9991_), .ZN(new_n10450_));
  NAND3_X1   g10165(.A1(new_n9982_), .A2(new_n9987_), .A3(new_n10450_), .ZN(new_n10451_));
  NAND2_X1   g10166(.A1(new_n9982_), .A2(new_n9987_), .ZN(new_n10452_));
  NAND2_X1   g10167(.A1(new_n10452_), .A2(new_n9991_), .ZN(new_n10453_));
  NAND2_X1   g10168(.A1(new_n10453_), .A2(new_n10451_), .ZN(new_n10454_));
  OAI21_X1   g10169(.A1(new_n10449_), .A2(new_n10446_), .B(new_n10454_), .ZN(new_n10455_));
  NOR2_X1    g10170(.A1(new_n10455_), .A2(new_n9992_), .ZN(new_n10456_));
  INV_X1     g10171(.I(new_n10452_), .ZN(new_n10457_));
  OAI21_X1   g10172(.A1(new_n10448_), .A2(new_n10447_), .B(new_n10077_), .ZN(new_n10458_));
  NAND3_X1   g10173(.A1(new_n10441_), .A2(new_n10445_), .A3(new_n10078_), .ZN(new_n10459_));
  NAND2_X1   g10174(.A1(new_n10458_), .A2(new_n10459_), .ZN(new_n10460_));
  NOR2_X1    g10175(.A1(new_n10457_), .A2(new_n9991_), .ZN(new_n10462_));
  OAI21_X1   g10176(.A1(new_n10456_), .A2(new_n10462_), .B(new_n10064_), .ZN(new_n10463_));
  NAND3_X1   g10177(.A1(new_n10460_), .A2(new_n10017_), .A3(new_n10454_), .ZN(new_n10464_));
  INV_X1     g10178(.I(new_n10462_), .ZN(new_n10465_));
  NAND3_X1   g10179(.A1(new_n10464_), .A2(new_n10062_), .A3(new_n10465_), .ZN(new_n10466_));
  OAI22_X1   g10180(.A1(new_n8948_), .A2(new_n341_), .B1(new_n404_), .B2(new_n9295_), .ZN(new_n10467_));
  OAI21_X1   g10181(.A1(new_n8563_), .A2(new_n366_), .B(new_n10467_), .ZN(new_n10468_));
  AOI21_X1   g10182(.A1(new_n10468_), .A2(new_n334_), .B(new_n341_), .ZN(new_n10469_));
  XNOR2_X1   g10183(.A1(new_n9299_), .A2(new_n10469_), .ZN(new_n10470_));
  AOI21_X1   g10184(.A1(new_n10463_), .A2(new_n10466_), .B(new_n10470_), .ZN(new_n10471_));
  XOR2_X1    g10185(.A1(new_n10073_), .A2(new_n10471_), .Z(new_n10472_));
  XOR2_X1    g10186(.A1(new_n10472_), .A2(new_n10066_), .Z(new_n10473_));
  XNOR2_X1   g10187(.A1(\b[51] ), .A2(\b[53] ), .ZN(new_n10474_));
  NOR2_X1    g10188(.A1(new_n10474_), .A2(new_n10030_), .ZN(new_n10475_));
  XOR2_X1    g10189(.A1(new_n10029_), .A2(new_n10475_), .Z(new_n10476_));
  INV_X1     g10190(.I(\b[53] ), .ZN(new_n10477_));
  OAI22_X1   g10191(.A1(new_n330_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n263_), .ZN(new_n10478_));
  OAI21_X1   g10192(.A1(new_n10025_), .A2(new_n289_), .B(new_n10478_), .ZN(new_n10479_));
  AOI21_X1   g10193(.A1(new_n10479_), .A2(new_n260_), .B(new_n426_), .ZN(new_n10480_));
  XOR2_X1    g10194(.A1(new_n10476_), .A2(new_n10480_), .Z(new_n10481_));
  INV_X1     g10195(.I(new_n10481_), .ZN(new_n10482_));
  XOR2_X1    g10196(.A1(new_n10473_), .A2(new_n10482_), .Z(new_n10483_));
  INV_X1     g10197(.I(new_n10473_), .ZN(new_n10484_));
  NAND2_X1   g10198(.A1(new_n10484_), .A2(new_n10482_), .ZN(new_n10485_));
  NAND2_X1   g10199(.A1(new_n10473_), .A2(new_n10481_), .ZN(new_n10486_));
  NAND2_X1   g10200(.A1(new_n10485_), .A2(new_n10486_), .ZN(new_n10487_));
  NAND2_X1   g10201(.A1(new_n10487_), .A2(new_n10061_), .ZN(new_n10488_));
  OAI21_X1   g10202(.A1(new_n10061_), .A2(new_n10483_), .B(new_n10488_), .ZN(\f[53] ));
  OAI22_X1   g10203(.A1(new_n9295_), .A2(new_n341_), .B1(new_n404_), .B2(new_n10025_), .ZN(new_n10490_));
  OAI21_X1   g10204(.A1(new_n8948_), .A2(new_n366_), .B(new_n10490_), .ZN(new_n10491_));
  AOI21_X1   g10205(.A1(new_n10491_), .A2(new_n334_), .B(new_n341_), .ZN(new_n10492_));
  XNOR2_X1   g10206(.A1(new_n9642_), .A2(new_n10492_), .ZN(new_n10493_));
  INV_X1     g10207(.I(new_n10493_), .ZN(new_n10494_));
  NAND2_X1   g10208(.A1(new_n10438_), .A2(new_n10436_), .ZN(new_n10495_));
  NOR2_X1    g10209(.A1(new_n10495_), .A2(new_n10429_), .ZN(new_n10496_));
  NOR2_X1    g10210(.A1(new_n10430_), .A2(new_n9979_), .ZN(new_n10497_));
  NOR2_X1    g10211(.A1(new_n10497_), .A2(new_n10442_), .ZN(new_n10498_));
  OAI21_X1   g10212(.A1(new_n10496_), .A2(new_n10498_), .B(new_n10077_), .ZN(new_n10499_));
  NAND2_X1   g10213(.A1(new_n10497_), .A2(new_n10442_), .ZN(new_n10500_));
  NAND2_X1   g10214(.A1(new_n10495_), .A2(new_n10429_), .ZN(new_n10501_));
  NAND3_X1   g10215(.A1(new_n10501_), .A2(new_n10500_), .A3(new_n10078_), .ZN(new_n10502_));
  AOI21_X1   g10216(.A1(new_n10499_), .A2(new_n10502_), .B(new_n10434_), .ZN(new_n10503_));
  AOI21_X1   g10217(.A1(new_n10460_), .A2(new_n10450_), .B(new_n10452_), .ZN(new_n10504_));
  OAI21_X1   g10218(.A1(new_n10460_), .A2(new_n10450_), .B(new_n10062_), .ZN(new_n10505_));
  NOR2_X1    g10219(.A1(new_n10429_), .A2(new_n10078_), .ZN(new_n10506_));
  NAND3_X1   g10220(.A1(new_n10427_), .A2(new_n9964_), .A3(new_n9673_), .ZN(new_n10507_));
  OAI21_X1   g10221(.A1(new_n10420_), .A2(new_n9972_), .B(new_n9969_), .ZN(new_n10508_));
  AOI21_X1   g10222(.A1(new_n10507_), .A2(new_n10508_), .B(new_n10077_), .ZN(new_n10509_));
  NOR3_X1    g10223(.A1(new_n10428_), .A2(new_n10421_), .A3(new_n10078_), .ZN(new_n10510_));
  OAI21_X1   g10224(.A1(new_n10509_), .A2(new_n10510_), .B(new_n9974_), .ZN(new_n10511_));
  NAND2_X1   g10225(.A1(new_n10511_), .A2(new_n9978_), .ZN(new_n10512_));
  INV_X1     g10226(.I(new_n10512_), .ZN(new_n10513_));
  OR2_X2     g10227(.A1(new_n10509_), .A2(new_n10510_), .Z(new_n10514_));
  OAI21_X1   g10228(.A1(new_n9974_), .A2(new_n10514_), .B(new_n9669_), .ZN(new_n10515_));
  AOI21_X1   g10229(.A1(new_n10426_), .A2(new_n10425_), .B(new_n10424_), .ZN(new_n10516_));
  OAI21_X1   g10230(.A1(new_n10516_), .A2(new_n9964_), .B(new_n9969_), .ZN(new_n10517_));
  OAI21_X1   g10231(.A1(new_n10397_), .A2(new_n10401_), .B(new_n10089_), .ZN(new_n10518_));
  AOI21_X1   g10232(.A1(new_n10518_), .A2(new_n10080_), .B(new_n9960_), .ZN(new_n10519_));
  AOI21_X1   g10233(.A1(new_n10390_), .A2(new_n10389_), .B(new_n10388_), .ZN(new_n10520_));
  OAI21_X1   g10234(.A1(new_n10520_), .A2(new_n9940_), .B(new_n9681_), .ZN(new_n10521_));
  OAI21_X1   g10235(.A1(new_n10364_), .A2(new_n10363_), .B(new_n10361_), .ZN(new_n10522_));
  OAI21_X1   g10236(.A1(new_n10366_), .A2(new_n10362_), .B(new_n10096_), .ZN(new_n10523_));
  AOI21_X1   g10237(.A1(new_n10523_), .A2(new_n9923_), .B(new_n9936_), .ZN(new_n10524_));
  OAI21_X1   g10238(.A1(new_n10343_), .A2(new_n10342_), .B(new_n10340_), .ZN(new_n10525_));
  INV_X1     g10239(.I(new_n10525_), .ZN(new_n10526_));
  INV_X1     g10240(.I(new_n10099_), .ZN(new_n10527_));
  AOI21_X1   g10241(.A1(new_n10350_), .A2(new_n9909_), .B(new_n10527_), .ZN(new_n10528_));
  OAI21_X1   g10242(.A1(new_n9909_), .A2(new_n10350_), .B(new_n9691_), .ZN(new_n10529_));
  NOR2_X1    g10243(.A1(new_n10325_), .A2(new_n10324_), .ZN(new_n10530_));
  NAND2_X1   g10244(.A1(new_n10530_), .A2(new_n10321_), .ZN(new_n10531_));
  AOI21_X1   g10245(.A1(new_n10326_), .A2(new_n10323_), .B(new_n10108_), .ZN(new_n10532_));
  OR2_X2     g10246(.A1(new_n10532_), .A2(new_n9893_), .Z(new_n10533_));
  XOR2_X1    g10247(.A1(new_n10299_), .A2(new_n10300_), .Z(new_n10534_));
  NAND2_X1   g10248(.A1(new_n10534_), .A2(new_n10283_), .ZN(new_n10535_));
  INV_X1     g10249(.I(new_n10535_), .ZN(new_n10536_));
  OAI21_X1   g10250(.A1(new_n10293_), .A2(new_n10289_), .B(new_n9859_), .ZN(new_n10537_));
  NAND2_X1   g10251(.A1(new_n10537_), .A2(new_n9865_), .ZN(new_n10538_));
  AOI22_X1   g10252(.A1(new_n10294_), .A2(new_n9858_), .B1(new_n9875_), .B2(new_n9870_), .ZN(new_n10539_));
  NAND2_X1   g10253(.A1(new_n10539_), .A2(new_n10538_), .ZN(new_n10540_));
  NAND3_X1   g10254(.A1(new_n10114_), .A2(new_n10113_), .A3(new_n10260_), .ZN(new_n10541_));
  NOR2_X1    g10255(.A1(new_n10234_), .A2(new_n10235_), .ZN(new_n10542_));
  NAND2_X1   g10256(.A1(new_n10117_), .A2(new_n9777_), .ZN(new_n10543_));
  INV_X1     g10257(.I(new_n10235_), .ZN(new_n10544_));
  NOR2_X1    g10258(.A1(new_n10543_), .A2(new_n10544_), .ZN(new_n10545_));
  OAI21_X1   g10259(.A1(new_n10542_), .A2(new_n10545_), .B(new_n10224_), .ZN(new_n10546_));
  INV_X1     g10260(.I(new_n10546_), .ZN(new_n10547_));
  OAI21_X1   g10261(.A1(new_n10232_), .A2(new_n9796_), .B(new_n10115_), .ZN(new_n10548_));
  NOR3_X1    g10262(.A1(new_n10231_), .A2(new_n10226_), .A3(new_n9800_), .ZN(new_n10549_));
  INV_X1     g10263(.I(new_n10549_), .ZN(new_n10550_));
  NAND3_X1   g10264(.A1(new_n10548_), .A2(new_n10550_), .A3(new_n10240_), .ZN(new_n10551_));
  AOI21_X1   g10265(.A1(new_n10209_), .A2(new_n10205_), .B(new_n10200_), .ZN(new_n10552_));
  INV_X1     g10266(.I(new_n10552_), .ZN(new_n10553_));
  NAND2_X1   g10267(.A1(new_n10118_), .A2(new_n9769_), .ZN(new_n10554_));
  AOI21_X1   g10268(.A1(new_n10554_), .A2(new_n10207_), .B(new_n10192_), .ZN(new_n10555_));
  NOR2_X1    g10269(.A1(new_n10171_), .A2(new_n10169_), .ZN(new_n10556_));
  INV_X1     g10270(.I(new_n10166_), .ZN(new_n10557_));
  OAI21_X1   g10271(.A1(new_n10556_), .A2(new_n10557_), .B(new_n10161_), .ZN(new_n10558_));
  NAND2_X1   g10272(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n10559_));
  NOR2_X1    g10273(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n10560_));
  INV_X1     g10274(.I(new_n10560_), .ZN(new_n10561_));
  NAND2_X1   g10275(.A1(new_n10561_), .A2(new_n10559_), .ZN(new_n10562_));
  NAND3_X1   g10276(.A1(new_n10130_), .A2(new_n10148_), .A3(new_n10140_), .ZN(new_n10563_));
  NAND2_X1   g10277(.A1(\b[2] ), .A2(\b[3] ), .ZN(new_n10564_));
  OAI21_X1   g10278(.A1(new_n10126_), .A2(new_n10124_), .B(new_n10564_), .ZN(new_n10565_));
  NAND2_X1   g10279(.A1(new_n10145_), .A2(\b[1] ), .ZN(new_n10566_));
  AOI21_X1   g10280(.A1(new_n10566_), .A2(new_n10565_), .B(\a[53] ), .ZN(new_n10567_));
  NOR3_X1    g10281(.A1(new_n10567_), .A2(new_n403_), .A3(new_n9712_), .ZN(new_n10568_));
  INV_X1     g10282(.I(new_n10564_), .ZN(new_n10569_));
  AOI21_X1   g10283(.A1(new_n9717_), .A2(new_n9715_), .B(new_n10569_), .ZN(new_n10570_));
  NOR2_X1    g10284(.A1(new_n10137_), .A2(new_n269_), .ZN(new_n10571_));
  OAI21_X1   g10285(.A1(new_n10570_), .A2(new_n10571_), .B(new_n9718_), .ZN(new_n10572_));
  AOI21_X1   g10286(.A1(new_n10572_), .A2(new_n301_), .B(new_n9713_), .ZN(new_n10573_));
  NOR2_X1    g10287(.A1(new_n10568_), .A2(new_n10573_), .ZN(new_n10574_));
  NOR3_X1    g10288(.A1(new_n10563_), .A2(new_n10574_), .A3(new_n10562_), .ZN(new_n10575_));
  INV_X1     g10289(.I(new_n10575_), .ZN(new_n10576_));
  OAI21_X1   g10290(.A1(new_n10563_), .A2(new_n10574_), .B(new_n10562_), .ZN(new_n10577_));
  AOI21_X1   g10291(.A1(new_n10576_), .A2(new_n10577_), .B(\b[0] ), .ZN(new_n10578_));
  INV_X1     g10292(.I(new_n10577_), .ZN(new_n10579_));
  NOR3_X1    g10293(.A1(new_n10579_), .A2(new_n258_), .A3(new_n10575_), .ZN(new_n10580_));
  NOR2_X1    g10294(.A1(new_n10578_), .A2(new_n10580_), .ZN(new_n10581_));
  AOI22_X1   g10295(.A1(new_n8631_), .A2(\b[5] ), .B1(\b[6] ), .B2(new_n9382_), .ZN(new_n10582_));
  AOI21_X1   g10296(.A1(\b[4] ), .A2(new_n9731_), .B(new_n10582_), .ZN(new_n10583_));
  OAI21_X1   g10297(.A1(new_n10583_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n10584_));
  XOR2_X1    g10298(.A1(new_n556_), .A2(new_n10584_), .Z(new_n10585_));
  NOR2_X1    g10299(.A1(new_n10581_), .A2(new_n10585_), .ZN(new_n10586_));
  OAI21_X1   g10300(.A1(new_n10579_), .A2(new_n10575_), .B(new_n258_), .ZN(new_n10587_));
  NAND3_X1   g10301(.A1(new_n10576_), .A2(\b[0] ), .A3(new_n10577_), .ZN(new_n10588_));
  NAND2_X1   g10302(.A1(new_n10587_), .A2(new_n10588_), .ZN(new_n10589_));
  XOR2_X1    g10303(.A1(new_n425_), .A2(new_n10584_), .Z(new_n10590_));
  NOR2_X1    g10304(.A1(new_n10589_), .A2(new_n10590_), .ZN(new_n10591_));
  OAI21_X1   g10305(.A1(new_n10586_), .A2(new_n10591_), .B(new_n10558_), .ZN(new_n10592_));
  NAND2_X1   g10306(.A1(new_n10122_), .A2(new_n10120_), .ZN(new_n10593_));
  INV_X1     g10307(.I(new_n10161_), .ZN(new_n10594_));
  AOI21_X1   g10308(.A1(new_n10593_), .A2(new_n10166_), .B(new_n10594_), .ZN(new_n10595_));
  NOR2_X1    g10309(.A1(new_n10589_), .A2(new_n10585_), .ZN(new_n10596_));
  AOI21_X1   g10310(.A1(new_n10587_), .A2(new_n10588_), .B(new_n10590_), .ZN(new_n10597_));
  OAI21_X1   g10311(.A1(new_n10596_), .A2(new_n10597_), .B(new_n10595_), .ZN(new_n10598_));
  NAND2_X1   g10312(.A1(new_n10592_), .A2(new_n10598_), .ZN(new_n10599_));
  OAI22_X1   g10313(.A1(new_n7619_), .A2(new_n515_), .B1(new_n565_), .B2(new_n8309_), .ZN(new_n10600_));
  OAI21_X1   g10314(.A1(new_n472_), .A2(new_n7947_), .B(new_n10600_), .ZN(new_n10601_));
  AOI21_X1   g10315(.A1(new_n10601_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n10602_));
  XOR2_X1    g10316(.A1(new_n759_), .A2(new_n10602_), .Z(new_n10603_));
  INV_X1     g10317(.I(new_n10603_), .ZN(new_n10604_));
  NAND2_X1   g10318(.A1(new_n10599_), .A2(new_n10604_), .ZN(new_n10605_));
  NAND3_X1   g10319(.A1(new_n10592_), .A2(new_n10598_), .A3(new_n10603_), .ZN(new_n10606_));
  AOI21_X1   g10320(.A1(new_n10605_), .A2(new_n10606_), .B(new_n10555_), .ZN(new_n10607_));
  NOR2_X1    g10321(.A1(new_n10191_), .A2(new_n9768_), .ZN(new_n10608_));
  OAI21_X1   g10322(.A1(new_n10608_), .A2(new_n10193_), .B(new_n10206_), .ZN(new_n10609_));
  NOR2_X1    g10323(.A1(new_n10599_), .A2(new_n10603_), .ZN(new_n10610_));
  AOI21_X1   g10324(.A1(new_n10592_), .A2(new_n10598_), .B(new_n10604_), .ZN(new_n10611_));
  NOR2_X1    g10325(.A1(new_n10610_), .A2(new_n10611_), .ZN(new_n10612_));
  NOR2_X1    g10326(.A1(new_n10612_), .A2(new_n10609_), .ZN(new_n10613_));
  OAI22_X1   g10327(.A1(new_n6644_), .A2(new_n706_), .B1(new_n780_), .B2(new_n6647_), .ZN(new_n10614_));
  OAI21_X1   g10328(.A1(new_n656_), .A2(new_n7284_), .B(new_n10614_), .ZN(new_n10615_));
  AOI21_X1   g10329(.A1(new_n10615_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n10616_));
  XOR2_X1    g10330(.A1(new_n785_), .A2(new_n10616_), .Z(new_n10617_));
  INV_X1     g10331(.I(new_n10617_), .ZN(new_n10618_));
  OAI21_X1   g10332(.A1(new_n10607_), .A2(new_n10613_), .B(new_n10618_), .ZN(new_n10619_));
  AOI21_X1   g10333(.A1(new_n10234_), .A2(new_n10544_), .B(new_n10619_), .ZN(new_n10620_));
  NAND2_X1   g10334(.A1(new_n10605_), .A2(new_n10606_), .ZN(new_n10621_));
  NAND2_X1   g10335(.A1(new_n10621_), .A2(new_n10609_), .ZN(new_n10622_));
  OAI21_X1   g10336(.A1(new_n10610_), .A2(new_n10611_), .B(new_n10555_), .ZN(new_n10623_));
  AOI21_X1   g10337(.A1(new_n10623_), .A2(new_n10622_), .B(new_n10617_), .ZN(new_n10624_));
  NOR4_X1    g10338(.A1(new_n10624_), .A2(new_n10227_), .A3(new_n9776_), .A4(new_n10235_), .ZN(new_n10625_));
  OAI21_X1   g10339(.A1(new_n10620_), .A2(new_n10625_), .B(new_n10553_), .ZN(new_n10626_));
  OAI21_X1   g10340(.A1(new_n10543_), .A2(new_n10235_), .B(new_n10624_), .ZN(new_n10627_));
  NAND4_X1   g10341(.A1(new_n10619_), .A2(new_n10117_), .A3(new_n10544_), .A4(new_n9777_), .ZN(new_n10628_));
  NAND3_X1   g10342(.A1(new_n10627_), .A2(new_n10552_), .A3(new_n10628_), .ZN(new_n10629_));
  OAI22_X1   g10343(.A1(new_n5993_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n5991_), .ZN(new_n10630_));
  OAI21_X1   g10344(.A1(new_n861_), .A2(new_n5997_), .B(new_n10630_), .ZN(new_n10631_));
  AOI21_X1   g10345(.A1(new_n10631_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n10632_));
  XOR2_X1    g10346(.A1(new_n1024_), .A2(new_n10632_), .Z(new_n10633_));
  AOI21_X1   g10347(.A1(new_n10626_), .A2(new_n10629_), .B(new_n10633_), .ZN(new_n10634_));
  NAND2_X1   g10348(.A1(new_n10551_), .A2(new_n10634_), .ZN(new_n10635_));
  NOR2_X1    g10349(.A1(new_n9702_), .A2(new_n10549_), .ZN(new_n10636_));
  AOI21_X1   g10350(.A1(new_n10627_), .A2(new_n10628_), .B(new_n10552_), .ZN(new_n10637_));
  NOR3_X1    g10351(.A1(new_n10620_), .A2(new_n10553_), .A3(new_n10625_), .ZN(new_n10638_));
  INV_X1     g10352(.I(new_n10633_), .ZN(new_n10639_));
  OAI21_X1   g10353(.A1(new_n10638_), .A2(new_n10637_), .B(new_n10639_), .ZN(new_n10640_));
  NAND3_X1   g10354(.A1(new_n10640_), .A2(new_n10636_), .A3(new_n10548_), .ZN(new_n10641_));
  AOI21_X1   g10355(.A1(new_n10635_), .A2(new_n10641_), .B(new_n10547_), .ZN(new_n10642_));
  INV_X1     g10356(.I(new_n10115_), .ZN(new_n10643_));
  AOI21_X1   g10357(.A1(new_n10248_), .A2(new_n9800_), .B(new_n10643_), .ZN(new_n10644_));
  NOR3_X1    g10358(.A1(new_n10644_), .A2(new_n9702_), .A3(new_n10549_), .ZN(new_n10645_));
  NOR2_X1    g10359(.A1(new_n10645_), .A2(new_n10640_), .ZN(new_n10646_));
  NOR2_X1    g10360(.A1(new_n10551_), .A2(new_n10634_), .ZN(new_n10647_));
  NOR3_X1    g10361(.A1(new_n10646_), .A2(new_n10647_), .A3(new_n10546_), .ZN(new_n10648_));
  OAI22_X1   g10362(.A1(new_n5420_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n5107_), .ZN(new_n10649_));
  OAI21_X1   g10363(.A1(new_n1109_), .A2(new_n5112_), .B(new_n10649_), .ZN(new_n10650_));
  AOI21_X1   g10364(.A1(new_n10650_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n10651_));
  XOR2_X1    g10365(.A1(new_n1299_), .A2(new_n10651_), .Z(new_n10652_));
  INV_X1     g10366(.I(new_n10652_), .ZN(new_n10653_));
  OAI21_X1   g10367(.A1(new_n10648_), .A2(new_n10642_), .B(new_n10653_), .ZN(new_n10654_));
  OAI21_X1   g10368(.A1(new_n10646_), .A2(new_n10647_), .B(new_n10546_), .ZN(new_n10655_));
  NAND3_X1   g10369(.A1(new_n10635_), .A2(new_n10641_), .A3(new_n10547_), .ZN(new_n10656_));
  NAND3_X1   g10370(.A1(new_n10655_), .A2(new_n10656_), .A3(new_n10652_), .ZN(new_n10657_));
  AOI22_X1   g10371(.A1(new_n10541_), .A2(new_n10257_), .B1(new_n10654_), .B2(new_n10657_), .ZN(new_n10658_));
  NOR3_X1    g10372(.A1(new_n10263_), .A2(new_n10112_), .A3(new_n10274_), .ZN(new_n10659_));
  NOR3_X1    g10373(.A1(new_n10648_), .A2(new_n10642_), .A3(new_n10652_), .ZN(new_n10660_));
  AOI21_X1   g10374(.A1(new_n10655_), .A2(new_n10656_), .B(new_n10653_), .ZN(new_n10661_));
  NOR2_X1    g10375(.A1(new_n10660_), .A2(new_n10661_), .ZN(new_n10662_));
  NOR3_X1    g10376(.A1(new_n10662_), .A2(new_n10659_), .A3(new_n10273_), .ZN(new_n10663_));
  OAI22_X1   g10377(.A1(new_n4072_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n4067_), .ZN(new_n10664_));
  OAI21_X1   g10378(.A1(new_n1518_), .A2(new_n4318_), .B(new_n10664_), .ZN(new_n10665_));
  AOI21_X1   g10379(.A1(new_n10665_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n10666_));
  XNOR2_X1   g10380(.A1(new_n1638_), .A2(new_n10666_), .ZN(new_n10667_));
  INV_X1     g10381(.I(new_n10667_), .ZN(new_n10668_));
  OAI21_X1   g10382(.A1(new_n10663_), .A2(new_n10658_), .B(new_n10668_), .ZN(new_n10669_));
  AOI21_X1   g10383(.A1(new_n10299_), .A2(new_n10300_), .B(new_n10669_), .ZN(new_n10670_));
  NAND2_X1   g10384(.A1(new_n10286_), .A2(new_n10287_), .ZN(new_n10671_));
  NAND2_X1   g10385(.A1(new_n10654_), .A2(new_n10657_), .ZN(new_n10672_));
  OAI21_X1   g10386(.A1(new_n10273_), .A2(new_n10659_), .B(new_n10672_), .ZN(new_n10673_));
  NAND3_X1   g10387(.A1(new_n10655_), .A2(new_n10656_), .A3(new_n10653_), .ZN(new_n10674_));
  OAI21_X1   g10388(.A1(new_n10648_), .A2(new_n10642_), .B(new_n10652_), .ZN(new_n10675_));
  NAND2_X1   g10389(.A1(new_n10675_), .A2(new_n10674_), .ZN(new_n10676_));
  NAND3_X1   g10390(.A1(new_n10676_), .A2(new_n10541_), .A3(new_n10257_), .ZN(new_n10677_));
  AOI21_X1   g10391(.A1(new_n10673_), .A2(new_n10677_), .B(new_n10667_), .ZN(new_n10678_));
  NOR3_X1    g10392(.A1(new_n10290_), .A2(new_n10671_), .A3(new_n10678_), .ZN(new_n10679_));
  OAI21_X1   g10393(.A1(new_n10679_), .A2(new_n10670_), .B(new_n10287_), .ZN(new_n10680_));
  OAI21_X1   g10394(.A1(new_n10290_), .A2(new_n10671_), .B(new_n10678_), .ZN(new_n10681_));
  NAND3_X1   g10395(.A1(new_n10299_), .A2(new_n10669_), .A3(new_n10300_), .ZN(new_n10682_));
  NAND3_X1   g10396(.A1(new_n10681_), .A2(new_n10682_), .A3(new_n10279_), .ZN(new_n10683_));
  NAND2_X1   g10397(.A1(new_n10680_), .A2(new_n10683_), .ZN(new_n10684_));
  OAI22_X1   g10398(.A1(new_n1936_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n2102_), .ZN(new_n10685_));
  OAI21_X1   g10399(.A1(new_n1803_), .A2(new_n3569_), .B(new_n10685_), .ZN(new_n10686_));
  AOI21_X1   g10400(.A1(new_n10686_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n10687_));
  XOR2_X1    g10401(.A1(new_n2106_), .A2(new_n10687_), .Z(new_n10688_));
  INV_X1     g10402(.I(new_n10688_), .ZN(new_n10689_));
  NAND3_X1   g10403(.A1(new_n10540_), .A2(new_n10684_), .A3(new_n10689_), .ZN(new_n10690_));
  AOI21_X1   g10404(.A1(new_n10311_), .A2(new_n9859_), .B(new_n9854_), .ZN(new_n10691_));
  NAND3_X1   g10405(.A1(new_n10310_), .A2(new_n10307_), .A3(new_n9858_), .ZN(new_n10692_));
  INV_X1     g10406(.I(new_n10692_), .ZN(new_n10693_));
  NOR3_X1    g10407(.A1(new_n10691_), .A2(new_n10105_), .A3(new_n10693_), .ZN(new_n10694_));
  NAND2_X1   g10408(.A1(new_n10684_), .A2(new_n10689_), .ZN(new_n10695_));
  NAND2_X1   g10409(.A1(new_n10694_), .A2(new_n10695_), .ZN(new_n10696_));
  AOI21_X1   g10410(.A1(new_n10690_), .A2(new_n10696_), .B(new_n10536_), .ZN(new_n10697_));
  NAND3_X1   g10411(.A1(new_n10690_), .A2(new_n10696_), .A3(new_n10536_), .ZN(new_n10698_));
  INV_X1     g10412(.I(new_n10698_), .ZN(new_n10699_));
  OAI22_X1   g10413(.A1(new_n2439_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n2643_), .ZN(new_n10700_));
  OAI21_X1   g10414(.A1(new_n2281_), .A2(new_n2884_), .B(new_n10700_), .ZN(new_n10701_));
  AOI21_X1   g10415(.A1(new_n10701_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n10702_));
  XNOR2_X1   g10416(.A1(new_n2647_), .A2(new_n10702_), .ZN(new_n10703_));
  INV_X1     g10417(.I(new_n10703_), .ZN(new_n10704_));
  OAI21_X1   g10418(.A1(new_n10699_), .A2(new_n10697_), .B(new_n10704_), .ZN(new_n10705_));
  AOI21_X1   g10419(.A1(new_n10533_), .A2(new_n10329_), .B(new_n10705_), .ZN(new_n10706_));
  OAI21_X1   g10420(.A1(new_n10532_), .A2(new_n9893_), .B(new_n10329_), .ZN(new_n10707_));
  INV_X1     g10421(.I(new_n10697_), .ZN(new_n10708_));
  AOI21_X1   g10422(.A1(new_n10708_), .A2(new_n10698_), .B(new_n10703_), .ZN(new_n10709_));
  NOR2_X1    g10423(.A1(new_n10709_), .A2(new_n10707_), .ZN(new_n10710_));
  OAI21_X1   g10424(.A1(new_n10706_), .A2(new_n10710_), .B(new_n10531_), .ZN(new_n10711_));
  INV_X1     g10425(.I(new_n10531_), .ZN(new_n10712_));
  NAND2_X1   g10426(.A1(new_n10709_), .A2(new_n10707_), .ZN(new_n10713_));
  NAND3_X1   g10427(.A1(new_n10533_), .A2(new_n10705_), .A3(new_n10329_), .ZN(new_n10714_));
  NAND3_X1   g10428(.A1(new_n10714_), .A2(new_n10713_), .A3(new_n10712_), .ZN(new_n10715_));
  OAI22_X1   g10429(.A1(new_n2171_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n2166_), .ZN(new_n10716_));
  OAI21_X1   g10430(.A1(new_n2842_), .A2(new_n2322_), .B(new_n10716_), .ZN(new_n10717_));
  AOI21_X1   g10431(.A1(new_n10717_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n10718_));
  XNOR2_X1   g10432(.A1(new_n3264_), .A2(new_n10718_), .ZN(new_n10719_));
  AOI21_X1   g10433(.A1(new_n10711_), .A2(new_n10715_), .B(new_n10719_), .ZN(new_n10720_));
  OAI21_X1   g10434(.A1(new_n10529_), .A2(new_n10528_), .B(new_n10720_), .ZN(new_n10721_));
  OAI21_X1   g10435(.A1(new_n10345_), .A2(new_n10341_), .B(new_n9909_), .ZN(new_n10722_));
  NAND2_X1   g10436(.A1(new_n10722_), .A2(new_n10099_), .ZN(new_n10723_));
  NOR2_X1    g10437(.A1(new_n10350_), .A2(new_n9909_), .ZN(new_n10724_));
  NOR2_X1    g10438(.A1(new_n10724_), .A2(new_n10098_), .ZN(new_n10725_));
  AOI21_X1   g10439(.A1(new_n10714_), .A2(new_n10713_), .B(new_n10712_), .ZN(new_n10726_));
  NOR3_X1    g10440(.A1(new_n10706_), .A2(new_n10531_), .A3(new_n10710_), .ZN(new_n10727_));
  INV_X1     g10441(.I(new_n10719_), .ZN(new_n10728_));
  OAI21_X1   g10442(.A1(new_n10727_), .A2(new_n10726_), .B(new_n10728_), .ZN(new_n10729_));
  NAND3_X1   g10443(.A1(new_n10725_), .A2(new_n10729_), .A3(new_n10723_), .ZN(new_n10730_));
  AOI21_X1   g10444(.A1(new_n10730_), .A2(new_n10721_), .B(new_n10526_), .ZN(new_n10731_));
  AOI21_X1   g10445(.A1(new_n10725_), .A2(new_n10723_), .B(new_n10729_), .ZN(new_n10732_));
  NOR3_X1    g10446(.A1(new_n10529_), .A2(new_n10720_), .A3(new_n10528_), .ZN(new_n10733_));
  NOR3_X1    g10447(.A1(new_n10732_), .A2(new_n10733_), .A3(new_n10525_), .ZN(new_n10734_));
  OAI22_X1   g10448(.A1(new_n1712_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n1707_), .ZN(new_n10735_));
  OAI21_X1   g10449(.A1(new_n3709_), .A2(new_n1850_), .B(new_n10735_), .ZN(new_n10736_));
  AOI21_X1   g10450(.A1(new_n10736_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n10737_));
  XNOR2_X1   g10451(.A1(new_n3993_), .A2(new_n10737_), .ZN(new_n10738_));
  INV_X1     g10452(.I(new_n10738_), .ZN(new_n10739_));
  OAI21_X1   g10453(.A1(new_n10731_), .A2(new_n10734_), .B(new_n10739_), .ZN(new_n10740_));
  NOR2_X1    g10454(.A1(new_n10524_), .A2(new_n10740_), .ZN(new_n10741_));
  AOI21_X1   g10455(.A1(new_n10371_), .A2(new_n10372_), .B(new_n10370_), .ZN(new_n10742_));
  OAI21_X1   g10456(.A1(new_n10742_), .A2(new_n9930_), .B(new_n9686_), .ZN(new_n10743_));
  OAI21_X1   g10457(.A1(new_n10732_), .A2(new_n10733_), .B(new_n10525_), .ZN(new_n10744_));
  NAND3_X1   g10458(.A1(new_n10730_), .A2(new_n10721_), .A3(new_n10526_), .ZN(new_n10745_));
  AOI21_X1   g10459(.A1(new_n10744_), .A2(new_n10745_), .B(new_n10738_), .ZN(new_n10746_));
  NOR2_X1    g10460(.A1(new_n10743_), .A2(new_n10746_), .ZN(new_n10747_));
  OAI21_X1   g10461(.A1(new_n10741_), .A2(new_n10747_), .B(new_n10522_), .ZN(new_n10748_));
  INV_X1     g10462(.I(new_n10522_), .ZN(new_n10749_));
  NAND2_X1   g10463(.A1(new_n10743_), .A2(new_n10746_), .ZN(new_n10750_));
  NAND2_X1   g10464(.A1(new_n10524_), .A2(new_n10740_), .ZN(new_n10751_));
  NAND3_X1   g10465(.A1(new_n10751_), .A2(new_n10750_), .A3(new_n10749_), .ZN(new_n10752_));
  OAI22_X1   g10466(.A1(new_n1347_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n1344_), .ZN(new_n10753_));
  OAI21_X1   g10467(.A1(new_n4253_), .A2(new_n1457_), .B(new_n10753_), .ZN(new_n10754_));
  AOI21_X1   g10468(.A1(new_n10754_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n10755_));
  XNOR2_X1   g10469(.A1(new_n4778_), .A2(new_n10755_), .ZN(new_n10756_));
  AOI21_X1   g10470(.A1(new_n10748_), .A2(new_n10752_), .B(new_n10756_), .ZN(new_n10757_));
  NAND2_X1   g10471(.A1(new_n10521_), .A2(new_n10757_), .ZN(new_n10758_));
  OAI21_X1   g10472(.A1(new_n10379_), .A2(new_n10383_), .B(new_n10092_), .ZN(new_n10759_));
  AOI21_X1   g10473(.A1(new_n10759_), .A2(new_n10087_), .B(new_n10085_), .ZN(new_n10760_));
  AOI21_X1   g10474(.A1(new_n10751_), .A2(new_n10750_), .B(new_n10749_), .ZN(new_n10761_));
  NOR3_X1    g10475(.A1(new_n10741_), .A2(new_n10747_), .A3(new_n10522_), .ZN(new_n10762_));
  INV_X1     g10476(.I(new_n10756_), .ZN(new_n10763_));
  OAI21_X1   g10477(.A1(new_n10761_), .A2(new_n10762_), .B(new_n10763_), .ZN(new_n10764_));
  NAND2_X1   g10478(.A1(new_n10760_), .A2(new_n10764_), .ZN(new_n10765_));
  AOI21_X1   g10479(.A1(new_n10765_), .A2(new_n10758_), .B(new_n10383_), .ZN(new_n10766_));
  NOR2_X1    g10480(.A1(new_n10760_), .A2(new_n10764_), .ZN(new_n10767_));
  NOR2_X1    g10481(.A1(new_n10521_), .A2(new_n10757_), .ZN(new_n10768_));
  NOR3_X1    g10482(.A1(new_n10767_), .A2(new_n10768_), .A3(new_n10390_), .ZN(new_n10769_));
  OAI22_X1   g10483(.A1(new_n1055_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n1061_), .ZN(new_n10770_));
  OAI21_X1   g10484(.A1(new_n5068_), .A2(new_n1332_), .B(new_n10770_), .ZN(new_n10771_));
  AOI21_X1   g10485(.A1(new_n10771_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n10772_));
  XNOR2_X1   g10486(.A1(new_n5600_), .A2(new_n10772_), .ZN(new_n10773_));
  INV_X1     g10487(.I(new_n10773_), .ZN(new_n10774_));
  OAI21_X1   g10488(.A1(new_n10766_), .A2(new_n10769_), .B(new_n10774_), .ZN(new_n10775_));
  NOR2_X1    g10489(.A1(new_n10519_), .A2(new_n10775_), .ZN(new_n10776_));
  AOI21_X1   g10490(.A1(new_n10408_), .A2(new_n10407_), .B(new_n10406_), .ZN(new_n10777_));
  OAI21_X1   g10491(.A1(new_n10777_), .A2(new_n9951_), .B(new_n9677_), .ZN(new_n10778_));
  OAI21_X1   g10492(.A1(new_n10767_), .A2(new_n10768_), .B(new_n10390_), .ZN(new_n10779_));
  NAND3_X1   g10493(.A1(new_n10765_), .A2(new_n10758_), .A3(new_n10383_), .ZN(new_n10780_));
  AOI21_X1   g10494(.A1(new_n10779_), .A2(new_n10780_), .B(new_n10773_), .ZN(new_n10781_));
  NOR2_X1    g10495(.A1(new_n10778_), .A2(new_n10781_), .ZN(new_n10782_));
  OAI21_X1   g10496(.A1(new_n10776_), .A2(new_n10782_), .B(new_n10408_), .ZN(new_n10783_));
  NAND2_X1   g10497(.A1(new_n10778_), .A2(new_n10781_), .ZN(new_n10784_));
  NAND2_X1   g10498(.A1(new_n10519_), .A2(new_n10775_), .ZN(new_n10785_));
  NAND3_X1   g10499(.A1(new_n10785_), .A2(new_n10784_), .A3(new_n10401_), .ZN(new_n10786_));
  NAND2_X1   g10500(.A1(new_n10783_), .A2(new_n10786_), .ZN(new_n10787_));
  OAI22_X1   g10501(.A1(new_n970_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n820_), .ZN(new_n10788_));
  OAI21_X1   g10502(.A1(new_n5921_), .A2(new_n894_), .B(new_n10788_), .ZN(new_n10789_));
  AOI21_X1   g10503(.A1(new_n10789_), .A2(new_n827_), .B(new_n970_), .ZN(new_n10790_));
  XOR2_X1    g10504(.A1(new_n6543_), .A2(new_n10790_), .Z(new_n10791_));
  INV_X1     g10505(.I(new_n10791_), .ZN(new_n10792_));
  NAND3_X1   g10506(.A1(new_n10517_), .A2(new_n10787_), .A3(new_n10792_), .ZN(new_n10793_));
  INV_X1     g10507(.I(new_n10793_), .ZN(new_n10794_));
  AOI21_X1   g10508(.A1(new_n10787_), .A2(new_n10792_), .B(new_n10517_), .ZN(new_n10795_));
  OAI21_X1   g10509(.A1(new_n10794_), .A2(new_n10795_), .B(new_n10426_), .ZN(new_n10796_));
  OAI21_X1   g10510(.A1(new_n10415_), .A2(new_n10419_), .B(new_n10082_), .ZN(new_n10797_));
  AOI21_X1   g10511(.A1(new_n10797_), .A2(new_n9972_), .B(new_n9673_), .ZN(new_n10798_));
  AOI21_X1   g10512(.A1(new_n10785_), .A2(new_n10784_), .B(new_n10401_), .ZN(new_n10799_));
  NOR3_X1    g10513(.A1(new_n10776_), .A2(new_n10782_), .A3(new_n10408_), .ZN(new_n10800_));
  NOR2_X1    g10514(.A1(new_n10799_), .A2(new_n10800_), .ZN(new_n10801_));
  OAI21_X1   g10515(.A1(new_n10801_), .A2(new_n10791_), .B(new_n10798_), .ZN(new_n10802_));
  NAND3_X1   g10516(.A1(new_n10802_), .A2(new_n10793_), .A3(new_n10419_), .ZN(new_n10803_));
  OAI22_X1   g10517(.A1(new_n607_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n610_), .ZN(new_n10804_));
  OAI21_X1   g10518(.A1(new_n6847_), .A2(new_n684_), .B(new_n10804_), .ZN(new_n10805_));
  AOI21_X1   g10519(.A1(new_n10805_), .A2(new_n612_), .B(new_n607_), .ZN(new_n10806_));
  XOR2_X1    g10520(.A1(new_n7516_), .A2(new_n10806_), .Z(new_n10807_));
  AOI21_X1   g10521(.A1(new_n10796_), .A2(new_n10803_), .B(new_n10807_), .ZN(new_n10808_));
  OAI21_X1   g10522(.A1(new_n10515_), .A2(new_n10513_), .B(new_n10808_), .ZN(new_n10809_));
  NOR3_X1    g10523(.A1(new_n10509_), .A2(new_n10510_), .A3(new_n9974_), .ZN(new_n10810_));
  NOR2_X1    g10524(.A1(new_n9985_), .A2(new_n10810_), .ZN(new_n10811_));
  AOI21_X1   g10525(.A1(new_n10802_), .A2(new_n10793_), .B(new_n10419_), .ZN(new_n10812_));
  NOR3_X1    g10526(.A1(new_n10794_), .A2(new_n10795_), .A3(new_n10426_), .ZN(new_n10813_));
  INV_X1     g10527(.I(new_n10807_), .ZN(new_n10814_));
  OAI21_X1   g10528(.A1(new_n10813_), .A2(new_n10812_), .B(new_n10814_), .ZN(new_n10815_));
  NAND3_X1   g10529(.A1(new_n10811_), .A2(new_n10815_), .A3(new_n10512_), .ZN(new_n10816_));
  AOI21_X1   g10530(.A1(new_n10809_), .A2(new_n10816_), .B(new_n10506_), .ZN(new_n10817_));
  INV_X1     g10531(.I(new_n10506_), .ZN(new_n10818_));
  AOI21_X1   g10532(.A1(new_n10811_), .A2(new_n10512_), .B(new_n10815_), .ZN(new_n10819_));
  NOR3_X1    g10533(.A1(new_n10515_), .A2(new_n10513_), .A3(new_n10808_), .ZN(new_n10820_));
  NOR3_X1    g10534(.A1(new_n10820_), .A2(new_n10819_), .A3(new_n10818_), .ZN(new_n10821_));
  NOR2_X1    g10535(.A1(new_n10821_), .A2(new_n10817_), .ZN(new_n10822_));
  OAI22_X1   g10536(.A1(new_n448_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n450_), .ZN(new_n10823_));
  OAI21_X1   g10537(.A1(new_n7870_), .A2(new_n496_), .B(new_n10823_), .ZN(new_n10824_));
  AOI21_X1   g10538(.A1(new_n10824_), .A2(new_n452_), .B(new_n448_), .ZN(new_n10825_));
  XOR2_X1    g10539(.A1(new_n8568_), .A2(new_n10825_), .Z(new_n10826_));
  NOR2_X1    g10540(.A1(new_n10822_), .A2(new_n10826_), .ZN(new_n10827_));
  OAI21_X1   g10541(.A1(new_n10504_), .A2(new_n10505_), .B(new_n10827_), .ZN(new_n10828_));
  OAI21_X1   g10542(.A1(new_n10449_), .A2(new_n10446_), .B(new_n10450_), .ZN(new_n10829_));
  NAND2_X1   g10543(.A1(new_n10829_), .A2(new_n10457_), .ZN(new_n10830_));
  NOR3_X1    g10544(.A1(new_n10449_), .A2(new_n10446_), .A3(new_n10450_), .ZN(new_n10831_));
  NOR2_X1    g10545(.A1(new_n10831_), .A2(new_n10064_), .ZN(new_n10832_));
  OAI21_X1   g10546(.A1(new_n10820_), .A2(new_n10819_), .B(new_n10818_), .ZN(new_n10833_));
  NAND3_X1   g10547(.A1(new_n10809_), .A2(new_n10816_), .A3(new_n10506_), .ZN(new_n10834_));
  NAND2_X1   g10548(.A1(new_n10833_), .A2(new_n10834_), .ZN(new_n10835_));
  INV_X1     g10549(.I(new_n10826_), .ZN(new_n10836_));
  NAND2_X1   g10550(.A1(new_n10835_), .A2(new_n10836_), .ZN(new_n10837_));
  NAND3_X1   g10551(.A1(new_n10832_), .A2(new_n10830_), .A3(new_n10837_), .ZN(new_n10838_));
  AOI21_X1   g10552(.A1(new_n10838_), .A2(new_n10828_), .B(new_n10503_), .ZN(new_n10839_));
  AOI21_X1   g10553(.A1(new_n10501_), .A2(new_n10500_), .B(new_n10078_), .ZN(new_n10840_));
  NOR3_X1    g10554(.A1(new_n10496_), .A2(new_n10498_), .A3(new_n10077_), .ZN(new_n10841_));
  OAI21_X1   g10555(.A1(new_n10841_), .A2(new_n10840_), .B(new_n10439_), .ZN(new_n10842_));
  AOI21_X1   g10556(.A1(new_n10832_), .A2(new_n10830_), .B(new_n10837_), .ZN(new_n10843_));
  NOR3_X1    g10557(.A1(new_n10504_), .A2(new_n10505_), .A3(new_n10827_), .ZN(new_n10844_));
  NOR3_X1    g10558(.A1(new_n10843_), .A2(new_n10844_), .A3(new_n10842_), .ZN(new_n10845_));
  NOR2_X1    g10559(.A1(new_n10839_), .A2(new_n10845_), .ZN(new_n10846_));
  AOI21_X1   g10560(.A1(new_n10464_), .A2(new_n10465_), .B(new_n10062_), .ZN(new_n10847_));
  NOR3_X1    g10561(.A1(new_n10456_), .A2(new_n10064_), .A3(new_n10462_), .ZN(new_n10848_));
  OAI21_X1   g10562(.A1(new_n10848_), .A2(new_n10847_), .B(new_n10066_), .ZN(new_n10849_));
  NOR3_X1    g10563(.A1(new_n10848_), .A2(new_n10847_), .A3(new_n10066_), .ZN(new_n10850_));
  INV_X1     g10564(.I(new_n10071_), .ZN(new_n10851_));
  INV_X1     g10565(.I(new_n10470_), .ZN(new_n10852_));
  NAND4_X1   g10566(.A1(new_n9320_), .A2(new_n10069_), .A3(new_n10851_), .A4(new_n10852_), .ZN(new_n10853_));
  OAI21_X1   g10567(.A1(new_n10853_), .A2(new_n10850_), .B(new_n10849_), .ZN(new_n10854_));
  NOR2_X1    g10568(.A1(\b[52] ), .A2(\b[53] ), .ZN(new_n10855_));
  AOI21_X1   g10569(.A1(new_n10029_), .A2(new_n10855_), .B(new_n10025_), .ZN(new_n10856_));
  NOR2_X1    g10570(.A1(new_n10031_), .A2(new_n10477_), .ZN(new_n10857_));
  INV_X1     g10571(.I(new_n10857_), .ZN(new_n10858_));
  NOR2_X1    g10572(.A1(new_n10029_), .A2(new_n10858_), .ZN(new_n10859_));
  NOR2_X1    g10573(.A1(new_n10856_), .A2(new_n10859_), .ZN(new_n10860_));
  XNOR2_X1   g10574(.A1(\b[53] ), .A2(\b[54] ), .ZN(new_n10861_));
  INV_X1     g10575(.I(\b[54] ), .ZN(new_n10862_));
  NOR2_X1    g10576(.A1(new_n10477_), .A2(new_n10862_), .ZN(new_n10863_));
  NOR2_X1    g10577(.A1(\b[53] ), .A2(\b[54] ), .ZN(new_n10864_));
  OAI21_X1   g10578(.A1(new_n10863_), .A2(new_n10864_), .B(new_n10860_), .ZN(new_n10865_));
  OAI21_X1   g10579(.A1(new_n10860_), .A2(new_n10861_), .B(new_n10865_), .ZN(new_n10866_));
  OAI22_X1   g10580(.A1(new_n330_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n263_), .ZN(new_n10867_));
  OAI21_X1   g10581(.A1(new_n10031_), .A2(new_n289_), .B(new_n10867_), .ZN(new_n10868_));
  AOI21_X1   g10582(.A1(new_n10868_), .A2(new_n260_), .B(new_n426_), .ZN(new_n10869_));
  XNOR2_X1   g10583(.A1(new_n10866_), .A2(new_n10869_), .ZN(new_n10870_));
  NOR2_X1    g10584(.A1(new_n10854_), .A2(new_n10870_), .ZN(new_n10871_));
  INV_X1     g10585(.I(new_n10066_), .ZN(new_n10872_));
  NAND3_X1   g10586(.A1(new_n10463_), .A2(new_n10466_), .A3(new_n10872_), .ZN(new_n10873_));
  NAND4_X1   g10587(.A1(new_n10873_), .A2(new_n10072_), .A3(new_n10069_), .A4(new_n10852_), .ZN(new_n10874_));
  INV_X1     g10588(.I(new_n10870_), .ZN(new_n10875_));
  AOI21_X1   g10589(.A1(new_n10874_), .A2(new_n10849_), .B(new_n10875_), .ZN(new_n10876_));
  OAI21_X1   g10590(.A1(new_n10871_), .A2(new_n10876_), .B(new_n10846_), .ZN(new_n10877_));
  OAI21_X1   g10591(.A1(new_n10843_), .A2(new_n10844_), .B(new_n10842_), .ZN(new_n10878_));
  NAND3_X1   g10592(.A1(new_n10838_), .A2(new_n10828_), .A3(new_n10503_), .ZN(new_n10879_));
  NAND2_X1   g10593(.A1(new_n10878_), .A2(new_n10879_), .ZN(new_n10880_));
  NAND3_X1   g10594(.A1(new_n10874_), .A2(new_n10849_), .A3(new_n10875_), .ZN(new_n10881_));
  NAND2_X1   g10595(.A1(new_n10854_), .A2(new_n10870_), .ZN(new_n10882_));
  NAND3_X1   g10596(.A1(new_n10882_), .A2(new_n10881_), .A3(new_n10880_), .ZN(new_n10883_));
  AOI21_X1   g10597(.A1(new_n10877_), .A2(new_n10883_), .B(new_n10494_), .ZN(new_n10884_));
  INV_X1     g10598(.I(new_n10884_), .ZN(new_n10885_));
  NAND3_X1   g10599(.A1(new_n10877_), .A2(new_n10883_), .A3(new_n10494_), .ZN(new_n10886_));
  AOI21_X1   g10600(.A1(new_n10885_), .A2(new_n10886_), .B(new_n10483_), .ZN(new_n10887_));
  XOR2_X1    g10601(.A1(new_n10887_), .A2(new_n10485_), .Z(new_n10888_));
  XOR2_X1    g10602(.A1(new_n10888_), .A2(new_n10061_), .Z(\f[54] ));
  NOR2_X1    g10603(.A1(new_n10822_), .A2(new_n10842_), .ZN(new_n10890_));
  NOR2_X1    g10604(.A1(new_n10503_), .A2(new_n10835_), .ZN(new_n10891_));
  NOR4_X1    g10605(.A1(new_n10504_), .A2(new_n10505_), .A3(new_n10826_), .A4(new_n10891_), .ZN(new_n10892_));
  AOI21_X1   g10606(.A1(new_n10796_), .A2(new_n10803_), .B(new_n10818_), .ZN(new_n10893_));
  INV_X1     g10607(.I(new_n10893_), .ZN(new_n10894_));
  NAND3_X1   g10608(.A1(new_n10796_), .A2(new_n10818_), .A3(new_n10803_), .ZN(new_n10895_));
  NAND4_X1   g10609(.A1(new_n10811_), .A2(new_n10895_), .A3(new_n10512_), .A4(new_n10814_), .ZN(new_n10896_));
  NAND2_X1   g10610(.A1(new_n10787_), .A2(new_n10419_), .ZN(new_n10897_));
  NAND3_X1   g10611(.A1(new_n10783_), .A2(new_n10786_), .A3(new_n10426_), .ZN(new_n10898_));
  NAND3_X1   g10612(.A1(new_n10798_), .A2(new_n10898_), .A3(new_n10792_), .ZN(new_n10899_));
  NAND2_X1   g10613(.A1(new_n10779_), .A2(new_n10780_), .ZN(new_n10900_));
  NAND2_X1   g10614(.A1(new_n10900_), .A2(new_n10401_), .ZN(new_n10901_));
  NAND3_X1   g10615(.A1(new_n10779_), .A2(new_n10780_), .A3(new_n10408_), .ZN(new_n10902_));
  NAND3_X1   g10616(.A1(new_n10519_), .A2(new_n10902_), .A3(new_n10774_), .ZN(new_n10903_));
  NOR2_X1    g10617(.A1(new_n10761_), .A2(new_n10762_), .ZN(new_n10904_));
  INV_X1     g10618(.I(new_n10904_), .ZN(new_n10905_));
  AOI21_X1   g10619(.A1(new_n10904_), .A2(new_n10390_), .B(new_n10756_), .ZN(new_n10906_));
  AOI22_X1   g10620(.A1(new_n10906_), .A2(new_n10760_), .B1(new_n10383_), .B2(new_n10905_), .ZN(new_n10907_));
  NOR2_X1    g10621(.A1(new_n10731_), .A2(new_n10734_), .ZN(new_n10908_));
  NAND3_X1   g10622(.A1(new_n10744_), .A2(new_n10745_), .A3(new_n10522_), .ZN(new_n10909_));
  NAND2_X1   g10623(.A1(new_n10909_), .A2(new_n10739_), .ZN(new_n10910_));
  OAI22_X1   g10624(.A1(new_n10910_), .A2(new_n10743_), .B1(new_n10522_), .B2(new_n10908_), .ZN(new_n10911_));
  NAND2_X1   g10625(.A1(new_n10711_), .A2(new_n10715_), .ZN(new_n10912_));
  NAND2_X1   g10626(.A1(new_n10912_), .A2(new_n10526_), .ZN(new_n10913_));
  NOR2_X1    g10627(.A1(new_n10529_), .A2(new_n10528_), .ZN(new_n10914_));
  NAND3_X1   g10628(.A1(new_n10711_), .A2(new_n10715_), .A3(new_n10525_), .ZN(new_n10915_));
  NAND3_X1   g10629(.A1(new_n10914_), .A2(new_n10728_), .A3(new_n10915_), .ZN(new_n10916_));
  NAND2_X1   g10630(.A1(new_n10916_), .A2(new_n10913_), .ZN(new_n10917_));
  OAI22_X1   g10631(.A1(new_n2102_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n2281_), .ZN(new_n10918_));
  OAI21_X1   g10632(.A1(new_n1936_), .A2(new_n3569_), .B(new_n10918_), .ZN(new_n10919_));
  AOI21_X1   g10633(.A1(new_n10919_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n10920_));
  XNOR2_X1   g10634(.A1(new_n2280_), .A2(new_n10920_), .ZN(new_n10921_));
  NOR2_X1    g10635(.A1(new_n10659_), .A2(new_n10273_), .ZN(new_n10922_));
  OAI21_X1   g10636(.A1(new_n10922_), .A2(new_n10661_), .B(new_n10674_), .ZN(new_n10923_));
  OAI22_X1   g10637(.A1(new_n5993_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n5991_), .ZN(new_n10924_));
  OAI21_X1   g10638(.A1(new_n930_), .A2(new_n5997_), .B(new_n10924_), .ZN(new_n10925_));
  AOI21_X1   g10639(.A1(new_n10925_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n10926_));
  XOR2_X1    g10640(.A1(new_n1114_), .A2(new_n10926_), .Z(new_n10927_));
  INV_X1     g10641(.I(new_n10927_), .ZN(new_n10928_));
  NAND2_X1   g10642(.A1(new_n10234_), .A2(new_n10544_), .ZN(new_n10929_));
  NAND2_X1   g10643(.A1(new_n10623_), .A2(new_n10622_), .ZN(new_n10930_));
  NAND2_X1   g10644(.A1(new_n10930_), .A2(new_n10552_), .ZN(new_n10931_));
  OAI21_X1   g10645(.A1(new_n10930_), .A2(new_n10552_), .B(new_n10618_), .ZN(new_n10932_));
  OAI21_X1   g10646(.A1(new_n10929_), .A2(new_n10932_), .B(new_n10931_), .ZN(new_n10933_));
  INV_X1     g10647(.I(new_n10933_), .ZN(new_n10934_));
  NOR2_X1    g10648(.A1(new_n10638_), .A2(new_n10637_), .ZN(new_n10935_));
  NOR2_X1    g10649(.A1(new_n10551_), .A2(new_n10935_), .ZN(new_n10936_));
  XOR2_X1    g10650(.A1(new_n10543_), .A2(new_n10235_), .Z(new_n10937_));
  NAND3_X1   g10651(.A1(new_n10937_), .A2(new_n10224_), .A3(new_n10639_), .ZN(new_n10938_));
  AOI21_X1   g10652(.A1(new_n10551_), .A2(new_n10935_), .B(new_n10938_), .ZN(new_n10939_));
  INV_X1     g10653(.I(new_n10611_), .ZN(new_n10940_));
  AOI21_X1   g10654(.A1(new_n10609_), .A2(new_n10940_), .B(new_n10610_), .ZN(new_n10941_));
  NAND2_X1   g10655(.A1(new_n10581_), .A2(new_n10590_), .ZN(new_n10942_));
  OAI21_X1   g10656(.A1(new_n10578_), .A2(new_n10580_), .B(new_n10585_), .ZN(new_n10943_));
  NAND2_X1   g10657(.A1(new_n10558_), .A2(new_n10943_), .ZN(new_n10944_));
  AND3_X2    g10658(.A1(new_n10148_), .A2(new_n10130_), .A3(new_n10140_), .Z(new_n10945_));
  OR2_X2     g10659(.A1(new_n10568_), .A2(new_n10573_), .Z(new_n10946_));
  NAND2_X1   g10660(.A1(new_n10945_), .A2(new_n10946_), .ZN(new_n10947_));
  INV_X1     g10661(.I(new_n10559_), .ZN(new_n10948_));
  NOR2_X1    g10662(.A1(new_n10948_), .A2(new_n10560_), .ZN(new_n10949_));
  NOR2_X1    g10663(.A1(new_n10949_), .A2(new_n258_), .ZN(new_n10950_));
  OAI21_X1   g10664(.A1(new_n10945_), .A2(new_n10946_), .B(new_n10950_), .ZN(new_n10951_));
  NAND2_X1   g10665(.A1(new_n10951_), .A2(new_n10947_), .ZN(new_n10952_));
  AOI21_X1   g10666(.A1(new_n9717_), .A2(new_n9715_), .B(new_n326_), .ZN(new_n10953_));
  NOR2_X1    g10667(.A1(new_n10137_), .A2(new_n280_), .ZN(new_n10954_));
  OAI21_X1   g10668(.A1(new_n10953_), .A2(new_n10954_), .B(new_n9718_), .ZN(new_n10955_));
  NAND3_X1   g10669(.A1(new_n10955_), .A2(new_n807_), .A3(new_n9712_), .ZN(new_n10956_));
  INV_X1     g10670(.I(new_n326_), .ZN(new_n10957_));
  OAI21_X1   g10671(.A1(new_n10126_), .A2(new_n10124_), .B(new_n10957_), .ZN(new_n10958_));
  NAND2_X1   g10672(.A1(new_n10145_), .A2(\b[2] ), .ZN(new_n10959_));
  AOI21_X1   g10673(.A1(new_n10959_), .A2(new_n10958_), .B(\a[53] ), .ZN(new_n10960_));
  OAI21_X1   g10674(.A1(new_n10960_), .A2(new_n9713_), .B(new_n329_), .ZN(new_n10961_));
  NAND2_X1   g10675(.A1(new_n10961_), .A2(new_n10956_), .ZN(new_n10962_));
  XOR2_X1    g10676(.A1(\a[55] ), .A2(\a[56] ), .Z(new_n10963_));
  NAND2_X1   g10677(.A1(new_n10949_), .A2(new_n10963_), .ZN(new_n10964_));
  INV_X1     g10678(.I(\a[55] ), .ZN(new_n10965_));
  NAND3_X1   g10679(.A1(new_n10965_), .A2(\a[53] ), .A3(\a[54] ), .ZN(new_n10966_));
  OAI21_X1   g10680(.A1(new_n10965_), .A2(new_n10561_), .B(new_n10966_), .ZN(new_n10967_));
  XNOR2_X1   g10681(.A1(\a[55] ), .A2(\a[56] ), .ZN(new_n10968_));
  NAND3_X1   g10682(.A1(new_n10967_), .A2(new_n10949_), .A3(new_n10968_), .ZN(new_n10969_));
  NOR2_X1    g10683(.A1(new_n319_), .A2(\a[56] ), .ZN(new_n10970_));
  AOI21_X1   g10684(.A1(new_n10969_), .A2(new_n10970_), .B(new_n10964_), .ZN(new_n10971_));
  NOR2_X1    g10685(.A1(new_n10971_), .A2(new_n444_), .ZN(new_n10972_));
  INV_X1     g10686(.I(\a[56] ), .ZN(new_n10973_));
  XNOR2_X1   g10687(.A1(\a[55] ), .A2(\a[56] ), .ZN(new_n10974_));
  NOR2_X1    g10688(.A1(new_n10562_), .A2(new_n10974_), .ZN(new_n10975_));
  NOR3_X1    g10689(.A1(new_n10965_), .A2(\a[53] ), .A3(\a[54] ), .ZN(new_n10976_));
  AOI21_X1   g10690(.A1(new_n10965_), .A2(new_n10948_), .B(new_n10976_), .ZN(new_n10977_));
  XOR2_X1    g10691(.A1(\a[55] ), .A2(\a[56] ), .Z(new_n10978_));
  NOR3_X1    g10692(.A1(new_n10977_), .A2(new_n10562_), .A3(new_n10978_), .ZN(new_n10979_));
  INV_X1     g10693(.I(new_n10970_), .ZN(new_n10980_));
  OAI21_X1   g10694(.A1(new_n10979_), .A2(new_n10980_), .B(new_n10975_), .ZN(new_n10981_));
  OAI21_X1   g10695(.A1(new_n10981_), .A2(new_n271_), .B(new_n10973_), .ZN(new_n10982_));
  NOR2_X1    g10696(.A1(new_n10982_), .A2(new_n10972_), .ZN(new_n10983_));
  NOR3_X1    g10697(.A1(new_n10983_), .A2(new_n258_), .A3(new_n10562_), .ZN(new_n10984_));
  NAND2_X1   g10698(.A1(new_n10981_), .A2(new_n271_), .ZN(new_n10985_));
  AOI21_X1   g10699(.A1(new_n10971_), .A2(new_n444_), .B(\a[56] ), .ZN(new_n10986_));
  NAND2_X1   g10700(.A1(new_n10986_), .A2(new_n10985_), .ZN(new_n10987_));
  AOI21_X1   g10701(.A1(new_n10987_), .A2(\b[0] ), .B(new_n10949_), .ZN(new_n10988_));
  OAI21_X1   g10702(.A1(new_n10984_), .A2(new_n10988_), .B(new_n10962_), .ZN(new_n10989_));
  NOR3_X1    g10703(.A1(new_n10960_), .A2(new_n329_), .A3(new_n9713_), .ZN(new_n10990_));
  AOI21_X1   g10704(.A1(new_n10955_), .A2(new_n9712_), .B(new_n807_), .ZN(new_n10991_));
  NOR2_X1    g10705(.A1(new_n10990_), .A2(new_n10991_), .ZN(new_n10992_));
  NAND3_X1   g10706(.A1(new_n10987_), .A2(\b[0] ), .A3(new_n10949_), .ZN(new_n10993_));
  OAI21_X1   g10707(.A1(new_n10983_), .A2(new_n258_), .B(new_n10562_), .ZN(new_n10994_));
  NAND3_X1   g10708(.A1(new_n10994_), .A2(new_n10993_), .A3(new_n10992_), .ZN(new_n10995_));
  NAND2_X1   g10709(.A1(new_n10989_), .A2(new_n10995_), .ZN(new_n10996_));
  NAND2_X1   g10710(.A1(new_n10952_), .A2(new_n10996_), .ZN(new_n10997_));
  NOR2_X1    g10711(.A1(new_n10563_), .A2(new_n10574_), .ZN(new_n10998_));
  INV_X1     g10712(.I(new_n10950_), .ZN(new_n10999_));
  AOI21_X1   g10713(.A1(new_n10563_), .A2(new_n10574_), .B(new_n10999_), .ZN(new_n11000_));
  NOR2_X1    g10714(.A1(new_n11000_), .A2(new_n10998_), .ZN(new_n11001_));
  AOI21_X1   g10715(.A1(new_n10994_), .A2(new_n10993_), .B(new_n10962_), .ZN(new_n11002_));
  NAND3_X1   g10716(.A1(new_n10994_), .A2(new_n10993_), .A3(new_n10962_), .ZN(new_n11003_));
  INV_X1     g10717(.I(new_n11003_), .ZN(new_n11004_));
  OAI21_X1   g10718(.A1(new_n11002_), .A2(new_n11004_), .B(new_n11001_), .ZN(new_n11005_));
  NAND2_X1   g10719(.A1(new_n10997_), .A2(new_n11005_), .ZN(new_n11006_));
  AOI22_X1   g10720(.A1(new_n8631_), .A2(\b[6] ), .B1(\b[7] ), .B2(new_n9382_), .ZN(new_n11007_));
  AOI21_X1   g10721(.A1(\b[5] ), .A2(new_n9731_), .B(new_n11007_), .ZN(new_n11008_));
  OAI21_X1   g10722(.A1(new_n11008_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n11009_));
  XNOR2_X1   g10723(.A1(new_n471_), .A2(new_n11009_), .ZN(new_n11010_));
  INV_X1     g10724(.I(new_n11010_), .ZN(new_n11011_));
  NAND2_X1   g10725(.A1(new_n11006_), .A2(new_n11011_), .ZN(new_n11012_));
  AOI21_X1   g10726(.A1(new_n10989_), .A2(new_n10995_), .B(new_n11001_), .ZN(new_n11013_));
  OAI21_X1   g10727(.A1(new_n10984_), .A2(new_n10988_), .B(new_n10992_), .ZN(new_n11014_));
  AOI21_X1   g10728(.A1(new_n11014_), .A2(new_n11003_), .B(new_n10952_), .ZN(new_n11015_));
  NOR2_X1    g10729(.A1(new_n11015_), .A2(new_n11013_), .ZN(new_n11016_));
  NAND2_X1   g10730(.A1(new_n11016_), .A2(new_n11010_), .ZN(new_n11017_));
  AOI22_X1   g10731(.A1(new_n11017_), .A2(new_n11012_), .B1(new_n10944_), .B2(new_n10942_), .ZN(new_n11018_));
  NAND2_X1   g10732(.A1(new_n10944_), .A2(new_n10942_), .ZN(new_n11019_));
  NOR3_X1    g10733(.A1(new_n11015_), .A2(new_n11013_), .A3(new_n11010_), .ZN(new_n11020_));
  AOI21_X1   g10734(.A1(new_n10997_), .A2(new_n11005_), .B(new_n11011_), .ZN(new_n11021_));
  NOR2_X1    g10735(.A1(new_n11020_), .A2(new_n11021_), .ZN(new_n11022_));
  NOR2_X1    g10736(.A1(new_n11019_), .A2(new_n11022_), .ZN(new_n11023_));
  NOR2_X1    g10737(.A1(new_n11023_), .A2(new_n11018_), .ZN(new_n11024_));
  OAI22_X1   g10738(.A1(new_n7619_), .A2(new_n565_), .B1(new_n656_), .B2(new_n8309_), .ZN(new_n11025_));
  OAI21_X1   g10739(.A1(new_n515_), .A2(new_n7947_), .B(new_n11025_), .ZN(new_n11026_));
  AOI21_X1   g10740(.A1(new_n11026_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n11027_));
  XNOR2_X1   g10741(.A1(new_n660_), .A2(new_n11027_), .ZN(new_n11028_));
  NOR2_X1    g10742(.A1(new_n11024_), .A2(new_n11028_), .ZN(new_n11029_));
  INV_X1     g10743(.I(new_n11029_), .ZN(new_n11030_));
  NAND2_X1   g10744(.A1(new_n11024_), .A2(new_n11028_), .ZN(new_n11031_));
  AOI21_X1   g10745(.A1(new_n11030_), .A2(new_n11031_), .B(new_n10941_), .ZN(new_n11032_));
  NOR2_X1    g10746(.A1(new_n10595_), .A2(new_n10597_), .ZN(new_n11033_));
  NOR2_X1    g10747(.A1(new_n11016_), .A2(new_n11010_), .ZN(new_n11034_));
  NOR2_X1    g10748(.A1(new_n11006_), .A2(new_n11011_), .ZN(new_n11035_));
  OAI22_X1   g10749(.A1(new_n11034_), .A2(new_n11035_), .B1(new_n11033_), .B2(new_n10596_), .ZN(new_n11036_));
  NOR2_X1    g10750(.A1(new_n11033_), .A2(new_n10596_), .ZN(new_n11037_));
  NAND3_X1   g10751(.A1(new_n10997_), .A2(new_n11005_), .A3(new_n11011_), .ZN(new_n11038_));
  OAI21_X1   g10752(.A1(new_n11015_), .A2(new_n11013_), .B(new_n11010_), .ZN(new_n11039_));
  NAND2_X1   g10753(.A1(new_n11039_), .A2(new_n11038_), .ZN(new_n11040_));
  NAND2_X1   g10754(.A1(new_n11037_), .A2(new_n11040_), .ZN(new_n11041_));
  INV_X1     g10755(.I(new_n11028_), .ZN(new_n11042_));
  NAND3_X1   g10756(.A1(new_n11041_), .A2(new_n11036_), .A3(new_n11042_), .ZN(new_n11043_));
  OAI21_X1   g10757(.A1(new_n11023_), .A2(new_n11018_), .B(new_n11028_), .ZN(new_n11044_));
  NAND2_X1   g10758(.A1(new_n11044_), .A2(new_n11043_), .ZN(new_n11045_));
  NAND2_X1   g10759(.A1(new_n10941_), .A2(new_n11045_), .ZN(new_n11046_));
  INV_X1     g10760(.I(new_n11046_), .ZN(new_n11047_));
  NOR2_X1    g10761(.A1(new_n11047_), .A2(new_n11032_), .ZN(new_n11048_));
  OAI22_X1   g10762(.A1(new_n6644_), .A2(new_n780_), .B1(new_n861_), .B2(new_n6647_), .ZN(new_n11049_));
  OAI21_X1   g10763(.A1(new_n706_), .A2(new_n7284_), .B(new_n11049_), .ZN(new_n11050_));
  AOI21_X1   g10764(.A1(new_n11050_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n11051_));
  XNOR2_X1   g10765(.A1(new_n860_), .A2(new_n11051_), .ZN(new_n11052_));
  NOR2_X1    g10766(.A1(new_n11048_), .A2(new_n11052_), .ZN(new_n11053_));
  INV_X1     g10767(.I(new_n11053_), .ZN(new_n11054_));
  NAND2_X1   g10768(.A1(new_n11048_), .A2(new_n11052_), .ZN(new_n11055_));
  NAND2_X1   g10769(.A1(new_n11054_), .A2(new_n11055_), .ZN(new_n11056_));
  INV_X1     g10770(.I(new_n11056_), .ZN(new_n11057_));
  NOR3_X1    g10771(.A1(new_n10939_), .A2(new_n10936_), .A3(new_n11057_), .ZN(new_n11058_));
  NAND2_X1   g10772(.A1(new_n10626_), .A2(new_n10629_), .ZN(new_n11059_));
  NAND2_X1   g10773(.A1(new_n10645_), .A2(new_n11059_), .ZN(new_n11060_));
  NOR2_X1    g10774(.A1(new_n10546_), .A2(new_n10633_), .ZN(new_n11061_));
  OAI21_X1   g10775(.A1(new_n10645_), .A2(new_n11059_), .B(new_n11061_), .ZN(new_n11062_));
  AOI21_X1   g10776(.A1(new_n11062_), .A2(new_n11060_), .B(new_n11056_), .ZN(new_n11063_));
  OAI21_X1   g10777(.A1(new_n11063_), .A2(new_n11058_), .B(new_n10934_), .ZN(new_n11064_));
  NAND3_X1   g10778(.A1(new_n11062_), .A2(new_n11060_), .A3(new_n11056_), .ZN(new_n11065_));
  OAI21_X1   g10779(.A1(new_n10939_), .A2(new_n10936_), .B(new_n11057_), .ZN(new_n11066_));
  NAND3_X1   g10780(.A1(new_n11065_), .A2(new_n11066_), .A3(new_n10933_), .ZN(new_n11067_));
  AOI21_X1   g10781(.A1(new_n11064_), .A2(new_n11067_), .B(new_n10928_), .ZN(new_n11068_));
  AOI21_X1   g10782(.A1(new_n11065_), .A2(new_n11066_), .B(new_n10933_), .ZN(new_n11069_));
  NOR3_X1    g10783(.A1(new_n11063_), .A2(new_n11058_), .A3(new_n10934_), .ZN(new_n11070_));
  NOR3_X1    g10784(.A1(new_n11069_), .A2(new_n11070_), .A3(new_n10927_), .ZN(new_n11071_));
  OAI22_X1   g10785(.A1(new_n5420_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n5107_), .ZN(new_n11072_));
  OAI21_X1   g10786(.A1(new_n1189_), .A2(new_n5112_), .B(new_n11072_), .ZN(new_n11073_));
  AOI21_X1   g10787(.A1(new_n11073_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n11074_));
  XNOR2_X1   g10788(.A1(new_n1421_), .A2(new_n11074_), .ZN(new_n11075_));
  NOR3_X1    g10789(.A1(new_n11071_), .A2(new_n11068_), .A3(new_n11075_), .ZN(new_n11076_));
  OAI21_X1   g10790(.A1(new_n11069_), .A2(new_n11070_), .B(new_n10927_), .ZN(new_n11077_));
  NAND3_X1   g10791(.A1(new_n11064_), .A2(new_n11067_), .A3(new_n10928_), .ZN(new_n11078_));
  INV_X1     g10792(.I(new_n11075_), .ZN(new_n11079_));
  AOI21_X1   g10793(.A1(new_n11077_), .A2(new_n11078_), .B(new_n11079_), .ZN(new_n11080_));
  OAI21_X1   g10794(.A1(new_n11076_), .A2(new_n11080_), .B(new_n10923_), .ZN(new_n11081_));
  NAND2_X1   g10795(.A1(new_n10541_), .A2(new_n10257_), .ZN(new_n11082_));
  AOI21_X1   g10796(.A1(new_n11082_), .A2(new_n10675_), .B(new_n10660_), .ZN(new_n11083_));
  NOR2_X1    g10797(.A1(new_n11071_), .A2(new_n11068_), .ZN(new_n11084_));
  NOR2_X1    g10798(.A1(new_n11084_), .A2(new_n11075_), .ZN(new_n11085_));
  NAND2_X1   g10799(.A1(new_n11077_), .A2(new_n11078_), .ZN(new_n11086_));
  NOR2_X1    g10800(.A1(new_n11086_), .A2(new_n11079_), .ZN(new_n11087_));
  OAI21_X1   g10801(.A1(new_n11085_), .A2(new_n11087_), .B(new_n11083_), .ZN(new_n11088_));
  OAI22_X1   g10802(.A1(new_n4072_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n4067_), .ZN(new_n11089_));
  OAI21_X1   g10803(.A1(new_n1525_), .A2(new_n4318_), .B(new_n11089_), .ZN(new_n11090_));
  AOI21_X1   g10804(.A1(new_n11090_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n11091_));
  XOR2_X1    g10805(.A1(new_n1808_), .A2(new_n11091_), .Z(new_n11092_));
  AOI21_X1   g10806(.A1(new_n11088_), .A2(new_n11081_), .B(new_n11092_), .ZN(new_n11093_));
  NAND3_X1   g10807(.A1(new_n11077_), .A2(new_n11078_), .A3(new_n11079_), .ZN(new_n11094_));
  OAI21_X1   g10808(.A1(new_n11071_), .A2(new_n11068_), .B(new_n11075_), .ZN(new_n11095_));
  AOI21_X1   g10809(.A1(new_n11094_), .A2(new_n11095_), .B(new_n11083_), .ZN(new_n11096_));
  NAND2_X1   g10810(.A1(new_n11086_), .A2(new_n11079_), .ZN(new_n11097_));
  NAND2_X1   g10811(.A1(new_n11084_), .A2(new_n11075_), .ZN(new_n11098_));
  AOI21_X1   g10812(.A1(new_n11098_), .A2(new_n11097_), .B(new_n10923_), .ZN(new_n11099_));
  INV_X1     g10813(.I(new_n11092_), .ZN(new_n11100_));
  NOR3_X1    g10814(.A1(new_n11099_), .A2(new_n11096_), .A3(new_n11100_), .ZN(new_n11101_));
  NOR2_X1    g10815(.A1(new_n11093_), .A2(new_n11101_), .ZN(new_n11102_));
  INV_X1     g10816(.I(new_n11102_), .ZN(new_n11103_));
  NAND4_X1   g10817(.A1(new_n10538_), .A2(new_n10684_), .A3(new_n9888_), .A4(new_n10692_), .ZN(new_n11104_));
  NAND3_X1   g10818(.A1(new_n10534_), .A2(new_n10283_), .A3(new_n10689_), .ZN(new_n11105_));
  INV_X1     g10819(.I(new_n11105_), .ZN(new_n11106_));
  OAI21_X1   g10820(.A1(new_n10694_), .A2(new_n10684_), .B(new_n11106_), .ZN(new_n11107_));
  NAND2_X1   g10821(.A1(new_n10299_), .A2(new_n10300_), .ZN(new_n11108_));
  NOR2_X1    g10822(.A1(new_n10663_), .A2(new_n10658_), .ZN(new_n11109_));
  NAND2_X1   g10823(.A1(new_n10673_), .A2(new_n10677_), .ZN(new_n11110_));
  OAI21_X1   g10824(.A1(new_n11110_), .A2(new_n10279_), .B(new_n10668_), .ZN(new_n11111_));
  OAI22_X1   g10825(.A1(new_n11108_), .A2(new_n11111_), .B1(new_n10287_), .B2(new_n11109_), .ZN(new_n11112_));
  NAND3_X1   g10826(.A1(new_n11107_), .A2(new_n11104_), .A3(new_n11112_), .ZN(new_n11113_));
  AOI21_X1   g10827(.A1(new_n10539_), .A2(new_n10538_), .B(new_n10684_), .ZN(new_n11114_));
  OAI21_X1   g10828(.A1(new_n11114_), .A2(new_n11105_), .B(new_n11104_), .ZN(new_n11115_));
  NOR2_X1    g10829(.A1(new_n10290_), .A2(new_n10671_), .ZN(new_n11116_));
  AOI21_X1   g10830(.A1(new_n11109_), .A2(new_n10287_), .B(new_n10667_), .ZN(new_n11117_));
  AOI22_X1   g10831(.A1(new_n11116_), .A2(new_n11117_), .B1(new_n10279_), .B2(new_n11110_), .ZN(new_n11118_));
  NAND2_X1   g10832(.A1(new_n11115_), .A2(new_n11118_), .ZN(new_n11119_));
  AOI21_X1   g10833(.A1(new_n11119_), .A2(new_n11113_), .B(new_n11103_), .ZN(new_n11120_));
  NOR2_X1    g10834(.A1(new_n11115_), .A2(new_n11118_), .ZN(new_n11121_));
  NAND2_X1   g10835(.A1(new_n9888_), .A2(new_n10692_), .ZN(new_n11122_));
  AOI21_X1   g10836(.A1(new_n10681_), .A2(new_n10682_), .B(new_n10279_), .ZN(new_n11123_));
  NOR3_X1    g10837(.A1(new_n10679_), .A2(new_n10670_), .A3(new_n10287_), .ZN(new_n11124_));
  NOR2_X1    g10838(.A1(new_n11124_), .A2(new_n11123_), .ZN(new_n11125_));
  NOR3_X1    g10839(.A1(new_n11122_), .A2(new_n10691_), .A3(new_n11125_), .ZN(new_n11126_));
  OAI21_X1   g10840(.A1(new_n11122_), .A2(new_n10691_), .B(new_n11125_), .ZN(new_n11127_));
  AOI21_X1   g10841(.A1(new_n11127_), .A2(new_n11106_), .B(new_n11126_), .ZN(new_n11128_));
  NOR2_X1    g10842(.A1(new_n11128_), .A2(new_n11112_), .ZN(new_n11129_));
  NOR3_X1    g10843(.A1(new_n11129_), .A2(new_n11121_), .A3(new_n11102_), .ZN(new_n11130_));
  OAI21_X1   g10844(.A1(new_n11130_), .A2(new_n11120_), .B(new_n10921_), .ZN(new_n11131_));
  INV_X1     g10845(.I(new_n10921_), .ZN(new_n11132_));
  OAI21_X1   g10846(.A1(new_n11129_), .A2(new_n11121_), .B(new_n11102_), .ZN(new_n11133_));
  NAND3_X1   g10847(.A1(new_n11119_), .A2(new_n11113_), .A3(new_n11103_), .ZN(new_n11134_));
  NAND3_X1   g10848(.A1(new_n11133_), .A2(new_n11134_), .A3(new_n11132_), .ZN(new_n11135_));
  OAI22_X1   g10849(.A1(new_n2643_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n2842_), .ZN(new_n11136_));
  OAI21_X1   g10850(.A1(new_n2439_), .A2(new_n2884_), .B(new_n11136_), .ZN(new_n11137_));
  AOI21_X1   g10851(.A1(new_n11137_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n11138_));
  XNOR2_X1   g10852(.A1(new_n2846_), .A2(new_n11138_), .ZN(new_n11139_));
  INV_X1     g10853(.I(new_n11139_), .ZN(new_n11140_));
  NAND3_X1   g10854(.A1(new_n11131_), .A2(new_n11135_), .A3(new_n11140_), .ZN(new_n11141_));
  AOI21_X1   g10855(.A1(new_n11133_), .A2(new_n11134_), .B(new_n11132_), .ZN(new_n11142_));
  NOR3_X1    g10856(.A1(new_n11130_), .A2(new_n11120_), .A3(new_n10921_), .ZN(new_n11143_));
  OAI21_X1   g10857(.A1(new_n11142_), .A2(new_n11143_), .B(new_n11139_), .ZN(new_n11144_));
  NAND2_X1   g10858(.A1(new_n11144_), .A2(new_n11141_), .ZN(new_n11145_));
  OAI21_X1   g10859(.A1(new_n10699_), .A2(new_n10697_), .B(new_n10712_), .ZN(new_n11146_));
  NAND3_X1   g10860(.A1(new_n10708_), .A2(new_n10531_), .A3(new_n10698_), .ZN(new_n11147_));
  NAND4_X1   g10861(.A1(new_n10533_), .A2(new_n11147_), .A3(new_n10329_), .A4(new_n10704_), .ZN(new_n11148_));
  NAND2_X1   g10862(.A1(new_n11148_), .A2(new_n11146_), .ZN(new_n11149_));
  OAI22_X1   g10863(.A1(new_n2171_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n2166_), .ZN(new_n11150_));
  OAI21_X1   g10864(.A1(new_n3018_), .A2(new_n2322_), .B(new_n11150_), .ZN(new_n11151_));
  AOI21_X1   g10865(.A1(new_n11151_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n11152_));
  XNOR2_X1   g10866(.A1(new_n3514_), .A2(new_n11152_), .ZN(new_n11153_));
  INV_X1     g10867(.I(new_n11153_), .ZN(new_n11154_));
  NAND2_X1   g10868(.A1(new_n11149_), .A2(new_n11154_), .ZN(new_n11155_));
  INV_X1     g10869(.I(new_n11155_), .ZN(new_n11156_));
  NOR2_X1    g10870(.A1(new_n11149_), .A2(new_n11154_), .ZN(new_n11157_));
  OAI21_X1   g10871(.A1(new_n11156_), .A2(new_n11157_), .B(new_n11145_), .ZN(new_n11158_));
  NOR3_X1    g10872(.A1(new_n11142_), .A2(new_n11143_), .A3(new_n11139_), .ZN(new_n11159_));
  AOI21_X1   g10873(.A1(new_n11131_), .A2(new_n11135_), .B(new_n11140_), .ZN(new_n11160_));
  NOR2_X1    g10874(.A1(new_n11159_), .A2(new_n11160_), .ZN(new_n11161_));
  NOR2_X1    g10875(.A1(new_n11149_), .A2(new_n11153_), .ZN(new_n11162_));
  INV_X1     g10876(.I(new_n11149_), .ZN(new_n11163_));
  NOR2_X1    g10877(.A1(new_n11163_), .A2(new_n11154_), .ZN(new_n11164_));
  OAI21_X1   g10878(.A1(new_n11164_), .A2(new_n11162_), .B(new_n11161_), .ZN(new_n11165_));
  NAND2_X1   g10879(.A1(new_n11165_), .A2(new_n11158_), .ZN(new_n11166_));
  OAI22_X1   g10880(.A1(new_n1712_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n1707_), .ZN(new_n11167_));
  OAI21_X1   g10881(.A1(new_n3717_), .A2(new_n1850_), .B(new_n11167_), .ZN(new_n11168_));
  AOI21_X1   g10882(.A1(new_n11168_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n11169_));
  XNOR2_X1   g10883(.A1(new_n4257_), .A2(new_n11169_), .ZN(new_n11170_));
  INV_X1     g10884(.I(new_n11170_), .ZN(new_n11171_));
  NAND2_X1   g10885(.A1(new_n11166_), .A2(new_n11171_), .ZN(new_n11172_));
  INV_X1     g10886(.I(new_n11172_), .ZN(new_n11173_));
  NOR2_X1    g10887(.A1(new_n11166_), .A2(new_n11171_), .ZN(new_n11174_));
  OAI21_X1   g10888(.A1(new_n11173_), .A2(new_n11174_), .B(new_n10917_), .ZN(new_n11175_));
  AND2_X2    g10889(.A1(new_n10915_), .A2(new_n10728_), .Z(new_n11176_));
  AOI22_X1   g10890(.A1(new_n11176_), .A2(new_n10914_), .B1(new_n10526_), .B2(new_n10912_), .ZN(new_n11177_));
  NOR2_X1    g10891(.A1(new_n11166_), .A2(new_n11170_), .ZN(new_n11178_));
  AOI21_X1   g10892(.A1(new_n11165_), .A2(new_n11158_), .B(new_n11171_), .ZN(new_n11179_));
  OAI21_X1   g10893(.A1(new_n11178_), .A2(new_n11179_), .B(new_n11177_), .ZN(new_n11180_));
  OAI22_X1   g10894(.A1(new_n1347_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n1344_), .ZN(new_n11181_));
  OAI21_X1   g10895(.A1(new_n4500_), .A2(new_n1457_), .B(new_n11181_), .ZN(new_n11182_));
  AOI21_X1   g10896(.A1(new_n11182_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n11183_));
  XOR2_X1    g10897(.A1(new_n5067_), .A2(new_n11183_), .Z(new_n11184_));
  AOI21_X1   g10898(.A1(new_n11175_), .A2(new_n11180_), .B(new_n11184_), .ZN(new_n11185_));
  INV_X1     g10899(.I(new_n11174_), .ZN(new_n11186_));
  AOI21_X1   g10900(.A1(new_n11186_), .A2(new_n11172_), .B(new_n11177_), .ZN(new_n11187_));
  INV_X1     g10901(.I(new_n11180_), .ZN(new_n11188_));
  INV_X1     g10902(.I(new_n11184_), .ZN(new_n11189_));
  NOR3_X1    g10903(.A1(new_n11187_), .A2(new_n11188_), .A3(new_n11189_), .ZN(new_n11190_));
  OAI21_X1   g10904(.A1(new_n11190_), .A2(new_n11185_), .B(new_n10911_), .ZN(new_n11191_));
  NOR2_X1    g10905(.A1(new_n10908_), .A2(new_n10522_), .ZN(new_n11192_));
  NOR2_X1    g10906(.A1(new_n10910_), .A2(new_n10743_), .ZN(new_n11193_));
  NOR2_X1    g10907(.A1(new_n11193_), .A2(new_n11192_), .ZN(new_n11194_));
  NAND2_X1   g10908(.A1(new_n11175_), .A2(new_n11180_), .ZN(new_n11195_));
  NOR2_X1    g10909(.A1(new_n11195_), .A2(new_n11184_), .ZN(new_n11196_));
  AOI21_X1   g10910(.A1(new_n11175_), .A2(new_n11180_), .B(new_n11189_), .ZN(new_n11197_));
  OAI21_X1   g10911(.A1(new_n11196_), .A2(new_n11197_), .B(new_n11194_), .ZN(new_n11198_));
  NAND2_X1   g10912(.A1(new_n11198_), .A2(new_n11191_), .ZN(new_n11199_));
  OAI22_X1   g10913(.A1(new_n1055_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n1061_), .ZN(new_n11200_));
  OAI21_X1   g10914(.A1(new_n5353_), .A2(new_n1332_), .B(new_n11200_), .ZN(new_n11201_));
  AOI21_X1   g10915(.A1(new_n11201_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n11202_));
  XOR2_X1    g10916(.A1(new_n5926_), .A2(new_n11202_), .Z(new_n11203_));
  INV_X1     g10917(.I(new_n11203_), .ZN(new_n11204_));
  XOR2_X1    g10918(.A1(new_n11199_), .A2(new_n11204_), .Z(new_n11205_));
  NOR2_X1    g10919(.A1(new_n11199_), .A2(new_n11203_), .ZN(new_n11206_));
  INV_X1     g10920(.I(new_n11191_), .ZN(new_n11207_));
  NOR2_X1    g10921(.A1(new_n11187_), .A2(new_n11188_), .ZN(new_n11208_));
  NAND2_X1   g10922(.A1(new_n11208_), .A2(new_n11189_), .ZN(new_n11209_));
  INV_X1     g10923(.I(new_n11197_), .ZN(new_n11210_));
  AOI21_X1   g10924(.A1(new_n11209_), .A2(new_n11210_), .B(new_n10911_), .ZN(new_n11211_));
  NOR2_X1    g10925(.A1(new_n11211_), .A2(new_n11207_), .ZN(new_n11212_));
  NOR2_X1    g10926(.A1(new_n11212_), .A2(new_n11204_), .ZN(new_n11213_));
  OAI21_X1   g10927(.A1(new_n11213_), .A2(new_n11206_), .B(new_n10907_), .ZN(new_n11214_));
  OAI21_X1   g10928(.A1(new_n10907_), .A2(new_n11205_), .B(new_n11214_), .ZN(new_n11215_));
  NAND3_X1   g10929(.A1(new_n11215_), .A2(new_n10903_), .A3(new_n10901_), .ZN(new_n11216_));
  NAND2_X1   g10930(.A1(new_n10903_), .A2(new_n10901_), .ZN(new_n11217_));
  NOR2_X1    g10931(.A1(new_n11205_), .A2(new_n10907_), .ZN(new_n11218_));
  NAND3_X1   g10932(.A1(new_n10748_), .A2(new_n10752_), .A3(new_n10390_), .ZN(new_n11219_));
  NAND2_X1   g10933(.A1(new_n11219_), .A2(new_n10763_), .ZN(new_n11220_));
  OAI22_X1   g10934(.A1(new_n11220_), .A2(new_n10521_), .B1(new_n10390_), .B2(new_n10904_), .ZN(new_n11221_));
  NOR2_X1    g10935(.A1(new_n11213_), .A2(new_n11206_), .ZN(new_n11222_));
  NOR2_X1    g10936(.A1(new_n11222_), .A2(new_n11221_), .ZN(new_n11223_));
  NOR2_X1    g10937(.A1(new_n11218_), .A2(new_n11223_), .ZN(new_n11224_));
  NAND2_X1   g10938(.A1(new_n11224_), .A2(new_n11217_), .ZN(new_n11225_));
  OAI22_X1   g10939(.A1(new_n970_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n820_), .ZN(new_n11226_));
  OAI21_X1   g10940(.A1(new_n6229_), .A2(new_n894_), .B(new_n11226_), .ZN(new_n11227_));
  AOI21_X1   g10941(.A1(new_n11227_), .A2(new_n827_), .B(new_n970_), .ZN(new_n11228_));
  XOR2_X1    g10942(.A1(new_n6851_), .A2(new_n11228_), .Z(new_n11229_));
  INV_X1     g10943(.I(new_n11229_), .ZN(new_n11230_));
  NAND3_X1   g10944(.A1(new_n11225_), .A2(new_n11216_), .A3(new_n11230_), .ZN(new_n11231_));
  INV_X1     g10945(.I(new_n11216_), .ZN(new_n11232_));
  AOI21_X1   g10946(.A1(new_n10901_), .A2(new_n10903_), .B(new_n11215_), .ZN(new_n11233_));
  OAI21_X1   g10947(.A1(new_n11232_), .A2(new_n11233_), .B(new_n11229_), .ZN(new_n11234_));
  AOI22_X1   g10948(.A1(new_n10899_), .A2(new_n10897_), .B1(new_n11234_), .B2(new_n11231_), .ZN(new_n11235_));
  NOR2_X1    g10949(.A1(new_n10801_), .A2(new_n10426_), .ZN(new_n11236_));
  NOR3_X1    g10950(.A1(new_n10799_), .A2(new_n10800_), .A3(new_n10419_), .ZN(new_n11237_));
  NOR3_X1    g10951(.A1(new_n10517_), .A2(new_n11237_), .A3(new_n10791_), .ZN(new_n11238_));
  AOI21_X1   g10952(.A1(new_n11225_), .A2(new_n11216_), .B(new_n11229_), .ZN(new_n11239_));
  NOR3_X1    g10953(.A1(new_n11232_), .A2(new_n11233_), .A3(new_n11230_), .ZN(new_n11240_));
  NOR2_X1    g10954(.A1(new_n11240_), .A2(new_n11239_), .ZN(new_n11241_));
  NOR3_X1    g10955(.A1(new_n11241_), .A2(new_n11236_), .A3(new_n11238_), .ZN(new_n11242_));
  OAI22_X1   g10956(.A1(new_n607_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n610_), .ZN(new_n11243_));
  OAI21_X1   g10957(.A1(new_n7198_), .A2(new_n684_), .B(new_n11243_), .ZN(new_n11244_));
  AOI21_X1   g10958(.A1(new_n11244_), .A2(new_n612_), .B(new_n607_), .ZN(new_n11245_));
  XNOR2_X1   g10959(.A1(new_n7874_), .A2(new_n11245_), .ZN(new_n11246_));
  NOR3_X1    g10960(.A1(new_n11242_), .A2(new_n11235_), .A3(new_n11246_), .ZN(new_n11247_));
  INV_X1     g10961(.I(new_n11247_), .ZN(new_n11248_));
  OAI21_X1   g10962(.A1(new_n11242_), .A2(new_n11235_), .B(new_n11246_), .ZN(new_n11249_));
  AOI22_X1   g10963(.A1(new_n10896_), .A2(new_n10894_), .B1(new_n11248_), .B2(new_n11249_), .ZN(new_n11250_));
  NAND2_X1   g10964(.A1(new_n10896_), .A2(new_n10894_), .ZN(new_n11251_));
  INV_X1     g10965(.I(new_n11246_), .ZN(new_n11252_));
  OAI21_X1   g10966(.A1(new_n11242_), .A2(new_n11235_), .B(new_n11252_), .ZN(new_n11253_));
  INV_X1     g10967(.I(new_n11253_), .ZN(new_n11254_));
  NOR3_X1    g10968(.A1(new_n11242_), .A2(new_n11235_), .A3(new_n11252_), .ZN(new_n11255_));
  NOR2_X1    g10969(.A1(new_n11254_), .A2(new_n11255_), .ZN(new_n11256_));
  NOR2_X1    g10970(.A1(new_n11251_), .A2(new_n11256_), .ZN(new_n11257_));
  OAI22_X1   g10971(.A1(new_n448_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n450_), .ZN(new_n11258_));
  OAI21_X1   g10972(.A1(new_n8218_), .A2(new_n496_), .B(new_n11258_), .ZN(new_n11259_));
  AOI21_X1   g10973(.A1(new_n11259_), .A2(new_n452_), .B(new_n448_), .ZN(new_n11260_));
  XOR2_X1    g10974(.A1(new_n8952_), .A2(new_n11260_), .Z(new_n11261_));
  INV_X1     g10975(.I(new_n11261_), .ZN(new_n11262_));
  OAI21_X1   g10976(.A1(new_n11257_), .A2(new_n11250_), .B(new_n11262_), .ZN(new_n11263_));
  NAND2_X1   g10977(.A1(new_n10895_), .A2(new_n10814_), .ZN(new_n11264_));
  NOR3_X1    g10978(.A1(new_n11264_), .A2(new_n10513_), .A3(new_n10515_), .ZN(new_n11265_));
  NAND2_X1   g10979(.A1(new_n11248_), .A2(new_n11249_), .ZN(new_n11266_));
  OAI21_X1   g10980(.A1(new_n11265_), .A2(new_n10893_), .B(new_n11266_), .ZN(new_n11267_));
  INV_X1     g10981(.I(new_n11255_), .ZN(new_n11268_));
  NAND2_X1   g10982(.A1(new_n11268_), .A2(new_n11253_), .ZN(new_n11269_));
  NAND3_X1   g10983(.A1(new_n11269_), .A2(new_n10896_), .A3(new_n10894_), .ZN(new_n11270_));
  NAND3_X1   g10984(.A1(new_n11267_), .A2(new_n11270_), .A3(new_n11261_), .ZN(new_n11271_));
  OAI22_X1   g10985(.A1(new_n10025_), .A2(new_n341_), .B1(new_n404_), .B2(new_n10031_), .ZN(new_n11272_));
  OAI21_X1   g10986(.A1(new_n9295_), .A2(new_n366_), .B(new_n11272_), .ZN(new_n11273_));
  AOI21_X1   g10987(.A1(new_n11273_), .A2(new_n334_), .B(new_n341_), .ZN(new_n11274_));
  XNOR2_X1   g10988(.A1(new_n10035_), .A2(new_n11274_), .ZN(new_n11275_));
  INV_X1     g10989(.I(new_n11275_), .ZN(new_n11276_));
  NAND3_X1   g10990(.A1(new_n11263_), .A2(new_n11271_), .A3(new_n11276_), .ZN(new_n11277_));
  INV_X1     g10991(.I(new_n11277_), .ZN(new_n11278_));
  AOI21_X1   g10992(.A1(new_n11263_), .A2(new_n11271_), .B(new_n11276_), .ZN(new_n11279_));
  OAI22_X1   g10993(.A1(new_n10892_), .A2(new_n10890_), .B1(new_n11278_), .B2(new_n11279_), .ZN(new_n11280_));
  INV_X1     g10994(.I(new_n10890_), .ZN(new_n11281_));
  AOI21_X1   g10995(.A1(new_n10822_), .A2(new_n10842_), .B(new_n10826_), .ZN(new_n11282_));
  NAND3_X1   g10996(.A1(new_n10832_), .A2(new_n10830_), .A3(new_n11282_), .ZN(new_n11283_));
  AOI21_X1   g10997(.A1(new_n11267_), .A2(new_n11270_), .B(new_n11261_), .ZN(new_n11284_));
  NOR3_X1    g10998(.A1(new_n11257_), .A2(new_n11250_), .A3(new_n11262_), .ZN(new_n11285_));
  OAI21_X1   g10999(.A1(new_n11285_), .A2(new_n11284_), .B(new_n11276_), .ZN(new_n11286_));
  NAND3_X1   g11000(.A1(new_n11263_), .A2(new_n11271_), .A3(new_n11275_), .ZN(new_n11287_));
  NAND2_X1   g11001(.A1(new_n11286_), .A2(new_n11287_), .ZN(new_n11288_));
  NAND3_X1   g11002(.A1(new_n11288_), .A2(new_n11283_), .A3(new_n11281_), .ZN(new_n11289_));
  NAND2_X1   g11003(.A1(new_n11280_), .A2(new_n11289_), .ZN(new_n11290_));
  NAND2_X1   g11004(.A1(new_n10846_), .A2(new_n10494_), .ZN(new_n11291_));
  OAI21_X1   g11005(.A1(new_n10839_), .A2(new_n10845_), .B(new_n10493_), .ZN(new_n11292_));
  NAND2_X1   g11006(.A1(new_n10854_), .A2(new_n11292_), .ZN(new_n11293_));
  XNOR2_X1   g11007(.A1(\b[53] ), .A2(\b[55] ), .ZN(new_n11294_));
  NOR4_X1    g11008(.A1(new_n10856_), .A2(new_n10859_), .A3(new_n10861_), .A4(new_n11294_), .ZN(new_n11295_));
  NOR2_X1    g11009(.A1(new_n11294_), .A2(new_n10861_), .ZN(new_n11296_));
  NOR2_X1    g11010(.A1(new_n10860_), .A2(new_n11296_), .ZN(new_n11297_));
  NOR2_X1    g11011(.A1(new_n11297_), .A2(new_n11295_), .ZN(new_n11298_));
  INV_X1     g11012(.I(new_n11298_), .ZN(new_n11299_));
  NOR2_X1    g11013(.A1(new_n330_), .A2(new_n10862_), .ZN(new_n11300_));
  INV_X1     g11014(.I(new_n11300_), .ZN(new_n11301_));
  AOI22_X1   g11015(.A1(new_n304_), .A2(\b[53] ), .B1(new_n262_), .B2(\b[55] ), .ZN(new_n11302_));
  AOI21_X1   g11016(.A1(new_n11301_), .A2(new_n11302_), .B(new_n426_), .ZN(new_n11303_));
  NAND2_X1   g11017(.A1(new_n11299_), .A2(new_n11303_), .ZN(new_n11304_));
  INV_X1     g11018(.I(new_n11304_), .ZN(new_n11305_));
  NAND3_X1   g11019(.A1(new_n11293_), .A2(new_n11291_), .A3(new_n11305_), .ZN(new_n11306_));
  NOR2_X1    g11020(.A1(new_n10880_), .A2(new_n10493_), .ZN(new_n11307_));
  AOI22_X1   g11021(.A1(new_n10874_), .A2(new_n10849_), .B1(new_n10880_), .B2(new_n10493_), .ZN(new_n11308_));
  OAI21_X1   g11022(.A1(new_n11308_), .A2(new_n11307_), .B(new_n11304_), .ZN(new_n11309_));
  AOI21_X1   g11023(.A1(new_n11309_), .A2(new_n11306_), .B(new_n11290_), .ZN(new_n11310_));
  INV_X1     g11024(.I(new_n11279_), .ZN(new_n11311_));
  AOI22_X1   g11025(.A1(new_n11283_), .A2(new_n11281_), .B1(new_n11311_), .B2(new_n11277_), .ZN(new_n11312_));
  AOI21_X1   g11026(.A1(new_n11263_), .A2(new_n11271_), .B(new_n11275_), .ZN(new_n11313_));
  NOR3_X1    g11027(.A1(new_n11285_), .A2(new_n11284_), .A3(new_n11276_), .ZN(new_n11314_));
  NOR2_X1    g11028(.A1(new_n11314_), .A2(new_n11313_), .ZN(new_n11315_));
  NOR3_X1    g11029(.A1(new_n11315_), .A2(new_n10892_), .A3(new_n10890_), .ZN(new_n11316_));
  NOR2_X1    g11030(.A1(new_n11312_), .A2(new_n11316_), .ZN(new_n11317_));
  NOR3_X1    g11031(.A1(new_n11308_), .A2(new_n11307_), .A3(new_n11304_), .ZN(new_n11318_));
  AOI21_X1   g11032(.A1(new_n11293_), .A2(new_n11291_), .B(new_n11305_), .ZN(new_n11319_));
  NOR3_X1    g11033(.A1(new_n11318_), .A2(new_n11319_), .A3(new_n11317_), .ZN(new_n11320_));
  OAI21_X1   g11034(.A1(new_n11320_), .A2(new_n11310_), .B(new_n260_), .ZN(new_n11321_));
  OAI21_X1   g11035(.A1(new_n11318_), .A2(new_n11319_), .B(new_n11317_), .ZN(new_n11322_));
  NAND3_X1   g11036(.A1(new_n11309_), .A2(new_n11306_), .A3(new_n11290_), .ZN(new_n11323_));
  NAND3_X1   g11037(.A1(new_n11322_), .A2(new_n11323_), .A3(\a[2] ), .ZN(new_n11324_));
  NAND2_X1   g11038(.A1(new_n11321_), .A2(new_n11324_), .ZN(new_n11325_));
  AOI21_X1   g11039(.A1(new_n10882_), .A2(new_n10881_), .B(new_n10880_), .ZN(new_n11326_));
  NOR3_X1    g11040(.A1(new_n10871_), .A2(new_n10876_), .A3(new_n10846_), .ZN(new_n11327_));
  NOR3_X1    g11041(.A1(new_n11327_), .A2(new_n11326_), .A3(new_n10493_), .ZN(new_n11328_));
  OAI21_X1   g11042(.A1(new_n11328_), .A2(new_n10884_), .B(new_n10482_), .ZN(new_n11329_));
  NAND2_X1   g11043(.A1(new_n11329_), .A2(new_n10473_), .ZN(new_n11330_));
  NAND3_X1   g11044(.A1(new_n10885_), .A2(new_n10886_), .A3(new_n10481_), .ZN(new_n11331_));
  NAND3_X1   g11045(.A1(new_n11330_), .A2(new_n10060_), .A3(new_n11331_), .ZN(new_n11332_));
  INV_X1     g11046(.I(new_n11332_), .ZN(new_n11333_));
  XOR2_X1    g11047(.A1(new_n10880_), .A2(new_n10493_), .Z(new_n11334_));
  NAND2_X1   g11048(.A1(new_n11334_), .A2(new_n10854_), .ZN(new_n11335_));
  INV_X1     g11049(.I(new_n10854_), .ZN(new_n11336_));
  NAND2_X1   g11050(.A1(new_n11291_), .A2(new_n11292_), .ZN(new_n11337_));
  NAND2_X1   g11051(.A1(new_n11337_), .A2(new_n11336_), .ZN(new_n11338_));
  AOI21_X1   g11052(.A1(new_n11335_), .A2(new_n11338_), .B(new_n10875_), .ZN(new_n11339_));
  NOR2_X1    g11053(.A1(new_n11333_), .A2(new_n11339_), .ZN(new_n11340_));
  INV_X1     g11054(.I(new_n11339_), .ZN(new_n11341_));
  NAND2_X1   g11055(.A1(new_n11325_), .A2(new_n11341_), .ZN(new_n11342_));
  OAI22_X1   g11056(.A1(new_n11340_), .A2(new_n11325_), .B1(new_n11333_), .B2(new_n11342_), .ZN(\f[55] ));
  XOR2_X1    g11057(.A1(new_n11290_), .A2(new_n260_), .Z(new_n11344_));
  AOI21_X1   g11058(.A1(new_n11309_), .A2(new_n11306_), .B(new_n11344_), .ZN(new_n11345_));
  AOI21_X1   g11059(.A1(new_n11325_), .A2(new_n11345_), .B(new_n11339_), .ZN(new_n11346_));
  NOR2_X1    g11060(.A1(new_n11346_), .A2(new_n11332_), .ZN(new_n11347_));
  OAI22_X1   g11061(.A1(new_n10892_), .A2(new_n10890_), .B1(new_n11284_), .B2(new_n11285_), .ZN(new_n11348_));
  NOR2_X1    g11062(.A1(new_n10892_), .A2(new_n10890_), .ZN(new_n11349_));
  NAND3_X1   g11063(.A1(new_n11349_), .A2(new_n11263_), .A3(new_n11271_), .ZN(new_n11350_));
  AOI21_X1   g11064(.A1(new_n11350_), .A2(new_n11348_), .B(new_n11276_), .ZN(new_n11351_));
  INV_X1     g11065(.I(new_n11351_), .ZN(new_n11352_));
  AOI21_X1   g11066(.A1(new_n11290_), .A2(new_n10880_), .B(new_n10494_), .ZN(new_n11353_));
  NOR2_X1    g11067(.A1(new_n11290_), .A2(new_n10880_), .ZN(new_n11354_));
  NOR3_X1    g11068(.A1(new_n11336_), .A2(new_n11353_), .A3(new_n11354_), .ZN(new_n11355_));
  NAND2_X1   g11069(.A1(new_n11283_), .A2(new_n11281_), .ZN(new_n11356_));
  INV_X1     g11070(.I(new_n11251_), .ZN(new_n11357_));
  OAI22_X1   g11071(.A1(new_n970_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n820_), .ZN(new_n11358_));
  OAI21_X1   g11072(.A1(new_n6538_), .A2(new_n894_), .B(new_n11358_), .ZN(new_n11359_));
  AOI21_X1   g11073(.A1(new_n11359_), .A2(new_n827_), .B(new_n970_), .ZN(new_n11360_));
  XNOR2_X1   g11074(.A1(new_n7202_), .A2(new_n11360_), .ZN(new_n11361_));
  INV_X1     g11075(.I(new_n11361_), .ZN(new_n11362_));
  INV_X1     g11076(.I(new_n11217_), .ZN(new_n11363_));
  XOR2_X1    g11077(.A1(new_n11221_), .A2(new_n11199_), .Z(new_n11364_));
  NAND2_X1   g11078(.A1(new_n11364_), .A2(new_n11203_), .ZN(new_n11365_));
  NOR2_X1    g11079(.A1(new_n11208_), .A2(new_n10911_), .ZN(new_n11366_));
  NOR2_X1    g11080(.A1(new_n11194_), .A2(new_n11195_), .ZN(new_n11367_));
  OAI21_X1   g11081(.A1(new_n11367_), .A2(new_n11366_), .B(new_n11184_), .ZN(new_n11368_));
  AND2_X2    g11082(.A1(new_n11165_), .A2(new_n11158_), .Z(new_n11369_));
  NOR2_X1    g11083(.A1(new_n11369_), .A2(new_n10917_), .ZN(new_n11370_));
  NOR2_X1    g11084(.A1(new_n11177_), .A2(new_n11166_), .ZN(new_n11371_));
  OAI21_X1   g11085(.A1(new_n11370_), .A2(new_n11371_), .B(new_n11170_), .ZN(new_n11372_));
  NOR2_X1    g11086(.A1(new_n11145_), .A2(new_n11163_), .ZN(new_n11373_));
  NOR2_X1    g11087(.A1(new_n11161_), .A2(new_n11149_), .ZN(new_n11374_));
  OAI21_X1   g11088(.A1(new_n11373_), .A2(new_n11374_), .B(new_n11153_), .ZN(new_n11375_));
  OAI22_X1   g11089(.A1(new_n2281_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n2439_), .ZN(new_n11376_));
  OAI21_X1   g11090(.A1(new_n2102_), .A2(new_n3569_), .B(new_n11376_), .ZN(new_n11377_));
  AOI21_X1   g11091(.A1(new_n11377_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n11378_));
  XNOR2_X1   g11092(.A1(new_n2443_), .A2(new_n11378_), .ZN(new_n11379_));
  INV_X1     g11093(.I(new_n11379_), .ZN(new_n11380_));
  NAND3_X1   g11094(.A1(new_n11088_), .A2(new_n11081_), .A3(new_n11092_), .ZN(new_n11381_));
  AOI21_X1   g11095(.A1(new_n11112_), .A2(new_n11381_), .B(new_n11093_), .ZN(new_n11382_));
  AOI21_X1   g11096(.A1(new_n10923_), .A2(new_n11095_), .B(new_n11076_), .ZN(new_n11383_));
  OAI21_X1   g11097(.A1(new_n10939_), .A2(new_n10936_), .B(new_n10928_), .ZN(new_n11384_));
  NOR3_X1    g11098(.A1(new_n10939_), .A2(new_n10936_), .A3(new_n10928_), .ZN(new_n11385_));
  XOR2_X1    g11099(.A1(new_n11056_), .A2(new_n10933_), .Z(new_n11386_));
  INV_X1     g11100(.I(new_n11386_), .ZN(new_n11387_));
  OAI21_X1   g11101(.A1(new_n11387_), .A2(new_n11385_), .B(new_n11384_), .ZN(new_n11388_));
  OAI21_X1   g11102(.A1(new_n10998_), .A2(new_n11000_), .B(new_n11014_), .ZN(new_n11389_));
  AOI21_X1   g11103(.A1(new_n10986_), .A2(new_n10985_), .B(new_n10999_), .ZN(new_n11390_));
  XNOR2_X1   g11104(.A1(\a[53] ), .A2(\a[55] ), .ZN(new_n11391_));
  XNOR2_X1   g11105(.A1(\a[53] ), .A2(\a[56] ), .ZN(new_n11392_));
  XNOR2_X1   g11106(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n11393_));
  NOR3_X1    g11107(.A1(new_n11391_), .A2(new_n11392_), .A3(new_n11393_), .ZN(new_n11394_));
  AOI22_X1   g11108(.A1(new_n10969_), .A2(new_n10131_), .B1(new_n11394_), .B2(\b[0] ), .ZN(new_n11395_));
  NOR2_X1    g11109(.A1(new_n11395_), .A2(\a[56] ), .ZN(new_n11396_));
  NOR3_X1    g11110(.A1(new_n11396_), .A2(new_n490_), .A3(new_n10975_), .ZN(new_n11397_));
  XOR2_X1    g11111(.A1(\a[53] ), .A2(\a[55] ), .Z(new_n11398_));
  XOR2_X1    g11112(.A1(\a[53] ), .A2(\a[56] ), .Z(new_n11399_));
  XOR2_X1    g11113(.A1(\a[53] ), .A2(\a[54] ), .Z(new_n11400_));
  NAND3_X1   g11114(.A1(new_n11398_), .A2(new_n11399_), .A3(new_n11400_), .ZN(new_n11401_));
  OAI22_X1   g11115(.A1(new_n10979_), .A2(new_n10132_), .B1(new_n258_), .B2(new_n11401_), .ZN(new_n11402_));
  NAND2_X1   g11116(.A1(new_n11402_), .A2(new_n10973_), .ZN(new_n11403_));
  AOI21_X1   g11117(.A1(new_n11403_), .A2(new_n282_), .B(new_n10964_), .ZN(new_n11404_));
  OAI21_X1   g11118(.A1(new_n11397_), .A2(new_n11404_), .B(new_n11390_), .ZN(new_n11405_));
  OAI21_X1   g11119(.A1(new_n10982_), .A2(new_n10972_), .B(new_n10950_), .ZN(new_n11406_));
  NAND3_X1   g11120(.A1(new_n11403_), .A2(new_n282_), .A3(new_n10964_), .ZN(new_n11407_));
  OAI21_X1   g11121(.A1(new_n11396_), .A2(new_n490_), .B(new_n10975_), .ZN(new_n11408_));
  NAND3_X1   g11122(.A1(new_n11406_), .A2(new_n11407_), .A3(new_n11408_), .ZN(new_n11409_));
  INV_X1     g11123(.I(new_n413_), .ZN(new_n11410_));
  NOR2_X1    g11124(.A1(new_n10126_), .A2(new_n10124_), .ZN(new_n11411_));
  OAI22_X1   g11125(.A1(new_n11411_), .A2(new_n11410_), .B1(new_n298_), .B2(new_n10137_), .ZN(new_n11412_));
  NAND2_X1   g11126(.A1(new_n11412_), .A2(new_n9718_), .ZN(new_n11413_));
  NAND3_X1   g11127(.A1(new_n11413_), .A2(new_n2333_), .A3(new_n9712_), .ZN(new_n11414_));
  NAND2_X1   g11128(.A1(new_n9717_), .A2(new_n9715_), .ZN(new_n11415_));
  NAND2_X1   g11129(.A1(new_n11415_), .A2(new_n413_), .ZN(new_n11416_));
  NAND2_X1   g11130(.A1(new_n10145_), .A2(\b[3] ), .ZN(new_n11417_));
  AOI21_X1   g11131(.A1(new_n11416_), .A2(new_n11417_), .B(\a[53] ), .ZN(new_n11418_));
  OAI21_X1   g11132(.A1(new_n11418_), .A2(new_n9713_), .B(new_n378_), .ZN(new_n11419_));
  NAND2_X1   g11133(.A1(new_n11414_), .A2(new_n11419_), .ZN(new_n11420_));
  NAND3_X1   g11134(.A1(new_n11405_), .A2(new_n11409_), .A3(new_n11420_), .ZN(new_n11421_));
  AOI21_X1   g11135(.A1(new_n11405_), .A2(new_n11409_), .B(new_n11420_), .ZN(new_n11422_));
  INV_X1     g11136(.I(new_n11422_), .ZN(new_n11423_));
  AOI22_X1   g11137(.A1(new_n11389_), .A2(new_n11003_), .B1(new_n11423_), .B2(new_n11421_), .ZN(new_n11424_));
  OAI21_X1   g11138(.A1(new_n11001_), .A2(new_n11002_), .B(new_n11003_), .ZN(new_n11425_));
  NOR3_X1    g11139(.A1(new_n11418_), .A2(new_n378_), .A3(new_n9713_), .ZN(new_n11426_));
  AOI21_X1   g11140(.A1(new_n11413_), .A2(new_n9712_), .B(new_n2333_), .ZN(new_n11427_));
  NOR2_X1    g11141(.A1(new_n11427_), .A2(new_n11426_), .ZN(new_n11428_));
  AOI21_X1   g11142(.A1(new_n11405_), .A2(new_n11409_), .B(new_n11428_), .ZN(new_n11429_));
  AOI21_X1   g11143(.A1(new_n11407_), .A2(new_n11408_), .B(new_n11406_), .ZN(new_n11430_));
  NOR3_X1    g11144(.A1(new_n11390_), .A2(new_n11404_), .A3(new_n11397_), .ZN(new_n11431_));
  NOR3_X1    g11145(.A1(new_n11430_), .A2(new_n11431_), .A3(new_n11420_), .ZN(new_n11432_));
  NOR2_X1    g11146(.A1(new_n11432_), .A2(new_n11429_), .ZN(new_n11433_));
  NOR2_X1    g11147(.A1(new_n11425_), .A2(new_n11433_), .ZN(new_n11434_));
  OAI22_X1   g11148(.A1(new_n8644_), .A2(new_n472_), .B1(new_n515_), .B2(new_n9388_), .ZN(new_n11435_));
  OAI21_X1   g11149(.A1(new_n420_), .A2(new_n10154_), .B(new_n11435_), .ZN(new_n11436_));
  AOI21_X1   g11150(.A1(new_n11436_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n11437_));
  XOR2_X1    g11151(.A1(new_n700_), .A2(new_n11437_), .Z(new_n11438_));
  NOR3_X1    g11152(.A1(new_n11434_), .A2(new_n11424_), .A3(new_n11438_), .ZN(new_n11439_));
  AOI21_X1   g11153(.A1(new_n10951_), .A2(new_n10947_), .B(new_n11002_), .ZN(new_n11440_));
  INV_X1     g11154(.I(new_n11421_), .ZN(new_n11441_));
  OAI22_X1   g11155(.A1(new_n11440_), .A2(new_n11004_), .B1(new_n11441_), .B2(new_n11422_), .ZN(new_n11442_));
  OAI21_X1   g11156(.A1(new_n11430_), .A2(new_n11431_), .B(new_n11420_), .ZN(new_n11443_));
  NAND3_X1   g11157(.A1(new_n11405_), .A2(new_n11409_), .A3(new_n11428_), .ZN(new_n11444_));
  NAND2_X1   g11158(.A1(new_n11443_), .A2(new_n11444_), .ZN(new_n11445_));
  NAND3_X1   g11159(.A1(new_n11445_), .A2(new_n11389_), .A3(new_n11003_), .ZN(new_n11446_));
  XOR2_X1    g11160(.A1(new_n522_), .A2(new_n11437_), .Z(new_n11447_));
  AOI21_X1   g11161(.A1(new_n11442_), .A2(new_n11446_), .B(new_n11447_), .ZN(new_n11448_));
  NOR2_X1    g11162(.A1(new_n11439_), .A2(new_n11448_), .ZN(new_n11449_));
  NOR3_X1    g11163(.A1(new_n11449_), .A2(new_n11034_), .A3(new_n11022_), .ZN(new_n11450_));
  NOR2_X1    g11164(.A1(new_n11016_), .A2(new_n11010_), .ZN(new_n11452_));
  OAI21_X1   g11165(.A1(new_n11450_), .A2(new_n11452_), .B(new_n11037_), .ZN(new_n11453_));
  NAND3_X1   g11166(.A1(new_n11442_), .A2(new_n11446_), .A3(new_n11447_), .ZN(new_n11454_));
  OAI21_X1   g11167(.A1(new_n11434_), .A2(new_n11424_), .B(new_n11438_), .ZN(new_n11455_));
  NAND2_X1   g11168(.A1(new_n11455_), .A2(new_n11454_), .ZN(new_n11456_));
  NAND3_X1   g11169(.A1(new_n11456_), .A2(new_n11012_), .A3(new_n11040_), .ZN(new_n11457_));
  INV_X1     g11170(.I(new_n11452_), .ZN(new_n11458_));
  NAND3_X1   g11171(.A1(new_n11457_), .A2(new_n11019_), .A3(new_n11458_), .ZN(new_n11459_));
  OAI22_X1   g11172(.A1(new_n7619_), .A2(new_n656_), .B1(new_n706_), .B2(new_n8309_), .ZN(new_n11460_));
  OAI21_X1   g11173(.A1(new_n565_), .A2(new_n7947_), .B(new_n11460_), .ZN(new_n11461_));
  AOI21_X1   g11174(.A1(new_n11461_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n11462_));
  XNOR2_X1   g11175(.A1(new_n710_), .A2(new_n11462_), .ZN(new_n11463_));
  AOI21_X1   g11176(.A1(new_n11453_), .A2(new_n11459_), .B(new_n11463_), .ZN(new_n11464_));
  AOI21_X1   g11177(.A1(new_n11457_), .A2(new_n11458_), .B(new_n11019_), .ZN(new_n11465_));
  NOR3_X1    g11178(.A1(new_n11450_), .A2(new_n11037_), .A3(new_n11452_), .ZN(new_n11466_));
  INV_X1     g11179(.I(new_n11463_), .ZN(new_n11467_));
  NOR3_X1    g11180(.A1(new_n11466_), .A2(new_n11465_), .A3(new_n11467_), .ZN(new_n11468_));
  OAI21_X1   g11181(.A1(new_n11468_), .A2(new_n11464_), .B(new_n11045_), .ZN(new_n11469_));
  NOR2_X1    g11182(.A1(new_n11469_), .A2(new_n11029_), .ZN(new_n11470_));
  OAI21_X1   g11183(.A1(new_n11466_), .A2(new_n11465_), .B(new_n11467_), .ZN(new_n11471_));
  NAND3_X1   g11184(.A1(new_n11453_), .A2(new_n11459_), .A3(new_n11463_), .ZN(new_n11472_));
  NAND2_X1   g11185(.A1(new_n11471_), .A2(new_n11472_), .ZN(new_n11473_));
  NOR2_X1    g11186(.A1(new_n11024_), .A2(new_n11028_), .ZN(new_n11475_));
  OAI21_X1   g11187(.A1(new_n11470_), .A2(new_n11475_), .B(new_n10941_), .ZN(new_n11476_));
  INV_X1     g11188(.I(new_n10941_), .ZN(new_n11477_));
  NAND3_X1   g11189(.A1(new_n11473_), .A2(new_n11030_), .A3(new_n11045_), .ZN(new_n11478_));
  INV_X1     g11190(.I(new_n11475_), .ZN(new_n11479_));
  NAND3_X1   g11191(.A1(new_n11478_), .A2(new_n11477_), .A3(new_n11479_), .ZN(new_n11480_));
  OAI22_X1   g11192(.A1(new_n6644_), .A2(new_n861_), .B1(new_n930_), .B2(new_n6647_), .ZN(new_n11481_));
  OAI21_X1   g11193(.A1(new_n780_), .A2(new_n7284_), .B(new_n11481_), .ZN(new_n11482_));
  AOI21_X1   g11194(.A1(new_n11482_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n11483_));
  XNOR2_X1   g11195(.A1(new_n937_), .A2(new_n11483_), .ZN(new_n11484_));
  INV_X1     g11196(.I(new_n11484_), .ZN(new_n11485_));
  NAND3_X1   g11197(.A1(new_n11476_), .A2(new_n11480_), .A3(new_n11485_), .ZN(new_n11486_));
  AOI21_X1   g11198(.A1(new_n11478_), .A2(new_n11479_), .B(new_n11477_), .ZN(new_n11487_));
  NOR3_X1    g11199(.A1(new_n11470_), .A2(new_n10941_), .A3(new_n11475_), .ZN(new_n11488_));
  OAI21_X1   g11200(.A1(new_n11488_), .A2(new_n11487_), .B(new_n11484_), .ZN(new_n11489_));
  NAND2_X1   g11201(.A1(new_n11489_), .A2(new_n11486_), .ZN(new_n11490_));
  INV_X1     g11202(.I(new_n11052_), .ZN(new_n11491_));
  NAND2_X1   g11203(.A1(new_n11048_), .A2(new_n11491_), .ZN(new_n11492_));
  OAI21_X1   g11204(.A1(new_n11047_), .A2(new_n11032_), .B(new_n11052_), .ZN(new_n11493_));
  NAND2_X1   g11205(.A1(new_n11492_), .A2(new_n11493_), .ZN(new_n11494_));
  NAND3_X1   g11206(.A1(new_n11490_), .A2(new_n11054_), .A3(new_n11494_), .ZN(new_n11495_));
  NOR2_X1    g11207(.A1(new_n11048_), .A2(new_n11052_), .ZN(new_n11497_));
  INV_X1     g11208(.I(new_n11497_), .ZN(new_n11498_));
  AOI21_X1   g11209(.A1(new_n11495_), .A2(new_n11498_), .B(new_n10933_), .ZN(new_n11499_));
  NOR3_X1    g11210(.A1(new_n11488_), .A2(new_n11487_), .A3(new_n11484_), .ZN(new_n11500_));
  AOI21_X1   g11211(.A1(new_n11476_), .A2(new_n11480_), .B(new_n11485_), .ZN(new_n11501_));
  OAI21_X1   g11212(.A1(new_n11500_), .A2(new_n11501_), .B(new_n11494_), .ZN(new_n11502_));
  NOR2_X1    g11213(.A1(new_n11502_), .A2(new_n11053_), .ZN(new_n11503_));
  NOR3_X1    g11214(.A1(new_n11503_), .A2(new_n10934_), .A3(new_n11497_), .ZN(new_n11504_));
  OAI22_X1   g11215(.A1(new_n5993_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n5991_), .ZN(new_n11505_));
  OAI21_X1   g11216(.A1(new_n1017_), .A2(new_n5997_), .B(new_n11505_), .ZN(new_n11506_));
  AOI21_X1   g11217(.A1(new_n11506_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n11507_));
  XNOR2_X1   g11218(.A1(new_n1196_), .A2(new_n11507_), .ZN(new_n11508_));
  NOR3_X1    g11219(.A1(new_n11504_), .A2(new_n11499_), .A3(new_n11508_), .ZN(new_n11509_));
  OAI21_X1   g11220(.A1(new_n11503_), .A2(new_n11497_), .B(new_n10934_), .ZN(new_n11510_));
  NAND3_X1   g11221(.A1(new_n11495_), .A2(new_n10933_), .A3(new_n11498_), .ZN(new_n11511_));
  INV_X1     g11222(.I(new_n11508_), .ZN(new_n11512_));
  AOI21_X1   g11223(.A1(new_n11510_), .A2(new_n11511_), .B(new_n11512_), .ZN(new_n11513_));
  OAI21_X1   g11224(.A1(new_n11509_), .A2(new_n11513_), .B(new_n11388_), .ZN(new_n11514_));
  AOI21_X1   g11225(.A1(new_n11062_), .A2(new_n11060_), .B(new_n10927_), .ZN(new_n11515_));
  NAND3_X1   g11226(.A1(new_n11062_), .A2(new_n11060_), .A3(new_n10927_), .ZN(new_n11516_));
  AOI21_X1   g11227(.A1(new_n11516_), .A2(new_n11386_), .B(new_n11515_), .ZN(new_n11517_));
  OAI21_X1   g11228(.A1(new_n11504_), .A2(new_n11499_), .B(new_n11512_), .ZN(new_n11518_));
  NAND3_X1   g11229(.A1(new_n11510_), .A2(new_n11511_), .A3(new_n11508_), .ZN(new_n11519_));
  NAND2_X1   g11230(.A1(new_n11518_), .A2(new_n11519_), .ZN(new_n11520_));
  NAND2_X1   g11231(.A1(new_n11520_), .A2(new_n11517_), .ZN(new_n11521_));
  OAI22_X1   g11232(.A1(new_n5420_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n5107_), .ZN(new_n11522_));
  OAI21_X1   g11233(.A1(new_n1294_), .A2(new_n5112_), .B(new_n11522_), .ZN(new_n11523_));
  AOI21_X1   g11234(.A1(new_n11523_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n11524_));
  XOR2_X1    g11235(.A1(new_n1530_), .A2(new_n11524_), .Z(new_n11525_));
  AOI21_X1   g11236(.A1(new_n11521_), .A2(new_n11514_), .B(new_n11525_), .ZN(new_n11526_));
  NAND2_X1   g11237(.A1(new_n11516_), .A2(new_n11386_), .ZN(new_n11527_));
  NAND3_X1   g11238(.A1(new_n11510_), .A2(new_n11511_), .A3(new_n11512_), .ZN(new_n11528_));
  OAI21_X1   g11239(.A1(new_n11504_), .A2(new_n11499_), .B(new_n11508_), .ZN(new_n11529_));
  AOI22_X1   g11240(.A1(new_n11384_), .A2(new_n11527_), .B1(new_n11529_), .B2(new_n11528_), .ZN(new_n11530_));
  AOI21_X1   g11241(.A1(new_n11518_), .A2(new_n11519_), .B(new_n11388_), .ZN(new_n11531_));
  INV_X1     g11242(.I(new_n11525_), .ZN(new_n11532_));
  NOR3_X1    g11243(.A1(new_n11531_), .A2(new_n11530_), .A3(new_n11532_), .ZN(new_n11533_));
  NOR2_X1    g11244(.A1(new_n11526_), .A2(new_n11533_), .ZN(new_n11534_));
  NOR2_X1    g11245(.A1(new_n11383_), .A2(new_n11534_), .ZN(new_n11535_));
  OAI21_X1   g11246(.A1(new_n11083_), .A2(new_n11080_), .B(new_n11094_), .ZN(new_n11536_));
  NOR3_X1    g11247(.A1(new_n11531_), .A2(new_n11530_), .A3(new_n11525_), .ZN(new_n11537_));
  AOI21_X1   g11248(.A1(new_n11521_), .A2(new_n11514_), .B(new_n11532_), .ZN(new_n11538_));
  NOR2_X1    g11249(.A1(new_n11538_), .A2(new_n11537_), .ZN(new_n11539_));
  NOR2_X1    g11250(.A1(new_n11536_), .A2(new_n11539_), .ZN(new_n11540_));
  OAI22_X1   g11251(.A1(new_n4072_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n4067_), .ZN(new_n11541_));
  OAI21_X1   g11252(.A1(new_n1634_), .A2(new_n4318_), .B(new_n11541_), .ZN(new_n11542_));
  AOI21_X1   g11253(.A1(new_n11542_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n11543_));
  XNOR2_X1   g11254(.A1(new_n1940_), .A2(new_n11543_), .ZN(new_n11544_));
  NOR3_X1    g11255(.A1(new_n11535_), .A2(new_n11540_), .A3(new_n11544_), .ZN(new_n11545_));
  OAI21_X1   g11256(.A1(new_n11531_), .A2(new_n11530_), .B(new_n11532_), .ZN(new_n11546_));
  NAND3_X1   g11257(.A1(new_n11521_), .A2(new_n11514_), .A3(new_n11525_), .ZN(new_n11547_));
  NAND2_X1   g11258(.A1(new_n11547_), .A2(new_n11546_), .ZN(new_n11548_));
  NAND2_X1   g11259(.A1(new_n11536_), .A2(new_n11548_), .ZN(new_n11549_));
  NAND3_X1   g11260(.A1(new_n11521_), .A2(new_n11514_), .A3(new_n11532_), .ZN(new_n11550_));
  OAI21_X1   g11261(.A1(new_n11531_), .A2(new_n11530_), .B(new_n11525_), .ZN(new_n11551_));
  NAND2_X1   g11262(.A1(new_n11550_), .A2(new_n11551_), .ZN(new_n11552_));
  NAND2_X1   g11263(.A1(new_n11383_), .A2(new_n11552_), .ZN(new_n11553_));
  INV_X1     g11264(.I(new_n11544_), .ZN(new_n11554_));
  AOI21_X1   g11265(.A1(new_n11553_), .A2(new_n11549_), .B(new_n11554_), .ZN(new_n11555_));
  NOR2_X1    g11266(.A1(new_n11545_), .A2(new_n11555_), .ZN(new_n11556_));
  NOR2_X1    g11267(.A1(new_n11556_), .A2(new_n11382_), .ZN(new_n11557_));
  OAI21_X1   g11268(.A1(new_n11099_), .A2(new_n11096_), .B(new_n11100_), .ZN(new_n11558_));
  OAI21_X1   g11269(.A1(new_n11118_), .A2(new_n11101_), .B(new_n11558_), .ZN(new_n11559_));
  NAND3_X1   g11270(.A1(new_n11553_), .A2(new_n11549_), .A3(new_n11554_), .ZN(new_n11560_));
  OAI21_X1   g11271(.A1(new_n11535_), .A2(new_n11540_), .B(new_n11544_), .ZN(new_n11561_));
  NAND2_X1   g11272(.A1(new_n11561_), .A2(new_n11560_), .ZN(new_n11562_));
  NOR2_X1    g11273(.A1(new_n11562_), .A2(new_n11559_), .ZN(new_n11563_));
  NOR2_X1    g11274(.A1(new_n11563_), .A2(new_n11557_), .ZN(new_n11564_));
  AOI21_X1   g11275(.A1(new_n11107_), .A2(new_n11104_), .B(new_n10921_), .ZN(new_n11565_));
  NOR2_X1    g11276(.A1(new_n11102_), .A2(new_n11112_), .ZN(new_n11566_));
  NOR3_X1    g11277(.A1(new_n11118_), .A2(new_n11093_), .A3(new_n11101_), .ZN(new_n11567_));
  NOR2_X1    g11278(.A1(new_n11566_), .A2(new_n11567_), .ZN(new_n11568_));
  AOI21_X1   g11279(.A1(new_n11128_), .A2(new_n10921_), .B(new_n11568_), .ZN(new_n11569_));
  OAI22_X1   g11280(.A1(new_n2842_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n3018_), .ZN(new_n11570_));
  OAI21_X1   g11281(.A1(new_n2643_), .A2(new_n2884_), .B(new_n11570_), .ZN(new_n11571_));
  AOI21_X1   g11282(.A1(new_n11571_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n11572_));
  XNOR2_X1   g11283(.A1(new_n3022_), .A2(new_n11572_), .ZN(new_n11573_));
  NOR3_X1    g11284(.A1(new_n11569_), .A2(new_n11565_), .A3(new_n11573_), .ZN(new_n11574_));
  NAND2_X1   g11285(.A1(new_n11115_), .A2(new_n11132_), .ZN(new_n11575_));
  INV_X1     g11286(.I(new_n11568_), .ZN(new_n11576_));
  OAI21_X1   g11287(.A1(new_n11115_), .A2(new_n11132_), .B(new_n11576_), .ZN(new_n11577_));
  INV_X1     g11288(.I(new_n11573_), .ZN(new_n11578_));
  AOI21_X1   g11289(.A1(new_n11577_), .A2(new_n11575_), .B(new_n11578_), .ZN(new_n11579_));
  OAI21_X1   g11290(.A1(new_n11574_), .A2(new_n11579_), .B(new_n11564_), .ZN(new_n11580_));
  INV_X1     g11291(.I(new_n11564_), .ZN(new_n11581_));
  NAND3_X1   g11292(.A1(new_n11577_), .A2(new_n11575_), .A3(new_n11578_), .ZN(new_n11582_));
  OAI21_X1   g11293(.A1(new_n11569_), .A2(new_n11565_), .B(new_n11573_), .ZN(new_n11583_));
  NAND3_X1   g11294(.A1(new_n11583_), .A2(new_n11582_), .A3(new_n11581_), .ZN(new_n11584_));
  AOI21_X1   g11295(.A1(new_n11580_), .A2(new_n11584_), .B(new_n11380_), .ZN(new_n11585_));
  AOI21_X1   g11296(.A1(new_n11583_), .A2(new_n11582_), .B(new_n11581_), .ZN(new_n11586_));
  NOR3_X1    g11297(.A1(new_n11574_), .A2(new_n11579_), .A3(new_n11564_), .ZN(new_n11587_));
  NOR3_X1    g11298(.A1(new_n11587_), .A2(new_n11586_), .A3(new_n11379_), .ZN(new_n11588_));
  NOR3_X1    g11299(.A1(new_n11588_), .A2(new_n11585_), .A3(new_n11160_), .ZN(new_n11589_));
  NOR3_X1    g11300(.A1(new_n11589_), .A2(new_n11163_), .A3(new_n11145_), .ZN(new_n11590_));
  OAI21_X1   g11301(.A1(new_n11587_), .A2(new_n11586_), .B(new_n11379_), .ZN(new_n11591_));
  NAND3_X1   g11302(.A1(new_n11580_), .A2(new_n11584_), .A3(new_n11380_), .ZN(new_n11592_));
  NAND3_X1   g11303(.A1(new_n11591_), .A2(new_n11592_), .A3(new_n11144_), .ZN(new_n11593_));
  AOI21_X1   g11304(.A1(new_n11593_), .A2(new_n11149_), .B(new_n11161_), .ZN(new_n11594_));
  OAI22_X1   g11305(.A1(new_n2171_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n2166_), .ZN(new_n11595_));
  OAI21_X1   g11306(.A1(new_n3260_), .A2(new_n2322_), .B(new_n11595_), .ZN(new_n11596_));
  AOI21_X1   g11307(.A1(new_n11596_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n11597_));
  XOR2_X1    g11308(.A1(new_n3722_), .A2(new_n11597_), .Z(new_n11598_));
  INV_X1     g11309(.I(new_n11598_), .ZN(new_n11599_));
  OAI21_X1   g11310(.A1(new_n11590_), .A2(new_n11594_), .B(new_n11599_), .ZN(new_n11600_));
  NAND3_X1   g11311(.A1(new_n11593_), .A2(new_n11161_), .A3(new_n11149_), .ZN(new_n11601_));
  OAI21_X1   g11312(.A1(new_n11589_), .A2(new_n11163_), .B(new_n11145_), .ZN(new_n11602_));
  NAND3_X1   g11313(.A1(new_n11602_), .A2(new_n11601_), .A3(new_n11598_), .ZN(new_n11603_));
  NAND3_X1   g11314(.A1(new_n11600_), .A2(new_n11603_), .A3(new_n11375_), .ZN(new_n11604_));
  NAND3_X1   g11315(.A1(new_n11604_), .A2(new_n11166_), .A3(new_n11177_), .ZN(new_n11605_));
  NAND2_X1   g11316(.A1(new_n11161_), .A2(new_n11149_), .ZN(new_n11606_));
  NAND2_X1   g11317(.A1(new_n11145_), .A2(new_n11163_), .ZN(new_n11607_));
  AOI21_X1   g11318(.A1(new_n11607_), .A2(new_n11606_), .B(new_n11154_), .ZN(new_n11608_));
  AOI21_X1   g11319(.A1(new_n11602_), .A2(new_n11601_), .B(new_n11598_), .ZN(new_n11609_));
  NOR3_X1    g11320(.A1(new_n11590_), .A2(new_n11594_), .A3(new_n11599_), .ZN(new_n11610_));
  NOR3_X1    g11321(.A1(new_n11610_), .A2(new_n11609_), .A3(new_n11608_), .ZN(new_n11611_));
  OAI21_X1   g11322(.A1(new_n11611_), .A2(new_n11369_), .B(new_n10917_), .ZN(new_n11612_));
  OAI22_X1   g11323(.A1(new_n1712_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n1707_), .ZN(new_n11613_));
  OAI21_X1   g11324(.A1(new_n3989_), .A2(new_n1850_), .B(new_n11613_), .ZN(new_n11614_));
  AOI21_X1   g11325(.A1(new_n11614_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n11615_));
  XOR2_X1    g11326(.A1(new_n4499_), .A2(new_n11615_), .Z(new_n11616_));
  INV_X1     g11327(.I(new_n11616_), .ZN(new_n11617_));
  NAND3_X1   g11328(.A1(new_n11612_), .A2(new_n11605_), .A3(new_n11617_), .ZN(new_n11618_));
  NOR3_X1    g11329(.A1(new_n11611_), .A2(new_n11369_), .A3(new_n10917_), .ZN(new_n11619_));
  AOI21_X1   g11330(.A1(new_n11604_), .A2(new_n11166_), .B(new_n11177_), .ZN(new_n11620_));
  OAI21_X1   g11331(.A1(new_n11619_), .A2(new_n11620_), .B(new_n11616_), .ZN(new_n11621_));
  NAND3_X1   g11332(.A1(new_n11621_), .A2(new_n11618_), .A3(new_n11372_), .ZN(new_n11622_));
  NAND3_X1   g11333(.A1(new_n11622_), .A2(new_n11194_), .A3(new_n11195_), .ZN(new_n11623_));
  NAND2_X1   g11334(.A1(new_n11177_), .A2(new_n11166_), .ZN(new_n11624_));
  NAND2_X1   g11335(.A1(new_n11369_), .A2(new_n10917_), .ZN(new_n11625_));
  AOI21_X1   g11336(.A1(new_n11625_), .A2(new_n11624_), .B(new_n11171_), .ZN(new_n11626_));
  NOR3_X1    g11337(.A1(new_n11619_), .A2(new_n11620_), .A3(new_n11616_), .ZN(new_n11627_));
  AOI21_X1   g11338(.A1(new_n11612_), .A2(new_n11605_), .B(new_n11617_), .ZN(new_n11628_));
  NOR3_X1    g11339(.A1(new_n11627_), .A2(new_n11628_), .A3(new_n11626_), .ZN(new_n11629_));
  OAI21_X1   g11340(.A1(new_n11629_), .A2(new_n11208_), .B(new_n10911_), .ZN(new_n11630_));
  OAI22_X1   g11341(.A1(new_n1347_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n1344_), .ZN(new_n11631_));
  OAI21_X1   g11342(.A1(new_n4774_), .A2(new_n1457_), .B(new_n11631_), .ZN(new_n11632_));
  AOI21_X1   g11343(.A1(new_n11632_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n11633_));
  XNOR2_X1   g11344(.A1(new_n5357_), .A2(new_n11633_), .ZN(new_n11634_));
  INV_X1     g11345(.I(new_n11634_), .ZN(new_n11635_));
  NAND3_X1   g11346(.A1(new_n11630_), .A2(new_n11623_), .A3(new_n11635_), .ZN(new_n11636_));
  NOR3_X1    g11347(.A1(new_n11629_), .A2(new_n10911_), .A3(new_n11208_), .ZN(new_n11637_));
  AOI21_X1   g11348(.A1(new_n11622_), .A2(new_n11195_), .B(new_n11194_), .ZN(new_n11638_));
  OAI21_X1   g11349(.A1(new_n11637_), .A2(new_n11638_), .B(new_n11634_), .ZN(new_n11639_));
  NAND3_X1   g11350(.A1(new_n11639_), .A2(new_n11636_), .A3(new_n11368_), .ZN(new_n11640_));
  NAND3_X1   g11351(.A1(new_n11640_), .A2(new_n10907_), .A3(new_n11199_), .ZN(new_n11641_));
  NAND2_X1   g11352(.A1(new_n11194_), .A2(new_n11195_), .ZN(new_n11642_));
  NAND2_X1   g11353(.A1(new_n11208_), .A2(new_n10911_), .ZN(new_n11643_));
  AOI21_X1   g11354(.A1(new_n11642_), .A2(new_n11643_), .B(new_n11189_), .ZN(new_n11644_));
  NOR3_X1    g11355(.A1(new_n11637_), .A2(new_n11638_), .A3(new_n11634_), .ZN(new_n11645_));
  AOI21_X1   g11356(.A1(new_n11630_), .A2(new_n11623_), .B(new_n11635_), .ZN(new_n11646_));
  NOR3_X1    g11357(.A1(new_n11645_), .A2(new_n11646_), .A3(new_n11644_), .ZN(new_n11647_));
  OAI21_X1   g11358(.A1(new_n11647_), .A2(new_n11212_), .B(new_n11221_), .ZN(new_n11648_));
  OAI22_X1   g11359(.A1(new_n1055_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n1061_), .ZN(new_n11649_));
  OAI21_X1   g11360(.A1(new_n5913_), .A2(new_n1332_), .B(new_n11649_), .ZN(new_n11650_));
  AOI21_X1   g11361(.A1(new_n11650_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n11651_));
  XOR2_X1    g11362(.A1(new_n6233_), .A2(new_n11651_), .Z(new_n11652_));
  INV_X1     g11363(.I(new_n11652_), .ZN(new_n11653_));
  NAND3_X1   g11364(.A1(new_n11648_), .A2(new_n11641_), .A3(new_n11653_), .ZN(new_n11654_));
  INV_X1     g11365(.I(new_n11641_), .ZN(new_n11655_));
  AOI21_X1   g11366(.A1(new_n11640_), .A2(new_n11199_), .B(new_n10907_), .ZN(new_n11656_));
  OAI21_X1   g11367(.A1(new_n11655_), .A2(new_n11656_), .B(new_n11652_), .ZN(new_n11657_));
  NAND3_X1   g11368(.A1(new_n11657_), .A2(new_n11365_), .A3(new_n11654_), .ZN(new_n11658_));
  NAND3_X1   g11369(.A1(new_n11658_), .A2(new_n11363_), .A3(new_n11215_), .ZN(new_n11659_));
  XOR2_X1    g11370(.A1(new_n11221_), .A2(new_n11212_), .Z(new_n11660_));
  NOR2_X1    g11371(.A1(new_n11660_), .A2(new_n11204_), .ZN(new_n11661_));
  NOR3_X1    g11372(.A1(new_n11655_), .A2(new_n11656_), .A3(new_n11652_), .ZN(new_n11662_));
  AOI21_X1   g11373(.A1(new_n11648_), .A2(new_n11641_), .B(new_n11653_), .ZN(new_n11663_));
  NOR3_X1    g11374(.A1(new_n11662_), .A2(new_n11661_), .A3(new_n11663_), .ZN(new_n11664_));
  OAI21_X1   g11375(.A1(new_n11664_), .A2(new_n11224_), .B(new_n11217_), .ZN(new_n11665_));
  NAND2_X1   g11376(.A1(new_n11665_), .A2(new_n11659_), .ZN(new_n11666_));
  INV_X1     g11377(.I(new_n11666_), .ZN(new_n11667_));
  INV_X1     g11378(.I(new_n11231_), .ZN(new_n11668_));
  AOI21_X1   g11379(.A1(new_n11225_), .A2(new_n11216_), .B(new_n11230_), .ZN(new_n11669_));
  AOI21_X1   g11380(.A1(new_n10899_), .A2(new_n10897_), .B(new_n11669_), .ZN(new_n11670_));
  OAI22_X1   g11381(.A1(new_n607_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n610_), .ZN(new_n11671_));
  OAI21_X1   g11382(.A1(new_n7864_), .A2(new_n684_), .B(new_n11671_), .ZN(new_n11672_));
  AOI21_X1   g11383(.A1(new_n11672_), .A2(new_n612_), .B(new_n607_), .ZN(new_n11673_));
  XOR2_X1    g11384(.A1(new_n8217_), .A2(new_n11673_), .Z(new_n11674_));
  NOR3_X1    g11385(.A1(new_n11670_), .A2(new_n11668_), .A3(new_n11674_), .ZN(new_n11675_));
  OAI21_X1   g11386(.A1(new_n11238_), .A2(new_n11236_), .B(new_n11234_), .ZN(new_n11676_));
  INV_X1     g11387(.I(new_n11674_), .ZN(new_n11677_));
  AOI21_X1   g11388(.A1(new_n11676_), .A2(new_n11231_), .B(new_n11677_), .ZN(new_n11678_));
  OAI21_X1   g11389(.A1(new_n11678_), .A2(new_n11675_), .B(new_n11667_), .ZN(new_n11679_));
  NAND3_X1   g11390(.A1(new_n11676_), .A2(new_n11231_), .A3(new_n11677_), .ZN(new_n11680_));
  OAI21_X1   g11391(.A1(new_n11670_), .A2(new_n11668_), .B(new_n11674_), .ZN(new_n11681_));
  NAND3_X1   g11392(.A1(new_n11680_), .A2(new_n11681_), .A3(new_n11666_), .ZN(new_n11682_));
  AOI21_X1   g11393(.A1(new_n11679_), .A2(new_n11682_), .B(new_n11362_), .ZN(new_n11683_));
  AOI21_X1   g11394(.A1(new_n11680_), .A2(new_n11681_), .B(new_n11666_), .ZN(new_n11684_));
  NOR3_X1    g11395(.A1(new_n11678_), .A2(new_n11675_), .A3(new_n11667_), .ZN(new_n11685_));
  NOR3_X1    g11396(.A1(new_n11684_), .A2(new_n11685_), .A3(new_n11361_), .ZN(new_n11686_));
  OAI21_X1   g11397(.A1(new_n11686_), .A2(new_n11683_), .B(new_n11266_), .ZN(new_n11687_));
  NOR2_X1    g11398(.A1(new_n11687_), .A2(new_n11254_), .ZN(new_n11688_));
  NOR2_X1    g11399(.A1(new_n11242_), .A2(new_n11235_), .ZN(new_n11689_));
  OAI21_X1   g11400(.A1(new_n11684_), .A2(new_n11685_), .B(new_n11361_), .ZN(new_n11690_));
  NAND3_X1   g11401(.A1(new_n11679_), .A2(new_n11682_), .A3(new_n11362_), .ZN(new_n11691_));
  NAND2_X1   g11402(.A1(new_n11690_), .A2(new_n11691_), .ZN(new_n11692_));
  NOR2_X1    g11403(.A1(new_n11689_), .A2(new_n11246_), .ZN(new_n11694_));
  OAI21_X1   g11404(.A1(new_n11688_), .A2(new_n11694_), .B(new_n11357_), .ZN(new_n11695_));
  NAND3_X1   g11405(.A1(new_n11692_), .A2(new_n11266_), .A3(new_n11253_), .ZN(new_n11696_));
  INV_X1     g11406(.I(new_n11694_), .ZN(new_n11697_));
  NAND3_X1   g11407(.A1(new_n11696_), .A2(new_n11251_), .A3(new_n11697_), .ZN(new_n11698_));
  OAI22_X1   g11408(.A1(new_n448_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n450_), .ZN(new_n11699_));
  OAI21_X1   g11409(.A1(new_n8563_), .A2(new_n496_), .B(new_n11699_), .ZN(new_n11700_));
  AOI21_X1   g11410(.A1(new_n11700_), .A2(new_n452_), .B(new_n448_), .ZN(new_n11701_));
  XNOR2_X1   g11411(.A1(new_n9299_), .A2(new_n11701_), .ZN(new_n11702_));
  INV_X1     g11412(.I(new_n11702_), .ZN(new_n11703_));
  NAND3_X1   g11413(.A1(new_n11695_), .A2(new_n11698_), .A3(new_n11703_), .ZN(new_n11704_));
  AOI21_X1   g11414(.A1(new_n11696_), .A2(new_n11697_), .B(new_n11251_), .ZN(new_n11705_));
  NOR3_X1    g11415(.A1(new_n11688_), .A2(new_n11357_), .A3(new_n11694_), .ZN(new_n11706_));
  OAI21_X1   g11416(.A1(new_n11706_), .A2(new_n11705_), .B(new_n11702_), .ZN(new_n11707_));
  NAND2_X1   g11417(.A1(new_n11707_), .A2(new_n11704_), .ZN(new_n11708_));
  NOR2_X1    g11418(.A1(new_n11257_), .A2(new_n11250_), .ZN(new_n11709_));
  XOR2_X1    g11419(.A1(new_n11709_), .A2(new_n11261_), .Z(new_n11710_));
  NAND3_X1   g11420(.A1(new_n11708_), .A2(new_n11263_), .A3(new_n11710_), .ZN(new_n11711_));
  NOR2_X1    g11421(.A1(new_n11709_), .A2(new_n11261_), .ZN(new_n11713_));
  INV_X1     g11422(.I(new_n11713_), .ZN(new_n11714_));
  AOI21_X1   g11423(.A1(new_n11711_), .A2(new_n11714_), .B(new_n11356_), .ZN(new_n11715_));
  NAND3_X1   g11424(.A1(new_n11711_), .A2(new_n11356_), .A3(new_n11714_), .ZN(new_n11716_));
  INV_X1     g11425(.I(new_n11716_), .ZN(new_n11717_));
  OAI22_X1   g11426(.A1(new_n10031_), .A2(new_n341_), .B1(new_n404_), .B2(new_n10477_), .ZN(new_n11718_));
  OAI21_X1   g11427(.A1(new_n10025_), .A2(new_n366_), .B(new_n11718_), .ZN(new_n11719_));
  AOI21_X1   g11428(.A1(new_n11719_), .A2(new_n334_), .B(new_n341_), .ZN(new_n11720_));
  XOR2_X1    g11429(.A1(new_n10476_), .A2(new_n11720_), .Z(new_n11721_));
  INV_X1     g11430(.I(new_n11721_), .ZN(new_n11722_));
  OAI21_X1   g11431(.A1(new_n11717_), .A2(new_n11715_), .B(new_n11722_), .ZN(new_n11723_));
  NOR2_X1    g11432(.A1(new_n11723_), .A2(new_n11355_), .ZN(new_n11724_));
  OAI21_X1   g11433(.A1(new_n11317_), .A2(new_n10846_), .B(new_n10493_), .ZN(new_n11725_));
  NAND2_X1   g11434(.A1(new_n11317_), .A2(new_n10846_), .ZN(new_n11726_));
  NAND3_X1   g11435(.A1(new_n11725_), .A2(new_n11726_), .A3(new_n10854_), .ZN(new_n11727_));
  INV_X1     g11436(.I(new_n11715_), .ZN(new_n11728_));
  NAND2_X1   g11437(.A1(new_n11728_), .A2(new_n11716_), .ZN(new_n11729_));
  AOI21_X1   g11438(.A1(new_n11729_), .A2(new_n11722_), .B(new_n11727_), .ZN(new_n11730_));
  OAI21_X1   g11439(.A1(new_n11730_), .A2(new_n11724_), .B(new_n11352_), .ZN(new_n11731_));
  NAND3_X1   g11440(.A1(new_n11729_), .A2(new_n11727_), .A3(new_n11722_), .ZN(new_n11732_));
  NAND2_X1   g11441(.A1(new_n11723_), .A2(new_n11355_), .ZN(new_n11733_));
  NAND3_X1   g11442(.A1(new_n11732_), .A2(new_n11733_), .A3(new_n11351_), .ZN(new_n11734_));
  NAND2_X1   g11443(.A1(new_n11731_), .A2(new_n11734_), .ZN(new_n11735_));
  NOR2_X1    g11444(.A1(\b[54] ), .A2(\b[55] ), .ZN(new_n11736_));
  AOI21_X1   g11445(.A1(new_n10860_), .A2(new_n11736_), .B(new_n10477_), .ZN(new_n11737_));
  INV_X1     g11446(.I(\b[55] ), .ZN(new_n11738_));
  NOR2_X1    g11447(.A1(new_n10862_), .A2(new_n11738_), .ZN(new_n11739_));
  INV_X1     g11448(.I(new_n11739_), .ZN(new_n11740_));
  NOR2_X1    g11449(.A1(new_n10860_), .A2(new_n11740_), .ZN(new_n11741_));
  NOR2_X1    g11450(.A1(new_n11737_), .A2(new_n11741_), .ZN(new_n11742_));
  XNOR2_X1   g11451(.A1(\b[55] ), .A2(\b[56] ), .ZN(new_n11743_));
  INV_X1     g11452(.I(\b[56] ), .ZN(new_n11744_));
  NOR2_X1    g11453(.A1(new_n11738_), .A2(new_n11744_), .ZN(new_n11745_));
  NOR2_X1    g11454(.A1(\b[55] ), .A2(\b[56] ), .ZN(new_n11746_));
  OAI21_X1   g11455(.A1(new_n11745_), .A2(new_n11746_), .B(new_n11742_), .ZN(new_n11747_));
  OAI21_X1   g11456(.A1(new_n11742_), .A2(new_n11743_), .B(new_n11747_), .ZN(new_n11748_));
  OAI22_X1   g11457(.A1(new_n330_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n263_), .ZN(new_n11749_));
  OAI21_X1   g11458(.A1(new_n10862_), .A2(new_n289_), .B(new_n11749_), .ZN(new_n11750_));
  AOI21_X1   g11459(.A1(new_n11750_), .A2(new_n260_), .B(new_n426_), .ZN(new_n11751_));
  XNOR2_X1   g11460(.A1(new_n11748_), .A2(new_n11751_), .ZN(new_n11752_));
  INV_X1     g11461(.I(new_n11752_), .ZN(new_n11753_));
  NAND2_X1   g11462(.A1(new_n11735_), .A2(new_n11753_), .ZN(new_n11754_));
  INV_X1     g11463(.I(new_n11735_), .ZN(new_n11755_));
  NAND2_X1   g11464(.A1(new_n11755_), .A2(new_n11752_), .ZN(new_n11756_));
  NAND2_X1   g11465(.A1(new_n11756_), .A2(new_n11754_), .ZN(new_n11757_));
  NAND2_X1   g11466(.A1(new_n11757_), .A2(new_n11347_), .ZN(new_n11758_));
  XOR2_X1    g11467(.A1(new_n11735_), .A2(new_n11752_), .Z(new_n11759_));
  OAI21_X1   g11468(.A1(new_n11347_), .A2(new_n11759_), .B(new_n11758_), .ZN(\f[56] ));
  NAND2_X1   g11469(.A1(new_n11729_), .A2(new_n11351_), .ZN(new_n11761_));
  NAND3_X1   g11470(.A1(new_n11352_), .A2(new_n11728_), .A3(new_n11716_), .ZN(new_n11762_));
  NOR4_X1    g11471(.A1(new_n11336_), .A2(new_n11353_), .A3(new_n11354_), .A4(new_n11721_), .ZN(new_n11763_));
  NAND2_X1   g11472(.A1(new_n11762_), .A2(new_n11763_), .ZN(new_n11764_));
  NAND2_X1   g11473(.A1(new_n11764_), .A2(new_n11761_), .ZN(new_n11765_));
  INV_X1     g11474(.I(new_n11709_), .ZN(new_n11766_));
  NOR3_X1    g11475(.A1(new_n11706_), .A2(new_n11705_), .A3(new_n11702_), .ZN(new_n11767_));
  AOI21_X1   g11476(.A1(new_n11695_), .A2(new_n11698_), .B(new_n11703_), .ZN(new_n11768_));
  OAI21_X1   g11477(.A1(new_n11767_), .A2(new_n11768_), .B(new_n11766_), .ZN(new_n11769_));
  NAND2_X1   g11478(.A1(new_n11769_), .A2(new_n11261_), .ZN(new_n11770_));
  NOR3_X1    g11479(.A1(new_n11767_), .A2(new_n11768_), .A3(new_n11766_), .ZN(new_n11771_));
  NOR2_X1    g11480(.A1(new_n11771_), .A2(new_n11349_), .ZN(new_n11772_));
  NOR2_X1    g11481(.A1(new_n11670_), .A2(new_n11668_), .ZN(new_n11773_));
  XOR2_X1    g11482(.A1(new_n11773_), .A2(new_n11666_), .Z(new_n11774_));
  NOR2_X1    g11483(.A1(new_n11774_), .A2(new_n11362_), .ZN(new_n11775_));
  XOR2_X1    g11484(.A1(new_n11773_), .A2(new_n11667_), .Z(new_n11776_));
  NOR2_X1    g11485(.A1(new_n11776_), .A2(new_n11361_), .ZN(new_n11777_));
  OAI21_X1   g11486(.A1(new_n11775_), .A2(new_n11777_), .B(new_n11677_), .ZN(new_n11778_));
  INV_X1     g11487(.I(new_n11778_), .ZN(new_n11779_));
  INV_X1     g11488(.I(new_n11689_), .ZN(new_n11780_));
  AOI21_X1   g11489(.A1(new_n11692_), .A2(new_n11252_), .B(new_n11780_), .ZN(new_n11781_));
  NAND3_X1   g11490(.A1(new_n11690_), .A2(new_n11691_), .A3(new_n11246_), .ZN(new_n11782_));
  NAND2_X1   g11491(.A1(new_n11782_), .A2(new_n11251_), .ZN(new_n11783_));
  NAND2_X1   g11492(.A1(new_n11666_), .A2(new_n11361_), .ZN(new_n11784_));
  NAND2_X1   g11493(.A1(new_n11676_), .A2(new_n11231_), .ZN(new_n11785_));
  NOR3_X1    g11494(.A1(new_n11664_), .A2(new_n11217_), .A3(new_n11224_), .ZN(new_n11786_));
  AOI21_X1   g11495(.A1(new_n11658_), .A2(new_n11215_), .B(new_n11363_), .ZN(new_n11787_));
  OAI21_X1   g11496(.A1(new_n11787_), .A2(new_n11786_), .B(new_n11362_), .ZN(new_n11788_));
  NAND3_X1   g11497(.A1(new_n11665_), .A2(new_n11659_), .A3(new_n11361_), .ZN(new_n11789_));
  NAND2_X1   g11498(.A1(new_n11788_), .A2(new_n11789_), .ZN(new_n11790_));
  INV_X1     g11499(.I(new_n11790_), .ZN(new_n11791_));
  NOR2_X1    g11500(.A1(new_n11791_), .A2(new_n11785_), .ZN(new_n11792_));
  AOI21_X1   g11501(.A1(new_n11657_), .A2(new_n11654_), .B(new_n11365_), .ZN(new_n11793_));
  OAI21_X1   g11502(.A1(new_n11793_), .A2(new_n11215_), .B(new_n11217_), .ZN(new_n11794_));
  OAI21_X1   g11503(.A1(new_n11645_), .A2(new_n11646_), .B(new_n11644_), .ZN(new_n11795_));
  AOI21_X1   g11504(.A1(new_n11795_), .A2(new_n11212_), .B(new_n10907_), .ZN(new_n11796_));
  AOI21_X1   g11505(.A1(new_n11621_), .A2(new_n11618_), .B(new_n11372_), .ZN(new_n11797_));
  OAI21_X1   g11506(.A1(new_n11797_), .A2(new_n11195_), .B(new_n10911_), .ZN(new_n11798_));
  AOI21_X1   g11507(.A1(new_n11602_), .A2(new_n11601_), .B(new_n11599_), .ZN(new_n11799_));
  INV_X1     g11508(.I(new_n11799_), .ZN(new_n11800_));
  OAI21_X1   g11509(.A1(new_n11610_), .A2(new_n11609_), .B(new_n11608_), .ZN(new_n11801_));
  AOI21_X1   g11510(.A1(new_n11801_), .A2(new_n11369_), .B(new_n11177_), .ZN(new_n11802_));
  NAND3_X1   g11511(.A1(new_n11107_), .A2(new_n10921_), .A3(new_n11104_), .ZN(new_n11803_));
  AOI21_X1   g11512(.A1(new_n11803_), .A2(new_n11576_), .B(new_n11565_), .ZN(new_n11804_));
  NAND2_X1   g11513(.A1(new_n11804_), .A2(new_n11581_), .ZN(new_n11805_));
  NAND2_X1   g11514(.A1(new_n11577_), .A2(new_n11575_), .ZN(new_n11806_));
  NAND2_X1   g11515(.A1(new_n11806_), .A2(new_n11564_), .ZN(new_n11807_));
  AOI21_X1   g11516(.A1(new_n11805_), .A2(new_n11807_), .B(new_n11380_), .ZN(new_n11808_));
  INV_X1     g11517(.I(new_n11808_), .ZN(new_n11809_));
  NAND3_X1   g11518(.A1(new_n11805_), .A2(new_n11807_), .A3(new_n11380_), .ZN(new_n11810_));
  AOI21_X1   g11519(.A1(new_n11809_), .A2(new_n11810_), .B(new_n11573_), .ZN(new_n11811_));
  AOI21_X1   g11520(.A1(new_n11591_), .A2(new_n11592_), .B(new_n11144_), .ZN(new_n11812_));
  OAI21_X1   g11521(.A1(new_n11812_), .A2(new_n11149_), .B(new_n11145_), .ZN(new_n11813_));
  OAI21_X1   g11522(.A1(new_n11563_), .A2(new_n11557_), .B(new_n11380_), .ZN(new_n11814_));
  NAND2_X1   g11523(.A1(new_n11562_), .A2(new_n11559_), .ZN(new_n11815_));
  NAND2_X1   g11524(.A1(new_n11556_), .A2(new_n11382_), .ZN(new_n11816_));
  NAND3_X1   g11525(.A1(new_n11815_), .A2(new_n11816_), .A3(new_n11379_), .ZN(new_n11817_));
  NAND2_X1   g11526(.A1(new_n11814_), .A2(new_n11817_), .ZN(new_n11818_));
  NAND3_X1   g11527(.A1(new_n11577_), .A2(new_n11575_), .A3(new_n11818_), .ZN(new_n11819_));
  NOR2_X1    g11528(.A1(new_n11564_), .A2(new_n11380_), .ZN(new_n11820_));
  NAND3_X1   g11529(.A1(new_n11553_), .A2(new_n11549_), .A3(new_n11544_), .ZN(new_n11821_));
  INV_X1     g11530(.I(new_n11821_), .ZN(new_n11822_));
  NOR2_X1    g11531(.A1(new_n11383_), .A2(new_n11533_), .ZN(new_n11823_));
  INV_X1     g11532(.I(new_n11048_), .ZN(new_n11824_));
  OAI21_X1   g11533(.A1(new_n11500_), .A2(new_n11501_), .B(new_n11824_), .ZN(new_n11825_));
  NAND2_X1   g11534(.A1(new_n11825_), .A2(new_n11052_), .ZN(new_n11826_));
  NOR3_X1    g11535(.A1(new_n11500_), .A2(new_n11501_), .A3(new_n11824_), .ZN(new_n11827_));
  NOR2_X1    g11536(.A1(new_n11827_), .A2(new_n10934_), .ZN(new_n11828_));
  AOI21_X1   g11537(.A1(new_n11453_), .A2(new_n11459_), .B(new_n11467_), .ZN(new_n11829_));
  INV_X1     g11538(.I(new_n11024_), .ZN(new_n11830_));
  AOI21_X1   g11539(.A1(new_n11473_), .A2(new_n11830_), .B(new_n11042_), .ZN(new_n11831_));
  OAI21_X1   g11540(.A1(new_n11473_), .A2(new_n11830_), .B(new_n11477_), .ZN(new_n11832_));
  NOR3_X1    g11541(.A1(new_n11434_), .A2(new_n11424_), .A3(new_n11447_), .ZN(new_n11833_));
  INV_X1     g11542(.I(new_n11833_), .ZN(new_n11834_));
  OAI21_X1   g11543(.A1(new_n11449_), .A2(new_n11016_), .B(new_n11010_), .ZN(new_n11835_));
  AOI21_X1   g11544(.A1(new_n11016_), .A2(new_n11449_), .B(new_n11037_), .ZN(new_n11836_));
  AOI21_X1   g11545(.A1(new_n11389_), .A2(new_n11003_), .B(new_n11422_), .ZN(new_n11837_));
  NOR2_X1    g11546(.A1(new_n11837_), .A2(new_n11441_), .ZN(new_n11838_));
  NAND2_X1   g11547(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n11839_));
  NOR2_X1    g11548(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n11840_));
  INV_X1     g11549(.I(new_n11840_), .ZN(new_n11841_));
  NAND2_X1   g11550(.A1(new_n11841_), .A2(new_n11839_), .ZN(new_n11842_));
  NOR3_X1    g11551(.A1(new_n11406_), .A2(new_n11404_), .A3(new_n11397_), .ZN(new_n11843_));
  INV_X1     g11552(.I(new_n11843_), .ZN(new_n11844_));
  OAI22_X1   g11553(.A1(new_n10979_), .A2(new_n10569_), .B1(new_n269_), .B2(new_n11401_), .ZN(new_n11845_));
  AOI21_X1   g11554(.A1(new_n11845_), .A2(new_n10973_), .B(new_n403_), .ZN(new_n11846_));
  XOR2_X1    g11555(.A1(new_n11846_), .A2(new_n10964_), .Z(new_n11847_));
  NOR3_X1    g11556(.A1(new_n11844_), .A2(new_n11842_), .A3(new_n11847_), .ZN(new_n11848_));
  INV_X1     g11557(.I(new_n11839_), .ZN(new_n11849_));
  NOR2_X1    g11558(.A1(new_n11849_), .A2(new_n11840_), .ZN(new_n11850_));
  INV_X1     g11559(.I(new_n11847_), .ZN(new_n11851_));
  AOI21_X1   g11560(.A1(new_n11851_), .A2(new_n11843_), .B(new_n11850_), .ZN(new_n11852_));
  OAI21_X1   g11561(.A1(new_n11852_), .A2(new_n11848_), .B(new_n258_), .ZN(new_n11853_));
  NAND3_X1   g11562(.A1(new_n11851_), .A2(new_n11843_), .A3(new_n11850_), .ZN(new_n11854_));
  OAI21_X1   g11563(.A1(new_n11844_), .A2(new_n11847_), .B(new_n11842_), .ZN(new_n11855_));
  NAND3_X1   g11564(.A1(new_n11854_), .A2(new_n11855_), .A3(\b[0] ), .ZN(new_n11856_));
  OAI22_X1   g11565(.A1(new_n11411_), .A2(new_n421_), .B1(new_n325_), .B2(new_n10137_), .ZN(new_n11857_));
  AOI21_X1   g11566(.A1(new_n11857_), .A2(new_n9718_), .B(new_n9713_), .ZN(new_n11858_));
  XOR2_X1    g11567(.A1(new_n425_), .A2(new_n11858_), .Z(new_n11859_));
  INV_X1     g11568(.I(new_n11859_), .ZN(new_n11860_));
  NAND3_X1   g11569(.A1(new_n11853_), .A2(new_n11856_), .A3(new_n11860_), .ZN(new_n11861_));
  AOI21_X1   g11570(.A1(new_n11853_), .A2(new_n11856_), .B(new_n11860_), .ZN(new_n11862_));
  INV_X1     g11571(.I(new_n11862_), .ZN(new_n11863_));
  AOI21_X1   g11572(.A1(new_n11863_), .A2(new_n11861_), .B(new_n11838_), .ZN(new_n11864_));
  AOI21_X1   g11573(.A1(new_n11853_), .A2(new_n11856_), .B(new_n11859_), .ZN(new_n11865_));
  AND3_X2    g11574(.A1(new_n11853_), .A2(new_n11856_), .A3(new_n11859_), .Z(new_n11866_));
  OAI21_X1   g11575(.A1(new_n11866_), .A2(new_n11865_), .B(new_n11838_), .ZN(new_n11867_));
  INV_X1     g11576(.I(new_n11867_), .ZN(new_n11868_));
  OAI22_X1   g11577(.A1(new_n8644_), .A2(new_n515_), .B1(new_n565_), .B2(new_n9388_), .ZN(new_n11869_));
  OAI21_X1   g11578(.A1(new_n472_), .A2(new_n10154_), .B(new_n11869_), .ZN(new_n11870_));
  AOI21_X1   g11579(.A1(new_n11870_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n11871_));
  XOR2_X1    g11580(.A1(new_n759_), .A2(new_n11871_), .Z(new_n11872_));
  INV_X1     g11581(.I(new_n11872_), .ZN(new_n11873_));
  OAI21_X1   g11582(.A1(new_n11868_), .A2(new_n11864_), .B(new_n11873_), .ZN(new_n11874_));
  AOI21_X1   g11583(.A1(new_n11835_), .A2(new_n11836_), .B(new_n11874_), .ZN(new_n11875_));
  AOI21_X1   g11584(.A1(new_n11456_), .A2(new_n11006_), .B(new_n11011_), .ZN(new_n11876_));
  OAI21_X1   g11585(.A1(new_n11006_), .A2(new_n11456_), .B(new_n11019_), .ZN(new_n11877_));
  INV_X1     g11586(.I(new_n11838_), .ZN(new_n11878_));
  INV_X1     g11587(.I(new_n11861_), .ZN(new_n11879_));
  OAI21_X1   g11588(.A1(new_n11879_), .A2(new_n11862_), .B(new_n11878_), .ZN(new_n11880_));
  AOI21_X1   g11589(.A1(new_n11880_), .A2(new_n11867_), .B(new_n11872_), .ZN(new_n11881_));
  NOR3_X1    g11590(.A1(new_n11881_), .A2(new_n11877_), .A3(new_n11876_), .ZN(new_n11882_));
  OAI21_X1   g11591(.A1(new_n11875_), .A2(new_n11882_), .B(new_n11834_), .ZN(new_n11883_));
  OAI21_X1   g11592(.A1(new_n11876_), .A2(new_n11877_), .B(new_n11881_), .ZN(new_n11884_));
  NAND3_X1   g11593(.A1(new_n11874_), .A2(new_n11836_), .A3(new_n11835_), .ZN(new_n11885_));
  NAND3_X1   g11594(.A1(new_n11885_), .A2(new_n11884_), .A3(new_n11833_), .ZN(new_n11886_));
  OAI22_X1   g11595(.A1(new_n7619_), .A2(new_n706_), .B1(new_n780_), .B2(new_n8309_), .ZN(new_n11887_));
  OAI21_X1   g11596(.A1(new_n656_), .A2(new_n7947_), .B(new_n11887_), .ZN(new_n11888_));
  AOI21_X1   g11597(.A1(new_n11888_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n11889_));
  XOR2_X1    g11598(.A1(new_n785_), .A2(new_n11889_), .Z(new_n11890_));
  AOI21_X1   g11599(.A1(new_n11883_), .A2(new_n11886_), .B(new_n11890_), .ZN(new_n11891_));
  OAI21_X1   g11600(.A1(new_n11832_), .A2(new_n11831_), .B(new_n11891_), .ZN(new_n11892_));
  OAI21_X1   g11601(.A1(new_n11468_), .A2(new_n11464_), .B(new_n11830_), .ZN(new_n11893_));
  NAND2_X1   g11602(.A1(new_n11893_), .A2(new_n11028_), .ZN(new_n11894_));
  NOR3_X1    g11603(.A1(new_n11468_), .A2(new_n11464_), .A3(new_n11830_), .ZN(new_n11895_));
  NOR2_X1    g11604(.A1(new_n11895_), .A2(new_n10941_), .ZN(new_n11896_));
  AOI21_X1   g11605(.A1(new_n11885_), .A2(new_n11884_), .B(new_n11833_), .ZN(new_n11897_));
  NOR3_X1    g11606(.A1(new_n11875_), .A2(new_n11834_), .A3(new_n11882_), .ZN(new_n11898_));
  INV_X1     g11607(.I(new_n11890_), .ZN(new_n11899_));
  OAI21_X1   g11608(.A1(new_n11898_), .A2(new_n11897_), .B(new_n11899_), .ZN(new_n11900_));
  NAND3_X1   g11609(.A1(new_n11896_), .A2(new_n11900_), .A3(new_n11894_), .ZN(new_n11901_));
  AOI21_X1   g11610(.A1(new_n11892_), .A2(new_n11901_), .B(new_n11829_), .ZN(new_n11902_));
  INV_X1     g11611(.I(new_n11829_), .ZN(new_n11903_));
  AOI21_X1   g11612(.A1(new_n11894_), .A2(new_n11896_), .B(new_n11900_), .ZN(new_n11904_));
  NOR3_X1    g11613(.A1(new_n11891_), .A2(new_n11832_), .A3(new_n11831_), .ZN(new_n11905_));
  NOR3_X1    g11614(.A1(new_n11904_), .A2(new_n11905_), .A3(new_n11903_), .ZN(new_n11906_));
  OAI22_X1   g11615(.A1(new_n6644_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n6647_), .ZN(new_n11907_));
  OAI21_X1   g11616(.A1(new_n861_), .A2(new_n7284_), .B(new_n11907_), .ZN(new_n11908_));
  AOI21_X1   g11617(.A1(new_n11908_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n11909_));
  XOR2_X1    g11618(.A1(new_n1024_), .A2(new_n11909_), .Z(new_n11910_));
  INV_X1     g11619(.I(new_n11910_), .ZN(new_n11911_));
  OAI21_X1   g11620(.A1(new_n11902_), .A2(new_n11906_), .B(new_n11911_), .ZN(new_n11912_));
  AOI21_X1   g11621(.A1(new_n11828_), .A2(new_n11826_), .B(new_n11912_), .ZN(new_n11913_));
  AOI21_X1   g11622(.A1(new_n11490_), .A2(new_n11824_), .B(new_n11491_), .ZN(new_n11914_));
  NAND3_X1   g11623(.A1(new_n11489_), .A2(new_n11486_), .A3(new_n11048_), .ZN(new_n11915_));
  NAND2_X1   g11624(.A1(new_n11915_), .A2(new_n10933_), .ZN(new_n11916_));
  OAI21_X1   g11625(.A1(new_n11904_), .A2(new_n11905_), .B(new_n11903_), .ZN(new_n11917_));
  NAND3_X1   g11626(.A1(new_n11892_), .A2(new_n11901_), .A3(new_n11829_), .ZN(new_n11918_));
  AOI21_X1   g11627(.A1(new_n11917_), .A2(new_n11918_), .B(new_n11910_), .ZN(new_n11919_));
  NOR3_X1    g11628(.A1(new_n11914_), .A2(new_n11916_), .A3(new_n11919_), .ZN(new_n11920_));
  OAI21_X1   g11629(.A1(new_n11913_), .A2(new_n11920_), .B(new_n11489_), .ZN(new_n11921_));
  OAI21_X1   g11630(.A1(new_n11914_), .A2(new_n11916_), .B(new_n11919_), .ZN(new_n11922_));
  NAND3_X1   g11631(.A1(new_n11828_), .A2(new_n11826_), .A3(new_n11912_), .ZN(new_n11923_));
  NAND3_X1   g11632(.A1(new_n11923_), .A2(new_n11922_), .A3(new_n11501_), .ZN(new_n11924_));
  OAI22_X1   g11633(.A1(new_n5993_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n5991_), .ZN(new_n11925_));
  OAI21_X1   g11634(.A1(new_n1109_), .A2(new_n5997_), .B(new_n11925_), .ZN(new_n11926_));
  AOI21_X1   g11635(.A1(new_n11926_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n11927_));
  XOR2_X1    g11636(.A1(new_n1299_), .A2(new_n11927_), .Z(new_n11928_));
  INV_X1     g11637(.I(new_n11928_), .ZN(new_n11929_));
  NAND3_X1   g11638(.A1(new_n11921_), .A2(new_n11924_), .A3(new_n11929_), .ZN(new_n11930_));
  AOI21_X1   g11639(.A1(new_n11923_), .A2(new_n11922_), .B(new_n11501_), .ZN(new_n11931_));
  NOR3_X1    g11640(.A1(new_n11913_), .A2(new_n11920_), .A3(new_n11489_), .ZN(new_n11932_));
  OAI21_X1   g11641(.A1(new_n11931_), .A2(new_n11932_), .B(new_n11928_), .ZN(new_n11933_));
  OAI21_X1   g11642(.A1(new_n11517_), .A2(new_n11513_), .B(new_n11528_), .ZN(new_n11934_));
  NAND3_X1   g11643(.A1(new_n11934_), .A2(new_n11930_), .A3(new_n11933_), .ZN(new_n11935_));
  NAND2_X1   g11644(.A1(new_n11933_), .A2(new_n11930_), .ZN(new_n11936_));
  AOI21_X1   g11645(.A1(new_n11388_), .A2(new_n11529_), .B(new_n11509_), .ZN(new_n11937_));
  NAND2_X1   g11646(.A1(new_n11936_), .A2(new_n11937_), .ZN(new_n11938_));
  OAI22_X1   g11647(.A1(new_n5420_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n5107_), .ZN(new_n11939_));
  OAI21_X1   g11648(.A1(new_n1518_), .A2(new_n5112_), .B(new_n11939_), .ZN(new_n11940_));
  AOI21_X1   g11649(.A1(new_n11940_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n11941_));
  XNOR2_X1   g11650(.A1(new_n1638_), .A2(new_n11941_), .ZN(new_n11942_));
  AOI21_X1   g11651(.A1(new_n11938_), .A2(new_n11935_), .B(new_n11942_), .ZN(new_n11943_));
  NOR2_X1    g11652(.A1(new_n11936_), .A2(new_n11937_), .ZN(new_n11944_));
  AOI21_X1   g11653(.A1(new_n11930_), .A2(new_n11933_), .B(new_n11934_), .ZN(new_n11945_));
  INV_X1     g11654(.I(new_n11942_), .ZN(new_n11946_));
  NOR3_X1    g11655(.A1(new_n11944_), .A2(new_n11945_), .A3(new_n11946_), .ZN(new_n11947_));
  OAI22_X1   g11656(.A1(new_n11823_), .A2(new_n11526_), .B1(new_n11943_), .B2(new_n11947_), .ZN(new_n11948_));
  AOI21_X1   g11657(.A1(new_n11536_), .A2(new_n11547_), .B(new_n11526_), .ZN(new_n11949_));
  NAND3_X1   g11658(.A1(new_n11938_), .A2(new_n11935_), .A3(new_n11946_), .ZN(new_n11950_));
  OAI21_X1   g11659(.A1(new_n11944_), .A2(new_n11945_), .B(new_n11942_), .ZN(new_n11951_));
  NAND2_X1   g11660(.A1(new_n11951_), .A2(new_n11950_), .ZN(new_n11952_));
  NAND2_X1   g11661(.A1(new_n11949_), .A2(new_n11952_), .ZN(new_n11953_));
  OAI22_X1   g11662(.A1(new_n4072_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n4067_), .ZN(new_n11954_));
  OAI21_X1   g11663(.A1(new_n1803_), .A2(new_n4318_), .B(new_n11954_), .ZN(new_n11955_));
  AOI21_X1   g11664(.A1(new_n11955_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n11956_));
  XOR2_X1    g11665(.A1(new_n2106_), .A2(new_n11956_), .Z(new_n11957_));
  AOI21_X1   g11666(.A1(new_n11948_), .A2(new_n11953_), .B(new_n11957_), .ZN(new_n11958_));
  OAI21_X1   g11667(.A1(new_n11559_), .A2(new_n11556_), .B(new_n11958_), .ZN(new_n11959_));
  NOR2_X1    g11668(.A1(new_n11947_), .A2(new_n11943_), .ZN(new_n11960_));
  NOR2_X1    g11669(.A1(new_n11949_), .A2(new_n11960_), .ZN(new_n11961_));
  OAI21_X1   g11670(.A1(new_n11383_), .A2(new_n11533_), .B(new_n11546_), .ZN(new_n11962_));
  NOR3_X1    g11671(.A1(new_n11944_), .A2(new_n11945_), .A3(new_n11942_), .ZN(new_n11963_));
  AOI21_X1   g11672(.A1(new_n11938_), .A2(new_n11935_), .B(new_n11946_), .ZN(new_n11964_));
  NOR2_X1    g11673(.A1(new_n11963_), .A2(new_n11964_), .ZN(new_n11965_));
  NOR2_X1    g11674(.A1(new_n11962_), .A2(new_n11965_), .ZN(new_n11966_));
  INV_X1     g11675(.I(new_n11957_), .ZN(new_n11967_));
  OAI21_X1   g11676(.A1(new_n11966_), .A2(new_n11961_), .B(new_n11967_), .ZN(new_n11968_));
  NAND3_X1   g11677(.A1(new_n11968_), .A2(new_n11562_), .A3(new_n11382_), .ZN(new_n11969_));
  AOI21_X1   g11678(.A1(new_n11959_), .A2(new_n11969_), .B(new_n11822_), .ZN(new_n11970_));
  AOI21_X1   g11679(.A1(new_n11382_), .A2(new_n11562_), .B(new_n11968_), .ZN(new_n11971_));
  NOR3_X1    g11680(.A1(new_n11958_), .A2(new_n11556_), .A3(new_n11559_), .ZN(new_n11972_));
  NOR3_X1    g11681(.A1(new_n11971_), .A2(new_n11972_), .A3(new_n11821_), .ZN(new_n11973_));
  NOR2_X1    g11682(.A1(new_n11970_), .A2(new_n11973_), .ZN(new_n11974_));
  AOI22_X1   g11683(.A1(new_n3346_), .A2(\b[26] ), .B1(\b[27] ), .B2(new_n3351_), .ZN(new_n11975_));
  AOI21_X1   g11684(.A1(\b[25] ), .A2(new_n4331_), .B(new_n11975_), .ZN(new_n11976_));
  OAI21_X1   g11685(.A1(new_n11976_), .A2(\a[32] ), .B(new_n3346_), .ZN(new_n11977_));
  XOR2_X1    g11686(.A1(new_n2647_), .A2(new_n11977_), .Z(new_n11978_));
  NOR3_X1    g11687(.A1(new_n11974_), .A2(new_n11820_), .A3(new_n11978_), .ZN(new_n11979_));
  INV_X1     g11688(.I(new_n11820_), .ZN(new_n11980_));
  NOR2_X1    g11689(.A1(new_n11974_), .A2(new_n11978_), .ZN(new_n11981_));
  NOR2_X1    g11690(.A1(new_n11981_), .A2(new_n11980_), .ZN(new_n11982_));
  OAI21_X1   g11691(.A1(new_n11982_), .A2(new_n11979_), .B(new_n11819_), .ZN(new_n11983_));
  INV_X1     g11692(.I(new_n11983_), .ZN(new_n11984_));
  NOR3_X1    g11693(.A1(new_n11982_), .A2(new_n11819_), .A3(new_n11979_), .ZN(new_n11985_));
  OAI22_X1   g11694(.A1(new_n3018_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n3260_), .ZN(new_n11986_));
  OAI21_X1   g11695(.A1(new_n2842_), .A2(new_n2884_), .B(new_n11986_), .ZN(new_n11987_));
  AOI21_X1   g11696(.A1(new_n11987_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n11988_));
  XNOR2_X1   g11697(.A1(new_n3264_), .A2(new_n11988_), .ZN(new_n11989_));
  INV_X1     g11698(.I(new_n11989_), .ZN(new_n11990_));
  OAI21_X1   g11699(.A1(new_n11984_), .A2(new_n11985_), .B(new_n11990_), .ZN(new_n11991_));
  INV_X1     g11700(.I(new_n11991_), .ZN(new_n11992_));
  NAND2_X1   g11701(.A1(new_n11813_), .A2(new_n11992_), .ZN(new_n11993_));
  OAI21_X1   g11702(.A1(new_n11588_), .A2(new_n11585_), .B(new_n11160_), .ZN(new_n11994_));
  AOI21_X1   g11703(.A1(new_n11994_), .A2(new_n11163_), .B(new_n11161_), .ZN(new_n11995_));
  NAND2_X1   g11704(.A1(new_n11995_), .A2(new_n11991_), .ZN(new_n11996_));
  AOI21_X1   g11705(.A1(new_n11996_), .A2(new_n11993_), .B(new_n11811_), .ZN(new_n11997_));
  INV_X1     g11706(.I(new_n11810_), .ZN(new_n11998_));
  OAI21_X1   g11707(.A1(new_n11998_), .A2(new_n11808_), .B(new_n11578_), .ZN(new_n11999_));
  NOR2_X1    g11708(.A1(new_n11995_), .A2(new_n11991_), .ZN(new_n12000_));
  NOR2_X1    g11709(.A1(new_n11813_), .A2(new_n11992_), .ZN(new_n12001_));
  NOR3_X1    g11710(.A1(new_n12000_), .A2(new_n12001_), .A3(new_n11999_), .ZN(new_n12002_));
  OAI22_X1   g11711(.A1(new_n2171_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n2166_), .ZN(new_n12003_));
  OAI21_X1   g11712(.A1(new_n3709_), .A2(new_n2322_), .B(new_n12003_), .ZN(new_n12004_));
  AOI21_X1   g11713(.A1(new_n12004_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n12005_));
  XNOR2_X1   g11714(.A1(new_n3993_), .A2(new_n12005_), .ZN(new_n12006_));
  INV_X1     g11715(.I(new_n12006_), .ZN(new_n12007_));
  OAI21_X1   g11716(.A1(new_n11997_), .A2(new_n12002_), .B(new_n12007_), .ZN(new_n12008_));
  NOR2_X1    g11717(.A1(new_n11802_), .A2(new_n12008_), .ZN(new_n12009_));
  AOI21_X1   g11718(.A1(new_n11600_), .A2(new_n11603_), .B(new_n11375_), .ZN(new_n12010_));
  OAI21_X1   g11719(.A1(new_n12010_), .A2(new_n11166_), .B(new_n10917_), .ZN(new_n12011_));
  OAI21_X1   g11720(.A1(new_n12000_), .A2(new_n12001_), .B(new_n11999_), .ZN(new_n12012_));
  NAND3_X1   g11721(.A1(new_n11996_), .A2(new_n11993_), .A3(new_n11811_), .ZN(new_n12013_));
  AOI21_X1   g11722(.A1(new_n12012_), .A2(new_n12013_), .B(new_n12006_), .ZN(new_n12014_));
  NOR2_X1    g11723(.A1(new_n12011_), .A2(new_n12014_), .ZN(new_n12015_));
  OAI21_X1   g11724(.A1(new_n12009_), .A2(new_n12015_), .B(new_n11800_), .ZN(new_n12016_));
  NAND2_X1   g11725(.A1(new_n12011_), .A2(new_n12014_), .ZN(new_n12017_));
  NAND2_X1   g11726(.A1(new_n11802_), .A2(new_n12008_), .ZN(new_n12018_));
  NAND3_X1   g11727(.A1(new_n12018_), .A2(new_n12017_), .A3(new_n11799_), .ZN(new_n12019_));
  OAI22_X1   g11728(.A1(new_n1712_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n1707_), .ZN(new_n12020_));
  OAI21_X1   g11729(.A1(new_n4253_), .A2(new_n1850_), .B(new_n12020_), .ZN(new_n12021_));
  AOI21_X1   g11730(.A1(new_n12021_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n12022_));
  XNOR2_X1   g11731(.A1(new_n4778_), .A2(new_n12022_), .ZN(new_n12023_));
  AOI21_X1   g11732(.A1(new_n12016_), .A2(new_n12019_), .B(new_n12023_), .ZN(new_n12024_));
  NAND2_X1   g11733(.A1(new_n11798_), .A2(new_n12024_), .ZN(new_n12025_));
  OAI21_X1   g11734(.A1(new_n11627_), .A2(new_n11628_), .B(new_n11626_), .ZN(new_n12026_));
  AOI21_X1   g11735(.A1(new_n12026_), .A2(new_n11208_), .B(new_n11194_), .ZN(new_n12027_));
  AOI21_X1   g11736(.A1(new_n12018_), .A2(new_n12017_), .B(new_n11799_), .ZN(new_n12028_));
  NOR3_X1    g11737(.A1(new_n12009_), .A2(new_n12015_), .A3(new_n11800_), .ZN(new_n12029_));
  INV_X1     g11738(.I(new_n12023_), .ZN(new_n12030_));
  OAI21_X1   g11739(.A1(new_n12028_), .A2(new_n12029_), .B(new_n12030_), .ZN(new_n12031_));
  NAND2_X1   g11740(.A1(new_n12027_), .A2(new_n12031_), .ZN(new_n12032_));
  AOI21_X1   g11741(.A1(new_n12032_), .A2(new_n12025_), .B(new_n11628_), .ZN(new_n12033_));
  NOR2_X1    g11742(.A1(new_n12027_), .A2(new_n12031_), .ZN(new_n12034_));
  NOR2_X1    g11743(.A1(new_n11798_), .A2(new_n12024_), .ZN(new_n12035_));
  NOR3_X1    g11744(.A1(new_n12034_), .A2(new_n12035_), .A3(new_n11621_), .ZN(new_n12036_));
  OAI22_X1   g11745(.A1(new_n1347_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n1344_), .ZN(new_n12037_));
  OAI21_X1   g11746(.A1(new_n5068_), .A2(new_n1457_), .B(new_n12037_), .ZN(new_n12038_));
  AOI21_X1   g11747(.A1(new_n12038_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n12039_));
  XNOR2_X1   g11748(.A1(new_n5600_), .A2(new_n12039_), .ZN(new_n12040_));
  INV_X1     g11749(.I(new_n12040_), .ZN(new_n12041_));
  OAI21_X1   g11750(.A1(new_n12033_), .A2(new_n12036_), .B(new_n12041_), .ZN(new_n12042_));
  NOR2_X1    g11751(.A1(new_n11796_), .A2(new_n12042_), .ZN(new_n12043_));
  AOI21_X1   g11752(.A1(new_n11639_), .A2(new_n11636_), .B(new_n11368_), .ZN(new_n12044_));
  OAI21_X1   g11753(.A1(new_n12044_), .A2(new_n11199_), .B(new_n11221_), .ZN(new_n12045_));
  OAI21_X1   g11754(.A1(new_n12034_), .A2(new_n12035_), .B(new_n11621_), .ZN(new_n12046_));
  NAND3_X1   g11755(.A1(new_n12032_), .A2(new_n12025_), .A3(new_n11628_), .ZN(new_n12047_));
  AOI21_X1   g11756(.A1(new_n12046_), .A2(new_n12047_), .B(new_n12040_), .ZN(new_n12048_));
  NOR2_X1    g11757(.A1(new_n12048_), .A2(new_n12045_), .ZN(new_n12049_));
  OAI21_X1   g11758(.A1(new_n12043_), .A2(new_n12049_), .B(new_n11639_), .ZN(new_n12050_));
  NAND2_X1   g11759(.A1(new_n12048_), .A2(new_n12045_), .ZN(new_n12051_));
  NAND2_X1   g11760(.A1(new_n11796_), .A2(new_n12042_), .ZN(new_n12052_));
  NAND3_X1   g11761(.A1(new_n12052_), .A2(new_n12051_), .A3(new_n11646_), .ZN(new_n12053_));
  OAI22_X1   g11762(.A1(new_n1055_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n1061_), .ZN(new_n12054_));
  OAI21_X1   g11763(.A1(new_n5921_), .A2(new_n1332_), .B(new_n12054_), .ZN(new_n12055_));
  AOI21_X1   g11764(.A1(new_n12055_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n12056_));
  XOR2_X1    g11765(.A1(new_n6543_), .A2(new_n12056_), .Z(new_n12057_));
  AOI21_X1   g11766(.A1(new_n12050_), .A2(new_n12053_), .B(new_n12057_), .ZN(new_n12058_));
  NAND2_X1   g11767(.A1(new_n11794_), .A2(new_n12058_), .ZN(new_n12059_));
  OAI21_X1   g11768(.A1(new_n11662_), .A2(new_n11663_), .B(new_n11661_), .ZN(new_n12060_));
  AOI21_X1   g11769(.A1(new_n12060_), .A2(new_n11224_), .B(new_n11363_), .ZN(new_n12061_));
  INV_X1     g11770(.I(new_n12058_), .ZN(new_n12062_));
  NAND2_X1   g11771(.A1(new_n12062_), .A2(new_n12061_), .ZN(new_n12063_));
  AOI21_X1   g11772(.A1(new_n12063_), .A2(new_n12059_), .B(new_n11663_), .ZN(new_n12064_));
  NOR2_X1    g11773(.A1(new_n12062_), .A2(new_n12061_), .ZN(new_n12065_));
  NOR2_X1    g11774(.A1(new_n11794_), .A2(new_n12058_), .ZN(new_n12066_));
  NOR3_X1    g11775(.A1(new_n12065_), .A2(new_n12066_), .A3(new_n11657_), .ZN(new_n12067_));
  OAI22_X1   g11776(.A1(new_n970_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n820_), .ZN(new_n12068_));
  OAI21_X1   g11777(.A1(new_n6847_), .A2(new_n894_), .B(new_n12068_), .ZN(new_n12069_));
  AOI21_X1   g11778(.A1(new_n12069_), .A2(new_n827_), .B(new_n970_), .ZN(new_n12070_));
  XOR2_X1    g11779(.A1(new_n7516_), .A2(new_n12070_), .Z(new_n12071_));
  INV_X1     g11780(.I(new_n12071_), .ZN(new_n12072_));
  OAI21_X1   g11781(.A1(new_n12067_), .A2(new_n12064_), .B(new_n12072_), .ZN(new_n12073_));
  NOR2_X1    g11782(.A1(new_n11792_), .A2(new_n12073_), .ZN(new_n12074_));
  NAND2_X1   g11783(.A1(new_n11773_), .A2(new_n11790_), .ZN(new_n12075_));
  OAI21_X1   g11784(.A1(new_n12065_), .A2(new_n12066_), .B(new_n11657_), .ZN(new_n12076_));
  NAND3_X1   g11785(.A1(new_n12063_), .A2(new_n12059_), .A3(new_n11663_), .ZN(new_n12077_));
  AOI21_X1   g11786(.A1(new_n12076_), .A2(new_n12077_), .B(new_n12071_), .ZN(new_n12078_));
  NOR2_X1    g11787(.A1(new_n12078_), .A2(new_n12075_), .ZN(new_n12079_));
  OAI21_X1   g11788(.A1(new_n12074_), .A2(new_n12079_), .B(new_n11784_), .ZN(new_n12080_));
  INV_X1     g11789(.I(new_n11784_), .ZN(new_n12081_));
  NAND2_X1   g11790(.A1(new_n12078_), .A2(new_n12075_), .ZN(new_n12082_));
  NAND2_X1   g11791(.A1(new_n11792_), .A2(new_n12073_), .ZN(new_n12083_));
  NAND3_X1   g11792(.A1(new_n12083_), .A2(new_n12082_), .A3(new_n12081_), .ZN(new_n12084_));
  OAI22_X1   g11793(.A1(new_n607_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n610_), .ZN(new_n12085_));
  OAI21_X1   g11794(.A1(new_n7870_), .A2(new_n684_), .B(new_n12085_), .ZN(new_n12086_));
  AOI21_X1   g11795(.A1(new_n12086_), .A2(new_n612_), .B(new_n607_), .ZN(new_n12087_));
  XOR2_X1    g11796(.A1(new_n8568_), .A2(new_n12087_), .Z(new_n12088_));
  AOI21_X1   g11797(.A1(new_n12080_), .A2(new_n12084_), .B(new_n12088_), .ZN(new_n12089_));
  OAI21_X1   g11798(.A1(new_n11781_), .A2(new_n11783_), .B(new_n12089_), .ZN(new_n12090_));
  OR3_X2     g11799(.A1(new_n11781_), .A2(new_n11783_), .A3(new_n12089_), .Z(new_n12091_));
  AOI21_X1   g11800(.A1(new_n12091_), .A2(new_n12090_), .B(new_n11779_), .ZN(new_n12092_));
  INV_X1     g11801(.I(new_n12090_), .ZN(new_n12093_));
  OAI21_X1   g11802(.A1(new_n11686_), .A2(new_n11683_), .B(new_n11252_), .ZN(new_n12094_));
  NAND2_X1   g11803(.A1(new_n12094_), .A2(new_n11689_), .ZN(new_n12095_));
  NAND3_X1   g11804(.A1(new_n12095_), .A2(new_n11251_), .A3(new_n11782_), .ZN(new_n12096_));
  NOR2_X1    g11805(.A1(new_n12096_), .A2(new_n12089_), .ZN(new_n12097_));
  NOR3_X1    g11806(.A1(new_n12097_), .A2(new_n12093_), .A3(new_n11778_), .ZN(new_n12098_));
  OAI22_X1   g11807(.A1(new_n448_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n450_), .ZN(new_n12099_));
  OAI21_X1   g11808(.A1(new_n8948_), .A2(new_n496_), .B(new_n12099_), .ZN(new_n12100_));
  AOI21_X1   g11809(.A1(new_n12100_), .A2(new_n452_), .B(new_n448_), .ZN(new_n12101_));
  XNOR2_X1   g11810(.A1(new_n9642_), .A2(new_n12101_), .ZN(new_n12102_));
  INV_X1     g11811(.I(new_n12102_), .ZN(new_n12103_));
  OAI21_X1   g11812(.A1(new_n12098_), .A2(new_n12092_), .B(new_n12103_), .ZN(new_n12104_));
  AOI21_X1   g11813(.A1(new_n11772_), .A2(new_n11770_), .B(new_n12104_), .ZN(new_n12105_));
  AOI21_X1   g11814(.A1(new_n11708_), .A2(new_n11766_), .B(new_n11262_), .ZN(new_n12106_));
  NAND3_X1   g11815(.A1(new_n11707_), .A2(new_n11704_), .A3(new_n11709_), .ZN(new_n12107_));
  NAND2_X1   g11816(.A1(new_n12107_), .A2(new_n11356_), .ZN(new_n12108_));
  OAI21_X1   g11817(.A1(new_n12097_), .A2(new_n12093_), .B(new_n11778_), .ZN(new_n12109_));
  NAND3_X1   g11818(.A1(new_n12091_), .A2(new_n11779_), .A3(new_n12090_), .ZN(new_n12110_));
  AOI21_X1   g11819(.A1(new_n12109_), .A2(new_n12110_), .B(new_n12102_), .ZN(new_n12111_));
  NOR3_X1    g11820(.A1(new_n12106_), .A2(new_n12108_), .A3(new_n12111_), .ZN(new_n12112_));
  OAI21_X1   g11821(.A1(new_n12105_), .A2(new_n12112_), .B(new_n11707_), .ZN(new_n12113_));
  OAI21_X1   g11822(.A1(new_n12106_), .A2(new_n12108_), .B(new_n12111_), .ZN(new_n12114_));
  NAND3_X1   g11823(.A1(new_n11772_), .A2(new_n11770_), .A3(new_n12104_), .ZN(new_n12115_));
  NAND3_X1   g11824(.A1(new_n12115_), .A2(new_n12114_), .A3(new_n11768_), .ZN(new_n12116_));
  OAI22_X1   g11825(.A1(new_n10477_), .A2(new_n341_), .B1(new_n404_), .B2(new_n10862_), .ZN(new_n12117_));
  OAI21_X1   g11826(.A1(new_n10031_), .A2(new_n366_), .B(new_n12117_), .ZN(new_n12118_));
  AOI21_X1   g11827(.A1(new_n12118_), .A2(new_n334_), .B(new_n341_), .ZN(new_n12119_));
  XNOR2_X1   g11828(.A1(new_n10866_), .A2(new_n12119_), .ZN(new_n12120_));
  INV_X1     g11829(.I(new_n12120_), .ZN(new_n12121_));
  NAND3_X1   g11830(.A1(new_n12113_), .A2(new_n12116_), .A3(new_n12121_), .ZN(new_n12122_));
  AOI21_X1   g11831(.A1(new_n12115_), .A2(new_n12114_), .B(new_n11768_), .ZN(new_n12123_));
  NOR3_X1    g11832(.A1(new_n12105_), .A2(new_n12112_), .A3(new_n11707_), .ZN(new_n12124_));
  OAI21_X1   g11833(.A1(new_n12123_), .A2(new_n12124_), .B(new_n12120_), .ZN(new_n12125_));
  XNOR2_X1   g11834(.A1(\b[55] ), .A2(\b[57] ), .ZN(new_n12126_));
  NOR2_X1    g11835(.A1(new_n12126_), .A2(new_n11743_), .ZN(new_n12127_));
  XNOR2_X1   g11836(.A1(new_n11742_), .A2(new_n12127_), .ZN(new_n12128_));
  NAND2_X1   g11837(.A1(new_n286_), .A2(\b[56] ), .ZN(new_n12129_));
  AOI22_X1   g11838(.A1(new_n304_), .A2(\b[55] ), .B1(new_n262_), .B2(\b[57] ), .ZN(new_n12130_));
  AOI21_X1   g11839(.A1(new_n12129_), .A2(new_n12130_), .B(new_n426_), .ZN(new_n12131_));
  NAND2_X1   g11840(.A1(new_n12128_), .A2(new_n12131_), .ZN(new_n12132_));
  XOR2_X1    g11841(.A1(new_n12132_), .A2(\a[2] ), .Z(new_n12133_));
  AOI21_X1   g11842(.A1(new_n12125_), .A2(new_n12122_), .B(new_n12133_), .ZN(new_n12134_));
  NOR3_X1    g11843(.A1(new_n12123_), .A2(new_n12124_), .A3(new_n12120_), .ZN(new_n12135_));
  AOI21_X1   g11844(.A1(new_n12113_), .A2(new_n12116_), .B(new_n12121_), .ZN(new_n12136_));
  INV_X1     g11845(.I(new_n12133_), .ZN(new_n12137_));
  NOR3_X1    g11846(.A1(new_n12135_), .A2(new_n12136_), .A3(new_n12137_), .ZN(new_n12138_));
  OAI21_X1   g11847(.A1(new_n12138_), .A2(new_n12134_), .B(new_n11765_), .ZN(new_n12139_));
  AOI21_X1   g11848(.A1(new_n11728_), .A2(new_n11716_), .B(new_n11352_), .ZN(new_n12140_));
  AOI21_X1   g11849(.A1(new_n11762_), .A2(new_n11763_), .B(new_n12140_), .ZN(new_n12141_));
  NOR3_X1    g11850(.A1(new_n12135_), .A2(new_n12136_), .A3(new_n12133_), .ZN(new_n12142_));
  AOI21_X1   g11851(.A1(new_n12125_), .A2(new_n12122_), .B(new_n12137_), .ZN(new_n12143_));
  OAI21_X1   g11852(.A1(new_n12142_), .A2(new_n12143_), .B(new_n12141_), .ZN(new_n12144_));
  AOI21_X1   g11853(.A1(new_n12139_), .A2(new_n12144_), .B(new_n11759_), .ZN(new_n12145_));
  XNOR2_X1   g11854(.A1(new_n12145_), .A2(new_n11754_), .ZN(new_n12146_));
  XOR2_X1    g11855(.A1(new_n12146_), .A2(new_n11347_), .Z(\f[57] ));
  NOR2_X1    g11856(.A1(new_n12135_), .A2(new_n12136_), .ZN(new_n12148_));
  AOI21_X1   g11857(.A1(new_n12113_), .A2(new_n12116_), .B(new_n12120_), .ZN(new_n12149_));
  NOR2_X1    g11858(.A1(new_n12106_), .A2(new_n12108_), .ZN(new_n12150_));
  NAND2_X1   g11859(.A1(new_n12109_), .A2(new_n12110_), .ZN(new_n12151_));
  NOR2_X1    g11860(.A1(new_n12098_), .A2(new_n12092_), .ZN(new_n12152_));
  AOI21_X1   g11861(.A1(new_n12152_), .A2(new_n11707_), .B(new_n12102_), .ZN(new_n12153_));
  AOI22_X1   g11862(.A1(new_n12150_), .A2(new_n12153_), .B1(new_n11768_), .B2(new_n12151_), .ZN(new_n12154_));
  AOI21_X1   g11863(.A1(new_n12076_), .A2(new_n12077_), .B(new_n11784_), .ZN(new_n12155_));
  NAND3_X1   g11864(.A1(new_n12076_), .A2(new_n12077_), .A3(new_n11784_), .ZN(new_n12156_));
  NOR3_X1    g11865(.A1(new_n11791_), .A2(new_n11785_), .A3(new_n12071_), .ZN(new_n12157_));
  AOI21_X1   g11866(.A1(new_n12157_), .A2(new_n12156_), .B(new_n12155_), .ZN(new_n12158_));
  AOI21_X1   g11867(.A1(new_n12052_), .A2(new_n12051_), .B(new_n11646_), .ZN(new_n12159_));
  NOR3_X1    g11868(.A1(new_n12043_), .A2(new_n12049_), .A3(new_n11639_), .ZN(new_n12160_));
  NOR2_X1    g11869(.A1(new_n12159_), .A2(new_n12160_), .ZN(new_n12161_));
  NAND2_X1   g11870(.A1(new_n12050_), .A2(new_n12053_), .ZN(new_n12162_));
  INV_X1     g11871(.I(new_n12057_), .ZN(new_n12163_));
  OAI21_X1   g11872(.A1(new_n12162_), .A2(new_n11663_), .B(new_n12163_), .ZN(new_n12164_));
  OAI22_X1   g11873(.A1(new_n12164_), .A2(new_n11794_), .B1(new_n11657_), .B2(new_n12161_), .ZN(new_n12165_));
  OAI22_X1   g11874(.A1(new_n1347_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n1344_), .ZN(new_n12166_));
  OAI21_X1   g11875(.A1(new_n5353_), .A2(new_n1457_), .B(new_n12166_), .ZN(new_n12167_));
  AOI21_X1   g11876(.A1(new_n12167_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n12168_));
  XOR2_X1    g11877(.A1(new_n5926_), .A2(new_n12168_), .Z(new_n12169_));
  INV_X1     g11878(.I(new_n12169_), .ZN(new_n12170_));
  NOR2_X1    g11879(.A1(new_n12028_), .A2(new_n12029_), .ZN(new_n12171_));
  INV_X1     g11880(.I(new_n12171_), .ZN(new_n12172_));
  AOI21_X1   g11881(.A1(new_n12171_), .A2(new_n11621_), .B(new_n12023_), .ZN(new_n12173_));
  AOI22_X1   g11882(.A1(new_n12173_), .A2(new_n12027_), .B1(new_n11628_), .B2(new_n12172_), .ZN(new_n12174_));
  AOI21_X1   g11883(.A1(new_n12046_), .A2(new_n12047_), .B(new_n11639_), .ZN(new_n12175_));
  NOR3_X1    g11884(.A1(new_n12033_), .A2(new_n12036_), .A3(new_n11646_), .ZN(new_n12176_));
  NOR3_X1    g11885(.A1(new_n12176_), .A2(new_n12045_), .A3(new_n12040_), .ZN(new_n12177_));
  AOI21_X1   g11886(.A1(new_n11815_), .A2(new_n11816_), .B(new_n11379_), .ZN(new_n12178_));
  NOR3_X1    g11887(.A1(new_n11563_), .A2(new_n11557_), .A3(new_n11380_), .ZN(new_n12179_));
  NOR2_X1    g11888(.A1(new_n12178_), .A2(new_n12179_), .ZN(new_n12180_));
  NOR4_X1    g11889(.A1(new_n11974_), .A2(new_n11569_), .A3(new_n11565_), .A4(new_n12180_), .ZN(new_n12181_));
  NAND2_X1   g11890(.A1(new_n11819_), .A2(new_n11974_), .ZN(new_n12182_));
  NOR2_X1    g11891(.A1(new_n11980_), .A2(new_n11978_), .ZN(new_n12183_));
  AOI21_X1   g11892(.A1(new_n12182_), .A2(new_n12183_), .B(new_n12181_), .ZN(new_n12184_));
  AOI21_X1   g11893(.A1(new_n11921_), .A2(new_n11924_), .B(new_n11929_), .ZN(new_n12185_));
  NAND3_X1   g11894(.A1(new_n11937_), .A2(new_n11930_), .A3(new_n11933_), .ZN(new_n12186_));
  NAND2_X1   g11895(.A1(new_n11917_), .A2(new_n11918_), .ZN(new_n12187_));
  NAND2_X1   g11896(.A1(new_n12187_), .A2(new_n11501_), .ZN(new_n12188_));
  INV_X1     g11897(.I(new_n12188_), .ZN(new_n12189_));
  NAND3_X1   g11898(.A1(new_n11917_), .A2(new_n11918_), .A3(new_n11489_), .ZN(new_n12190_));
  NAND2_X1   g11899(.A1(new_n12190_), .A2(new_n11911_), .ZN(new_n12191_));
  NOR3_X1    g11900(.A1(new_n12191_), .A2(new_n11914_), .A3(new_n11916_), .ZN(new_n12192_));
  NAND2_X1   g11901(.A1(new_n11883_), .A2(new_n11886_), .ZN(new_n12193_));
  NAND2_X1   g11902(.A1(new_n12193_), .A2(new_n11829_), .ZN(new_n12194_));
  INV_X1     g11903(.I(new_n12194_), .ZN(new_n12195_));
  NAND2_X1   g11904(.A1(new_n11896_), .A2(new_n11894_), .ZN(new_n12196_));
  OAI21_X1   g11905(.A1(new_n12193_), .A2(new_n11829_), .B(new_n11899_), .ZN(new_n12197_));
  NOR2_X1    g11906(.A1(new_n12196_), .A2(new_n12197_), .ZN(new_n12198_));
  OAI21_X1   g11907(.A1(new_n11868_), .A2(new_n11864_), .B(new_n11833_), .ZN(new_n12199_));
  INV_X1     g11908(.I(new_n12199_), .ZN(new_n12200_));
  NAND2_X1   g11909(.A1(new_n11836_), .A2(new_n11835_), .ZN(new_n12201_));
  NOR3_X1    g11910(.A1(new_n11868_), .A2(new_n11864_), .A3(new_n11833_), .ZN(new_n12202_));
  NOR3_X1    g11911(.A1(new_n12201_), .A2(new_n11872_), .A3(new_n12202_), .ZN(new_n12203_));
  NAND2_X1   g11912(.A1(new_n11863_), .A2(new_n11878_), .ZN(new_n12204_));
  NAND2_X1   g11913(.A1(new_n11851_), .A2(new_n11843_), .ZN(new_n12205_));
  NOR2_X1    g11914(.A1(new_n11850_), .A2(new_n258_), .ZN(new_n12206_));
  OAI21_X1   g11915(.A1(new_n11851_), .A2(new_n11843_), .B(new_n12206_), .ZN(new_n12207_));
  NAND2_X1   g11916(.A1(new_n12207_), .A2(new_n12205_), .ZN(new_n12208_));
  AOI22_X1   g11917(.A1(new_n10969_), .A2(new_n10957_), .B1(new_n11394_), .B2(\b[2] ), .ZN(new_n12209_));
  OAI21_X1   g11918(.A1(new_n12209_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n12210_));
  XOR2_X1    g11919(.A1(new_n12210_), .A2(new_n329_), .Z(new_n12211_));
  INV_X1     g11920(.I(new_n12211_), .ZN(new_n12212_));
  XNOR2_X1   g11921(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n12213_));
  NOR2_X1    g11922(.A1(new_n11842_), .A2(new_n12213_), .ZN(new_n12214_));
  NAND2_X1   g11923(.A1(new_n11840_), .A2(\a[58] ), .ZN(new_n12215_));
  OAI21_X1   g11924(.A1(\a[58] ), .A2(new_n11839_), .B(new_n12215_), .ZN(new_n12216_));
  XNOR2_X1   g11925(.A1(\a[58] ), .A2(\a[59] ), .ZN(new_n12217_));
  NAND3_X1   g11926(.A1(new_n12216_), .A2(new_n11850_), .A3(new_n12217_), .ZN(new_n12218_));
  NOR2_X1    g11927(.A1(new_n319_), .A2(\a[59] ), .ZN(new_n12219_));
  NAND2_X1   g11928(.A1(new_n12218_), .A2(new_n12219_), .ZN(new_n12220_));
  AOI21_X1   g11929(.A1(new_n12220_), .A2(new_n12214_), .B(new_n444_), .ZN(new_n12221_));
  INV_X1     g11930(.I(\a[59] ), .ZN(new_n12222_));
  NOR2_X1    g11931(.A1(new_n11839_), .A2(\a[58] ), .ZN(new_n12223_));
  AOI21_X1   g11932(.A1(\a[58] ), .A2(new_n11840_), .B(new_n12223_), .ZN(new_n12224_));
  NAND2_X1   g11933(.A1(new_n11850_), .A2(new_n12217_), .ZN(new_n12225_));
  NOR2_X1    g11934(.A1(new_n12225_), .A2(new_n12224_), .ZN(new_n12226_));
  INV_X1     g11935(.I(new_n12219_), .ZN(new_n12227_));
  OAI21_X1   g11936(.A1(new_n12226_), .A2(new_n12227_), .B(new_n12214_), .ZN(new_n12228_));
  OAI21_X1   g11937(.A1(new_n12228_), .A2(new_n271_), .B(new_n12222_), .ZN(new_n12229_));
  NOR2_X1    g11938(.A1(new_n12229_), .A2(new_n12221_), .ZN(new_n12230_));
  INV_X1     g11939(.I(new_n12230_), .ZN(new_n12231_));
  NAND3_X1   g11940(.A1(new_n12231_), .A2(\b[0] ), .A3(new_n11850_), .ZN(new_n12232_));
  OAI21_X1   g11941(.A1(new_n12230_), .A2(new_n258_), .B(new_n11842_), .ZN(new_n12233_));
  NAND2_X1   g11942(.A1(new_n12232_), .A2(new_n12233_), .ZN(new_n12234_));
  NAND2_X1   g11943(.A1(new_n12234_), .A2(new_n12212_), .ZN(new_n12235_));
  NAND3_X1   g11944(.A1(new_n12232_), .A2(new_n12211_), .A3(new_n12233_), .ZN(new_n12236_));
  NAND2_X1   g11945(.A1(new_n12235_), .A2(new_n12236_), .ZN(new_n12237_));
  NAND2_X1   g11946(.A1(new_n12237_), .A2(new_n12208_), .ZN(new_n12238_));
  NAND2_X1   g11947(.A1(new_n12234_), .A2(new_n12211_), .ZN(new_n12239_));
  NOR2_X1    g11948(.A1(new_n12234_), .A2(new_n12211_), .ZN(new_n12240_));
  INV_X1     g11949(.I(new_n12240_), .ZN(new_n12241_));
  AOI21_X1   g11950(.A1(new_n12241_), .A2(new_n12239_), .B(new_n12208_), .ZN(new_n12242_));
  INV_X1     g11951(.I(new_n12242_), .ZN(new_n12243_));
  NAND2_X1   g11952(.A1(new_n12243_), .A2(new_n12238_), .ZN(new_n12244_));
  OAI22_X1   g11953(.A1(new_n11411_), .A2(new_n509_), .B1(new_n419_), .B2(new_n10137_), .ZN(new_n12245_));
  AOI21_X1   g11954(.A1(new_n12245_), .A2(new_n9718_), .B(new_n9713_), .ZN(new_n12246_));
  XOR2_X1    g11955(.A1(new_n471_), .A2(new_n12246_), .Z(new_n12247_));
  INV_X1     g11956(.I(new_n12247_), .ZN(new_n12248_));
  NAND2_X1   g11957(.A1(new_n12244_), .A2(new_n12248_), .ZN(new_n12249_));
  NAND3_X1   g11958(.A1(new_n12243_), .A2(new_n12238_), .A3(new_n12247_), .ZN(new_n12250_));
  AOI22_X1   g11959(.A1(new_n12249_), .A2(new_n12250_), .B1(new_n12204_), .B2(new_n11861_), .ZN(new_n12251_));
  NAND2_X1   g11960(.A1(new_n12204_), .A2(new_n11861_), .ZN(new_n12252_));
  NAND3_X1   g11961(.A1(new_n12243_), .A2(new_n12238_), .A3(new_n12248_), .ZN(new_n12253_));
  INV_X1     g11962(.I(new_n12238_), .ZN(new_n12254_));
  OAI21_X1   g11963(.A1(new_n12254_), .A2(new_n12242_), .B(new_n12247_), .ZN(new_n12255_));
  AOI21_X1   g11964(.A1(new_n12253_), .A2(new_n12255_), .B(new_n12252_), .ZN(new_n12256_));
  NOR2_X1    g11965(.A1(new_n12256_), .A2(new_n12251_), .ZN(new_n12257_));
  OAI22_X1   g11966(.A1(new_n8644_), .A2(new_n565_), .B1(new_n656_), .B2(new_n9388_), .ZN(new_n12258_));
  OAI21_X1   g11967(.A1(new_n515_), .A2(new_n10154_), .B(new_n12258_), .ZN(new_n12259_));
  AOI21_X1   g11968(.A1(new_n12259_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n12260_));
  XNOR2_X1   g11969(.A1(new_n660_), .A2(new_n12260_), .ZN(new_n12261_));
  NOR2_X1    g11970(.A1(new_n12257_), .A2(new_n12261_), .ZN(new_n12262_));
  INV_X1     g11971(.I(new_n12261_), .ZN(new_n12263_));
  NOR3_X1    g11972(.A1(new_n12256_), .A2(new_n12251_), .A3(new_n12263_), .ZN(new_n12264_));
  OAI22_X1   g11973(.A1(new_n12262_), .A2(new_n12264_), .B1(new_n12200_), .B2(new_n12203_), .ZN(new_n12265_));
  NOR2_X1    g11974(.A1(new_n12203_), .A2(new_n12200_), .ZN(new_n12266_));
  INV_X1     g11975(.I(new_n12251_), .ZN(new_n12267_));
  NAND2_X1   g11976(.A1(new_n12253_), .A2(new_n12255_), .ZN(new_n12268_));
  NAND3_X1   g11977(.A1(new_n12268_), .A2(new_n11861_), .A3(new_n12204_), .ZN(new_n12269_));
  NAND3_X1   g11978(.A1(new_n12267_), .A2(new_n12269_), .A3(new_n12263_), .ZN(new_n12270_));
  OAI21_X1   g11979(.A1(new_n12256_), .A2(new_n12251_), .B(new_n12261_), .ZN(new_n12271_));
  NAND2_X1   g11980(.A1(new_n12270_), .A2(new_n12271_), .ZN(new_n12272_));
  NAND2_X1   g11981(.A1(new_n12272_), .A2(new_n12266_), .ZN(new_n12273_));
  OAI22_X1   g11982(.A1(new_n7619_), .A2(new_n780_), .B1(new_n861_), .B2(new_n8309_), .ZN(new_n12274_));
  OAI21_X1   g11983(.A1(new_n706_), .A2(new_n7947_), .B(new_n12274_), .ZN(new_n12275_));
  AOI21_X1   g11984(.A1(new_n12275_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n12276_));
  XNOR2_X1   g11985(.A1(new_n860_), .A2(new_n12276_), .ZN(new_n12277_));
  INV_X1     g11986(.I(new_n12277_), .ZN(new_n12278_));
  NAND3_X1   g11987(.A1(new_n12273_), .A2(new_n12265_), .A3(new_n12278_), .ZN(new_n12279_));
  NAND2_X1   g11988(.A1(new_n12267_), .A2(new_n12269_), .ZN(new_n12280_));
  NAND2_X1   g11989(.A1(new_n12280_), .A2(new_n12263_), .ZN(new_n12281_));
  INV_X1     g11990(.I(new_n12264_), .ZN(new_n12282_));
  AOI21_X1   g11991(.A1(new_n12281_), .A2(new_n12282_), .B(new_n12266_), .ZN(new_n12283_));
  INV_X1     g11992(.I(new_n12266_), .ZN(new_n12284_));
  NOR3_X1    g11993(.A1(new_n12256_), .A2(new_n12251_), .A3(new_n12261_), .ZN(new_n12285_));
  AOI21_X1   g11994(.A1(new_n12267_), .A2(new_n12269_), .B(new_n12263_), .ZN(new_n12286_));
  NOR2_X1    g11995(.A1(new_n12286_), .A2(new_n12285_), .ZN(new_n12287_));
  NOR2_X1    g11996(.A1(new_n12284_), .A2(new_n12287_), .ZN(new_n12288_));
  OAI21_X1   g11997(.A1(new_n12288_), .A2(new_n12283_), .B(new_n12277_), .ZN(new_n12289_));
  NAND2_X1   g11998(.A1(new_n12289_), .A2(new_n12279_), .ZN(new_n12290_));
  OAI21_X1   g11999(.A1(new_n12195_), .A2(new_n12198_), .B(new_n12290_), .ZN(new_n12291_));
  OR2_X2     g12000(.A1(new_n12196_), .A2(new_n12197_), .Z(new_n12292_));
  OAI21_X1   g12001(.A1(new_n12288_), .A2(new_n12283_), .B(new_n12278_), .ZN(new_n12293_));
  NAND3_X1   g12002(.A1(new_n12273_), .A2(new_n12265_), .A3(new_n12277_), .ZN(new_n12294_));
  NAND2_X1   g12003(.A1(new_n12293_), .A2(new_n12294_), .ZN(new_n12295_));
  NAND3_X1   g12004(.A1(new_n12295_), .A2(new_n12292_), .A3(new_n12194_), .ZN(new_n12296_));
  NAND2_X1   g12005(.A1(new_n12291_), .A2(new_n12296_), .ZN(new_n12297_));
  OAI22_X1   g12006(.A1(new_n6644_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n6647_), .ZN(new_n12298_));
  OAI21_X1   g12007(.A1(new_n930_), .A2(new_n7284_), .B(new_n12298_), .ZN(new_n12299_));
  AOI21_X1   g12008(.A1(new_n12299_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n12300_));
  XOR2_X1    g12009(.A1(new_n1114_), .A2(new_n12300_), .Z(new_n12301_));
  NOR2_X1    g12010(.A1(new_n12297_), .A2(new_n12301_), .ZN(new_n12302_));
  AOI22_X1   g12011(.A1(new_n12292_), .A2(new_n12194_), .B1(new_n12279_), .B2(new_n12289_), .ZN(new_n12303_));
  AOI21_X1   g12012(.A1(new_n12273_), .A2(new_n12265_), .B(new_n12277_), .ZN(new_n12304_));
  NOR3_X1    g12013(.A1(new_n12288_), .A2(new_n12283_), .A3(new_n12278_), .ZN(new_n12305_));
  NOR2_X1    g12014(.A1(new_n12305_), .A2(new_n12304_), .ZN(new_n12306_));
  NOR3_X1    g12015(.A1(new_n12306_), .A2(new_n12195_), .A3(new_n12198_), .ZN(new_n12307_));
  NOR2_X1    g12016(.A1(new_n12303_), .A2(new_n12307_), .ZN(new_n12308_));
  INV_X1     g12017(.I(new_n12301_), .ZN(new_n12309_));
  NOR2_X1    g12018(.A1(new_n12308_), .A2(new_n12309_), .ZN(new_n12310_));
  OAI22_X1   g12019(.A1(new_n12302_), .A2(new_n12310_), .B1(new_n12192_), .B2(new_n12189_), .ZN(new_n12311_));
  NOR2_X1    g12020(.A1(new_n12192_), .A2(new_n12189_), .ZN(new_n12312_));
  NAND2_X1   g12021(.A1(new_n12297_), .A2(new_n12309_), .ZN(new_n12313_));
  NAND2_X1   g12022(.A1(new_n12308_), .A2(new_n12301_), .ZN(new_n12314_));
  NAND2_X1   g12023(.A1(new_n12313_), .A2(new_n12314_), .ZN(new_n12315_));
  NAND2_X1   g12024(.A1(new_n12315_), .A2(new_n12312_), .ZN(new_n12316_));
  OAI22_X1   g12025(.A1(new_n5993_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n5991_), .ZN(new_n12317_));
  OAI21_X1   g12026(.A1(new_n1189_), .A2(new_n5997_), .B(new_n12317_), .ZN(new_n12318_));
  AOI21_X1   g12027(.A1(new_n12318_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n12319_));
  XNOR2_X1   g12028(.A1(new_n1421_), .A2(new_n12319_), .ZN(new_n12320_));
  AOI21_X1   g12029(.A1(new_n12316_), .A2(new_n12311_), .B(new_n12320_), .ZN(new_n12321_));
  NAND2_X1   g12030(.A1(new_n12186_), .A2(new_n12321_), .ZN(new_n12322_));
  OR3_X2     g12031(.A1(new_n11936_), .A2(new_n12321_), .A3(new_n11934_), .Z(new_n12323_));
  AOI21_X1   g12032(.A1(new_n12323_), .A2(new_n12322_), .B(new_n12185_), .ZN(new_n12324_));
  INV_X1     g12033(.I(new_n12322_), .ZN(new_n12325_));
  NOR2_X1    g12034(.A1(new_n12186_), .A2(new_n12321_), .ZN(new_n12326_));
  NOR3_X1    g12035(.A1(new_n12325_), .A2(new_n11933_), .A3(new_n12326_), .ZN(new_n12327_));
  OAI22_X1   g12036(.A1(new_n5420_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n5107_), .ZN(new_n12328_));
  OAI21_X1   g12037(.A1(new_n1525_), .A2(new_n5112_), .B(new_n12328_), .ZN(new_n12329_));
  AOI21_X1   g12038(.A1(new_n12329_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n12330_));
  XOR2_X1    g12039(.A1(new_n1808_), .A2(new_n12330_), .Z(new_n12331_));
  INV_X1     g12040(.I(new_n12331_), .ZN(new_n12332_));
  OAI21_X1   g12041(.A1(new_n12327_), .A2(new_n12324_), .B(new_n12332_), .ZN(new_n12333_));
  OAI21_X1   g12042(.A1(new_n12325_), .A2(new_n12326_), .B(new_n11933_), .ZN(new_n12334_));
  NAND3_X1   g12043(.A1(new_n12323_), .A2(new_n12185_), .A3(new_n12322_), .ZN(new_n12335_));
  NAND3_X1   g12044(.A1(new_n12334_), .A2(new_n12335_), .A3(new_n12331_), .ZN(new_n12336_));
  NAND2_X1   g12045(.A1(new_n12333_), .A2(new_n12336_), .ZN(new_n12337_));
  OAI21_X1   g12046(.A1(new_n11949_), .A2(new_n11964_), .B(new_n11950_), .ZN(new_n12338_));
  OAI22_X1   g12047(.A1(new_n4072_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n4067_), .ZN(new_n12339_));
  OAI21_X1   g12048(.A1(new_n1936_), .A2(new_n4318_), .B(new_n12339_), .ZN(new_n12340_));
  AOI21_X1   g12049(.A1(new_n12340_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n12341_));
  XNOR2_X1   g12050(.A1(new_n2280_), .A2(new_n12341_), .ZN(new_n12342_));
  XOR2_X1    g12051(.A1(new_n12338_), .A2(new_n12342_), .Z(new_n12343_));
  NAND2_X1   g12052(.A1(new_n12343_), .A2(new_n12337_), .ZN(new_n12344_));
  XOR2_X1    g12053(.A1(new_n12338_), .A2(new_n12342_), .Z(new_n12345_));
  OAI21_X1   g12054(.A1(new_n12337_), .A2(new_n12345_), .B(new_n12344_), .ZN(new_n12346_));
  NAND2_X1   g12055(.A1(new_n11562_), .A2(new_n11382_), .ZN(new_n12347_));
  INV_X1     g12056(.I(new_n12347_), .ZN(new_n12348_));
  NOR2_X1    g12057(.A1(new_n11966_), .A2(new_n11961_), .ZN(new_n12349_));
  NOR2_X1    g12058(.A1(new_n12349_), .A2(new_n11821_), .ZN(new_n12350_));
  AOI21_X1   g12059(.A1(new_n12349_), .A2(new_n11821_), .B(new_n11957_), .ZN(new_n12351_));
  AOI21_X1   g12060(.A1(new_n12348_), .A2(new_n12351_), .B(new_n12350_), .ZN(new_n12352_));
  OAI22_X1   g12061(.A1(new_n2643_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n2842_), .ZN(new_n12353_));
  OAI21_X1   g12062(.A1(new_n2439_), .A2(new_n3569_), .B(new_n12353_), .ZN(new_n12354_));
  AOI21_X1   g12063(.A1(new_n12354_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n12355_));
  XNOR2_X1   g12064(.A1(new_n2846_), .A2(new_n12355_), .ZN(new_n12356_));
  XOR2_X1    g12065(.A1(new_n12352_), .A2(new_n12356_), .Z(new_n12357_));
  INV_X1     g12066(.I(new_n12356_), .ZN(new_n12358_));
  XOR2_X1    g12067(.A1(new_n12352_), .A2(new_n12358_), .Z(new_n12359_));
  MUX2_X1    g12068(.I0(new_n12359_), .I1(new_n12357_), .S(new_n12346_), .Z(new_n12360_));
  XOR2_X1    g12069(.A1(new_n12360_), .A2(new_n12184_), .Z(new_n12361_));
  OAI22_X1   g12070(.A1(new_n3260_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n3709_), .ZN(new_n12362_));
  OAI21_X1   g12071(.A1(new_n3018_), .A2(new_n2884_), .B(new_n12362_), .ZN(new_n12363_));
  AOI21_X1   g12072(.A1(new_n12363_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n12364_));
  XNOR2_X1   g12073(.A1(new_n3514_), .A2(new_n12364_), .ZN(new_n12365_));
  XOR2_X1    g12074(.A1(new_n12361_), .A2(new_n12365_), .Z(new_n12366_));
  NOR2_X1    g12075(.A1(new_n11984_), .A2(new_n11985_), .ZN(new_n12367_));
  INV_X1     g12076(.I(new_n12367_), .ZN(new_n12368_));
  NAND2_X1   g12077(.A1(new_n11995_), .A2(new_n12368_), .ZN(new_n12369_));
  NOR2_X1    g12078(.A1(new_n11999_), .A2(new_n11989_), .ZN(new_n12370_));
  OAI21_X1   g12079(.A1(new_n11995_), .A2(new_n12368_), .B(new_n12370_), .ZN(new_n12371_));
  NAND2_X1   g12080(.A1(new_n12371_), .A2(new_n12369_), .ZN(new_n12372_));
  OAI22_X1   g12081(.A1(new_n2171_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n2166_), .ZN(new_n12373_));
  OAI21_X1   g12082(.A1(new_n3717_), .A2(new_n2322_), .B(new_n12373_), .ZN(new_n12374_));
  AOI21_X1   g12083(.A1(new_n12374_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n12375_));
  XNOR2_X1   g12084(.A1(new_n4257_), .A2(new_n12375_), .ZN(new_n12376_));
  INV_X1     g12085(.I(new_n12376_), .ZN(new_n12377_));
  XOR2_X1    g12086(.A1(new_n12372_), .A2(new_n12377_), .Z(new_n12378_));
  AOI21_X1   g12087(.A1(new_n12371_), .A2(new_n12369_), .B(new_n12376_), .ZN(new_n12379_));
  INV_X1     g12088(.I(new_n12379_), .ZN(new_n12380_));
  NAND3_X1   g12089(.A1(new_n12371_), .A2(new_n12369_), .A3(new_n12376_), .ZN(new_n12381_));
  AOI21_X1   g12090(.A1(new_n12380_), .A2(new_n12381_), .B(new_n12366_), .ZN(new_n12382_));
  AOI21_X1   g12091(.A1(new_n12378_), .A2(new_n12366_), .B(new_n12382_), .ZN(new_n12383_));
  NOR2_X1    g12092(.A1(new_n11997_), .A2(new_n12002_), .ZN(new_n12384_));
  NAND3_X1   g12093(.A1(new_n12012_), .A2(new_n12013_), .A3(new_n11800_), .ZN(new_n12385_));
  NAND2_X1   g12094(.A1(new_n12385_), .A2(new_n12007_), .ZN(new_n12386_));
  OAI22_X1   g12095(.A1(new_n12386_), .A2(new_n12011_), .B1(new_n11800_), .B2(new_n12384_), .ZN(new_n12387_));
  OAI22_X1   g12096(.A1(new_n1712_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n1707_), .ZN(new_n12388_));
  OAI21_X1   g12097(.A1(new_n4500_), .A2(new_n1850_), .B(new_n12388_), .ZN(new_n12389_));
  AOI21_X1   g12098(.A1(new_n12389_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n12390_));
  XOR2_X1    g12099(.A1(new_n5067_), .A2(new_n12390_), .Z(new_n12391_));
  INV_X1     g12100(.I(new_n12391_), .ZN(new_n12392_));
  NAND2_X1   g12101(.A1(new_n12387_), .A2(new_n12392_), .ZN(new_n12393_));
  INV_X1     g12102(.I(new_n12384_), .ZN(new_n12394_));
  AOI21_X1   g12103(.A1(new_n12384_), .A2(new_n11800_), .B(new_n12006_), .ZN(new_n12395_));
  AOI22_X1   g12104(.A1(new_n12395_), .A2(new_n11802_), .B1(new_n11799_), .B2(new_n12394_), .ZN(new_n12396_));
  NAND2_X1   g12105(.A1(new_n12396_), .A2(new_n12391_), .ZN(new_n12397_));
  AOI21_X1   g12106(.A1(new_n12397_), .A2(new_n12393_), .B(new_n12383_), .ZN(new_n12398_));
  XNOR2_X1   g12107(.A1(new_n12361_), .A2(new_n12365_), .ZN(new_n12399_));
  XOR2_X1    g12108(.A1(new_n12372_), .A2(new_n12376_), .Z(new_n12400_));
  INV_X1     g12109(.I(new_n12381_), .ZN(new_n12401_));
  OAI21_X1   g12110(.A1(new_n12401_), .A2(new_n12379_), .B(new_n12399_), .ZN(new_n12402_));
  OAI21_X1   g12111(.A1(new_n12400_), .A2(new_n12399_), .B(new_n12402_), .ZN(new_n12403_));
  NAND2_X1   g12112(.A1(new_n12396_), .A2(new_n12392_), .ZN(new_n12404_));
  NAND2_X1   g12113(.A1(new_n12387_), .A2(new_n12391_), .ZN(new_n12405_));
  AOI21_X1   g12114(.A1(new_n12404_), .A2(new_n12405_), .B(new_n12403_), .ZN(new_n12406_));
  NOR2_X1    g12115(.A1(new_n12398_), .A2(new_n12406_), .ZN(new_n12407_));
  NOR3_X1    g12116(.A1(new_n12177_), .A2(new_n12175_), .A3(new_n12407_), .ZN(new_n12408_));
  INV_X1     g12117(.I(new_n12175_), .ZN(new_n12409_));
  NAND3_X1   g12118(.A1(new_n12046_), .A2(new_n12047_), .A3(new_n11639_), .ZN(new_n12410_));
  NAND3_X1   g12119(.A1(new_n11796_), .A2(new_n12410_), .A3(new_n12041_), .ZN(new_n12411_));
  OR2_X2     g12120(.A1(new_n12398_), .A2(new_n12406_), .Z(new_n12412_));
  AOI21_X1   g12121(.A1(new_n12411_), .A2(new_n12409_), .B(new_n12412_), .ZN(new_n12413_));
  OAI21_X1   g12122(.A1(new_n12408_), .A2(new_n12413_), .B(new_n12174_), .ZN(new_n12414_));
  NAND3_X1   g12123(.A1(new_n12016_), .A2(new_n12019_), .A3(new_n11621_), .ZN(new_n12415_));
  NAND2_X1   g12124(.A1(new_n12415_), .A2(new_n12030_), .ZN(new_n12416_));
  OAI22_X1   g12125(.A1(new_n12416_), .A2(new_n11798_), .B1(new_n11621_), .B2(new_n12171_), .ZN(new_n12417_));
  NAND3_X1   g12126(.A1(new_n12411_), .A2(new_n12409_), .A3(new_n12412_), .ZN(new_n12418_));
  OAI21_X1   g12127(.A1(new_n12177_), .A2(new_n12175_), .B(new_n12407_), .ZN(new_n12419_));
  NAND3_X1   g12128(.A1(new_n12419_), .A2(new_n12418_), .A3(new_n12417_), .ZN(new_n12420_));
  AOI21_X1   g12129(.A1(new_n12414_), .A2(new_n12420_), .B(new_n12170_), .ZN(new_n12421_));
  AOI21_X1   g12130(.A1(new_n12419_), .A2(new_n12418_), .B(new_n12417_), .ZN(new_n12422_));
  NOR3_X1    g12131(.A1(new_n12408_), .A2(new_n12413_), .A3(new_n12174_), .ZN(new_n12423_));
  NOR3_X1    g12132(.A1(new_n12423_), .A2(new_n12422_), .A3(new_n12169_), .ZN(new_n12424_));
  OAI22_X1   g12133(.A1(new_n1055_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n1061_), .ZN(new_n12425_));
  OAI21_X1   g12134(.A1(new_n6229_), .A2(new_n1332_), .B(new_n12425_), .ZN(new_n12426_));
  AOI21_X1   g12135(.A1(new_n12426_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n12427_));
  XOR2_X1    g12136(.A1(new_n6851_), .A2(new_n12427_), .Z(new_n12428_));
  NOR3_X1    g12137(.A1(new_n12424_), .A2(new_n12421_), .A3(new_n12428_), .ZN(new_n12429_));
  OAI21_X1   g12138(.A1(new_n12423_), .A2(new_n12422_), .B(new_n12169_), .ZN(new_n12430_));
  NAND3_X1   g12139(.A1(new_n12414_), .A2(new_n12420_), .A3(new_n12170_), .ZN(new_n12431_));
  INV_X1     g12140(.I(new_n12428_), .ZN(new_n12432_));
  AOI21_X1   g12141(.A1(new_n12430_), .A2(new_n12431_), .B(new_n12432_), .ZN(new_n12433_));
  OAI21_X1   g12142(.A1(new_n12429_), .A2(new_n12433_), .B(new_n12165_), .ZN(new_n12434_));
  AOI21_X1   g12143(.A1(new_n12161_), .A2(new_n11657_), .B(new_n12057_), .ZN(new_n12435_));
  AOI22_X1   g12144(.A1(new_n12435_), .A2(new_n12061_), .B1(new_n11663_), .B2(new_n12162_), .ZN(new_n12436_));
  AOI21_X1   g12145(.A1(new_n12430_), .A2(new_n12431_), .B(new_n12428_), .ZN(new_n12437_));
  NOR3_X1    g12146(.A1(new_n12424_), .A2(new_n12421_), .A3(new_n12432_), .ZN(new_n12438_));
  OAI21_X1   g12147(.A1(new_n12437_), .A2(new_n12438_), .B(new_n12436_), .ZN(new_n12439_));
  OAI22_X1   g12148(.A1(new_n970_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n820_), .ZN(new_n12440_));
  OAI21_X1   g12149(.A1(new_n7198_), .A2(new_n894_), .B(new_n12440_), .ZN(new_n12441_));
  AOI21_X1   g12150(.A1(new_n12441_), .A2(new_n827_), .B(new_n970_), .ZN(new_n12442_));
  XNOR2_X1   g12151(.A1(new_n7874_), .A2(new_n12442_), .ZN(new_n12443_));
  INV_X1     g12152(.I(new_n12443_), .ZN(new_n12444_));
  NAND3_X1   g12153(.A1(new_n12439_), .A2(new_n12434_), .A3(new_n12444_), .ZN(new_n12445_));
  NAND3_X1   g12154(.A1(new_n12430_), .A2(new_n12431_), .A3(new_n12432_), .ZN(new_n12446_));
  OAI21_X1   g12155(.A1(new_n12424_), .A2(new_n12421_), .B(new_n12428_), .ZN(new_n12447_));
  AOI21_X1   g12156(.A1(new_n12447_), .A2(new_n12446_), .B(new_n12436_), .ZN(new_n12448_));
  OAI21_X1   g12157(.A1(new_n12424_), .A2(new_n12421_), .B(new_n12432_), .ZN(new_n12449_));
  NAND3_X1   g12158(.A1(new_n12430_), .A2(new_n12431_), .A3(new_n12428_), .ZN(new_n12450_));
  AOI21_X1   g12159(.A1(new_n12449_), .A2(new_n12450_), .B(new_n12165_), .ZN(new_n12451_));
  OAI21_X1   g12160(.A1(new_n12448_), .A2(new_n12451_), .B(new_n12443_), .ZN(new_n12452_));
  AOI21_X1   g12161(.A1(new_n12445_), .A2(new_n12452_), .B(new_n12158_), .ZN(new_n12453_));
  OAI21_X1   g12162(.A1(new_n12067_), .A2(new_n12064_), .B(new_n12081_), .ZN(new_n12454_));
  INV_X1     g12163(.I(new_n12156_), .ZN(new_n12455_));
  NAND3_X1   g12164(.A1(new_n11773_), .A2(new_n11790_), .A3(new_n12072_), .ZN(new_n12456_));
  OAI21_X1   g12165(.A1(new_n12455_), .A2(new_n12456_), .B(new_n12454_), .ZN(new_n12457_));
  NAND2_X1   g12166(.A1(new_n12439_), .A2(new_n12434_), .ZN(new_n12458_));
  NAND2_X1   g12167(.A1(new_n12458_), .A2(new_n12444_), .ZN(new_n12459_));
  NOR2_X1    g12168(.A1(new_n12448_), .A2(new_n12451_), .ZN(new_n12460_));
  NAND2_X1   g12169(.A1(new_n12460_), .A2(new_n12443_), .ZN(new_n12461_));
  AOI21_X1   g12170(.A1(new_n12459_), .A2(new_n12461_), .B(new_n12457_), .ZN(new_n12462_));
  OAI22_X1   g12171(.A1(new_n607_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n610_), .ZN(new_n12463_));
  OAI21_X1   g12172(.A1(new_n8218_), .A2(new_n684_), .B(new_n12463_), .ZN(new_n12464_));
  AOI21_X1   g12173(.A1(new_n12464_), .A2(new_n612_), .B(new_n607_), .ZN(new_n12465_));
  XOR2_X1    g12174(.A1(new_n8952_), .A2(new_n12465_), .Z(new_n12466_));
  INV_X1     g12175(.I(new_n12466_), .ZN(new_n12467_));
  OAI21_X1   g12176(.A1(new_n12462_), .A2(new_n12453_), .B(new_n12467_), .ZN(new_n12468_));
  NOR2_X1    g12177(.A1(new_n12462_), .A2(new_n12453_), .ZN(new_n12469_));
  NAND2_X1   g12178(.A1(new_n12469_), .A2(new_n12466_), .ZN(new_n12470_));
  NAND2_X1   g12179(.A1(new_n12470_), .A2(new_n12468_), .ZN(new_n12471_));
  AOI21_X1   g12180(.A1(new_n12083_), .A2(new_n12082_), .B(new_n12081_), .ZN(new_n12472_));
  NOR3_X1    g12181(.A1(new_n12074_), .A2(new_n12079_), .A3(new_n11784_), .ZN(new_n12473_));
  NOR2_X1    g12182(.A1(new_n12473_), .A2(new_n12472_), .ZN(new_n12474_));
  NOR3_X1    g12183(.A1(new_n11781_), .A2(new_n11783_), .A3(new_n12474_), .ZN(new_n12475_));
  XOR2_X1    g12184(.A1(new_n11774_), .A2(new_n11361_), .Z(new_n12476_));
  INV_X1     g12185(.I(new_n12088_), .ZN(new_n12477_));
  NAND3_X1   g12186(.A1(new_n12476_), .A2(new_n11677_), .A3(new_n12477_), .ZN(new_n12478_));
  AOI21_X1   g12187(.A1(new_n12096_), .A2(new_n12474_), .B(new_n12478_), .ZN(new_n12479_));
  OAI22_X1   g12188(.A1(new_n448_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n450_), .ZN(new_n12480_));
  OAI21_X1   g12189(.A1(new_n9295_), .A2(new_n496_), .B(new_n12480_), .ZN(new_n12481_));
  AOI21_X1   g12190(.A1(new_n12481_), .A2(new_n452_), .B(new_n448_), .ZN(new_n12482_));
  XNOR2_X1   g12191(.A1(new_n10035_), .A2(new_n12482_), .ZN(new_n12483_));
  INV_X1     g12192(.I(new_n12483_), .ZN(new_n12484_));
  OAI21_X1   g12193(.A1(new_n12479_), .A2(new_n12475_), .B(new_n12484_), .ZN(new_n12485_));
  INV_X1     g12194(.I(new_n12485_), .ZN(new_n12486_));
  NOR3_X1    g12195(.A1(new_n12479_), .A2(new_n12475_), .A3(new_n12484_), .ZN(new_n12487_));
  OAI21_X1   g12196(.A1(new_n12486_), .A2(new_n12487_), .B(new_n12471_), .ZN(new_n12488_));
  AND2_X2    g12197(.A1(new_n12470_), .A2(new_n12468_), .Z(new_n12489_));
  NOR3_X1    g12198(.A1(new_n12479_), .A2(new_n12475_), .A3(new_n12483_), .ZN(new_n12490_));
  OAI21_X1   g12199(.A1(new_n11781_), .A2(new_n11783_), .B(new_n12474_), .ZN(new_n12491_));
  NOR2_X1    g12200(.A1(new_n11778_), .A2(new_n12088_), .ZN(new_n12492_));
  AOI21_X1   g12201(.A1(new_n12491_), .A2(new_n12492_), .B(new_n12475_), .ZN(new_n12493_));
  NOR2_X1    g12202(.A1(new_n12493_), .A2(new_n12484_), .ZN(new_n12494_));
  OAI21_X1   g12203(.A1(new_n12494_), .A2(new_n12490_), .B(new_n12489_), .ZN(new_n12495_));
  NAND2_X1   g12204(.A1(new_n12488_), .A2(new_n12495_), .ZN(new_n12496_));
  OAI22_X1   g12205(.A1(new_n10862_), .A2(new_n341_), .B1(new_n404_), .B2(new_n11738_), .ZN(new_n12497_));
  OAI21_X1   g12206(.A1(new_n10477_), .A2(new_n366_), .B(new_n12497_), .ZN(new_n12498_));
  AOI21_X1   g12207(.A1(new_n12498_), .A2(new_n334_), .B(new_n341_), .ZN(new_n12499_));
  XOR2_X1    g12208(.A1(new_n11298_), .A2(new_n12499_), .Z(new_n12500_));
  INV_X1     g12209(.I(new_n12500_), .ZN(new_n12501_));
  NAND2_X1   g12210(.A1(new_n12496_), .A2(new_n12501_), .ZN(new_n12502_));
  INV_X1     g12211(.I(new_n12487_), .ZN(new_n12503_));
  AOI21_X1   g12212(.A1(new_n12503_), .A2(new_n12485_), .B(new_n12489_), .ZN(new_n12504_));
  INV_X1     g12213(.I(new_n12490_), .ZN(new_n12505_));
  OAI21_X1   g12214(.A1(new_n12479_), .A2(new_n12475_), .B(new_n12483_), .ZN(new_n12506_));
  AOI21_X1   g12215(.A1(new_n12505_), .A2(new_n12506_), .B(new_n12471_), .ZN(new_n12507_));
  NOR2_X1    g12216(.A1(new_n12504_), .A2(new_n12507_), .ZN(new_n12508_));
  NAND2_X1   g12217(.A1(new_n12508_), .A2(new_n12500_), .ZN(new_n12509_));
  AOI21_X1   g12218(.A1(new_n12509_), .A2(new_n12502_), .B(new_n12154_), .ZN(new_n12510_));
  NAND2_X1   g12219(.A1(new_n11772_), .A2(new_n11770_), .ZN(new_n12511_));
  OAI21_X1   g12220(.A1(new_n12151_), .A2(new_n11768_), .B(new_n12103_), .ZN(new_n12512_));
  OAI22_X1   g12221(.A1(new_n12511_), .A2(new_n12512_), .B1(new_n11707_), .B2(new_n12152_), .ZN(new_n12513_));
  NAND3_X1   g12222(.A1(new_n12488_), .A2(new_n12495_), .A3(new_n12501_), .ZN(new_n12514_));
  OAI21_X1   g12223(.A1(new_n12504_), .A2(new_n12507_), .B(new_n12500_), .ZN(new_n12515_));
  AOI21_X1   g12224(.A1(new_n12514_), .A2(new_n12515_), .B(new_n12513_), .ZN(new_n12516_));
  NOR2_X1    g12225(.A1(new_n12510_), .A2(new_n12516_), .ZN(new_n12517_));
  NOR3_X1    g12226(.A1(new_n12517_), .A2(new_n12148_), .A3(new_n12149_), .ZN(new_n12518_));
  NAND2_X1   g12227(.A1(new_n12113_), .A2(new_n12116_), .ZN(new_n12519_));
  NAND2_X1   g12228(.A1(new_n12519_), .A2(new_n12121_), .ZN(new_n12520_));
  INV_X1     g12229(.I(new_n12520_), .ZN(new_n12521_));
  OAI21_X1   g12230(.A1(new_n12518_), .A2(new_n12521_), .B(new_n12141_), .ZN(new_n12522_));
  NAND2_X1   g12231(.A1(new_n12125_), .A2(new_n12122_), .ZN(new_n12523_));
  INV_X1     g12232(.I(new_n12149_), .ZN(new_n12524_));
  NOR2_X1    g12233(.A1(new_n12508_), .A2(new_n12500_), .ZN(new_n12525_));
  NOR2_X1    g12234(.A1(new_n12496_), .A2(new_n12501_), .ZN(new_n12526_));
  OAI21_X1   g12235(.A1(new_n12525_), .A2(new_n12526_), .B(new_n12513_), .ZN(new_n12527_));
  NAND2_X1   g12236(.A1(new_n12515_), .A2(new_n12514_), .ZN(new_n12528_));
  NAND2_X1   g12237(.A1(new_n12528_), .A2(new_n12154_), .ZN(new_n12529_));
  NAND2_X1   g12238(.A1(new_n12527_), .A2(new_n12529_), .ZN(new_n12530_));
  NAND3_X1   g12239(.A1(new_n12530_), .A2(new_n12523_), .A3(new_n12524_), .ZN(new_n12531_));
  NAND3_X1   g12240(.A1(new_n12531_), .A2(new_n11765_), .A3(new_n12520_), .ZN(new_n12532_));
  NAND2_X1   g12241(.A1(new_n12522_), .A2(new_n12532_), .ZN(new_n12533_));
  NOR2_X1    g12242(.A1(\b[56] ), .A2(\b[57] ), .ZN(new_n12534_));
  AOI21_X1   g12243(.A1(new_n11742_), .A2(new_n12534_), .B(new_n11738_), .ZN(new_n12535_));
  INV_X1     g12244(.I(\b[57] ), .ZN(new_n12536_));
  NOR2_X1    g12245(.A1(new_n11744_), .A2(new_n12536_), .ZN(new_n12537_));
  INV_X1     g12246(.I(new_n12537_), .ZN(new_n12538_));
  NOR2_X1    g12247(.A1(new_n11742_), .A2(new_n12538_), .ZN(new_n12539_));
  NOR2_X1    g12248(.A1(new_n12535_), .A2(new_n12539_), .ZN(new_n12540_));
  XNOR2_X1   g12249(.A1(\b[57] ), .A2(\b[58] ), .ZN(new_n12541_));
  INV_X1     g12250(.I(\b[58] ), .ZN(new_n12542_));
  NOR2_X1    g12251(.A1(new_n12536_), .A2(new_n12542_), .ZN(new_n12543_));
  NOR2_X1    g12252(.A1(\b[57] ), .A2(\b[58] ), .ZN(new_n12544_));
  OAI21_X1   g12253(.A1(new_n12543_), .A2(new_n12544_), .B(new_n12540_), .ZN(new_n12545_));
  OAI21_X1   g12254(.A1(new_n12540_), .A2(new_n12541_), .B(new_n12545_), .ZN(new_n12546_));
  OAI22_X1   g12255(.A1(new_n330_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n263_), .ZN(new_n12547_));
  OAI21_X1   g12256(.A1(new_n11744_), .A2(new_n289_), .B(new_n12547_), .ZN(new_n12548_));
  AOI21_X1   g12257(.A1(new_n12548_), .A2(new_n260_), .B(new_n426_), .ZN(new_n12549_));
  XNOR2_X1   g12258(.A1(new_n12546_), .A2(new_n12549_), .ZN(new_n12550_));
  XOR2_X1    g12259(.A1(new_n12533_), .A2(new_n12550_), .Z(new_n12551_));
  NAND2_X1   g12260(.A1(new_n12139_), .A2(new_n12144_), .ZN(new_n12552_));
  AOI21_X1   g12261(.A1(new_n12552_), .A2(new_n11735_), .B(new_n11753_), .ZN(new_n12553_));
  NOR2_X1    g12262(.A1(new_n12552_), .A2(new_n11735_), .ZN(new_n12554_));
  NOR4_X1    g12263(.A1(new_n12553_), .A2(new_n12554_), .A3(new_n11332_), .A4(new_n11346_), .ZN(new_n12555_));
  NOR2_X1    g12264(.A1(new_n11765_), .A2(new_n12148_), .ZN(new_n12556_));
  NOR2_X1    g12265(.A1(new_n12523_), .A2(new_n12141_), .ZN(new_n12557_));
  OAI21_X1   g12266(.A1(new_n12556_), .A2(new_n12557_), .B(new_n12133_), .ZN(new_n12558_));
  INV_X1     g12267(.I(new_n12558_), .ZN(new_n12559_));
  NOR2_X1    g12268(.A1(new_n12555_), .A2(new_n12559_), .ZN(new_n12560_));
  NAND2_X1   g12269(.A1(new_n12551_), .A2(new_n12558_), .ZN(new_n12561_));
  OAI22_X1   g12270(.A1(new_n12561_), .A2(new_n12555_), .B1(new_n12551_), .B2(new_n12560_), .ZN(\f[58] ));
  OAI21_X1   g12271(.A1(new_n12135_), .A2(new_n12136_), .B(new_n12137_), .ZN(new_n12563_));
  NAND3_X1   g12272(.A1(new_n12125_), .A2(new_n12122_), .A3(new_n12133_), .ZN(new_n12564_));
  AOI21_X1   g12273(.A1(new_n12563_), .A2(new_n12564_), .B(new_n12141_), .ZN(new_n12565_));
  NAND3_X1   g12274(.A1(new_n12125_), .A2(new_n12122_), .A3(new_n12137_), .ZN(new_n12566_));
  OAI21_X1   g12275(.A1(new_n12135_), .A2(new_n12136_), .B(new_n12133_), .ZN(new_n12567_));
  AOI21_X1   g12276(.A1(new_n12567_), .A2(new_n12566_), .B(new_n11765_), .ZN(new_n12568_));
  OAI21_X1   g12277(.A1(new_n12568_), .A2(new_n12565_), .B(new_n11735_), .ZN(new_n12569_));
  NAND2_X1   g12278(.A1(new_n12569_), .A2(new_n11752_), .ZN(new_n12570_));
  NAND3_X1   g12279(.A1(new_n11755_), .A2(new_n12139_), .A3(new_n12144_), .ZN(new_n12571_));
  NAND3_X1   g12280(.A1(new_n11347_), .A2(new_n12570_), .A3(new_n12571_), .ZN(new_n12572_));
  NAND2_X1   g12281(.A1(new_n12533_), .A2(new_n12559_), .ZN(new_n12573_));
  INV_X1     g12282(.I(new_n12550_), .ZN(new_n12574_));
  OAI21_X1   g12283(.A1(new_n12533_), .A2(new_n12559_), .B(new_n12574_), .ZN(new_n12575_));
  OAI21_X1   g12284(.A1(new_n12572_), .A2(new_n12575_), .B(new_n12573_), .ZN(new_n12576_));
  AOI21_X1   g12285(.A1(new_n11765_), .A2(new_n12125_), .B(new_n12135_), .ZN(new_n12577_));
  XOR2_X1    g12286(.A1(new_n12513_), .A2(new_n12496_), .Z(new_n12578_));
  NOR2_X1    g12287(.A1(new_n12578_), .A2(new_n12500_), .ZN(new_n12579_));
  NOR2_X1    g12288(.A1(new_n12489_), .A2(new_n12493_), .ZN(new_n12580_));
  NOR3_X1    g12289(.A1(new_n12479_), .A2(new_n12471_), .A3(new_n12475_), .ZN(new_n12581_));
  NOR2_X1    g12290(.A1(new_n12580_), .A2(new_n12581_), .ZN(new_n12582_));
  NOR2_X1    g12291(.A1(new_n12582_), .A2(new_n12483_), .ZN(new_n12583_));
  NAND2_X1   g12292(.A1(new_n12469_), .A2(new_n12467_), .ZN(new_n12584_));
  OAI22_X1   g12293(.A1(new_n12479_), .A2(new_n12475_), .B1(new_n12469_), .B2(new_n12467_), .ZN(new_n12585_));
  NAND2_X1   g12294(.A1(new_n12452_), .A2(new_n12445_), .ZN(new_n12586_));
  OAI21_X1   g12295(.A1(new_n12436_), .A2(new_n12433_), .B(new_n12446_), .ZN(new_n12587_));
  AOI21_X1   g12296(.A1(new_n12411_), .A2(new_n12409_), .B(new_n12169_), .ZN(new_n12588_));
  INV_X1     g12297(.I(new_n12588_), .ZN(new_n12589_));
  NAND3_X1   g12298(.A1(new_n12411_), .A2(new_n12169_), .A3(new_n12409_), .ZN(new_n12590_));
  XOR2_X1    g12299(.A1(new_n12417_), .A2(new_n12407_), .Z(new_n12591_));
  INV_X1     g12300(.I(new_n12591_), .ZN(new_n12592_));
  NAND2_X1   g12301(.A1(new_n12590_), .A2(new_n12592_), .ZN(new_n12593_));
  NAND2_X1   g12302(.A1(new_n12387_), .A2(new_n12383_), .ZN(new_n12594_));
  NAND2_X1   g12303(.A1(new_n12396_), .A2(new_n12403_), .ZN(new_n12595_));
  AOI21_X1   g12304(.A1(new_n12595_), .A2(new_n12594_), .B(new_n12392_), .ZN(new_n12596_));
  NAND2_X1   g12305(.A1(new_n12372_), .A2(new_n12366_), .ZN(new_n12597_));
  NAND3_X1   g12306(.A1(new_n12399_), .A2(new_n12369_), .A3(new_n12371_), .ZN(new_n12598_));
  AOI21_X1   g12307(.A1(new_n12598_), .A2(new_n12597_), .B(new_n12377_), .ZN(new_n12599_));
  NOR2_X1    g12308(.A1(new_n12361_), .A2(new_n12365_), .ZN(new_n12600_));
  INV_X1     g12309(.I(new_n12600_), .ZN(new_n12601_));
  NOR2_X1    g12310(.A1(new_n11813_), .A2(new_n12367_), .ZN(new_n12602_));
  NAND2_X1   g12311(.A1(new_n11811_), .A2(new_n11990_), .ZN(new_n12603_));
  AOI21_X1   g12312(.A1(new_n11813_), .A2(new_n12367_), .B(new_n12603_), .ZN(new_n12604_));
  NAND2_X1   g12313(.A1(new_n12361_), .A2(new_n12365_), .ZN(new_n12605_));
  OAI21_X1   g12314(.A1(new_n12604_), .A2(new_n12602_), .B(new_n12605_), .ZN(new_n12606_));
  OAI22_X1   g12315(.A1(new_n2842_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n3018_), .ZN(new_n12607_));
  OAI21_X1   g12316(.A1(new_n2643_), .A2(new_n3569_), .B(new_n12607_), .ZN(new_n12608_));
  AOI21_X1   g12317(.A1(new_n12608_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n12609_));
  XNOR2_X1   g12318(.A1(new_n3022_), .A2(new_n12609_), .ZN(new_n12610_));
  NAND2_X1   g12319(.A1(new_n12316_), .A2(new_n12311_), .ZN(new_n12611_));
  INV_X1     g12320(.I(new_n12611_), .ZN(new_n12612_));
  NOR2_X1    g12321(.A1(new_n12612_), .A2(new_n11933_), .ZN(new_n12613_));
  INV_X1     g12322(.I(new_n12320_), .ZN(new_n12614_));
  OAI21_X1   g12323(.A1(new_n12611_), .A2(new_n12185_), .B(new_n12614_), .ZN(new_n12615_));
  NOR2_X1    g12324(.A1(new_n12615_), .A2(new_n12186_), .ZN(new_n12616_));
  NOR2_X1    g12325(.A1(new_n12616_), .A2(new_n12613_), .ZN(new_n12617_));
  OAI22_X1   g12326(.A1(new_n6644_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n6647_), .ZN(new_n12618_));
  OAI21_X1   g12327(.A1(new_n1017_), .A2(new_n7284_), .B(new_n12618_), .ZN(new_n12619_));
  AOI21_X1   g12328(.A1(new_n12619_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n12620_));
  XNOR2_X1   g12329(.A1(new_n1196_), .A2(new_n12620_), .ZN(new_n12621_));
  INV_X1     g12330(.I(new_n12621_), .ZN(new_n12622_));
  OAI21_X1   g12331(.A1(new_n12198_), .A2(new_n12195_), .B(new_n12289_), .ZN(new_n12623_));
  NAND2_X1   g12332(.A1(new_n12623_), .A2(new_n12279_), .ZN(new_n12624_));
  INV_X1     g12333(.I(new_n12624_), .ZN(new_n12625_));
  INV_X1     g12334(.I(new_n12313_), .ZN(new_n12626_));
  NAND4_X1   g12335(.A1(new_n11828_), .A2(new_n11826_), .A3(new_n11911_), .A4(new_n12190_), .ZN(new_n12627_));
  AOI22_X1   g12336(.A1(new_n12627_), .A2(new_n12188_), .B1(new_n12308_), .B2(new_n12301_), .ZN(new_n12628_));
  INV_X1     g12337(.I(new_n12253_), .ZN(new_n12629_));
  AOI22_X1   g12338(.A1(new_n12204_), .A2(new_n11861_), .B1(new_n12244_), .B2(new_n12247_), .ZN(new_n12630_));
  NOR2_X1    g12339(.A1(new_n12630_), .A2(new_n12629_), .ZN(new_n12631_));
  NAND2_X1   g12340(.A1(new_n12208_), .A2(new_n12239_), .ZN(new_n12632_));
  NOR3_X1    g12341(.A1(new_n12230_), .A2(new_n258_), .A3(new_n11850_), .ZN(new_n12633_));
  XNOR2_X1   g12342(.A1(\a[56] ), .A2(\a[58] ), .ZN(new_n12634_));
  XNOR2_X1   g12343(.A1(\a[56] ), .A2(\a[59] ), .ZN(new_n12635_));
  XNOR2_X1   g12344(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n12636_));
  OR3_X2     g12345(.A1(new_n12634_), .A2(new_n12635_), .A3(new_n12636_), .Z(new_n12637_));
  OAI22_X1   g12346(.A1(new_n12226_), .A2(new_n10132_), .B1(new_n12637_), .B2(new_n258_), .ZN(new_n12638_));
  AOI21_X1   g12347(.A1(new_n12638_), .A2(new_n12222_), .B(new_n490_), .ZN(new_n12639_));
  XOR2_X1    g12348(.A1(new_n12639_), .A2(new_n12214_), .Z(new_n12640_));
  NAND2_X1   g12349(.A1(new_n12640_), .A2(new_n12633_), .ZN(new_n12641_));
  NAND2_X1   g12350(.A1(new_n12231_), .A2(new_n12206_), .ZN(new_n12642_));
  INV_X1     g12351(.I(new_n12214_), .ZN(new_n12643_));
  XOR2_X1    g12352(.A1(new_n12639_), .A2(new_n12643_), .Z(new_n12644_));
  NAND2_X1   g12353(.A1(new_n12644_), .A2(new_n12642_), .ZN(new_n12645_));
  NAND2_X1   g12354(.A1(new_n12645_), .A2(new_n12641_), .ZN(new_n12646_));
  AOI22_X1   g12355(.A1(new_n10969_), .A2(new_n413_), .B1(new_n11394_), .B2(\b[3] ), .ZN(new_n12647_));
  OAI21_X1   g12356(.A1(new_n12647_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n12648_));
  XOR2_X1    g12357(.A1(new_n12648_), .A2(new_n378_), .Z(new_n12649_));
  NOR2_X1    g12358(.A1(new_n12646_), .A2(new_n12649_), .ZN(new_n12650_));
  NOR2_X1    g12359(.A1(new_n12644_), .A2(new_n12642_), .ZN(new_n12651_));
  NOR2_X1    g12360(.A1(new_n12640_), .A2(new_n12633_), .ZN(new_n12652_));
  NOR2_X1    g12361(.A1(new_n12651_), .A2(new_n12652_), .ZN(new_n12653_));
  INV_X1     g12362(.I(new_n12649_), .ZN(new_n12654_));
  NOR2_X1    g12363(.A1(new_n12653_), .A2(new_n12654_), .ZN(new_n12655_));
  NOR2_X1    g12364(.A1(new_n12655_), .A2(new_n12650_), .ZN(new_n12656_));
  AOI21_X1   g12365(.A1(new_n12241_), .A2(new_n12632_), .B(new_n12656_), .ZN(new_n12657_));
  NAND2_X1   g12366(.A1(new_n12632_), .A2(new_n12241_), .ZN(new_n12658_));
  NOR2_X1    g12367(.A1(new_n12653_), .A2(new_n12649_), .ZN(new_n12659_));
  NOR2_X1    g12368(.A1(new_n12646_), .A2(new_n12654_), .ZN(new_n12660_));
  NOR2_X1    g12369(.A1(new_n12659_), .A2(new_n12660_), .ZN(new_n12661_));
  NOR2_X1    g12370(.A1(new_n12658_), .A2(new_n12661_), .ZN(new_n12662_));
  AOI22_X1   g12371(.A1(new_n11415_), .A2(new_n517_), .B1(\b[6] ), .B2(new_n10145_), .ZN(new_n12663_));
  OAI21_X1   g12372(.A1(new_n12663_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n12664_));
  XOR2_X1    g12373(.A1(new_n522_), .A2(new_n12664_), .Z(new_n12665_));
  NOR3_X1    g12374(.A1(new_n12657_), .A2(new_n12662_), .A3(new_n12665_), .ZN(new_n12666_));
  OAI21_X1   g12375(.A1(new_n12650_), .A2(new_n12655_), .B(new_n12658_), .ZN(new_n12667_));
  INV_X1     g12376(.I(new_n12662_), .ZN(new_n12668_));
  INV_X1     g12377(.I(new_n12665_), .ZN(new_n12669_));
  AOI21_X1   g12378(.A1(new_n12668_), .A2(new_n12667_), .B(new_n12669_), .ZN(new_n12670_));
  NOR2_X1    g12379(.A1(new_n12670_), .A2(new_n12666_), .ZN(new_n12671_));
  NOR2_X1    g12380(.A1(new_n12671_), .A2(new_n12631_), .ZN(new_n12672_));
  NAND3_X1   g12381(.A1(new_n12668_), .A2(new_n12667_), .A3(new_n12669_), .ZN(new_n12673_));
  OAI21_X1   g12382(.A1(new_n12657_), .A2(new_n12662_), .B(new_n12665_), .ZN(new_n12674_));
  NAND2_X1   g12383(.A1(new_n12673_), .A2(new_n12674_), .ZN(new_n12675_));
  NOR3_X1    g12384(.A1(new_n12675_), .A2(new_n12629_), .A3(new_n12630_), .ZN(new_n12676_));
  OAI22_X1   g12385(.A1(new_n8644_), .A2(new_n656_), .B1(new_n706_), .B2(new_n9388_), .ZN(new_n12677_));
  OAI21_X1   g12386(.A1(new_n565_), .A2(new_n10154_), .B(new_n12677_), .ZN(new_n12678_));
  AOI21_X1   g12387(.A1(new_n12678_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n12679_));
  XNOR2_X1   g12388(.A1(new_n710_), .A2(new_n12679_), .ZN(new_n12680_));
  INV_X1     g12389(.I(new_n12680_), .ZN(new_n12681_));
  OAI21_X1   g12390(.A1(new_n12672_), .A2(new_n12676_), .B(new_n12681_), .ZN(new_n12682_));
  OAI21_X1   g12391(.A1(new_n12629_), .A2(new_n12630_), .B(new_n12675_), .ZN(new_n12683_));
  NAND2_X1   g12392(.A1(new_n12671_), .A2(new_n12631_), .ZN(new_n12684_));
  NAND3_X1   g12393(.A1(new_n12683_), .A2(new_n12684_), .A3(new_n12680_), .ZN(new_n12685_));
  NAND2_X1   g12394(.A1(new_n12685_), .A2(new_n12682_), .ZN(new_n12686_));
  NAND3_X1   g12395(.A1(new_n12686_), .A2(new_n12281_), .A3(new_n12272_), .ZN(new_n12687_));
  NOR2_X1    g12396(.A1(new_n12672_), .A2(new_n12676_), .ZN(new_n12688_));
  NOR2_X1    g12397(.A1(new_n12257_), .A2(new_n12261_), .ZN(new_n12689_));
  INV_X1     g12398(.I(new_n12689_), .ZN(new_n12690_));
  AOI21_X1   g12399(.A1(new_n12687_), .A2(new_n12690_), .B(new_n12284_), .ZN(new_n12691_));
  AOI21_X1   g12400(.A1(new_n12683_), .A2(new_n12684_), .B(new_n12680_), .ZN(new_n12692_));
  NOR3_X1    g12401(.A1(new_n12672_), .A2(new_n12676_), .A3(new_n12681_), .ZN(new_n12693_));
  NOR2_X1    g12402(.A1(new_n12692_), .A2(new_n12693_), .ZN(new_n12694_));
  NOR3_X1    g12403(.A1(new_n12694_), .A2(new_n12262_), .A3(new_n12287_), .ZN(new_n12695_));
  NOR3_X1    g12404(.A1(new_n12695_), .A2(new_n12266_), .A3(new_n12689_), .ZN(new_n12696_));
  OAI22_X1   g12405(.A1(new_n7619_), .A2(new_n861_), .B1(new_n930_), .B2(new_n8309_), .ZN(new_n12697_));
  OAI21_X1   g12406(.A1(new_n780_), .A2(new_n7947_), .B(new_n12697_), .ZN(new_n12698_));
  AOI21_X1   g12407(.A1(new_n12698_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n12699_));
  XNOR2_X1   g12408(.A1(new_n937_), .A2(new_n12699_), .ZN(new_n12700_));
  NOR3_X1    g12409(.A1(new_n12696_), .A2(new_n12691_), .A3(new_n12700_), .ZN(new_n12701_));
  OAI21_X1   g12410(.A1(new_n12695_), .A2(new_n12689_), .B(new_n12266_), .ZN(new_n12702_));
  NAND3_X1   g12411(.A1(new_n12687_), .A2(new_n12284_), .A3(new_n12690_), .ZN(new_n12703_));
  INV_X1     g12412(.I(new_n12700_), .ZN(new_n12704_));
  AOI21_X1   g12413(.A1(new_n12702_), .A2(new_n12703_), .B(new_n12704_), .ZN(new_n12705_));
  NOR2_X1    g12414(.A1(new_n12701_), .A2(new_n12705_), .ZN(new_n12706_));
  NOR3_X1    g12415(.A1(new_n12628_), .A2(new_n12626_), .A3(new_n12706_), .ZN(new_n12707_));
  OAI21_X1   g12416(.A1(new_n12189_), .A2(new_n12192_), .B(new_n12314_), .ZN(new_n12708_));
  NAND3_X1   g12417(.A1(new_n12702_), .A2(new_n12703_), .A3(new_n12704_), .ZN(new_n12709_));
  OAI21_X1   g12418(.A1(new_n12696_), .A2(new_n12691_), .B(new_n12700_), .ZN(new_n12710_));
  NAND2_X1   g12419(.A1(new_n12710_), .A2(new_n12709_), .ZN(new_n12711_));
  AOI21_X1   g12420(.A1(new_n12708_), .A2(new_n12313_), .B(new_n12711_), .ZN(new_n12712_));
  OAI21_X1   g12421(.A1(new_n12712_), .A2(new_n12707_), .B(new_n12625_), .ZN(new_n12713_));
  NAND3_X1   g12422(.A1(new_n12708_), .A2(new_n12313_), .A3(new_n12711_), .ZN(new_n12714_));
  OAI21_X1   g12423(.A1(new_n12628_), .A2(new_n12626_), .B(new_n12706_), .ZN(new_n12715_));
  NAND3_X1   g12424(.A1(new_n12714_), .A2(new_n12715_), .A3(new_n12624_), .ZN(new_n12716_));
  AOI21_X1   g12425(.A1(new_n12713_), .A2(new_n12716_), .B(new_n12622_), .ZN(new_n12717_));
  AOI21_X1   g12426(.A1(new_n12714_), .A2(new_n12715_), .B(new_n12624_), .ZN(new_n12718_));
  NOR3_X1    g12427(.A1(new_n12712_), .A2(new_n12707_), .A3(new_n12625_), .ZN(new_n12719_));
  NOR3_X1    g12428(.A1(new_n12718_), .A2(new_n12719_), .A3(new_n12621_), .ZN(new_n12720_));
  OAI22_X1   g12429(.A1(new_n5993_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n5991_), .ZN(new_n12721_));
  OAI21_X1   g12430(.A1(new_n1294_), .A2(new_n5997_), .B(new_n12721_), .ZN(new_n12722_));
  AOI21_X1   g12431(.A1(new_n12722_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n12723_));
  XOR2_X1    g12432(.A1(new_n1530_), .A2(new_n12723_), .Z(new_n12724_));
  INV_X1     g12433(.I(new_n12724_), .ZN(new_n12725_));
  OAI21_X1   g12434(.A1(new_n12720_), .A2(new_n12717_), .B(new_n12725_), .ZN(new_n12726_));
  OAI21_X1   g12435(.A1(new_n12718_), .A2(new_n12719_), .B(new_n12621_), .ZN(new_n12727_));
  NAND3_X1   g12436(.A1(new_n12713_), .A2(new_n12716_), .A3(new_n12622_), .ZN(new_n12728_));
  NAND3_X1   g12437(.A1(new_n12727_), .A2(new_n12728_), .A3(new_n12724_), .ZN(new_n12729_));
  AOI21_X1   g12438(.A1(new_n12726_), .A2(new_n12729_), .B(new_n12617_), .ZN(new_n12730_));
  OAI22_X1   g12439(.A1(new_n12615_), .A2(new_n12186_), .B1(new_n11933_), .B2(new_n12612_), .ZN(new_n12731_));
  NAND3_X1   g12440(.A1(new_n12727_), .A2(new_n12728_), .A3(new_n12725_), .ZN(new_n12732_));
  OAI21_X1   g12441(.A1(new_n12720_), .A2(new_n12717_), .B(new_n12724_), .ZN(new_n12733_));
  AOI21_X1   g12442(.A1(new_n12733_), .A2(new_n12732_), .B(new_n12731_), .ZN(new_n12734_));
  OAI22_X1   g12443(.A1(new_n5420_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n5107_), .ZN(new_n12735_));
  OAI21_X1   g12444(.A1(new_n1634_), .A2(new_n5112_), .B(new_n12735_), .ZN(new_n12736_));
  AOI21_X1   g12445(.A1(new_n12736_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n12737_));
  XNOR2_X1   g12446(.A1(new_n1940_), .A2(new_n12737_), .ZN(new_n12738_));
  NOR3_X1    g12447(.A1(new_n12730_), .A2(new_n12734_), .A3(new_n12738_), .ZN(new_n12739_));
  AOI21_X1   g12448(.A1(new_n12727_), .A2(new_n12728_), .B(new_n12724_), .ZN(new_n12740_));
  NOR3_X1    g12449(.A1(new_n12720_), .A2(new_n12717_), .A3(new_n12725_), .ZN(new_n12741_));
  OAI21_X1   g12450(.A1(new_n12741_), .A2(new_n12740_), .B(new_n12731_), .ZN(new_n12742_));
  NOR3_X1    g12451(.A1(new_n12720_), .A2(new_n12717_), .A3(new_n12724_), .ZN(new_n12743_));
  AOI21_X1   g12452(.A1(new_n12727_), .A2(new_n12728_), .B(new_n12725_), .ZN(new_n12744_));
  OAI21_X1   g12453(.A1(new_n12743_), .A2(new_n12744_), .B(new_n12617_), .ZN(new_n12745_));
  INV_X1     g12454(.I(new_n12738_), .ZN(new_n12746_));
  AOI21_X1   g12455(.A1(new_n12742_), .A2(new_n12745_), .B(new_n12746_), .ZN(new_n12747_));
  NOR2_X1    g12456(.A1(new_n12747_), .A2(new_n12739_), .ZN(new_n12748_));
  NAND2_X1   g12457(.A1(new_n12338_), .A2(new_n12332_), .ZN(new_n12749_));
  OAI22_X1   g12458(.A1(new_n12338_), .A2(new_n12332_), .B1(new_n12324_), .B2(new_n12327_), .ZN(new_n12750_));
  OAI22_X1   g12459(.A1(new_n4072_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n4067_), .ZN(new_n12751_));
  OAI21_X1   g12460(.A1(new_n2102_), .A2(new_n4318_), .B(new_n12751_), .ZN(new_n12752_));
  AOI21_X1   g12461(.A1(new_n12752_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n12753_));
  XNOR2_X1   g12462(.A1(new_n2443_), .A2(new_n12753_), .ZN(new_n12754_));
  INV_X1     g12463(.I(new_n12754_), .ZN(new_n12755_));
  NAND3_X1   g12464(.A1(new_n12750_), .A2(new_n12749_), .A3(new_n12755_), .ZN(new_n12756_));
  AOI21_X1   g12465(.A1(new_n12750_), .A2(new_n12749_), .B(new_n12755_), .ZN(new_n12757_));
  INV_X1     g12466(.I(new_n12757_), .ZN(new_n12758_));
  AOI21_X1   g12467(.A1(new_n12758_), .A2(new_n12756_), .B(new_n12748_), .ZN(new_n12759_));
  OR2_X2     g12468(.A1(new_n12747_), .A2(new_n12739_), .Z(new_n12760_));
  AOI21_X1   g12469(.A1(new_n11962_), .A2(new_n11951_), .B(new_n11963_), .ZN(new_n12761_));
  NOR2_X1    g12470(.A1(new_n12761_), .A2(new_n12331_), .ZN(new_n12762_));
  NOR2_X1    g12471(.A1(new_n12327_), .A2(new_n12324_), .ZN(new_n12763_));
  AOI21_X1   g12472(.A1(new_n12761_), .A2(new_n12331_), .B(new_n12763_), .ZN(new_n12764_));
  OAI21_X1   g12473(.A1(new_n12764_), .A2(new_n12762_), .B(new_n12755_), .ZN(new_n12765_));
  NAND3_X1   g12474(.A1(new_n12750_), .A2(new_n12749_), .A3(new_n12754_), .ZN(new_n12766_));
  AOI21_X1   g12475(.A1(new_n12765_), .A2(new_n12766_), .B(new_n12760_), .ZN(new_n12767_));
  NOR2_X1    g12476(.A1(new_n12759_), .A2(new_n12767_), .ZN(new_n12768_));
  INV_X1     g12477(.I(new_n12342_), .ZN(new_n12769_));
  NAND3_X1   g12478(.A1(new_n11948_), .A2(new_n11821_), .A3(new_n11953_), .ZN(new_n12770_));
  NAND2_X1   g12479(.A1(new_n12770_), .A2(new_n11967_), .ZN(new_n12771_));
  NOR2_X1    g12480(.A1(new_n12771_), .A2(new_n12347_), .ZN(new_n12772_));
  OAI21_X1   g12481(.A1(new_n12772_), .A2(new_n12350_), .B(new_n12769_), .ZN(new_n12773_));
  OAI21_X1   g12482(.A1(new_n11961_), .A2(new_n11966_), .B(new_n11822_), .ZN(new_n12774_));
  NAND4_X1   g12483(.A1(new_n12770_), .A2(new_n11562_), .A3(new_n11382_), .A4(new_n11967_), .ZN(new_n12775_));
  NAND3_X1   g12484(.A1(new_n12775_), .A2(new_n12342_), .A3(new_n12774_), .ZN(new_n12776_));
  XOR2_X1    g12485(.A1(new_n12337_), .A2(new_n12338_), .Z(new_n12777_));
  NAND2_X1   g12486(.A1(new_n12776_), .A2(new_n12777_), .ZN(new_n12778_));
  NAND2_X1   g12487(.A1(new_n12778_), .A2(new_n12773_), .ZN(new_n12779_));
  NAND2_X1   g12488(.A1(new_n12779_), .A2(new_n12768_), .ZN(new_n12780_));
  INV_X1     g12489(.I(new_n12756_), .ZN(new_n12781_));
  OAI21_X1   g12490(.A1(new_n12781_), .A2(new_n12757_), .B(new_n12760_), .ZN(new_n12782_));
  AOI21_X1   g12491(.A1(new_n12750_), .A2(new_n12749_), .B(new_n12754_), .ZN(new_n12783_));
  NOR3_X1    g12492(.A1(new_n12764_), .A2(new_n12762_), .A3(new_n12755_), .ZN(new_n12784_));
  OAI21_X1   g12493(.A1(new_n12783_), .A2(new_n12784_), .B(new_n12748_), .ZN(new_n12785_));
  NAND2_X1   g12494(.A1(new_n12782_), .A2(new_n12785_), .ZN(new_n12786_));
  AOI21_X1   g12495(.A1(new_n12775_), .A2(new_n12774_), .B(new_n12342_), .ZN(new_n12787_));
  AOI21_X1   g12496(.A1(new_n12776_), .A2(new_n12777_), .B(new_n12787_), .ZN(new_n12788_));
  NAND2_X1   g12497(.A1(new_n12786_), .A2(new_n12788_), .ZN(new_n12789_));
  NAND2_X1   g12498(.A1(new_n12780_), .A2(new_n12789_), .ZN(new_n12790_));
  OAI21_X1   g12499(.A1(new_n11971_), .A2(new_n11972_), .B(new_n11821_), .ZN(new_n12791_));
  NAND3_X1   g12500(.A1(new_n11959_), .A2(new_n11969_), .A3(new_n11822_), .ZN(new_n12792_));
  NAND2_X1   g12501(.A1(new_n12791_), .A2(new_n12792_), .ZN(new_n12793_));
  NAND4_X1   g12502(.A1(new_n12793_), .A2(new_n11577_), .A3(new_n11575_), .A4(new_n11818_), .ZN(new_n12794_));
  AOI21_X1   g12503(.A1(new_n11804_), .A2(new_n11818_), .B(new_n12793_), .ZN(new_n12795_));
  INV_X1     g12504(.I(new_n12183_), .ZN(new_n12796_));
  OAI21_X1   g12505(.A1(new_n12795_), .A2(new_n12796_), .B(new_n12794_), .ZN(new_n12797_));
  NAND2_X1   g12506(.A1(new_n12797_), .A2(new_n12358_), .ZN(new_n12798_));
  XNOR2_X1   g12507(.A1(new_n12346_), .A2(new_n12352_), .ZN(new_n12799_));
  OAI21_X1   g12508(.A1(new_n12797_), .A2(new_n12358_), .B(new_n12799_), .ZN(new_n12800_));
  OAI22_X1   g12509(.A1(new_n3709_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n3717_), .ZN(new_n12801_));
  OAI21_X1   g12510(.A1(new_n3260_), .A2(new_n2884_), .B(new_n12801_), .ZN(new_n12802_));
  AOI21_X1   g12511(.A1(new_n12802_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n12803_));
  XOR2_X1    g12512(.A1(new_n3722_), .A2(new_n12803_), .Z(new_n12804_));
  INV_X1     g12513(.I(new_n12804_), .ZN(new_n12805_));
  NAND3_X1   g12514(.A1(new_n12800_), .A2(new_n12798_), .A3(new_n12805_), .ZN(new_n12806_));
  NOR2_X1    g12515(.A1(new_n12184_), .A2(new_n12356_), .ZN(new_n12807_));
  XOR2_X1    g12516(.A1(new_n12346_), .A2(new_n12352_), .Z(new_n12808_));
  AOI21_X1   g12517(.A1(new_n12184_), .A2(new_n12356_), .B(new_n12808_), .ZN(new_n12809_));
  OAI21_X1   g12518(.A1(new_n12809_), .A2(new_n12807_), .B(new_n12804_), .ZN(new_n12810_));
  AOI21_X1   g12519(.A1(new_n12806_), .A2(new_n12810_), .B(new_n12790_), .ZN(new_n12811_));
  NOR2_X1    g12520(.A1(new_n12786_), .A2(new_n12788_), .ZN(new_n12812_));
  NOR2_X1    g12521(.A1(new_n12779_), .A2(new_n12768_), .ZN(new_n12813_));
  NOR2_X1    g12522(.A1(new_n12813_), .A2(new_n12812_), .ZN(new_n12814_));
  NOR3_X1    g12523(.A1(new_n12809_), .A2(new_n12807_), .A3(new_n12804_), .ZN(new_n12815_));
  AOI21_X1   g12524(.A1(new_n12800_), .A2(new_n12798_), .B(new_n12805_), .ZN(new_n12816_));
  NOR3_X1    g12525(.A1(new_n12816_), .A2(new_n12815_), .A3(new_n12814_), .ZN(new_n12817_));
  OAI21_X1   g12526(.A1(new_n12811_), .A2(new_n12817_), .B(new_n12610_), .ZN(new_n12818_));
  INV_X1     g12527(.I(new_n12610_), .ZN(new_n12819_));
  OAI21_X1   g12528(.A1(new_n12816_), .A2(new_n12815_), .B(new_n12814_), .ZN(new_n12820_));
  NAND3_X1   g12529(.A1(new_n12806_), .A2(new_n12810_), .A3(new_n12790_), .ZN(new_n12821_));
  NAND3_X1   g12530(.A1(new_n12820_), .A2(new_n12821_), .A3(new_n12819_), .ZN(new_n12822_));
  AOI22_X1   g12531(.A1(new_n12606_), .A2(new_n12601_), .B1(new_n12818_), .B2(new_n12822_), .ZN(new_n12823_));
  AOI22_X1   g12532(.A1(new_n12371_), .A2(new_n12369_), .B1(new_n12361_), .B2(new_n12365_), .ZN(new_n12824_));
  NAND2_X1   g12533(.A1(new_n12818_), .A2(new_n12822_), .ZN(new_n12825_));
  NOR3_X1    g12534(.A1(new_n12825_), .A2(new_n12600_), .A3(new_n12824_), .ZN(new_n12826_));
  OAI22_X1   g12535(.A1(new_n2171_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n2166_), .ZN(new_n12827_));
  OAI21_X1   g12536(.A1(new_n3989_), .A2(new_n2322_), .B(new_n12827_), .ZN(new_n12828_));
  AOI21_X1   g12537(.A1(new_n12828_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n12829_));
  XOR2_X1    g12538(.A1(new_n4499_), .A2(new_n12829_), .Z(new_n12830_));
  NOR3_X1    g12539(.A1(new_n12826_), .A2(new_n12823_), .A3(new_n12830_), .ZN(new_n12831_));
  AOI21_X1   g12540(.A1(new_n12820_), .A2(new_n12821_), .B(new_n12819_), .ZN(new_n12832_));
  NOR3_X1    g12541(.A1(new_n12811_), .A2(new_n12817_), .A3(new_n12610_), .ZN(new_n12833_));
  OAI22_X1   g12542(.A1(new_n12824_), .A2(new_n12600_), .B1(new_n12832_), .B2(new_n12833_), .ZN(new_n12834_));
  NAND4_X1   g12543(.A1(new_n12606_), .A2(new_n12601_), .A3(new_n12818_), .A4(new_n12822_), .ZN(new_n12835_));
  INV_X1     g12544(.I(new_n12830_), .ZN(new_n12836_));
  AOI21_X1   g12545(.A1(new_n12834_), .A2(new_n12835_), .B(new_n12836_), .ZN(new_n12837_));
  NOR3_X1    g12546(.A1(new_n12831_), .A2(new_n12837_), .A3(new_n12599_), .ZN(new_n12838_));
  NOR3_X1    g12547(.A1(new_n12838_), .A2(new_n12403_), .A3(new_n12396_), .ZN(new_n12839_));
  AOI21_X1   g12548(.A1(new_n12369_), .A2(new_n12371_), .B(new_n12399_), .ZN(new_n12840_));
  NOR2_X1    g12549(.A1(new_n12372_), .A2(new_n12366_), .ZN(new_n12841_));
  OAI21_X1   g12550(.A1(new_n12840_), .A2(new_n12841_), .B(new_n12376_), .ZN(new_n12842_));
  NAND3_X1   g12551(.A1(new_n12834_), .A2(new_n12835_), .A3(new_n12836_), .ZN(new_n12843_));
  OAI21_X1   g12552(.A1(new_n12826_), .A2(new_n12823_), .B(new_n12830_), .ZN(new_n12844_));
  NAND3_X1   g12553(.A1(new_n12844_), .A2(new_n12843_), .A3(new_n12842_), .ZN(new_n12845_));
  AOI21_X1   g12554(.A1(new_n12845_), .A2(new_n12387_), .B(new_n12383_), .ZN(new_n12846_));
  OAI22_X1   g12555(.A1(new_n1712_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n1707_), .ZN(new_n12847_));
  OAI21_X1   g12556(.A1(new_n4774_), .A2(new_n1850_), .B(new_n12847_), .ZN(new_n12848_));
  AOI21_X1   g12557(.A1(new_n12848_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n12849_));
  XNOR2_X1   g12558(.A1(new_n5357_), .A2(new_n12849_), .ZN(new_n12850_));
  NOR3_X1    g12559(.A1(new_n12839_), .A2(new_n12846_), .A3(new_n12850_), .ZN(new_n12851_));
  NAND3_X1   g12560(.A1(new_n12845_), .A2(new_n12383_), .A3(new_n12387_), .ZN(new_n12852_));
  OAI21_X1   g12561(.A1(new_n12838_), .A2(new_n12396_), .B(new_n12403_), .ZN(new_n12853_));
  INV_X1     g12562(.I(new_n12850_), .ZN(new_n12854_));
  AOI21_X1   g12563(.A1(new_n12853_), .A2(new_n12852_), .B(new_n12854_), .ZN(new_n12855_));
  NOR3_X1    g12564(.A1(new_n12851_), .A2(new_n12855_), .A3(new_n12596_), .ZN(new_n12856_));
  NOR3_X1    g12565(.A1(new_n12856_), .A2(new_n12407_), .A3(new_n12417_), .ZN(new_n12857_));
  NOR2_X1    g12566(.A1(new_n12396_), .A2(new_n12403_), .ZN(new_n12858_));
  NOR2_X1    g12567(.A1(new_n12387_), .A2(new_n12383_), .ZN(new_n12859_));
  OAI21_X1   g12568(.A1(new_n12858_), .A2(new_n12859_), .B(new_n12391_), .ZN(new_n12860_));
  NAND3_X1   g12569(.A1(new_n12853_), .A2(new_n12852_), .A3(new_n12854_), .ZN(new_n12861_));
  OAI21_X1   g12570(.A1(new_n12839_), .A2(new_n12846_), .B(new_n12850_), .ZN(new_n12862_));
  NAND3_X1   g12571(.A1(new_n12862_), .A2(new_n12861_), .A3(new_n12860_), .ZN(new_n12863_));
  AOI21_X1   g12572(.A1(new_n12863_), .A2(new_n12412_), .B(new_n12174_), .ZN(new_n12864_));
  OAI22_X1   g12573(.A1(new_n1347_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n1344_), .ZN(new_n12865_));
  OAI21_X1   g12574(.A1(new_n5913_), .A2(new_n1457_), .B(new_n12865_), .ZN(new_n12866_));
  AOI21_X1   g12575(.A1(new_n12866_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n12867_));
  XOR2_X1    g12576(.A1(new_n6233_), .A2(new_n12867_), .Z(new_n12868_));
  NOR3_X1    g12577(.A1(new_n12857_), .A2(new_n12864_), .A3(new_n12868_), .ZN(new_n12869_));
  NAND3_X1   g12578(.A1(new_n12863_), .A2(new_n12412_), .A3(new_n12174_), .ZN(new_n12870_));
  OAI21_X1   g12579(.A1(new_n12856_), .A2(new_n12407_), .B(new_n12417_), .ZN(new_n12871_));
  INV_X1     g12580(.I(new_n12868_), .ZN(new_n12872_));
  AOI21_X1   g12581(.A1(new_n12871_), .A2(new_n12870_), .B(new_n12872_), .ZN(new_n12873_));
  NOR2_X1    g12582(.A1(new_n12869_), .A2(new_n12873_), .ZN(new_n12874_));
  AOI21_X1   g12583(.A1(new_n12593_), .A2(new_n12589_), .B(new_n12874_), .ZN(new_n12875_));
  NOR2_X1    g12584(.A1(new_n12177_), .A2(new_n12175_), .ZN(new_n12876_));
  AOI21_X1   g12585(.A1(new_n12876_), .A2(new_n12169_), .B(new_n12591_), .ZN(new_n12877_));
  OAI21_X1   g12586(.A1(new_n12857_), .A2(new_n12864_), .B(new_n12872_), .ZN(new_n12878_));
  NAND3_X1   g12587(.A1(new_n12871_), .A2(new_n12870_), .A3(new_n12868_), .ZN(new_n12879_));
  AND2_X2    g12588(.A1(new_n12878_), .A2(new_n12879_), .Z(new_n12880_));
  NOR3_X1    g12589(.A1(new_n12877_), .A2(new_n12880_), .A3(new_n12588_), .ZN(new_n12881_));
  OAI22_X1   g12590(.A1(new_n1055_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n1061_), .ZN(new_n12882_));
  OAI21_X1   g12591(.A1(new_n6538_), .A2(new_n1332_), .B(new_n12882_), .ZN(new_n12883_));
  AOI21_X1   g12592(.A1(new_n12883_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n12884_));
  XNOR2_X1   g12593(.A1(new_n7202_), .A2(new_n12884_), .ZN(new_n12885_));
  INV_X1     g12594(.I(new_n12885_), .ZN(new_n12886_));
  OAI21_X1   g12595(.A1(new_n12881_), .A2(new_n12875_), .B(new_n12886_), .ZN(new_n12887_));
  NAND3_X1   g12596(.A1(new_n12871_), .A2(new_n12870_), .A3(new_n12872_), .ZN(new_n12888_));
  OAI21_X1   g12597(.A1(new_n12857_), .A2(new_n12864_), .B(new_n12868_), .ZN(new_n12889_));
  NAND2_X1   g12598(.A1(new_n12889_), .A2(new_n12888_), .ZN(new_n12890_));
  OAI21_X1   g12599(.A1(new_n12877_), .A2(new_n12588_), .B(new_n12890_), .ZN(new_n12891_));
  NAND2_X1   g12600(.A1(new_n12878_), .A2(new_n12879_), .ZN(new_n12892_));
  NAND3_X1   g12601(.A1(new_n12593_), .A2(new_n12589_), .A3(new_n12892_), .ZN(new_n12893_));
  NAND3_X1   g12602(.A1(new_n12891_), .A2(new_n12893_), .A3(new_n12885_), .ZN(new_n12894_));
  OAI22_X1   g12603(.A1(new_n970_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n820_), .ZN(new_n12895_));
  OAI21_X1   g12604(.A1(new_n7864_), .A2(new_n894_), .B(new_n12895_), .ZN(new_n12896_));
  AOI21_X1   g12605(.A1(new_n12896_), .A2(new_n827_), .B(new_n970_), .ZN(new_n12897_));
  XOR2_X1    g12606(.A1(new_n8217_), .A2(new_n12897_), .Z(new_n12898_));
  INV_X1     g12607(.I(new_n12898_), .ZN(new_n12899_));
  NAND3_X1   g12608(.A1(new_n12887_), .A2(new_n12894_), .A3(new_n12899_), .ZN(new_n12900_));
  INV_X1     g12609(.I(new_n12900_), .ZN(new_n12901_));
  AOI21_X1   g12610(.A1(new_n12887_), .A2(new_n12894_), .B(new_n12899_), .ZN(new_n12902_));
  OAI21_X1   g12611(.A1(new_n12901_), .A2(new_n12902_), .B(new_n12587_), .ZN(new_n12903_));
  AOI21_X1   g12612(.A1(new_n12165_), .A2(new_n12447_), .B(new_n12429_), .ZN(new_n12904_));
  AOI21_X1   g12613(.A1(new_n12891_), .A2(new_n12893_), .B(new_n12885_), .ZN(new_n12905_));
  NOR3_X1    g12614(.A1(new_n12881_), .A2(new_n12875_), .A3(new_n12886_), .ZN(new_n12906_));
  OAI21_X1   g12615(.A1(new_n12906_), .A2(new_n12905_), .B(new_n12899_), .ZN(new_n12907_));
  NAND3_X1   g12616(.A1(new_n12887_), .A2(new_n12894_), .A3(new_n12898_), .ZN(new_n12908_));
  NAND2_X1   g12617(.A1(new_n12907_), .A2(new_n12908_), .ZN(new_n12909_));
  NAND2_X1   g12618(.A1(new_n12909_), .A2(new_n12904_), .ZN(new_n12910_));
  NAND2_X1   g12619(.A1(new_n12910_), .A2(new_n12903_), .ZN(new_n12911_));
  NAND3_X1   g12620(.A1(new_n12911_), .A2(new_n12586_), .A3(new_n12459_), .ZN(new_n12912_));
  NAND2_X1   g12621(.A1(new_n12447_), .A2(new_n12165_), .ZN(new_n12913_));
  OAI21_X1   g12622(.A1(new_n12906_), .A2(new_n12905_), .B(new_n12898_), .ZN(new_n12914_));
  AOI22_X1   g12623(.A1(new_n12913_), .A2(new_n12446_), .B1(new_n12914_), .B2(new_n12900_), .ZN(new_n12915_));
  AOI21_X1   g12624(.A1(new_n12907_), .A2(new_n12908_), .B(new_n12587_), .ZN(new_n12916_));
  NOR2_X1    g12625(.A1(new_n12916_), .A2(new_n12915_), .ZN(new_n12917_));
  NAND2_X1   g12626(.A1(new_n12458_), .A2(new_n12444_), .ZN(new_n12918_));
  AOI21_X1   g12627(.A1(new_n12912_), .A2(new_n12918_), .B(new_n12457_), .ZN(new_n12919_));
  NAND3_X1   g12628(.A1(new_n12912_), .A2(new_n12457_), .A3(new_n12918_), .ZN(new_n12920_));
  INV_X1     g12629(.I(new_n12920_), .ZN(new_n12921_));
  OAI22_X1   g12630(.A1(new_n607_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n610_), .ZN(new_n12922_));
  OAI21_X1   g12631(.A1(new_n8563_), .A2(new_n684_), .B(new_n12922_), .ZN(new_n12923_));
  AOI21_X1   g12632(.A1(new_n12923_), .A2(new_n612_), .B(new_n607_), .ZN(new_n12924_));
  XNOR2_X1   g12633(.A1(new_n9299_), .A2(new_n12924_), .ZN(new_n12925_));
  INV_X1     g12634(.I(new_n12925_), .ZN(new_n12926_));
  OAI21_X1   g12635(.A1(new_n12921_), .A2(new_n12919_), .B(new_n12926_), .ZN(new_n12927_));
  INV_X1     g12636(.I(new_n12919_), .ZN(new_n12928_));
  NAND3_X1   g12637(.A1(new_n12928_), .A2(new_n12920_), .A3(new_n12925_), .ZN(new_n12929_));
  AOI22_X1   g12638(.A1(new_n12585_), .A2(new_n12584_), .B1(new_n12927_), .B2(new_n12929_), .ZN(new_n12930_));
  NOR2_X1    g12639(.A1(new_n12469_), .A2(new_n12467_), .ZN(new_n12931_));
  OAI21_X1   g12640(.A1(new_n12493_), .A2(new_n12931_), .B(new_n12584_), .ZN(new_n12932_));
  NOR3_X1    g12641(.A1(new_n12921_), .A2(new_n12919_), .A3(new_n12925_), .ZN(new_n12933_));
  AOI21_X1   g12642(.A1(new_n12928_), .A2(new_n12920_), .B(new_n12926_), .ZN(new_n12934_));
  NOR2_X1    g12643(.A1(new_n12934_), .A2(new_n12933_), .ZN(new_n12935_));
  NOR2_X1    g12644(.A1(new_n12932_), .A2(new_n12935_), .ZN(new_n12936_));
  OAI22_X1   g12645(.A1(new_n448_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n450_), .ZN(new_n12937_));
  OAI21_X1   g12646(.A1(new_n10025_), .A2(new_n496_), .B(new_n12937_), .ZN(new_n12938_));
  AOI21_X1   g12647(.A1(new_n12938_), .A2(new_n452_), .B(new_n448_), .ZN(new_n12939_));
  XOR2_X1    g12648(.A1(new_n10476_), .A2(new_n12939_), .Z(new_n12940_));
  NOR3_X1    g12649(.A1(new_n12930_), .A2(new_n12936_), .A3(new_n12940_), .ZN(new_n12941_));
  NAND2_X1   g12650(.A1(new_n12929_), .A2(new_n12927_), .ZN(new_n12942_));
  NAND2_X1   g12651(.A1(new_n12932_), .A2(new_n12942_), .ZN(new_n12943_));
  NAND3_X1   g12652(.A1(new_n12928_), .A2(new_n12920_), .A3(new_n12926_), .ZN(new_n12944_));
  OAI21_X1   g12653(.A1(new_n12921_), .A2(new_n12919_), .B(new_n12925_), .ZN(new_n12945_));
  NAND2_X1   g12654(.A1(new_n12944_), .A2(new_n12945_), .ZN(new_n12946_));
  NAND3_X1   g12655(.A1(new_n12585_), .A2(new_n12946_), .A3(new_n12584_), .ZN(new_n12947_));
  INV_X1     g12656(.I(new_n12940_), .ZN(new_n12948_));
  AOI21_X1   g12657(.A1(new_n12947_), .A2(new_n12943_), .B(new_n12948_), .ZN(new_n12949_));
  OAI21_X1   g12658(.A1(new_n12580_), .A2(new_n12581_), .B(new_n12483_), .ZN(new_n12950_));
  OAI21_X1   g12659(.A1(new_n12479_), .A2(new_n12475_), .B(new_n12471_), .ZN(new_n12951_));
  NAND2_X1   g12660(.A1(new_n12489_), .A2(new_n12493_), .ZN(new_n12952_));
  NAND3_X1   g12661(.A1(new_n12952_), .A2(new_n12951_), .A3(new_n12484_), .ZN(new_n12953_));
  NAND2_X1   g12662(.A1(new_n12950_), .A2(new_n12953_), .ZN(new_n12954_));
  OAI21_X1   g12663(.A1(new_n12941_), .A2(new_n12949_), .B(new_n12954_), .ZN(new_n12955_));
  NOR2_X1    g12664(.A1(new_n12955_), .A2(new_n12583_), .ZN(new_n12956_));
  NAND3_X1   g12665(.A1(new_n12947_), .A2(new_n12943_), .A3(new_n12948_), .ZN(new_n12957_));
  OAI21_X1   g12666(.A1(new_n12930_), .A2(new_n12936_), .B(new_n12940_), .ZN(new_n12958_));
  NAND2_X1   g12667(.A1(new_n12958_), .A2(new_n12957_), .ZN(new_n12959_));
  NOR2_X1    g12668(.A1(new_n12582_), .A2(new_n12483_), .ZN(new_n12961_));
  OAI21_X1   g12669(.A1(new_n12956_), .A2(new_n12961_), .B(new_n12154_), .ZN(new_n12962_));
  INV_X1     g12670(.I(new_n12583_), .ZN(new_n12963_));
  NAND3_X1   g12671(.A1(new_n12959_), .A2(new_n12963_), .A3(new_n12954_), .ZN(new_n12964_));
  INV_X1     g12672(.I(new_n12961_), .ZN(new_n12965_));
  NAND3_X1   g12673(.A1(new_n12964_), .A2(new_n12513_), .A3(new_n12965_), .ZN(new_n12966_));
  XNOR2_X1   g12674(.A1(\b[57] ), .A2(\b[59] ), .ZN(new_n12967_));
  NOR2_X1    g12675(.A1(new_n12967_), .A2(new_n12541_), .ZN(new_n12968_));
  XOR2_X1    g12676(.A1(new_n12540_), .A2(new_n12968_), .Z(new_n12969_));
  INV_X1     g12677(.I(\b[59] ), .ZN(new_n12970_));
  OAI22_X1   g12678(.A1(new_n330_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n263_), .ZN(new_n12971_));
  OAI21_X1   g12679(.A1(new_n12536_), .A2(new_n289_), .B(new_n12971_), .ZN(new_n12972_));
  AOI21_X1   g12680(.A1(new_n12972_), .A2(new_n260_), .B(new_n426_), .ZN(new_n12973_));
  XOR2_X1    g12681(.A1(new_n12969_), .A2(new_n12973_), .Z(new_n12974_));
  OAI22_X1   g12682(.A1(new_n11738_), .A2(new_n341_), .B1(new_n404_), .B2(new_n11744_), .ZN(new_n12975_));
  OAI21_X1   g12683(.A1(new_n10862_), .A2(new_n366_), .B(new_n12975_), .ZN(new_n12976_));
  AOI21_X1   g12684(.A1(new_n12976_), .A2(new_n334_), .B(new_n341_), .ZN(new_n12977_));
  XNOR2_X1   g12685(.A1(new_n11748_), .A2(new_n12977_), .ZN(new_n12978_));
  NOR2_X1    g12686(.A1(new_n12974_), .A2(new_n12978_), .ZN(new_n12979_));
  INV_X1     g12687(.I(new_n12979_), .ZN(new_n12980_));
  INV_X1     g12688(.I(new_n12974_), .ZN(new_n12981_));
  INV_X1     g12689(.I(new_n12978_), .ZN(new_n12982_));
  NOR2_X1    g12690(.A1(new_n12981_), .A2(new_n12982_), .ZN(new_n12983_));
  INV_X1     g12691(.I(new_n12983_), .ZN(new_n12984_));
  AOI22_X1   g12692(.A1(new_n12962_), .A2(new_n12966_), .B1(new_n12980_), .B2(new_n12984_), .ZN(new_n12985_));
  AOI21_X1   g12693(.A1(new_n12964_), .A2(new_n12965_), .B(new_n12513_), .ZN(new_n12986_));
  NOR3_X1    g12694(.A1(new_n12956_), .A2(new_n12154_), .A3(new_n12961_), .ZN(new_n12987_));
  XOR2_X1    g12695(.A1(new_n12974_), .A2(new_n12982_), .Z(new_n12988_));
  NOR3_X1    g12696(.A1(new_n12987_), .A2(new_n12986_), .A3(new_n12988_), .ZN(new_n12989_));
  NOR2_X1    g12697(.A1(new_n12578_), .A2(new_n12501_), .ZN(new_n12990_));
  XOR2_X1    g12698(.A1(new_n12513_), .A2(new_n12508_), .Z(new_n12991_));
  NOR2_X1    g12699(.A1(new_n12991_), .A2(new_n12500_), .ZN(new_n12992_));
  OAI22_X1   g12700(.A1(new_n12985_), .A2(new_n12989_), .B1(new_n12990_), .B2(new_n12992_), .ZN(new_n12993_));
  NOR2_X1    g12701(.A1(new_n12993_), .A2(new_n12579_), .ZN(new_n12994_));
  OAI22_X1   g12702(.A1(new_n12987_), .A2(new_n12986_), .B1(new_n12979_), .B2(new_n12983_), .ZN(new_n12995_));
  INV_X1     g12703(.I(new_n12988_), .ZN(new_n12996_));
  NAND3_X1   g12704(.A1(new_n12962_), .A2(new_n12966_), .A3(new_n12996_), .ZN(new_n12997_));
  NAND2_X1   g12705(.A1(new_n12995_), .A2(new_n12997_), .ZN(new_n12998_));
  NOR2_X1    g12706(.A1(new_n12578_), .A2(new_n12500_), .ZN(new_n13000_));
  OAI21_X1   g12707(.A1(new_n12994_), .A2(new_n13000_), .B(new_n12577_), .ZN(new_n13001_));
  INV_X1     g12708(.I(new_n12577_), .ZN(new_n13002_));
  INV_X1     g12709(.I(new_n12579_), .ZN(new_n13003_));
  OR2_X2     g12710(.A1(new_n12990_), .A2(new_n12992_), .Z(new_n13004_));
  NAND3_X1   g12711(.A1(new_n13004_), .A2(new_n13003_), .A3(new_n12998_), .ZN(new_n13005_));
  INV_X1     g12712(.I(new_n13000_), .ZN(new_n13006_));
  NAND3_X1   g12713(.A1(new_n13005_), .A2(new_n13002_), .A3(new_n13006_), .ZN(new_n13007_));
  NAND2_X1   g12714(.A1(new_n13007_), .A2(new_n13001_), .ZN(new_n13008_));
  XOR2_X1    g12715(.A1(new_n12576_), .A2(new_n13008_), .Z(\f[59] ));
  AOI21_X1   g12716(.A1(new_n12531_), .A2(new_n12520_), .B(new_n11765_), .ZN(new_n13010_));
  NOR3_X1    g12717(.A1(new_n12518_), .A2(new_n12521_), .A3(new_n12141_), .ZN(new_n13011_));
  NOR2_X1    g12718(.A1(new_n13011_), .A2(new_n13010_), .ZN(new_n13012_));
  NOR2_X1    g12719(.A1(new_n13012_), .A2(new_n12558_), .ZN(new_n13013_));
  AOI21_X1   g12720(.A1(new_n13012_), .A2(new_n12558_), .B(new_n12550_), .ZN(new_n13014_));
  AOI21_X1   g12721(.A1(new_n12555_), .A2(new_n13014_), .B(new_n13013_), .ZN(new_n13015_));
  OAI21_X1   g12722(.A1(new_n12985_), .A2(new_n12989_), .B(new_n12991_), .ZN(new_n13016_));
  NAND2_X1   g12723(.A1(new_n13016_), .A2(new_n12500_), .ZN(new_n13017_));
  NAND3_X1   g12724(.A1(new_n12995_), .A2(new_n12997_), .A3(new_n12578_), .ZN(new_n13018_));
  NAND3_X1   g12725(.A1(new_n13017_), .A2(new_n13002_), .A3(new_n13018_), .ZN(new_n13019_));
  OAI22_X1   g12726(.A1(new_n11744_), .A2(new_n341_), .B1(new_n404_), .B2(new_n12536_), .ZN(new_n13020_));
  OAI21_X1   g12727(.A1(new_n11738_), .A2(new_n366_), .B(new_n13020_), .ZN(new_n13021_));
  AOI21_X1   g12728(.A1(new_n13021_), .A2(new_n334_), .B(new_n341_), .ZN(new_n13022_));
  XNOR2_X1   g12729(.A1(new_n12128_), .A2(new_n13022_), .ZN(new_n13023_));
  INV_X1     g12730(.I(new_n12582_), .ZN(new_n13024_));
  OAI21_X1   g12731(.A1(new_n12941_), .A2(new_n12949_), .B(new_n13024_), .ZN(new_n13025_));
  NAND2_X1   g12732(.A1(new_n13025_), .A2(new_n12483_), .ZN(new_n13026_));
  NOR3_X1    g12733(.A1(new_n12941_), .A2(new_n12949_), .A3(new_n13024_), .ZN(new_n13027_));
  NOR2_X1    g12734(.A1(new_n13027_), .A2(new_n12154_), .ZN(new_n13028_));
  AOI21_X1   g12735(.A1(new_n12932_), .A2(new_n12945_), .B(new_n12933_), .ZN(new_n13029_));
  NAND2_X1   g12736(.A1(new_n12887_), .A2(new_n12894_), .ZN(new_n13030_));
  XOR2_X1    g12737(.A1(new_n12587_), .A2(new_n13030_), .Z(new_n13031_));
  NAND2_X1   g12738(.A1(new_n13031_), .A2(new_n12898_), .ZN(new_n13032_));
  INV_X1     g12739(.I(new_n13032_), .ZN(new_n13033_));
  OAI21_X1   g12740(.A1(new_n12917_), .A2(new_n12443_), .B(new_n12460_), .ZN(new_n13034_));
  AOI21_X1   g12741(.A1(new_n12917_), .A2(new_n12443_), .B(new_n12158_), .ZN(new_n13035_));
  NAND2_X1   g12742(.A1(new_n13035_), .A2(new_n13034_), .ZN(new_n13036_));
  NAND2_X1   g12743(.A1(new_n12587_), .A2(new_n12894_), .ZN(new_n13037_));
  OAI21_X1   g12744(.A1(new_n12851_), .A2(new_n12855_), .B(new_n12596_), .ZN(new_n13038_));
  AOI21_X1   g12745(.A1(new_n13038_), .A2(new_n12407_), .B(new_n12174_), .ZN(new_n13039_));
  AOI21_X1   g12746(.A1(new_n12844_), .A2(new_n12843_), .B(new_n12842_), .ZN(new_n13040_));
  OAI21_X1   g12747(.A1(new_n13040_), .A2(new_n12387_), .B(new_n12403_), .ZN(new_n13041_));
  NOR2_X1    g12748(.A1(new_n12809_), .A2(new_n12807_), .ZN(new_n13042_));
  XOR2_X1    g12749(.A1(new_n13042_), .A2(new_n12814_), .Z(new_n13043_));
  NAND2_X1   g12750(.A1(new_n13043_), .A2(new_n12610_), .ZN(new_n13044_));
  XOR2_X1    g12751(.A1(new_n13042_), .A2(new_n12790_), .Z(new_n13045_));
  NAND2_X1   g12752(.A1(new_n13045_), .A2(new_n12819_), .ZN(new_n13046_));
  AOI21_X1   g12753(.A1(new_n13044_), .A2(new_n13046_), .B(new_n12804_), .ZN(new_n13047_));
  INV_X1     g12754(.I(new_n13047_), .ZN(new_n13048_));
  AOI21_X1   g12755(.A1(new_n12372_), .A2(new_n12605_), .B(new_n12600_), .ZN(new_n13049_));
  AOI21_X1   g12756(.A1(new_n12780_), .A2(new_n12789_), .B(new_n12610_), .ZN(new_n13050_));
  NOR3_X1    g12757(.A1(new_n12813_), .A2(new_n12812_), .A3(new_n12819_), .ZN(new_n13051_));
  NOR2_X1    g12758(.A1(new_n13051_), .A2(new_n13050_), .ZN(new_n13052_));
  NOR3_X1    g12759(.A1(new_n12809_), .A2(new_n12807_), .A3(new_n13052_), .ZN(new_n13053_));
  NAND2_X1   g12760(.A1(new_n12790_), .A2(new_n12610_), .ZN(new_n13054_));
  NOR2_X1    g12761(.A1(new_n12764_), .A2(new_n12762_), .ZN(new_n13055_));
  XOR2_X1    g12762(.A1(new_n13055_), .A2(new_n12748_), .Z(new_n13056_));
  NOR2_X1    g12763(.A1(new_n13056_), .A2(new_n12755_), .ZN(new_n13057_));
  INV_X1     g12764(.I(new_n13057_), .ZN(new_n13058_));
  NOR2_X1    g12765(.A1(new_n12779_), .A2(new_n12786_), .ZN(new_n13059_));
  NOR2_X1    g12766(.A1(new_n12741_), .A2(new_n12617_), .ZN(new_n13060_));
  NOR2_X1    g12767(.A1(new_n13060_), .A2(new_n12740_), .ZN(new_n13061_));
  NAND2_X1   g12768(.A1(new_n12708_), .A2(new_n12313_), .ZN(new_n13062_));
  NAND2_X1   g12769(.A1(new_n13062_), .A2(new_n12622_), .ZN(new_n13063_));
  XOR2_X1    g12770(.A1(new_n12711_), .A2(new_n12624_), .Z(new_n13064_));
  OAI21_X1   g12771(.A1(new_n13062_), .A2(new_n12622_), .B(new_n13064_), .ZN(new_n13065_));
  NAND2_X1   g12772(.A1(new_n13065_), .A2(new_n13063_), .ZN(new_n13066_));
  NOR2_X1    g12773(.A1(new_n12711_), .A2(new_n12624_), .ZN(new_n13067_));
  NOR2_X1    g12774(.A1(new_n12688_), .A2(new_n12681_), .ZN(new_n13068_));
  AOI21_X1   g12775(.A1(new_n12686_), .A2(new_n12280_), .B(new_n12263_), .ZN(new_n13069_));
  OAI21_X1   g12776(.A1(new_n12686_), .A2(new_n12280_), .B(new_n12284_), .ZN(new_n13070_));
  NOR3_X1    g12777(.A1(new_n12657_), .A2(new_n12662_), .A3(new_n12669_), .ZN(new_n13071_));
  INV_X1     g12778(.I(new_n13071_), .ZN(new_n13072_));
  AOI21_X1   g12779(.A1(new_n12632_), .A2(new_n12241_), .B(new_n12655_), .ZN(new_n13073_));
  NOR2_X1    g12780(.A1(new_n13073_), .A2(new_n12650_), .ZN(new_n13074_));
  NAND2_X1   g12781(.A1(\a[59] ), .A2(\a[60] ), .ZN(new_n13075_));
  OR2_X2     g12782(.A1(\a[59] ), .A2(\a[60] ), .Z(new_n13076_));
  NAND2_X1   g12783(.A1(new_n13076_), .A2(new_n13075_), .ZN(new_n13077_));
  INV_X1     g12784(.I(new_n12637_), .ZN(new_n13078_));
  AOI22_X1   g12785(.A1(new_n13078_), .A2(\b[1] ), .B1(new_n10564_), .B2(new_n12218_), .ZN(new_n13079_));
  OAI21_X1   g12786(.A1(new_n13079_), .A2(\a[59] ), .B(new_n301_), .ZN(new_n13080_));
  XOR2_X1    g12787(.A1(new_n13080_), .A2(new_n12643_), .Z(new_n13081_));
  NAND3_X1   g12788(.A1(new_n12644_), .A2(new_n13081_), .A3(new_n12633_), .ZN(new_n13082_));
  NOR2_X1    g12789(.A1(new_n13082_), .A2(new_n13077_), .ZN(new_n13083_));
  INV_X1     g12790(.I(new_n13077_), .ZN(new_n13084_));
  NAND2_X1   g12791(.A1(new_n12644_), .A2(new_n12633_), .ZN(new_n13085_));
  XOR2_X1    g12792(.A1(new_n13080_), .A2(new_n12214_), .Z(new_n13086_));
  NOR2_X1    g12793(.A1(new_n13085_), .A2(new_n13086_), .ZN(new_n13087_));
  NOR2_X1    g12794(.A1(new_n13087_), .A2(new_n13084_), .ZN(new_n13088_));
  OAI21_X1   g12795(.A1(new_n13088_), .A2(new_n13083_), .B(new_n258_), .ZN(new_n13089_));
  NAND2_X1   g12796(.A1(new_n13087_), .A2(new_n13084_), .ZN(new_n13090_));
  NAND2_X1   g12797(.A1(new_n13082_), .A2(new_n13077_), .ZN(new_n13091_));
  NAND3_X1   g12798(.A1(new_n13090_), .A2(new_n13091_), .A3(\b[0] ), .ZN(new_n13092_));
  OAI22_X1   g12799(.A1(new_n10979_), .A2(new_n421_), .B1(new_n325_), .B2(new_n11401_), .ZN(new_n13093_));
  AOI21_X1   g12800(.A1(new_n13093_), .A2(new_n10973_), .B(new_n10964_), .ZN(new_n13094_));
  XOR2_X1    g12801(.A1(new_n425_), .A2(new_n13094_), .Z(new_n13095_));
  INV_X1     g12802(.I(new_n13095_), .ZN(new_n13096_));
  NAND3_X1   g12803(.A1(new_n13089_), .A2(new_n13092_), .A3(new_n13096_), .ZN(new_n13097_));
  INV_X1     g12804(.I(new_n13089_), .ZN(new_n13098_));
  INV_X1     g12805(.I(new_n13092_), .ZN(new_n13099_));
  OAI21_X1   g12806(.A1(new_n13098_), .A2(new_n13099_), .B(new_n13095_), .ZN(new_n13100_));
  AOI21_X1   g12807(.A1(new_n13100_), .A2(new_n13097_), .B(new_n13074_), .ZN(new_n13101_));
  INV_X1     g12808(.I(new_n13074_), .ZN(new_n13102_));
  OAI21_X1   g12809(.A1(new_n13098_), .A2(new_n13099_), .B(new_n13096_), .ZN(new_n13103_));
  NAND3_X1   g12810(.A1(new_n13089_), .A2(new_n13092_), .A3(new_n13095_), .ZN(new_n13104_));
  AOI21_X1   g12811(.A1(new_n13103_), .A2(new_n13104_), .B(new_n13102_), .ZN(new_n13105_));
  AOI22_X1   g12812(.A1(new_n11415_), .A2(new_n650_), .B1(\b[7] ), .B2(new_n10145_), .ZN(new_n13106_));
  OAI21_X1   g12813(.A1(new_n13106_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n13107_));
  XOR2_X1    g12814(.A1(new_n569_), .A2(new_n13107_), .Z(new_n13108_));
  INV_X1     g12815(.I(new_n13108_), .ZN(new_n13109_));
  OAI21_X1   g12816(.A1(new_n13105_), .A2(new_n13101_), .B(new_n13109_), .ZN(new_n13110_));
  AOI21_X1   g12817(.A1(new_n12631_), .A2(new_n12675_), .B(new_n13110_), .ZN(new_n13111_));
  NAND2_X1   g12818(.A1(new_n12631_), .A2(new_n12675_), .ZN(new_n13112_));
  INV_X1     g12819(.I(new_n13101_), .ZN(new_n13113_));
  NAND2_X1   g12820(.A1(new_n13103_), .A2(new_n13104_), .ZN(new_n13114_));
  NAND2_X1   g12821(.A1(new_n13114_), .A2(new_n13074_), .ZN(new_n13115_));
  AOI21_X1   g12822(.A1(new_n13113_), .A2(new_n13115_), .B(new_n13108_), .ZN(new_n13116_));
  NOR2_X1    g12823(.A1(new_n13112_), .A2(new_n13116_), .ZN(new_n13117_));
  OAI21_X1   g12824(.A1(new_n13117_), .A2(new_n13111_), .B(new_n13072_), .ZN(new_n13118_));
  NAND2_X1   g12825(.A1(new_n13112_), .A2(new_n13116_), .ZN(new_n13119_));
  NAND3_X1   g12826(.A1(new_n13110_), .A2(new_n12631_), .A3(new_n12675_), .ZN(new_n13120_));
  NAND3_X1   g12827(.A1(new_n13119_), .A2(new_n13120_), .A3(new_n13071_), .ZN(new_n13121_));
  AOI22_X1   g12828(.A1(new_n8631_), .A2(\b[11] ), .B1(\b[12] ), .B2(new_n9382_), .ZN(new_n13122_));
  AOI21_X1   g12829(.A1(\b[10] ), .A2(new_n9731_), .B(new_n13122_), .ZN(new_n13123_));
  OAI21_X1   g12830(.A1(new_n13123_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n13124_));
  XNOR2_X1   g12831(.A1(new_n785_), .A2(new_n13124_), .ZN(new_n13125_));
  AOI21_X1   g12832(.A1(new_n13118_), .A2(new_n13121_), .B(new_n13125_), .ZN(new_n13126_));
  OAI21_X1   g12833(.A1(new_n13069_), .A2(new_n13070_), .B(new_n13126_), .ZN(new_n13127_));
  OAI21_X1   g12834(.A1(new_n12694_), .A2(new_n12257_), .B(new_n12261_), .ZN(new_n13128_));
  AOI21_X1   g12835(.A1(new_n12694_), .A2(new_n12257_), .B(new_n12266_), .ZN(new_n13129_));
  AOI21_X1   g12836(.A1(new_n13119_), .A2(new_n13120_), .B(new_n13071_), .ZN(new_n13130_));
  NOR3_X1    g12837(.A1(new_n13117_), .A2(new_n13111_), .A3(new_n13072_), .ZN(new_n13131_));
  INV_X1     g12838(.I(new_n13125_), .ZN(new_n13132_));
  OAI21_X1   g12839(.A1(new_n13131_), .A2(new_n13130_), .B(new_n13132_), .ZN(new_n13133_));
  NAND3_X1   g12840(.A1(new_n13128_), .A2(new_n13129_), .A3(new_n13133_), .ZN(new_n13134_));
  AOI21_X1   g12841(.A1(new_n13134_), .A2(new_n13127_), .B(new_n13068_), .ZN(new_n13135_));
  INV_X1     g12842(.I(new_n13068_), .ZN(new_n13136_));
  AOI21_X1   g12843(.A1(new_n13129_), .A2(new_n13128_), .B(new_n13133_), .ZN(new_n13137_));
  NOR3_X1    g12844(.A1(new_n13069_), .A2(new_n13070_), .A3(new_n13126_), .ZN(new_n13138_));
  NOR3_X1    g12845(.A1(new_n13137_), .A2(new_n13138_), .A3(new_n13136_), .ZN(new_n13139_));
  OAI22_X1   g12846(.A1(new_n7619_), .A2(new_n930_), .B1(new_n1017_), .B2(new_n8309_), .ZN(new_n13140_));
  OAI21_X1   g12847(.A1(new_n861_), .A2(new_n7947_), .B(new_n13140_), .ZN(new_n13141_));
  AOI21_X1   g12848(.A1(new_n13141_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n13142_));
  XOR2_X1    g12849(.A1(new_n1024_), .A2(new_n13142_), .Z(new_n13143_));
  INV_X1     g12850(.I(new_n13143_), .ZN(new_n13144_));
  OAI21_X1   g12851(.A1(new_n13135_), .A2(new_n13139_), .B(new_n13144_), .ZN(new_n13145_));
  NOR2_X1    g12852(.A1(new_n13067_), .A2(new_n13145_), .ZN(new_n13146_));
  OAI21_X1   g12853(.A1(new_n13137_), .A2(new_n13138_), .B(new_n13136_), .ZN(new_n13147_));
  NAND3_X1   g12854(.A1(new_n13134_), .A2(new_n13127_), .A3(new_n13068_), .ZN(new_n13148_));
  AOI21_X1   g12855(.A1(new_n13147_), .A2(new_n13148_), .B(new_n13143_), .ZN(new_n13149_));
  NOR3_X1    g12856(.A1(new_n13149_), .A2(new_n12624_), .A3(new_n12711_), .ZN(new_n13150_));
  OAI21_X1   g12857(.A1(new_n13146_), .A2(new_n13150_), .B(new_n12710_), .ZN(new_n13151_));
  OAI21_X1   g12858(.A1(new_n12624_), .A2(new_n12711_), .B(new_n13149_), .ZN(new_n13152_));
  NAND3_X1   g12859(.A1(new_n13145_), .A2(new_n12625_), .A3(new_n12706_), .ZN(new_n13153_));
  NAND3_X1   g12860(.A1(new_n13152_), .A2(new_n13153_), .A3(new_n12705_), .ZN(new_n13154_));
  OAI22_X1   g12861(.A1(new_n6644_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n6647_), .ZN(new_n13155_));
  OAI21_X1   g12862(.A1(new_n1109_), .A2(new_n7284_), .B(new_n13155_), .ZN(new_n13156_));
  AOI21_X1   g12863(.A1(new_n13156_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n13157_));
  XOR2_X1    g12864(.A1(new_n1299_), .A2(new_n13157_), .Z(new_n13158_));
  INV_X1     g12865(.I(new_n13158_), .ZN(new_n13159_));
  NAND3_X1   g12866(.A1(new_n13151_), .A2(new_n13154_), .A3(new_n13159_), .ZN(new_n13160_));
  AOI21_X1   g12867(.A1(new_n13152_), .A2(new_n13153_), .B(new_n12705_), .ZN(new_n13161_));
  NOR3_X1    g12868(.A1(new_n13146_), .A2(new_n13150_), .A3(new_n12710_), .ZN(new_n13162_));
  OAI21_X1   g12869(.A1(new_n13162_), .A2(new_n13161_), .B(new_n13158_), .ZN(new_n13163_));
  NAND2_X1   g12870(.A1(new_n13163_), .A2(new_n13160_), .ZN(new_n13164_));
  XOR2_X1    g12871(.A1(new_n13066_), .A2(new_n13164_), .Z(new_n13165_));
  OAI22_X1   g12872(.A1(new_n5993_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n5991_), .ZN(new_n13166_));
  OAI21_X1   g12873(.A1(new_n1518_), .A2(new_n5997_), .B(new_n13166_), .ZN(new_n13167_));
  AOI21_X1   g12874(.A1(new_n13167_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n13168_));
  XNOR2_X1   g12875(.A1(new_n1638_), .A2(new_n13168_), .ZN(new_n13169_));
  INV_X1     g12876(.I(new_n13169_), .ZN(new_n13170_));
  XOR2_X1    g12877(.A1(new_n13165_), .A2(new_n13170_), .Z(new_n13171_));
  NOR2_X1    g12878(.A1(new_n13165_), .A2(new_n13169_), .ZN(new_n13172_));
  XNOR2_X1   g12879(.A1(new_n13066_), .A2(new_n13164_), .ZN(new_n13173_));
  NOR2_X1    g12880(.A1(new_n13173_), .A2(new_n13170_), .ZN(new_n13174_));
  NOR2_X1    g12881(.A1(new_n13174_), .A2(new_n13172_), .ZN(new_n13175_));
  MUX2_X1    g12882(.I0(new_n13171_), .I1(new_n13175_), .S(new_n13061_), .Z(new_n13176_));
  NAND2_X1   g12883(.A1(new_n12742_), .A2(new_n12745_), .ZN(new_n13177_));
  NAND2_X1   g12884(.A1(new_n13177_), .A2(new_n12746_), .ZN(new_n13178_));
  INV_X1     g12885(.I(new_n13178_), .ZN(new_n13179_));
  NOR2_X1    g12886(.A1(new_n12730_), .A2(new_n12734_), .ZN(new_n13180_));
  AOI22_X1   g12887(.A1(new_n12750_), .A2(new_n12749_), .B1(new_n13180_), .B2(new_n12738_), .ZN(new_n13181_));
  OAI22_X1   g12888(.A1(new_n5420_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n5107_), .ZN(new_n13182_));
  OAI21_X1   g12889(.A1(new_n1803_), .A2(new_n5112_), .B(new_n13182_), .ZN(new_n13183_));
  AOI21_X1   g12890(.A1(new_n13183_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n13184_));
  XOR2_X1    g12891(.A1(new_n2106_), .A2(new_n13184_), .Z(new_n13185_));
  INV_X1     g12892(.I(new_n13185_), .ZN(new_n13186_));
  OAI21_X1   g12893(.A1(new_n13181_), .A2(new_n13179_), .B(new_n13186_), .ZN(new_n13187_));
  OAI22_X1   g12894(.A1(new_n12764_), .A2(new_n12762_), .B1(new_n13177_), .B2(new_n12746_), .ZN(new_n13188_));
  NAND3_X1   g12895(.A1(new_n13188_), .A2(new_n13178_), .A3(new_n13185_), .ZN(new_n13189_));
  AOI21_X1   g12896(.A1(new_n13187_), .A2(new_n13189_), .B(new_n13176_), .ZN(new_n13190_));
  OAI21_X1   g12897(.A1(new_n13172_), .A2(new_n13174_), .B(new_n13061_), .ZN(new_n13191_));
  OAI21_X1   g12898(.A1(new_n13061_), .A2(new_n13171_), .B(new_n13191_), .ZN(new_n13192_));
  NAND3_X1   g12899(.A1(new_n13188_), .A2(new_n13178_), .A3(new_n13186_), .ZN(new_n13193_));
  OAI21_X1   g12900(.A1(new_n13181_), .A2(new_n13179_), .B(new_n13185_), .ZN(new_n13194_));
  AOI21_X1   g12901(.A1(new_n13194_), .A2(new_n13193_), .B(new_n13192_), .ZN(new_n13195_));
  OAI22_X1   g12902(.A1(new_n2439_), .A2(new_n4072_), .B1(new_n4067_), .B2(new_n2643_), .ZN(new_n13196_));
  OAI21_X1   g12903(.A1(new_n2281_), .A2(new_n4318_), .B(new_n13196_), .ZN(new_n13197_));
  AOI21_X1   g12904(.A1(new_n13197_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n13198_));
  XOR2_X1    g12905(.A1(new_n2647_), .A2(new_n13198_), .Z(new_n13199_));
  OAI21_X1   g12906(.A1(new_n13195_), .A2(new_n13190_), .B(new_n13199_), .ZN(new_n13200_));
  NOR2_X1    g12907(.A1(new_n13059_), .A2(new_n13200_), .ZN(new_n13201_));
  NAND2_X1   g12908(.A1(new_n12768_), .A2(new_n12788_), .ZN(new_n13202_));
  AOI21_X1   g12909(.A1(new_n13188_), .A2(new_n13178_), .B(new_n13185_), .ZN(new_n13203_));
  NOR3_X1    g12910(.A1(new_n13181_), .A2(new_n13179_), .A3(new_n13186_), .ZN(new_n13204_));
  OAI21_X1   g12911(.A1(new_n13204_), .A2(new_n13203_), .B(new_n13192_), .ZN(new_n13205_));
  NOR3_X1    g12912(.A1(new_n13181_), .A2(new_n13179_), .A3(new_n13185_), .ZN(new_n13206_));
  AOI21_X1   g12913(.A1(new_n13188_), .A2(new_n13178_), .B(new_n13186_), .ZN(new_n13207_));
  OAI21_X1   g12914(.A1(new_n13206_), .A2(new_n13207_), .B(new_n13176_), .ZN(new_n13208_));
  NAND2_X1   g12915(.A1(new_n13205_), .A2(new_n13208_), .ZN(new_n13209_));
  AOI21_X1   g12916(.A1(new_n13209_), .A2(new_n13199_), .B(new_n13202_), .ZN(new_n13210_));
  OAI21_X1   g12917(.A1(new_n13210_), .A2(new_n13201_), .B(new_n13058_), .ZN(new_n13211_));
  NAND3_X1   g12918(.A1(new_n13202_), .A2(new_n13209_), .A3(new_n13199_), .ZN(new_n13212_));
  NAND2_X1   g12919(.A1(new_n13059_), .A2(new_n13200_), .ZN(new_n13213_));
  NAND3_X1   g12920(.A1(new_n13213_), .A2(new_n13212_), .A3(new_n13057_), .ZN(new_n13214_));
  NAND2_X1   g12921(.A1(new_n13211_), .A2(new_n13214_), .ZN(new_n13215_));
  OAI22_X1   g12922(.A1(new_n3018_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n3260_), .ZN(new_n13216_));
  OAI21_X1   g12923(.A1(new_n2842_), .A2(new_n3569_), .B(new_n13216_), .ZN(new_n13217_));
  AOI21_X1   g12924(.A1(new_n13217_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n13218_));
  XNOR2_X1   g12925(.A1(new_n3264_), .A2(new_n13218_), .ZN(new_n13219_));
  INV_X1     g12926(.I(new_n13219_), .ZN(new_n13220_));
  NAND3_X1   g12927(.A1(new_n13215_), .A2(new_n13054_), .A3(new_n13220_), .ZN(new_n13221_));
  INV_X1     g12928(.I(new_n13054_), .ZN(new_n13222_));
  AOI21_X1   g12929(.A1(new_n13213_), .A2(new_n13212_), .B(new_n13057_), .ZN(new_n13223_));
  NOR3_X1    g12930(.A1(new_n13210_), .A2(new_n13201_), .A3(new_n13058_), .ZN(new_n13224_));
  NOR2_X1    g12931(.A1(new_n13224_), .A2(new_n13223_), .ZN(new_n13225_));
  OAI21_X1   g12932(.A1(new_n13225_), .A2(new_n13219_), .B(new_n13222_), .ZN(new_n13226_));
  AOI21_X1   g12933(.A1(new_n13226_), .A2(new_n13221_), .B(new_n13053_), .ZN(new_n13227_));
  OAI21_X1   g12934(.A1(new_n12813_), .A2(new_n12812_), .B(new_n12819_), .ZN(new_n13228_));
  NAND3_X1   g12935(.A1(new_n12780_), .A2(new_n12789_), .A3(new_n12610_), .ZN(new_n13229_));
  NAND2_X1   g12936(.A1(new_n13228_), .A2(new_n13229_), .ZN(new_n13230_));
  NAND3_X1   g12937(.A1(new_n12800_), .A2(new_n12798_), .A3(new_n13230_), .ZN(new_n13231_));
  NOR3_X1    g12938(.A1(new_n13225_), .A2(new_n13222_), .A3(new_n13219_), .ZN(new_n13232_));
  AOI21_X1   g12939(.A1(new_n13215_), .A2(new_n13220_), .B(new_n13054_), .ZN(new_n13233_));
  NOR3_X1    g12940(.A1(new_n13232_), .A2(new_n13233_), .A3(new_n13231_), .ZN(new_n13234_));
  OAI22_X1   g12941(.A1(new_n3717_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n3989_), .ZN(new_n13235_));
  OAI21_X1   g12942(.A1(new_n3709_), .A2(new_n2884_), .B(new_n13235_), .ZN(new_n13236_));
  AOI21_X1   g12943(.A1(new_n13236_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n13237_));
  XNOR2_X1   g12944(.A1(new_n3993_), .A2(new_n13237_), .ZN(new_n13238_));
  INV_X1     g12945(.I(new_n13238_), .ZN(new_n13239_));
  OAI21_X1   g12946(.A1(new_n13234_), .A2(new_n13227_), .B(new_n13239_), .ZN(new_n13240_));
  AOI21_X1   g12947(.A1(new_n13049_), .A2(new_n12825_), .B(new_n13240_), .ZN(new_n13241_));
  NAND2_X1   g12948(.A1(new_n12606_), .A2(new_n12601_), .ZN(new_n13242_));
  NOR2_X1    g12949(.A1(new_n12833_), .A2(new_n12832_), .ZN(new_n13243_));
  INV_X1     g12950(.I(new_n13240_), .ZN(new_n13244_));
  NOR3_X1    g12951(.A1(new_n13244_), .A2(new_n13242_), .A3(new_n13243_), .ZN(new_n13245_));
  OAI21_X1   g12952(.A1(new_n13245_), .A2(new_n13241_), .B(new_n13048_), .ZN(new_n13246_));
  OAI21_X1   g12953(.A1(new_n13242_), .A2(new_n13243_), .B(new_n13244_), .ZN(new_n13247_));
  NAND3_X1   g12954(.A1(new_n13049_), .A2(new_n12825_), .A3(new_n13240_), .ZN(new_n13248_));
  NAND3_X1   g12955(.A1(new_n13247_), .A2(new_n13047_), .A3(new_n13248_), .ZN(new_n13249_));
  OAI22_X1   g12956(.A1(new_n2171_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n2166_), .ZN(new_n13250_));
  OAI21_X1   g12957(.A1(new_n4253_), .A2(new_n2322_), .B(new_n13250_), .ZN(new_n13251_));
  AOI21_X1   g12958(.A1(new_n13251_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n13252_));
  XNOR2_X1   g12959(.A1(new_n4778_), .A2(new_n13252_), .ZN(new_n13253_));
  AOI21_X1   g12960(.A1(new_n13246_), .A2(new_n13249_), .B(new_n13253_), .ZN(new_n13254_));
  NAND2_X1   g12961(.A1(new_n13041_), .A2(new_n13254_), .ZN(new_n13255_));
  OAI21_X1   g12962(.A1(new_n12831_), .A2(new_n12837_), .B(new_n12599_), .ZN(new_n13256_));
  AOI21_X1   g12963(.A1(new_n13256_), .A2(new_n12396_), .B(new_n12383_), .ZN(new_n13257_));
  AOI21_X1   g12964(.A1(new_n13247_), .A2(new_n13248_), .B(new_n13047_), .ZN(new_n13258_));
  NOR3_X1    g12965(.A1(new_n13245_), .A2(new_n13048_), .A3(new_n13241_), .ZN(new_n13259_));
  INV_X1     g12966(.I(new_n13253_), .ZN(new_n13260_));
  OAI21_X1   g12967(.A1(new_n13258_), .A2(new_n13259_), .B(new_n13260_), .ZN(new_n13261_));
  NAND2_X1   g12968(.A1(new_n13257_), .A2(new_n13261_), .ZN(new_n13262_));
  AOI21_X1   g12969(.A1(new_n13262_), .A2(new_n13255_), .B(new_n12837_), .ZN(new_n13263_));
  NOR2_X1    g12970(.A1(new_n13257_), .A2(new_n13261_), .ZN(new_n13264_));
  NOR2_X1    g12971(.A1(new_n13041_), .A2(new_n13254_), .ZN(new_n13265_));
  NOR3_X1    g12972(.A1(new_n13264_), .A2(new_n13265_), .A3(new_n12844_), .ZN(new_n13266_));
  OAI22_X1   g12973(.A1(new_n1712_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n1707_), .ZN(new_n13267_));
  OAI21_X1   g12974(.A1(new_n5068_), .A2(new_n1850_), .B(new_n13267_), .ZN(new_n13268_));
  AOI21_X1   g12975(.A1(new_n13268_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n13269_));
  XNOR2_X1   g12976(.A1(new_n5600_), .A2(new_n13269_), .ZN(new_n13270_));
  INV_X1     g12977(.I(new_n13270_), .ZN(new_n13271_));
  OAI21_X1   g12978(.A1(new_n13263_), .A2(new_n13266_), .B(new_n13271_), .ZN(new_n13272_));
  NOR2_X1    g12979(.A1(new_n13039_), .A2(new_n13272_), .ZN(new_n13273_));
  AOI21_X1   g12980(.A1(new_n12862_), .A2(new_n12861_), .B(new_n12860_), .ZN(new_n13274_));
  OAI21_X1   g12981(.A1(new_n13274_), .A2(new_n12412_), .B(new_n12417_), .ZN(new_n13275_));
  OAI21_X1   g12982(.A1(new_n13264_), .A2(new_n13265_), .B(new_n12844_), .ZN(new_n13276_));
  NAND3_X1   g12983(.A1(new_n13262_), .A2(new_n13255_), .A3(new_n12837_), .ZN(new_n13277_));
  AOI21_X1   g12984(.A1(new_n13276_), .A2(new_n13277_), .B(new_n13270_), .ZN(new_n13278_));
  NOR2_X1    g12985(.A1(new_n13275_), .A2(new_n13278_), .ZN(new_n13279_));
  OAI21_X1   g12986(.A1(new_n13273_), .A2(new_n13279_), .B(new_n12862_), .ZN(new_n13280_));
  NAND2_X1   g12987(.A1(new_n13275_), .A2(new_n13278_), .ZN(new_n13281_));
  NAND2_X1   g12988(.A1(new_n13039_), .A2(new_n13272_), .ZN(new_n13282_));
  NAND3_X1   g12989(.A1(new_n13282_), .A2(new_n13281_), .A3(new_n12855_), .ZN(new_n13283_));
  OAI22_X1   g12990(.A1(new_n1347_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n1344_), .ZN(new_n13284_));
  OAI21_X1   g12991(.A1(new_n5921_), .A2(new_n1457_), .B(new_n13284_), .ZN(new_n13285_));
  AOI21_X1   g12992(.A1(new_n13285_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n13286_));
  XOR2_X1    g12993(.A1(new_n6543_), .A2(new_n13286_), .Z(new_n13287_));
  AOI21_X1   g12994(.A1(new_n13280_), .A2(new_n13283_), .B(new_n13287_), .ZN(new_n13288_));
  NAND2_X1   g12995(.A1(new_n12893_), .A2(new_n13288_), .ZN(new_n13289_));
  AOI21_X1   g12996(.A1(new_n13282_), .A2(new_n13281_), .B(new_n12855_), .ZN(new_n13290_));
  NOR3_X1    g12997(.A1(new_n13273_), .A2(new_n13279_), .A3(new_n12862_), .ZN(new_n13291_));
  INV_X1     g12998(.I(new_n13287_), .ZN(new_n13292_));
  OAI21_X1   g12999(.A1(new_n13290_), .A2(new_n13291_), .B(new_n13292_), .ZN(new_n13293_));
  NAND4_X1   g13000(.A1(new_n13293_), .A2(new_n12589_), .A3(new_n12593_), .A4(new_n12892_), .ZN(new_n13294_));
  AOI21_X1   g13001(.A1(new_n13289_), .A2(new_n13294_), .B(new_n12873_), .ZN(new_n13295_));
  NOR2_X1    g13002(.A1(new_n12881_), .A2(new_n13293_), .ZN(new_n13296_));
  NOR2_X1    g13003(.A1(new_n12893_), .A2(new_n13288_), .ZN(new_n13297_));
  NOR3_X1    g13004(.A1(new_n13296_), .A2(new_n13297_), .A3(new_n12889_), .ZN(new_n13298_));
  OAI22_X1   g13005(.A1(new_n1055_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n1061_), .ZN(new_n13299_));
  OAI21_X1   g13006(.A1(new_n6847_), .A2(new_n1332_), .B(new_n13299_), .ZN(new_n13300_));
  AOI21_X1   g13007(.A1(new_n13300_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n13301_));
  XOR2_X1    g13008(.A1(new_n7516_), .A2(new_n13301_), .Z(new_n13302_));
  INV_X1     g13009(.I(new_n13302_), .ZN(new_n13303_));
  OAI21_X1   g13010(.A1(new_n13298_), .A2(new_n13295_), .B(new_n13303_), .ZN(new_n13304_));
  OAI21_X1   g13011(.A1(new_n13296_), .A2(new_n13297_), .B(new_n12889_), .ZN(new_n13305_));
  NAND3_X1   g13012(.A1(new_n13289_), .A2(new_n13294_), .A3(new_n12873_), .ZN(new_n13306_));
  NAND3_X1   g13013(.A1(new_n13305_), .A2(new_n13306_), .A3(new_n13302_), .ZN(new_n13307_));
  AOI22_X1   g13014(.A1(new_n13037_), .A2(new_n12887_), .B1(new_n13304_), .B2(new_n13307_), .ZN(new_n13308_));
  OAI21_X1   g13015(.A1(new_n12904_), .A2(new_n12906_), .B(new_n12887_), .ZN(new_n13309_));
  NOR3_X1    g13016(.A1(new_n13298_), .A2(new_n13295_), .A3(new_n13302_), .ZN(new_n13310_));
  AOI21_X1   g13017(.A1(new_n13305_), .A2(new_n13306_), .B(new_n13303_), .ZN(new_n13311_));
  NOR2_X1    g13018(.A1(new_n13310_), .A2(new_n13311_), .ZN(new_n13312_));
  NOR2_X1    g13019(.A1(new_n13312_), .A2(new_n13309_), .ZN(new_n13313_));
  NOR2_X1    g13020(.A1(new_n13313_), .A2(new_n13308_), .ZN(new_n13314_));
  OAI22_X1   g13021(.A1(new_n970_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n820_), .ZN(new_n13315_));
  OAI21_X1   g13022(.A1(new_n7870_), .A2(new_n894_), .B(new_n13315_), .ZN(new_n13316_));
  AOI21_X1   g13023(.A1(new_n13316_), .A2(new_n827_), .B(new_n970_), .ZN(new_n13317_));
  XOR2_X1    g13024(.A1(new_n8568_), .A2(new_n13317_), .Z(new_n13318_));
  NOR2_X1    g13025(.A1(new_n13314_), .A2(new_n13318_), .ZN(new_n13319_));
  NAND2_X1   g13026(.A1(new_n13036_), .A2(new_n13319_), .ZN(new_n13320_));
  NOR2_X1    g13027(.A1(new_n13036_), .A2(new_n13319_), .ZN(new_n13321_));
  INV_X1     g13028(.I(new_n13321_), .ZN(new_n13322_));
  AOI21_X1   g13029(.A1(new_n13322_), .A2(new_n13320_), .B(new_n13033_), .ZN(new_n13323_));
  INV_X1     g13030(.I(new_n13320_), .ZN(new_n13324_));
  NOR3_X1    g13031(.A1(new_n13324_), .A2(new_n13032_), .A3(new_n13321_), .ZN(new_n13325_));
  OAI22_X1   g13032(.A1(new_n607_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n610_), .ZN(new_n13326_));
  OAI21_X1   g13033(.A1(new_n8948_), .A2(new_n684_), .B(new_n13326_), .ZN(new_n13327_));
  AOI21_X1   g13034(.A1(new_n13327_), .A2(new_n612_), .B(new_n607_), .ZN(new_n13328_));
  XNOR2_X1   g13035(.A1(new_n9642_), .A2(new_n13328_), .ZN(new_n13329_));
  INV_X1     g13036(.I(new_n13329_), .ZN(new_n13330_));
  OAI21_X1   g13037(.A1(new_n13323_), .A2(new_n13325_), .B(new_n13330_), .ZN(new_n13331_));
  OAI21_X1   g13038(.A1(new_n13324_), .A2(new_n13321_), .B(new_n13032_), .ZN(new_n13332_));
  NAND3_X1   g13039(.A1(new_n13322_), .A2(new_n13033_), .A3(new_n13320_), .ZN(new_n13333_));
  NAND3_X1   g13040(.A1(new_n13332_), .A2(new_n13333_), .A3(new_n13329_), .ZN(new_n13334_));
  AOI21_X1   g13041(.A1(new_n13331_), .A2(new_n13334_), .B(new_n13029_), .ZN(new_n13335_));
  NAND3_X1   g13042(.A1(new_n13332_), .A2(new_n13333_), .A3(new_n13330_), .ZN(new_n13336_));
  INV_X1     g13043(.I(new_n13336_), .ZN(new_n13337_));
  AOI21_X1   g13044(.A1(new_n13332_), .A2(new_n13333_), .B(new_n13330_), .ZN(new_n13338_));
  OAI21_X1   g13045(.A1(new_n13337_), .A2(new_n13338_), .B(new_n13029_), .ZN(new_n13339_));
  INV_X1     g13046(.I(new_n13339_), .ZN(new_n13340_));
  OAI22_X1   g13047(.A1(new_n448_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n450_), .ZN(new_n13341_));
  OAI21_X1   g13048(.A1(new_n10031_), .A2(new_n496_), .B(new_n13341_), .ZN(new_n13342_));
  AOI21_X1   g13049(.A1(new_n13342_), .A2(new_n452_), .B(new_n448_), .ZN(new_n13343_));
  XNOR2_X1   g13050(.A1(new_n10866_), .A2(new_n13343_), .ZN(new_n13344_));
  INV_X1     g13051(.I(new_n13344_), .ZN(new_n13345_));
  OAI21_X1   g13052(.A1(new_n13340_), .A2(new_n13335_), .B(new_n13345_), .ZN(new_n13346_));
  AOI21_X1   g13053(.A1(new_n13028_), .A2(new_n13026_), .B(new_n13346_), .ZN(new_n13347_));
  AOI21_X1   g13054(.A1(new_n12959_), .A2(new_n13024_), .B(new_n12484_), .ZN(new_n13348_));
  NAND3_X1   g13055(.A1(new_n12958_), .A2(new_n12957_), .A3(new_n12582_), .ZN(new_n13349_));
  NAND2_X1   g13056(.A1(new_n13349_), .A2(new_n12513_), .ZN(new_n13350_));
  INV_X1     g13057(.I(new_n13335_), .ZN(new_n13351_));
  AOI21_X1   g13058(.A1(new_n13351_), .A2(new_n13339_), .B(new_n13344_), .ZN(new_n13352_));
  NOR3_X1    g13059(.A1(new_n13348_), .A2(new_n13350_), .A3(new_n13352_), .ZN(new_n13353_));
  OAI21_X1   g13060(.A1(new_n13347_), .A2(new_n13353_), .B(new_n12958_), .ZN(new_n13354_));
  OAI21_X1   g13061(.A1(new_n13348_), .A2(new_n13350_), .B(new_n13352_), .ZN(new_n13355_));
  NAND3_X1   g13062(.A1(new_n13028_), .A2(new_n13026_), .A3(new_n13346_), .ZN(new_n13356_));
  NAND3_X1   g13063(.A1(new_n13355_), .A2(new_n13356_), .A3(new_n12949_), .ZN(new_n13357_));
  NAND2_X1   g13064(.A1(new_n13354_), .A2(new_n13357_), .ZN(new_n13358_));
  OAI21_X1   g13065(.A1(new_n12987_), .A2(new_n12986_), .B(new_n12984_), .ZN(new_n13359_));
  NOR2_X1    g13066(.A1(\b[58] ), .A2(\b[59] ), .ZN(new_n13360_));
  AOI21_X1   g13067(.A1(new_n12540_), .A2(new_n13360_), .B(new_n12536_), .ZN(new_n13361_));
  NOR2_X1    g13068(.A1(new_n12542_), .A2(new_n12970_), .ZN(new_n13362_));
  INV_X1     g13069(.I(new_n13362_), .ZN(new_n13363_));
  NOR2_X1    g13070(.A1(new_n12540_), .A2(new_n13363_), .ZN(new_n13364_));
  NOR2_X1    g13071(.A1(new_n13361_), .A2(new_n13364_), .ZN(new_n13365_));
  XNOR2_X1   g13072(.A1(\b[59] ), .A2(\b[60] ), .ZN(new_n13366_));
  INV_X1     g13073(.I(\b[60] ), .ZN(new_n13367_));
  NOR2_X1    g13074(.A1(new_n12970_), .A2(new_n13367_), .ZN(new_n13368_));
  NOR2_X1    g13075(.A1(\b[59] ), .A2(\b[60] ), .ZN(new_n13369_));
  OAI21_X1   g13076(.A1(new_n13368_), .A2(new_n13369_), .B(new_n13365_), .ZN(new_n13370_));
  OAI21_X1   g13077(.A1(new_n13365_), .A2(new_n13366_), .B(new_n13370_), .ZN(new_n13371_));
  OAI22_X1   g13078(.A1(new_n330_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n263_), .ZN(new_n13372_));
  OAI21_X1   g13079(.A1(new_n12542_), .A2(new_n289_), .B(new_n13372_), .ZN(new_n13373_));
  AOI21_X1   g13080(.A1(new_n13373_), .A2(new_n260_), .B(new_n426_), .ZN(new_n13374_));
  XNOR2_X1   g13081(.A1(new_n13371_), .A2(new_n13374_), .ZN(new_n13375_));
  INV_X1     g13082(.I(new_n13375_), .ZN(new_n13376_));
  NAND3_X1   g13083(.A1(new_n13359_), .A2(new_n12980_), .A3(new_n13376_), .ZN(new_n13377_));
  AOI21_X1   g13084(.A1(new_n12962_), .A2(new_n12966_), .B(new_n12983_), .ZN(new_n13378_));
  OAI21_X1   g13085(.A1(new_n13378_), .A2(new_n12979_), .B(new_n13375_), .ZN(new_n13379_));
  AOI21_X1   g13086(.A1(new_n13377_), .A2(new_n13379_), .B(new_n13358_), .ZN(new_n13380_));
  AOI21_X1   g13087(.A1(new_n13355_), .A2(new_n13356_), .B(new_n12949_), .ZN(new_n13381_));
  NOR3_X1    g13088(.A1(new_n13347_), .A2(new_n13353_), .A3(new_n12958_), .ZN(new_n13382_));
  NOR2_X1    g13089(.A1(new_n13382_), .A2(new_n13381_), .ZN(new_n13383_));
  NOR3_X1    g13090(.A1(new_n13378_), .A2(new_n12979_), .A3(new_n13375_), .ZN(new_n13384_));
  AOI21_X1   g13091(.A1(new_n13359_), .A2(new_n12980_), .B(new_n13376_), .ZN(new_n13385_));
  NOR3_X1    g13092(.A1(new_n13383_), .A2(new_n13385_), .A3(new_n13384_), .ZN(new_n13386_));
  OAI21_X1   g13093(.A1(new_n13380_), .A2(new_n13386_), .B(new_n13023_), .ZN(new_n13387_));
  INV_X1     g13094(.I(new_n13023_), .ZN(new_n13388_));
  OAI21_X1   g13095(.A1(new_n13384_), .A2(new_n13385_), .B(new_n13383_), .ZN(new_n13389_));
  NAND3_X1   g13096(.A1(new_n13358_), .A2(new_n13379_), .A3(new_n13377_), .ZN(new_n13390_));
  NAND3_X1   g13097(.A1(new_n13389_), .A2(new_n13390_), .A3(new_n13388_), .ZN(new_n13391_));
  NAND3_X1   g13098(.A1(new_n13387_), .A2(new_n13391_), .A3(new_n13019_), .ZN(new_n13392_));
  NAND2_X1   g13099(.A1(new_n13392_), .A2(new_n13008_), .ZN(new_n13393_));
  XOR2_X1    g13100(.A1(new_n13393_), .A2(new_n13015_), .Z(\f[60] ));
  NAND2_X1   g13101(.A1(new_n13359_), .A2(new_n12980_), .ZN(new_n13395_));
  NAND2_X1   g13102(.A1(new_n13383_), .A2(new_n13376_), .ZN(new_n13396_));
  NAND2_X1   g13103(.A1(new_n13358_), .A2(new_n13375_), .ZN(new_n13397_));
  AOI21_X1   g13104(.A1(new_n13396_), .A2(new_n13397_), .B(new_n13388_), .ZN(new_n13398_));
  NOR2_X1    g13105(.A1(new_n13358_), .A2(new_n13375_), .ZN(new_n13399_));
  NOR2_X1    g13106(.A1(new_n13383_), .A2(new_n13376_), .ZN(new_n13400_));
  NOR3_X1    g13107(.A1(new_n13400_), .A2(new_n13399_), .A3(new_n13023_), .ZN(new_n13401_));
  OAI21_X1   g13108(.A1(new_n13398_), .A2(new_n13401_), .B(new_n13395_), .ZN(new_n13402_));
  AOI21_X1   g13109(.A1(new_n13387_), .A2(new_n13391_), .B(new_n13019_), .ZN(new_n13403_));
  OAI21_X1   g13110(.A1(new_n13403_), .A2(new_n13008_), .B(new_n12576_), .ZN(new_n13404_));
  OAI21_X1   g13111(.A1(new_n13029_), .A2(new_n13338_), .B(new_n13336_), .ZN(new_n13405_));
  INV_X1     g13112(.I(new_n13405_), .ZN(new_n13406_));
  NAND2_X1   g13113(.A1(new_n13304_), .A2(new_n13307_), .ZN(new_n13407_));
  NAND2_X1   g13114(.A1(new_n13407_), .A2(new_n13309_), .ZN(new_n13408_));
  OAI21_X1   g13115(.A1(new_n13309_), .A2(new_n13312_), .B(new_n13408_), .ZN(new_n13409_));
  NAND3_X1   g13116(.A1(new_n13409_), .A2(new_n13035_), .A3(new_n13034_), .ZN(new_n13410_));
  AOI21_X1   g13117(.A1(new_n13034_), .A2(new_n13035_), .B(new_n13409_), .ZN(new_n13411_));
  INV_X1     g13118(.I(new_n13318_), .ZN(new_n13412_));
  NAND3_X1   g13119(.A1(new_n13031_), .A2(new_n12898_), .A3(new_n13412_), .ZN(new_n13413_));
  OAI21_X1   g13120(.A1(new_n13411_), .A2(new_n13413_), .B(new_n13410_), .ZN(new_n13414_));
  AOI21_X1   g13121(.A1(new_n12587_), .A2(new_n12894_), .B(new_n12905_), .ZN(new_n13415_));
  INV_X1     g13122(.I(new_n13310_), .ZN(new_n13416_));
  OAI21_X1   g13123(.A1(new_n13415_), .A2(new_n13311_), .B(new_n13416_), .ZN(new_n13417_));
  AOI21_X1   g13124(.A1(new_n13280_), .A2(new_n13283_), .B(new_n12889_), .ZN(new_n13418_));
  INV_X1     g13125(.I(new_n13418_), .ZN(new_n13419_));
  NAND3_X1   g13126(.A1(new_n13280_), .A2(new_n13283_), .A3(new_n12889_), .ZN(new_n13420_));
  NAND2_X1   g13127(.A1(new_n13420_), .A2(new_n13292_), .ZN(new_n13421_));
  OAI21_X1   g13128(.A1(new_n13421_), .A2(new_n12893_), .B(new_n13419_), .ZN(new_n13422_));
  AOI21_X1   g13129(.A1(new_n13276_), .A2(new_n13277_), .B(new_n12862_), .ZN(new_n13423_));
  INV_X1     g13130(.I(new_n13423_), .ZN(new_n13424_));
  NAND3_X1   g13131(.A1(new_n13276_), .A2(new_n13277_), .A3(new_n12862_), .ZN(new_n13425_));
  NAND3_X1   g13132(.A1(new_n13039_), .A2(new_n13425_), .A3(new_n13271_), .ZN(new_n13426_));
  NAND2_X1   g13133(.A1(new_n13426_), .A2(new_n13424_), .ZN(new_n13427_));
  NOR2_X1    g13134(.A1(new_n13234_), .A2(new_n13227_), .ZN(new_n13428_));
  OR3_X2     g13135(.A1(new_n13242_), .A2(new_n13243_), .A3(new_n13428_), .Z(new_n13429_));
  NAND2_X1   g13136(.A1(new_n13049_), .A2(new_n12825_), .ZN(new_n13430_));
  AND2_X2    g13137(.A1(new_n13430_), .A2(new_n13428_), .Z(new_n13431_));
  NAND2_X1   g13138(.A1(new_n13047_), .A2(new_n13239_), .ZN(new_n13432_));
  OAI21_X1   g13139(.A1(new_n13431_), .A2(new_n13432_), .B(new_n13429_), .ZN(new_n13433_));
  OAI22_X1   g13140(.A1(new_n3260_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n3709_), .ZN(new_n13434_));
  OAI21_X1   g13141(.A1(new_n3018_), .A2(new_n3569_), .B(new_n13434_), .ZN(new_n13435_));
  AOI21_X1   g13142(.A1(new_n13435_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n13436_));
  XNOR2_X1   g13143(.A1(new_n3514_), .A2(new_n13436_), .ZN(new_n13437_));
  NAND2_X1   g13144(.A1(new_n13209_), .A2(new_n13057_), .ZN(new_n13438_));
  NOR2_X1    g13145(.A1(new_n13209_), .A2(new_n13057_), .ZN(new_n13439_));
  NAND2_X1   g13146(.A1(new_n13059_), .A2(new_n13199_), .ZN(new_n13440_));
  OAI21_X1   g13147(.A1(new_n13440_), .A2(new_n13439_), .B(new_n13438_), .ZN(new_n13441_));
  NAND2_X1   g13148(.A1(new_n13053_), .A2(new_n13215_), .ZN(new_n13442_));
  NOR2_X1    g13149(.A1(new_n13054_), .A2(new_n13219_), .ZN(new_n13443_));
  OAI21_X1   g13150(.A1(new_n13053_), .A2(new_n13215_), .B(new_n13443_), .ZN(new_n13444_));
  NOR2_X1    g13151(.A1(new_n13066_), .A2(new_n13164_), .ZN(new_n13445_));
  OAI21_X1   g13152(.A1(new_n13135_), .A2(new_n13139_), .B(new_n12705_), .ZN(new_n13446_));
  NAND3_X1   g13153(.A1(new_n13147_), .A2(new_n13148_), .A3(new_n12710_), .ZN(new_n13447_));
  NAND3_X1   g13154(.A1(new_n13067_), .A2(new_n13144_), .A3(new_n13447_), .ZN(new_n13448_));
  NAND2_X1   g13155(.A1(new_n13118_), .A2(new_n13121_), .ZN(new_n13449_));
  NAND2_X1   g13156(.A1(new_n13449_), .A2(new_n13068_), .ZN(new_n13450_));
  INV_X1     g13157(.I(new_n13450_), .ZN(new_n13451_));
  NOR2_X1    g13158(.A1(new_n13449_), .A2(new_n13068_), .ZN(new_n13452_));
  NOR4_X1    g13159(.A1(new_n13452_), .A2(new_n13069_), .A3(new_n13070_), .A4(new_n13125_), .ZN(new_n13453_));
  AOI21_X1   g13160(.A1(new_n13113_), .A2(new_n13115_), .B(new_n13072_), .ZN(new_n13454_));
  NOR3_X1    g13161(.A1(new_n13105_), .A2(new_n13071_), .A3(new_n13101_), .ZN(new_n13455_));
  NOR3_X1    g13162(.A1(new_n13112_), .A2(new_n13455_), .A3(new_n13108_), .ZN(new_n13456_));
  NOR2_X1    g13163(.A1(new_n13456_), .A2(new_n13454_), .ZN(new_n13457_));
  NAND2_X1   g13164(.A1(new_n13102_), .A2(new_n13100_), .ZN(new_n13458_));
  NOR2_X1    g13165(.A1(new_n13084_), .A2(new_n258_), .ZN(new_n13459_));
  INV_X1     g13166(.I(new_n13459_), .ZN(new_n13460_));
  AOI21_X1   g13167(.A1(new_n13085_), .A2(new_n13086_), .B(new_n13460_), .ZN(new_n13461_));
  AOI22_X1   g13168(.A1(new_n13078_), .A2(\b[2] ), .B1(new_n10957_), .B2(new_n12218_), .ZN(new_n13462_));
  OAI21_X1   g13169(.A1(new_n13462_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n13463_));
  XOR2_X1    g13170(.A1(new_n13463_), .A2(new_n329_), .Z(new_n13464_));
  XNOR2_X1   g13171(.A1(\a[61] ), .A2(\a[62] ), .ZN(new_n13465_));
  NOR2_X1    g13172(.A1(new_n13077_), .A2(new_n13465_), .ZN(new_n13466_));
  INV_X1     g13173(.I(\a[61] ), .ZN(new_n13467_));
  NAND3_X1   g13174(.A1(new_n13467_), .A2(\a[59] ), .A3(\a[60] ), .ZN(new_n13468_));
  OAI21_X1   g13175(.A1(new_n13467_), .A2(new_n13076_), .B(new_n13468_), .ZN(new_n13469_));
  XOR2_X1    g13176(.A1(\a[61] ), .A2(\a[62] ), .Z(new_n13470_));
  NOR2_X1    g13177(.A1(new_n13077_), .A2(new_n13470_), .ZN(new_n13471_));
  NAND2_X1   g13178(.A1(new_n13471_), .A2(new_n13469_), .ZN(new_n13472_));
  NOR2_X1    g13179(.A1(new_n319_), .A2(\a[62] ), .ZN(new_n13473_));
  NAND2_X1   g13180(.A1(new_n13472_), .A2(new_n13473_), .ZN(new_n13474_));
  AOI21_X1   g13181(.A1(new_n13474_), .A2(new_n13466_), .B(new_n444_), .ZN(new_n13475_));
  INV_X1     g13182(.I(\a[62] ), .ZN(new_n13476_));
  NAND3_X1   g13183(.A1(new_n13474_), .A2(new_n444_), .A3(new_n13466_), .ZN(new_n13477_));
  NAND2_X1   g13184(.A1(new_n13477_), .A2(new_n13476_), .ZN(new_n13478_));
  NOR2_X1    g13185(.A1(new_n13478_), .A2(new_n13475_), .ZN(new_n13479_));
  NOR2_X1    g13186(.A1(new_n13479_), .A2(new_n258_), .ZN(new_n13480_));
  XOR2_X1    g13187(.A1(new_n13480_), .A2(new_n13077_), .Z(new_n13481_));
  XOR2_X1    g13188(.A1(new_n13481_), .A2(new_n13464_), .Z(new_n13482_));
  OAI21_X1   g13189(.A1(new_n13087_), .A2(new_n13461_), .B(new_n13482_), .ZN(new_n13483_));
  NOR2_X1    g13190(.A1(new_n13461_), .A2(new_n13087_), .ZN(new_n13484_));
  INV_X1     g13191(.I(new_n13464_), .ZN(new_n13485_));
  XOR2_X1    g13192(.A1(new_n13480_), .A2(new_n13084_), .Z(new_n13486_));
  NOR2_X1    g13193(.A1(new_n13486_), .A2(new_n13485_), .ZN(new_n13487_));
  NOR2_X1    g13194(.A1(new_n13481_), .A2(new_n13464_), .ZN(new_n13488_));
  OAI21_X1   g13195(.A1(new_n13487_), .A2(new_n13488_), .B(new_n13484_), .ZN(new_n13489_));
  NAND2_X1   g13196(.A1(new_n13483_), .A2(new_n13489_), .ZN(new_n13490_));
  OAI22_X1   g13197(.A1(new_n10979_), .A2(new_n509_), .B1(new_n419_), .B2(new_n11401_), .ZN(new_n13491_));
  AOI21_X1   g13198(.A1(new_n13491_), .A2(new_n10973_), .B(new_n10964_), .ZN(new_n13492_));
  XOR2_X1    g13199(.A1(new_n471_), .A2(new_n13492_), .Z(new_n13493_));
  INV_X1     g13200(.I(new_n13493_), .ZN(new_n13494_));
  NAND2_X1   g13201(.A1(new_n13490_), .A2(new_n13494_), .ZN(new_n13495_));
  NAND3_X1   g13202(.A1(new_n13483_), .A2(new_n13489_), .A3(new_n13493_), .ZN(new_n13496_));
  AOI22_X1   g13203(.A1(new_n13495_), .A2(new_n13496_), .B1(new_n13097_), .B2(new_n13458_), .ZN(new_n13497_));
  NAND2_X1   g13204(.A1(new_n13458_), .A2(new_n13097_), .ZN(new_n13498_));
  NAND3_X1   g13205(.A1(new_n13483_), .A2(new_n13489_), .A3(new_n13494_), .ZN(new_n13499_));
  NAND2_X1   g13206(.A1(new_n13490_), .A2(new_n13493_), .ZN(new_n13500_));
  AOI21_X1   g13207(.A1(new_n13499_), .A2(new_n13500_), .B(new_n13498_), .ZN(new_n13501_));
  NOR2_X1    g13208(.A1(new_n13501_), .A2(new_n13497_), .ZN(new_n13502_));
  INV_X1     g13209(.I(new_n657_), .ZN(new_n13503_));
  AOI22_X1   g13210(.A1(new_n11415_), .A2(new_n13503_), .B1(\b[8] ), .B2(new_n10145_), .ZN(new_n13504_));
  OAI21_X1   g13211(.A1(new_n13504_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n13505_));
  XOR2_X1    g13212(.A1(new_n660_), .A2(new_n13505_), .Z(new_n13506_));
  NOR2_X1    g13213(.A1(new_n13502_), .A2(new_n13506_), .ZN(new_n13507_));
  INV_X1     g13214(.I(new_n13506_), .ZN(new_n13508_));
  NOR3_X1    g13215(.A1(new_n13501_), .A2(new_n13497_), .A3(new_n13508_), .ZN(new_n13509_));
  NOR2_X1    g13216(.A1(new_n13507_), .A2(new_n13509_), .ZN(new_n13510_));
  NOR2_X1    g13217(.A1(new_n13510_), .A2(new_n13457_), .ZN(new_n13511_));
  NOR3_X1    g13218(.A1(new_n13501_), .A2(new_n13497_), .A3(new_n13506_), .ZN(new_n13512_));
  OAI21_X1   g13219(.A1(new_n13501_), .A2(new_n13497_), .B(new_n13506_), .ZN(new_n13513_));
  INV_X1     g13220(.I(new_n13513_), .ZN(new_n13514_));
  OAI21_X1   g13221(.A1(new_n13514_), .A2(new_n13512_), .B(new_n13457_), .ZN(new_n13515_));
  INV_X1     g13222(.I(new_n13515_), .ZN(new_n13516_));
  AOI22_X1   g13223(.A1(new_n8631_), .A2(\b[12] ), .B1(\b[13] ), .B2(new_n9382_), .ZN(new_n13517_));
  AOI21_X1   g13224(.A1(\b[11] ), .A2(new_n9731_), .B(new_n13517_), .ZN(new_n13518_));
  OAI21_X1   g13225(.A1(new_n13518_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n13519_));
  XOR2_X1    g13226(.A1(new_n860_), .A2(new_n13519_), .Z(new_n13520_));
  NOR3_X1    g13227(.A1(new_n13516_), .A2(new_n13511_), .A3(new_n13520_), .ZN(new_n13521_));
  INV_X1     g13228(.I(new_n13457_), .ZN(new_n13522_));
  OAI21_X1   g13229(.A1(new_n13507_), .A2(new_n13509_), .B(new_n13522_), .ZN(new_n13523_));
  INV_X1     g13230(.I(new_n13520_), .ZN(new_n13524_));
  AOI21_X1   g13231(.A1(new_n13523_), .A2(new_n13515_), .B(new_n13524_), .ZN(new_n13525_));
  OAI22_X1   g13232(.A1(new_n13453_), .A2(new_n13451_), .B1(new_n13521_), .B2(new_n13525_), .ZN(new_n13526_));
  NOR2_X1    g13233(.A1(new_n13453_), .A2(new_n13451_), .ZN(new_n13527_));
  OAI21_X1   g13234(.A1(new_n13516_), .A2(new_n13511_), .B(new_n13524_), .ZN(new_n13528_));
  NAND3_X1   g13235(.A1(new_n13523_), .A2(new_n13515_), .A3(new_n13520_), .ZN(new_n13529_));
  NAND2_X1   g13236(.A1(new_n13528_), .A2(new_n13529_), .ZN(new_n13530_));
  NAND2_X1   g13237(.A1(new_n13527_), .A2(new_n13530_), .ZN(new_n13531_));
  OAI22_X1   g13238(.A1(new_n7619_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n8309_), .ZN(new_n13532_));
  OAI21_X1   g13239(.A1(new_n930_), .A2(new_n7947_), .B(new_n13532_), .ZN(new_n13533_));
  AOI21_X1   g13240(.A1(new_n13533_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n13534_));
  XOR2_X1    g13241(.A1(new_n1114_), .A2(new_n13534_), .Z(new_n13535_));
  INV_X1     g13242(.I(new_n13535_), .ZN(new_n13536_));
  NAND3_X1   g13243(.A1(new_n13531_), .A2(new_n13526_), .A3(new_n13536_), .ZN(new_n13537_));
  NAND2_X1   g13244(.A1(new_n13531_), .A2(new_n13526_), .ZN(new_n13538_));
  NAND2_X1   g13245(.A1(new_n13538_), .A2(new_n13535_), .ZN(new_n13539_));
  AOI22_X1   g13246(.A1(new_n13539_), .A2(new_n13537_), .B1(new_n13448_), .B2(new_n13446_), .ZN(new_n13540_));
  NAND2_X1   g13247(.A1(new_n13448_), .A2(new_n13446_), .ZN(new_n13541_));
  AOI21_X1   g13248(.A1(new_n13531_), .A2(new_n13526_), .B(new_n13535_), .ZN(new_n13542_));
  NOR2_X1    g13249(.A1(new_n13521_), .A2(new_n13525_), .ZN(new_n13543_));
  NOR2_X1    g13250(.A1(new_n13527_), .A2(new_n13543_), .ZN(new_n13544_));
  AOI21_X1   g13251(.A1(new_n13523_), .A2(new_n13515_), .B(new_n13520_), .ZN(new_n13545_));
  NOR3_X1    g13252(.A1(new_n13516_), .A2(new_n13511_), .A3(new_n13524_), .ZN(new_n13546_));
  NOR2_X1    g13253(.A1(new_n13546_), .A2(new_n13545_), .ZN(new_n13547_));
  NOR3_X1    g13254(.A1(new_n13547_), .A2(new_n13451_), .A3(new_n13453_), .ZN(new_n13548_));
  NOR3_X1    g13255(.A1(new_n13548_), .A2(new_n13544_), .A3(new_n13536_), .ZN(new_n13549_));
  NOR2_X1    g13256(.A1(new_n13549_), .A2(new_n13542_), .ZN(new_n13550_));
  NOR2_X1    g13257(.A1(new_n13541_), .A2(new_n13550_), .ZN(new_n13551_));
  OAI22_X1   g13258(.A1(new_n6644_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n6647_), .ZN(new_n13552_));
  OAI21_X1   g13259(.A1(new_n1189_), .A2(new_n7284_), .B(new_n13552_), .ZN(new_n13553_));
  AOI21_X1   g13260(.A1(new_n13553_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n13554_));
  XNOR2_X1   g13261(.A1(new_n1421_), .A2(new_n13554_), .ZN(new_n13555_));
  INV_X1     g13262(.I(new_n13555_), .ZN(new_n13556_));
  OAI21_X1   g13263(.A1(new_n13551_), .A2(new_n13540_), .B(new_n13556_), .ZN(new_n13557_));
  NOR2_X1    g13264(.A1(new_n13445_), .A2(new_n13557_), .ZN(new_n13558_));
  INV_X1     g13265(.I(new_n13557_), .ZN(new_n13559_));
  NOR3_X1    g13266(.A1(new_n13559_), .A2(new_n13066_), .A3(new_n13164_), .ZN(new_n13560_));
  OAI21_X1   g13267(.A1(new_n13558_), .A2(new_n13560_), .B(new_n13163_), .ZN(new_n13561_));
  AOI21_X1   g13268(.A1(new_n13151_), .A2(new_n13154_), .B(new_n13159_), .ZN(new_n13562_));
  OAI21_X1   g13269(.A1(new_n13066_), .A2(new_n13164_), .B(new_n13559_), .ZN(new_n13563_));
  INV_X1     g13270(.I(new_n13160_), .ZN(new_n13564_));
  NOR2_X1    g13271(.A1(new_n13564_), .A2(new_n13562_), .ZN(new_n13565_));
  NAND4_X1   g13272(.A1(new_n13565_), .A2(new_n13557_), .A3(new_n13063_), .A4(new_n13065_), .ZN(new_n13566_));
  NAND3_X1   g13273(.A1(new_n13563_), .A2(new_n13566_), .A3(new_n13562_), .ZN(new_n13567_));
  OAI22_X1   g13274(.A1(new_n5993_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n5991_), .ZN(new_n13568_));
  OAI21_X1   g13275(.A1(new_n1525_), .A2(new_n5997_), .B(new_n13568_), .ZN(new_n13569_));
  AOI21_X1   g13276(.A1(new_n13569_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n13570_));
  XOR2_X1    g13277(.A1(new_n1808_), .A2(new_n13570_), .Z(new_n13571_));
  AOI21_X1   g13278(.A1(new_n13561_), .A2(new_n13567_), .B(new_n13571_), .ZN(new_n13572_));
  AOI21_X1   g13279(.A1(new_n13563_), .A2(new_n13566_), .B(new_n13562_), .ZN(new_n13573_));
  NOR3_X1    g13280(.A1(new_n13558_), .A2(new_n13163_), .A3(new_n13560_), .ZN(new_n13574_));
  INV_X1     g13281(.I(new_n13571_), .ZN(new_n13575_));
  NOR3_X1    g13282(.A1(new_n13574_), .A2(new_n13573_), .A3(new_n13575_), .ZN(new_n13576_));
  NOR2_X1    g13283(.A1(new_n13576_), .A2(new_n13572_), .ZN(new_n13577_));
  NAND2_X1   g13284(.A1(new_n13173_), .A2(new_n13170_), .ZN(new_n13578_));
  OAI22_X1   g13285(.A1(new_n13060_), .A2(new_n12740_), .B1(new_n13173_), .B2(new_n13170_), .ZN(new_n13579_));
  NAND2_X1   g13286(.A1(new_n13579_), .A2(new_n13578_), .ZN(new_n13580_));
  OAI22_X1   g13287(.A1(new_n5420_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n5107_), .ZN(new_n13581_));
  OAI21_X1   g13288(.A1(new_n1936_), .A2(new_n5112_), .B(new_n13581_), .ZN(new_n13582_));
  AOI21_X1   g13289(.A1(new_n13582_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n13583_));
  XNOR2_X1   g13290(.A1(new_n2280_), .A2(new_n13583_), .ZN(new_n13584_));
  INV_X1     g13291(.I(new_n13584_), .ZN(new_n13585_));
  NAND2_X1   g13292(.A1(new_n13580_), .A2(new_n13585_), .ZN(new_n13586_));
  NAND2_X1   g13293(.A1(new_n12729_), .A2(new_n12731_), .ZN(new_n13587_));
  AOI22_X1   g13294(.A1(new_n13587_), .A2(new_n12726_), .B1(new_n13165_), .B2(new_n13169_), .ZN(new_n13588_));
  NOR2_X1    g13295(.A1(new_n13588_), .A2(new_n13172_), .ZN(new_n13589_));
  NAND2_X1   g13296(.A1(new_n13589_), .A2(new_n13584_), .ZN(new_n13590_));
  AND2_X2    g13297(.A1(new_n13586_), .A2(new_n13590_), .Z(new_n13591_));
  NOR2_X1    g13298(.A1(new_n13580_), .A2(new_n13584_), .ZN(new_n13592_));
  NOR2_X1    g13299(.A1(new_n13589_), .A2(new_n13585_), .ZN(new_n13593_));
  OAI21_X1   g13300(.A1(new_n13592_), .A2(new_n13593_), .B(new_n13577_), .ZN(new_n13594_));
  OAI21_X1   g13301(.A1(new_n13591_), .A2(new_n13577_), .B(new_n13594_), .ZN(new_n13595_));
  AOI21_X1   g13302(.A1(new_n13176_), .A2(new_n13189_), .B(new_n13203_), .ZN(new_n13596_));
  OAI22_X1   g13303(.A1(new_n4072_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n4067_), .ZN(new_n13597_));
  OAI21_X1   g13304(.A1(new_n2439_), .A2(new_n4318_), .B(new_n13597_), .ZN(new_n13598_));
  AOI21_X1   g13305(.A1(new_n13598_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n13599_));
  XNOR2_X1   g13306(.A1(new_n2846_), .A2(new_n13599_), .ZN(new_n13600_));
  NOR2_X1    g13307(.A1(new_n13596_), .A2(new_n13600_), .ZN(new_n13601_));
  OAI21_X1   g13308(.A1(new_n13192_), .A2(new_n13204_), .B(new_n13187_), .ZN(new_n13602_));
  INV_X1     g13309(.I(new_n13600_), .ZN(new_n13603_));
  NOR2_X1    g13310(.A1(new_n13602_), .A2(new_n13603_), .ZN(new_n13604_));
  OAI21_X1   g13311(.A1(new_n13604_), .A2(new_n13601_), .B(new_n13595_), .ZN(new_n13605_));
  NAND2_X1   g13312(.A1(new_n13596_), .A2(new_n13603_), .ZN(new_n13606_));
  NAND2_X1   g13313(.A1(new_n13602_), .A2(new_n13600_), .ZN(new_n13607_));
  AOI21_X1   g13314(.A1(new_n13607_), .A2(new_n13606_), .B(new_n13595_), .ZN(new_n13608_));
  INV_X1     g13315(.I(new_n13608_), .ZN(new_n13609_));
  NAND2_X1   g13316(.A1(new_n13609_), .A2(new_n13605_), .ZN(new_n13610_));
  NAND3_X1   g13317(.A1(new_n13444_), .A2(new_n13442_), .A3(new_n13610_), .ZN(new_n13611_));
  NOR2_X1    g13318(.A1(new_n13231_), .A2(new_n13225_), .ZN(new_n13612_));
  NAND2_X1   g13319(.A1(new_n13222_), .A2(new_n13220_), .ZN(new_n13613_));
  AOI21_X1   g13320(.A1(new_n13231_), .A2(new_n13225_), .B(new_n13613_), .ZN(new_n13614_));
  OR2_X2     g13321(.A1(new_n13604_), .A2(new_n13601_), .Z(new_n13615_));
  AOI21_X1   g13322(.A1(new_n13615_), .A2(new_n13595_), .B(new_n13608_), .ZN(new_n13616_));
  OAI21_X1   g13323(.A1(new_n13614_), .A2(new_n13612_), .B(new_n13616_), .ZN(new_n13617_));
  AOI21_X1   g13324(.A1(new_n13617_), .A2(new_n13611_), .B(new_n13441_), .ZN(new_n13618_));
  INV_X1     g13325(.I(new_n13441_), .ZN(new_n13619_));
  NOR3_X1    g13326(.A1(new_n13614_), .A2(new_n13612_), .A3(new_n13616_), .ZN(new_n13620_));
  AOI21_X1   g13327(.A1(new_n13444_), .A2(new_n13442_), .B(new_n13610_), .ZN(new_n13621_));
  NOR3_X1    g13328(.A1(new_n13620_), .A2(new_n13621_), .A3(new_n13619_), .ZN(new_n13622_));
  OAI21_X1   g13329(.A1(new_n13622_), .A2(new_n13618_), .B(new_n13437_), .ZN(new_n13623_));
  INV_X1     g13330(.I(new_n13437_), .ZN(new_n13624_));
  OAI21_X1   g13331(.A1(new_n13620_), .A2(new_n13621_), .B(new_n13619_), .ZN(new_n13625_));
  NAND3_X1   g13332(.A1(new_n13617_), .A2(new_n13611_), .A3(new_n13441_), .ZN(new_n13626_));
  NAND3_X1   g13333(.A1(new_n13625_), .A2(new_n13626_), .A3(new_n13624_), .ZN(new_n13627_));
  OAI22_X1   g13334(.A1(new_n3989_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n4253_), .ZN(new_n13628_));
  OAI21_X1   g13335(.A1(new_n3717_), .A2(new_n2884_), .B(new_n13628_), .ZN(new_n13629_));
  AOI21_X1   g13336(.A1(new_n13629_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n13630_));
  XNOR2_X1   g13337(.A1(new_n4257_), .A2(new_n13630_), .ZN(new_n13631_));
  INV_X1     g13338(.I(new_n13631_), .ZN(new_n13632_));
  NAND3_X1   g13339(.A1(new_n13623_), .A2(new_n13627_), .A3(new_n13632_), .ZN(new_n13633_));
  AOI21_X1   g13340(.A1(new_n13625_), .A2(new_n13626_), .B(new_n13624_), .ZN(new_n13634_));
  NOR3_X1    g13341(.A1(new_n13622_), .A2(new_n13618_), .A3(new_n13437_), .ZN(new_n13635_));
  OAI21_X1   g13342(.A1(new_n13635_), .A2(new_n13634_), .B(new_n13631_), .ZN(new_n13636_));
  NAND2_X1   g13343(.A1(new_n13636_), .A2(new_n13633_), .ZN(new_n13637_));
  NAND2_X1   g13344(.A1(new_n13433_), .A2(new_n13637_), .ZN(new_n13638_));
  NOR2_X1    g13345(.A1(new_n13430_), .A2(new_n13428_), .ZN(new_n13639_));
  NAND2_X1   g13346(.A1(new_n13430_), .A2(new_n13428_), .ZN(new_n13640_));
  INV_X1     g13347(.I(new_n13432_), .ZN(new_n13641_));
  AOI21_X1   g13348(.A1(new_n13641_), .A2(new_n13640_), .B(new_n13639_), .ZN(new_n13642_));
  NAND2_X1   g13349(.A1(new_n13623_), .A2(new_n13627_), .ZN(new_n13643_));
  NAND2_X1   g13350(.A1(new_n13643_), .A2(new_n13632_), .ZN(new_n13644_));
  NOR2_X1    g13351(.A1(new_n13635_), .A2(new_n13634_), .ZN(new_n13645_));
  NAND2_X1   g13352(.A1(new_n13645_), .A2(new_n13631_), .ZN(new_n13646_));
  NAND2_X1   g13353(.A1(new_n13646_), .A2(new_n13644_), .ZN(new_n13647_));
  NAND2_X1   g13354(.A1(new_n13647_), .A2(new_n13642_), .ZN(new_n13648_));
  OAI22_X1   g13355(.A1(new_n2171_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n2166_), .ZN(new_n13649_));
  OAI21_X1   g13356(.A1(new_n4500_), .A2(new_n2322_), .B(new_n13649_), .ZN(new_n13650_));
  AOI21_X1   g13357(.A1(new_n13650_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n13651_));
  XOR2_X1    g13358(.A1(new_n5067_), .A2(new_n13651_), .Z(new_n13652_));
  INV_X1     g13359(.I(new_n13652_), .ZN(new_n13653_));
  NAND3_X1   g13360(.A1(new_n13648_), .A2(new_n13638_), .A3(new_n13653_), .ZN(new_n13654_));
  INV_X1     g13361(.I(new_n13654_), .ZN(new_n13655_));
  AOI21_X1   g13362(.A1(new_n13648_), .A2(new_n13638_), .B(new_n13653_), .ZN(new_n13656_));
  NOR2_X1    g13363(.A1(new_n13655_), .A2(new_n13656_), .ZN(new_n13657_));
  AOI21_X1   g13364(.A1(new_n13246_), .A2(new_n13249_), .B(new_n12844_), .ZN(new_n13658_));
  INV_X1     g13365(.I(new_n13658_), .ZN(new_n13659_));
  NAND3_X1   g13366(.A1(new_n13246_), .A2(new_n13249_), .A3(new_n12844_), .ZN(new_n13660_));
  NAND3_X1   g13367(.A1(new_n13257_), .A2(new_n13260_), .A3(new_n13660_), .ZN(new_n13661_));
  NAND2_X1   g13368(.A1(new_n13661_), .A2(new_n13659_), .ZN(new_n13662_));
  OAI22_X1   g13369(.A1(new_n1712_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n1707_), .ZN(new_n13663_));
  OAI21_X1   g13370(.A1(new_n5353_), .A2(new_n1850_), .B(new_n13663_), .ZN(new_n13664_));
  AOI21_X1   g13371(.A1(new_n13664_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n13665_));
  XOR2_X1    g13372(.A1(new_n5926_), .A2(new_n13665_), .Z(new_n13666_));
  INV_X1     g13373(.I(new_n13666_), .ZN(new_n13667_));
  NAND2_X1   g13374(.A1(new_n13662_), .A2(new_n13667_), .ZN(new_n13668_));
  NOR2_X1    g13375(.A1(new_n13662_), .A2(new_n13667_), .ZN(new_n13669_));
  INV_X1     g13376(.I(new_n13669_), .ZN(new_n13670_));
  AOI21_X1   g13377(.A1(new_n13670_), .A2(new_n13668_), .B(new_n13657_), .ZN(new_n13671_));
  NOR3_X1    g13378(.A1(new_n13635_), .A2(new_n13634_), .A3(new_n13631_), .ZN(new_n13672_));
  AOI21_X1   g13379(.A1(new_n13623_), .A2(new_n13627_), .B(new_n13632_), .ZN(new_n13673_));
  NOR2_X1    g13380(.A1(new_n13672_), .A2(new_n13673_), .ZN(new_n13674_));
  NOR2_X1    g13381(.A1(new_n13642_), .A2(new_n13674_), .ZN(new_n13675_));
  AOI21_X1   g13382(.A1(new_n13644_), .A2(new_n13646_), .B(new_n13433_), .ZN(new_n13676_));
  OAI21_X1   g13383(.A1(new_n13676_), .A2(new_n13675_), .B(new_n13652_), .ZN(new_n13677_));
  NAND2_X1   g13384(.A1(new_n13677_), .A2(new_n13654_), .ZN(new_n13678_));
  NOR2_X1    g13385(.A1(new_n13662_), .A2(new_n13666_), .ZN(new_n13679_));
  INV_X1     g13386(.I(new_n13679_), .ZN(new_n13680_));
  NAND2_X1   g13387(.A1(new_n13662_), .A2(new_n13666_), .ZN(new_n13681_));
  AOI21_X1   g13388(.A1(new_n13680_), .A2(new_n13681_), .B(new_n13678_), .ZN(new_n13682_));
  NOR2_X1    g13389(.A1(new_n13671_), .A2(new_n13682_), .ZN(new_n13683_));
  NOR2_X1    g13390(.A1(new_n13683_), .A2(new_n13427_), .ZN(new_n13684_));
  NOR3_X1    g13391(.A1(new_n13263_), .A2(new_n13266_), .A3(new_n12855_), .ZN(new_n13685_));
  NOR2_X1    g13392(.A1(new_n13685_), .A2(new_n13270_), .ZN(new_n13686_));
  AOI21_X1   g13393(.A1(new_n13686_), .A2(new_n13039_), .B(new_n13423_), .ZN(new_n13687_));
  INV_X1     g13394(.I(new_n13668_), .ZN(new_n13688_));
  OAI21_X1   g13395(.A1(new_n13688_), .A2(new_n13669_), .B(new_n13678_), .ZN(new_n13689_));
  INV_X1     g13396(.I(new_n13681_), .ZN(new_n13690_));
  OAI21_X1   g13397(.A1(new_n13690_), .A2(new_n13679_), .B(new_n13657_), .ZN(new_n13691_));
  NAND2_X1   g13398(.A1(new_n13689_), .A2(new_n13691_), .ZN(new_n13692_));
  NOR2_X1    g13399(.A1(new_n13692_), .A2(new_n13687_), .ZN(new_n13693_));
  OAI22_X1   g13400(.A1(new_n1347_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n1344_), .ZN(new_n13694_));
  OAI21_X1   g13401(.A1(new_n6229_), .A2(new_n1457_), .B(new_n13694_), .ZN(new_n13695_));
  AOI21_X1   g13402(.A1(new_n13695_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n13696_));
  XOR2_X1    g13403(.A1(new_n6851_), .A2(new_n13696_), .Z(new_n13697_));
  NOR3_X1    g13404(.A1(new_n13684_), .A2(new_n13693_), .A3(new_n13697_), .ZN(new_n13698_));
  NAND2_X1   g13405(.A1(new_n13692_), .A2(new_n13687_), .ZN(new_n13699_));
  NAND2_X1   g13406(.A1(new_n13683_), .A2(new_n13427_), .ZN(new_n13700_));
  INV_X1     g13407(.I(new_n13697_), .ZN(new_n13701_));
  AOI21_X1   g13408(.A1(new_n13700_), .A2(new_n13699_), .B(new_n13701_), .ZN(new_n13702_));
  OAI21_X1   g13409(.A1(new_n13698_), .A2(new_n13702_), .B(new_n13422_), .ZN(new_n13703_));
  NOR3_X1    g13410(.A1(new_n13290_), .A2(new_n13291_), .A3(new_n12873_), .ZN(new_n13704_));
  NOR2_X1    g13411(.A1(new_n13704_), .A2(new_n13287_), .ZN(new_n13705_));
  AOI21_X1   g13412(.A1(new_n13705_), .A2(new_n12881_), .B(new_n13418_), .ZN(new_n13706_));
  OAI21_X1   g13413(.A1(new_n13684_), .A2(new_n13693_), .B(new_n13701_), .ZN(new_n13707_));
  NAND3_X1   g13414(.A1(new_n13700_), .A2(new_n13699_), .A3(new_n13697_), .ZN(new_n13708_));
  NAND2_X1   g13415(.A1(new_n13707_), .A2(new_n13708_), .ZN(new_n13709_));
  NAND2_X1   g13416(.A1(new_n13706_), .A2(new_n13709_), .ZN(new_n13710_));
  OAI22_X1   g13417(.A1(new_n1055_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n1061_), .ZN(new_n13711_));
  OAI21_X1   g13418(.A1(new_n7198_), .A2(new_n1332_), .B(new_n13711_), .ZN(new_n13712_));
  AOI21_X1   g13419(.A1(new_n13712_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n13713_));
  XNOR2_X1   g13420(.A1(new_n7874_), .A2(new_n13713_), .ZN(new_n13714_));
  INV_X1     g13421(.I(new_n13714_), .ZN(new_n13715_));
  NAND3_X1   g13422(.A1(new_n13703_), .A2(new_n13710_), .A3(new_n13715_), .ZN(new_n13716_));
  INV_X1     g13423(.I(new_n13698_), .ZN(new_n13717_));
  INV_X1     g13424(.I(new_n13702_), .ZN(new_n13718_));
  AOI21_X1   g13425(.A1(new_n13717_), .A2(new_n13718_), .B(new_n13706_), .ZN(new_n13719_));
  AOI21_X1   g13426(.A1(new_n13707_), .A2(new_n13708_), .B(new_n13422_), .ZN(new_n13720_));
  OAI21_X1   g13427(.A1(new_n13720_), .A2(new_n13719_), .B(new_n13714_), .ZN(new_n13721_));
  NAND2_X1   g13428(.A1(new_n13721_), .A2(new_n13716_), .ZN(new_n13722_));
  NAND2_X1   g13429(.A1(new_n13417_), .A2(new_n13722_), .ZN(new_n13723_));
  INV_X1     g13430(.I(new_n13723_), .ZN(new_n13724_));
  NAND2_X1   g13431(.A1(new_n13703_), .A2(new_n13710_), .ZN(new_n13725_));
  NAND2_X1   g13432(.A1(new_n13725_), .A2(new_n13715_), .ZN(new_n13726_));
  NAND3_X1   g13433(.A1(new_n13703_), .A2(new_n13710_), .A3(new_n13714_), .ZN(new_n13727_));
  AOI21_X1   g13434(.A1(new_n13726_), .A2(new_n13727_), .B(new_n13417_), .ZN(new_n13728_));
  OAI22_X1   g13435(.A1(new_n970_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n820_), .ZN(new_n13729_));
  OAI21_X1   g13436(.A1(new_n8218_), .A2(new_n894_), .B(new_n13729_), .ZN(new_n13730_));
  AOI21_X1   g13437(.A1(new_n13730_), .A2(new_n827_), .B(new_n970_), .ZN(new_n13731_));
  XOR2_X1    g13438(.A1(new_n8952_), .A2(new_n13731_), .Z(new_n13732_));
  INV_X1     g13439(.I(new_n13732_), .ZN(new_n13733_));
  OAI21_X1   g13440(.A1(new_n13724_), .A2(new_n13728_), .B(new_n13733_), .ZN(new_n13734_));
  NOR2_X1    g13441(.A1(new_n13415_), .A2(new_n13311_), .ZN(new_n13735_));
  NOR2_X1    g13442(.A1(new_n13735_), .A2(new_n13310_), .ZN(new_n13736_));
  NAND2_X1   g13443(.A1(new_n13726_), .A2(new_n13727_), .ZN(new_n13737_));
  NAND2_X1   g13444(.A1(new_n13736_), .A2(new_n13737_), .ZN(new_n13738_));
  NAND3_X1   g13445(.A1(new_n13738_), .A2(new_n13723_), .A3(new_n13732_), .ZN(new_n13739_));
  NAND2_X1   g13446(.A1(new_n13734_), .A2(new_n13739_), .ZN(new_n13740_));
  NAND2_X1   g13447(.A1(new_n13414_), .A2(new_n13740_), .ZN(new_n13741_));
  AOI21_X1   g13448(.A1(new_n12911_), .A2(new_n12444_), .B(new_n12458_), .ZN(new_n13742_));
  NAND3_X1   g13449(.A1(new_n12910_), .A2(new_n12903_), .A3(new_n12443_), .ZN(new_n13743_));
  NAND2_X1   g13450(.A1(new_n13743_), .A2(new_n12457_), .ZN(new_n13744_));
  NOR3_X1    g13451(.A1(new_n13742_), .A2(new_n13744_), .A3(new_n13314_), .ZN(new_n13745_));
  OAI21_X1   g13452(.A1(new_n13742_), .A2(new_n13744_), .B(new_n13314_), .ZN(new_n13746_));
  INV_X1     g13453(.I(new_n13413_), .ZN(new_n13747_));
  AOI21_X1   g13454(.A1(new_n13746_), .A2(new_n13747_), .B(new_n13745_), .ZN(new_n13748_));
  NAND3_X1   g13455(.A1(new_n13738_), .A2(new_n13723_), .A3(new_n13733_), .ZN(new_n13749_));
  OAI21_X1   g13456(.A1(new_n13724_), .A2(new_n13728_), .B(new_n13732_), .ZN(new_n13750_));
  NAND2_X1   g13457(.A1(new_n13750_), .A2(new_n13749_), .ZN(new_n13751_));
  NAND2_X1   g13458(.A1(new_n13751_), .A2(new_n13748_), .ZN(new_n13752_));
  NAND2_X1   g13459(.A1(new_n13741_), .A2(new_n13752_), .ZN(new_n13753_));
  OAI22_X1   g13460(.A1(new_n607_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n610_), .ZN(new_n13754_));
  OAI21_X1   g13461(.A1(new_n9295_), .A2(new_n684_), .B(new_n13754_), .ZN(new_n13755_));
  AOI21_X1   g13462(.A1(new_n13755_), .A2(new_n612_), .B(new_n607_), .ZN(new_n13756_));
  XNOR2_X1   g13463(.A1(new_n10035_), .A2(new_n13756_), .ZN(new_n13757_));
  INV_X1     g13464(.I(new_n13757_), .ZN(new_n13758_));
  NAND2_X1   g13465(.A1(new_n13753_), .A2(new_n13758_), .ZN(new_n13759_));
  INV_X1     g13466(.I(new_n13759_), .ZN(new_n13760_));
  NOR2_X1    g13467(.A1(new_n13753_), .A2(new_n13758_), .ZN(new_n13761_));
  NOR2_X1    g13468(.A1(new_n13760_), .A2(new_n13761_), .ZN(new_n13762_));
  XOR2_X1    g13469(.A1(new_n13753_), .A2(new_n13758_), .Z(new_n13763_));
  NAND2_X1   g13470(.A1(new_n13406_), .A2(new_n13763_), .ZN(new_n13764_));
  OAI21_X1   g13471(.A1(new_n13406_), .A2(new_n13762_), .B(new_n13764_), .ZN(new_n13765_));
  OAI22_X1   g13472(.A1(new_n448_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n450_), .ZN(new_n13766_));
  OAI21_X1   g13473(.A1(new_n10477_), .A2(new_n496_), .B(new_n13766_), .ZN(new_n13767_));
  AOI21_X1   g13474(.A1(new_n13767_), .A2(new_n452_), .B(new_n448_), .ZN(new_n13768_));
  XOR2_X1    g13475(.A1(new_n11298_), .A2(new_n13768_), .Z(new_n13769_));
  NOR2_X1    g13476(.A1(new_n13765_), .A2(new_n13769_), .ZN(new_n13770_));
  NOR2_X1    g13477(.A1(new_n13762_), .A2(new_n13406_), .ZN(new_n13771_));
  AOI21_X1   g13478(.A1(new_n13406_), .A2(new_n13763_), .B(new_n13771_), .ZN(new_n13772_));
  INV_X1     g13479(.I(new_n13769_), .ZN(new_n13773_));
  NOR2_X1    g13480(.A1(new_n13772_), .A2(new_n13773_), .ZN(new_n13774_));
  NOR2_X1    g13481(.A1(new_n13774_), .A2(new_n13770_), .ZN(new_n13775_));
  NOR2_X1    g13482(.A1(new_n13348_), .A2(new_n13350_), .ZN(new_n13776_));
  NOR2_X1    g13483(.A1(new_n13340_), .A2(new_n13335_), .ZN(new_n13777_));
  INV_X1     g13484(.I(new_n13777_), .ZN(new_n13778_));
  AOI21_X1   g13485(.A1(new_n13777_), .A2(new_n12958_), .B(new_n13344_), .ZN(new_n13779_));
  AOI22_X1   g13486(.A1(new_n13776_), .A2(new_n13779_), .B1(new_n12949_), .B2(new_n13778_), .ZN(new_n13780_));
  XNOR2_X1   g13487(.A1(new_n13775_), .A2(new_n13780_), .ZN(new_n13781_));
  XNOR2_X1   g13488(.A1(\b[59] ), .A2(\b[61] ), .ZN(new_n13782_));
  NOR2_X1    g13489(.A1(new_n13782_), .A2(new_n13366_), .ZN(new_n13783_));
  XOR2_X1    g13490(.A1(new_n13365_), .A2(new_n13783_), .Z(new_n13784_));
  INV_X1     g13491(.I(\b[61] ), .ZN(new_n13785_));
  OAI22_X1   g13492(.A1(new_n330_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n263_), .ZN(new_n13786_));
  OAI21_X1   g13493(.A1(new_n12970_), .A2(new_n289_), .B(new_n13786_), .ZN(new_n13787_));
  AOI21_X1   g13494(.A1(new_n13787_), .A2(new_n260_), .B(new_n426_), .ZN(new_n13788_));
  XOR2_X1    g13495(.A1(new_n13784_), .A2(new_n13788_), .Z(new_n13789_));
  OAI22_X1   g13496(.A1(new_n12536_), .A2(new_n341_), .B1(new_n404_), .B2(new_n12542_), .ZN(new_n13790_));
  OAI21_X1   g13497(.A1(new_n11744_), .A2(new_n366_), .B(new_n13790_), .ZN(new_n13791_));
  AOI21_X1   g13498(.A1(new_n13791_), .A2(new_n334_), .B(new_n341_), .ZN(new_n13792_));
  XNOR2_X1   g13499(.A1(new_n12546_), .A2(new_n13792_), .ZN(new_n13793_));
  XNOR2_X1   g13500(.A1(new_n13789_), .A2(new_n13793_), .ZN(new_n13794_));
  NOR2_X1    g13501(.A1(new_n13781_), .A2(new_n13794_), .ZN(new_n13795_));
  NOR2_X1    g13502(.A1(new_n13789_), .A2(new_n13793_), .ZN(new_n13796_));
  INV_X1     g13503(.I(new_n13796_), .ZN(new_n13797_));
  NAND2_X1   g13504(.A1(new_n13789_), .A2(new_n13793_), .ZN(new_n13798_));
  NAND2_X1   g13505(.A1(new_n13797_), .A2(new_n13798_), .ZN(new_n13799_));
  AOI21_X1   g13506(.A1(new_n13781_), .A2(new_n13799_), .B(new_n13795_), .ZN(new_n13800_));
  NOR2_X1    g13507(.A1(new_n13375_), .A2(new_n13023_), .ZN(new_n13801_));
  AOI21_X1   g13508(.A1(new_n13023_), .A2(new_n13375_), .B(new_n13358_), .ZN(new_n13802_));
  NOR2_X1    g13509(.A1(new_n13802_), .A2(new_n13801_), .ZN(new_n13803_));
  NOR2_X1    g13510(.A1(new_n13800_), .A2(new_n13803_), .ZN(new_n13804_));
  XOR2_X1    g13511(.A1(new_n13804_), .A2(new_n13404_), .Z(new_n13805_));
  XOR2_X1    g13512(.A1(new_n13805_), .A2(new_n13402_), .Z(\f[61] ));
  AOI21_X1   g13513(.A1(new_n13005_), .A2(new_n13006_), .B(new_n13002_), .ZN(new_n13807_));
  NOR3_X1    g13514(.A1(new_n12994_), .A2(new_n12577_), .A3(new_n13000_), .ZN(new_n13808_));
  NOR2_X1    g13515(.A1(new_n13807_), .A2(new_n13808_), .ZN(new_n13809_));
  NAND2_X1   g13516(.A1(new_n13018_), .A2(new_n13002_), .ZN(new_n13810_));
  AOI21_X1   g13517(.A1(new_n12500_), .A2(new_n13016_), .B(new_n13810_), .ZN(new_n13811_));
  AOI21_X1   g13518(.A1(new_n13389_), .A2(new_n13390_), .B(new_n13388_), .ZN(new_n13812_));
  NOR3_X1    g13519(.A1(new_n13380_), .A2(new_n13386_), .A3(new_n13023_), .ZN(new_n13813_));
  OAI21_X1   g13520(.A1(new_n13812_), .A2(new_n13813_), .B(new_n13811_), .ZN(new_n13814_));
  AOI21_X1   g13521(.A1(new_n13814_), .A2(new_n13809_), .B(new_n13015_), .ZN(new_n13815_));
  INV_X1     g13522(.I(new_n13800_), .ZN(new_n13816_));
  NAND2_X1   g13523(.A1(new_n13815_), .A2(new_n13816_), .ZN(new_n13817_));
  NOR2_X1    g13524(.A1(new_n13402_), .A2(new_n13803_), .ZN(new_n13818_));
  OAI21_X1   g13525(.A1(new_n13815_), .A2(new_n13816_), .B(new_n13818_), .ZN(new_n13819_));
  NAND2_X1   g13526(.A1(new_n13819_), .A2(new_n13817_), .ZN(new_n13820_));
  AOI21_X1   g13527(.A1(new_n13781_), .A2(new_n13798_), .B(new_n13796_), .ZN(new_n13821_));
  INV_X1     g13528(.I(new_n13821_), .ZN(new_n13822_));
  NAND2_X1   g13529(.A1(new_n13772_), .A2(new_n13773_), .ZN(new_n13823_));
  OAI21_X1   g13530(.A1(new_n13780_), .A2(new_n13774_), .B(new_n13823_), .ZN(new_n13824_));
  XOR2_X1    g13531(.A1(new_n13753_), .A2(new_n13757_), .Z(new_n13825_));
  AOI21_X1   g13532(.A1(new_n13036_), .A2(new_n13314_), .B(new_n13413_), .ZN(new_n13826_));
  OAI21_X1   g13533(.A1(new_n13826_), .A2(new_n13745_), .B(new_n13750_), .ZN(new_n13827_));
  NOR3_X1    g13534(.A1(new_n13720_), .A2(new_n13719_), .A3(new_n13714_), .ZN(new_n13828_));
  AOI21_X1   g13535(.A1(new_n13703_), .A2(new_n13710_), .B(new_n13715_), .ZN(new_n13829_));
  NOR2_X1    g13536(.A1(new_n13828_), .A2(new_n13829_), .ZN(new_n13830_));
  NOR2_X1    g13537(.A1(new_n13720_), .A2(new_n13719_), .ZN(new_n13831_));
  NOR2_X1    g13538(.A1(new_n13831_), .A2(new_n13714_), .ZN(new_n13832_));
  AOI21_X1   g13539(.A1(new_n13422_), .A2(new_n13718_), .B(new_n13698_), .ZN(new_n13833_));
  NAND2_X1   g13540(.A1(new_n13427_), .A2(new_n13667_), .ZN(new_n13834_));
  XOR2_X1    g13541(.A1(new_n13678_), .A2(new_n13662_), .Z(new_n13835_));
  OAI21_X1   g13542(.A1(new_n13427_), .A2(new_n13667_), .B(new_n13835_), .ZN(new_n13836_));
  NOR2_X1    g13543(.A1(new_n13645_), .A2(new_n13631_), .ZN(new_n13837_));
  OAI22_X1   g13544(.A1(new_n3709_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n3717_), .ZN(new_n13838_));
  OAI21_X1   g13545(.A1(new_n3260_), .A2(new_n3569_), .B(new_n13838_), .ZN(new_n13839_));
  AOI21_X1   g13546(.A1(new_n13839_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n13840_));
  XOR2_X1    g13547(.A1(new_n3722_), .A2(new_n13840_), .Z(new_n13841_));
  INV_X1     g13548(.I(new_n13841_), .ZN(new_n13842_));
  NAND2_X1   g13549(.A1(new_n13444_), .A2(new_n13442_), .ZN(new_n13843_));
  NAND2_X1   g13550(.A1(new_n13843_), .A2(new_n13624_), .ZN(new_n13844_));
  XOR2_X1    g13551(.A1(new_n13610_), .A2(new_n13441_), .Z(new_n13845_));
  OAI21_X1   g13552(.A1(new_n13843_), .A2(new_n13624_), .B(new_n13845_), .ZN(new_n13846_));
  NOR2_X1    g13553(.A1(new_n13595_), .A2(new_n13596_), .ZN(new_n13847_));
  AOI21_X1   g13554(.A1(new_n13586_), .A2(new_n13590_), .B(new_n13577_), .ZN(new_n13848_));
  OR2_X2     g13555(.A1(new_n13592_), .A2(new_n13593_), .Z(new_n13849_));
  AOI21_X1   g13556(.A1(new_n13849_), .A2(new_n13577_), .B(new_n13848_), .ZN(new_n13850_));
  NOR2_X1    g13557(.A1(new_n13850_), .A2(new_n13602_), .ZN(new_n13851_));
  OAI21_X1   g13558(.A1(new_n13851_), .A2(new_n13847_), .B(new_n13600_), .ZN(new_n13852_));
  OAI21_X1   g13559(.A1(new_n13574_), .A2(new_n13573_), .B(new_n13575_), .ZN(new_n13853_));
  NAND3_X1   g13560(.A1(new_n13561_), .A2(new_n13567_), .A3(new_n13571_), .ZN(new_n13854_));
  NAND2_X1   g13561(.A1(new_n13853_), .A2(new_n13854_), .ZN(new_n13855_));
  NOR2_X1    g13562(.A1(new_n13855_), .A2(new_n13589_), .ZN(new_n13856_));
  NOR2_X1    g13563(.A1(new_n13577_), .A2(new_n13580_), .ZN(new_n13857_));
  OAI21_X1   g13564(.A1(new_n13857_), .A2(new_n13856_), .B(new_n13584_), .ZN(new_n13858_));
  AOI21_X1   g13565(.A1(new_n13579_), .A2(new_n13578_), .B(new_n13576_), .ZN(new_n13859_));
  NOR2_X1    g13566(.A1(new_n13551_), .A2(new_n13540_), .ZN(new_n13860_));
  NOR2_X1    g13567(.A1(new_n13860_), .A2(new_n13163_), .ZN(new_n13861_));
  INV_X1     g13568(.I(new_n13861_), .ZN(new_n13862_));
  AOI21_X1   g13569(.A1(new_n13860_), .A2(new_n13163_), .B(new_n13555_), .ZN(new_n13863_));
  NAND2_X1   g13570(.A1(new_n13445_), .A2(new_n13863_), .ZN(new_n13864_));
  AOI21_X1   g13571(.A1(new_n13448_), .A2(new_n13446_), .B(new_n13549_), .ZN(new_n13865_));
  NOR2_X1    g13572(.A1(new_n13865_), .A2(new_n13542_), .ZN(new_n13866_));
  NAND3_X1   g13573(.A1(new_n13523_), .A2(new_n13515_), .A3(new_n13524_), .ZN(new_n13867_));
  OAI21_X1   g13574(.A1(new_n13527_), .A2(new_n13525_), .B(new_n13867_), .ZN(new_n13868_));
  INV_X1     g13575(.I(new_n13868_), .ZN(new_n13869_));
  INV_X1     g13576(.I(new_n13527_), .ZN(new_n13870_));
  OAI21_X1   g13577(.A1(new_n13516_), .A2(new_n13511_), .B(new_n13520_), .ZN(new_n13871_));
  NAND2_X1   g13578(.A1(new_n13870_), .A2(new_n13871_), .ZN(new_n13872_));
  AOI21_X1   g13579(.A1(new_n13522_), .A2(new_n13513_), .B(new_n13512_), .ZN(new_n13873_));
  INV_X1     g13580(.I(new_n13499_), .ZN(new_n13874_));
  AOI22_X1   g13581(.A1(new_n13458_), .A2(new_n13097_), .B1(new_n13490_), .B2(new_n13493_), .ZN(new_n13875_));
  NOR2_X1    g13582(.A1(new_n13487_), .A2(new_n13484_), .ZN(new_n13876_));
  NOR2_X1    g13583(.A1(new_n13876_), .A2(new_n13488_), .ZN(new_n13877_));
  NOR2_X1    g13584(.A1(new_n13479_), .A2(new_n13460_), .ZN(new_n13878_));
  INV_X1     g13585(.I(new_n13466_), .ZN(new_n13879_));
  INV_X1     g13586(.I(new_n13472_), .ZN(new_n13880_));
  XNOR2_X1   g13587(.A1(\a[59] ), .A2(\a[61] ), .ZN(new_n13881_));
  XNOR2_X1   g13588(.A1(\a[59] ), .A2(\a[62] ), .ZN(new_n13882_));
  XNOR2_X1   g13589(.A1(\a[59] ), .A2(\a[60] ), .ZN(new_n13883_));
  NOR3_X1    g13590(.A1(new_n13881_), .A2(new_n13882_), .A3(new_n13883_), .ZN(new_n13884_));
  INV_X1     g13591(.I(new_n13884_), .ZN(new_n13885_));
  OAI22_X1   g13592(.A1(new_n13880_), .A2(new_n10132_), .B1(new_n258_), .B2(new_n13885_), .ZN(new_n13886_));
  AOI21_X1   g13593(.A1(new_n13886_), .A2(new_n13476_), .B(new_n490_), .ZN(new_n13887_));
  XOR2_X1    g13594(.A1(new_n13887_), .A2(new_n13879_), .Z(new_n13888_));
  XOR2_X1    g13595(.A1(new_n13888_), .A2(new_n13878_), .Z(new_n13889_));
  AOI22_X1   g13596(.A1(new_n13078_), .A2(\b[3] ), .B1(new_n413_), .B2(new_n12218_), .ZN(new_n13890_));
  OAI21_X1   g13597(.A1(new_n13890_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n13891_));
  XOR2_X1    g13598(.A1(new_n13891_), .A2(new_n378_), .Z(new_n13892_));
  NOR2_X1    g13599(.A1(new_n13889_), .A2(new_n13892_), .ZN(new_n13893_));
  INV_X1     g13600(.I(new_n13893_), .ZN(new_n13894_));
  NAND2_X1   g13601(.A1(new_n13889_), .A2(new_n13892_), .ZN(new_n13895_));
  AOI21_X1   g13602(.A1(new_n13894_), .A2(new_n13895_), .B(new_n13877_), .ZN(new_n13896_));
  INV_X1     g13603(.I(new_n13877_), .ZN(new_n13897_));
  INV_X1     g13604(.I(new_n13892_), .ZN(new_n13898_));
  XOR2_X1    g13605(.A1(new_n13889_), .A2(new_n13898_), .Z(new_n13899_));
  NOR2_X1    g13606(.A1(new_n13897_), .A2(new_n13899_), .ZN(new_n13900_));
  AOI22_X1   g13607(.A1(new_n10969_), .A2(new_n517_), .B1(new_n11394_), .B2(\b[6] ), .ZN(new_n13901_));
  OAI21_X1   g13608(.A1(new_n13901_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n13902_));
  XOR2_X1    g13609(.A1(new_n522_), .A2(new_n13902_), .Z(new_n13903_));
  NOR3_X1    g13610(.A1(new_n13900_), .A2(new_n13896_), .A3(new_n13903_), .ZN(new_n13904_));
  NOR2_X1    g13611(.A1(new_n13900_), .A2(new_n13896_), .ZN(new_n13905_));
  INV_X1     g13612(.I(new_n13903_), .ZN(new_n13906_));
  NOR2_X1    g13613(.A1(new_n13905_), .A2(new_n13906_), .ZN(new_n13907_));
  OAI22_X1   g13614(.A1(new_n13907_), .A2(new_n13904_), .B1(new_n13875_), .B2(new_n13874_), .ZN(new_n13908_));
  NOR2_X1    g13615(.A1(new_n13875_), .A2(new_n13874_), .ZN(new_n13909_));
  OAI21_X1   g13616(.A1(new_n13900_), .A2(new_n13896_), .B(new_n13906_), .ZN(new_n13910_));
  INV_X1     g13617(.I(new_n13910_), .ZN(new_n13911_));
  NOR3_X1    g13618(.A1(new_n13900_), .A2(new_n13896_), .A3(new_n13906_), .ZN(new_n13912_));
  OAI21_X1   g13619(.A1(new_n13911_), .A2(new_n13912_), .B(new_n13909_), .ZN(new_n13913_));
  AOI22_X1   g13620(.A1(new_n11415_), .A2(new_n773_), .B1(\b[9] ), .B2(new_n10145_), .ZN(new_n13914_));
  OAI21_X1   g13621(.A1(new_n13914_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n13915_));
  XOR2_X1    g13622(.A1(new_n710_), .A2(new_n13915_), .Z(new_n13916_));
  AOI21_X1   g13623(.A1(new_n13913_), .A2(new_n13908_), .B(new_n13916_), .ZN(new_n13917_));
  INV_X1     g13624(.I(new_n13908_), .ZN(new_n13918_));
  NOR2_X1    g13625(.A1(new_n13911_), .A2(new_n13912_), .ZN(new_n13919_));
  NOR3_X1    g13626(.A1(new_n13919_), .A2(new_n13874_), .A3(new_n13875_), .ZN(new_n13920_));
  INV_X1     g13627(.I(new_n13916_), .ZN(new_n13921_));
  NOR3_X1    g13628(.A1(new_n13918_), .A2(new_n13920_), .A3(new_n13921_), .ZN(new_n13922_));
  NOR2_X1    g13629(.A1(new_n13922_), .A2(new_n13917_), .ZN(new_n13923_));
  NOR2_X1    g13630(.A1(new_n13873_), .A2(new_n13923_), .ZN(new_n13924_));
  INV_X1     g13631(.I(new_n13512_), .ZN(new_n13925_));
  OAI21_X1   g13632(.A1(new_n13457_), .A2(new_n13514_), .B(new_n13925_), .ZN(new_n13926_));
  OAI21_X1   g13633(.A1(new_n13918_), .A2(new_n13920_), .B(new_n13921_), .ZN(new_n13927_));
  NAND3_X1   g13634(.A1(new_n13913_), .A2(new_n13908_), .A3(new_n13916_), .ZN(new_n13928_));
  NAND2_X1   g13635(.A1(new_n13927_), .A2(new_n13928_), .ZN(new_n13929_));
  NOR2_X1    g13636(.A1(new_n13929_), .A2(new_n13926_), .ZN(new_n13930_));
  OAI22_X1   g13637(.A1(new_n8644_), .A2(new_n861_), .B1(new_n930_), .B2(new_n9388_), .ZN(new_n13931_));
  OAI21_X1   g13638(.A1(new_n780_), .A2(new_n10154_), .B(new_n13931_), .ZN(new_n13932_));
  AOI21_X1   g13639(.A1(new_n13932_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n13933_));
  XNOR2_X1   g13640(.A1(new_n937_), .A2(new_n13933_), .ZN(new_n13934_));
  NOR3_X1    g13641(.A1(new_n13924_), .A2(new_n13930_), .A3(new_n13934_), .ZN(new_n13935_));
  NAND2_X1   g13642(.A1(new_n13929_), .A2(new_n13926_), .ZN(new_n13936_));
  NAND2_X1   g13643(.A1(new_n13873_), .A2(new_n13923_), .ZN(new_n13937_));
  INV_X1     g13644(.I(new_n13934_), .ZN(new_n13938_));
  AOI21_X1   g13645(.A1(new_n13937_), .A2(new_n13936_), .B(new_n13938_), .ZN(new_n13939_));
  OAI22_X1   g13646(.A1(new_n7619_), .A2(new_n1109_), .B1(new_n1189_), .B2(new_n8309_), .ZN(new_n13940_));
  OAI21_X1   g13647(.A1(new_n1017_), .A2(new_n7947_), .B(new_n13940_), .ZN(new_n13941_));
  AOI21_X1   g13648(.A1(new_n13941_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n13942_));
  XNOR2_X1   g13649(.A1(new_n1196_), .A2(new_n13942_), .ZN(new_n13943_));
  INV_X1     g13650(.I(new_n13943_), .ZN(new_n13944_));
  OAI21_X1   g13651(.A1(new_n13935_), .A2(new_n13939_), .B(new_n13944_), .ZN(new_n13945_));
  NAND3_X1   g13652(.A1(new_n13937_), .A2(new_n13936_), .A3(new_n13938_), .ZN(new_n13946_));
  OAI21_X1   g13653(.A1(new_n13924_), .A2(new_n13930_), .B(new_n13934_), .ZN(new_n13947_));
  NAND3_X1   g13654(.A1(new_n13947_), .A2(new_n13946_), .A3(new_n13943_), .ZN(new_n13948_));
  AOI22_X1   g13655(.A1(new_n13872_), .A2(new_n13867_), .B1(new_n13945_), .B2(new_n13948_), .ZN(new_n13949_));
  NAND2_X1   g13656(.A1(new_n13947_), .A2(new_n13946_), .ZN(new_n13950_));
  XOR2_X1    g13657(.A1(new_n13950_), .A2(new_n13944_), .Z(new_n13951_));
  AOI21_X1   g13658(.A1(new_n13869_), .A2(new_n13951_), .B(new_n13949_), .ZN(new_n13952_));
  NOR2_X1    g13659(.A1(new_n13866_), .A2(new_n13952_), .ZN(new_n13953_));
  NAND2_X1   g13660(.A1(new_n13945_), .A2(new_n13948_), .ZN(new_n13954_));
  NAND2_X1   g13661(.A1(new_n13954_), .A2(new_n13868_), .ZN(new_n13955_));
  XOR2_X1    g13662(.A1(new_n13950_), .A2(new_n13943_), .Z(new_n13956_));
  OAI21_X1   g13663(.A1(new_n13956_), .A2(new_n13868_), .B(new_n13955_), .ZN(new_n13957_));
  NOR3_X1    g13664(.A1(new_n13957_), .A2(new_n13542_), .A3(new_n13865_), .ZN(new_n13958_));
  OAI22_X1   g13665(.A1(new_n6644_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n6647_), .ZN(new_n13959_));
  OAI21_X1   g13666(.A1(new_n1294_), .A2(new_n7284_), .B(new_n13959_), .ZN(new_n13960_));
  AOI21_X1   g13667(.A1(new_n13960_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n13961_));
  XOR2_X1    g13668(.A1(new_n1530_), .A2(new_n13961_), .Z(new_n13962_));
  INV_X1     g13669(.I(new_n13962_), .ZN(new_n13963_));
  OAI21_X1   g13670(.A1(new_n13953_), .A2(new_n13958_), .B(new_n13963_), .ZN(new_n13964_));
  OAI21_X1   g13671(.A1(new_n13865_), .A2(new_n13542_), .B(new_n13957_), .ZN(new_n13965_));
  NAND2_X1   g13672(.A1(new_n13866_), .A2(new_n13952_), .ZN(new_n13966_));
  NAND3_X1   g13673(.A1(new_n13966_), .A2(new_n13965_), .A3(new_n13962_), .ZN(new_n13967_));
  OAI22_X1   g13674(.A1(new_n5993_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n5991_), .ZN(new_n13968_));
  OAI21_X1   g13675(.A1(new_n1634_), .A2(new_n5997_), .B(new_n13968_), .ZN(new_n13969_));
  AOI21_X1   g13676(.A1(new_n13969_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n13970_));
  XNOR2_X1   g13677(.A1(new_n1940_), .A2(new_n13970_), .ZN(new_n13971_));
  INV_X1     g13678(.I(new_n13971_), .ZN(new_n13972_));
  NAND3_X1   g13679(.A1(new_n13967_), .A2(new_n13964_), .A3(new_n13972_), .ZN(new_n13973_));
  AOI21_X1   g13680(.A1(new_n13966_), .A2(new_n13965_), .B(new_n13962_), .ZN(new_n13974_));
  NOR3_X1    g13681(.A1(new_n13953_), .A2(new_n13958_), .A3(new_n13963_), .ZN(new_n13975_));
  OAI21_X1   g13682(.A1(new_n13974_), .A2(new_n13975_), .B(new_n13971_), .ZN(new_n13976_));
  AOI22_X1   g13683(.A1(new_n13976_), .A2(new_n13973_), .B1(new_n13862_), .B2(new_n13864_), .ZN(new_n13977_));
  INV_X1     g13684(.I(new_n13977_), .ZN(new_n13978_));
  OAI21_X1   g13685(.A1(new_n13974_), .A2(new_n13975_), .B(new_n13972_), .ZN(new_n13979_));
  NAND3_X1   g13686(.A1(new_n13967_), .A2(new_n13964_), .A3(new_n13971_), .ZN(new_n13980_));
  NAND2_X1   g13687(.A1(new_n13979_), .A2(new_n13980_), .ZN(new_n13981_));
  NAND3_X1   g13688(.A1(new_n13981_), .A2(new_n13862_), .A3(new_n13864_), .ZN(new_n13982_));
  NAND2_X1   g13689(.A1(new_n13978_), .A2(new_n13982_), .ZN(new_n13983_));
  OAI21_X1   g13690(.A1(new_n13859_), .A2(new_n13572_), .B(new_n13983_), .ZN(new_n13984_));
  OAI21_X1   g13691(.A1(new_n13172_), .A2(new_n13588_), .B(new_n13854_), .ZN(new_n13985_));
  INV_X1     g13692(.I(new_n13864_), .ZN(new_n13986_));
  NOR2_X1    g13693(.A1(new_n13986_), .A2(new_n13861_), .ZN(new_n13987_));
  AOI21_X1   g13694(.A1(new_n13987_), .A2(new_n13981_), .B(new_n13977_), .ZN(new_n13988_));
  NAND3_X1   g13695(.A1(new_n13985_), .A2(new_n13853_), .A3(new_n13988_), .ZN(new_n13989_));
  OAI22_X1   g13696(.A1(new_n5420_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n5107_), .ZN(new_n13990_));
  OAI21_X1   g13697(.A1(new_n2102_), .A2(new_n5112_), .B(new_n13990_), .ZN(new_n13991_));
  AOI21_X1   g13698(.A1(new_n13991_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n13992_));
  XNOR2_X1   g13699(.A1(new_n2443_), .A2(new_n13992_), .ZN(new_n13993_));
  INV_X1     g13700(.I(new_n13993_), .ZN(new_n13994_));
  NAND3_X1   g13701(.A1(new_n13984_), .A2(new_n13989_), .A3(new_n13994_), .ZN(new_n13995_));
  AOI21_X1   g13702(.A1(new_n13985_), .A2(new_n13853_), .B(new_n13988_), .ZN(new_n13996_));
  NOR3_X1    g13703(.A1(new_n13859_), .A2(new_n13983_), .A3(new_n13572_), .ZN(new_n13997_));
  OAI21_X1   g13704(.A1(new_n13997_), .A2(new_n13996_), .B(new_n13993_), .ZN(new_n13998_));
  NAND3_X1   g13705(.A1(new_n13998_), .A2(new_n13995_), .A3(new_n13858_), .ZN(new_n13999_));
  NAND3_X1   g13706(.A1(new_n13999_), .A2(new_n13602_), .A3(new_n13850_), .ZN(new_n14000_));
  NAND2_X1   g13707(.A1(new_n13577_), .A2(new_n13580_), .ZN(new_n14001_));
  NAND2_X1   g13708(.A1(new_n13855_), .A2(new_n13589_), .ZN(new_n14002_));
  AOI21_X1   g13709(.A1(new_n14001_), .A2(new_n14002_), .B(new_n13585_), .ZN(new_n14003_));
  NOR3_X1    g13710(.A1(new_n13997_), .A2(new_n13996_), .A3(new_n13993_), .ZN(new_n14004_));
  AOI21_X1   g13711(.A1(new_n13984_), .A2(new_n13989_), .B(new_n13994_), .ZN(new_n14005_));
  NOR3_X1    g13712(.A1(new_n14004_), .A2(new_n14005_), .A3(new_n14003_), .ZN(new_n14006_));
  OAI21_X1   g13713(.A1(new_n14006_), .A2(new_n13596_), .B(new_n13595_), .ZN(new_n14007_));
  OAI22_X1   g13714(.A1(new_n4072_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n4067_), .ZN(new_n14008_));
  OAI21_X1   g13715(.A1(new_n2643_), .A2(new_n4318_), .B(new_n14008_), .ZN(new_n14009_));
  AOI21_X1   g13716(.A1(new_n14009_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n14010_));
  XNOR2_X1   g13717(.A1(new_n3022_), .A2(new_n14010_), .ZN(new_n14011_));
  INV_X1     g13718(.I(new_n14011_), .ZN(new_n14012_));
  NAND3_X1   g13719(.A1(new_n14007_), .A2(new_n14000_), .A3(new_n14012_), .ZN(new_n14013_));
  NOR3_X1    g13720(.A1(new_n14006_), .A2(new_n13595_), .A3(new_n13596_), .ZN(new_n14014_));
  AOI21_X1   g13721(.A1(new_n13999_), .A2(new_n13602_), .B(new_n13850_), .ZN(new_n14015_));
  OAI21_X1   g13722(.A1(new_n14014_), .A2(new_n14015_), .B(new_n14011_), .ZN(new_n14016_));
  NAND3_X1   g13723(.A1(new_n14016_), .A2(new_n14013_), .A3(new_n13852_), .ZN(new_n14017_));
  NAND3_X1   g13724(.A1(new_n14017_), .A2(new_n13619_), .A3(new_n13610_), .ZN(new_n14018_));
  NAND2_X1   g13725(.A1(new_n13850_), .A2(new_n13602_), .ZN(new_n14019_));
  NAND2_X1   g13726(.A1(new_n13595_), .A2(new_n13596_), .ZN(new_n14020_));
  AOI21_X1   g13727(.A1(new_n14019_), .A2(new_n14020_), .B(new_n13603_), .ZN(new_n14021_));
  NOR3_X1    g13728(.A1(new_n14014_), .A2(new_n14015_), .A3(new_n14011_), .ZN(new_n14022_));
  AOI21_X1   g13729(.A1(new_n14007_), .A2(new_n14000_), .B(new_n14012_), .ZN(new_n14023_));
  NOR3_X1    g13730(.A1(new_n14022_), .A2(new_n14023_), .A3(new_n14021_), .ZN(new_n14024_));
  OAI21_X1   g13731(.A1(new_n14024_), .A2(new_n13616_), .B(new_n13441_), .ZN(new_n14025_));
  OAI22_X1   g13732(.A1(new_n4253_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n4500_), .ZN(new_n14026_));
  OAI21_X1   g13733(.A1(new_n3989_), .A2(new_n2884_), .B(new_n14026_), .ZN(new_n14027_));
  AOI21_X1   g13734(.A1(new_n14027_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n14028_));
  XOR2_X1    g13735(.A1(new_n4499_), .A2(new_n14028_), .Z(new_n14029_));
  INV_X1     g13736(.I(new_n14029_), .ZN(new_n14030_));
  NAND3_X1   g13737(.A1(new_n14025_), .A2(new_n14018_), .A3(new_n14030_), .ZN(new_n14031_));
  NOR3_X1    g13738(.A1(new_n14024_), .A2(new_n13616_), .A3(new_n13441_), .ZN(new_n14032_));
  AOI21_X1   g13739(.A1(new_n14017_), .A2(new_n13610_), .B(new_n13619_), .ZN(new_n14033_));
  OAI21_X1   g13740(.A1(new_n14032_), .A2(new_n14033_), .B(new_n14029_), .ZN(new_n14034_));
  NAND2_X1   g13741(.A1(new_n14034_), .A2(new_n14031_), .ZN(new_n14035_));
  NAND3_X1   g13742(.A1(new_n13846_), .A2(new_n13844_), .A3(new_n14035_), .ZN(new_n14036_));
  NOR2_X1    g13743(.A1(new_n13614_), .A2(new_n13612_), .ZN(new_n14037_));
  NOR2_X1    g13744(.A1(new_n14037_), .A2(new_n13437_), .ZN(new_n14038_));
  XOR2_X1    g13745(.A1(new_n13616_), .A2(new_n13441_), .Z(new_n14039_));
  AOI21_X1   g13746(.A1(new_n14037_), .A2(new_n13437_), .B(new_n14039_), .ZN(new_n14040_));
  NOR3_X1    g13747(.A1(new_n14032_), .A2(new_n14033_), .A3(new_n14029_), .ZN(new_n14041_));
  AOI21_X1   g13748(.A1(new_n14025_), .A2(new_n14018_), .B(new_n14030_), .ZN(new_n14042_));
  NOR2_X1    g13749(.A1(new_n14041_), .A2(new_n14042_), .ZN(new_n14043_));
  OAI21_X1   g13750(.A1(new_n14040_), .A2(new_n14038_), .B(new_n14043_), .ZN(new_n14044_));
  AOI21_X1   g13751(.A1(new_n14044_), .A2(new_n14036_), .B(new_n13842_), .ZN(new_n14045_));
  NOR3_X1    g13752(.A1(new_n14040_), .A2(new_n14038_), .A3(new_n14043_), .ZN(new_n14046_));
  AOI21_X1   g13753(.A1(new_n13846_), .A2(new_n13844_), .B(new_n14035_), .ZN(new_n14047_));
  NOR3_X1    g13754(.A1(new_n14046_), .A2(new_n14047_), .A3(new_n13841_), .ZN(new_n14048_));
  NOR2_X1    g13755(.A1(new_n14048_), .A2(new_n14045_), .ZN(new_n14049_));
  NOR3_X1    g13756(.A1(new_n13674_), .A2(new_n13837_), .A3(new_n14049_), .ZN(new_n14050_));
  NOR2_X1    g13757(.A1(new_n13645_), .A2(new_n13631_), .ZN(new_n14052_));
  OAI21_X1   g13758(.A1(new_n14050_), .A2(new_n14052_), .B(new_n13642_), .ZN(new_n14053_));
  OAI21_X1   g13759(.A1(new_n14046_), .A2(new_n14047_), .B(new_n13841_), .ZN(new_n14054_));
  NAND3_X1   g13760(.A1(new_n14044_), .A2(new_n14036_), .A3(new_n13842_), .ZN(new_n14055_));
  NAND2_X1   g13761(.A1(new_n14054_), .A2(new_n14055_), .ZN(new_n14056_));
  NAND3_X1   g13762(.A1(new_n13637_), .A2(new_n13644_), .A3(new_n14056_), .ZN(new_n14057_));
  INV_X1     g13763(.I(new_n14052_), .ZN(new_n14058_));
  NAND3_X1   g13764(.A1(new_n14057_), .A2(new_n13433_), .A3(new_n14058_), .ZN(new_n14059_));
  OAI22_X1   g13765(.A1(new_n2171_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n2166_), .ZN(new_n14060_));
  OAI21_X1   g13766(.A1(new_n4774_), .A2(new_n2322_), .B(new_n14060_), .ZN(new_n14061_));
  AOI21_X1   g13767(.A1(new_n14061_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n14062_));
  XNOR2_X1   g13768(.A1(new_n5357_), .A2(new_n14062_), .ZN(new_n14063_));
  INV_X1     g13769(.I(new_n14063_), .ZN(new_n14064_));
  NAND3_X1   g13770(.A1(new_n14053_), .A2(new_n14059_), .A3(new_n14064_), .ZN(new_n14065_));
  AOI21_X1   g13771(.A1(new_n14057_), .A2(new_n14058_), .B(new_n13433_), .ZN(new_n14066_));
  NOR3_X1    g13772(.A1(new_n14050_), .A2(new_n13642_), .A3(new_n14052_), .ZN(new_n14067_));
  OAI21_X1   g13773(.A1(new_n14067_), .A2(new_n14066_), .B(new_n14063_), .ZN(new_n14068_));
  NAND3_X1   g13774(.A1(new_n14068_), .A2(new_n14065_), .A3(new_n13677_), .ZN(new_n14069_));
  NAND3_X1   g13775(.A1(new_n14069_), .A2(new_n13657_), .A3(new_n13662_), .ZN(new_n14070_));
  INV_X1     g13776(.I(new_n13662_), .ZN(new_n14071_));
  NOR3_X1    g13777(.A1(new_n14067_), .A2(new_n14066_), .A3(new_n14063_), .ZN(new_n14072_));
  AOI21_X1   g13778(.A1(new_n14053_), .A2(new_n14059_), .B(new_n14064_), .ZN(new_n14073_));
  NOR3_X1    g13779(.A1(new_n14072_), .A2(new_n14073_), .A3(new_n13656_), .ZN(new_n14074_));
  OAI21_X1   g13780(.A1(new_n14074_), .A2(new_n14071_), .B(new_n13678_), .ZN(new_n14075_));
  OAI22_X1   g13781(.A1(new_n1712_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n1707_), .ZN(new_n14076_));
  OAI21_X1   g13782(.A1(new_n5913_), .A2(new_n1850_), .B(new_n14076_), .ZN(new_n14077_));
  AOI21_X1   g13783(.A1(new_n14077_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n14078_));
  XOR2_X1    g13784(.A1(new_n6233_), .A2(new_n14078_), .Z(new_n14079_));
  INV_X1     g13785(.I(new_n14079_), .ZN(new_n14080_));
  NAND3_X1   g13786(.A1(new_n14075_), .A2(new_n14070_), .A3(new_n14080_), .ZN(new_n14081_));
  NOR3_X1    g13787(.A1(new_n14074_), .A2(new_n13678_), .A3(new_n14071_), .ZN(new_n14082_));
  AOI21_X1   g13788(.A1(new_n14069_), .A2(new_n13662_), .B(new_n13657_), .ZN(new_n14083_));
  OAI21_X1   g13789(.A1(new_n14082_), .A2(new_n14083_), .B(new_n14079_), .ZN(new_n14084_));
  AOI22_X1   g13790(.A1(new_n13836_), .A2(new_n13834_), .B1(new_n14081_), .B2(new_n14084_), .ZN(new_n14085_));
  NOR2_X1    g13791(.A1(new_n13687_), .A2(new_n13666_), .ZN(new_n14086_));
  XOR2_X1    g13792(.A1(new_n13678_), .A2(new_n14071_), .Z(new_n14087_));
  AOI21_X1   g13793(.A1(new_n13687_), .A2(new_n13666_), .B(new_n14087_), .ZN(new_n14088_));
  AOI21_X1   g13794(.A1(new_n14075_), .A2(new_n14070_), .B(new_n14079_), .ZN(new_n14089_));
  NOR3_X1    g13795(.A1(new_n14082_), .A2(new_n14083_), .A3(new_n14080_), .ZN(new_n14090_));
  NOR2_X1    g13796(.A1(new_n14090_), .A2(new_n14089_), .ZN(new_n14091_));
  NOR3_X1    g13797(.A1(new_n14091_), .A2(new_n14086_), .A3(new_n14088_), .ZN(new_n14092_));
  OAI22_X1   g13798(.A1(new_n1347_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n1344_), .ZN(new_n14093_));
  OAI21_X1   g13799(.A1(new_n6538_), .A2(new_n1457_), .B(new_n14093_), .ZN(new_n14094_));
  AOI21_X1   g13800(.A1(new_n14094_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n14095_));
  XNOR2_X1   g13801(.A1(new_n7202_), .A2(new_n14095_), .ZN(new_n14096_));
  INV_X1     g13802(.I(new_n14096_), .ZN(new_n14097_));
  OAI21_X1   g13803(.A1(new_n14092_), .A2(new_n14085_), .B(new_n14097_), .ZN(new_n14098_));
  NOR3_X1    g13804(.A1(new_n14082_), .A2(new_n14083_), .A3(new_n14079_), .ZN(new_n14099_));
  AOI21_X1   g13805(.A1(new_n14075_), .A2(new_n14070_), .B(new_n14080_), .ZN(new_n14100_));
  OAI22_X1   g13806(.A1(new_n14088_), .A2(new_n14086_), .B1(new_n14099_), .B2(new_n14100_), .ZN(new_n14101_));
  OAI21_X1   g13807(.A1(new_n14082_), .A2(new_n14083_), .B(new_n14080_), .ZN(new_n14102_));
  NAND3_X1   g13808(.A1(new_n14075_), .A2(new_n14070_), .A3(new_n14079_), .ZN(new_n14103_));
  NAND2_X1   g13809(.A1(new_n14102_), .A2(new_n14103_), .ZN(new_n14104_));
  NAND3_X1   g13810(.A1(new_n14104_), .A2(new_n13836_), .A3(new_n13834_), .ZN(new_n14105_));
  NAND3_X1   g13811(.A1(new_n14105_), .A2(new_n14101_), .A3(new_n14096_), .ZN(new_n14106_));
  OAI22_X1   g13812(.A1(new_n1055_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n1061_), .ZN(new_n14107_));
  OAI21_X1   g13813(.A1(new_n7864_), .A2(new_n1332_), .B(new_n14107_), .ZN(new_n14108_));
  AOI21_X1   g13814(.A1(new_n14108_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n14109_));
  XOR2_X1    g13815(.A1(new_n8217_), .A2(new_n14109_), .Z(new_n14110_));
  INV_X1     g13816(.I(new_n14110_), .ZN(new_n14111_));
  NAND3_X1   g13817(.A1(new_n14098_), .A2(new_n14106_), .A3(new_n14111_), .ZN(new_n14112_));
  AOI21_X1   g13818(.A1(new_n14105_), .A2(new_n14101_), .B(new_n14096_), .ZN(new_n14113_));
  NOR3_X1    g13819(.A1(new_n14092_), .A2(new_n14085_), .A3(new_n14097_), .ZN(new_n14114_));
  OAI21_X1   g13820(.A1(new_n14114_), .A2(new_n14113_), .B(new_n14110_), .ZN(new_n14115_));
  AOI21_X1   g13821(.A1(new_n14115_), .A2(new_n14112_), .B(new_n13833_), .ZN(new_n14116_));
  OAI21_X1   g13822(.A1(new_n13706_), .A2(new_n13702_), .B(new_n13717_), .ZN(new_n14117_));
  OAI21_X1   g13823(.A1(new_n14114_), .A2(new_n14113_), .B(new_n14111_), .ZN(new_n14118_));
  NAND3_X1   g13824(.A1(new_n14098_), .A2(new_n14106_), .A3(new_n14110_), .ZN(new_n14119_));
  AOI21_X1   g13825(.A1(new_n14118_), .A2(new_n14119_), .B(new_n14117_), .ZN(new_n14120_));
  NOR2_X1    g13826(.A1(new_n14116_), .A2(new_n14120_), .ZN(new_n14121_));
  NOR3_X1    g13827(.A1(new_n14121_), .A2(new_n13830_), .A3(new_n13832_), .ZN(new_n14122_));
  NAND2_X1   g13828(.A1(new_n14098_), .A2(new_n14106_), .ZN(new_n14123_));
  NOR2_X1    g13829(.A1(new_n13831_), .A2(new_n13714_), .ZN(new_n14125_));
  OAI21_X1   g13830(.A1(new_n14122_), .A2(new_n14125_), .B(new_n13736_), .ZN(new_n14126_));
  NOR3_X1    g13831(.A1(new_n14114_), .A2(new_n14113_), .A3(new_n14110_), .ZN(new_n14127_));
  AOI21_X1   g13832(.A1(new_n14098_), .A2(new_n14106_), .B(new_n14111_), .ZN(new_n14128_));
  OAI21_X1   g13833(.A1(new_n14127_), .A2(new_n14128_), .B(new_n14117_), .ZN(new_n14129_));
  AOI21_X1   g13834(.A1(new_n14098_), .A2(new_n14106_), .B(new_n14110_), .ZN(new_n14130_));
  NOR3_X1    g13835(.A1(new_n14114_), .A2(new_n14113_), .A3(new_n14111_), .ZN(new_n14131_));
  OAI21_X1   g13836(.A1(new_n14131_), .A2(new_n14130_), .B(new_n13833_), .ZN(new_n14132_));
  NAND2_X1   g13837(.A1(new_n14129_), .A2(new_n14132_), .ZN(new_n14133_));
  NAND3_X1   g13838(.A1(new_n14133_), .A2(new_n13722_), .A3(new_n13726_), .ZN(new_n14134_));
  INV_X1     g13839(.I(new_n14125_), .ZN(new_n14135_));
  NAND3_X1   g13840(.A1(new_n14134_), .A2(new_n13417_), .A3(new_n14135_), .ZN(new_n14136_));
  OAI22_X1   g13841(.A1(new_n970_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n820_), .ZN(new_n14137_));
  OAI21_X1   g13842(.A1(new_n8563_), .A2(new_n894_), .B(new_n14137_), .ZN(new_n14138_));
  AOI21_X1   g13843(.A1(new_n14138_), .A2(new_n827_), .B(new_n970_), .ZN(new_n14139_));
  XNOR2_X1   g13844(.A1(new_n9299_), .A2(new_n14139_), .ZN(new_n14140_));
  INV_X1     g13845(.I(new_n14140_), .ZN(new_n14141_));
  NAND3_X1   g13846(.A1(new_n14126_), .A2(new_n14136_), .A3(new_n14141_), .ZN(new_n14142_));
  AOI21_X1   g13847(.A1(new_n14134_), .A2(new_n14135_), .B(new_n13417_), .ZN(new_n14143_));
  NOR3_X1    g13848(.A1(new_n14122_), .A2(new_n13736_), .A3(new_n14125_), .ZN(new_n14144_));
  OAI21_X1   g13849(.A1(new_n14144_), .A2(new_n14143_), .B(new_n14140_), .ZN(new_n14145_));
  OAI22_X1   g13850(.A1(new_n607_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n610_), .ZN(new_n14146_));
  OAI21_X1   g13851(.A1(new_n10025_), .A2(new_n684_), .B(new_n14146_), .ZN(new_n14147_));
  AOI21_X1   g13852(.A1(new_n14147_), .A2(new_n612_), .B(new_n607_), .ZN(new_n14148_));
  XOR2_X1    g13853(.A1(new_n10476_), .A2(new_n14148_), .Z(new_n14149_));
  INV_X1     g13854(.I(new_n14149_), .ZN(new_n14150_));
  NAND3_X1   g13855(.A1(new_n14145_), .A2(new_n14142_), .A3(new_n14150_), .ZN(new_n14151_));
  NOR3_X1    g13856(.A1(new_n14144_), .A2(new_n14143_), .A3(new_n14140_), .ZN(new_n14152_));
  AOI21_X1   g13857(.A1(new_n14126_), .A2(new_n14136_), .B(new_n14141_), .ZN(new_n14153_));
  OAI21_X1   g13858(.A1(new_n14152_), .A2(new_n14153_), .B(new_n14149_), .ZN(new_n14154_));
  AOI22_X1   g13859(.A1(new_n14154_), .A2(new_n14151_), .B1(new_n13827_), .B2(new_n13749_), .ZN(new_n14155_));
  AOI21_X1   g13860(.A1(new_n13738_), .A2(new_n13723_), .B(new_n13733_), .ZN(new_n14156_));
  OAI21_X1   g13861(.A1(new_n13748_), .A2(new_n14156_), .B(new_n13749_), .ZN(new_n14157_));
  OAI21_X1   g13862(.A1(new_n14152_), .A2(new_n14153_), .B(new_n14150_), .ZN(new_n14158_));
  NAND3_X1   g13863(.A1(new_n14145_), .A2(new_n14142_), .A3(new_n14149_), .ZN(new_n14159_));
  AOI21_X1   g13864(.A1(new_n14158_), .A2(new_n14159_), .B(new_n14157_), .ZN(new_n14160_));
  NOR2_X1    g13865(.A1(new_n14160_), .A2(new_n14155_), .ZN(new_n14161_));
  NOR3_X1    g13866(.A1(new_n13825_), .A2(new_n14161_), .A3(new_n13760_), .ZN(new_n14162_));
  AOI21_X1   g13867(.A1(new_n13734_), .A2(new_n13739_), .B(new_n13748_), .ZN(new_n14163_));
  NOR3_X1    g13868(.A1(new_n13724_), .A2(new_n13728_), .A3(new_n13732_), .ZN(new_n14164_));
  NOR2_X1    g13869(.A1(new_n14164_), .A2(new_n14156_), .ZN(new_n14165_));
  NOR2_X1    g13870(.A1(new_n13414_), .A2(new_n14165_), .ZN(new_n14166_));
  NOR2_X1    g13871(.A1(new_n14163_), .A2(new_n14166_), .ZN(new_n14167_));
  NOR2_X1    g13872(.A1(new_n14167_), .A2(new_n13757_), .ZN(new_n14168_));
  OAI21_X1   g13873(.A1(new_n14162_), .A2(new_n14168_), .B(new_n13406_), .ZN(new_n14169_));
  NOR3_X1    g13874(.A1(new_n14152_), .A2(new_n14153_), .A3(new_n14149_), .ZN(new_n14170_));
  AOI21_X1   g13875(.A1(new_n14145_), .A2(new_n14142_), .B(new_n14150_), .ZN(new_n14171_));
  OAI21_X1   g13876(.A1(new_n14170_), .A2(new_n14171_), .B(new_n14157_), .ZN(new_n14172_));
  AOI21_X1   g13877(.A1(new_n13414_), .A2(new_n13750_), .B(new_n14164_), .ZN(new_n14173_));
  AOI21_X1   g13878(.A1(new_n14145_), .A2(new_n14142_), .B(new_n14149_), .ZN(new_n14174_));
  NOR3_X1    g13879(.A1(new_n14152_), .A2(new_n14153_), .A3(new_n14150_), .ZN(new_n14175_));
  OAI21_X1   g13880(.A1(new_n14174_), .A2(new_n14175_), .B(new_n14173_), .ZN(new_n14176_));
  NAND2_X1   g13881(.A1(new_n14176_), .A2(new_n14172_), .ZN(new_n14177_));
  NAND3_X1   g13882(.A1(new_n13763_), .A2(new_n13759_), .A3(new_n14177_), .ZN(new_n14178_));
  INV_X1     g13883(.I(new_n14168_), .ZN(new_n14179_));
  NAND3_X1   g13884(.A1(new_n14178_), .A2(new_n13405_), .A3(new_n14179_), .ZN(new_n14180_));
  OAI22_X1   g13885(.A1(new_n12542_), .A2(new_n341_), .B1(new_n404_), .B2(new_n12970_), .ZN(new_n14181_));
  OAI21_X1   g13886(.A1(new_n12536_), .A2(new_n366_), .B(new_n14181_), .ZN(new_n14182_));
  AOI21_X1   g13887(.A1(new_n14182_), .A2(new_n334_), .B(new_n341_), .ZN(new_n14183_));
  XOR2_X1    g13888(.A1(new_n12969_), .A2(new_n14183_), .Z(new_n14184_));
  OAI22_X1   g13889(.A1(new_n448_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n450_), .ZN(new_n14185_));
  OAI21_X1   g13890(.A1(new_n10862_), .A2(new_n496_), .B(new_n14185_), .ZN(new_n14186_));
  AOI21_X1   g13891(.A1(new_n14186_), .A2(new_n452_), .B(new_n448_), .ZN(new_n14187_));
  XNOR2_X1   g13892(.A1(new_n11748_), .A2(new_n14187_), .ZN(new_n14188_));
  INV_X1     g13893(.I(new_n14188_), .ZN(new_n14189_));
  XOR2_X1    g13894(.A1(new_n14184_), .A2(new_n14189_), .Z(new_n14190_));
  AOI21_X1   g13895(.A1(new_n14169_), .A2(new_n14180_), .B(new_n14190_), .ZN(new_n14191_));
  AOI21_X1   g13896(.A1(new_n14178_), .A2(new_n14179_), .B(new_n13405_), .ZN(new_n14192_));
  NOR3_X1    g13897(.A1(new_n14162_), .A2(new_n13406_), .A3(new_n14168_), .ZN(new_n14193_));
  NOR2_X1    g13898(.A1(new_n14184_), .A2(new_n14188_), .ZN(new_n14194_));
  NAND2_X1   g13899(.A1(new_n14184_), .A2(new_n14188_), .ZN(new_n14195_));
  INV_X1     g13900(.I(new_n14195_), .ZN(new_n14196_));
  NOR2_X1    g13901(.A1(new_n14196_), .A2(new_n14194_), .ZN(new_n14197_));
  NOR3_X1    g13902(.A1(new_n14193_), .A2(new_n14192_), .A3(new_n14197_), .ZN(new_n14198_));
  NOR2_X1    g13903(.A1(\b[60] ), .A2(\b[61] ), .ZN(new_n14199_));
  AOI21_X1   g13904(.A1(new_n13365_), .A2(new_n14199_), .B(new_n12970_), .ZN(new_n14200_));
  NOR2_X1    g13905(.A1(new_n13367_), .A2(new_n13785_), .ZN(new_n14201_));
  INV_X1     g13906(.I(new_n14201_), .ZN(new_n14202_));
  NOR2_X1    g13907(.A1(new_n13365_), .A2(new_n14202_), .ZN(new_n14203_));
  NOR2_X1    g13908(.A1(new_n14200_), .A2(new_n14203_), .ZN(new_n14204_));
  XNOR2_X1   g13909(.A1(\b[61] ), .A2(\b[62] ), .ZN(new_n14205_));
  NOR2_X1    g13910(.A1(new_n14204_), .A2(new_n14205_), .ZN(new_n14206_));
  INV_X1     g13911(.I(new_n14204_), .ZN(new_n14207_));
  INV_X1     g13912(.I(\b[62] ), .ZN(new_n14208_));
  NOR2_X1    g13913(.A1(new_n13785_), .A2(new_n14208_), .ZN(new_n14209_));
  NOR2_X1    g13914(.A1(\b[61] ), .A2(\b[62] ), .ZN(new_n14210_));
  NOR2_X1    g13915(.A1(new_n14209_), .A2(new_n14210_), .ZN(new_n14211_));
  NOR2_X1    g13916(.A1(new_n14207_), .A2(new_n14211_), .ZN(new_n14212_));
  NOR2_X1    g13917(.A1(new_n14212_), .A2(new_n14206_), .ZN(new_n14213_));
  OAI22_X1   g13918(.A1(new_n330_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n263_), .ZN(new_n14214_));
  OAI21_X1   g13919(.A1(new_n13367_), .A2(new_n289_), .B(new_n14214_), .ZN(new_n14215_));
  AOI21_X1   g13920(.A1(new_n14215_), .A2(new_n260_), .B(new_n426_), .ZN(new_n14216_));
  XOR2_X1    g13921(.A1(new_n14213_), .A2(new_n14216_), .Z(new_n14217_));
  NOR3_X1    g13922(.A1(new_n14198_), .A2(new_n14191_), .A3(new_n14217_), .ZN(new_n14218_));
  INV_X1     g13923(.I(new_n14190_), .ZN(new_n14219_));
  OAI21_X1   g13924(.A1(new_n14193_), .A2(new_n14192_), .B(new_n14219_), .ZN(new_n14220_));
  INV_X1     g13925(.I(new_n14197_), .ZN(new_n14221_));
  NAND3_X1   g13926(.A1(new_n14169_), .A2(new_n14180_), .A3(new_n14221_), .ZN(new_n14222_));
  INV_X1     g13927(.I(new_n14217_), .ZN(new_n14223_));
  AOI21_X1   g13928(.A1(new_n14220_), .A2(new_n14222_), .B(new_n14223_), .ZN(new_n14224_));
  OAI21_X1   g13929(.A1(new_n14218_), .A2(new_n14224_), .B(new_n13824_), .ZN(new_n14225_));
  INV_X1     g13930(.I(new_n13824_), .ZN(new_n14226_));
  OAI21_X1   g13931(.A1(new_n14198_), .A2(new_n14191_), .B(new_n14223_), .ZN(new_n14227_));
  NAND3_X1   g13932(.A1(new_n14220_), .A2(new_n14222_), .A3(new_n14217_), .ZN(new_n14228_));
  NAND2_X1   g13933(.A1(new_n14227_), .A2(new_n14228_), .ZN(new_n14229_));
  NAND2_X1   g13934(.A1(new_n14226_), .A2(new_n14229_), .ZN(new_n14230_));
  NAND2_X1   g13935(.A1(new_n14230_), .A2(new_n14225_), .ZN(new_n14231_));
  NAND2_X1   g13936(.A1(new_n13822_), .A2(new_n14231_), .ZN(new_n14232_));
  AND2_X2    g13937(.A1(new_n14230_), .A2(new_n14225_), .Z(new_n14233_));
  NAND2_X1   g13938(.A1(new_n14233_), .A2(new_n13821_), .ZN(new_n14234_));
  NAND2_X1   g13939(.A1(new_n14232_), .A2(new_n14234_), .ZN(new_n14235_));
  XNOR2_X1   g13940(.A1(new_n13821_), .A2(new_n14231_), .ZN(new_n14236_));
  MUX2_X1    g13941(.I0(new_n14236_), .I1(new_n14235_), .S(new_n13820_), .Z(\f[62] ));
  OAI22_X1   g13942(.A1(new_n12970_), .A2(new_n341_), .B1(new_n404_), .B2(new_n13367_), .ZN(new_n14238_));
  OAI21_X1   g13943(.A1(new_n12542_), .A2(new_n366_), .B(new_n14238_), .ZN(new_n14239_));
  AOI21_X1   g13944(.A1(new_n14239_), .A2(new_n334_), .B(new_n341_), .ZN(new_n14240_));
  XNOR2_X1   g13945(.A1(new_n13371_), .A2(new_n14240_), .ZN(new_n14241_));
  INV_X1     g13946(.I(new_n14194_), .ZN(new_n14242_));
  NAND3_X1   g13947(.A1(new_n14169_), .A2(new_n14180_), .A3(new_n14195_), .ZN(new_n14243_));
  NAND2_X1   g13948(.A1(new_n14243_), .A2(new_n14242_), .ZN(new_n14244_));
  NOR2_X1    g13949(.A1(new_n14152_), .A2(new_n14153_), .ZN(new_n14245_));
  XOR2_X1    g13950(.A1(new_n14123_), .A2(new_n14117_), .Z(new_n14246_));
  NAND2_X1   g13951(.A1(new_n14246_), .A2(new_n14110_), .ZN(new_n14247_));
  INV_X1     g13952(.I(new_n14247_), .ZN(new_n14248_));
  OAI21_X1   g13953(.A1(new_n14121_), .A2(new_n13714_), .B(new_n13831_), .ZN(new_n14249_));
  INV_X1     g13954(.I(new_n14249_), .ZN(new_n14250_));
  OAI21_X1   g13955(.A1(new_n14133_), .A2(new_n13715_), .B(new_n13417_), .ZN(new_n14251_));
  OAI21_X1   g13956(.A1(new_n13833_), .A2(new_n14114_), .B(new_n14098_), .ZN(new_n14252_));
  OAI21_X1   g13957(.A1(new_n14072_), .A2(new_n14073_), .B(new_n13656_), .ZN(new_n14253_));
  AOI21_X1   g13958(.A1(new_n14253_), .A2(new_n14071_), .B(new_n13657_), .ZN(new_n14254_));
  NAND2_X1   g13959(.A1(new_n13846_), .A2(new_n13844_), .ZN(new_n14255_));
  NAND2_X1   g13960(.A1(new_n14025_), .A2(new_n14018_), .ZN(new_n14256_));
  XOR2_X1    g13961(.A1(new_n14256_), .A2(new_n13842_), .Z(new_n14257_));
  NOR2_X1    g13962(.A1(new_n14255_), .A2(new_n14257_), .ZN(new_n14258_));
  NAND2_X1   g13963(.A1(new_n14256_), .A2(new_n13841_), .ZN(new_n14259_));
  OAI21_X1   g13964(.A1(new_n14022_), .A2(new_n14023_), .B(new_n14021_), .ZN(new_n14260_));
  AOI21_X1   g13965(.A1(new_n14260_), .A2(new_n13616_), .B(new_n13619_), .ZN(new_n14261_));
  INV_X1     g13966(.I(new_n14261_), .ZN(new_n14262_));
  OAI21_X1   g13967(.A1(new_n14004_), .A2(new_n14005_), .B(new_n14003_), .ZN(new_n14263_));
  NAND2_X1   g13968(.A1(new_n14263_), .A2(new_n13596_), .ZN(new_n14264_));
  NOR2_X1    g13969(.A1(new_n13974_), .A2(new_n13975_), .ZN(new_n14265_));
  XOR2_X1    g13970(.A1(new_n13987_), .A2(new_n14265_), .Z(new_n14266_));
  NAND2_X1   g13971(.A1(new_n13985_), .A2(new_n13853_), .ZN(new_n14267_));
  AOI21_X1   g13972(.A1(new_n13864_), .A2(new_n13862_), .B(new_n13975_), .ZN(new_n14268_));
  XOR2_X1    g13973(.A1(new_n13868_), .A2(new_n13950_), .Z(new_n14269_));
  NAND2_X1   g13974(.A1(new_n14269_), .A2(new_n13943_), .ZN(new_n14270_));
  AOI21_X1   g13975(.A1(new_n13913_), .A2(new_n13908_), .B(new_n13921_), .ZN(new_n14271_));
  INV_X1     g13976(.I(new_n14271_), .ZN(new_n14272_));
  INV_X1     g13977(.I(new_n13912_), .ZN(new_n14273_));
  OAI21_X1   g13978(.A1(new_n13875_), .A2(new_n13874_), .B(new_n14273_), .ZN(new_n14274_));
  AOI21_X1   g13979(.A1(new_n13897_), .A2(new_n13895_), .B(new_n13893_), .ZN(new_n14275_));
  NAND2_X1   g13980(.A1(new_n13888_), .A2(new_n13878_), .ZN(new_n14276_));
  OAI22_X1   g13981(.A1(new_n13880_), .A2(new_n10569_), .B1(new_n269_), .B2(new_n13885_), .ZN(new_n14277_));
  AOI21_X1   g13982(.A1(new_n14277_), .A2(new_n13476_), .B(new_n403_), .ZN(new_n14278_));
  XOR2_X1    g13983(.A1(new_n14278_), .A2(new_n13466_), .Z(new_n14279_));
  INV_X1     g13984(.I(\a[63] ), .ZN(new_n14280_));
  NOR2_X1    g13985(.A1(new_n14280_), .A2(\a[62] ), .ZN(new_n14281_));
  NOR2_X1    g13986(.A1(new_n13476_), .A2(\a[63] ), .ZN(new_n14282_));
  OAI21_X1   g13987(.A1(new_n14281_), .A2(new_n14282_), .B(\b[0] ), .ZN(new_n14283_));
  INV_X1     g13988(.I(new_n14283_), .ZN(new_n14284_));
  XOR2_X1    g13989(.A1(new_n14279_), .A2(new_n14284_), .Z(new_n14285_));
  NOR2_X1    g13990(.A1(new_n14285_), .A2(new_n14276_), .ZN(new_n14286_));
  OR2_X2     g13991(.A1(new_n14279_), .A2(new_n14283_), .Z(new_n14287_));
  NAND2_X1   g13992(.A1(new_n14279_), .A2(new_n14283_), .ZN(new_n14288_));
  NAND2_X1   g13993(.A1(new_n14287_), .A2(new_n14288_), .ZN(new_n14289_));
  AOI21_X1   g13994(.A1(new_n14276_), .A2(new_n14289_), .B(new_n14286_), .ZN(new_n14290_));
  OAI22_X1   g13995(.A1(new_n12226_), .A2(new_n421_), .B1(new_n12637_), .B2(new_n325_), .ZN(new_n14291_));
  AOI21_X1   g13996(.A1(new_n14291_), .A2(new_n12222_), .B(new_n12643_), .ZN(new_n14292_));
  XOR2_X1    g13997(.A1(new_n425_), .A2(new_n14292_), .Z(new_n14293_));
  INV_X1     g13998(.I(new_n14293_), .ZN(new_n14294_));
  NAND2_X1   g13999(.A1(new_n14290_), .A2(new_n14294_), .ZN(new_n14295_));
  NAND2_X1   g14000(.A1(new_n14289_), .A2(new_n14276_), .ZN(new_n14296_));
  OAI21_X1   g14001(.A1(new_n14276_), .A2(new_n14285_), .B(new_n14296_), .ZN(new_n14297_));
  NAND2_X1   g14002(.A1(new_n14297_), .A2(new_n14293_), .ZN(new_n14298_));
  AOI21_X1   g14003(.A1(new_n14295_), .A2(new_n14298_), .B(new_n14275_), .ZN(new_n14299_));
  INV_X1     g14004(.I(new_n14275_), .ZN(new_n14300_));
  NOR2_X1    g14005(.A1(new_n14290_), .A2(new_n14293_), .ZN(new_n14301_));
  NOR2_X1    g14006(.A1(new_n14297_), .A2(new_n14294_), .ZN(new_n14302_));
  NOR2_X1    g14007(.A1(new_n14302_), .A2(new_n14301_), .ZN(new_n14303_));
  NOR2_X1    g14008(.A1(new_n14300_), .A2(new_n14303_), .ZN(new_n14304_));
  AOI22_X1   g14009(.A1(new_n10969_), .A2(new_n650_), .B1(new_n11394_), .B2(\b[7] ), .ZN(new_n14305_));
  OAI21_X1   g14010(.A1(new_n14305_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n14306_));
  XOR2_X1    g14011(.A1(new_n569_), .A2(new_n14306_), .Z(new_n14307_));
  NOR3_X1    g14012(.A1(new_n14304_), .A2(new_n14299_), .A3(new_n14307_), .ZN(new_n14308_));
  NAND2_X1   g14013(.A1(new_n14298_), .A2(new_n14295_), .ZN(new_n14309_));
  NAND2_X1   g14014(.A1(new_n14300_), .A2(new_n14309_), .ZN(new_n14310_));
  OAI21_X1   g14015(.A1(new_n14301_), .A2(new_n14302_), .B(new_n14275_), .ZN(new_n14311_));
  INV_X1     g14016(.I(new_n14307_), .ZN(new_n14312_));
  AOI21_X1   g14017(.A1(new_n14310_), .A2(new_n14311_), .B(new_n14312_), .ZN(new_n14313_));
  NOR2_X1    g14018(.A1(new_n14308_), .A2(new_n14313_), .ZN(new_n14314_));
  AOI21_X1   g14019(.A1(new_n13910_), .A2(new_n14274_), .B(new_n14314_), .ZN(new_n14315_));
  NAND2_X1   g14020(.A1(new_n14274_), .A2(new_n13910_), .ZN(new_n14316_));
  OAI21_X1   g14021(.A1(new_n14304_), .A2(new_n14299_), .B(new_n14312_), .ZN(new_n14317_));
  NAND3_X1   g14022(.A1(new_n14310_), .A2(new_n14311_), .A3(new_n14307_), .ZN(new_n14318_));
  AOI21_X1   g14023(.A1(new_n14317_), .A2(new_n14318_), .B(new_n14316_), .ZN(new_n14319_));
  INV_X1     g14024(.I(new_n781_), .ZN(new_n14320_));
  AOI22_X1   g14025(.A1(new_n11415_), .A2(new_n14320_), .B1(\b[10] ), .B2(new_n10145_), .ZN(new_n14321_));
  OAI21_X1   g14026(.A1(new_n14321_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n14322_));
  XNOR2_X1   g14027(.A1(new_n785_), .A2(new_n14322_), .ZN(new_n14323_));
  INV_X1     g14028(.I(new_n14323_), .ZN(new_n14324_));
  OAI21_X1   g14029(.A1(new_n14319_), .A2(new_n14315_), .B(new_n14324_), .ZN(new_n14325_));
  AOI21_X1   g14030(.A1(new_n13873_), .A2(new_n13929_), .B(new_n14325_), .ZN(new_n14326_));
  OAI21_X1   g14031(.A1(new_n14308_), .A2(new_n14313_), .B(new_n14316_), .ZN(new_n14327_));
  NAND2_X1   g14032(.A1(new_n14317_), .A2(new_n14318_), .ZN(new_n14328_));
  NAND3_X1   g14033(.A1(new_n14328_), .A2(new_n13910_), .A3(new_n14274_), .ZN(new_n14329_));
  AOI21_X1   g14034(.A1(new_n14327_), .A2(new_n14329_), .B(new_n14323_), .ZN(new_n14330_));
  NOR3_X1    g14035(.A1(new_n14330_), .A2(new_n13923_), .A3(new_n13926_), .ZN(new_n14331_));
  OAI21_X1   g14036(.A1(new_n14326_), .A2(new_n14331_), .B(new_n14272_), .ZN(new_n14332_));
  OAI21_X1   g14037(.A1(new_n13926_), .A2(new_n13923_), .B(new_n14330_), .ZN(new_n14333_));
  NAND3_X1   g14038(.A1(new_n14325_), .A2(new_n13929_), .A3(new_n13873_), .ZN(new_n14334_));
  NAND3_X1   g14039(.A1(new_n14333_), .A2(new_n14334_), .A3(new_n14271_), .ZN(new_n14335_));
  AOI22_X1   g14040(.A1(new_n8631_), .A2(\b[14] ), .B1(\b[15] ), .B2(new_n9382_), .ZN(new_n14336_));
  AOI21_X1   g14041(.A1(\b[13] ), .A2(new_n9731_), .B(new_n14336_), .ZN(new_n14337_));
  OAI21_X1   g14042(.A1(new_n14337_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n14338_));
  XNOR2_X1   g14043(.A1(new_n1024_), .A2(new_n14338_), .ZN(new_n14339_));
  AOI21_X1   g14044(.A1(new_n14332_), .A2(new_n14335_), .B(new_n14339_), .ZN(new_n14340_));
  OAI21_X1   g14045(.A1(new_n13868_), .A2(new_n13950_), .B(new_n14340_), .ZN(new_n14341_));
  NOR2_X1    g14046(.A1(new_n13868_), .A2(new_n13950_), .ZN(new_n14342_));
  AOI21_X1   g14047(.A1(new_n14333_), .A2(new_n14334_), .B(new_n14271_), .ZN(new_n14343_));
  NOR3_X1    g14048(.A1(new_n14326_), .A2(new_n14272_), .A3(new_n14331_), .ZN(new_n14344_));
  INV_X1     g14049(.I(new_n14339_), .ZN(new_n14345_));
  OAI21_X1   g14050(.A1(new_n14344_), .A2(new_n14343_), .B(new_n14345_), .ZN(new_n14346_));
  NAND2_X1   g14051(.A1(new_n14342_), .A2(new_n14346_), .ZN(new_n14347_));
  AOI21_X1   g14052(.A1(new_n14341_), .A2(new_n14347_), .B(new_n13939_), .ZN(new_n14348_));
  NOR2_X1    g14053(.A1(new_n14342_), .A2(new_n14346_), .ZN(new_n14349_));
  NOR3_X1    g14054(.A1(new_n14340_), .A2(new_n13868_), .A3(new_n13950_), .ZN(new_n14350_));
  NOR3_X1    g14055(.A1(new_n14349_), .A2(new_n14350_), .A3(new_n13947_), .ZN(new_n14351_));
  OAI22_X1   g14056(.A1(new_n7619_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n8309_), .ZN(new_n14352_));
  OAI21_X1   g14057(.A1(new_n1109_), .A2(new_n7947_), .B(new_n14352_), .ZN(new_n14353_));
  AOI21_X1   g14058(.A1(new_n14353_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n14354_));
  XOR2_X1    g14059(.A1(new_n1299_), .A2(new_n14354_), .Z(new_n14355_));
  INV_X1     g14060(.I(new_n14355_), .ZN(new_n14356_));
  OAI21_X1   g14061(.A1(new_n14348_), .A2(new_n14351_), .B(new_n14356_), .ZN(new_n14357_));
  NOR2_X1    g14062(.A1(new_n14357_), .A2(new_n13958_), .ZN(new_n14358_));
  OAI21_X1   g14063(.A1(new_n14349_), .A2(new_n14350_), .B(new_n13947_), .ZN(new_n14359_));
  NAND3_X1   g14064(.A1(new_n14341_), .A2(new_n14347_), .A3(new_n13939_), .ZN(new_n14360_));
  AOI21_X1   g14065(.A1(new_n14360_), .A2(new_n14359_), .B(new_n14355_), .ZN(new_n14361_));
  NOR2_X1    g14066(.A1(new_n13966_), .A2(new_n14361_), .ZN(new_n14362_));
  OAI21_X1   g14067(.A1(new_n14362_), .A2(new_n14358_), .B(new_n14270_), .ZN(new_n14363_));
  INV_X1     g14068(.I(new_n14270_), .ZN(new_n14364_));
  NAND2_X1   g14069(.A1(new_n13966_), .A2(new_n14361_), .ZN(new_n14365_));
  NAND2_X1   g14070(.A1(new_n14357_), .A2(new_n13958_), .ZN(new_n14366_));
  NAND3_X1   g14071(.A1(new_n14365_), .A2(new_n14366_), .A3(new_n14364_), .ZN(new_n14367_));
  OAI22_X1   g14072(.A1(new_n6644_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n6647_), .ZN(new_n14368_));
  OAI21_X1   g14073(.A1(new_n1518_), .A2(new_n7284_), .B(new_n14368_), .ZN(new_n14369_));
  AOI21_X1   g14074(.A1(new_n14369_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n14370_));
  XNOR2_X1   g14075(.A1(new_n1638_), .A2(new_n14370_), .ZN(new_n14371_));
  AOI21_X1   g14076(.A1(new_n14363_), .A2(new_n14367_), .B(new_n14371_), .ZN(new_n14372_));
  AOI21_X1   g14077(.A1(new_n14365_), .A2(new_n14366_), .B(new_n14364_), .ZN(new_n14373_));
  NOR3_X1    g14078(.A1(new_n14362_), .A2(new_n14358_), .A3(new_n14270_), .ZN(new_n14374_));
  INV_X1     g14079(.I(new_n14371_), .ZN(new_n14375_));
  NOR3_X1    g14080(.A1(new_n14373_), .A2(new_n14374_), .A3(new_n14375_), .ZN(new_n14376_));
  OAI22_X1   g14081(.A1(new_n14376_), .A2(new_n14372_), .B1(new_n14268_), .B2(new_n13974_), .ZN(new_n14377_));
  NOR2_X1    g14082(.A1(new_n14268_), .A2(new_n13974_), .ZN(new_n14378_));
  NOR3_X1    g14083(.A1(new_n14373_), .A2(new_n14374_), .A3(new_n14371_), .ZN(new_n14379_));
  AOI21_X1   g14084(.A1(new_n14363_), .A2(new_n14367_), .B(new_n14375_), .ZN(new_n14380_));
  OAI21_X1   g14085(.A1(new_n14379_), .A2(new_n14380_), .B(new_n14378_), .ZN(new_n14381_));
  OAI22_X1   g14086(.A1(new_n5993_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n5991_), .ZN(new_n14382_));
  OAI21_X1   g14087(.A1(new_n1803_), .A2(new_n5997_), .B(new_n14382_), .ZN(new_n14383_));
  AOI21_X1   g14088(.A1(new_n14383_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n14384_));
  XOR2_X1    g14089(.A1(new_n2106_), .A2(new_n14384_), .Z(new_n14385_));
  AOI21_X1   g14090(.A1(new_n14381_), .A2(new_n14377_), .B(new_n14385_), .ZN(new_n14386_));
  OAI21_X1   g14091(.A1(new_n14267_), .A2(new_n13988_), .B(new_n14386_), .ZN(new_n14387_));
  NOR2_X1    g14092(.A1(new_n14267_), .A2(new_n13988_), .ZN(new_n14388_));
  INV_X1     g14093(.I(new_n14377_), .ZN(new_n14389_));
  INV_X1     g14094(.I(new_n14268_), .ZN(new_n14390_));
  NAND2_X1   g14095(.A1(new_n14390_), .A2(new_n13964_), .ZN(new_n14391_));
  NOR2_X1    g14096(.A1(new_n14379_), .A2(new_n14380_), .ZN(new_n14392_));
  NOR2_X1    g14097(.A1(new_n14391_), .A2(new_n14392_), .ZN(new_n14393_));
  INV_X1     g14098(.I(new_n14385_), .ZN(new_n14394_));
  OAI21_X1   g14099(.A1(new_n14393_), .A2(new_n14389_), .B(new_n14394_), .ZN(new_n14395_));
  NAND2_X1   g14100(.A1(new_n14388_), .A2(new_n14395_), .ZN(new_n14396_));
  AOI22_X1   g14101(.A1(new_n14396_), .A2(new_n14387_), .B1(new_n13971_), .B2(new_n14266_), .ZN(new_n14397_));
  NAND2_X1   g14102(.A1(new_n14266_), .A2(new_n13971_), .ZN(new_n14398_));
  NOR2_X1    g14103(.A1(new_n14388_), .A2(new_n14395_), .ZN(new_n14399_));
  NOR3_X1    g14104(.A1(new_n14386_), .A2(new_n14267_), .A3(new_n13988_), .ZN(new_n14400_));
  NOR3_X1    g14105(.A1(new_n14399_), .A2(new_n14400_), .A3(new_n14398_), .ZN(new_n14401_));
  OAI22_X1   g14106(.A1(new_n5420_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n5107_), .ZN(new_n14402_));
  OAI21_X1   g14107(.A1(new_n2281_), .A2(new_n5112_), .B(new_n14402_), .ZN(new_n14403_));
  AOI21_X1   g14108(.A1(new_n14403_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n14404_));
  XNOR2_X1   g14109(.A1(new_n2647_), .A2(new_n14404_), .ZN(new_n14405_));
  INV_X1     g14110(.I(new_n14405_), .ZN(new_n14406_));
  OAI21_X1   g14111(.A1(new_n14397_), .A2(new_n14401_), .B(new_n14406_), .ZN(new_n14407_));
  AOI21_X1   g14112(.A1(new_n13595_), .A2(new_n14264_), .B(new_n14407_), .ZN(new_n14408_));
  NAND2_X1   g14113(.A1(new_n14264_), .A2(new_n13595_), .ZN(new_n14409_));
  OAI21_X1   g14114(.A1(new_n14399_), .A2(new_n14400_), .B(new_n14398_), .ZN(new_n14410_));
  NAND4_X1   g14115(.A1(new_n14396_), .A2(new_n13971_), .A3(new_n14266_), .A4(new_n14387_), .ZN(new_n14411_));
  AOI21_X1   g14116(.A1(new_n14411_), .A2(new_n14410_), .B(new_n14405_), .ZN(new_n14412_));
  NOR2_X1    g14117(.A1(new_n14409_), .A2(new_n14412_), .ZN(new_n14413_));
  OAI21_X1   g14118(.A1(new_n14408_), .A2(new_n14413_), .B(new_n13998_), .ZN(new_n14414_));
  NAND2_X1   g14119(.A1(new_n14409_), .A2(new_n14412_), .ZN(new_n14415_));
  NAND3_X1   g14120(.A1(new_n14407_), .A2(new_n13595_), .A3(new_n14264_), .ZN(new_n14416_));
  NAND3_X1   g14121(.A1(new_n14415_), .A2(new_n14416_), .A3(new_n14005_), .ZN(new_n14417_));
  OAI22_X1   g14122(.A1(new_n4072_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n4067_), .ZN(new_n14418_));
  OAI21_X1   g14123(.A1(new_n2842_), .A2(new_n4318_), .B(new_n14418_), .ZN(new_n14419_));
  AOI21_X1   g14124(.A1(new_n14419_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n14420_));
  XNOR2_X1   g14125(.A1(new_n3264_), .A2(new_n14420_), .ZN(new_n14421_));
  AOI21_X1   g14126(.A1(new_n14414_), .A2(new_n14417_), .B(new_n14421_), .ZN(new_n14422_));
  NAND2_X1   g14127(.A1(new_n14262_), .A2(new_n14422_), .ZN(new_n14423_));
  AOI21_X1   g14128(.A1(new_n14415_), .A2(new_n14416_), .B(new_n14005_), .ZN(new_n14424_));
  NOR3_X1    g14129(.A1(new_n14408_), .A2(new_n14413_), .A3(new_n13998_), .ZN(new_n14425_));
  INV_X1     g14130(.I(new_n14421_), .ZN(new_n14426_));
  OAI21_X1   g14131(.A1(new_n14425_), .A2(new_n14424_), .B(new_n14426_), .ZN(new_n14427_));
  NAND2_X1   g14132(.A1(new_n14427_), .A2(new_n14261_), .ZN(new_n14428_));
  AOI21_X1   g14133(.A1(new_n14423_), .A2(new_n14428_), .B(new_n14023_), .ZN(new_n14429_));
  NOR2_X1    g14134(.A1(new_n14427_), .A2(new_n14261_), .ZN(new_n14430_));
  NOR2_X1    g14135(.A1(new_n14262_), .A2(new_n14422_), .ZN(new_n14431_));
  NOR3_X1    g14136(.A1(new_n14431_), .A2(new_n14430_), .A3(new_n14016_), .ZN(new_n14432_));
  NOR2_X1    g14137(.A1(new_n14432_), .A2(new_n14429_), .ZN(new_n14433_));
  OAI22_X1   g14138(.A1(new_n3717_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n3989_), .ZN(new_n14434_));
  OAI21_X1   g14139(.A1(new_n3709_), .A2(new_n3569_), .B(new_n14434_), .ZN(new_n14435_));
  AOI21_X1   g14140(.A1(new_n14435_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n14436_));
  XNOR2_X1   g14141(.A1(new_n3993_), .A2(new_n14436_), .ZN(new_n14437_));
  INV_X1     g14142(.I(new_n14437_), .ZN(new_n14438_));
  NAND2_X1   g14143(.A1(new_n14433_), .A2(new_n14438_), .ZN(new_n14439_));
  OAI21_X1   g14144(.A1(new_n14431_), .A2(new_n14430_), .B(new_n14016_), .ZN(new_n14440_));
  NAND3_X1   g14145(.A1(new_n14423_), .A2(new_n14428_), .A3(new_n14023_), .ZN(new_n14441_));
  NAND2_X1   g14146(.A1(new_n14440_), .A2(new_n14441_), .ZN(new_n14442_));
  NAND2_X1   g14147(.A1(new_n14442_), .A2(new_n14437_), .ZN(new_n14443_));
  NAND2_X1   g14148(.A1(new_n14439_), .A2(new_n14443_), .ZN(new_n14444_));
  OAI22_X1   g14149(.A1(new_n4500_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n4774_), .ZN(new_n14445_));
  OAI21_X1   g14150(.A1(new_n4253_), .A2(new_n2884_), .B(new_n14445_), .ZN(new_n14446_));
  AOI21_X1   g14151(.A1(new_n14446_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n14447_));
  XNOR2_X1   g14152(.A1(new_n4778_), .A2(new_n14447_), .ZN(new_n14448_));
  INV_X1     g14153(.I(new_n14448_), .ZN(new_n14449_));
  NAND3_X1   g14154(.A1(new_n14444_), .A2(new_n14259_), .A3(new_n14449_), .ZN(new_n14450_));
  INV_X1     g14155(.I(new_n14259_), .ZN(new_n14451_));
  NOR2_X1    g14156(.A1(new_n14442_), .A2(new_n14437_), .ZN(new_n14452_));
  NOR2_X1    g14157(.A1(new_n14433_), .A2(new_n14438_), .ZN(new_n14453_));
  OAI21_X1   g14158(.A1(new_n14453_), .A2(new_n14452_), .B(new_n14449_), .ZN(new_n14454_));
  NAND2_X1   g14159(.A1(new_n14454_), .A2(new_n14451_), .ZN(new_n14455_));
  AOI21_X1   g14160(.A1(new_n14455_), .A2(new_n14450_), .B(new_n14258_), .ZN(new_n14456_));
  INV_X1     g14161(.I(new_n14258_), .ZN(new_n14457_));
  NOR2_X1    g14162(.A1(new_n14454_), .A2(new_n14451_), .ZN(new_n14458_));
  AOI21_X1   g14163(.A1(new_n14444_), .A2(new_n14449_), .B(new_n14259_), .ZN(new_n14459_));
  NOR3_X1    g14164(.A1(new_n14458_), .A2(new_n14459_), .A3(new_n14457_), .ZN(new_n14460_));
  NOR2_X1    g14165(.A1(new_n14460_), .A2(new_n14456_), .ZN(new_n14461_));
  AOI21_X1   g14166(.A1(new_n14056_), .A2(new_n13632_), .B(new_n13643_), .ZN(new_n14462_));
  NAND2_X1   g14167(.A1(new_n14049_), .A2(new_n13631_), .ZN(new_n14463_));
  NAND2_X1   g14168(.A1(new_n14463_), .A2(new_n13433_), .ZN(new_n14464_));
  NOR2_X1    g14169(.A1(new_n14464_), .A2(new_n14462_), .ZN(new_n14465_));
  INV_X1     g14170(.I(new_n14465_), .ZN(new_n14466_));
  XNOR2_X1   g14171(.A1(new_n14255_), .A2(new_n14256_), .ZN(new_n14467_));
  NOR2_X1    g14172(.A1(new_n14467_), .A2(new_n13842_), .ZN(new_n14468_));
  XOR2_X1    g14173(.A1(new_n14255_), .A2(new_n14256_), .Z(new_n14469_));
  NOR2_X1    g14174(.A1(new_n14469_), .A2(new_n13841_), .ZN(new_n14470_));
  OAI21_X1   g14175(.A1(new_n14468_), .A2(new_n14470_), .B(new_n14030_), .ZN(new_n14471_));
  NAND2_X1   g14176(.A1(new_n14466_), .A2(new_n14471_), .ZN(new_n14472_));
  INV_X1     g14177(.I(new_n14471_), .ZN(new_n14473_));
  NOR2_X1    g14178(.A1(new_n14461_), .A2(new_n14473_), .ZN(new_n14474_));
  AOI22_X1   g14179(.A1(new_n14472_), .A2(new_n14461_), .B1(new_n14474_), .B2(new_n14466_), .ZN(new_n14475_));
  OAI22_X1   g14180(.A1(new_n2171_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n2166_), .ZN(new_n14476_));
  OAI21_X1   g14181(.A1(new_n5068_), .A2(new_n2322_), .B(new_n14476_), .ZN(new_n14477_));
  AOI21_X1   g14182(.A1(new_n14477_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n14478_));
  XNOR2_X1   g14183(.A1(new_n5600_), .A2(new_n14478_), .ZN(new_n14479_));
  NOR3_X1    g14184(.A1(new_n14254_), .A2(new_n14475_), .A3(new_n14479_), .ZN(new_n14480_));
  AOI21_X1   g14185(.A1(new_n14068_), .A2(new_n14065_), .B(new_n13677_), .ZN(new_n14481_));
  OAI21_X1   g14186(.A1(new_n14481_), .A2(new_n13662_), .B(new_n13678_), .ZN(new_n14482_));
  OAI21_X1   g14187(.A1(new_n14465_), .A2(new_n14473_), .B(new_n14461_), .ZN(new_n14483_));
  OAI21_X1   g14188(.A1(new_n14458_), .A2(new_n14459_), .B(new_n14457_), .ZN(new_n14484_));
  NAND3_X1   g14189(.A1(new_n14455_), .A2(new_n14450_), .A3(new_n14258_), .ZN(new_n14485_));
  NAND2_X1   g14190(.A1(new_n14484_), .A2(new_n14485_), .ZN(new_n14486_));
  NAND3_X1   g14191(.A1(new_n14466_), .A2(new_n14486_), .A3(new_n14471_), .ZN(new_n14487_));
  AOI21_X1   g14192(.A1(new_n14487_), .A2(new_n14483_), .B(new_n14479_), .ZN(new_n14488_));
  NOR2_X1    g14193(.A1(new_n14482_), .A2(new_n14488_), .ZN(new_n14489_));
  OAI21_X1   g14194(.A1(new_n14480_), .A2(new_n14489_), .B(new_n14068_), .ZN(new_n14490_));
  NAND2_X1   g14195(.A1(new_n14482_), .A2(new_n14488_), .ZN(new_n14491_));
  OAI21_X1   g14196(.A1(new_n14475_), .A2(new_n14479_), .B(new_n14254_), .ZN(new_n14492_));
  NAND3_X1   g14197(.A1(new_n14492_), .A2(new_n14073_), .A3(new_n14491_), .ZN(new_n14493_));
  NAND2_X1   g14198(.A1(new_n14493_), .A2(new_n14490_), .ZN(new_n14494_));
  AOI22_X1   g14199(.A1(\b[42] ), .A2(new_n2725_), .B1(new_n1702_), .B2(\b[41] ), .ZN(new_n14495_));
  AOI21_X1   g14200(.A1(\b[40] ), .A2(new_n1851_), .B(new_n14495_), .ZN(new_n14496_));
  OAI21_X1   g14201(.A1(new_n14496_), .A2(\a[23] ), .B(new_n1702_), .ZN(new_n14497_));
  XOR2_X1    g14202(.A1(new_n6543_), .A2(new_n14497_), .Z(new_n14498_));
  NAND3_X1   g14203(.A1(new_n14494_), .A2(new_n14084_), .A3(new_n14498_), .ZN(new_n14499_));
  AOI21_X1   g14204(.A1(new_n14492_), .A2(new_n14491_), .B(new_n14073_), .ZN(new_n14500_));
  NOR3_X1    g14205(.A1(new_n14480_), .A2(new_n14489_), .A3(new_n14068_), .ZN(new_n14501_));
  OAI21_X1   g14206(.A1(new_n14500_), .A2(new_n14501_), .B(new_n14498_), .ZN(new_n14502_));
  NAND2_X1   g14207(.A1(new_n14502_), .A2(new_n14100_), .ZN(new_n14503_));
  AOI21_X1   g14208(.A1(new_n14503_), .A2(new_n14499_), .B(new_n14092_), .ZN(new_n14504_));
  NOR2_X1    g14209(.A1(new_n14502_), .A2(new_n14100_), .ZN(new_n14505_));
  AOI21_X1   g14210(.A1(new_n14494_), .A2(new_n14498_), .B(new_n14084_), .ZN(new_n14506_));
  NOR3_X1    g14211(.A1(new_n14505_), .A2(new_n14506_), .A3(new_n14105_), .ZN(new_n14507_));
  OAI22_X1   g14212(.A1(new_n1347_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n1344_), .ZN(new_n14508_));
  OAI21_X1   g14213(.A1(new_n6847_), .A2(new_n1457_), .B(new_n14508_), .ZN(new_n14509_));
  AOI21_X1   g14214(.A1(new_n14509_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n14510_));
  XOR2_X1    g14215(.A1(new_n7516_), .A2(new_n14510_), .Z(new_n14511_));
  INV_X1     g14216(.I(new_n14511_), .ZN(new_n14512_));
  OAI21_X1   g14217(.A1(new_n14507_), .A2(new_n14504_), .B(new_n14512_), .ZN(new_n14513_));
  OAI21_X1   g14218(.A1(new_n14505_), .A2(new_n14506_), .B(new_n14105_), .ZN(new_n14514_));
  NAND3_X1   g14219(.A1(new_n14503_), .A2(new_n14499_), .A3(new_n14092_), .ZN(new_n14515_));
  NAND3_X1   g14220(.A1(new_n14514_), .A2(new_n14515_), .A3(new_n14511_), .ZN(new_n14516_));
  NAND2_X1   g14221(.A1(new_n14513_), .A2(new_n14516_), .ZN(new_n14517_));
  NAND2_X1   g14222(.A1(new_n14517_), .A2(new_n14252_), .ZN(new_n14518_));
  INV_X1     g14223(.I(new_n14252_), .ZN(new_n14519_));
  NOR3_X1    g14224(.A1(new_n14507_), .A2(new_n14504_), .A3(new_n14511_), .ZN(new_n14520_));
  AOI21_X1   g14225(.A1(new_n14514_), .A2(new_n14515_), .B(new_n14512_), .ZN(new_n14521_));
  OAI21_X1   g14226(.A1(new_n14520_), .A2(new_n14521_), .B(new_n14519_), .ZN(new_n14522_));
  OAI22_X1   g14227(.A1(new_n1055_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n1061_), .ZN(new_n14523_));
  OAI21_X1   g14228(.A1(new_n7870_), .A2(new_n1332_), .B(new_n14523_), .ZN(new_n14524_));
  AOI21_X1   g14229(.A1(new_n14524_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n14525_));
  XOR2_X1    g14230(.A1(new_n8568_), .A2(new_n14525_), .Z(new_n14526_));
  AOI21_X1   g14231(.A1(new_n14518_), .A2(new_n14522_), .B(new_n14526_), .ZN(new_n14527_));
  OAI21_X1   g14232(.A1(new_n14250_), .A2(new_n14251_), .B(new_n14527_), .ZN(new_n14528_));
  NOR2_X1    g14233(.A1(new_n14133_), .A2(new_n13715_), .ZN(new_n14529_));
  NOR2_X1    g14234(.A1(new_n14529_), .A2(new_n13736_), .ZN(new_n14530_));
  AOI21_X1   g14235(.A1(new_n14513_), .A2(new_n14516_), .B(new_n14519_), .ZN(new_n14531_));
  NAND3_X1   g14236(.A1(new_n14514_), .A2(new_n14515_), .A3(new_n14512_), .ZN(new_n14532_));
  OAI21_X1   g14237(.A1(new_n14507_), .A2(new_n14504_), .B(new_n14511_), .ZN(new_n14533_));
  AOI21_X1   g14238(.A1(new_n14533_), .A2(new_n14532_), .B(new_n14252_), .ZN(new_n14534_));
  INV_X1     g14239(.I(new_n14526_), .ZN(new_n14535_));
  OAI21_X1   g14240(.A1(new_n14531_), .A2(new_n14534_), .B(new_n14535_), .ZN(new_n14536_));
  NAND3_X1   g14241(.A1(new_n14530_), .A2(new_n14536_), .A3(new_n14249_), .ZN(new_n14537_));
  AOI21_X1   g14242(.A1(new_n14528_), .A2(new_n14537_), .B(new_n14248_), .ZN(new_n14538_));
  AOI21_X1   g14243(.A1(new_n14530_), .A2(new_n14249_), .B(new_n14536_), .ZN(new_n14539_));
  NOR3_X1    g14244(.A1(new_n14527_), .A2(new_n14250_), .A3(new_n14251_), .ZN(new_n14540_));
  NOR3_X1    g14245(.A1(new_n14539_), .A2(new_n14540_), .A3(new_n14247_), .ZN(new_n14541_));
  OAI22_X1   g14246(.A1(new_n970_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n820_), .ZN(new_n14542_));
  OAI21_X1   g14247(.A1(new_n8948_), .A2(new_n894_), .B(new_n14542_), .ZN(new_n14543_));
  AOI21_X1   g14248(.A1(new_n14543_), .A2(new_n827_), .B(new_n970_), .ZN(new_n14544_));
  XNOR2_X1   g14249(.A1(new_n9642_), .A2(new_n14544_), .ZN(new_n14545_));
  INV_X1     g14250(.I(new_n14545_), .ZN(new_n14546_));
  OAI21_X1   g14251(.A1(new_n14538_), .A2(new_n14541_), .B(new_n14546_), .ZN(new_n14547_));
  AOI21_X1   g14252(.A1(new_n14173_), .A2(new_n14245_), .B(new_n14547_), .ZN(new_n14548_));
  NAND2_X1   g14253(.A1(new_n14173_), .A2(new_n14245_), .ZN(new_n14549_));
  OAI21_X1   g14254(.A1(new_n14539_), .A2(new_n14540_), .B(new_n14247_), .ZN(new_n14550_));
  NAND3_X1   g14255(.A1(new_n14528_), .A2(new_n14537_), .A3(new_n14248_), .ZN(new_n14551_));
  AOI21_X1   g14256(.A1(new_n14550_), .A2(new_n14551_), .B(new_n14545_), .ZN(new_n14552_));
  NOR2_X1    g14257(.A1(new_n14549_), .A2(new_n14552_), .ZN(new_n14553_));
  OAI21_X1   g14258(.A1(new_n14548_), .A2(new_n14553_), .B(new_n14145_), .ZN(new_n14554_));
  NAND2_X1   g14259(.A1(new_n14549_), .A2(new_n14552_), .ZN(new_n14555_));
  NAND3_X1   g14260(.A1(new_n14547_), .A2(new_n14173_), .A3(new_n14245_), .ZN(new_n14556_));
  NAND3_X1   g14261(.A1(new_n14555_), .A2(new_n14556_), .A3(new_n14153_), .ZN(new_n14557_));
  OAI22_X1   g14262(.A1(new_n607_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n610_), .ZN(new_n14558_));
  OAI21_X1   g14263(.A1(new_n10031_), .A2(new_n684_), .B(new_n14558_), .ZN(new_n14559_));
  AOI21_X1   g14264(.A1(new_n14559_), .A2(new_n612_), .B(new_n607_), .ZN(new_n14560_));
  XNOR2_X1   g14265(.A1(new_n10866_), .A2(new_n14560_), .ZN(new_n14561_));
  INV_X1     g14266(.I(new_n14561_), .ZN(new_n14562_));
  NAND3_X1   g14267(.A1(new_n14554_), .A2(new_n14557_), .A3(new_n14562_), .ZN(new_n14563_));
  AOI21_X1   g14268(.A1(new_n14555_), .A2(new_n14556_), .B(new_n14153_), .ZN(new_n14564_));
  NOR3_X1    g14269(.A1(new_n14548_), .A2(new_n14553_), .A3(new_n14145_), .ZN(new_n14565_));
  OAI21_X1   g14270(.A1(new_n14565_), .A2(new_n14564_), .B(new_n14561_), .ZN(new_n14566_));
  NAND2_X1   g14271(.A1(new_n14566_), .A2(new_n14563_), .ZN(new_n14567_));
  AOI21_X1   g14272(.A1(new_n14177_), .A2(new_n13753_), .B(new_n13758_), .ZN(new_n14568_));
  NAND3_X1   g14273(.A1(new_n14176_), .A2(new_n14172_), .A3(new_n14167_), .ZN(new_n14569_));
  NAND2_X1   g14274(.A1(new_n13405_), .A2(new_n14569_), .ZN(new_n14570_));
  XOR2_X1    g14275(.A1(new_n14173_), .A2(new_n14245_), .Z(new_n14571_));
  NAND2_X1   g14276(.A1(new_n14571_), .A2(new_n14149_), .ZN(new_n14572_));
  OAI21_X1   g14277(.A1(new_n14570_), .A2(new_n14568_), .B(new_n14572_), .ZN(new_n14573_));
  OAI22_X1   g14278(.A1(new_n448_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n450_), .ZN(new_n14574_));
  OAI21_X1   g14279(.A1(new_n11738_), .A2(new_n496_), .B(new_n14574_), .ZN(new_n14575_));
  AOI21_X1   g14280(.A1(new_n14575_), .A2(new_n452_), .B(new_n448_), .ZN(new_n14576_));
  XNOR2_X1   g14281(.A1(new_n12128_), .A2(new_n14576_), .ZN(new_n14577_));
  NOR2_X1    g14282(.A1(new_n14573_), .A2(new_n14577_), .ZN(new_n14578_));
  OAI21_X1   g14283(.A1(new_n14161_), .A2(new_n14167_), .B(new_n13757_), .ZN(new_n14579_));
  NAND3_X1   g14284(.A1(new_n14579_), .A2(new_n13405_), .A3(new_n14569_), .ZN(new_n14580_));
  INV_X1     g14285(.I(new_n14577_), .ZN(new_n14581_));
  AOI21_X1   g14286(.A1(new_n14580_), .A2(new_n14572_), .B(new_n14581_), .ZN(new_n14582_));
  OAI21_X1   g14287(.A1(new_n14578_), .A2(new_n14582_), .B(new_n14567_), .ZN(new_n14583_));
  NOR3_X1    g14288(.A1(new_n14565_), .A2(new_n14564_), .A3(new_n14561_), .ZN(new_n14584_));
  AOI21_X1   g14289(.A1(new_n14554_), .A2(new_n14557_), .B(new_n14562_), .ZN(new_n14585_));
  NOR2_X1    g14290(.A1(new_n14584_), .A2(new_n14585_), .ZN(new_n14586_));
  AOI21_X1   g14291(.A1(new_n14580_), .A2(new_n14572_), .B(new_n14577_), .ZN(new_n14587_));
  NOR2_X1    g14292(.A1(new_n14573_), .A2(new_n14581_), .ZN(new_n14588_));
  OAI21_X1   g14293(.A1(new_n14588_), .A2(new_n14587_), .B(new_n14586_), .ZN(new_n14589_));
  INV_X1     g14294(.I(new_n14209_), .ZN(new_n14590_));
  AOI21_X1   g14295(.A1(new_n14207_), .A2(new_n14590_), .B(new_n14210_), .ZN(new_n14591_));
  INV_X1     g14296(.I(\b[63] ), .ZN(new_n14592_));
  NOR2_X1    g14297(.A1(new_n14592_), .A2(\b[62] ), .ZN(new_n14593_));
  NOR2_X1    g14298(.A1(new_n14208_), .A2(\b[63] ), .ZN(new_n14594_));
  NOR2_X1    g14299(.A1(new_n14593_), .A2(new_n14594_), .ZN(new_n14595_));
  NOR2_X1    g14300(.A1(new_n14208_), .A2(new_n14592_), .ZN(new_n14596_));
  NOR2_X1    g14301(.A1(\b[62] ), .A2(\b[63] ), .ZN(new_n14597_));
  OAI21_X1   g14302(.A1(new_n14596_), .A2(new_n14597_), .B(new_n14591_), .ZN(new_n14598_));
  OAI21_X1   g14303(.A1(new_n14591_), .A2(new_n14595_), .B(new_n14598_), .ZN(new_n14599_));
  NAND2_X1   g14304(.A1(new_n286_), .A2(\b[62] ), .ZN(new_n14600_));
  AOI22_X1   g14305(.A1(new_n304_), .A2(\b[61] ), .B1(new_n262_), .B2(\b[63] ), .ZN(new_n14601_));
  AOI21_X1   g14306(.A1(new_n14600_), .A2(new_n14601_), .B(new_n426_), .ZN(new_n14602_));
  NAND2_X1   g14307(.A1(new_n14599_), .A2(new_n14602_), .ZN(new_n14603_));
  XOR2_X1    g14308(.A1(new_n14603_), .A2(\a[2] ), .Z(new_n14604_));
  INV_X1     g14309(.I(new_n14604_), .ZN(new_n14605_));
  NAND3_X1   g14310(.A1(new_n14583_), .A2(new_n14589_), .A3(new_n14605_), .ZN(new_n14606_));
  NAND3_X1   g14311(.A1(new_n14580_), .A2(new_n14572_), .A3(new_n14581_), .ZN(new_n14607_));
  NAND2_X1   g14312(.A1(new_n14573_), .A2(new_n14577_), .ZN(new_n14608_));
  AOI21_X1   g14313(.A1(new_n14608_), .A2(new_n14607_), .B(new_n14586_), .ZN(new_n14609_));
  NAND2_X1   g14314(.A1(new_n14573_), .A2(new_n14581_), .ZN(new_n14610_));
  NAND3_X1   g14315(.A1(new_n14580_), .A2(new_n14572_), .A3(new_n14577_), .ZN(new_n14611_));
  AOI21_X1   g14316(.A1(new_n14610_), .A2(new_n14611_), .B(new_n14567_), .ZN(new_n14612_));
  OAI21_X1   g14317(.A1(new_n14609_), .A2(new_n14612_), .B(new_n14604_), .ZN(new_n14613_));
  AOI21_X1   g14318(.A1(new_n14613_), .A2(new_n14606_), .B(new_n14244_), .ZN(new_n14614_));
  NOR3_X1    g14319(.A1(new_n14193_), .A2(new_n14192_), .A3(new_n14196_), .ZN(new_n14615_));
  NOR2_X1    g14320(.A1(new_n14615_), .A2(new_n14194_), .ZN(new_n14616_));
  NOR3_X1    g14321(.A1(new_n14609_), .A2(new_n14612_), .A3(new_n14604_), .ZN(new_n14617_));
  AOI21_X1   g14322(.A1(new_n14583_), .A2(new_n14589_), .B(new_n14605_), .ZN(new_n14618_));
  NOR3_X1    g14323(.A1(new_n14618_), .A2(new_n14617_), .A3(new_n14616_), .ZN(new_n14619_));
  OAI21_X1   g14324(.A1(new_n14614_), .A2(new_n14619_), .B(new_n14241_), .ZN(new_n14620_));
  INV_X1     g14325(.I(new_n14241_), .ZN(new_n14621_));
  OAI21_X1   g14326(.A1(new_n14618_), .A2(new_n14617_), .B(new_n14616_), .ZN(new_n14622_));
  NAND3_X1   g14327(.A1(new_n14613_), .A2(new_n14606_), .A3(new_n14244_), .ZN(new_n14623_));
  NAND3_X1   g14328(.A1(new_n14622_), .A2(new_n14623_), .A3(new_n14621_), .ZN(new_n14624_));
  INV_X1     g14329(.I(new_n14227_), .ZN(new_n14625_));
  AOI21_X1   g14330(.A1(new_n13824_), .A2(new_n14228_), .B(new_n14625_), .ZN(new_n14626_));
  AOI21_X1   g14331(.A1(new_n14620_), .A2(new_n14624_), .B(new_n14626_), .ZN(new_n14627_));
  AOI21_X1   g14332(.A1(new_n14622_), .A2(new_n14623_), .B(new_n14621_), .ZN(new_n14628_));
  NOR3_X1    g14333(.A1(new_n14614_), .A2(new_n14619_), .A3(new_n14241_), .ZN(new_n14629_));
  NAND2_X1   g14334(.A1(new_n13824_), .A2(new_n14228_), .ZN(new_n14630_));
  NAND2_X1   g14335(.A1(new_n14630_), .A2(new_n14227_), .ZN(new_n14631_));
  NOR3_X1    g14336(.A1(new_n14629_), .A2(new_n14628_), .A3(new_n14631_), .ZN(new_n14632_));
  OAI21_X1   g14337(.A1(new_n14627_), .A2(new_n14632_), .B(new_n14236_), .ZN(new_n14633_));
  XOR2_X1    g14338(.A1(new_n14633_), .A2(new_n14232_), .Z(new_n14634_));
  XOR2_X1    g14339(.A1(new_n14634_), .A2(new_n13820_), .Z(\f[63] ));
  NOR2_X1    g14340(.A1(new_n13404_), .A2(new_n13800_), .ZN(new_n14636_));
  OAI21_X1   g14341(.A1(new_n13400_), .A2(new_n13399_), .B(new_n13023_), .ZN(new_n14637_));
  NAND3_X1   g14342(.A1(new_n13396_), .A2(new_n13397_), .A3(new_n13388_), .ZN(new_n14638_));
  NAND2_X1   g14343(.A1(new_n14637_), .A2(new_n14638_), .ZN(new_n14639_));
  INV_X1     g14344(.I(new_n13803_), .ZN(new_n14640_));
  NAND3_X1   g14345(.A1(new_n14639_), .A2(new_n14640_), .A3(new_n13395_), .ZN(new_n14641_));
  AOI21_X1   g14346(.A1(new_n13404_), .A2(new_n13800_), .B(new_n14641_), .ZN(new_n14642_));
  NOR3_X1    g14347(.A1(new_n14632_), .A2(new_n14627_), .A3(new_n14231_), .ZN(new_n14643_));
  OAI21_X1   g14348(.A1(new_n14632_), .A2(new_n14627_), .B(new_n14231_), .ZN(new_n14644_));
  AOI21_X1   g14349(.A1(new_n13821_), .A2(new_n14644_), .B(new_n14643_), .ZN(new_n14645_));
  OAI21_X1   g14350(.A1(new_n14642_), .A2(new_n14636_), .B(new_n14645_), .ZN(new_n14646_));
  OAI22_X1   g14351(.A1(new_n13367_), .A2(new_n341_), .B1(new_n404_), .B2(new_n13785_), .ZN(new_n14647_));
  OAI21_X1   g14352(.A1(new_n12970_), .A2(new_n366_), .B(new_n14647_), .ZN(new_n14648_));
  AOI21_X1   g14353(.A1(new_n14648_), .A2(new_n334_), .B(new_n341_), .ZN(new_n14649_));
  XOR2_X1    g14354(.A1(new_n13784_), .A2(new_n14649_), .Z(new_n14650_));
  NAND2_X1   g14355(.A1(new_n14621_), .A2(new_n14581_), .ZN(new_n14651_));
  XOR2_X1    g14356(.A1(new_n14586_), .A2(new_n14573_), .Z(new_n14652_));
  OAI21_X1   g14357(.A1(new_n14621_), .A2(new_n14581_), .B(new_n14652_), .ZN(new_n14653_));
  NAND2_X1   g14358(.A1(new_n14653_), .A2(new_n14651_), .ZN(new_n14654_));
  OAI21_X1   g14359(.A1(new_n14573_), .A2(new_n14585_), .B(new_n14563_), .ZN(new_n14655_));
  AOI21_X1   g14360(.A1(new_n14550_), .A2(new_n14551_), .B(new_n14145_), .ZN(new_n14656_));
  NOR3_X1    g14361(.A1(new_n14538_), .A2(new_n14541_), .A3(new_n14153_), .ZN(new_n14657_));
  NOR3_X1    g14362(.A1(new_n14549_), .A2(new_n14545_), .A3(new_n14657_), .ZN(new_n14658_));
  NOR2_X1    g14363(.A1(new_n14658_), .A2(new_n14656_), .ZN(new_n14659_));
  NAND2_X1   g14364(.A1(new_n14518_), .A2(new_n14522_), .ZN(new_n14660_));
  NAND3_X1   g14365(.A1(new_n14530_), .A2(new_n14660_), .A3(new_n14249_), .ZN(new_n14661_));
  INV_X1     g14366(.I(new_n14661_), .ZN(new_n14662_));
  AOI21_X1   g14367(.A1(new_n14530_), .A2(new_n14249_), .B(new_n14660_), .ZN(new_n14663_));
  NAND2_X1   g14368(.A1(new_n14248_), .A2(new_n14535_), .ZN(new_n14664_));
  NOR2_X1    g14369(.A1(new_n14663_), .A2(new_n14664_), .ZN(new_n14665_));
  NOR2_X1    g14370(.A1(new_n14665_), .A2(new_n14662_), .ZN(new_n14666_));
  AOI21_X1   g14371(.A1(new_n14252_), .A2(new_n14533_), .B(new_n14520_), .ZN(new_n14667_));
  INV_X1     g14372(.I(new_n14667_), .ZN(new_n14668_));
  OAI22_X1   g14373(.A1(new_n1712_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n1707_), .ZN(new_n14669_));
  OAI21_X1   g14374(.A1(new_n6229_), .A2(new_n1850_), .B(new_n14669_), .ZN(new_n14670_));
  AOI21_X1   g14375(.A1(new_n14670_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n14671_));
  XOR2_X1    g14376(.A1(new_n6851_), .A2(new_n14671_), .Z(new_n14672_));
  INV_X1     g14377(.I(new_n14672_), .ZN(new_n14673_));
  OAI22_X1   g14378(.A1(new_n2171_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n2166_), .ZN(new_n14674_));
  OAI21_X1   g14379(.A1(new_n5353_), .A2(new_n2322_), .B(new_n14674_), .ZN(new_n14675_));
  AOI21_X1   g14380(.A1(new_n14675_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n14676_));
  XOR2_X1    g14381(.A1(new_n5926_), .A2(new_n14676_), .Z(new_n14677_));
  INV_X1     g14382(.I(new_n14677_), .ZN(new_n14678_));
  NOR2_X1    g14383(.A1(new_n14258_), .A2(new_n14451_), .ZN(new_n14679_));
  NAND2_X1   g14384(.A1(new_n14444_), .A2(new_n14259_), .ZN(new_n14680_));
  OAI22_X1   g14385(.A1(new_n14680_), .A2(new_n14258_), .B1(new_n14444_), .B2(new_n14679_), .ZN(new_n14681_));
  NAND2_X1   g14386(.A1(new_n14465_), .A2(new_n14681_), .ZN(new_n14682_));
  NOR2_X1    g14387(.A1(new_n14465_), .A2(new_n14681_), .ZN(new_n14683_));
  NAND2_X1   g14388(.A1(new_n14473_), .A2(new_n14449_), .ZN(new_n14684_));
  OAI21_X1   g14389(.A1(new_n14683_), .A2(new_n14684_), .B(new_n14682_), .ZN(new_n14685_));
  INV_X1     g14390(.I(new_n14685_), .ZN(new_n14686_));
  NOR2_X1    g14391(.A1(new_n14482_), .A2(new_n14475_), .ZN(new_n14687_));
  NOR2_X1    g14392(.A1(new_n14068_), .A2(new_n14479_), .ZN(new_n14688_));
  INV_X1     g14393(.I(new_n14688_), .ZN(new_n14689_));
  AOI21_X1   g14394(.A1(new_n14482_), .A2(new_n14475_), .B(new_n14689_), .ZN(new_n14690_));
  OAI22_X1   g14395(.A1(new_n5420_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n5107_), .ZN(new_n14691_));
  OAI21_X1   g14396(.A1(new_n2439_), .A2(new_n5112_), .B(new_n14691_), .ZN(new_n14692_));
  AOI21_X1   g14397(.A1(new_n14692_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n14693_));
  XNOR2_X1   g14398(.A1(new_n2846_), .A2(new_n14693_), .ZN(new_n14694_));
  INV_X1     g14399(.I(new_n14694_), .ZN(new_n14695_));
  NAND2_X1   g14400(.A1(new_n14381_), .A2(new_n14377_), .ZN(new_n14696_));
  NAND2_X1   g14401(.A1(new_n14388_), .A2(new_n14696_), .ZN(new_n14697_));
  NOR2_X1    g14402(.A1(new_n14398_), .A2(new_n14385_), .ZN(new_n14698_));
  OAI21_X1   g14403(.A1(new_n14388_), .A2(new_n14696_), .B(new_n14698_), .ZN(new_n14699_));
  NAND2_X1   g14404(.A1(new_n14699_), .A2(new_n14697_), .ZN(new_n14700_));
  INV_X1     g14405(.I(new_n14700_), .ZN(new_n14701_));
  OAI21_X1   g14406(.A1(new_n14397_), .A2(new_n14401_), .B(new_n14005_), .ZN(new_n14702_));
  NOR2_X1    g14407(.A1(new_n14397_), .A2(new_n14401_), .ZN(new_n14703_));
  NAND2_X1   g14408(.A1(new_n14703_), .A2(new_n13998_), .ZN(new_n14704_));
  NAND4_X1   g14409(.A1(new_n14704_), .A2(new_n13595_), .A3(new_n14264_), .A4(new_n14406_), .ZN(new_n14705_));
  NAND2_X1   g14410(.A1(new_n14705_), .A2(new_n14702_), .ZN(new_n14706_));
  OAI21_X1   g14411(.A1(new_n14373_), .A2(new_n14374_), .B(new_n14371_), .ZN(new_n14707_));
  AOI21_X1   g14412(.A1(new_n14391_), .A2(new_n14707_), .B(new_n14379_), .ZN(new_n14708_));
  INV_X1     g14413(.I(new_n14708_), .ZN(new_n14709_));
  OAI22_X1   g14414(.A1(new_n8644_), .A2(new_n1017_), .B1(new_n1109_), .B2(new_n9388_), .ZN(new_n14710_));
  OAI21_X1   g14415(.A1(new_n930_), .A2(new_n10154_), .B(new_n14710_), .ZN(new_n14711_));
  AOI21_X1   g14416(.A1(new_n14711_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n14712_));
  XOR2_X1    g14417(.A1(new_n1114_), .A2(new_n14712_), .Z(new_n14713_));
  INV_X1     g14418(.I(new_n14713_), .ZN(new_n14714_));
  OAI21_X1   g14419(.A1(new_n14319_), .A2(new_n14315_), .B(new_n14271_), .ZN(new_n14715_));
  NAND3_X1   g14420(.A1(new_n14272_), .A2(new_n14327_), .A3(new_n14329_), .ZN(new_n14716_));
  NAND4_X1   g14421(.A1(new_n14716_), .A2(new_n13873_), .A3(new_n13929_), .A4(new_n14324_), .ZN(new_n14717_));
  NAND2_X1   g14422(.A1(new_n14717_), .A2(new_n14715_), .ZN(new_n14718_));
  INV_X1     g14423(.I(new_n14718_), .ZN(new_n14719_));
  NOR2_X1    g14424(.A1(new_n14344_), .A2(new_n14343_), .ZN(new_n14720_));
  NOR2_X1    g14425(.A1(new_n14720_), .A2(new_n13947_), .ZN(new_n14721_));
  INV_X1     g14426(.I(new_n14721_), .ZN(new_n14722_));
  NAND2_X1   g14427(.A1(new_n14720_), .A2(new_n13947_), .ZN(new_n14723_));
  NAND3_X1   g14428(.A1(new_n14723_), .A2(new_n14342_), .A3(new_n14345_), .ZN(new_n14724_));
  NAND2_X1   g14429(.A1(new_n14724_), .A2(new_n14722_), .ZN(new_n14725_));
  AOI21_X1   g14430(.A1(new_n14274_), .A2(new_n13910_), .B(new_n14313_), .ZN(new_n14726_));
  NOR2_X1    g14431(.A1(new_n14726_), .A2(new_n14308_), .ZN(new_n14727_));
  NOR2_X1    g14432(.A1(new_n14275_), .A2(new_n14302_), .ZN(new_n14728_));
  NOR2_X1    g14433(.A1(new_n14728_), .A2(new_n14301_), .ZN(new_n14729_));
  NAND2_X1   g14434(.A1(new_n14287_), .A2(new_n14276_), .ZN(new_n14730_));
  NAND2_X1   g14435(.A1(new_n14730_), .A2(new_n14288_), .ZN(new_n14731_));
  AOI22_X1   g14436(.A1(new_n13472_), .A2(new_n10957_), .B1(\b[2] ), .B2(new_n13884_), .ZN(new_n14732_));
  OAI21_X1   g14437(.A1(new_n14732_), .A2(\a[62] ), .B(new_n13466_), .ZN(new_n14733_));
  XOR2_X1    g14438(.A1(new_n14733_), .A2(new_n329_), .Z(new_n14734_));
  NOR2_X1    g14439(.A1(new_n13476_), .A2(new_n258_), .ZN(new_n14735_));
  NAND2_X1   g14440(.A1(\a[62] ), .A2(\a[63] ), .ZN(new_n14736_));
  XOR2_X1    g14441(.A1(new_n14736_), .A2(new_n258_), .Z(new_n14737_));
  NAND2_X1   g14442(.A1(new_n14737_), .A2(\b[1] ), .ZN(new_n14738_));
  XOR2_X1    g14443(.A1(new_n14738_), .A2(new_n14735_), .Z(new_n14739_));
  XNOR2_X1   g14444(.A1(new_n14734_), .A2(new_n14739_), .ZN(new_n14740_));
  INV_X1     g14445(.I(new_n14740_), .ZN(new_n14741_));
  NAND2_X1   g14446(.A1(new_n14731_), .A2(new_n14741_), .ZN(new_n14742_));
  INV_X1     g14447(.I(new_n14742_), .ZN(new_n14743_));
  NOR2_X1    g14448(.A1(new_n14734_), .A2(new_n14739_), .ZN(new_n14744_));
  INV_X1     g14449(.I(new_n14744_), .ZN(new_n14745_));
  NAND2_X1   g14450(.A1(new_n14734_), .A2(new_n14739_), .ZN(new_n14746_));
  AOI21_X1   g14451(.A1(new_n14745_), .A2(new_n14746_), .B(new_n14731_), .ZN(new_n14747_));
  NOR2_X1    g14452(.A1(new_n14743_), .A2(new_n14747_), .ZN(new_n14748_));
  OAI22_X1   g14453(.A1(new_n12226_), .A2(new_n509_), .B1(new_n12637_), .B2(new_n419_), .ZN(new_n14749_));
  AOI21_X1   g14454(.A1(new_n14749_), .A2(new_n12222_), .B(new_n12643_), .ZN(new_n14750_));
  XOR2_X1    g14455(.A1(new_n471_), .A2(new_n14750_), .Z(new_n14751_));
  XOR2_X1    g14456(.A1(new_n14748_), .A2(new_n14751_), .Z(new_n14752_));
  NOR2_X1    g14457(.A1(new_n14752_), .A2(new_n14729_), .ZN(new_n14753_));
  INV_X1     g14458(.I(new_n14729_), .ZN(new_n14754_));
  INV_X1     g14459(.I(new_n14751_), .ZN(new_n14755_));
  NAND2_X1   g14460(.A1(new_n14748_), .A2(new_n14755_), .ZN(new_n14756_));
  OAI21_X1   g14461(.A1(new_n14743_), .A2(new_n14747_), .B(new_n14751_), .ZN(new_n14757_));
  AOI21_X1   g14462(.A1(new_n14756_), .A2(new_n14757_), .B(new_n14754_), .ZN(new_n14758_));
  NOR2_X1    g14463(.A1(new_n14758_), .A2(new_n14753_), .ZN(new_n14759_));
  AOI22_X1   g14464(.A1(new_n10969_), .A2(new_n13503_), .B1(new_n11394_), .B2(\b[8] ), .ZN(new_n14760_));
  OAI21_X1   g14465(.A1(new_n14760_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n14761_));
  XOR2_X1    g14466(.A1(new_n660_), .A2(new_n14761_), .Z(new_n14762_));
  XOR2_X1    g14467(.A1(new_n14759_), .A2(new_n14762_), .Z(new_n14763_));
  NOR2_X1    g14468(.A1(new_n14763_), .A2(new_n14727_), .ZN(new_n14764_));
  INV_X1     g14469(.I(new_n14727_), .ZN(new_n14765_));
  INV_X1     g14470(.I(new_n14762_), .ZN(new_n14766_));
  NAND2_X1   g14471(.A1(new_n14759_), .A2(new_n14766_), .ZN(new_n14767_));
  INV_X1     g14472(.I(new_n14759_), .ZN(new_n14768_));
  NAND2_X1   g14473(.A1(new_n14768_), .A2(new_n14762_), .ZN(new_n14769_));
  AOI21_X1   g14474(.A1(new_n14769_), .A2(new_n14767_), .B(new_n14765_), .ZN(new_n14770_));
  NOR2_X1    g14475(.A1(new_n14764_), .A2(new_n14770_), .ZN(new_n14771_));
  AOI22_X1   g14476(.A1(new_n11415_), .A2(new_n927_), .B1(\b[11] ), .B2(new_n10145_), .ZN(new_n14772_));
  OAI21_X1   g14477(.A1(new_n14772_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n14773_));
  XOR2_X1    g14478(.A1(new_n860_), .A2(new_n14773_), .Z(new_n14774_));
  XOR2_X1    g14479(.A1(new_n14771_), .A2(new_n14774_), .Z(new_n14775_));
  NOR2_X1    g14480(.A1(new_n14725_), .A2(new_n14775_), .ZN(new_n14776_));
  NAND2_X1   g14481(.A1(new_n14725_), .A2(new_n14775_), .ZN(new_n14777_));
  INV_X1     g14482(.I(new_n14777_), .ZN(new_n14778_));
  OAI21_X1   g14483(.A1(new_n14778_), .A2(new_n14776_), .B(new_n14719_), .ZN(new_n14779_));
  INV_X1     g14484(.I(new_n14776_), .ZN(new_n14780_));
  NAND3_X1   g14485(.A1(new_n14780_), .A2(new_n14718_), .A3(new_n14777_), .ZN(new_n14781_));
  AOI21_X1   g14486(.A1(new_n14779_), .A2(new_n14781_), .B(new_n14714_), .ZN(new_n14782_));
  AOI21_X1   g14487(.A1(new_n14780_), .A2(new_n14777_), .B(new_n14718_), .ZN(new_n14783_));
  NOR3_X1    g14488(.A1(new_n14778_), .A2(new_n14719_), .A3(new_n14776_), .ZN(new_n14784_));
  NOR3_X1    g14489(.A1(new_n14783_), .A2(new_n14784_), .A3(new_n14713_), .ZN(new_n14785_));
  OAI22_X1   g14490(.A1(new_n7619_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n8309_), .ZN(new_n14786_));
  OAI21_X1   g14491(.A1(new_n1189_), .A2(new_n7947_), .B(new_n14786_), .ZN(new_n14787_));
  AOI21_X1   g14492(.A1(new_n14787_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n14788_));
  XNOR2_X1   g14493(.A1(new_n1421_), .A2(new_n14788_), .ZN(new_n14789_));
  INV_X1     g14494(.I(new_n14789_), .ZN(new_n14790_));
  OAI21_X1   g14495(.A1(new_n14782_), .A2(new_n14785_), .B(new_n14790_), .ZN(new_n14791_));
  OAI21_X1   g14496(.A1(new_n14783_), .A2(new_n14784_), .B(new_n14713_), .ZN(new_n14792_));
  NAND3_X1   g14497(.A1(new_n14779_), .A2(new_n14781_), .A3(new_n14714_), .ZN(new_n14793_));
  NAND3_X1   g14498(.A1(new_n14792_), .A2(new_n14793_), .A3(new_n14789_), .ZN(new_n14794_));
  NAND2_X1   g14499(.A1(new_n14360_), .A2(new_n14359_), .ZN(new_n14795_));
  NAND2_X1   g14500(.A1(new_n13958_), .A2(new_n14795_), .ZN(new_n14796_));
  NOR2_X1    g14501(.A1(new_n14270_), .A2(new_n14355_), .ZN(new_n14797_));
  OAI21_X1   g14502(.A1(new_n13958_), .A2(new_n14795_), .B(new_n14797_), .ZN(new_n14798_));
  NAND2_X1   g14503(.A1(new_n14798_), .A2(new_n14796_), .ZN(new_n14799_));
  OAI22_X1   g14504(.A1(new_n6644_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n6647_), .ZN(new_n14800_));
  OAI21_X1   g14505(.A1(new_n1525_), .A2(new_n7284_), .B(new_n14800_), .ZN(new_n14801_));
  AOI21_X1   g14506(.A1(new_n14801_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n14802_));
  XOR2_X1    g14507(.A1(new_n1808_), .A2(new_n14802_), .Z(new_n14803_));
  XOR2_X1    g14508(.A1(new_n14799_), .A2(new_n14803_), .Z(new_n14804_));
  AOI21_X1   g14509(.A1(new_n14791_), .A2(new_n14794_), .B(new_n14804_), .ZN(new_n14805_));
  NAND2_X1   g14510(.A1(new_n14791_), .A2(new_n14794_), .ZN(new_n14806_));
  INV_X1     g14511(.I(new_n14803_), .ZN(new_n14807_));
  XOR2_X1    g14512(.A1(new_n14799_), .A2(new_n14807_), .Z(new_n14808_));
  NOR2_X1    g14513(.A1(new_n14806_), .A2(new_n14808_), .ZN(new_n14809_));
  NOR2_X1    g14514(.A1(new_n14809_), .A2(new_n14805_), .ZN(new_n14810_));
  OAI22_X1   g14515(.A1(new_n5993_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n5991_), .ZN(new_n14811_));
  OAI21_X1   g14516(.A1(new_n1936_), .A2(new_n5997_), .B(new_n14811_), .ZN(new_n14812_));
  AOI21_X1   g14517(.A1(new_n14812_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n14813_));
  XNOR2_X1   g14518(.A1(new_n2280_), .A2(new_n14813_), .ZN(new_n14814_));
  NOR2_X1    g14519(.A1(new_n14810_), .A2(new_n14814_), .ZN(new_n14815_));
  INV_X1     g14520(.I(new_n14814_), .ZN(new_n14816_));
  NOR3_X1    g14521(.A1(new_n14809_), .A2(new_n14805_), .A3(new_n14816_), .ZN(new_n14817_));
  OAI21_X1   g14522(.A1(new_n14815_), .A2(new_n14817_), .B(new_n14709_), .ZN(new_n14818_));
  XOR2_X1    g14523(.A1(new_n14810_), .A2(new_n14816_), .Z(new_n14819_));
  OAI21_X1   g14524(.A1(new_n14819_), .A2(new_n14709_), .B(new_n14818_), .ZN(new_n14820_));
  INV_X1     g14525(.I(new_n14820_), .ZN(new_n14821_));
  NOR2_X1    g14526(.A1(new_n14706_), .A2(new_n14821_), .ZN(new_n14822_));
  NAND2_X1   g14527(.A1(new_n14706_), .A2(new_n14821_), .ZN(new_n14823_));
  INV_X1     g14528(.I(new_n14823_), .ZN(new_n14824_));
  OAI21_X1   g14529(.A1(new_n14824_), .A2(new_n14822_), .B(new_n14701_), .ZN(new_n14825_));
  INV_X1     g14530(.I(new_n14822_), .ZN(new_n14826_));
  NAND3_X1   g14531(.A1(new_n14826_), .A2(new_n14700_), .A3(new_n14823_), .ZN(new_n14827_));
  AOI21_X1   g14532(.A1(new_n14825_), .A2(new_n14827_), .B(new_n14695_), .ZN(new_n14828_));
  AOI21_X1   g14533(.A1(new_n14826_), .A2(new_n14823_), .B(new_n14700_), .ZN(new_n14829_));
  NOR3_X1    g14534(.A1(new_n14824_), .A2(new_n14701_), .A3(new_n14822_), .ZN(new_n14830_));
  NOR3_X1    g14535(.A1(new_n14829_), .A2(new_n14830_), .A3(new_n14694_), .ZN(new_n14831_));
  OAI22_X1   g14536(.A1(new_n4072_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n4067_), .ZN(new_n14832_));
  OAI21_X1   g14537(.A1(new_n3018_), .A2(new_n4318_), .B(new_n14832_), .ZN(new_n14833_));
  AOI21_X1   g14538(.A1(new_n14833_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n14834_));
  XNOR2_X1   g14539(.A1(new_n3514_), .A2(new_n14834_), .ZN(new_n14835_));
  INV_X1     g14540(.I(new_n14835_), .ZN(new_n14836_));
  OAI21_X1   g14541(.A1(new_n14828_), .A2(new_n14831_), .B(new_n14836_), .ZN(new_n14837_));
  OAI21_X1   g14542(.A1(new_n14829_), .A2(new_n14830_), .B(new_n14694_), .ZN(new_n14838_));
  NAND3_X1   g14543(.A1(new_n14825_), .A2(new_n14827_), .A3(new_n14695_), .ZN(new_n14839_));
  NAND3_X1   g14544(.A1(new_n14838_), .A2(new_n14839_), .A3(new_n14835_), .ZN(new_n14840_));
  AOI21_X1   g14545(.A1(new_n14414_), .A2(new_n14417_), .B(new_n14016_), .ZN(new_n14841_));
  NOR3_X1    g14546(.A1(new_n14425_), .A2(new_n14424_), .A3(new_n14023_), .ZN(new_n14842_));
  NOR3_X1    g14547(.A1(new_n14262_), .A2(new_n14842_), .A3(new_n14421_), .ZN(new_n14843_));
  NOR2_X1    g14548(.A1(new_n14843_), .A2(new_n14841_), .ZN(new_n14844_));
  OAI22_X1   g14549(.A1(new_n3989_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n4253_), .ZN(new_n14845_));
  OAI21_X1   g14550(.A1(new_n3717_), .A2(new_n3569_), .B(new_n14845_), .ZN(new_n14846_));
  AOI21_X1   g14551(.A1(new_n14846_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n14847_));
  XNOR2_X1   g14552(.A1(new_n4257_), .A2(new_n14847_), .ZN(new_n14848_));
  INV_X1     g14553(.I(new_n14848_), .ZN(new_n14849_));
  XOR2_X1    g14554(.A1(new_n14844_), .A2(new_n14849_), .Z(new_n14850_));
  AOI21_X1   g14555(.A1(new_n14837_), .A2(new_n14840_), .B(new_n14850_), .ZN(new_n14851_));
  AOI21_X1   g14556(.A1(new_n14838_), .A2(new_n14839_), .B(new_n14835_), .ZN(new_n14852_));
  NOR3_X1    g14557(.A1(new_n14828_), .A2(new_n14831_), .A3(new_n14836_), .ZN(new_n14853_));
  XOR2_X1    g14558(.A1(new_n14844_), .A2(new_n14848_), .Z(new_n14854_));
  NOR3_X1    g14559(.A1(new_n14854_), .A2(new_n14853_), .A3(new_n14852_), .ZN(new_n14855_));
  NOR2_X1    g14560(.A1(new_n14851_), .A2(new_n14855_), .ZN(new_n14856_));
  NAND2_X1   g14561(.A1(new_n14258_), .A2(new_n14442_), .ZN(new_n14857_));
  NOR2_X1    g14562(.A1(new_n14259_), .A2(new_n14437_), .ZN(new_n14858_));
  OAI21_X1   g14563(.A1(new_n14258_), .A2(new_n14442_), .B(new_n14858_), .ZN(new_n14859_));
  NAND2_X1   g14564(.A1(new_n14859_), .A2(new_n14857_), .ZN(new_n14860_));
  OAI22_X1   g14565(.A1(new_n4774_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n5068_), .ZN(new_n14861_));
  OAI21_X1   g14566(.A1(new_n4500_), .A2(new_n2884_), .B(new_n14861_), .ZN(new_n14862_));
  AOI21_X1   g14567(.A1(new_n14862_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n14863_));
  XOR2_X1    g14568(.A1(new_n5067_), .A2(new_n14863_), .Z(new_n14864_));
  INV_X1     g14569(.I(new_n14864_), .ZN(new_n14865_));
  XOR2_X1    g14570(.A1(new_n14860_), .A2(new_n14865_), .Z(new_n14866_));
  NOR2_X1    g14571(.A1(new_n14860_), .A2(new_n14864_), .ZN(new_n14867_));
  INV_X1     g14572(.I(new_n14860_), .ZN(new_n14868_));
  NOR2_X1    g14573(.A1(new_n14868_), .A2(new_n14865_), .ZN(new_n14869_));
  OAI21_X1   g14574(.A1(new_n14869_), .A2(new_n14867_), .B(new_n14856_), .ZN(new_n14870_));
  OAI21_X1   g14575(.A1(new_n14856_), .A2(new_n14866_), .B(new_n14870_), .ZN(new_n14871_));
  INV_X1     g14576(.I(new_n14871_), .ZN(new_n14872_));
  NOR3_X1    g14577(.A1(new_n14690_), .A2(new_n14687_), .A3(new_n14872_), .ZN(new_n14873_));
  NAND2_X1   g14578(.A1(new_n14487_), .A2(new_n14483_), .ZN(new_n14874_));
  NAND2_X1   g14579(.A1(new_n14254_), .A2(new_n14874_), .ZN(new_n14875_));
  OAI21_X1   g14580(.A1(new_n14254_), .A2(new_n14874_), .B(new_n14688_), .ZN(new_n14876_));
  AOI21_X1   g14581(.A1(new_n14876_), .A2(new_n14875_), .B(new_n14871_), .ZN(new_n14877_));
  OAI21_X1   g14582(.A1(new_n14877_), .A2(new_n14873_), .B(new_n14686_), .ZN(new_n14878_));
  NAND3_X1   g14583(.A1(new_n14876_), .A2(new_n14875_), .A3(new_n14871_), .ZN(new_n14879_));
  OAI21_X1   g14584(.A1(new_n14690_), .A2(new_n14687_), .B(new_n14872_), .ZN(new_n14880_));
  NAND3_X1   g14585(.A1(new_n14880_), .A2(new_n14879_), .A3(new_n14685_), .ZN(new_n14881_));
  AOI21_X1   g14586(.A1(new_n14878_), .A2(new_n14881_), .B(new_n14678_), .ZN(new_n14882_));
  AOI21_X1   g14587(.A1(new_n14880_), .A2(new_n14879_), .B(new_n14685_), .ZN(new_n14883_));
  NOR3_X1    g14588(.A1(new_n14877_), .A2(new_n14873_), .A3(new_n14686_), .ZN(new_n14884_));
  NOR3_X1    g14589(.A1(new_n14883_), .A2(new_n14884_), .A3(new_n14677_), .ZN(new_n14885_));
  NOR2_X1    g14590(.A1(new_n14885_), .A2(new_n14882_), .ZN(new_n14886_));
  NOR2_X1    g14591(.A1(new_n14500_), .A2(new_n14501_), .ZN(new_n14887_));
  NOR2_X1    g14592(.A1(new_n14887_), .A2(new_n14105_), .ZN(new_n14888_));
  NAND2_X1   g14593(.A1(new_n14100_), .A2(new_n14498_), .ZN(new_n14889_));
  AOI21_X1   g14594(.A1(new_n14887_), .A2(new_n14105_), .B(new_n14889_), .ZN(new_n14890_));
  OAI22_X1   g14595(.A1(new_n1347_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n1344_), .ZN(new_n14891_));
  OAI21_X1   g14596(.A1(new_n7198_), .A2(new_n1457_), .B(new_n14891_), .ZN(new_n14892_));
  AOI21_X1   g14597(.A1(new_n14892_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n14893_));
  XNOR2_X1   g14598(.A1(new_n7874_), .A2(new_n14893_), .ZN(new_n14894_));
  NOR3_X1    g14599(.A1(new_n14890_), .A2(new_n14888_), .A3(new_n14894_), .ZN(new_n14895_));
  OAI21_X1   g14600(.A1(new_n14890_), .A2(new_n14888_), .B(new_n14894_), .ZN(new_n14896_));
  INV_X1     g14601(.I(new_n14896_), .ZN(new_n14897_));
  OAI21_X1   g14602(.A1(new_n14897_), .A2(new_n14895_), .B(new_n14886_), .ZN(new_n14898_));
  OAI21_X1   g14603(.A1(new_n14883_), .A2(new_n14884_), .B(new_n14677_), .ZN(new_n14899_));
  NAND3_X1   g14604(.A1(new_n14878_), .A2(new_n14881_), .A3(new_n14678_), .ZN(new_n14900_));
  NAND2_X1   g14605(.A1(new_n14899_), .A2(new_n14900_), .ZN(new_n14901_));
  INV_X1     g14606(.I(new_n14895_), .ZN(new_n14902_));
  NAND3_X1   g14607(.A1(new_n14902_), .A2(new_n14901_), .A3(new_n14896_), .ZN(new_n14903_));
  AOI21_X1   g14608(.A1(new_n14898_), .A2(new_n14903_), .B(new_n14673_), .ZN(new_n14904_));
  AOI21_X1   g14609(.A1(new_n14902_), .A2(new_n14896_), .B(new_n14901_), .ZN(new_n14905_));
  NOR3_X1    g14610(.A1(new_n14897_), .A2(new_n14886_), .A3(new_n14895_), .ZN(new_n14906_));
  NOR3_X1    g14611(.A1(new_n14905_), .A2(new_n14906_), .A3(new_n14672_), .ZN(new_n14907_));
  NOR2_X1    g14612(.A1(new_n14907_), .A2(new_n14904_), .ZN(new_n14908_));
  OAI22_X1   g14613(.A1(new_n1055_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n1061_), .ZN(new_n14909_));
  OAI21_X1   g14614(.A1(new_n8218_), .A2(new_n1332_), .B(new_n14909_), .ZN(new_n14910_));
  AOI21_X1   g14615(.A1(new_n14910_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n14911_));
  XOR2_X1    g14616(.A1(new_n8952_), .A2(new_n14911_), .Z(new_n14912_));
  NOR2_X1    g14617(.A1(new_n14908_), .A2(new_n14912_), .ZN(new_n14913_));
  OAI21_X1   g14618(.A1(new_n14905_), .A2(new_n14906_), .B(new_n14672_), .ZN(new_n14914_));
  NAND3_X1   g14619(.A1(new_n14898_), .A2(new_n14903_), .A3(new_n14673_), .ZN(new_n14915_));
  NAND2_X1   g14620(.A1(new_n14914_), .A2(new_n14915_), .ZN(new_n14916_));
  INV_X1     g14621(.I(new_n14912_), .ZN(new_n14917_));
  NOR2_X1    g14622(.A1(new_n14916_), .A2(new_n14917_), .ZN(new_n14918_));
  OAI21_X1   g14623(.A1(new_n14913_), .A2(new_n14918_), .B(new_n14668_), .ZN(new_n14919_));
  NOR2_X1    g14624(.A1(new_n14916_), .A2(new_n14912_), .ZN(new_n14920_));
  NOR2_X1    g14625(.A1(new_n14908_), .A2(new_n14917_), .ZN(new_n14921_));
  OAI21_X1   g14626(.A1(new_n14921_), .A2(new_n14920_), .B(new_n14667_), .ZN(new_n14922_));
  NAND2_X1   g14627(.A1(new_n14919_), .A2(new_n14922_), .ZN(new_n14923_));
  NAND2_X1   g14628(.A1(new_n14923_), .A2(new_n14666_), .ZN(new_n14924_));
  OAI21_X1   g14629(.A1(new_n14663_), .A2(new_n14664_), .B(new_n14661_), .ZN(new_n14925_));
  NAND2_X1   g14630(.A1(new_n14916_), .A2(new_n14917_), .ZN(new_n14926_));
  NAND2_X1   g14631(.A1(new_n14908_), .A2(new_n14912_), .ZN(new_n14927_));
  AOI21_X1   g14632(.A1(new_n14927_), .A2(new_n14926_), .B(new_n14667_), .ZN(new_n14928_));
  NAND2_X1   g14633(.A1(new_n14908_), .A2(new_n14917_), .ZN(new_n14929_));
  NAND2_X1   g14634(.A1(new_n14916_), .A2(new_n14912_), .ZN(new_n14930_));
  AOI21_X1   g14635(.A1(new_n14929_), .A2(new_n14930_), .B(new_n14668_), .ZN(new_n14931_));
  NOR2_X1    g14636(.A1(new_n14928_), .A2(new_n14931_), .ZN(new_n14932_));
  NAND2_X1   g14637(.A1(new_n14932_), .A2(new_n14925_), .ZN(new_n14933_));
  NAND2_X1   g14638(.A1(new_n14924_), .A2(new_n14933_), .ZN(new_n14934_));
  OAI22_X1   g14639(.A1(new_n970_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n820_), .ZN(new_n14935_));
  OAI21_X1   g14640(.A1(new_n9295_), .A2(new_n894_), .B(new_n14935_), .ZN(new_n14936_));
  AOI21_X1   g14641(.A1(new_n14936_), .A2(new_n827_), .B(new_n970_), .ZN(new_n14937_));
  XNOR2_X1   g14642(.A1(new_n10035_), .A2(new_n14937_), .ZN(new_n14938_));
  INV_X1     g14643(.I(new_n14938_), .ZN(new_n14939_));
  NAND2_X1   g14644(.A1(new_n14934_), .A2(new_n14939_), .ZN(new_n14940_));
  NAND3_X1   g14645(.A1(new_n14924_), .A2(new_n14933_), .A3(new_n14938_), .ZN(new_n14941_));
  AOI21_X1   g14646(.A1(new_n14940_), .A2(new_n14941_), .B(new_n14659_), .ZN(new_n14942_));
  NAND3_X1   g14647(.A1(new_n14924_), .A2(new_n14933_), .A3(new_n14939_), .ZN(new_n14943_));
  NOR2_X1    g14648(.A1(new_n14932_), .A2(new_n14925_), .ZN(new_n14944_));
  NOR2_X1    g14649(.A1(new_n14923_), .A2(new_n14666_), .ZN(new_n14945_));
  OAI21_X1   g14650(.A1(new_n14945_), .A2(new_n14944_), .B(new_n14938_), .ZN(new_n14946_));
  NAND2_X1   g14651(.A1(new_n14946_), .A2(new_n14943_), .ZN(new_n14947_));
  NAND2_X1   g14652(.A1(new_n14947_), .A2(new_n14659_), .ZN(new_n14948_));
  INV_X1     g14653(.I(new_n14948_), .ZN(new_n14949_));
  OAI22_X1   g14654(.A1(new_n607_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n610_), .ZN(new_n14950_));
  OAI21_X1   g14655(.A1(new_n10477_), .A2(new_n684_), .B(new_n14950_), .ZN(new_n14951_));
  AOI21_X1   g14656(.A1(new_n14951_), .A2(new_n612_), .B(new_n607_), .ZN(new_n14952_));
  XOR2_X1    g14657(.A1(new_n11298_), .A2(new_n14952_), .Z(new_n14953_));
  INV_X1     g14658(.I(new_n14953_), .ZN(new_n14954_));
  OAI21_X1   g14659(.A1(new_n14949_), .A2(new_n14942_), .B(new_n14954_), .ZN(new_n14955_));
  INV_X1     g14660(.I(new_n14659_), .ZN(new_n14956_));
  NAND2_X1   g14661(.A1(new_n14940_), .A2(new_n14941_), .ZN(new_n14957_));
  NAND2_X1   g14662(.A1(new_n14957_), .A2(new_n14956_), .ZN(new_n14958_));
  NAND3_X1   g14663(.A1(new_n14958_), .A2(new_n14948_), .A3(new_n14953_), .ZN(new_n14959_));
  NAND2_X1   g14664(.A1(new_n14955_), .A2(new_n14959_), .ZN(new_n14960_));
  OAI22_X1   g14665(.A1(new_n448_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n450_), .ZN(new_n14961_));
  OAI21_X1   g14666(.A1(new_n11744_), .A2(new_n496_), .B(new_n14961_), .ZN(new_n14962_));
  AOI21_X1   g14667(.A1(new_n14962_), .A2(new_n452_), .B(new_n448_), .ZN(new_n14963_));
  XNOR2_X1   g14668(.A1(new_n12546_), .A2(new_n14963_), .ZN(new_n14964_));
  NOR2_X1    g14669(.A1(new_n14960_), .A2(new_n14964_), .ZN(new_n14965_));
  AOI21_X1   g14670(.A1(new_n14958_), .A2(new_n14948_), .B(new_n14953_), .ZN(new_n14966_));
  NOR3_X1    g14671(.A1(new_n14949_), .A2(new_n14942_), .A3(new_n14954_), .ZN(new_n14967_));
  NOR2_X1    g14672(.A1(new_n14967_), .A2(new_n14966_), .ZN(new_n14968_));
  INV_X1     g14673(.I(new_n14964_), .ZN(new_n14969_));
  NOR2_X1    g14674(.A1(new_n14968_), .A2(new_n14969_), .ZN(new_n14970_));
  OAI21_X1   g14675(.A1(new_n14970_), .A2(new_n14965_), .B(new_n14655_), .ZN(new_n14971_));
  INV_X1     g14676(.I(new_n14655_), .ZN(new_n14972_));
  NOR2_X1    g14677(.A1(new_n14968_), .A2(new_n14964_), .ZN(new_n14973_));
  NOR2_X1    g14678(.A1(new_n14960_), .A2(new_n14969_), .ZN(new_n14974_));
  OAI21_X1   g14679(.A1(new_n14973_), .A2(new_n14974_), .B(new_n14972_), .ZN(new_n14975_));
  INV_X1     g14680(.I(new_n14593_), .ZN(new_n14976_));
  NAND2_X1   g14681(.A1(new_n14591_), .A2(new_n14594_), .ZN(new_n14977_));
  OAI21_X1   g14682(.A1(new_n14591_), .A2(new_n14976_), .B(new_n14977_), .ZN(new_n14978_));
  AOI21_X1   g14683(.A1(\b[62] ), .A2(\b[63] ), .B(\a[2] ), .ZN(new_n14979_));
  NOR2_X1    g14684(.A1(new_n426_), .A2(new_n14979_), .ZN(new_n14980_));
  XOR2_X1    g14685(.A1(new_n14978_), .A2(new_n14980_), .Z(new_n14981_));
  INV_X1     g14686(.I(new_n14981_), .ZN(new_n14982_));
  NAND3_X1   g14687(.A1(new_n14971_), .A2(new_n14975_), .A3(new_n14982_), .ZN(new_n14983_));
  NAND2_X1   g14688(.A1(new_n14968_), .A2(new_n14969_), .ZN(new_n14984_));
  NAND2_X1   g14689(.A1(new_n14960_), .A2(new_n14964_), .ZN(new_n14985_));
  AOI21_X1   g14690(.A1(new_n14984_), .A2(new_n14985_), .B(new_n14972_), .ZN(new_n14986_));
  NAND2_X1   g14691(.A1(new_n14960_), .A2(new_n14969_), .ZN(new_n14987_));
  NAND2_X1   g14692(.A1(new_n14968_), .A2(new_n14964_), .ZN(new_n14988_));
  AOI21_X1   g14693(.A1(new_n14988_), .A2(new_n14987_), .B(new_n14655_), .ZN(new_n14989_));
  OAI21_X1   g14694(.A1(new_n14986_), .A2(new_n14989_), .B(new_n14981_), .ZN(new_n14990_));
  AOI21_X1   g14695(.A1(new_n14990_), .A2(new_n14983_), .B(new_n14654_), .ZN(new_n14991_));
  INV_X1     g14696(.I(new_n14654_), .ZN(new_n14992_));
  NOR3_X1    g14697(.A1(new_n14986_), .A2(new_n14989_), .A3(new_n14981_), .ZN(new_n14993_));
  AOI21_X1   g14698(.A1(new_n14971_), .A2(new_n14975_), .B(new_n14982_), .ZN(new_n14994_));
  NOR3_X1    g14699(.A1(new_n14992_), .A2(new_n14994_), .A3(new_n14993_), .ZN(new_n14995_));
  OAI21_X1   g14700(.A1(new_n14995_), .A2(new_n14991_), .B(new_n14650_), .ZN(new_n14996_));
  INV_X1     g14701(.I(new_n14650_), .ZN(new_n14997_));
  OAI21_X1   g14702(.A1(new_n14993_), .A2(new_n14994_), .B(new_n14992_), .ZN(new_n14998_));
  NAND3_X1   g14703(.A1(new_n14990_), .A2(new_n14983_), .A3(new_n14654_), .ZN(new_n14999_));
  NAND3_X1   g14704(.A1(new_n14998_), .A2(new_n14997_), .A3(new_n14999_), .ZN(new_n15000_));
  NAND2_X1   g14705(.A1(new_n15000_), .A2(new_n14996_), .ZN(new_n15001_));
  NOR2_X1    g14706(.A1(new_n14616_), .A2(new_n14604_), .ZN(new_n15002_));
  INV_X1     g14707(.I(new_n15002_), .ZN(new_n15003_));
  NOR2_X1    g14708(.A1(new_n14609_), .A2(new_n14612_), .ZN(new_n15004_));
  XOR2_X1    g14709(.A1(new_n15004_), .A2(new_n14241_), .Z(new_n15005_));
  OAI21_X1   g14710(.A1(new_n14244_), .A2(new_n14605_), .B(new_n15005_), .ZN(new_n15006_));
  NAND2_X1   g14711(.A1(new_n15006_), .A2(new_n15003_), .ZN(new_n15007_));
  NAND2_X1   g14712(.A1(new_n15001_), .A2(new_n15007_), .ZN(new_n15008_));
  XOR2_X1    g14713(.A1(new_n14646_), .A2(new_n15008_), .Z(new_n15009_));
  XOR2_X1    g14714(.A1(new_n15009_), .A2(new_n14632_), .Z(\f[64] ));
  OAI21_X1   g14715(.A1(new_n14629_), .A2(new_n14628_), .B(new_n14631_), .ZN(new_n15011_));
  NAND3_X1   g14716(.A1(new_n14620_), .A2(new_n14624_), .A3(new_n14626_), .ZN(new_n15012_));
  NAND3_X1   g14717(.A1(new_n14233_), .A2(new_n15011_), .A3(new_n15012_), .ZN(new_n15013_));
  AOI21_X1   g14718(.A1(new_n15011_), .A2(new_n15012_), .B(new_n14233_), .ZN(new_n15014_));
  OAI21_X1   g14719(.A1(new_n15014_), .A2(new_n13822_), .B(new_n15013_), .ZN(new_n15015_));
  AOI21_X1   g14720(.A1(new_n13819_), .A2(new_n13817_), .B(new_n15015_), .ZN(new_n15016_));
  AOI21_X1   g14721(.A1(new_n14998_), .A2(new_n14999_), .B(new_n14997_), .ZN(new_n15017_));
  NOR3_X1    g14722(.A1(new_n14995_), .A2(new_n14991_), .A3(new_n14650_), .ZN(new_n15018_));
  NOR2_X1    g14723(.A1(new_n15017_), .A2(new_n15018_), .ZN(new_n15019_));
  NOR2_X1    g14724(.A1(new_n15019_), .A2(new_n15012_), .ZN(new_n15020_));
  AOI22_X1   g14725(.A1(new_n15019_), .A2(new_n15012_), .B1(new_n15003_), .B2(new_n15006_), .ZN(new_n15021_));
  AOI21_X1   g14726(.A1(new_n15016_), .A2(new_n15021_), .B(new_n15020_), .ZN(new_n15022_));
  OAI22_X1   g14727(.A1(new_n13785_), .A2(new_n341_), .B1(new_n404_), .B2(new_n14208_), .ZN(new_n15023_));
  OAI21_X1   g14728(.A1(new_n13367_), .A2(new_n366_), .B(new_n15023_), .ZN(new_n15024_));
  AOI21_X1   g14729(.A1(new_n15024_), .A2(new_n334_), .B(new_n341_), .ZN(new_n15025_));
  XOR2_X1    g14730(.A1(new_n14213_), .A2(new_n15025_), .Z(new_n15026_));
  NOR2_X1    g14731(.A1(new_n14650_), .A2(new_n14964_), .ZN(new_n15027_));
  NOR2_X1    g14732(.A1(new_n14997_), .A2(new_n14969_), .ZN(new_n15028_));
  NAND2_X1   g14733(.A1(new_n14960_), .A2(new_n14972_), .ZN(new_n15029_));
  NAND2_X1   g14734(.A1(new_n14968_), .A2(new_n14655_), .ZN(new_n15030_));
  AOI21_X1   g14735(.A1(new_n15030_), .A2(new_n15029_), .B(new_n15028_), .ZN(new_n15031_));
  NOR2_X1    g14736(.A1(new_n15031_), .A2(new_n15027_), .ZN(new_n15032_));
  INV_X1     g14737(.I(new_n15032_), .ZN(new_n15033_));
  NAND3_X1   g14738(.A1(new_n14958_), .A2(new_n14948_), .A3(new_n14954_), .ZN(new_n15034_));
  OAI21_X1   g14739(.A1(new_n14949_), .A2(new_n14942_), .B(new_n14953_), .ZN(new_n15035_));
  NAND2_X1   g14740(.A1(new_n15035_), .A2(new_n14655_), .ZN(new_n15036_));
  NAND2_X1   g14741(.A1(new_n15036_), .A2(new_n15034_), .ZN(new_n15037_));
  INV_X1     g14742(.I(new_n15037_), .ZN(new_n15038_));
  INV_X1     g14743(.I(new_n14940_), .ZN(new_n15039_));
  XOR2_X1    g14744(.A1(new_n14916_), .A2(new_n14668_), .Z(new_n15040_));
  NAND2_X1   g14745(.A1(new_n15040_), .A2(new_n14912_), .ZN(new_n15041_));
  OAI21_X1   g14746(.A1(new_n14923_), .A2(new_n14925_), .B(new_n15041_), .ZN(new_n15042_));
  NOR2_X1    g14747(.A1(new_n14890_), .A2(new_n14888_), .ZN(new_n15043_));
  NAND2_X1   g14748(.A1(new_n14901_), .A2(new_n15043_), .ZN(new_n15044_));
  INV_X1     g14749(.I(new_n15044_), .ZN(new_n15045_));
  NOR2_X1    g14750(.A1(new_n14901_), .A2(new_n15043_), .ZN(new_n15046_));
  OAI21_X1   g14751(.A1(new_n15045_), .A2(new_n15046_), .B(new_n14672_), .ZN(new_n15047_));
  INV_X1     g14752(.I(new_n15046_), .ZN(new_n15048_));
  NAND3_X1   g14753(.A1(new_n15048_), .A2(new_n14673_), .A3(new_n15044_), .ZN(new_n15049_));
  AOI21_X1   g14754(.A1(new_n15047_), .A2(new_n15049_), .B(new_n14894_), .ZN(new_n15050_));
  INV_X1     g14755(.I(new_n15050_), .ZN(new_n15051_));
  NOR2_X1    g14756(.A1(new_n14886_), .A2(new_n14672_), .ZN(new_n15052_));
  OAI22_X1   g14757(.A1(new_n2171_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n2166_), .ZN(new_n15053_));
  OAI21_X1   g14758(.A1(new_n5913_), .A2(new_n2322_), .B(new_n15053_), .ZN(new_n15054_));
  AOI21_X1   g14759(.A1(new_n15054_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n15055_));
  XOR2_X1    g14760(.A1(new_n6233_), .A2(new_n15055_), .Z(new_n15056_));
  INV_X1     g14761(.I(new_n15056_), .ZN(new_n15057_));
  NOR2_X1    g14762(.A1(new_n14828_), .A2(new_n14831_), .ZN(new_n15058_));
  NAND2_X1   g14763(.A1(new_n15058_), .A2(new_n14836_), .ZN(new_n15059_));
  INV_X1     g14764(.I(new_n14844_), .ZN(new_n15060_));
  OAI21_X1   g14765(.A1(new_n15058_), .A2(new_n14836_), .B(new_n15060_), .ZN(new_n15061_));
  NAND2_X1   g14766(.A1(new_n15061_), .A2(new_n15059_), .ZN(new_n15062_));
  INV_X1     g14767(.I(new_n15062_), .ZN(new_n15063_));
  NAND2_X1   g14768(.A1(new_n14706_), .A2(new_n14695_), .ZN(new_n15064_));
  INV_X1     g14769(.I(new_n15064_), .ZN(new_n15065_));
  NOR2_X1    g14770(.A1(new_n14706_), .A2(new_n14695_), .ZN(new_n15066_));
  XNOR2_X1   g14771(.A1(new_n14820_), .A2(new_n14700_), .ZN(new_n15067_));
  NOR2_X1    g14772(.A1(new_n15066_), .A2(new_n15067_), .ZN(new_n15068_));
  NOR2_X1    g14773(.A1(new_n15068_), .A2(new_n15065_), .ZN(new_n15069_));
  INV_X1     g14774(.I(new_n15069_), .ZN(new_n15070_));
  NOR2_X1    g14775(.A1(new_n14701_), .A2(new_n14814_), .ZN(new_n15071_));
  INV_X1     g14776(.I(new_n15071_), .ZN(new_n15072_));
  NAND2_X1   g14777(.A1(new_n14701_), .A2(new_n14814_), .ZN(new_n15073_));
  XOR2_X1    g14778(.A1(new_n14810_), .A2(new_n14708_), .Z(new_n15074_));
  NAND2_X1   g14779(.A1(new_n15073_), .A2(new_n15074_), .ZN(new_n15075_));
  NAND2_X1   g14780(.A1(new_n15075_), .A2(new_n15072_), .ZN(new_n15076_));
  OAI22_X1   g14781(.A1(new_n6644_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n6647_), .ZN(new_n15077_));
  OAI21_X1   g14782(.A1(new_n1634_), .A2(new_n7284_), .B(new_n15077_), .ZN(new_n15078_));
  AOI21_X1   g14783(.A1(new_n15078_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n15079_));
  XNOR2_X1   g14784(.A1(new_n1940_), .A2(new_n15079_), .ZN(new_n15080_));
  NAND3_X1   g14785(.A1(new_n14792_), .A2(new_n14793_), .A3(new_n14790_), .ZN(new_n15081_));
  OAI21_X1   g14786(.A1(new_n14782_), .A2(new_n14785_), .B(new_n14789_), .ZN(new_n15082_));
  NAND2_X1   g14787(.A1(new_n15082_), .A2(new_n14799_), .ZN(new_n15083_));
  NAND2_X1   g14788(.A1(new_n15083_), .A2(new_n15081_), .ZN(new_n15084_));
  NOR2_X1    g14789(.A1(new_n14708_), .A2(new_n14803_), .ZN(new_n15085_));
  NAND3_X1   g14790(.A1(new_n14791_), .A2(new_n14794_), .A3(new_n14799_), .ZN(new_n15086_));
  INV_X1     g14791(.I(new_n14799_), .ZN(new_n15087_));
  NAND2_X1   g14792(.A1(new_n14806_), .A2(new_n15087_), .ZN(new_n15088_));
  AOI22_X1   g14793(.A1(new_n15086_), .A2(new_n15088_), .B1(new_n14708_), .B2(new_n14803_), .ZN(new_n15089_));
  NOR2_X1    g14794(.A1(new_n15089_), .A2(new_n15085_), .ZN(new_n15090_));
  NAND2_X1   g14795(.A1(new_n14725_), .A2(new_n14714_), .ZN(new_n15091_));
  XOR2_X1    g14796(.A1(new_n14775_), .A2(new_n14719_), .Z(new_n15092_));
  OAI21_X1   g14797(.A1(new_n14725_), .A2(new_n14714_), .B(new_n15092_), .ZN(new_n15093_));
  NAND2_X1   g14798(.A1(new_n15093_), .A2(new_n15091_), .ZN(new_n15094_));
  INV_X1     g14799(.I(new_n14771_), .ZN(new_n15095_));
  NOR2_X1    g14800(.A1(new_n15095_), .A2(new_n14774_), .ZN(new_n15096_));
  NAND2_X1   g14801(.A1(new_n15095_), .A2(new_n14774_), .ZN(new_n15097_));
  AOI21_X1   g14802(.A1(new_n14718_), .A2(new_n15097_), .B(new_n15096_), .ZN(new_n15098_));
  INV_X1     g14803(.I(new_n14767_), .ZN(new_n15099_));
  AOI21_X1   g14804(.A1(new_n14765_), .A2(new_n14769_), .B(new_n15099_), .ZN(new_n15100_));
  INV_X1     g14805(.I(new_n14757_), .ZN(new_n15101_));
  OAI21_X1   g14806(.A1(new_n14729_), .A2(new_n15101_), .B(new_n14756_), .ZN(new_n15102_));
  AOI21_X1   g14807(.A1(new_n14731_), .A2(new_n14746_), .B(new_n14744_), .ZN(new_n15103_));
  AOI22_X1   g14808(.A1(new_n13472_), .A2(new_n413_), .B1(\b[3] ), .B2(new_n13884_), .ZN(new_n15104_));
  OAI21_X1   g14809(.A1(new_n15104_), .A2(\a[62] ), .B(new_n13466_), .ZN(new_n15105_));
  XOR2_X1    g14810(.A1(new_n15105_), .A2(new_n378_), .Z(new_n15106_));
  NOR2_X1    g14811(.A1(new_n13476_), .A2(new_n269_), .ZN(new_n15107_));
  XOR2_X1    g14812(.A1(new_n14736_), .A2(new_n269_), .Z(new_n15108_));
  NAND2_X1   g14813(.A1(new_n15108_), .A2(\b[2] ), .ZN(new_n15109_));
  XOR2_X1    g14814(.A1(new_n15109_), .A2(new_n15107_), .Z(new_n15110_));
  XNOR2_X1   g14815(.A1(new_n15106_), .A2(new_n15110_), .ZN(new_n15111_));
  NOR2_X1    g14816(.A1(new_n15106_), .A2(new_n15110_), .ZN(new_n15112_));
  NAND2_X1   g14817(.A1(new_n15106_), .A2(new_n15110_), .ZN(new_n15113_));
  INV_X1     g14818(.I(new_n15113_), .ZN(new_n15114_));
  OAI21_X1   g14819(.A1(new_n15112_), .A2(new_n15114_), .B(new_n15103_), .ZN(new_n15115_));
  OAI21_X1   g14820(.A1(new_n15103_), .A2(new_n15111_), .B(new_n15115_), .ZN(new_n15116_));
  AOI22_X1   g14821(.A1(new_n13078_), .A2(\b[6] ), .B1(new_n517_), .B2(new_n12218_), .ZN(new_n15117_));
  OAI21_X1   g14822(.A1(new_n15117_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n15118_));
  XOR2_X1    g14823(.A1(new_n522_), .A2(new_n15118_), .Z(new_n15119_));
  NOR2_X1    g14824(.A1(new_n15116_), .A2(new_n15119_), .ZN(new_n15120_));
  NAND2_X1   g14825(.A1(new_n15116_), .A2(new_n15119_), .ZN(new_n15121_));
  INV_X1     g14826(.I(new_n15121_), .ZN(new_n15122_));
  OAI21_X1   g14827(.A1(new_n15120_), .A2(new_n15122_), .B(new_n15102_), .ZN(new_n15123_));
  XOR2_X1    g14828(.A1(new_n15116_), .A2(new_n15119_), .Z(new_n15124_));
  INV_X1     g14829(.I(new_n15124_), .ZN(new_n15125_));
  OAI21_X1   g14830(.A1(new_n15102_), .A2(new_n15125_), .B(new_n15123_), .ZN(new_n15126_));
  AOI22_X1   g14831(.A1(new_n10969_), .A2(new_n773_), .B1(new_n11394_), .B2(\b[9] ), .ZN(new_n15127_));
  OAI21_X1   g14832(.A1(new_n15127_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n15128_));
  XOR2_X1    g14833(.A1(new_n710_), .A2(new_n15128_), .Z(new_n15129_));
  XOR2_X1    g14834(.A1(new_n15126_), .A2(new_n15129_), .Z(new_n15130_));
  OR2_X2     g14835(.A1(new_n15130_), .A2(new_n15100_), .Z(new_n15131_));
  INV_X1     g14836(.I(new_n15129_), .ZN(new_n15132_));
  AND2_X2    g14837(.A1(new_n15126_), .A2(new_n15132_), .Z(new_n15133_));
  NOR2_X1    g14838(.A1(new_n15126_), .A2(new_n15132_), .ZN(new_n15134_));
  OAI21_X1   g14839(.A1(new_n15133_), .A2(new_n15134_), .B(new_n15100_), .ZN(new_n15135_));
  AOI22_X1   g14840(.A1(new_n11415_), .A2(new_n932_), .B1(\b[12] ), .B2(new_n10145_), .ZN(new_n15136_));
  OAI21_X1   g14841(.A1(new_n15136_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n15137_));
  XOR2_X1    g14842(.A1(new_n937_), .A2(new_n15137_), .Z(new_n15138_));
  INV_X1     g14843(.I(new_n15138_), .ZN(new_n15139_));
  NAND3_X1   g14844(.A1(new_n15131_), .A2(new_n15135_), .A3(new_n15139_), .ZN(new_n15140_));
  INV_X1     g14845(.I(new_n15140_), .ZN(new_n15141_));
  AOI21_X1   g14846(.A1(new_n15131_), .A2(new_n15135_), .B(new_n15139_), .ZN(new_n15142_));
  NOR2_X1    g14847(.A1(new_n15141_), .A2(new_n15142_), .ZN(new_n15143_));
  NOR2_X1    g14848(.A1(new_n15143_), .A2(new_n15098_), .ZN(new_n15144_));
  INV_X1     g14849(.I(new_n15098_), .ZN(new_n15145_));
  NAND2_X1   g14850(.A1(new_n15131_), .A2(new_n15135_), .ZN(new_n15146_));
  XOR2_X1    g14851(.A1(new_n15146_), .A2(new_n15139_), .Z(new_n15147_));
  NOR2_X1    g14852(.A1(new_n15145_), .A2(new_n15147_), .ZN(new_n15148_));
  NOR2_X1    g14853(.A1(new_n15148_), .A2(new_n15144_), .ZN(new_n15149_));
  AOI22_X1   g14854(.A1(new_n8631_), .A2(\b[16] ), .B1(\b[17] ), .B2(new_n9382_), .ZN(new_n15150_));
  AOI21_X1   g14855(.A1(\b[15] ), .A2(new_n9731_), .B(new_n15150_), .ZN(new_n15151_));
  OAI21_X1   g14856(.A1(new_n15151_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n15152_));
  XOR2_X1    g14857(.A1(new_n1196_), .A2(new_n15152_), .Z(new_n15153_));
  XOR2_X1    g14858(.A1(new_n15149_), .A2(new_n15153_), .Z(new_n15154_));
  NAND2_X1   g14859(.A1(new_n15154_), .A2(new_n15094_), .ZN(new_n15155_));
  INV_X1     g14860(.I(new_n15153_), .ZN(new_n15156_));
  OAI21_X1   g14861(.A1(new_n15148_), .A2(new_n15144_), .B(new_n15156_), .ZN(new_n15157_));
  NAND2_X1   g14862(.A1(new_n15149_), .A2(new_n15153_), .ZN(new_n15158_));
  AND2_X2    g14863(.A1(new_n15158_), .A2(new_n15157_), .Z(new_n15159_));
  NOR2_X1    g14864(.A1(new_n15159_), .A2(new_n15094_), .ZN(new_n15160_));
  INV_X1     g14865(.I(new_n15160_), .ZN(new_n15161_));
  OAI22_X1   g14866(.A1(new_n7619_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n8309_), .ZN(new_n15162_));
  OAI21_X1   g14867(.A1(new_n1294_), .A2(new_n7947_), .B(new_n15162_), .ZN(new_n15163_));
  AOI21_X1   g14868(.A1(new_n15163_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n15164_));
  XOR2_X1    g14869(.A1(new_n1530_), .A2(new_n15164_), .Z(new_n15165_));
  INV_X1     g14870(.I(new_n15165_), .ZN(new_n15166_));
  NAND3_X1   g14871(.A1(new_n15161_), .A2(new_n15155_), .A3(new_n15166_), .ZN(new_n15167_));
  INV_X1     g14872(.I(new_n15155_), .ZN(new_n15168_));
  OAI21_X1   g14873(.A1(new_n15168_), .A2(new_n15160_), .B(new_n15165_), .ZN(new_n15169_));
  NAND2_X1   g14874(.A1(new_n15167_), .A2(new_n15169_), .ZN(new_n15170_));
  NAND2_X1   g14875(.A1(new_n15090_), .A2(new_n15170_), .ZN(new_n15171_));
  INV_X1     g14876(.I(new_n15170_), .ZN(new_n15172_));
  OAI21_X1   g14877(.A1(new_n15089_), .A2(new_n15085_), .B(new_n15172_), .ZN(new_n15173_));
  AOI21_X1   g14878(.A1(new_n15171_), .A2(new_n15173_), .B(new_n15084_), .ZN(new_n15174_));
  NAND3_X1   g14879(.A1(new_n15171_), .A2(new_n15173_), .A3(new_n15084_), .ZN(new_n15175_));
  INV_X1     g14880(.I(new_n15175_), .ZN(new_n15176_));
  OAI21_X1   g14881(.A1(new_n15176_), .A2(new_n15174_), .B(new_n15080_), .ZN(new_n15177_));
  INV_X1     g14882(.I(new_n15080_), .ZN(new_n15178_));
  INV_X1     g14883(.I(new_n15174_), .ZN(new_n15179_));
  NAND3_X1   g14884(.A1(new_n15179_), .A2(new_n15175_), .A3(new_n15178_), .ZN(new_n15180_));
  OAI22_X1   g14885(.A1(new_n5993_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n5991_), .ZN(new_n15181_));
  OAI21_X1   g14886(.A1(new_n2102_), .A2(new_n5997_), .B(new_n15181_), .ZN(new_n15182_));
  AOI21_X1   g14887(.A1(new_n15182_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n15183_));
  XNOR2_X1   g14888(.A1(new_n2443_), .A2(new_n15183_), .ZN(new_n15184_));
  AOI21_X1   g14889(.A1(new_n15180_), .A2(new_n15177_), .B(new_n15184_), .ZN(new_n15185_));
  NAND3_X1   g14890(.A1(new_n15180_), .A2(new_n15177_), .A3(new_n15184_), .ZN(new_n15186_));
  INV_X1     g14891(.I(new_n15186_), .ZN(new_n15187_));
  OAI21_X1   g14892(.A1(new_n15187_), .A2(new_n15185_), .B(new_n15076_), .ZN(new_n15188_));
  INV_X1     g14893(.I(new_n15076_), .ZN(new_n15189_));
  INV_X1     g14894(.I(new_n15184_), .ZN(new_n15190_));
  NAND3_X1   g14895(.A1(new_n15180_), .A2(new_n15177_), .A3(new_n15190_), .ZN(new_n15191_));
  INV_X1     g14896(.I(new_n15191_), .ZN(new_n15192_));
  AOI21_X1   g14897(.A1(new_n15180_), .A2(new_n15177_), .B(new_n15190_), .ZN(new_n15193_));
  OAI21_X1   g14898(.A1(new_n15192_), .A2(new_n15193_), .B(new_n15189_), .ZN(new_n15194_));
  OAI22_X1   g14899(.A1(new_n5420_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n5107_), .ZN(new_n15195_));
  OAI21_X1   g14900(.A1(new_n2643_), .A2(new_n5112_), .B(new_n15195_), .ZN(new_n15196_));
  AOI21_X1   g14901(.A1(new_n15196_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n15197_));
  XNOR2_X1   g14902(.A1(new_n3022_), .A2(new_n15197_), .ZN(new_n15198_));
  AOI21_X1   g14903(.A1(new_n15194_), .A2(new_n15188_), .B(new_n15198_), .ZN(new_n15199_));
  NAND3_X1   g14904(.A1(new_n15194_), .A2(new_n15188_), .A3(new_n15198_), .ZN(new_n15200_));
  INV_X1     g14905(.I(new_n15200_), .ZN(new_n15201_));
  OAI21_X1   g14906(.A1(new_n15201_), .A2(new_n15199_), .B(new_n15070_), .ZN(new_n15202_));
  INV_X1     g14907(.I(new_n15198_), .ZN(new_n15203_));
  NAND3_X1   g14908(.A1(new_n15194_), .A2(new_n15188_), .A3(new_n15203_), .ZN(new_n15204_));
  NAND2_X1   g14909(.A1(new_n15180_), .A2(new_n15177_), .ZN(new_n15205_));
  NAND2_X1   g14910(.A1(new_n15205_), .A2(new_n15190_), .ZN(new_n15206_));
  AOI22_X1   g14911(.A1(new_n15206_), .A2(new_n15186_), .B1(new_n15072_), .B2(new_n15075_), .ZN(new_n15207_));
  INV_X1     g14912(.I(new_n15193_), .ZN(new_n15208_));
  AOI21_X1   g14913(.A1(new_n15208_), .A2(new_n15191_), .B(new_n15076_), .ZN(new_n15209_));
  OAI21_X1   g14914(.A1(new_n15207_), .A2(new_n15209_), .B(new_n15198_), .ZN(new_n15210_));
  NAND2_X1   g14915(.A1(new_n15204_), .A2(new_n15210_), .ZN(new_n15211_));
  NAND2_X1   g14916(.A1(new_n15211_), .A2(new_n15069_), .ZN(new_n15212_));
  OAI22_X1   g14917(.A1(new_n4072_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n4067_), .ZN(new_n15213_));
  OAI21_X1   g14918(.A1(new_n3260_), .A2(new_n4318_), .B(new_n15213_), .ZN(new_n15214_));
  AOI21_X1   g14919(.A1(new_n15214_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n15215_));
  XOR2_X1    g14920(.A1(new_n3722_), .A2(new_n15215_), .Z(new_n15216_));
  INV_X1     g14921(.I(new_n15216_), .ZN(new_n15217_));
  NAND3_X1   g14922(.A1(new_n15212_), .A2(new_n15202_), .A3(new_n15217_), .ZN(new_n15218_));
  INV_X1     g14923(.I(new_n15199_), .ZN(new_n15219_));
  AOI21_X1   g14924(.A1(new_n15219_), .A2(new_n15200_), .B(new_n15069_), .ZN(new_n15220_));
  AOI21_X1   g14925(.A1(new_n15204_), .A2(new_n15210_), .B(new_n15070_), .ZN(new_n15221_));
  OAI21_X1   g14926(.A1(new_n15220_), .A2(new_n15221_), .B(new_n15216_), .ZN(new_n15222_));
  AOI22_X1   g14927(.A1(new_n15218_), .A2(new_n15222_), .B1(new_n15061_), .B2(new_n15059_), .ZN(new_n15223_));
  OAI21_X1   g14928(.A1(new_n15220_), .A2(new_n15221_), .B(new_n15217_), .ZN(new_n15224_));
  NAND3_X1   g14929(.A1(new_n15212_), .A2(new_n15202_), .A3(new_n15216_), .ZN(new_n15225_));
  NAND2_X1   g14930(.A1(new_n15224_), .A2(new_n15225_), .ZN(new_n15226_));
  AOI21_X1   g14931(.A1(new_n15063_), .A2(new_n15226_), .B(new_n15223_), .ZN(new_n15227_));
  NAND2_X1   g14932(.A1(new_n14860_), .A2(new_n14849_), .ZN(new_n15228_));
  INV_X1     g14933(.I(new_n15228_), .ZN(new_n15229_));
  NAND3_X1   g14934(.A1(new_n14837_), .A2(new_n14840_), .A3(new_n15060_), .ZN(new_n15230_));
  OAI21_X1   g14935(.A1(new_n14853_), .A2(new_n14852_), .B(new_n14844_), .ZN(new_n15231_));
  AOI22_X1   g14936(.A1(new_n14868_), .A2(new_n14848_), .B1(new_n15230_), .B2(new_n15231_), .ZN(new_n15232_));
  NOR2_X1    g14937(.A1(new_n15232_), .A2(new_n15229_), .ZN(new_n15233_));
  OAI22_X1   g14938(.A1(new_n4253_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n4500_), .ZN(new_n15234_));
  OAI21_X1   g14939(.A1(new_n3989_), .A2(new_n3569_), .B(new_n15234_), .ZN(new_n15235_));
  AOI21_X1   g14940(.A1(new_n15235_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n15236_));
  XOR2_X1    g14941(.A1(new_n4499_), .A2(new_n15236_), .Z(new_n15237_));
  INV_X1     g14942(.I(new_n15237_), .ZN(new_n15238_));
  NAND2_X1   g14943(.A1(new_n15233_), .A2(new_n15238_), .ZN(new_n15239_));
  NAND2_X1   g14944(.A1(new_n15231_), .A2(new_n15230_), .ZN(new_n15240_));
  OAI21_X1   g14945(.A1(new_n14849_), .A2(new_n14860_), .B(new_n15240_), .ZN(new_n15241_));
  NAND2_X1   g14946(.A1(new_n15241_), .A2(new_n15228_), .ZN(new_n15242_));
  NAND2_X1   g14947(.A1(new_n15242_), .A2(new_n15237_), .ZN(new_n15243_));
  AOI21_X1   g14948(.A1(new_n15243_), .A2(new_n15239_), .B(new_n15227_), .ZN(new_n15244_));
  INV_X1     g14949(.I(new_n15223_), .ZN(new_n15245_));
  NAND3_X1   g14950(.A1(new_n15226_), .A2(new_n15059_), .A3(new_n15061_), .ZN(new_n15246_));
  NAND2_X1   g14951(.A1(new_n15245_), .A2(new_n15246_), .ZN(new_n15247_));
  NAND2_X1   g14952(.A1(new_n15242_), .A2(new_n15238_), .ZN(new_n15248_));
  NAND2_X1   g14953(.A1(new_n15233_), .A2(new_n15237_), .ZN(new_n15249_));
  AOI21_X1   g14954(.A1(new_n15248_), .A2(new_n15249_), .B(new_n15247_), .ZN(new_n15250_));
  OAI22_X1   g14955(.A1(new_n5068_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n5353_), .ZN(new_n15251_));
  OAI21_X1   g14956(.A1(new_n4774_), .A2(new_n2884_), .B(new_n15251_), .ZN(new_n15252_));
  AOI21_X1   g14957(.A1(new_n15252_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n15253_));
  XNOR2_X1   g14958(.A1(new_n5357_), .A2(new_n15253_), .ZN(new_n15254_));
  NOR3_X1    g14959(.A1(new_n15244_), .A2(new_n15250_), .A3(new_n15254_), .ZN(new_n15255_));
  NOR2_X1    g14960(.A1(new_n15242_), .A2(new_n15237_), .ZN(new_n15256_));
  NOR2_X1    g14961(.A1(new_n15233_), .A2(new_n15238_), .ZN(new_n15257_));
  OAI21_X1   g14962(.A1(new_n15256_), .A2(new_n15257_), .B(new_n15247_), .ZN(new_n15258_));
  NOR2_X1    g14963(.A1(new_n15233_), .A2(new_n15237_), .ZN(new_n15259_));
  NOR2_X1    g14964(.A1(new_n15242_), .A2(new_n15238_), .ZN(new_n15260_));
  OAI21_X1   g14965(.A1(new_n15260_), .A2(new_n15259_), .B(new_n15227_), .ZN(new_n15261_));
  INV_X1     g14966(.I(new_n15254_), .ZN(new_n15262_));
  AOI21_X1   g14967(.A1(new_n15258_), .A2(new_n15261_), .B(new_n15262_), .ZN(new_n15263_));
  NOR2_X1    g14968(.A1(new_n15263_), .A2(new_n15255_), .ZN(new_n15264_));
  NAND2_X1   g14969(.A1(new_n14685_), .A2(new_n14865_), .ZN(new_n15265_));
  NOR2_X1    g14970(.A1(new_n14685_), .A2(new_n14865_), .ZN(new_n15266_));
  XOR2_X1    g14971(.A1(new_n14856_), .A2(new_n14860_), .Z(new_n15267_));
  OAI21_X1   g14972(.A1(new_n15266_), .A2(new_n15267_), .B(new_n15265_), .ZN(new_n15268_));
  XOR2_X1    g14973(.A1(new_n15264_), .A2(new_n15268_), .Z(new_n15269_));
  OAI21_X1   g14974(.A1(new_n14690_), .A2(new_n14687_), .B(new_n14678_), .ZN(new_n15270_));
  INV_X1     g14975(.I(new_n15270_), .ZN(new_n15271_));
  NOR2_X1    g14976(.A1(new_n14690_), .A2(new_n14687_), .ZN(new_n15272_));
  XNOR2_X1   g14977(.A1(new_n14685_), .A2(new_n14871_), .ZN(new_n15273_));
  AOI21_X1   g14978(.A1(new_n15272_), .A2(new_n14677_), .B(new_n15273_), .ZN(new_n15274_));
  OAI22_X1   g14979(.A1(new_n1712_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n1707_), .ZN(new_n15275_));
  OAI21_X1   g14980(.A1(new_n6538_), .A2(new_n1850_), .B(new_n15275_), .ZN(new_n15276_));
  AOI21_X1   g14981(.A1(new_n15276_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n15277_));
  XNOR2_X1   g14982(.A1(new_n7202_), .A2(new_n15277_), .ZN(new_n15278_));
  NOR3_X1    g14983(.A1(new_n15274_), .A2(new_n15271_), .A3(new_n15278_), .ZN(new_n15279_));
  NAND3_X1   g14984(.A1(new_n14876_), .A2(new_n14875_), .A3(new_n14677_), .ZN(new_n15280_));
  XOR2_X1    g14985(.A1(new_n14685_), .A2(new_n14871_), .Z(new_n15281_));
  NAND2_X1   g14986(.A1(new_n15280_), .A2(new_n15281_), .ZN(new_n15282_));
  INV_X1     g14987(.I(new_n15278_), .ZN(new_n15283_));
  AOI21_X1   g14988(.A1(new_n15282_), .A2(new_n15270_), .B(new_n15283_), .ZN(new_n15284_));
  OAI21_X1   g14989(.A1(new_n15279_), .A2(new_n15284_), .B(new_n15269_), .ZN(new_n15285_));
  NAND2_X1   g14990(.A1(new_n15264_), .A2(new_n15268_), .ZN(new_n15286_));
  NAND3_X1   g14991(.A1(new_n15258_), .A2(new_n15261_), .A3(new_n15262_), .ZN(new_n15287_));
  OAI21_X1   g14992(.A1(new_n15244_), .A2(new_n15250_), .B(new_n15254_), .ZN(new_n15288_));
  NAND2_X1   g14993(.A1(new_n15288_), .A2(new_n15287_), .ZN(new_n15289_));
  INV_X1     g14994(.I(new_n15268_), .ZN(new_n15290_));
  NAND2_X1   g14995(.A1(new_n15290_), .A2(new_n15289_), .ZN(new_n15291_));
  NAND2_X1   g14996(.A1(new_n15291_), .A2(new_n15286_), .ZN(new_n15292_));
  NAND3_X1   g14997(.A1(new_n15282_), .A2(new_n15270_), .A3(new_n15283_), .ZN(new_n15293_));
  OAI21_X1   g14998(.A1(new_n15274_), .A2(new_n15271_), .B(new_n15278_), .ZN(new_n15294_));
  NAND3_X1   g14999(.A1(new_n15294_), .A2(new_n15293_), .A3(new_n15292_), .ZN(new_n15295_));
  AOI21_X1   g15000(.A1(new_n15285_), .A2(new_n15295_), .B(new_n15057_), .ZN(new_n15296_));
  AOI21_X1   g15001(.A1(new_n15294_), .A2(new_n15293_), .B(new_n15292_), .ZN(new_n15297_));
  NOR3_X1    g15002(.A1(new_n15279_), .A2(new_n15284_), .A3(new_n15269_), .ZN(new_n15298_));
  NOR3_X1    g15003(.A1(new_n15298_), .A2(new_n15297_), .A3(new_n15056_), .ZN(new_n15299_));
  NOR2_X1    g15004(.A1(new_n15299_), .A2(new_n15296_), .ZN(new_n15300_));
  NAND3_X1   g15005(.A1(new_n14899_), .A2(new_n14900_), .A3(new_n14673_), .ZN(new_n15301_));
  INV_X1     g15006(.I(new_n15301_), .ZN(new_n15302_));
  AOI21_X1   g15007(.A1(new_n14899_), .A2(new_n14900_), .B(new_n14673_), .ZN(new_n15303_));
  NOR2_X1    g15008(.A1(new_n15302_), .A2(new_n15303_), .ZN(new_n15304_));
  NOR3_X1    g15009(.A1(new_n15300_), .A2(new_n15052_), .A3(new_n15304_), .ZN(new_n15305_));
  NOR2_X1    g15010(.A1(new_n14886_), .A2(new_n14672_), .ZN(new_n15307_));
  OAI21_X1   g15011(.A1(new_n15305_), .A2(new_n15307_), .B(new_n15043_), .ZN(new_n15308_));
  INV_X1     g15012(.I(new_n15043_), .ZN(new_n15309_));
  INV_X1     g15013(.I(new_n15052_), .ZN(new_n15310_));
  OAI21_X1   g15014(.A1(new_n15298_), .A2(new_n15297_), .B(new_n15056_), .ZN(new_n15311_));
  NAND3_X1   g15015(.A1(new_n15285_), .A2(new_n15295_), .A3(new_n15057_), .ZN(new_n15312_));
  NAND2_X1   g15016(.A1(new_n15311_), .A2(new_n15312_), .ZN(new_n15313_));
  OAI21_X1   g15017(.A1(new_n14885_), .A2(new_n14882_), .B(new_n14672_), .ZN(new_n15314_));
  NAND2_X1   g15018(.A1(new_n15314_), .A2(new_n15301_), .ZN(new_n15315_));
  NAND3_X1   g15019(.A1(new_n15313_), .A2(new_n15310_), .A3(new_n15315_), .ZN(new_n15316_));
  INV_X1     g15020(.I(new_n15307_), .ZN(new_n15317_));
  NAND3_X1   g15021(.A1(new_n15316_), .A2(new_n15309_), .A3(new_n15317_), .ZN(new_n15318_));
  OAI22_X1   g15022(.A1(new_n1347_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n1344_), .ZN(new_n15319_));
  OAI21_X1   g15023(.A1(new_n7864_), .A2(new_n1457_), .B(new_n15319_), .ZN(new_n15320_));
  AOI21_X1   g15024(.A1(new_n15320_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n15321_));
  XOR2_X1    g15025(.A1(new_n8217_), .A2(new_n15321_), .Z(new_n15322_));
  INV_X1     g15026(.I(new_n15322_), .ZN(new_n15323_));
  NAND3_X1   g15027(.A1(new_n15308_), .A2(new_n15318_), .A3(new_n15323_), .ZN(new_n15324_));
  AOI21_X1   g15028(.A1(new_n15316_), .A2(new_n15317_), .B(new_n15309_), .ZN(new_n15325_));
  NOR3_X1    g15029(.A1(new_n15305_), .A2(new_n15043_), .A3(new_n15307_), .ZN(new_n15326_));
  OAI21_X1   g15030(.A1(new_n15326_), .A2(new_n15325_), .B(new_n15322_), .ZN(new_n15327_));
  NAND3_X1   g15031(.A1(new_n15327_), .A2(new_n15324_), .A3(new_n15051_), .ZN(new_n15328_));
  NAND3_X1   g15032(.A1(new_n15328_), .A2(new_n14667_), .A3(new_n14916_), .ZN(new_n15329_));
  NOR3_X1    g15033(.A1(new_n15326_), .A2(new_n15325_), .A3(new_n15322_), .ZN(new_n15330_));
  AOI21_X1   g15034(.A1(new_n15308_), .A2(new_n15318_), .B(new_n15323_), .ZN(new_n15331_));
  NOR3_X1    g15035(.A1(new_n15330_), .A2(new_n15331_), .A3(new_n15050_), .ZN(new_n15332_));
  OAI21_X1   g15036(.A1(new_n15332_), .A2(new_n14908_), .B(new_n14668_), .ZN(new_n15333_));
  OAI22_X1   g15037(.A1(new_n1055_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n1061_), .ZN(new_n15334_));
  OAI21_X1   g15038(.A1(new_n8563_), .A2(new_n1332_), .B(new_n15334_), .ZN(new_n15335_));
  AOI21_X1   g15039(.A1(new_n15335_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n15336_));
  XNOR2_X1   g15040(.A1(new_n9299_), .A2(new_n15336_), .ZN(new_n15337_));
  INV_X1     g15041(.I(new_n15337_), .ZN(new_n15338_));
  NAND3_X1   g15042(.A1(new_n15333_), .A2(new_n15329_), .A3(new_n15338_), .ZN(new_n15339_));
  NOR3_X1    g15043(.A1(new_n15332_), .A2(new_n14668_), .A3(new_n14908_), .ZN(new_n15340_));
  AOI21_X1   g15044(.A1(new_n15328_), .A2(new_n14916_), .B(new_n14667_), .ZN(new_n15341_));
  OAI21_X1   g15045(.A1(new_n15340_), .A2(new_n15341_), .B(new_n15337_), .ZN(new_n15342_));
  AOI21_X1   g15046(.A1(new_n15342_), .A2(new_n15339_), .B(new_n15042_), .ZN(new_n15343_));
  AOI22_X1   g15047(.A1(new_n14932_), .A2(new_n14666_), .B1(new_n14912_), .B2(new_n15040_), .ZN(new_n15344_));
  OAI21_X1   g15048(.A1(new_n15340_), .A2(new_n15341_), .B(new_n15338_), .ZN(new_n15345_));
  NAND3_X1   g15049(.A1(new_n15333_), .A2(new_n15329_), .A3(new_n15337_), .ZN(new_n15346_));
  AOI21_X1   g15050(.A1(new_n15345_), .A2(new_n15346_), .B(new_n15344_), .ZN(new_n15347_));
  OAI22_X1   g15051(.A1(new_n970_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n820_), .ZN(new_n15348_));
  OAI21_X1   g15052(.A1(new_n10025_), .A2(new_n894_), .B(new_n15348_), .ZN(new_n15349_));
  AOI21_X1   g15053(.A1(new_n15349_), .A2(new_n827_), .B(new_n970_), .ZN(new_n15350_));
  XOR2_X1    g15054(.A1(new_n10476_), .A2(new_n15350_), .Z(new_n15351_));
  NOR3_X1    g15055(.A1(new_n15343_), .A2(new_n15347_), .A3(new_n15351_), .ZN(new_n15352_));
  NOR3_X1    g15056(.A1(new_n15340_), .A2(new_n15341_), .A3(new_n15337_), .ZN(new_n15353_));
  AOI21_X1   g15057(.A1(new_n15333_), .A2(new_n15329_), .B(new_n15338_), .ZN(new_n15354_));
  OAI21_X1   g15058(.A1(new_n15353_), .A2(new_n15354_), .B(new_n15344_), .ZN(new_n15355_));
  AOI21_X1   g15059(.A1(new_n15333_), .A2(new_n15329_), .B(new_n15337_), .ZN(new_n15356_));
  NOR3_X1    g15060(.A1(new_n15340_), .A2(new_n15341_), .A3(new_n15338_), .ZN(new_n15357_));
  OAI21_X1   g15061(.A1(new_n15357_), .A2(new_n15356_), .B(new_n15042_), .ZN(new_n15358_));
  INV_X1     g15062(.I(new_n15351_), .ZN(new_n15359_));
  AOI21_X1   g15063(.A1(new_n15358_), .A2(new_n15355_), .B(new_n15359_), .ZN(new_n15360_));
  OAI21_X1   g15064(.A1(new_n15360_), .A2(new_n15352_), .B(new_n14947_), .ZN(new_n15361_));
  NOR2_X1    g15065(.A1(new_n15361_), .A2(new_n15039_), .ZN(new_n15362_));
  NAND3_X1   g15066(.A1(new_n15358_), .A2(new_n15355_), .A3(new_n15359_), .ZN(new_n15363_));
  OAI21_X1   g15067(.A1(new_n15343_), .A2(new_n15347_), .B(new_n15351_), .ZN(new_n15364_));
  NAND2_X1   g15068(.A1(new_n15363_), .A2(new_n15364_), .ZN(new_n15365_));
  NAND2_X1   g15069(.A1(new_n14934_), .A2(new_n14939_), .ZN(new_n15367_));
  INV_X1     g15070(.I(new_n15367_), .ZN(new_n15368_));
  OAI21_X1   g15071(.A1(new_n15362_), .A2(new_n15368_), .B(new_n14659_), .ZN(new_n15369_));
  NAND3_X1   g15072(.A1(new_n15365_), .A2(new_n14940_), .A3(new_n14947_), .ZN(new_n15370_));
  NAND3_X1   g15073(.A1(new_n15370_), .A2(new_n14956_), .A3(new_n15367_), .ZN(new_n15371_));
  OAI22_X1   g15074(.A1(new_n448_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n450_), .ZN(new_n15372_));
  OAI21_X1   g15075(.A1(new_n12536_), .A2(new_n496_), .B(new_n15372_), .ZN(new_n15373_));
  AOI21_X1   g15076(.A1(new_n15373_), .A2(new_n452_), .B(new_n448_), .ZN(new_n15374_));
  XOR2_X1    g15077(.A1(new_n12969_), .A2(new_n15374_), .Z(new_n15375_));
  OAI22_X1   g15078(.A1(new_n607_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n610_), .ZN(new_n15376_));
  OAI21_X1   g15079(.A1(new_n10862_), .A2(new_n684_), .B(new_n15376_), .ZN(new_n15377_));
  AOI21_X1   g15080(.A1(new_n15377_), .A2(new_n612_), .B(new_n607_), .ZN(new_n15378_));
  XNOR2_X1   g15081(.A1(new_n11748_), .A2(new_n15378_), .ZN(new_n15379_));
  INV_X1     g15082(.I(new_n15379_), .ZN(new_n15380_));
  XOR2_X1    g15083(.A1(new_n15375_), .A2(new_n15380_), .Z(new_n15381_));
  AOI21_X1   g15084(.A1(new_n15369_), .A2(new_n15371_), .B(new_n15381_), .ZN(new_n15382_));
  AOI21_X1   g15085(.A1(new_n15370_), .A2(new_n15367_), .B(new_n14956_), .ZN(new_n15383_));
  NOR3_X1    g15086(.A1(new_n15362_), .A2(new_n14659_), .A3(new_n15368_), .ZN(new_n15384_));
  NOR2_X1    g15087(.A1(new_n15375_), .A2(new_n15379_), .ZN(new_n15385_));
  NAND2_X1   g15088(.A1(new_n15375_), .A2(new_n15379_), .ZN(new_n15386_));
  INV_X1     g15089(.I(new_n15386_), .ZN(new_n15387_));
  NOR2_X1    g15090(.A1(new_n15387_), .A2(new_n15385_), .ZN(new_n15388_));
  NOR3_X1    g15091(.A1(new_n15384_), .A2(new_n15383_), .A3(new_n15388_), .ZN(new_n15389_));
  OAI21_X1   g15092(.A1(new_n15389_), .A2(new_n15382_), .B(new_n15038_), .ZN(new_n15390_));
  INV_X1     g15093(.I(new_n15381_), .ZN(new_n15391_));
  OAI21_X1   g15094(.A1(new_n15384_), .A2(new_n15383_), .B(new_n15391_), .ZN(new_n15392_));
  INV_X1     g15095(.I(new_n15388_), .ZN(new_n15393_));
  NAND3_X1   g15096(.A1(new_n15369_), .A2(new_n15371_), .A3(new_n15393_), .ZN(new_n15394_));
  NAND3_X1   g15097(.A1(new_n15392_), .A2(new_n15394_), .A3(new_n15037_), .ZN(new_n15395_));
  NOR3_X1    g15098(.A1(new_n426_), .A2(new_n14592_), .A3(new_n289_), .ZN(new_n15396_));
  NOR2_X1    g15099(.A1(new_n14591_), .A2(\b[62] ), .ZN(new_n15397_));
  NOR2_X1    g15100(.A1(new_n15397_), .A2(new_n14592_), .ZN(new_n15398_));
  OAI21_X1   g15101(.A1(new_n15398_), .A2(new_n15396_), .B(new_n260_), .ZN(new_n15399_));
  XOR2_X1    g15102(.A1(new_n15399_), .A2(new_n15396_), .Z(new_n15400_));
  INV_X1     g15103(.I(new_n15400_), .ZN(new_n15401_));
  NAND3_X1   g15104(.A1(new_n15390_), .A2(new_n15395_), .A3(new_n15401_), .ZN(new_n15402_));
  AOI21_X1   g15105(.A1(new_n15392_), .A2(new_n15394_), .B(new_n15037_), .ZN(new_n15403_));
  NOR3_X1    g15106(.A1(new_n15389_), .A2(new_n15382_), .A3(new_n15038_), .ZN(new_n15404_));
  OAI21_X1   g15107(.A1(new_n15404_), .A2(new_n15403_), .B(new_n15400_), .ZN(new_n15405_));
  AOI21_X1   g15108(.A1(new_n15405_), .A2(new_n15402_), .B(new_n15033_), .ZN(new_n15406_));
  NOR3_X1    g15109(.A1(new_n15404_), .A2(new_n15403_), .A3(new_n15400_), .ZN(new_n15407_));
  AOI21_X1   g15110(.A1(new_n15390_), .A2(new_n15395_), .B(new_n15401_), .ZN(new_n15408_));
  NOR3_X1    g15111(.A1(new_n15407_), .A2(new_n15408_), .A3(new_n15032_), .ZN(new_n15409_));
  OAI21_X1   g15112(.A1(new_n15409_), .A2(new_n15406_), .B(new_n15026_), .ZN(new_n15410_));
  OR3_X2     g15113(.A1(new_n15409_), .A2(new_n15406_), .A3(new_n15026_), .Z(new_n15411_));
  NAND2_X1   g15114(.A1(new_n15411_), .A2(new_n15410_), .ZN(new_n15412_));
  NOR2_X1    g15115(.A1(new_n14992_), .A2(new_n14981_), .ZN(new_n15413_));
  NAND2_X1   g15116(.A1(new_n14992_), .A2(new_n14981_), .ZN(new_n15414_));
  NOR2_X1    g15117(.A1(new_n14986_), .A2(new_n14989_), .ZN(new_n15415_));
  XOR2_X1    g15118(.A1(new_n15415_), .A2(new_n14650_), .Z(new_n15416_));
  AOI21_X1   g15119(.A1(new_n15416_), .A2(new_n15414_), .B(new_n15413_), .ZN(new_n15417_));
  XOR2_X1    g15120(.A1(new_n15412_), .A2(new_n15417_), .Z(new_n15418_));
  INV_X1     g15121(.I(new_n15417_), .ZN(new_n15419_));
  NAND2_X1   g15122(.A1(new_n15412_), .A2(new_n15419_), .ZN(new_n15420_));
  INV_X1     g15123(.I(new_n15412_), .ZN(new_n15421_));
  NAND2_X1   g15124(.A1(new_n15421_), .A2(new_n15417_), .ZN(new_n15422_));
  NAND2_X1   g15125(.A1(new_n15422_), .A2(new_n15420_), .ZN(new_n15423_));
  NAND2_X1   g15126(.A1(new_n15423_), .A2(new_n15022_), .ZN(new_n15424_));
  OAI21_X1   g15127(.A1(new_n15022_), .A2(new_n15418_), .B(new_n15424_), .ZN(\f[65] ));
  AOI21_X1   g15128(.A1(new_n15392_), .A2(new_n15394_), .B(new_n15026_), .ZN(new_n15426_));
  INV_X1     g15129(.I(new_n15026_), .ZN(new_n15427_));
  NOR3_X1    g15130(.A1(new_n15389_), .A2(new_n15382_), .A3(new_n15427_), .ZN(new_n15428_));
  NOR2_X1    g15131(.A1(new_n15428_), .A2(new_n15038_), .ZN(new_n15429_));
  OAI22_X1   g15132(.A1(new_n14208_), .A2(new_n341_), .B1(new_n404_), .B2(new_n14592_), .ZN(new_n15430_));
  OAI21_X1   g15133(.A1(new_n13785_), .A2(new_n366_), .B(new_n15430_), .ZN(new_n15431_));
  AOI21_X1   g15134(.A1(new_n15431_), .A2(new_n334_), .B(new_n341_), .ZN(new_n15432_));
  XNOR2_X1   g15135(.A1(new_n14599_), .A2(new_n15432_), .ZN(new_n15433_));
  INV_X1     g15136(.I(new_n15433_), .ZN(new_n15434_));
  OAI21_X1   g15137(.A1(new_n15429_), .A2(new_n15426_), .B(new_n15434_), .ZN(new_n15435_));
  INV_X1     g15138(.I(new_n15426_), .ZN(new_n15436_));
  NAND3_X1   g15139(.A1(new_n15392_), .A2(new_n15394_), .A3(new_n15026_), .ZN(new_n15437_));
  NAND2_X1   g15140(.A1(new_n15437_), .A2(new_n15037_), .ZN(new_n15438_));
  NAND3_X1   g15141(.A1(new_n15438_), .A2(new_n15436_), .A3(new_n15433_), .ZN(new_n15439_));
  NAND2_X1   g15142(.A1(new_n15435_), .A2(new_n15439_), .ZN(new_n15440_));
  NOR2_X1    g15143(.A1(new_n15032_), .A2(new_n15400_), .ZN(new_n15441_));
  NOR3_X1    g15144(.A1(new_n15031_), .A2(new_n15027_), .A3(new_n15401_), .ZN(new_n15442_));
  NAND3_X1   g15145(.A1(new_n15390_), .A2(new_n15395_), .A3(new_n15427_), .ZN(new_n15443_));
  OAI21_X1   g15146(.A1(new_n15404_), .A2(new_n15403_), .B(new_n15026_), .ZN(new_n15444_));
  AOI21_X1   g15147(.A1(new_n15444_), .A2(new_n15443_), .B(new_n15442_), .ZN(new_n15445_));
  OAI21_X1   g15148(.A1(new_n15360_), .A2(new_n15352_), .B(new_n14934_), .ZN(new_n15446_));
  NAND2_X1   g15149(.A1(new_n15446_), .A2(new_n14938_), .ZN(new_n15447_));
  NOR3_X1    g15150(.A1(new_n15360_), .A2(new_n15352_), .A3(new_n14934_), .ZN(new_n15448_));
  NOR2_X1    g15151(.A1(new_n15448_), .A2(new_n14659_), .ZN(new_n15449_));
  AOI21_X1   g15152(.A1(new_n15327_), .A2(new_n15324_), .B(new_n15051_), .ZN(new_n15450_));
  OAI21_X1   g15153(.A1(new_n15450_), .A2(new_n14916_), .B(new_n14668_), .ZN(new_n15451_));
  NAND2_X1   g15154(.A1(new_n15282_), .A2(new_n15270_), .ZN(new_n15452_));
  XOR2_X1    g15155(.A1(new_n15452_), .A2(new_n15292_), .Z(new_n15453_));
  XOR2_X1    g15156(.A1(new_n15453_), .A2(new_n15057_), .Z(new_n15454_));
  NAND2_X1   g15157(.A1(new_n15454_), .A2(new_n15283_), .ZN(new_n15455_));
  OAI21_X1   g15158(.A1(new_n15300_), .A2(new_n14672_), .B(new_n14886_), .ZN(new_n15456_));
  AOI21_X1   g15159(.A1(new_n15300_), .A2(new_n14672_), .B(new_n15043_), .ZN(new_n15457_));
  INV_X1     g15160(.I(new_n15452_), .ZN(new_n15458_));
  XOR2_X1    g15161(.A1(new_n15292_), .A2(new_n15056_), .Z(new_n15459_));
  NAND2_X1   g15162(.A1(new_n15292_), .A2(new_n15056_), .ZN(new_n15460_));
  XOR2_X1    g15163(.A1(new_n15227_), .A2(new_n15237_), .Z(new_n15461_));
  NAND2_X1   g15164(.A1(new_n15227_), .A2(new_n15237_), .ZN(new_n15462_));
  INV_X1     g15165(.I(new_n15218_), .ZN(new_n15463_));
  NAND2_X1   g15166(.A1(new_n15212_), .A2(new_n15202_), .ZN(new_n15464_));
  AOI22_X1   g15167(.A1(new_n15061_), .A2(new_n15059_), .B1(new_n15464_), .B2(new_n15216_), .ZN(new_n15465_));
  NOR2_X1    g15168(.A1(new_n15465_), .A2(new_n15463_), .ZN(new_n15466_));
  INV_X1     g15169(.I(new_n15466_), .ZN(new_n15467_));
  INV_X1     g15170(.I(new_n15204_), .ZN(new_n15468_));
  NAND2_X1   g15171(.A1(new_n15194_), .A2(new_n15188_), .ZN(new_n15469_));
  AOI21_X1   g15172(.A1(new_n15469_), .A2(new_n15198_), .B(new_n15069_), .ZN(new_n15470_));
  AOI22_X1   g15173(.A1(new_n15205_), .A2(new_n15184_), .B1(new_n15075_), .B2(new_n15072_), .ZN(new_n15471_));
  NOR2_X1    g15174(.A1(new_n15471_), .A2(new_n15192_), .ZN(new_n15472_));
  NOR2_X1    g15175(.A1(new_n15090_), .A2(new_n15080_), .ZN(new_n15473_));
  NAND2_X1   g15176(.A1(new_n15090_), .A2(new_n15080_), .ZN(new_n15474_));
  XOR2_X1    g15177(.A1(new_n15170_), .A2(new_n15084_), .Z(new_n15475_));
  NAND2_X1   g15178(.A1(new_n15475_), .A2(new_n15474_), .ZN(new_n15476_));
  INV_X1     g15179(.I(new_n15476_), .ZN(new_n15477_));
  NAND2_X1   g15180(.A1(new_n15169_), .A2(new_n15084_), .ZN(new_n15478_));
  INV_X1     g15181(.I(new_n15157_), .ZN(new_n15479_));
  AOI22_X1   g15182(.A1(new_n15093_), .A2(new_n15091_), .B1(new_n15149_), .B2(new_n15153_), .ZN(new_n15480_));
  NOR2_X1    g15183(.A1(new_n15480_), .A2(new_n15479_), .ZN(new_n15481_));
  NOR2_X1    g15184(.A1(new_n15098_), .A2(new_n15142_), .ZN(new_n15482_));
  NOR2_X1    g15185(.A1(new_n15100_), .A2(new_n15134_), .ZN(new_n15483_));
  NOR2_X1    g15186(.A1(new_n15483_), .A2(new_n15133_), .ZN(new_n15484_));
  AOI21_X1   g15187(.A1(new_n15102_), .A2(new_n15121_), .B(new_n15120_), .ZN(new_n15485_));
  INV_X1     g15188(.I(new_n15112_), .ZN(new_n15486_));
  OAI21_X1   g15189(.A1(new_n15103_), .A2(new_n15114_), .B(new_n15486_), .ZN(new_n15487_));
  OAI22_X1   g15190(.A1(new_n13880_), .A2(new_n421_), .B1(new_n325_), .B2(new_n13885_), .ZN(new_n15488_));
  AOI21_X1   g15191(.A1(new_n15488_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n15489_));
  XOR2_X1    g15192(.A1(new_n556_), .A2(new_n15489_), .Z(new_n15490_));
  INV_X1     g15193(.I(new_n15490_), .ZN(new_n15491_));
  NOR2_X1    g15194(.A1(new_n13476_), .A2(new_n280_), .ZN(new_n15492_));
  XOR2_X1    g15195(.A1(new_n14736_), .A2(new_n280_), .Z(new_n15493_));
  NAND2_X1   g15196(.A1(new_n15493_), .A2(\b[3] ), .ZN(new_n15494_));
  XOR2_X1    g15197(.A1(new_n15494_), .A2(new_n15492_), .Z(new_n15495_));
  XOR2_X1    g15198(.A1(new_n15495_), .A2(new_n260_), .Z(new_n15496_));
  NOR2_X1    g15199(.A1(new_n15491_), .A2(new_n15496_), .ZN(new_n15497_));
  AND2_X2    g15200(.A1(new_n15495_), .A2(\a[2] ), .Z(new_n15498_));
  NOR2_X1    g15201(.A1(new_n15495_), .A2(\a[2] ), .ZN(new_n15499_));
  NOR2_X1    g15202(.A1(new_n15498_), .A2(new_n15499_), .ZN(new_n15500_));
  NOR2_X1    g15203(.A1(new_n15490_), .A2(new_n15500_), .ZN(new_n15501_));
  AOI22_X1   g15204(.A1(new_n13078_), .A2(\b[7] ), .B1(new_n650_), .B2(new_n12218_), .ZN(new_n15502_));
  OAI21_X1   g15205(.A1(new_n15502_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n15503_));
  XOR2_X1    g15206(.A1(new_n569_), .A2(new_n15503_), .Z(new_n15504_));
  NOR3_X1    g15207(.A1(new_n15504_), .A2(new_n15497_), .A3(new_n15501_), .ZN(new_n15505_));
  NOR2_X1    g15208(.A1(new_n15497_), .A2(new_n15501_), .ZN(new_n15506_));
  INV_X1     g15209(.I(new_n15504_), .ZN(new_n15507_));
  NOR2_X1    g15210(.A1(new_n15506_), .A2(new_n15507_), .ZN(new_n15508_));
  OAI21_X1   g15211(.A1(new_n15505_), .A2(new_n15508_), .B(new_n15487_), .ZN(new_n15509_));
  INV_X1     g15212(.I(new_n15487_), .ZN(new_n15510_));
  XOR2_X1    g15213(.A1(new_n15506_), .A2(new_n15507_), .Z(new_n15511_));
  NAND2_X1   g15214(.A1(new_n15510_), .A2(new_n15511_), .ZN(new_n15512_));
  NAND2_X1   g15215(.A1(new_n15512_), .A2(new_n15509_), .ZN(new_n15513_));
  AOI22_X1   g15216(.A1(new_n10969_), .A2(new_n14320_), .B1(new_n11394_), .B2(\b[10] ), .ZN(new_n15514_));
  OAI21_X1   g15217(.A1(new_n15514_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n15515_));
  XNOR2_X1   g15218(.A1(new_n785_), .A2(new_n15515_), .ZN(new_n15516_));
  XOR2_X1    g15219(.A1(new_n15513_), .A2(new_n15516_), .Z(new_n15517_));
  NOR2_X1    g15220(.A1(new_n15517_), .A2(new_n15485_), .ZN(new_n15518_));
  INV_X1     g15221(.I(new_n15518_), .ZN(new_n15519_));
  INV_X1     g15222(.I(new_n15513_), .ZN(new_n15520_));
  NOR2_X1    g15223(.A1(new_n15520_), .A2(new_n15516_), .ZN(new_n15521_));
  NAND2_X1   g15224(.A1(new_n15520_), .A2(new_n15516_), .ZN(new_n15522_));
  INV_X1     g15225(.I(new_n15522_), .ZN(new_n15523_));
  OAI21_X1   g15226(.A1(new_n15523_), .A2(new_n15521_), .B(new_n15485_), .ZN(new_n15524_));
  NAND2_X1   g15227(.A1(new_n15519_), .A2(new_n15524_), .ZN(new_n15525_));
  AOI22_X1   g15228(.A1(new_n11415_), .A2(new_n1105_), .B1(\b[13] ), .B2(new_n10145_), .ZN(new_n15526_));
  OAI21_X1   g15229(.A1(new_n15526_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n15527_));
  XNOR2_X1   g15230(.A1(new_n1024_), .A2(new_n15527_), .ZN(new_n15528_));
  NOR2_X1    g15231(.A1(new_n15525_), .A2(new_n15528_), .ZN(new_n15529_));
  INV_X1     g15232(.I(new_n15529_), .ZN(new_n15530_));
  NAND2_X1   g15233(.A1(new_n15525_), .A2(new_n15528_), .ZN(new_n15531_));
  AOI21_X1   g15234(.A1(new_n15530_), .A2(new_n15531_), .B(new_n15484_), .ZN(new_n15532_));
  AOI21_X1   g15235(.A1(new_n15519_), .A2(new_n15524_), .B(new_n15528_), .ZN(new_n15533_));
  NAND3_X1   g15236(.A1(new_n15519_), .A2(new_n15524_), .A3(new_n15528_), .ZN(new_n15534_));
  INV_X1     g15237(.I(new_n15534_), .ZN(new_n15535_));
  OAI21_X1   g15238(.A1(new_n15533_), .A2(new_n15535_), .B(new_n15484_), .ZN(new_n15536_));
  INV_X1     g15239(.I(new_n15536_), .ZN(new_n15537_));
  NOR2_X1    g15240(.A1(new_n15537_), .A2(new_n15532_), .ZN(new_n15538_));
  OAI22_X1   g15241(.A1(new_n8644_), .A2(new_n1189_), .B1(new_n1294_), .B2(new_n9388_), .ZN(new_n15539_));
  OAI21_X1   g15242(.A1(new_n1109_), .A2(new_n10154_), .B(new_n15539_), .ZN(new_n15540_));
  AOI21_X1   g15243(.A1(new_n15540_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n15541_));
  XOR2_X1    g15244(.A1(new_n1299_), .A2(new_n15541_), .Z(new_n15542_));
  NOR2_X1    g15245(.A1(new_n15538_), .A2(new_n15542_), .ZN(new_n15543_));
  INV_X1     g15246(.I(new_n15532_), .ZN(new_n15544_));
  NAND2_X1   g15247(.A1(new_n15544_), .A2(new_n15536_), .ZN(new_n15545_));
  INV_X1     g15248(.I(new_n15542_), .ZN(new_n15546_));
  NOR2_X1    g15249(.A1(new_n15545_), .A2(new_n15546_), .ZN(new_n15547_));
  OAI22_X1   g15250(.A1(new_n15543_), .A2(new_n15547_), .B1(new_n15141_), .B2(new_n15482_), .ZN(new_n15548_));
  NOR2_X1    g15251(.A1(new_n15482_), .A2(new_n15141_), .ZN(new_n15549_));
  NOR2_X1    g15252(.A1(new_n15545_), .A2(new_n15542_), .ZN(new_n15550_));
  NOR2_X1    g15253(.A1(new_n15538_), .A2(new_n15546_), .ZN(new_n15551_));
  OAI21_X1   g15254(.A1(new_n15550_), .A2(new_n15551_), .B(new_n15549_), .ZN(new_n15552_));
  OAI22_X1   g15255(.A1(new_n7619_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n8309_), .ZN(new_n15553_));
  OAI21_X1   g15256(.A1(new_n1518_), .A2(new_n7947_), .B(new_n15553_), .ZN(new_n15554_));
  AOI21_X1   g15257(.A1(new_n15554_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n15555_));
  XNOR2_X1   g15258(.A1(new_n1638_), .A2(new_n15555_), .ZN(new_n15556_));
  INV_X1     g15259(.I(new_n15556_), .ZN(new_n15557_));
  NAND3_X1   g15260(.A1(new_n15552_), .A2(new_n15548_), .A3(new_n15557_), .ZN(new_n15558_));
  NAND2_X1   g15261(.A1(new_n15552_), .A2(new_n15548_), .ZN(new_n15559_));
  NAND2_X1   g15262(.A1(new_n15559_), .A2(new_n15556_), .ZN(new_n15560_));
  AOI21_X1   g15263(.A1(new_n15558_), .A2(new_n15560_), .B(new_n15481_), .ZN(new_n15561_));
  INV_X1     g15264(.I(new_n15561_), .ZN(new_n15562_));
  AOI21_X1   g15265(.A1(new_n15552_), .A2(new_n15548_), .B(new_n15556_), .ZN(new_n15563_));
  NOR2_X1    g15266(.A1(new_n15559_), .A2(new_n15557_), .ZN(new_n15564_));
  OAI21_X1   g15267(.A1(new_n15563_), .A2(new_n15564_), .B(new_n15481_), .ZN(new_n15565_));
  OAI22_X1   g15268(.A1(new_n6644_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n6647_), .ZN(new_n15566_));
  OAI21_X1   g15269(.A1(new_n1803_), .A2(new_n7284_), .B(new_n15566_), .ZN(new_n15567_));
  AOI21_X1   g15270(.A1(new_n15567_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n15568_));
  XOR2_X1    g15271(.A1(new_n2106_), .A2(new_n15568_), .Z(new_n15569_));
  INV_X1     g15272(.I(new_n15569_), .ZN(new_n15570_));
  NAND3_X1   g15273(.A1(new_n15562_), .A2(new_n15565_), .A3(new_n15570_), .ZN(new_n15571_));
  INV_X1     g15274(.I(new_n15565_), .ZN(new_n15572_));
  OAI21_X1   g15275(.A1(new_n15572_), .A2(new_n15561_), .B(new_n15569_), .ZN(new_n15573_));
  AOI22_X1   g15276(.A1(new_n15478_), .A2(new_n15167_), .B1(new_n15571_), .B2(new_n15573_), .ZN(new_n15574_));
  INV_X1     g15277(.I(new_n15574_), .ZN(new_n15575_));
  OAI21_X1   g15278(.A1(new_n15572_), .A2(new_n15561_), .B(new_n15570_), .ZN(new_n15576_));
  NAND3_X1   g15279(.A1(new_n15562_), .A2(new_n15565_), .A3(new_n15569_), .ZN(new_n15577_));
  NAND2_X1   g15280(.A1(new_n15576_), .A2(new_n15577_), .ZN(new_n15578_));
  NAND3_X1   g15281(.A1(new_n15578_), .A2(new_n15478_), .A3(new_n15167_), .ZN(new_n15579_));
  OAI22_X1   g15282(.A1(new_n5993_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n5991_), .ZN(new_n15580_));
  OAI21_X1   g15283(.A1(new_n2281_), .A2(new_n5997_), .B(new_n15580_), .ZN(new_n15581_));
  AOI21_X1   g15284(.A1(new_n15581_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n15582_));
  XNOR2_X1   g15285(.A1(new_n2647_), .A2(new_n15582_), .ZN(new_n15583_));
  AOI21_X1   g15286(.A1(new_n15575_), .A2(new_n15579_), .B(new_n15583_), .ZN(new_n15584_));
  INV_X1     g15287(.I(new_n15579_), .ZN(new_n15585_));
  INV_X1     g15288(.I(new_n15583_), .ZN(new_n15586_));
  NOR3_X1    g15289(.A1(new_n15585_), .A2(new_n15574_), .A3(new_n15586_), .ZN(new_n15587_));
  OAI22_X1   g15290(.A1(new_n15477_), .A2(new_n15473_), .B1(new_n15584_), .B2(new_n15587_), .ZN(new_n15588_));
  INV_X1     g15291(.I(new_n15588_), .ZN(new_n15589_));
  NOR3_X1    g15292(.A1(new_n15585_), .A2(new_n15574_), .A3(new_n15583_), .ZN(new_n15590_));
  AOI21_X1   g15293(.A1(new_n15575_), .A2(new_n15579_), .B(new_n15586_), .ZN(new_n15591_));
  NOR2_X1    g15294(.A1(new_n15590_), .A2(new_n15591_), .ZN(new_n15592_));
  NOR3_X1    g15295(.A1(new_n15592_), .A2(new_n15473_), .A3(new_n15477_), .ZN(new_n15593_));
  OAI22_X1   g15296(.A1(new_n5420_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n5107_), .ZN(new_n15594_));
  OAI21_X1   g15297(.A1(new_n2842_), .A2(new_n5112_), .B(new_n15594_), .ZN(new_n15595_));
  AOI21_X1   g15298(.A1(new_n15595_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n15596_));
  XNOR2_X1   g15299(.A1(new_n3264_), .A2(new_n15596_), .ZN(new_n15597_));
  NOR3_X1    g15300(.A1(new_n15589_), .A2(new_n15593_), .A3(new_n15597_), .ZN(new_n15598_));
  INV_X1     g15301(.I(new_n15593_), .ZN(new_n15599_));
  INV_X1     g15302(.I(new_n15597_), .ZN(new_n15600_));
  AOI21_X1   g15303(.A1(new_n15599_), .A2(new_n15588_), .B(new_n15600_), .ZN(new_n15601_));
  NOR2_X1    g15304(.A1(new_n15601_), .A2(new_n15598_), .ZN(new_n15602_));
  NOR2_X1    g15305(.A1(new_n15472_), .A2(new_n15602_), .ZN(new_n15603_));
  AOI21_X1   g15306(.A1(new_n15599_), .A2(new_n15588_), .B(new_n15597_), .ZN(new_n15604_));
  NOR3_X1    g15307(.A1(new_n15589_), .A2(new_n15593_), .A3(new_n15600_), .ZN(new_n15605_));
  NOR2_X1    g15308(.A1(new_n15604_), .A2(new_n15605_), .ZN(new_n15606_));
  NOR3_X1    g15309(.A1(new_n15606_), .A2(new_n15192_), .A3(new_n15471_), .ZN(new_n15607_));
  OAI22_X1   g15310(.A1(new_n4072_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n4067_), .ZN(new_n15608_));
  OAI21_X1   g15311(.A1(new_n3709_), .A2(new_n4318_), .B(new_n15608_), .ZN(new_n15609_));
  AOI21_X1   g15312(.A1(new_n15609_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n15610_));
  XNOR2_X1   g15313(.A1(new_n3993_), .A2(new_n15610_), .ZN(new_n15611_));
  NOR3_X1    g15314(.A1(new_n15607_), .A2(new_n15603_), .A3(new_n15611_), .ZN(new_n15612_));
  OAI22_X1   g15315(.A1(new_n15471_), .A2(new_n15192_), .B1(new_n15601_), .B2(new_n15598_), .ZN(new_n15613_));
  OAI21_X1   g15316(.A1(new_n15589_), .A2(new_n15593_), .B(new_n15600_), .ZN(new_n15614_));
  NAND3_X1   g15317(.A1(new_n15599_), .A2(new_n15588_), .A3(new_n15597_), .ZN(new_n15615_));
  NAND2_X1   g15318(.A1(new_n15615_), .A2(new_n15614_), .ZN(new_n15616_));
  NAND2_X1   g15319(.A1(new_n15472_), .A2(new_n15616_), .ZN(new_n15617_));
  INV_X1     g15320(.I(new_n15611_), .ZN(new_n15618_));
  AOI21_X1   g15321(.A1(new_n15617_), .A2(new_n15613_), .B(new_n15618_), .ZN(new_n15619_));
  OAI22_X1   g15322(.A1(new_n15470_), .A2(new_n15468_), .B1(new_n15612_), .B2(new_n15619_), .ZN(new_n15620_));
  OAI21_X1   g15323(.A1(new_n15068_), .A2(new_n15065_), .B(new_n15210_), .ZN(new_n15621_));
  OAI21_X1   g15324(.A1(new_n15607_), .A2(new_n15603_), .B(new_n15618_), .ZN(new_n15622_));
  NAND3_X1   g15325(.A1(new_n15617_), .A2(new_n15613_), .A3(new_n15611_), .ZN(new_n15623_));
  NAND2_X1   g15326(.A1(new_n15622_), .A2(new_n15623_), .ZN(new_n15624_));
  NAND3_X1   g15327(.A1(new_n15624_), .A2(new_n15204_), .A3(new_n15621_), .ZN(new_n15625_));
  OAI22_X1   g15328(.A1(new_n4500_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n4774_), .ZN(new_n15626_));
  OAI21_X1   g15329(.A1(new_n4253_), .A2(new_n3569_), .B(new_n15626_), .ZN(new_n15627_));
  AOI21_X1   g15330(.A1(new_n15627_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n15628_));
  XNOR2_X1   g15331(.A1(new_n4778_), .A2(new_n15628_), .ZN(new_n15629_));
  AOI21_X1   g15332(.A1(new_n15625_), .A2(new_n15620_), .B(new_n15629_), .ZN(new_n15630_));
  NAND3_X1   g15333(.A1(new_n15617_), .A2(new_n15613_), .A3(new_n15618_), .ZN(new_n15631_));
  OAI21_X1   g15334(.A1(new_n15607_), .A2(new_n15603_), .B(new_n15611_), .ZN(new_n15632_));
  AOI22_X1   g15335(.A1(new_n15621_), .A2(new_n15204_), .B1(new_n15632_), .B2(new_n15631_), .ZN(new_n15633_));
  NAND2_X1   g15336(.A1(new_n15621_), .A2(new_n15204_), .ZN(new_n15634_));
  AOI21_X1   g15337(.A1(new_n15617_), .A2(new_n15613_), .B(new_n15611_), .ZN(new_n15635_));
  NOR3_X1    g15338(.A1(new_n15607_), .A2(new_n15603_), .A3(new_n15618_), .ZN(new_n15636_));
  NOR2_X1    g15339(.A1(new_n15636_), .A2(new_n15635_), .ZN(new_n15637_));
  NOR2_X1    g15340(.A1(new_n15634_), .A2(new_n15637_), .ZN(new_n15638_));
  INV_X1     g15341(.I(new_n15629_), .ZN(new_n15639_));
  NOR3_X1    g15342(.A1(new_n15638_), .A2(new_n15633_), .A3(new_n15639_), .ZN(new_n15640_));
  OAI22_X1   g15343(.A1(new_n15465_), .A2(new_n15463_), .B1(new_n15640_), .B2(new_n15630_), .ZN(new_n15641_));
  NOR3_X1    g15344(.A1(new_n15638_), .A2(new_n15633_), .A3(new_n15629_), .ZN(new_n15642_));
  AOI21_X1   g15345(.A1(new_n15625_), .A2(new_n15620_), .B(new_n15639_), .ZN(new_n15643_));
  NOR2_X1    g15346(.A1(new_n15642_), .A2(new_n15643_), .ZN(new_n15644_));
  OAI21_X1   g15347(.A1(new_n15467_), .A2(new_n15644_), .B(new_n15641_), .ZN(new_n15645_));
  OAI22_X1   g15348(.A1(new_n5913_), .A2(new_n2700_), .B1(new_n2705_), .B2(new_n5353_), .ZN(new_n15646_));
  OAI21_X1   g15349(.A1(new_n5068_), .A2(new_n2884_), .B(new_n15646_), .ZN(new_n15647_));
  AOI21_X1   g15350(.A1(new_n15647_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n15648_));
  XOR2_X1    g15351(.A1(new_n5600_), .A2(new_n15648_), .Z(new_n15649_));
  NAND3_X1   g15352(.A1(new_n15645_), .A2(new_n15462_), .A3(new_n15649_), .ZN(new_n15650_));
  NOR2_X1    g15353(.A1(new_n15247_), .A2(new_n15238_), .ZN(new_n15651_));
  NOR2_X1    g15354(.A1(new_n15640_), .A2(new_n15630_), .ZN(new_n15652_));
  NOR2_X1    g15355(.A1(new_n15466_), .A2(new_n15652_), .ZN(new_n15653_));
  NOR3_X1    g15356(.A1(new_n15644_), .A2(new_n15463_), .A3(new_n15465_), .ZN(new_n15654_));
  OAI21_X1   g15357(.A1(new_n15653_), .A2(new_n15654_), .B(new_n15649_), .ZN(new_n15655_));
  NAND2_X1   g15358(.A1(new_n15655_), .A2(new_n15651_), .ZN(new_n15656_));
  AOI22_X1   g15359(.A1(new_n15656_), .A2(new_n15650_), .B1(new_n15461_), .B2(new_n15233_), .ZN(new_n15657_));
  XOR2_X1    g15360(.A1(new_n15227_), .A2(new_n15238_), .Z(new_n15658_));
  NOR2_X1    g15361(.A1(new_n15655_), .A2(new_n15651_), .ZN(new_n15659_));
  AOI21_X1   g15362(.A1(new_n15645_), .A2(new_n15649_), .B(new_n15462_), .ZN(new_n15660_));
  NOR4_X1    g15363(.A1(new_n15659_), .A2(new_n15658_), .A3(new_n15660_), .A4(new_n15242_), .ZN(new_n15661_));
  OAI22_X1   g15364(.A1(new_n2171_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n2166_), .ZN(new_n15662_));
  OAI21_X1   g15365(.A1(new_n5921_), .A2(new_n2322_), .B(new_n15662_), .ZN(new_n15663_));
  AOI21_X1   g15366(.A1(new_n15663_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n15664_));
  XOR2_X1    g15367(.A1(new_n6543_), .A2(new_n15664_), .Z(new_n15665_));
  INV_X1     g15368(.I(new_n15665_), .ZN(new_n15666_));
  OAI21_X1   g15369(.A1(new_n15657_), .A2(new_n15661_), .B(new_n15666_), .ZN(new_n15667_));
  AOI21_X1   g15370(.A1(new_n15290_), .A2(new_n15264_), .B(new_n15667_), .ZN(new_n15668_));
  OAI22_X1   g15371(.A1(new_n15659_), .A2(new_n15660_), .B1(new_n15658_), .B2(new_n15242_), .ZN(new_n15669_));
  NAND4_X1   g15372(.A1(new_n15656_), .A2(new_n15461_), .A3(new_n15650_), .A4(new_n15233_), .ZN(new_n15670_));
  AOI21_X1   g15373(.A1(new_n15669_), .A2(new_n15670_), .B(new_n15665_), .ZN(new_n15671_));
  NOR3_X1    g15374(.A1(new_n15671_), .A2(new_n15289_), .A3(new_n15268_), .ZN(new_n15672_));
  OAI21_X1   g15375(.A1(new_n15668_), .A2(new_n15672_), .B(new_n15288_), .ZN(new_n15673_));
  OAI21_X1   g15376(.A1(new_n15289_), .A2(new_n15268_), .B(new_n15671_), .ZN(new_n15674_));
  NAND3_X1   g15377(.A1(new_n15290_), .A2(new_n15667_), .A3(new_n15264_), .ZN(new_n15675_));
  NAND3_X1   g15378(.A1(new_n15674_), .A2(new_n15675_), .A3(new_n15263_), .ZN(new_n15676_));
  NAND2_X1   g15379(.A1(new_n15673_), .A2(new_n15676_), .ZN(new_n15677_));
  OAI22_X1   g15380(.A1(new_n1712_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n1707_), .ZN(new_n15678_));
  OAI21_X1   g15381(.A1(new_n6847_), .A2(new_n1850_), .B(new_n15678_), .ZN(new_n15679_));
  AOI21_X1   g15382(.A1(new_n15679_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n15680_));
  XOR2_X1    g15383(.A1(new_n7516_), .A2(new_n15680_), .Z(new_n15681_));
  INV_X1     g15384(.I(new_n15681_), .ZN(new_n15682_));
  NAND3_X1   g15385(.A1(new_n15677_), .A2(new_n15460_), .A3(new_n15682_), .ZN(new_n15683_));
  INV_X1     g15386(.I(new_n15460_), .ZN(new_n15684_));
  AOI21_X1   g15387(.A1(new_n15674_), .A2(new_n15675_), .B(new_n15263_), .ZN(new_n15685_));
  NOR3_X1    g15388(.A1(new_n15668_), .A2(new_n15672_), .A3(new_n15288_), .ZN(new_n15686_));
  OAI21_X1   g15389(.A1(new_n15686_), .A2(new_n15685_), .B(new_n15682_), .ZN(new_n15687_));
  NAND2_X1   g15390(.A1(new_n15687_), .A2(new_n15684_), .ZN(new_n15688_));
  AOI22_X1   g15391(.A1(new_n15688_), .A2(new_n15683_), .B1(new_n15459_), .B2(new_n15458_), .ZN(new_n15689_));
  NAND2_X1   g15392(.A1(new_n15459_), .A2(new_n15458_), .ZN(new_n15690_));
  NOR2_X1    g15393(.A1(new_n15687_), .A2(new_n15684_), .ZN(new_n15691_));
  AOI21_X1   g15394(.A1(new_n15677_), .A2(new_n15682_), .B(new_n15460_), .ZN(new_n15692_));
  NOR3_X1    g15395(.A1(new_n15690_), .A2(new_n15691_), .A3(new_n15692_), .ZN(new_n15693_));
  OAI22_X1   g15396(.A1(new_n1347_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n1344_), .ZN(new_n15694_));
  OAI21_X1   g15397(.A1(new_n7870_), .A2(new_n1457_), .B(new_n15694_), .ZN(new_n15695_));
  AOI21_X1   g15398(.A1(new_n15695_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n15696_));
  XOR2_X1    g15399(.A1(new_n8568_), .A2(new_n15696_), .Z(new_n15697_));
  INV_X1     g15400(.I(new_n15697_), .ZN(new_n15698_));
  OAI21_X1   g15401(.A1(new_n15693_), .A2(new_n15689_), .B(new_n15698_), .ZN(new_n15699_));
  AOI21_X1   g15402(.A1(new_n15456_), .A2(new_n15457_), .B(new_n15699_), .ZN(new_n15700_));
  AOI21_X1   g15403(.A1(new_n15313_), .A2(new_n14673_), .B(new_n14901_), .ZN(new_n15701_));
  OAI21_X1   g15404(.A1(new_n15313_), .A2(new_n14673_), .B(new_n15309_), .ZN(new_n15702_));
  XOR2_X1    g15405(.A1(new_n15292_), .A2(new_n15057_), .Z(new_n15703_));
  OAI22_X1   g15406(.A1(new_n15691_), .A2(new_n15692_), .B1(new_n15703_), .B2(new_n15452_), .ZN(new_n15704_));
  NAND4_X1   g15407(.A1(new_n15688_), .A2(new_n15683_), .A3(new_n15459_), .A4(new_n15458_), .ZN(new_n15705_));
  AOI21_X1   g15408(.A1(new_n15704_), .A2(new_n15705_), .B(new_n15697_), .ZN(new_n15706_));
  NOR3_X1    g15409(.A1(new_n15706_), .A2(new_n15701_), .A3(new_n15702_), .ZN(new_n15707_));
  OAI21_X1   g15410(.A1(new_n15700_), .A2(new_n15707_), .B(new_n15455_), .ZN(new_n15708_));
  INV_X1     g15411(.I(new_n15455_), .ZN(new_n15709_));
  OAI21_X1   g15412(.A1(new_n15701_), .A2(new_n15702_), .B(new_n15706_), .ZN(new_n15710_));
  NAND3_X1   g15413(.A1(new_n15699_), .A2(new_n15457_), .A3(new_n15456_), .ZN(new_n15711_));
  NAND3_X1   g15414(.A1(new_n15710_), .A2(new_n15711_), .A3(new_n15709_), .ZN(new_n15712_));
  OAI22_X1   g15415(.A1(new_n1055_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n1061_), .ZN(new_n15713_));
  OAI21_X1   g15416(.A1(new_n8948_), .A2(new_n1332_), .B(new_n15713_), .ZN(new_n15714_));
  AOI21_X1   g15417(.A1(new_n15714_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n15715_));
  XNOR2_X1   g15418(.A1(new_n9642_), .A2(new_n15715_), .ZN(new_n15716_));
  AOI21_X1   g15419(.A1(new_n15708_), .A2(new_n15712_), .B(new_n15716_), .ZN(new_n15717_));
  NAND2_X1   g15420(.A1(new_n15451_), .A2(new_n15717_), .ZN(new_n15718_));
  OAI21_X1   g15421(.A1(new_n15330_), .A2(new_n15331_), .B(new_n15050_), .ZN(new_n15719_));
  NAND2_X1   g15422(.A1(new_n15719_), .A2(new_n14908_), .ZN(new_n15720_));
  AOI21_X1   g15423(.A1(new_n15710_), .A2(new_n15711_), .B(new_n15709_), .ZN(new_n15721_));
  NOR3_X1    g15424(.A1(new_n15700_), .A2(new_n15707_), .A3(new_n15455_), .ZN(new_n15722_));
  INV_X1     g15425(.I(new_n15716_), .ZN(new_n15723_));
  OAI21_X1   g15426(.A1(new_n15722_), .A2(new_n15721_), .B(new_n15723_), .ZN(new_n15724_));
  NAND3_X1   g15427(.A1(new_n15720_), .A2(new_n14668_), .A3(new_n15724_), .ZN(new_n15725_));
  AOI21_X1   g15428(.A1(new_n15718_), .A2(new_n15725_), .B(new_n15331_), .ZN(new_n15726_));
  AOI21_X1   g15429(.A1(new_n15720_), .A2(new_n14668_), .B(new_n15724_), .ZN(new_n15727_));
  NOR2_X1    g15430(.A1(new_n15451_), .A2(new_n15717_), .ZN(new_n15728_));
  NOR3_X1    g15431(.A1(new_n15727_), .A2(new_n15728_), .A3(new_n15327_), .ZN(new_n15729_));
  NOR2_X1    g15432(.A1(new_n15729_), .A2(new_n15726_), .ZN(new_n15730_));
  NOR2_X1    g15433(.A1(new_n15357_), .A2(new_n15042_), .ZN(new_n15731_));
  OAI22_X1   g15434(.A1(new_n970_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n820_), .ZN(new_n15732_));
  OAI21_X1   g15435(.A1(new_n10031_), .A2(new_n894_), .B(new_n15732_), .ZN(new_n15733_));
  AOI21_X1   g15436(.A1(new_n15733_), .A2(new_n827_), .B(new_n970_), .ZN(new_n15734_));
  XNOR2_X1   g15437(.A1(new_n10866_), .A2(new_n15734_), .ZN(new_n15735_));
  INV_X1     g15438(.I(new_n15735_), .ZN(new_n15736_));
  OAI21_X1   g15439(.A1(new_n15731_), .A2(new_n15356_), .B(new_n15736_), .ZN(new_n15737_));
  NAND2_X1   g15440(.A1(new_n15346_), .A2(new_n15344_), .ZN(new_n15738_));
  NAND3_X1   g15441(.A1(new_n15738_), .A2(new_n15345_), .A3(new_n15735_), .ZN(new_n15739_));
  AOI21_X1   g15442(.A1(new_n15737_), .A2(new_n15739_), .B(new_n15730_), .ZN(new_n15740_));
  OAI21_X1   g15443(.A1(new_n15727_), .A2(new_n15728_), .B(new_n15327_), .ZN(new_n15741_));
  NAND3_X1   g15444(.A1(new_n15718_), .A2(new_n15725_), .A3(new_n15331_), .ZN(new_n15742_));
  NAND2_X1   g15445(.A1(new_n15741_), .A2(new_n15742_), .ZN(new_n15743_));
  NAND3_X1   g15446(.A1(new_n15738_), .A2(new_n15345_), .A3(new_n15736_), .ZN(new_n15744_));
  OAI21_X1   g15447(.A1(new_n15731_), .A2(new_n15356_), .B(new_n15735_), .ZN(new_n15745_));
  AOI21_X1   g15448(.A1(new_n15745_), .A2(new_n15744_), .B(new_n15743_), .ZN(new_n15746_));
  OAI22_X1   g15449(.A1(new_n607_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n610_), .ZN(new_n15747_));
  OAI21_X1   g15450(.A1(new_n11738_), .A2(new_n684_), .B(new_n15747_), .ZN(new_n15748_));
  AOI21_X1   g15451(.A1(new_n15748_), .A2(new_n612_), .B(new_n607_), .ZN(new_n15749_));
  XNOR2_X1   g15452(.A1(new_n12128_), .A2(new_n15749_), .ZN(new_n15750_));
  INV_X1     g15453(.I(new_n15750_), .ZN(new_n15751_));
  OAI21_X1   g15454(.A1(new_n15740_), .A2(new_n15746_), .B(new_n15751_), .ZN(new_n15752_));
  AOI21_X1   g15455(.A1(new_n15447_), .A2(new_n15449_), .B(new_n15752_), .ZN(new_n15753_));
  AOI21_X1   g15456(.A1(new_n15365_), .A2(new_n14934_), .B(new_n14939_), .ZN(new_n15754_));
  OAI21_X1   g15457(.A1(new_n15365_), .A2(new_n14934_), .B(new_n14956_), .ZN(new_n15755_));
  AOI21_X1   g15458(.A1(new_n15738_), .A2(new_n15345_), .B(new_n15735_), .ZN(new_n15756_));
  NOR3_X1    g15459(.A1(new_n15731_), .A2(new_n15356_), .A3(new_n15736_), .ZN(new_n15757_));
  OAI21_X1   g15460(.A1(new_n15757_), .A2(new_n15756_), .B(new_n15743_), .ZN(new_n15758_));
  NOR3_X1    g15461(.A1(new_n15731_), .A2(new_n15356_), .A3(new_n15735_), .ZN(new_n15759_));
  AOI21_X1   g15462(.A1(new_n15738_), .A2(new_n15345_), .B(new_n15736_), .ZN(new_n15760_));
  OAI21_X1   g15463(.A1(new_n15759_), .A2(new_n15760_), .B(new_n15730_), .ZN(new_n15761_));
  AOI21_X1   g15464(.A1(new_n15761_), .A2(new_n15758_), .B(new_n15750_), .ZN(new_n15762_));
  NOR3_X1    g15465(.A1(new_n15754_), .A2(new_n15755_), .A3(new_n15762_), .ZN(new_n15763_));
  OAI21_X1   g15466(.A1(new_n15753_), .A2(new_n15763_), .B(new_n15364_), .ZN(new_n15764_));
  OAI21_X1   g15467(.A1(new_n15754_), .A2(new_n15755_), .B(new_n15762_), .ZN(new_n15765_));
  NAND3_X1   g15468(.A1(new_n15449_), .A2(new_n15752_), .A3(new_n15447_), .ZN(new_n15766_));
  NAND3_X1   g15469(.A1(new_n15765_), .A2(new_n15766_), .A3(new_n15360_), .ZN(new_n15767_));
  NOR3_X1    g15470(.A1(new_n15384_), .A2(new_n15383_), .A3(new_n15387_), .ZN(new_n15768_));
  OAI22_X1   g15471(.A1(new_n448_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n450_), .ZN(new_n15769_));
  OAI21_X1   g15472(.A1(new_n12542_), .A2(new_n496_), .B(new_n15769_), .ZN(new_n15770_));
  AOI21_X1   g15473(.A1(new_n15770_), .A2(new_n452_), .B(new_n448_), .ZN(new_n15771_));
  XNOR2_X1   g15474(.A1(new_n13371_), .A2(new_n15771_), .ZN(new_n15772_));
  INV_X1     g15475(.I(new_n15772_), .ZN(new_n15773_));
  OAI21_X1   g15476(.A1(new_n15768_), .A2(new_n15385_), .B(new_n15773_), .ZN(new_n15774_));
  INV_X1     g15477(.I(new_n15385_), .ZN(new_n15775_));
  NAND3_X1   g15478(.A1(new_n15369_), .A2(new_n15371_), .A3(new_n15386_), .ZN(new_n15776_));
  NAND3_X1   g15479(.A1(new_n15776_), .A2(new_n15775_), .A3(new_n15772_), .ZN(new_n15777_));
  AOI22_X1   g15480(.A1(new_n15774_), .A2(new_n15777_), .B1(new_n15764_), .B2(new_n15767_), .ZN(new_n15778_));
  NAND2_X1   g15481(.A1(new_n15764_), .A2(new_n15767_), .ZN(new_n15779_));
  NAND3_X1   g15482(.A1(new_n15776_), .A2(new_n15775_), .A3(new_n15773_), .ZN(new_n15780_));
  OAI21_X1   g15483(.A1(new_n15768_), .A2(new_n15385_), .B(new_n15772_), .ZN(new_n15781_));
  AOI21_X1   g15484(.A1(new_n15780_), .A2(new_n15781_), .B(new_n15779_), .ZN(new_n15782_));
  NOR2_X1    g15485(.A1(new_n15782_), .A2(new_n15778_), .ZN(new_n15783_));
  NOR3_X1    g15486(.A1(new_n15445_), .A2(new_n15783_), .A3(new_n15441_), .ZN(new_n15784_));
  INV_X1     g15487(.I(new_n15441_), .ZN(new_n15785_));
  INV_X1     g15488(.I(new_n15442_), .ZN(new_n15786_));
  NOR3_X1    g15489(.A1(new_n15404_), .A2(new_n15403_), .A3(new_n15026_), .ZN(new_n15787_));
  AOI21_X1   g15490(.A1(new_n15390_), .A2(new_n15395_), .B(new_n15427_), .ZN(new_n15788_));
  OAI21_X1   g15491(.A1(new_n15787_), .A2(new_n15788_), .B(new_n15786_), .ZN(new_n15789_));
  AOI21_X1   g15492(.A1(new_n15765_), .A2(new_n15766_), .B(new_n15360_), .ZN(new_n15790_));
  NOR3_X1    g15493(.A1(new_n15753_), .A2(new_n15763_), .A3(new_n15364_), .ZN(new_n15791_));
  AOI21_X1   g15494(.A1(new_n15776_), .A2(new_n15775_), .B(new_n15772_), .ZN(new_n15792_));
  NOR3_X1    g15495(.A1(new_n15768_), .A2(new_n15385_), .A3(new_n15773_), .ZN(new_n15793_));
  OAI22_X1   g15496(.A1(new_n15793_), .A2(new_n15792_), .B1(new_n15790_), .B2(new_n15791_), .ZN(new_n15794_));
  NOR2_X1    g15497(.A1(new_n15791_), .A2(new_n15790_), .ZN(new_n15795_));
  NOR3_X1    g15498(.A1(new_n15768_), .A2(new_n15385_), .A3(new_n15772_), .ZN(new_n15796_));
  AOI21_X1   g15499(.A1(new_n15776_), .A2(new_n15775_), .B(new_n15773_), .ZN(new_n15797_));
  OAI21_X1   g15500(.A1(new_n15796_), .A2(new_n15797_), .B(new_n15795_), .ZN(new_n15798_));
  NAND2_X1   g15501(.A1(new_n15798_), .A2(new_n15794_), .ZN(new_n15799_));
  AOI21_X1   g15502(.A1(new_n15785_), .A2(new_n15789_), .B(new_n15799_), .ZN(new_n15800_));
  OAI21_X1   g15503(.A1(new_n15800_), .A2(new_n15784_), .B(new_n15440_), .ZN(new_n15801_));
  AOI21_X1   g15504(.A1(new_n15438_), .A2(new_n15436_), .B(new_n15433_), .ZN(new_n15802_));
  NOR3_X1    g15505(.A1(new_n15429_), .A2(new_n15426_), .A3(new_n15434_), .ZN(new_n15803_));
  NOR2_X1    g15506(.A1(new_n15803_), .A2(new_n15802_), .ZN(new_n15804_));
  AOI21_X1   g15507(.A1(new_n15789_), .A2(new_n15785_), .B(new_n15783_), .ZN(new_n15805_));
  NOR3_X1    g15508(.A1(new_n15445_), .A2(new_n15799_), .A3(new_n15441_), .ZN(new_n15806_));
  OAI21_X1   g15509(.A1(new_n15805_), .A2(new_n15806_), .B(new_n15804_), .ZN(new_n15807_));
  AOI21_X1   g15510(.A1(new_n15801_), .A2(new_n15807_), .B(new_n15418_), .ZN(new_n15808_));
  XOR2_X1    g15511(.A1(new_n15808_), .A2(new_n15420_), .Z(new_n15809_));
  XOR2_X1    g15512(.A1(new_n15809_), .A2(new_n15022_), .Z(\f[66] ));
  NOR2_X1    g15513(.A1(new_n15445_), .A2(new_n15441_), .ZN(new_n15811_));
  NOR2_X1    g15514(.A1(new_n15440_), .A2(new_n15783_), .ZN(new_n15812_));
  NOR2_X1    g15515(.A1(new_n15804_), .A2(new_n15799_), .ZN(new_n15813_));
  OAI21_X1   g15516(.A1(new_n15813_), .A2(new_n15812_), .B(new_n15811_), .ZN(new_n15814_));
  NAND2_X1   g15517(.A1(new_n15001_), .A2(new_n14632_), .ZN(new_n15815_));
  OAI21_X1   g15518(.A1(new_n15001_), .A2(new_n14632_), .B(new_n15007_), .ZN(new_n15816_));
  OAI21_X1   g15519(.A1(new_n14646_), .A2(new_n15816_), .B(new_n15815_), .ZN(new_n15817_));
  NAND3_X1   g15520(.A1(new_n15789_), .A2(new_n15799_), .A3(new_n15785_), .ZN(new_n15818_));
  OAI21_X1   g15521(.A1(new_n15441_), .A2(new_n15445_), .B(new_n15783_), .ZN(new_n15819_));
  AOI21_X1   g15522(.A1(new_n15819_), .A2(new_n15818_), .B(new_n15804_), .ZN(new_n15820_));
  OAI22_X1   g15523(.A1(new_n15445_), .A2(new_n15441_), .B1(new_n15778_), .B2(new_n15782_), .ZN(new_n15821_));
  NAND3_X1   g15524(.A1(new_n15789_), .A2(new_n15783_), .A3(new_n15785_), .ZN(new_n15822_));
  AOI21_X1   g15525(.A1(new_n15821_), .A2(new_n15822_), .B(new_n15440_), .ZN(new_n15823_));
  OAI21_X1   g15526(.A1(new_n15820_), .A2(new_n15823_), .B(new_n15419_), .ZN(new_n15824_));
  NAND2_X1   g15527(.A1(new_n15824_), .A2(new_n15421_), .ZN(new_n15825_));
  NAND3_X1   g15528(.A1(new_n15807_), .A2(new_n15801_), .A3(new_n15417_), .ZN(new_n15826_));
  NAND3_X1   g15529(.A1(new_n15825_), .A2(new_n15817_), .A3(new_n15826_), .ZN(new_n15827_));
  NOR2_X1    g15530(.A1(new_n15783_), .A2(new_n15433_), .ZN(new_n15828_));
  AOI22_X1   g15531(.A1(new_n15783_), .A2(new_n15433_), .B1(new_n15436_), .B2(new_n15438_), .ZN(new_n15829_));
  NOR2_X1    g15532(.A1(new_n15829_), .A2(new_n15828_), .ZN(new_n15830_));
  NAND2_X1   g15533(.A1(new_n15761_), .A2(new_n15758_), .ZN(new_n15831_));
  NAND2_X1   g15534(.A1(new_n15831_), .A2(new_n15360_), .ZN(new_n15832_));
  INV_X1     g15535(.I(new_n15832_), .ZN(new_n15833_));
  OAI21_X1   g15536(.A1(new_n15831_), .A2(new_n15360_), .B(new_n15751_), .ZN(new_n15834_));
  NOR3_X1    g15537(.A1(new_n15834_), .A2(new_n15754_), .A3(new_n15755_), .ZN(new_n15835_));
  NOR2_X1    g15538(.A1(new_n15835_), .A2(new_n15833_), .ZN(new_n15836_));
  INV_X1     g15539(.I(new_n15451_), .ZN(new_n15837_));
  AOI21_X1   g15540(.A1(new_n15708_), .A2(new_n15712_), .B(new_n15327_), .ZN(new_n15838_));
  NOR3_X1    g15541(.A1(new_n15722_), .A2(new_n15721_), .A3(new_n15331_), .ZN(new_n15839_));
  NOR2_X1    g15542(.A1(new_n15839_), .A2(new_n15716_), .ZN(new_n15840_));
  AOI21_X1   g15543(.A1(new_n15837_), .A2(new_n15840_), .B(new_n15838_), .ZN(new_n15841_));
  INV_X1     g15544(.I(new_n15677_), .ZN(new_n15842_));
  NOR2_X1    g15545(.A1(new_n15690_), .A2(new_n15842_), .ZN(new_n15843_));
  NAND2_X1   g15546(.A1(new_n15684_), .A2(new_n15682_), .ZN(new_n15844_));
  AOI21_X1   g15547(.A1(new_n15690_), .A2(new_n15842_), .B(new_n15844_), .ZN(new_n15845_));
  NOR2_X1    g15548(.A1(new_n15845_), .A2(new_n15843_), .ZN(new_n15846_));
  AOI21_X1   g15549(.A1(new_n15669_), .A2(new_n15670_), .B(new_n15288_), .ZN(new_n15847_));
  NAND2_X1   g15550(.A1(new_n15669_), .A2(new_n15670_), .ZN(new_n15848_));
  NOR2_X1    g15551(.A1(new_n15848_), .A2(new_n15263_), .ZN(new_n15849_));
  NOR4_X1    g15552(.A1(new_n15849_), .A2(new_n15289_), .A3(new_n15268_), .A4(new_n15665_), .ZN(new_n15850_));
  NOR2_X1    g15553(.A1(new_n15850_), .A2(new_n15847_), .ZN(new_n15851_));
  INV_X1     g15554(.I(new_n15851_), .ZN(new_n15852_));
  NAND2_X1   g15555(.A1(new_n15461_), .A2(new_n15233_), .ZN(new_n15853_));
  INV_X1     g15556(.I(new_n15645_), .ZN(new_n15854_));
  NOR2_X1    g15557(.A1(new_n15853_), .A2(new_n15854_), .ZN(new_n15855_));
  NAND2_X1   g15558(.A1(new_n15651_), .A2(new_n15649_), .ZN(new_n15856_));
  AOI21_X1   g15559(.A1(new_n15853_), .A2(new_n15854_), .B(new_n15856_), .ZN(new_n15857_));
  NOR2_X1    g15560(.A1(new_n15857_), .A2(new_n15855_), .ZN(new_n15858_));
  NOR2_X1    g15561(.A1(new_n15466_), .A2(new_n15640_), .ZN(new_n15859_));
  NAND2_X1   g15562(.A1(new_n15634_), .A2(new_n15632_), .ZN(new_n15860_));
  OAI21_X1   g15563(.A1(new_n15471_), .A2(new_n15192_), .B(new_n15615_), .ZN(new_n15861_));
  INV_X1     g15564(.I(new_n15473_), .ZN(new_n15862_));
  AOI21_X1   g15565(.A1(new_n15476_), .A2(new_n15862_), .B(new_n15587_), .ZN(new_n15863_));
  NOR2_X1    g15566(.A1(new_n15863_), .A2(new_n15584_), .ZN(new_n15864_));
  INV_X1     g15567(.I(new_n15864_), .ZN(new_n15865_));
  NAND2_X1   g15568(.A1(new_n15478_), .A2(new_n15167_), .ZN(new_n15866_));
  NAND2_X1   g15569(.A1(new_n15866_), .A2(new_n15573_), .ZN(new_n15867_));
  NOR2_X1    g15570(.A1(new_n15481_), .A2(new_n15564_), .ZN(new_n15868_));
  NOR2_X1    g15571(.A1(new_n15868_), .A2(new_n15563_), .ZN(new_n15869_));
  INV_X1     g15572(.I(new_n15869_), .ZN(new_n15870_));
  NOR2_X1    g15573(.A1(new_n15549_), .A2(new_n15547_), .ZN(new_n15871_));
  NOR2_X1    g15574(.A1(new_n15871_), .A2(new_n15543_), .ZN(new_n15872_));
  INV_X1     g15575(.I(new_n15484_), .ZN(new_n15873_));
  AOI21_X1   g15576(.A1(new_n15873_), .A2(new_n15531_), .B(new_n15529_), .ZN(new_n15874_));
  NOR2_X1    g15577(.A1(new_n15523_), .A2(new_n15485_), .ZN(new_n15875_));
  NOR2_X1    g15578(.A1(new_n15875_), .A2(new_n15521_), .ZN(new_n15876_));
  NOR2_X1    g15579(.A1(new_n15510_), .A2(new_n15508_), .ZN(new_n15877_));
  OAI22_X1   g15580(.A1(new_n13880_), .A2(new_n509_), .B1(new_n419_), .B2(new_n13885_), .ZN(new_n15878_));
  AOI21_X1   g15581(.A1(new_n15878_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n15879_));
  XOR2_X1    g15582(.A1(new_n471_), .A2(new_n15879_), .Z(new_n15880_));
  NOR2_X1    g15583(.A1(new_n13476_), .A2(new_n298_), .ZN(new_n15881_));
  XOR2_X1    g15584(.A1(new_n14736_), .A2(new_n298_), .Z(new_n15882_));
  NAND2_X1   g15585(.A1(new_n15882_), .A2(\b[4] ), .ZN(new_n15883_));
  XOR2_X1    g15586(.A1(new_n15883_), .A2(new_n15881_), .Z(new_n15884_));
  AND2_X2    g15587(.A1(new_n15884_), .A2(\a[2] ), .Z(new_n15885_));
  NOR2_X1    g15588(.A1(new_n15884_), .A2(\a[2] ), .ZN(new_n15886_));
  NOR2_X1    g15589(.A1(new_n15885_), .A2(new_n15886_), .ZN(new_n15887_));
  NOR2_X1    g15590(.A1(new_n15880_), .A2(new_n15887_), .ZN(new_n15888_));
  XOR2_X1    g15591(.A1(new_n15884_), .A2(new_n260_), .Z(new_n15889_));
  INV_X1     g15592(.I(new_n15889_), .ZN(new_n15890_));
  AOI21_X1   g15593(.A1(new_n15880_), .A2(new_n15890_), .B(new_n15888_), .ZN(new_n15891_));
  INV_X1     g15594(.I(new_n15891_), .ZN(new_n15892_));
  INV_X1     g15595(.I(new_n15498_), .ZN(new_n15893_));
  AOI21_X1   g15596(.A1(new_n15490_), .A2(new_n15893_), .B(new_n15499_), .ZN(new_n15894_));
  AOI22_X1   g15597(.A1(new_n13078_), .A2(\b[8] ), .B1(new_n13503_), .B2(new_n12218_), .ZN(new_n15895_));
  OAI21_X1   g15598(.A1(new_n15895_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n15896_));
  XOR2_X1    g15599(.A1(new_n660_), .A2(new_n15896_), .Z(new_n15897_));
  NOR2_X1    g15600(.A1(new_n15897_), .A2(new_n15894_), .ZN(new_n15898_));
  AND2_X2    g15601(.A1(new_n15897_), .A2(new_n15894_), .Z(new_n15899_));
  OAI21_X1   g15602(.A1(new_n15899_), .A2(new_n15898_), .B(new_n15892_), .ZN(new_n15900_));
  XOR2_X1    g15603(.A1(new_n15897_), .A2(new_n15894_), .Z(new_n15901_));
  NAND2_X1   g15604(.A1(new_n15901_), .A2(new_n15891_), .ZN(new_n15902_));
  NAND2_X1   g15605(.A1(new_n15902_), .A2(new_n15900_), .ZN(new_n15903_));
  AOI22_X1   g15606(.A1(new_n10969_), .A2(new_n927_), .B1(new_n11394_), .B2(\b[11] ), .ZN(new_n15904_));
  OAI21_X1   g15607(.A1(new_n15904_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n15905_));
  XNOR2_X1   g15608(.A1(new_n860_), .A2(new_n15905_), .ZN(new_n15906_));
  INV_X1     g15609(.I(new_n15906_), .ZN(new_n15907_));
  NOR2_X1    g15610(.A1(new_n15903_), .A2(new_n15907_), .ZN(new_n15908_));
  INV_X1     g15611(.I(new_n15903_), .ZN(new_n15909_));
  NOR2_X1    g15612(.A1(new_n15909_), .A2(new_n15906_), .ZN(new_n15910_));
  OAI22_X1   g15613(.A1(new_n15910_), .A2(new_n15908_), .B1(new_n15505_), .B2(new_n15877_), .ZN(new_n15911_));
  NOR2_X1    g15614(.A1(new_n15877_), .A2(new_n15505_), .ZN(new_n15912_));
  NOR2_X1    g15615(.A1(new_n15909_), .A2(new_n15907_), .ZN(new_n15913_));
  NOR2_X1    g15616(.A1(new_n15903_), .A2(new_n15906_), .ZN(new_n15914_));
  OAI21_X1   g15617(.A1(new_n15913_), .A2(new_n15914_), .B(new_n15912_), .ZN(new_n15915_));
  AOI22_X1   g15618(.A1(new_n11415_), .A2(new_n1111_), .B1(\b[14] ), .B2(new_n10145_), .ZN(new_n15916_));
  OAI21_X1   g15619(.A1(new_n15916_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n15917_));
  XOR2_X1    g15620(.A1(new_n1114_), .A2(new_n15917_), .Z(new_n15918_));
  NAND3_X1   g15621(.A1(new_n15911_), .A2(new_n15915_), .A3(new_n15918_), .ZN(new_n15919_));
  NAND2_X1   g15622(.A1(new_n15911_), .A2(new_n15915_), .ZN(new_n15920_));
  INV_X1     g15623(.I(new_n15918_), .ZN(new_n15921_));
  NAND2_X1   g15624(.A1(new_n15920_), .A2(new_n15921_), .ZN(new_n15922_));
  AOI21_X1   g15625(.A1(new_n15922_), .A2(new_n15919_), .B(new_n15876_), .ZN(new_n15923_));
  INV_X1     g15626(.I(new_n15876_), .ZN(new_n15924_));
  XOR2_X1    g15627(.A1(new_n15920_), .A2(new_n15918_), .Z(new_n15925_));
  NOR2_X1    g15628(.A1(new_n15925_), .A2(new_n15924_), .ZN(new_n15926_));
  NOR2_X1    g15629(.A1(new_n15926_), .A2(new_n15923_), .ZN(new_n15927_));
  OAI22_X1   g15630(.A1(new_n8644_), .A2(new_n1294_), .B1(new_n1518_), .B2(new_n9388_), .ZN(new_n15928_));
  OAI21_X1   g15631(.A1(new_n1189_), .A2(new_n10154_), .B(new_n15928_), .ZN(new_n15929_));
  AOI21_X1   g15632(.A1(new_n15929_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n15930_));
  XNOR2_X1   g15633(.A1(new_n1421_), .A2(new_n15930_), .ZN(new_n15931_));
  NOR2_X1    g15634(.A1(new_n15927_), .A2(new_n15931_), .ZN(new_n15932_));
  NAND2_X1   g15635(.A1(new_n15927_), .A2(new_n15931_), .ZN(new_n15933_));
  INV_X1     g15636(.I(new_n15933_), .ZN(new_n15934_));
  NOR2_X1    g15637(.A1(new_n15934_), .A2(new_n15932_), .ZN(new_n15935_));
  NOR2_X1    g15638(.A1(new_n15935_), .A2(new_n15874_), .ZN(new_n15936_));
  INV_X1     g15639(.I(new_n15874_), .ZN(new_n15937_));
  XNOR2_X1   g15640(.A1(new_n15927_), .A2(new_n15931_), .ZN(new_n15938_));
  NOR2_X1    g15641(.A1(new_n15938_), .A2(new_n15937_), .ZN(new_n15939_));
  NOR2_X1    g15642(.A1(new_n15936_), .A2(new_n15939_), .ZN(new_n15940_));
  OAI22_X1   g15643(.A1(new_n7619_), .A2(new_n1634_), .B1(new_n1803_), .B2(new_n8309_), .ZN(new_n15941_));
  OAI21_X1   g15644(.A1(new_n1525_), .A2(new_n7947_), .B(new_n15941_), .ZN(new_n15942_));
  AOI21_X1   g15645(.A1(new_n15942_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n15943_));
  XOR2_X1    g15646(.A1(new_n1808_), .A2(new_n15943_), .Z(new_n15944_));
  NOR2_X1    g15647(.A1(new_n15940_), .A2(new_n15944_), .ZN(new_n15945_));
  INV_X1     g15648(.I(new_n15945_), .ZN(new_n15946_));
  NAND2_X1   g15649(.A1(new_n15940_), .A2(new_n15944_), .ZN(new_n15947_));
  AOI21_X1   g15650(.A1(new_n15946_), .A2(new_n15947_), .B(new_n15872_), .ZN(new_n15948_));
  INV_X1     g15651(.I(new_n15872_), .ZN(new_n15949_));
  XNOR2_X1   g15652(.A1(new_n15940_), .A2(new_n15944_), .ZN(new_n15950_));
  NOR2_X1    g15653(.A1(new_n15950_), .A2(new_n15949_), .ZN(new_n15951_));
  NOR2_X1    g15654(.A1(new_n15951_), .A2(new_n15948_), .ZN(new_n15952_));
  OAI22_X1   g15655(.A1(new_n6644_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n6647_), .ZN(new_n15953_));
  OAI21_X1   g15656(.A1(new_n1936_), .A2(new_n7284_), .B(new_n15953_), .ZN(new_n15954_));
  AOI21_X1   g15657(.A1(new_n15954_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n15955_));
  XNOR2_X1   g15658(.A1(new_n2280_), .A2(new_n15955_), .ZN(new_n15956_));
  NOR2_X1    g15659(.A1(new_n15952_), .A2(new_n15956_), .ZN(new_n15957_));
  NAND2_X1   g15660(.A1(new_n15952_), .A2(new_n15956_), .ZN(new_n15958_));
  INV_X1     g15661(.I(new_n15958_), .ZN(new_n15959_));
  OAI21_X1   g15662(.A1(new_n15959_), .A2(new_n15957_), .B(new_n15870_), .ZN(new_n15960_));
  XNOR2_X1   g15663(.A1(new_n15952_), .A2(new_n15956_), .ZN(new_n15961_));
  OAI21_X1   g15664(.A1(new_n15870_), .A2(new_n15961_), .B(new_n15960_), .ZN(new_n15962_));
  OAI22_X1   g15665(.A1(new_n5993_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n5991_), .ZN(new_n15963_));
  OAI21_X1   g15666(.A1(new_n2439_), .A2(new_n5997_), .B(new_n15963_), .ZN(new_n15964_));
  AOI21_X1   g15667(.A1(new_n15964_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n15965_));
  XNOR2_X1   g15668(.A1(new_n2846_), .A2(new_n15965_), .ZN(new_n15966_));
  INV_X1     g15669(.I(new_n15966_), .ZN(new_n15967_));
  NAND2_X1   g15670(.A1(new_n15962_), .A2(new_n15967_), .ZN(new_n15968_));
  INV_X1     g15671(.I(new_n15960_), .ZN(new_n15969_));
  NOR2_X1    g15672(.A1(new_n15961_), .A2(new_n15870_), .ZN(new_n15970_));
  OR3_X2     g15673(.A1(new_n15970_), .A2(new_n15969_), .A3(new_n15967_), .Z(new_n15971_));
  AOI22_X1   g15674(.A1(new_n15971_), .A2(new_n15968_), .B1(new_n15571_), .B2(new_n15867_), .ZN(new_n15972_));
  NAND2_X1   g15675(.A1(new_n15867_), .A2(new_n15571_), .ZN(new_n15973_));
  XOR2_X1    g15676(.A1(new_n15962_), .A2(new_n15966_), .Z(new_n15974_));
  NOR2_X1    g15677(.A1(new_n15974_), .A2(new_n15973_), .ZN(new_n15975_));
  OR2_X2     g15678(.A1(new_n15975_), .A2(new_n15972_), .Z(new_n15976_));
  OAI22_X1   g15679(.A1(new_n5420_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n5107_), .ZN(new_n15977_));
  OAI21_X1   g15680(.A1(new_n3018_), .A2(new_n5112_), .B(new_n15977_), .ZN(new_n15978_));
  AOI21_X1   g15681(.A1(new_n15978_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n15979_));
  XNOR2_X1   g15682(.A1(new_n3514_), .A2(new_n15979_), .ZN(new_n15980_));
  NOR2_X1    g15683(.A1(new_n15976_), .A2(new_n15980_), .ZN(new_n15981_));
  NOR2_X1    g15684(.A1(new_n15975_), .A2(new_n15972_), .ZN(new_n15982_));
  INV_X1     g15685(.I(new_n15980_), .ZN(new_n15983_));
  NOR2_X1    g15686(.A1(new_n15982_), .A2(new_n15983_), .ZN(new_n15984_));
  OAI21_X1   g15687(.A1(new_n15981_), .A2(new_n15984_), .B(new_n15865_), .ZN(new_n15985_));
  NOR2_X1    g15688(.A1(new_n15982_), .A2(new_n15980_), .ZN(new_n15986_));
  NOR2_X1    g15689(.A1(new_n15976_), .A2(new_n15983_), .ZN(new_n15987_));
  OAI21_X1   g15690(.A1(new_n15987_), .A2(new_n15986_), .B(new_n15864_), .ZN(new_n15988_));
  NAND2_X1   g15691(.A1(new_n15988_), .A2(new_n15985_), .ZN(new_n15989_));
  OAI22_X1   g15692(.A1(new_n4072_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n4067_), .ZN(new_n15990_));
  OAI21_X1   g15693(.A1(new_n3717_), .A2(new_n4318_), .B(new_n15990_), .ZN(new_n15991_));
  AOI21_X1   g15694(.A1(new_n15991_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n15992_));
  XNOR2_X1   g15695(.A1(new_n4257_), .A2(new_n15992_), .ZN(new_n15993_));
  NOR2_X1    g15696(.A1(new_n15989_), .A2(new_n15993_), .ZN(new_n15994_));
  INV_X1     g15697(.I(new_n15994_), .ZN(new_n15995_));
  NAND2_X1   g15698(.A1(new_n15989_), .A2(new_n15993_), .ZN(new_n15996_));
  AOI22_X1   g15699(.A1(new_n15995_), .A2(new_n15996_), .B1(new_n15614_), .B2(new_n15861_), .ZN(new_n15997_));
  NAND2_X1   g15700(.A1(new_n15861_), .A2(new_n15614_), .ZN(new_n15998_));
  INV_X1     g15701(.I(new_n15993_), .ZN(new_n15999_));
  XOR2_X1    g15702(.A1(new_n15989_), .A2(new_n15999_), .Z(new_n16000_));
  NOR2_X1    g15703(.A1(new_n16000_), .A2(new_n15998_), .ZN(new_n16001_));
  NOR2_X1    g15704(.A1(new_n16001_), .A2(new_n15997_), .ZN(new_n16002_));
  OAI22_X1   g15705(.A1(new_n4774_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n5068_), .ZN(new_n16003_));
  OAI21_X1   g15706(.A1(new_n4500_), .A2(new_n3569_), .B(new_n16003_), .ZN(new_n16004_));
  AOI21_X1   g15707(.A1(new_n16004_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n16005_));
  XOR2_X1    g15708(.A1(new_n5067_), .A2(new_n16005_), .Z(new_n16006_));
  INV_X1     g15709(.I(new_n16006_), .ZN(new_n16007_));
  NAND2_X1   g15710(.A1(new_n16002_), .A2(new_n16007_), .ZN(new_n16008_));
  INV_X1     g15711(.I(new_n15996_), .ZN(new_n16009_));
  OAI21_X1   g15712(.A1(new_n16009_), .A2(new_n15994_), .B(new_n15998_), .ZN(new_n16010_));
  XOR2_X1    g15713(.A1(new_n15989_), .A2(new_n15993_), .Z(new_n16011_));
  NAND3_X1   g15714(.A1(new_n16011_), .A2(new_n15614_), .A3(new_n15861_), .ZN(new_n16012_));
  NAND2_X1   g15715(.A1(new_n16012_), .A2(new_n16010_), .ZN(new_n16013_));
  NAND2_X1   g15716(.A1(new_n16013_), .A2(new_n16006_), .ZN(new_n16014_));
  AOI22_X1   g15717(.A1(new_n16014_), .A2(new_n16008_), .B1(new_n15631_), .B2(new_n15860_), .ZN(new_n16015_));
  NAND2_X1   g15718(.A1(new_n15860_), .A2(new_n15631_), .ZN(new_n16016_));
  NAND2_X1   g15719(.A1(new_n16013_), .A2(new_n16007_), .ZN(new_n16017_));
  NAND3_X1   g15720(.A1(new_n16012_), .A2(new_n16010_), .A3(new_n16006_), .ZN(new_n16018_));
  AOI21_X1   g15721(.A1(new_n16017_), .A2(new_n16018_), .B(new_n16016_), .ZN(new_n16019_));
  OAI22_X1   g15722(.A1(new_n5913_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n5921_), .ZN(new_n16020_));
  OAI21_X1   g15723(.A1(new_n5353_), .A2(new_n2884_), .B(new_n16020_), .ZN(new_n16021_));
  AOI21_X1   g15724(.A1(new_n16021_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n16022_));
  XOR2_X1    g15725(.A1(new_n5926_), .A2(new_n16022_), .Z(new_n16023_));
  NOR3_X1    g15726(.A1(new_n16015_), .A2(new_n16019_), .A3(new_n16023_), .ZN(new_n16024_));
  NAND2_X1   g15727(.A1(new_n16014_), .A2(new_n16008_), .ZN(new_n16025_));
  NAND2_X1   g15728(.A1(new_n16025_), .A2(new_n16016_), .ZN(new_n16026_));
  INV_X1     g15729(.I(new_n16019_), .ZN(new_n16027_));
  INV_X1     g15730(.I(new_n16023_), .ZN(new_n16028_));
  AOI21_X1   g15731(.A1(new_n16026_), .A2(new_n16027_), .B(new_n16028_), .ZN(new_n16029_));
  OAI22_X1   g15732(.A1(new_n16029_), .A2(new_n16024_), .B1(new_n15630_), .B2(new_n15859_), .ZN(new_n16030_));
  NOR2_X1    g15733(.A1(new_n15859_), .A2(new_n15630_), .ZN(new_n16031_));
  AOI21_X1   g15734(.A1(new_n16026_), .A2(new_n16027_), .B(new_n16023_), .ZN(new_n16032_));
  NOR3_X1    g15735(.A1(new_n16015_), .A2(new_n16019_), .A3(new_n16028_), .ZN(new_n16033_));
  OAI21_X1   g15736(.A1(new_n16032_), .A2(new_n16033_), .B(new_n16031_), .ZN(new_n16034_));
  OAI22_X1   g15737(.A1(new_n2171_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n2166_), .ZN(new_n16035_));
  OAI21_X1   g15738(.A1(new_n6229_), .A2(new_n2322_), .B(new_n16035_), .ZN(new_n16036_));
  AOI21_X1   g15739(.A1(new_n16036_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n16037_));
  XOR2_X1    g15740(.A1(new_n6851_), .A2(new_n16037_), .Z(new_n16038_));
  AOI21_X1   g15741(.A1(new_n16030_), .A2(new_n16034_), .B(new_n16038_), .ZN(new_n16039_));
  INV_X1     g15742(.I(new_n16039_), .ZN(new_n16040_));
  NAND3_X1   g15743(.A1(new_n16030_), .A2(new_n16034_), .A3(new_n16038_), .ZN(new_n16041_));
  AOI21_X1   g15744(.A1(new_n16040_), .A2(new_n16041_), .B(new_n15858_), .ZN(new_n16042_));
  INV_X1     g15745(.I(new_n15858_), .ZN(new_n16043_));
  INV_X1     g15746(.I(new_n16038_), .ZN(new_n16044_));
  NAND3_X1   g15747(.A1(new_n16030_), .A2(new_n16034_), .A3(new_n16044_), .ZN(new_n16045_));
  AOI21_X1   g15748(.A1(new_n16030_), .A2(new_n16034_), .B(new_n16044_), .ZN(new_n16046_));
  INV_X1     g15749(.I(new_n16046_), .ZN(new_n16047_));
  AOI21_X1   g15750(.A1(new_n16047_), .A2(new_n16045_), .B(new_n16043_), .ZN(new_n16048_));
  NOR2_X1    g15751(.A1(new_n16048_), .A2(new_n16042_), .ZN(new_n16049_));
  OAI22_X1   g15752(.A1(new_n1712_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n1707_), .ZN(new_n16050_));
  OAI21_X1   g15753(.A1(new_n7198_), .A2(new_n1850_), .B(new_n16050_), .ZN(new_n16051_));
  AOI21_X1   g15754(.A1(new_n16051_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n16052_));
  XNOR2_X1   g15755(.A1(new_n7874_), .A2(new_n16052_), .ZN(new_n16053_));
  NOR2_X1    g15756(.A1(new_n16049_), .A2(new_n16053_), .ZN(new_n16054_));
  INV_X1     g15757(.I(new_n16041_), .ZN(new_n16055_));
  OAI21_X1   g15758(.A1(new_n16055_), .A2(new_n16039_), .B(new_n16043_), .ZN(new_n16056_));
  INV_X1     g15759(.I(new_n16045_), .ZN(new_n16057_));
  OAI21_X1   g15760(.A1(new_n16057_), .A2(new_n16046_), .B(new_n15858_), .ZN(new_n16058_));
  NAND2_X1   g15761(.A1(new_n16056_), .A2(new_n16058_), .ZN(new_n16059_));
  INV_X1     g15762(.I(new_n16053_), .ZN(new_n16060_));
  NOR2_X1    g15763(.A1(new_n16059_), .A2(new_n16060_), .ZN(new_n16061_));
  OAI21_X1   g15764(.A1(new_n16054_), .A2(new_n16061_), .B(new_n15852_), .ZN(new_n16062_));
  NOR2_X1    g15765(.A1(new_n16059_), .A2(new_n16053_), .ZN(new_n16063_));
  NOR2_X1    g15766(.A1(new_n16049_), .A2(new_n16060_), .ZN(new_n16064_));
  OAI21_X1   g15767(.A1(new_n16064_), .A2(new_n16063_), .B(new_n15851_), .ZN(new_n16065_));
  OAI22_X1   g15768(.A1(new_n1347_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n1344_), .ZN(new_n16066_));
  OAI21_X1   g15769(.A1(new_n8218_), .A2(new_n1457_), .B(new_n16066_), .ZN(new_n16067_));
  AOI21_X1   g15770(.A1(new_n16067_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n16068_));
  XOR2_X1    g15771(.A1(new_n8952_), .A2(new_n16068_), .Z(new_n16069_));
  AOI21_X1   g15772(.A1(new_n16062_), .A2(new_n16065_), .B(new_n16069_), .ZN(new_n16070_));
  NAND2_X1   g15773(.A1(new_n16062_), .A2(new_n16065_), .ZN(new_n16071_));
  INV_X1     g15774(.I(new_n16069_), .ZN(new_n16072_));
  NOR2_X1    g15775(.A1(new_n16071_), .A2(new_n16072_), .ZN(new_n16073_));
  NOR2_X1    g15776(.A1(new_n16073_), .A2(new_n16070_), .ZN(new_n16074_));
  NOR2_X1    g15777(.A1(new_n16074_), .A2(new_n15846_), .ZN(new_n16075_));
  XOR2_X1    g15778(.A1(new_n16071_), .A2(new_n16072_), .Z(new_n16076_));
  AOI21_X1   g15779(.A1(new_n15846_), .A2(new_n16076_), .B(new_n16075_), .ZN(new_n16077_));
  NAND2_X1   g15780(.A1(new_n15457_), .A2(new_n15456_), .ZN(new_n16078_));
  NOR2_X1    g15781(.A1(new_n15693_), .A2(new_n15689_), .ZN(new_n16079_));
  OR2_X2     g15782(.A1(new_n16078_), .A2(new_n16079_), .Z(new_n16080_));
  NAND2_X1   g15783(.A1(new_n16078_), .A2(new_n16079_), .ZN(new_n16081_));
  NOR2_X1    g15784(.A1(new_n15455_), .A2(new_n15697_), .ZN(new_n16082_));
  NAND2_X1   g15785(.A1(new_n16081_), .A2(new_n16082_), .ZN(new_n16083_));
  NAND2_X1   g15786(.A1(new_n16083_), .A2(new_n16080_), .ZN(new_n16084_));
  OAI22_X1   g15787(.A1(new_n1055_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n1061_), .ZN(new_n16085_));
  OAI21_X1   g15788(.A1(new_n9295_), .A2(new_n1332_), .B(new_n16085_), .ZN(new_n16086_));
  AOI21_X1   g15789(.A1(new_n16086_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n16087_));
  XNOR2_X1   g15790(.A1(new_n10035_), .A2(new_n16087_), .ZN(new_n16088_));
  INV_X1     g15791(.I(new_n16088_), .ZN(new_n16089_));
  NAND2_X1   g15792(.A1(new_n16084_), .A2(new_n16089_), .ZN(new_n16090_));
  NOR2_X1    g15793(.A1(new_n16084_), .A2(new_n16089_), .ZN(new_n16091_));
  INV_X1     g15794(.I(new_n16091_), .ZN(new_n16092_));
  AOI21_X1   g15795(.A1(new_n16092_), .A2(new_n16090_), .B(new_n16077_), .ZN(new_n16093_));
  INV_X1     g15796(.I(new_n16077_), .ZN(new_n16094_));
  XOR2_X1    g15797(.A1(new_n16084_), .A2(new_n16088_), .Z(new_n16095_));
  NOR2_X1    g15798(.A1(new_n16095_), .A2(new_n16094_), .ZN(new_n16096_));
  OAI22_X1   g15799(.A1(new_n970_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n820_), .ZN(new_n16097_));
  OAI21_X1   g15800(.A1(new_n10477_), .A2(new_n894_), .B(new_n16097_), .ZN(new_n16098_));
  AOI21_X1   g15801(.A1(new_n16098_), .A2(new_n827_), .B(new_n970_), .ZN(new_n16099_));
  XOR2_X1    g15802(.A1(new_n11298_), .A2(new_n16099_), .Z(new_n16100_));
  INV_X1     g15803(.I(new_n16100_), .ZN(new_n16101_));
  OAI21_X1   g15804(.A1(new_n16096_), .A2(new_n16093_), .B(new_n16101_), .ZN(new_n16102_));
  INV_X1     g15805(.I(new_n16090_), .ZN(new_n16103_));
  OAI21_X1   g15806(.A1(new_n16103_), .A2(new_n16091_), .B(new_n16094_), .ZN(new_n16104_));
  XOR2_X1    g15807(.A1(new_n16084_), .A2(new_n16089_), .Z(new_n16105_));
  NAND2_X1   g15808(.A1(new_n16105_), .A2(new_n16077_), .ZN(new_n16106_));
  NAND3_X1   g15809(.A1(new_n16106_), .A2(new_n16104_), .A3(new_n16100_), .ZN(new_n16107_));
  AOI21_X1   g15810(.A1(new_n16102_), .A2(new_n16107_), .B(new_n15841_), .ZN(new_n16108_));
  INV_X1     g15811(.I(new_n15841_), .ZN(new_n16109_));
  NAND3_X1   g15812(.A1(new_n16106_), .A2(new_n16104_), .A3(new_n16101_), .ZN(new_n16110_));
  OAI21_X1   g15813(.A1(new_n16096_), .A2(new_n16093_), .B(new_n16100_), .ZN(new_n16111_));
  AOI21_X1   g15814(.A1(new_n16111_), .A2(new_n16110_), .B(new_n16109_), .ZN(new_n16112_));
  NOR2_X1    g15815(.A1(new_n16108_), .A2(new_n16112_), .ZN(new_n16113_));
  INV_X1     g15816(.I(new_n16113_), .ZN(new_n16114_));
  NAND2_X1   g15817(.A1(new_n15743_), .A2(new_n15739_), .ZN(new_n16115_));
  OAI22_X1   g15818(.A1(new_n607_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n610_), .ZN(new_n16116_));
  OAI21_X1   g15819(.A1(new_n11744_), .A2(new_n684_), .B(new_n16116_), .ZN(new_n16117_));
  AOI21_X1   g15820(.A1(new_n16117_), .A2(new_n612_), .B(new_n607_), .ZN(new_n16118_));
  XNOR2_X1   g15821(.A1(new_n12546_), .A2(new_n16118_), .ZN(new_n16119_));
  AOI21_X1   g15822(.A1(new_n16115_), .A2(new_n15737_), .B(new_n16119_), .ZN(new_n16120_));
  NAND2_X1   g15823(.A1(new_n16115_), .A2(new_n15737_), .ZN(new_n16121_));
  INV_X1     g15824(.I(new_n16119_), .ZN(new_n16122_));
  NOR2_X1    g15825(.A1(new_n16121_), .A2(new_n16122_), .ZN(new_n16123_));
  OAI21_X1   g15826(.A1(new_n16123_), .A2(new_n16120_), .B(new_n16114_), .ZN(new_n16124_));
  NAND3_X1   g15827(.A1(new_n16115_), .A2(new_n15737_), .A3(new_n16122_), .ZN(new_n16125_));
  NAND2_X1   g15828(.A1(new_n16121_), .A2(new_n16119_), .ZN(new_n16126_));
  NAND2_X1   g15829(.A1(new_n16126_), .A2(new_n16125_), .ZN(new_n16127_));
  NAND2_X1   g15830(.A1(new_n16127_), .A2(new_n16113_), .ZN(new_n16128_));
  OAI22_X1   g15831(.A1(new_n448_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n450_), .ZN(new_n16129_));
  OAI21_X1   g15832(.A1(new_n12970_), .A2(new_n496_), .B(new_n16129_), .ZN(new_n16130_));
  AOI21_X1   g15833(.A1(new_n16130_), .A2(new_n452_), .B(new_n448_), .ZN(new_n16131_));
  XOR2_X1    g15834(.A1(new_n13784_), .A2(new_n16131_), .Z(new_n16132_));
  AOI21_X1   g15835(.A1(new_n16124_), .A2(new_n16128_), .B(new_n16132_), .ZN(new_n16133_));
  INV_X1     g15836(.I(new_n16133_), .ZN(new_n16134_));
  NAND3_X1   g15837(.A1(new_n16124_), .A2(new_n16128_), .A3(new_n16132_), .ZN(new_n16135_));
  AOI21_X1   g15838(.A1(new_n16134_), .A2(new_n16135_), .B(new_n15836_), .ZN(new_n16136_));
  INV_X1     g15839(.I(new_n15836_), .ZN(new_n16137_));
  INV_X1     g15840(.I(new_n16132_), .ZN(new_n16138_));
  NAND3_X1   g15841(.A1(new_n16124_), .A2(new_n16128_), .A3(new_n16138_), .ZN(new_n16139_));
  NOR2_X1    g15842(.A1(new_n16123_), .A2(new_n16120_), .ZN(new_n16140_));
  NOR2_X1    g15843(.A1(new_n16140_), .A2(new_n16113_), .ZN(new_n16141_));
  AOI21_X1   g15844(.A1(new_n16126_), .A2(new_n16125_), .B(new_n16114_), .ZN(new_n16142_));
  OAI21_X1   g15845(.A1(new_n16142_), .A2(new_n16141_), .B(new_n16132_), .ZN(new_n16143_));
  AOI21_X1   g15846(.A1(new_n16139_), .A2(new_n16143_), .B(new_n16137_), .ZN(new_n16144_));
  NOR2_X1    g15847(.A1(new_n16136_), .A2(new_n16144_), .ZN(new_n16145_));
  AOI21_X1   g15848(.A1(new_n15779_), .A2(new_n15777_), .B(new_n15792_), .ZN(new_n16146_));
  NOR2_X1    g15849(.A1(new_n366_), .A2(new_n404_), .ZN(new_n16147_));
  INV_X1     g15850(.I(new_n14596_), .ZN(new_n16148_));
  NAND2_X1   g15851(.A1(new_n16148_), .A2(new_n334_), .ZN(new_n16149_));
  OAI21_X1   g15852(.A1(new_n16147_), .A2(new_n16149_), .B(new_n340_), .ZN(new_n16150_));
  XNOR2_X1   g15853(.A1(new_n14978_), .A2(new_n16150_), .ZN(new_n16151_));
  INV_X1     g15854(.I(new_n16151_), .ZN(new_n16152_));
  NAND2_X1   g15855(.A1(new_n16146_), .A2(new_n16152_), .ZN(new_n16153_));
  NOR2_X1    g15856(.A1(new_n16146_), .A2(new_n16152_), .ZN(new_n16154_));
  INV_X1     g15857(.I(new_n16154_), .ZN(new_n16155_));
  AOI21_X1   g15858(.A1(new_n16155_), .A2(new_n16153_), .B(new_n16145_), .ZN(new_n16156_));
  INV_X1     g15859(.I(new_n16135_), .ZN(new_n16157_));
  OAI21_X1   g15860(.A1(new_n16157_), .A2(new_n16133_), .B(new_n16137_), .ZN(new_n16158_));
  AND2_X2    g15861(.A1(new_n16143_), .A2(new_n16139_), .Z(new_n16159_));
  OAI21_X1   g15862(.A1(new_n16159_), .A2(new_n16137_), .B(new_n16158_), .ZN(new_n16160_));
  NOR2_X1    g15863(.A1(new_n16146_), .A2(new_n16151_), .ZN(new_n16161_));
  INV_X1     g15864(.I(new_n16161_), .ZN(new_n16162_));
  NAND2_X1   g15865(.A1(new_n16146_), .A2(new_n16151_), .ZN(new_n16163_));
  AOI21_X1   g15866(.A1(new_n16163_), .A2(new_n16162_), .B(new_n16160_), .ZN(new_n16164_));
  NOR2_X1    g15867(.A1(new_n16164_), .A2(new_n16156_), .ZN(new_n16165_));
  NOR2_X1    g15868(.A1(new_n16165_), .A2(new_n15830_), .ZN(new_n16166_));
  XOR2_X1    g15869(.A1(new_n15827_), .A2(new_n16166_), .Z(new_n16167_));
  XOR2_X1    g15870(.A1(new_n16167_), .A2(new_n15814_), .Z(\f[67] ));
  NAND2_X1   g15871(.A1(new_n15807_), .A2(new_n15801_), .ZN(new_n16169_));
  AOI21_X1   g15872(.A1(new_n16169_), .A2(new_n15419_), .B(new_n15412_), .ZN(new_n16170_));
  NOR3_X1    g15873(.A1(new_n15820_), .A2(new_n15823_), .A3(new_n15419_), .ZN(new_n16171_));
  INV_X1     g15874(.I(new_n15814_), .ZN(new_n16172_));
  INV_X1     g15875(.I(new_n16153_), .ZN(new_n16173_));
  OAI21_X1   g15876(.A1(new_n16154_), .A2(new_n16173_), .B(new_n16160_), .ZN(new_n16174_));
  INV_X1     g15877(.I(new_n16163_), .ZN(new_n16175_));
  OAI21_X1   g15878(.A1(new_n16175_), .A2(new_n16161_), .B(new_n16145_), .ZN(new_n16176_));
  NAND3_X1   g15879(.A1(new_n15830_), .A2(new_n16174_), .A3(new_n16176_), .ZN(new_n16177_));
  NAND2_X1   g15880(.A1(new_n16172_), .A2(new_n16177_), .ZN(new_n16178_));
  NOR4_X1    g15881(.A1(new_n16170_), .A2(new_n15022_), .A3(new_n16178_), .A4(new_n16171_), .ZN(new_n16179_));
  NOR2_X1    g15882(.A1(new_n16179_), .A2(new_n16166_), .ZN(new_n16180_));
  INV_X1     g15883(.I(new_n16180_), .ZN(new_n16181_));
  AOI21_X1   g15884(.A1(new_n16160_), .A2(new_n16163_), .B(new_n16161_), .ZN(new_n16182_));
  INV_X1     g15885(.I(new_n16182_), .ZN(new_n16183_));
  AOI21_X1   g15886(.A1(new_n16106_), .A2(new_n16104_), .B(new_n16100_), .ZN(new_n16184_));
  AOI21_X1   g15887(.A1(new_n16109_), .A2(new_n16107_), .B(new_n16184_), .ZN(new_n16185_));
  NOR2_X1    g15888(.A1(new_n16091_), .A2(new_n16077_), .ZN(new_n16186_));
  NOR2_X1    g15889(.A1(new_n16186_), .A2(new_n16103_), .ZN(new_n16187_));
  NOR2_X1    g15890(.A1(new_n16073_), .A2(new_n15846_), .ZN(new_n16188_));
  NOR2_X1    g15891(.A1(new_n16188_), .A2(new_n16070_), .ZN(new_n16189_));
  INV_X1     g15892(.I(new_n16189_), .ZN(new_n16190_));
  NOR2_X1    g15893(.A1(new_n16061_), .A2(new_n15851_), .ZN(new_n16191_));
  NOR2_X1    g15894(.A1(new_n16191_), .A2(new_n16054_), .ZN(new_n16192_));
  NOR2_X1    g15895(.A1(new_n16055_), .A2(new_n15858_), .ZN(new_n16193_));
  NOR2_X1    g15896(.A1(new_n16029_), .A2(new_n16031_), .ZN(new_n16194_));
  NOR2_X1    g15897(.A1(new_n16002_), .A2(new_n16006_), .ZN(new_n16195_));
  AOI21_X1   g15898(.A1(new_n16016_), .A2(new_n16018_), .B(new_n16195_), .ZN(new_n16196_));
  AOI21_X1   g15899(.A1(new_n15998_), .A2(new_n15996_), .B(new_n15994_), .ZN(new_n16197_));
  INV_X1     g15900(.I(new_n16197_), .ZN(new_n16198_));
  NAND2_X1   g15901(.A1(new_n15976_), .A2(new_n15983_), .ZN(new_n16199_));
  OAI21_X1   g15902(.A1(new_n15976_), .A2(new_n15983_), .B(new_n15865_), .ZN(new_n16200_));
  NAND2_X1   g15903(.A1(new_n16200_), .A2(new_n16199_), .ZN(new_n16201_));
  NAND2_X1   g15904(.A1(new_n15971_), .A2(new_n15973_), .ZN(new_n16202_));
  NAND2_X1   g15905(.A1(new_n16202_), .A2(new_n15968_), .ZN(new_n16203_));
  INV_X1     g15906(.I(new_n16203_), .ZN(new_n16204_));
  AOI21_X1   g15907(.A1(new_n15870_), .A2(new_n15958_), .B(new_n15957_), .ZN(new_n16205_));
  INV_X1     g15908(.I(new_n16205_), .ZN(new_n16206_));
  AOI21_X1   g15909(.A1(new_n15937_), .A2(new_n15933_), .B(new_n15932_), .ZN(new_n16207_));
  NAND2_X1   g15910(.A1(new_n15922_), .A2(new_n15924_), .ZN(new_n16208_));
  AND2_X2    g15911(.A1(new_n16208_), .A2(new_n15919_), .Z(new_n16209_));
  INV_X1     g15912(.I(new_n16209_), .ZN(new_n16210_));
  NOR2_X1    g15913(.A1(new_n15914_), .A2(new_n15912_), .ZN(new_n16211_));
  AOI22_X1   g15914(.A1(new_n10969_), .A2(new_n932_), .B1(new_n11394_), .B2(\b[12] ), .ZN(new_n16212_));
  OAI21_X1   g15915(.A1(new_n16212_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n16213_));
  XOR2_X1    g15916(.A1(new_n937_), .A2(new_n16213_), .Z(new_n16214_));
  INV_X1     g15917(.I(new_n16214_), .ZN(new_n16215_));
  OAI22_X1   g15918(.A1(new_n13880_), .A2(new_n516_), .B1(new_n420_), .B2(new_n13885_), .ZN(new_n16216_));
  AOI21_X1   g15919(.A1(new_n16216_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n16217_));
  XOR2_X1    g15920(.A1(new_n522_), .A2(new_n16217_), .Z(new_n16218_));
  NOR2_X1    g15921(.A1(new_n13476_), .A2(new_n325_), .ZN(new_n16219_));
  XOR2_X1    g15922(.A1(new_n14736_), .A2(new_n325_), .Z(new_n16220_));
  NAND2_X1   g15923(.A1(new_n16220_), .A2(\b[5] ), .ZN(new_n16221_));
  XOR2_X1    g15924(.A1(new_n16221_), .A2(new_n16219_), .Z(new_n16222_));
  INV_X1     g15925(.I(new_n16222_), .ZN(new_n16223_));
  NOR2_X1    g15926(.A1(new_n16223_), .A2(new_n260_), .ZN(new_n16224_));
  NOR2_X1    g15927(.A1(new_n16222_), .A2(\a[2] ), .ZN(new_n16225_));
  NOR2_X1    g15928(.A1(new_n16224_), .A2(new_n16225_), .ZN(new_n16226_));
  INV_X1     g15929(.I(new_n16226_), .ZN(new_n16227_));
  XOR2_X1    g15930(.A1(new_n16222_), .A2(new_n260_), .Z(new_n16228_));
  NOR2_X1    g15931(.A1(new_n16218_), .A2(new_n16228_), .ZN(new_n16229_));
  AOI21_X1   g15932(.A1(new_n16218_), .A2(new_n16227_), .B(new_n16229_), .ZN(new_n16230_));
  INV_X1     g15933(.I(new_n16230_), .ZN(new_n16231_));
  NOR2_X1    g15934(.A1(new_n15880_), .A2(new_n15885_), .ZN(new_n16232_));
  NOR2_X1    g15935(.A1(new_n16232_), .A2(new_n15886_), .ZN(new_n16233_));
  AOI22_X1   g15936(.A1(new_n13078_), .A2(\b[9] ), .B1(new_n773_), .B2(new_n12218_), .ZN(new_n16234_));
  OAI21_X1   g15937(.A1(new_n16234_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n16235_));
  XOR2_X1    g15938(.A1(new_n710_), .A2(new_n16235_), .Z(new_n16236_));
  XOR2_X1    g15939(.A1(new_n16236_), .A2(new_n16233_), .Z(new_n16237_));
  NAND2_X1   g15940(.A1(new_n16237_), .A2(new_n16231_), .ZN(new_n16238_));
  NOR2_X1    g15941(.A1(new_n16236_), .A2(new_n16233_), .ZN(new_n16239_));
  AND2_X2    g15942(.A1(new_n16236_), .A2(new_n16233_), .Z(new_n16240_));
  OAI21_X1   g15943(.A1(new_n16240_), .A2(new_n16239_), .B(new_n16230_), .ZN(new_n16241_));
  NAND2_X1   g15944(.A1(new_n16238_), .A2(new_n16241_), .ZN(new_n16242_));
  NOR2_X1    g15945(.A1(new_n15899_), .A2(new_n15891_), .ZN(new_n16243_));
  NOR2_X1    g15946(.A1(new_n16243_), .A2(new_n15898_), .ZN(new_n16244_));
  NOR2_X1    g15947(.A1(new_n16242_), .A2(new_n16244_), .ZN(new_n16245_));
  AND2_X2    g15948(.A1(new_n16242_), .A2(new_n16244_), .Z(new_n16246_));
  OAI21_X1   g15949(.A1(new_n16246_), .A2(new_n16245_), .B(new_n16215_), .ZN(new_n16247_));
  XOR2_X1    g15950(.A1(new_n16242_), .A2(new_n16244_), .Z(new_n16248_));
  NAND2_X1   g15951(.A1(new_n16248_), .A2(new_n16214_), .ZN(new_n16249_));
  NAND2_X1   g15952(.A1(new_n16249_), .A2(new_n16247_), .ZN(new_n16250_));
  AOI22_X1   g15953(.A1(new_n11415_), .A2(new_n1292_), .B1(\b[15] ), .B2(new_n10145_), .ZN(new_n16251_));
  OAI21_X1   g15954(.A1(new_n16251_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n16252_));
  XOR2_X1    g15955(.A1(new_n1196_), .A2(new_n16252_), .Z(new_n16253_));
  INV_X1     g15956(.I(new_n16253_), .ZN(new_n16254_));
  NAND2_X1   g15957(.A1(new_n16250_), .A2(new_n16254_), .ZN(new_n16255_));
  INV_X1     g15958(.I(new_n16255_), .ZN(new_n16256_));
  NOR2_X1    g15959(.A1(new_n16250_), .A2(new_n16254_), .ZN(new_n16257_));
  OAI22_X1   g15960(.A1(new_n16256_), .A2(new_n16257_), .B1(new_n15913_), .B2(new_n16211_), .ZN(new_n16258_));
  NOR2_X1    g15961(.A1(new_n16211_), .A2(new_n15913_), .ZN(new_n16259_));
  XOR2_X1    g15962(.A1(new_n16250_), .A2(new_n16254_), .Z(new_n16260_));
  NAND2_X1   g15963(.A1(new_n16260_), .A2(new_n16259_), .ZN(new_n16261_));
  NAND2_X1   g15964(.A1(new_n16261_), .A2(new_n16258_), .ZN(new_n16262_));
  OAI22_X1   g15965(.A1(new_n8644_), .A2(new_n1518_), .B1(new_n1525_), .B2(new_n9388_), .ZN(new_n16263_));
  OAI21_X1   g15966(.A1(new_n1294_), .A2(new_n10154_), .B(new_n16263_), .ZN(new_n16264_));
  AOI21_X1   g15967(.A1(new_n16264_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n16265_));
  XOR2_X1    g15968(.A1(new_n1530_), .A2(new_n16265_), .Z(new_n16266_));
  INV_X1     g15969(.I(new_n16266_), .ZN(new_n16267_));
  XOR2_X1    g15970(.A1(new_n16262_), .A2(new_n16267_), .Z(new_n16268_));
  NAND2_X1   g15971(.A1(new_n16268_), .A2(new_n16210_), .ZN(new_n16269_));
  NAND2_X1   g15972(.A1(new_n16262_), .A2(new_n16267_), .ZN(new_n16270_));
  INV_X1     g15973(.I(new_n16270_), .ZN(new_n16271_));
  NOR2_X1    g15974(.A1(new_n16262_), .A2(new_n16267_), .ZN(new_n16272_));
  OAI21_X1   g15975(.A1(new_n16271_), .A2(new_n16272_), .B(new_n16209_), .ZN(new_n16273_));
  OAI22_X1   g15976(.A1(new_n7619_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n8309_), .ZN(new_n16274_));
  OAI21_X1   g15977(.A1(new_n1634_), .A2(new_n7947_), .B(new_n16274_), .ZN(new_n16275_));
  AOI21_X1   g15978(.A1(new_n16275_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n16276_));
  XNOR2_X1   g15979(.A1(new_n1940_), .A2(new_n16276_), .ZN(new_n16277_));
  INV_X1     g15980(.I(new_n16277_), .ZN(new_n16278_));
  NAND3_X1   g15981(.A1(new_n16269_), .A2(new_n16273_), .A3(new_n16278_), .ZN(new_n16279_));
  NAND2_X1   g15982(.A1(new_n16269_), .A2(new_n16273_), .ZN(new_n16280_));
  NAND2_X1   g15983(.A1(new_n16280_), .A2(new_n16277_), .ZN(new_n16281_));
  AOI21_X1   g15984(.A1(new_n16281_), .A2(new_n16279_), .B(new_n16207_), .ZN(new_n16282_));
  INV_X1     g15985(.I(new_n16207_), .ZN(new_n16283_));
  XOR2_X1    g15986(.A1(new_n16280_), .A2(new_n16278_), .Z(new_n16284_));
  NOR2_X1    g15987(.A1(new_n16284_), .A2(new_n16283_), .ZN(new_n16285_));
  NOR2_X1    g15988(.A1(new_n16285_), .A2(new_n16282_), .ZN(new_n16286_));
  AOI21_X1   g15989(.A1(new_n15949_), .A2(new_n15947_), .B(new_n15945_), .ZN(new_n16287_));
  OAI22_X1   g15990(.A1(new_n6644_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n6647_), .ZN(new_n16288_));
  OAI21_X1   g15991(.A1(new_n2102_), .A2(new_n7284_), .B(new_n16288_), .ZN(new_n16289_));
  AOI21_X1   g15992(.A1(new_n2443_), .A2(new_n6631_), .B(new_n16289_), .ZN(new_n16290_));
  XNOR2_X1   g15993(.A1(new_n16287_), .A2(new_n16290_), .ZN(new_n16291_));
  NAND2_X1   g15994(.A1(new_n16291_), .A2(new_n16286_), .ZN(new_n16292_));
  INV_X1     g15995(.I(new_n16286_), .ZN(new_n16293_));
  XOR2_X1    g15996(.A1(new_n16287_), .A2(new_n16290_), .Z(new_n16294_));
  NAND2_X1   g15997(.A1(new_n16294_), .A2(new_n16293_), .ZN(new_n16295_));
  AOI21_X1   g15998(.A1(new_n16295_), .A2(new_n16292_), .B(\a[44] ), .ZN(new_n16296_));
  INV_X1     g15999(.I(new_n16296_), .ZN(new_n16297_));
  NAND3_X1   g16000(.A1(new_n16295_), .A2(new_n16292_), .A3(\a[44] ), .ZN(new_n16298_));
  OAI22_X1   g16001(.A1(new_n5993_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n5991_), .ZN(new_n16299_));
  OAI21_X1   g16002(.A1(new_n2643_), .A2(new_n5997_), .B(new_n16299_), .ZN(new_n16300_));
  AOI21_X1   g16003(.A1(new_n16300_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n16301_));
  XNOR2_X1   g16004(.A1(new_n3022_), .A2(new_n16301_), .ZN(new_n16302_));
  AOI21_X1   g16005(.A1(new_n16297_), .A2(new_n16298_), .B(new_n16302_), .ZN(new_n16303_));
  NAND3_X1   g16006(.A1(new_n16297_), .A2(new_n16298_), .A3(new_n16302_), .ZN(new_n16304_));
  INV_X1     g16007(.I(new_n16304_), .ZN(new_n16305_));
  OAI21_X1   g16008(.A1(new_n16305_), .A2(new_n16303_), .B(new_n16206_), .ZN(new_n16306_));
  INV_X1     g16009(.I(new_n16302_), .ZN(new_n16307_));
  NAND3_X1   g16010(.A1(new_n16297_), .A2(new_n16298_), .A3(new_n16307_), .ZN(new_n16308_));
  INV_X1     g16011(.I(new_n16308_), .ZN(new_n16309_));
  AOI21_X1   g16012(.A1(new_n16297_), .A2(new_n16298_), .B(new_n16307_), .ZN(new_n16310_));
  OAI21_X1   g16013(.A1(new_n16309_), .A2(new_n16310_), .B(new_n16205_), .ZN(new_n16311_));
  OAI22_X1   g16014(.A1(new_n5420_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n5107_), .ZN(new_n16312_));
  OAI21_X1   g16015(.A1(new_n3260_), .A2(new_n5112_), .B(new_n16312_), .ZN(new_n16313_));
  AOI21_X1   g16016(.A1(new_n16313_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n16314_));
  XOR2_X1    g16017(.A1(new_n3722_), .A2(new_n16314_), .Z(new_n16315_));
  INV_X1     g16018(.I(new_n16315_), .ZN(new_n16316_));
  NAND3_X1   g16019(.A1(new_n16306_), .A2(new_n16311_), .A3(new_n16316_), .ZN(new_n16317_));
  INV_X1     g16020(.I(new_n16303_), .ZN(new_n16318_));
  AOI21_X1   g16021(.A1(new_n16318_), .A2(new_n16304_), .B(new_n16205_), .ZN(new_n16319_));
  INV_X1     g16022(.I(new_n16310_), .ZN(new_n16320_));
  AOI21_X1   g16023(.A1(new_n16320_), .A2(new_n16308_), .B(new_n16206_), .ZN(new_n16321_));
  OAI21_X1   g16024(.A1(new_n16319_), .A2(new_n16321_), .B(new_n16315_), .ZN(new_n16322_));
  AOI21_X1   g16025(.A1(new_n16322_), .A2(new_n16317_), .B(new_n16204_), .ZN(new_n16323_));
  AOI21_X1   g16026(.A1(new_n16306_), .A2(new_n16311_), .B(new_n16315_), .ZN(new_n16324_));
  INV_X1     g16027(.I(new_n16324_), .ZN(new_n16325_));
  NAND3_X1   g16028(.A1(new_n16306_), .A2(new_n16311_), .A3(new_n16315_), .ZN(new_n16326_));
  AOI21_X1   g16029(.A1(new_n16325_), .A2(new_n16326_), .B(new_n16203_), .ZN(new_n16327_));
  OAI22_X1   g16030(.A1(new_n4072_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n4067_), .ZN(new_n16328_));
  OAI21_X1   g16031(.A1(new_n3989_), .A2(new_n4318_), .B(new_n16328_), .ZN(new_n16329_));
  AOI21_X1   g16032(.A1(new_n16329_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n16330_));
  XOR2_X1    g16033(.A1(new_n4499_), .A2(new_n16330_), .Z(new_n16331_));
  NOR3_X1    g16034(.A1(new_n16327_), .A2(new_n16323_), .A3(new_n16331_), .ZN(new_n16332_));
  NOR3_X1    g16035(.A1(new_n16319_), .A2(new_n16321_), .A3(new_n16315_), .ZN(new_n16333_));
  AOI21_X1   g16036(.A1(new_n16306_), .A2(new_n16311_), .B(new_n16316_), .ZN(new_n16334_));
  OAI21_X1   g16037(.A1(new_n16333_), .A2(new_n16334_), .B(new_n16203_), .ZN(new_n16335_));
  NOR3_X1    g16038(.A1(new_n16319_), .A2(new_n16321_), .A3(new_n16316_), .ZN(new_n16336_));
  OAI21_X1   g16039(.A1(new_n16324_), .A2(new_n16336_), .B(new_n16204_), .ZN(new_n16337_));
  INV_X1     g16040(.I(new_n16331_), .ZN(new_n16338_));
  AOI21_X1   g16041(.A1(new_n16337_), .A2(new_n16335_), .B(new_n16338_), .ZN(new_n16339_));
  OAI21_X1   g16042(.A1(new_n16332_), .A2(new_n16339_), .B(new_n16201_), .ZN(new_n16340_));
  OAI21_X1   g16043(.A1(new_n16327_), .A2(new_n16323_), .B(new_n16338_), .ZN(new_n16341_));
  NAND3_X1   g16044(.A1(new_n16337_), .A2(new_n16335_), .A3(new_n16331_), .ZN(new_n16342_));
  NAND2_X1   g16045(.A1(new_n16341_), .A2(new_n16342_), .ZN(new_n16343_));
  NAND3_X1   g16046(.A1(new_n16343_), .A2(new_n16199_), .A3(new_n16200_), .ZN(new_n16344_));
  NAND2_X1   g16047(.A1(new_n16344_), .A2(new_n16340_), .ZN(new_n16345_));
  OAI22_X1   g16048(.A1(new_n5068_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n5353_), .ZN(new_n16346_));
  OAI21_X1   g16049(.A1(new_n4774_), .A2(new_n3569_), .B(new_n16346_), .ZN(new_n16347_));
  AOI21_X1   g16050(.A1(new_n16347_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n16348_));
  XNOR2_X1   g16051(.A1(new_n5357_), .A2(new_n16348_), .ZN(new_n16349_));
  INV_X1     g16052(.I(new_n16349_), .ZN(new_n16350_));
  NAND2_X1   g16053(.A1(new_n16345_), .A2(new_n16350_), .ZN(new_n16351_));
  NAND3_X1   g16054(.A1(new_n16344_), .A2(new_n16340_), .A3(new_n16349_), .ZN(new_n16352_));
  NAND2_X1   g16055(.A1(new_n16351_), .A2(new_n16352_), .ZN(new_n16353_));
  NAND2_X1   g16056(.A1(new_n16353_), .A2(new_n16198_), .ZN(new_n16354_));
  NAND3_X1   g16057(.A1(new_n16344_), .A2(new_n16340_), .A3(new_n16350_), .ZN(new_n16355_));
  NAND2_X1   g16058(.A1(new_n16345_), .A2(new_n16349_), .ZN(new_n16356_));
  NAND2_X1   g16059(.A1(new_n16356_), .A2(new_n16355_), .ZN(new_n16357_));
  NAND2_X1   g16060(.A1(new_n16357_), .A2(new_n16197_), .ZN(new_n16358_));
  OAI22_X1   g16061(.A1(new_n5921_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n6229_), .ZN(new_n16359_));
  OAI21_X1   g16062(.A1(new_n5913_), .A2(new_n2884_), .B(new_n16359_), .ZN(new_n16360_));
  AOI21_X1   g16063(.A1(new_n16360_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n16361_));
  XOR2_X1    g16064(.A1(new_n6233_), .A2(new_n16361_), .Z(new_n16362_));
  AOI21_X1   g16065(.A1(new_n16354_), .A2(new_n16358_), .B(new_n16362_), .ZN(new_n16363_));
  AOI21_X1   g16066(.A1(new_n16351_), .A2(new_n16352_), .B(new_n16197_), .ZN(new_n16364_));
  AOI21_X1   g16067(.A1(new_n16355_), .A2(new_n16356_), .B(new_n16198_), .ZN(new_n16365_));
  INV_X1     g16068(.I(new_n16362_), .ZN(new_n16366_));
  NOR3_X1    g16069(.A1(new_n16365_), .A2(new_n16364_), .A3(new_n16366_), .ZN(new_n16367_));
  NOR2_X1    g16070(.A1(new_n16367_), .A2(new_n16363_), .ZN(new_n16368_));
  NOR2_X1    g16071(.A1(new_n16368_), .A2(new_n16196_), .ZN(new_n16369_));
  NAND2_X1   g16072(.A1(new_n16018_), .A2(new_n16016_), .ZN(new_n16370_));
  NAND2_X1   g16073(.A1(new_n16370_), .A2(new_n16017_), .ZN(new_n16371_));
  NOR3_X1    g16074(.A1(new_n16365_), .A2(new_n16364_), .A3(new_n16362_), .ZN(new_n16372_));
  AOI21_X1   g16075(.A1(new_n16358_), .A2(new_n16354_), .B(new_n16366_), .ZN(new_n16373_));
  NOR2_X1    g16076(.A1(new_n16372_), .A2(new_n16373_), .ZN(new_n16374_));
  NOR2_X1    g16077(.A1(new_n16374_), .A2(new_n16371_), .ZN(new_n16375_));
  OAI22_X1   g16078(.A1(new_n2171_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n2166_), .ZN(new_n16376_));
  OAI21_X1   g16079(.A1(new_n6538_), .A2(new_n2322_), .B(new_n16376_), .ZN(new_n16377_));
  AOI21_X1   g16080(.A1(new_n16377_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n16378_));
  XNOR2_X1   g16081(.A1(new_n7202_), .A2(new_n16378_), .ZN(new_n16379_));
  INV_X1     g16082(.I(new_n16379_), .ZN(new_n16380_));
  OAI21_X1   g16083(.A1(new_n16369_), .A2(new_n16375_), .B(new_n16380_), .ZN(new_n16381_));
  OAI21_X1   g16084(.A1(new_n16363_), .A2(new_n16367_), .B(new_n16371_), .ZN(new_n16382_));
  OAI21_X1   g16085(.A1(new_n16372_), .A2(new_n16373_), .B(new_n16196_), .ZN(new_n16383_));
  NAND3_X1   g16086(.A1(new_n16383_), .A2(new_n16382_), .A3(new_n16379_), .ZN(new_n16384_));
  NAND2_X1   g16087(.A1(new_n16384_), .A2(new_n16381_), .ZN(new_n16385_));
  OAI21_X1   g16088(.A1(new_n16194_), .A2(new_n16024_), .B(new_n16385_), .ZN(new_n16386_));
  NOR2_X1    g16089(.A1(new_n16194_), .A2(new_n16024_), .ZN(new_n16387_));
  NAND3_X1   g16090(.A1(new_n16383_), .A2(new_n16382_), .A3(new_n16380_), .ZN(new_n16388_));
  OAI21_X1   g16091(.A1(new_n16369_), .A2(new_n16375_), .B(new_n16379_), .ZN(new_n16389_));
  NAND2_X1   g16092(.A1(new_n16388_), .A2(new_n16389_), .ZN(new_n16390_));
  NAND2_X1   g16093(.A1(new_n16387_), .A2(new_n16390_), .ZN(new_n16391_));
  OAI22_X1   g16094(.A1(new_n1712_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n1707_), .ZN(new_n16392_));
  OAI21_X1   g16095(.A1(new_n7864_), .A2(new_n1850_), .B(new_n16392_), .ZN(new_n16393_));
  AOI21_X1   g16096(.A1(new_n16393_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n16394_));
  XOR2_X1    g16097(.A1(new_n8217_), .A2(new_n16394_), .Z(new_n16395_));
  AOI21_X1   g16098(.A1(new_n16386_), .A2(new_n16391_), .B(new_n16395_), .ZN(new_n16396_));
  AOI21_X1   g16099(.A1(new_n16381_), .A2(new_n16384_), .B(new_n16387_), .ZN(new_n16397_));
  NOR3_X1    g16100(.A1(new_n16369_), .A2(new_n16375_), .A3(new_n16379_), .ZN(new_n16398_));
  AOI21_X1   g16101(.A1(new_n16383_), .A2(new_n16382_), .B(new_n16380_), .ZN(new_n16399_));
  NOR2_X1    g16102(.A1(new_n16399_), .A2(new_n16398_), .ZN(new_n16400_));
  NOR3_X1    g16103(.A1(new_n16400_), .A2(new_n16024_), .A3(new_n16194_), .ZN(new_n16401_));
  INV_X1     g16104(.I(new_n16395_), .ZN(new_n16402_));
  NOR3_X1    g16105(.A1(new_n16397_), .A2(new_n16401_), .A3(new_n16402_), .ZN(new_n16403_));
  OAI22_X1   g16106(.A1(new_n16403_), .A2(new_n16396_), .B1(new_n16193_), .B2(new_n16039_), .ZN(new_n16404_));
  NOR2_X1    g16107(.A1(new_n16193_), .A2(new_n16039_), .ZN(new_n16405_));
  NAND3_X1   g16108(.A1(new_n16386_), .A2(new_n16391_), .A3(new_n16402_), .ZN(new_n16406_));
  OAI21_X1   g16109(.A1(new_n16397_), .A2(new_n16401_), .B(new_n16395_), .ZN(new_n16407_));
  NAND2_X1   g16110(.A1(new_n16407_), .A2(new_n16406_), .ZN(new_n16408_));
  NAND2_X1   g16111(.A1(new_n16408_), .A2(new_n16405_), .ZN(new_n16409_));
  OAI22_X1   g16112(.A1(new_n1347_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n1344_), .ZN(new_n16410_));
  OAI21_X1   g16113(.A1(new_n8563_), .A2(new_n1457_), .B(new_n16410_), .ZN(new_n16411_));
  AOI21_X1   g16114(.A1(new_n16411_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n16412_));
  XNOR2_X1   g16115(.A1(new_n9299_), .A2(new_n16412_), .ZN(new_n16413_));
  AOI21_X1   g16116(.A1(new_n16409_), .A2(new_n16404_), .B(new_n16413_), .ZN(new_n16414_));
  NAND2_X1   g16117(.A1(new_n16409_), .A2(new_n16404_), .ZN(new_n16415_));
  INV_X1     g16118(.I(new_n16413_), .ZN(new_n16416_));
  NOR2_X1    g16119(.A1(new_n16415_), .A2(new_n16416_), .ZN(new_n16417_));
  NOR2_X1    g16120(.A1(new_n16417_), .A2(new_n16414_), .ZN(new_n16418_));
  NOR2_X1    g16121(.A1(new_n16418_), .A2(new_n16192_), .ZN(new_n16419_));
  INV_X1     g16122(.I(new_n16054_), .ZN(new_n16420_));
  OAI21_X1   g16123(.A1(new_n15851_), .A2(new_n16061_), .B(new_n16420_), .ZN(new_n16421_));
  NAND3_X1   g16124(.A1(new_n16409_), .A2(new_n16404_), .A3(new_n16416_), .ZN(new_n16422_));
  NAND2_X1   g16125(.A1(new_n16415_), .A2(new_n16413_), .ZN(new_n16423_));
  AOI21_X1   g16126(.A1(new_n16422_), .A2(new_n16423_), .B(new_n16421_), .ZN(new_n16424_));
  NOR2_X1    g16127(.A1(new_n16419_), .A2(new_n16424_), .ZN(new_n16425_));
  OAI22_X1   g16128(.A1(new_n1055_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n1061_), .ZN(new_n16426_));
  OAI21_X1   g16129(.A1(new_n10025_), .A2(new_n1332_), .B(new_n16426_), .ZN(new_n16427_));
  AOI21_X1   g16130(.A1(new_n16427_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n16428_));
  XOR2_X1    g16131(.A1(new_n10476_), .A2(new_n16428_), .Z(new_n16429_));
  NOR2_X1    g16132(.A1(new_n16425_), .A2(new_n16429_), .ZN(new_n16430_));
  INV_X1     g16133(.I(new_n16429_), .ZN(new_n16431_));
  NOR3_X1    g16134(.A1(new_n16419_), .A2(new_n16424_), .A3(new_n16431_), .ZN(new_n16432_));
  OAI21_X1   g16135(.A1(new_n16430_), .A2(new_n16432_), .B(new_n16190_), .ZN(new_n16433_));
  NOR3_X1    g16136(.A1(new_n16419_), .A2(new_n16424_), .A3(new_n16429_), .ZN(new_n16434_));
  NOR2_X1    g16137(.A1(new_n16425_), .A2(new_n16431_), .ZN(new_n16435_));
  OAI21_X1   g16138(.A1(new_n16435_), .A2(new_n16434_), .B(new_n16189_), .ZN(new_n16436_));
  OAI22_X1   g16139(.A1(new_n970_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n820_), .ZN(new_n16437_));
  OAI21_X1   g16140(.A1(new_n10862_), .A2(new_n894_), .B(new_n16437_), .ZN(new_n16438_));
  AOI21_X1   g16141(.A1(new_n16438_), .A2(new_n827_), .B(new_n970_), .ZN(new_n16439_));
  XNOR2_X1   g16142(.A1(new_n11748_), .A2(new_n16439_), .ZN(new_n16440_));
  AOI21_X1   g16143(.A1(new_n16433_), .A2(new_n16436_), .B(new_n16440_), .ZN(new_n16441_));
  INV_X1     g16144(.I(new_n16441_), .ZN(new_n16442_));
  NAND3_X1   g16145(.A1(new_n16433_), .A2(new_n16436_), .A3(new_n16440_), .ZN(new_n16443_));
  AOI21_X1   g16146(.A1(new_n16442_), .A2(new_n16443_), .B(new_n16187_), .ZN(new_n16444_));
  NOR2_X1    g16147(.A1(new_n16430_), .A2(new_n16432_), .ZN(new_n16445_));
  NOR2_X1    g16148(.A1(new_n16445_), .A2(new_n16189_), .ZN(new_n16446_));
  INV_X1     g16149(.I(new_n16436_), .ZN(new_n16447_));
  NOR3_X1    g16150(.A1(new_n16446_), .A2(new_n16447_), .A3(new_n16440_), .ZN(new_n16448_));
  INV_X1     g16151(.I(new_n16440_), .ZN(new_n16449_));
  AOI21_X1   g16152(.A1(new_n16433_), .A2(new_n16436_), .B(new_n16449_), .ZN(new_n16450_));
  NOR2_X1    g16153(.A1(new_n16448_), .A2(new_n16450_), .ZN(new_n16451_));
  NOR3_X1    g16154(.A1(new_n16451_), .A2(new_n16103_), .A3(new_n16186_), .ZN(new_n16452_));
  OAI22_X1   g16155(.A1(new_n607_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n610_), .ZN(new_n16453_));
  OAI21_X1   g16156(.A1(new_n12536_), .A2(new_n684_), .B(new_n16453_), .ZN(new_n16454_));
  AOI21_X1   g16157(.A1(new_n16454_), .A2(new_n612_), .B(new_n607_), .ZN(new_n16455_));
  XOR2_X1    g16158(.A1(new_n12969_), .A2(new_n16455_), .Z(new_n16456_));
  INV_X1     g16159(.I(new_n16456_), .ZN(new_n16457_));
  OAI21_X1   g16160(.A1(new_n16452_), .A2(new_n16444_), .B(new_n16457_), .ZN(new_n16458_));
  NOR3_X1    g16161(.A1(new_n16452_), .A2(new_n16444_), .A3(new_n16457_), .ZN(new_n16459_));
  INV_X1     g16162(.I(new_n16459_), .ZN(new_n16460_));
  AOI21_X1   g16163(.A1(new_n16460_), .A2(new_n16458_), .B(new_n16185_), .ZN(new_n16461_));
  NAND2_X1   g16164(.A1(new_n16107_), .A2(new_n16109_), .ZN(new_n16462_));
  NAND2_X1   g16165(.A1(new_n16462_), .A2(new_n16102_), .ZN(new_n16463_));
  NOR2_X1    g16166(.A1(new_n16452_), .A2(new_n16444_), .ZN(new_n16464_));
  XOR2_X1    g16167(.A1(new_n16464_), .A2(new_n16457_), .Z(new_n16465_));
  NOR2_X1    g16168(.A1(new_n16465_), .A2(new_n16463_), .ZN(new_n16466_));
  NOR2_X1    g16169(.A1(new_n16466_), .A2(new_n16461_), .ZN(new_n16467_));
  NOR2_X1    g16170(.A1(new_n16123_), .A2(new_n16113_), .ZN(new_n16468_));
  OAI22_X1   g16171(.A1(new_n448_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n450_), .ZN(new_n16469_));
  OAI21_X1   g16172(.A1(new_n13367_), .A2(new_n496_), .B(new_n16469_), .ZN(new_n16470_));
  AOI21_X1   g16173(.A1(new_n16470_), .A2(new_n452_), .B(new_n448_), .ZN(new_n16471_));
  XOR2_X1    g16174(.A1(new_n14213_), .A2(new_n16471_), .Z(new_n16472_));
  NOR3_X1    g16175(.A1(new_n16468_), .A2(new_n16120_), .A3(new_n16472_), .ZN(new_n16473_));
  INV_X1     g16176(.I(new_n16473_), .ZN(new_n16474_));
  OAI21_X1   g16177(.A1(new_n16468_), .A2(new_n16120_), .B(new_n16472_), .ZN(new_n16475_));
  AOI21_X1   g16178(.A1(new_n16474_), .A2(new_n16475_), .B(new_n16467_), .ZN(new_n16476_));
  INV_X1     g16179(.I(new_n16461_), .ZN(new_n16477_));
  OAI21_X1   g16180(.A1(new_n16465_), .A2(new_n16463_), .B(new_n16477_), .ZN(new_n16478_));
  INV_X1     g16181(.I(new_n16472_), .ZN(new_n16479_));
  OAI21_X1   g16182(.A1(new_n16468_), .A2(new_n16120_), .B(new_n16479_), .ZN(new_n16480_));
  NOR2_X1    g16183(.A1(new_n16468_), .A2(new_n16120_), .ZN(new_n16481_));
  NAND2_X1   g16184(.A1(new_n16481_), .A2(new_n16472_), .ZN(new_n16482_));
  AOI21_X1   g16185(.A1(new_n16482_), .A2(new_n16480_), .B(new_n16478_), .ZN(new_n16483_));
  NOR2_X1    g16186(.A1(new_n16476_), .A2(new_n16483_), .ZN(new_n16484_));
  AOI21_X1   g16187(.A1(new_n16137_), .A2(new_n16135_), .B(new_n16133_), .ZN(new_n16485_));
  NOR2_X1    g16188(.A1(new_n15397_), .A2(new_n14592_), .ZN(new_n16486_));
  INV_X1     g16189(.I(new_n16486_), .ZN(new_n16487_));
  OAI21_X1   g16190(.A1(new_n341_), .A2(new_n366_), .B(new_n16487_), .ZN(new_n16488_));
  NAND2_X1   g16191(.A1(new_n16485_), .A2(new_n16488_), .ZN(new_n16489_));
  INV_X1     g16192(.I(new_n16489_), .ZN(new_n16490_));
  NOR2_X1    g16193(.A1(new_n16485_), .A2(new_n16488_), .ZN(new_n16491_));
  OAI21_X1   g16194(.A1(new_n16490_), .A2(new_n16491_), .B(new_n16484_), .ZN(new_n16492_));
  OR2_X2     g16195(.A1(new_n16476_), .A2(new_n16483_), .Z(new_n16493_));
  INV_X1     g16196(.I(new_n16491_), .ZN(new_n16494_));
  NAND3_X1   g16197(.A1(new_n16494_), .A2(new_n16493_), .A3(new_n16489_), .ZN(new_n16495_));
  AOI21_X1   g16198(.A1(new_n16492_), .A2(new_n16495_), .B(\a[5] ), .ZN(new_n16496_));
  AOI21_X1   g16199(.A1(new_n16494_), .A2(new_n16489_), .B(new_n16493_), .ZN(new_n16497_));
  NOR3_X1    g16200(.A1(new_n16490_), .A2(new_n16484_), .A3(new_n16491_), .ZN(new_n16498_));
  NOR3_X1    g16201(.A1(new_n16497_), .A2(new_n16498_), .A3(new_n334_), .ZN(new_n16499_));
  OAI21_X1   g16202(.A1(new_n16496_), .A2(new_n16499_), .B(new_n16183_), .ZN(new_n16500_));
  NOR2_X1    g16203(.A1(new_n16496_), .A2(new_n16499_), .ZN(new_n16501_));
  NAND2_X1   g16204(.A1(new_n16501_), .A2(new_n16182_), .ZN(new_n16502_));
  NAND2_X1   g16205(.A1(new_n16502_), .A2(new_n16500_), .ZN(new_n16503_));
  NAND2_X1   g16206(.A1(new_n16181_), .A2(new_n16503_), .ZN(new_n16504_));
  XOR2_X1    g16207(.A1(new_n16501_), .A2(new_n16182_), .Z(new_n16505_));
  NAND2_X1   g16208(.A1(new_n16180_), .A2(new_n16505_), .ZN(new_n16506_));
  NAND2_X1   g16209(.A1(new_n16504_), .A2(new_n16506_), .ZN(\f[68] ));
  INV_X1     g16210(.I(new_n16485_), .ZN(new_n16508_));
  NAND2_X1   g16211(.A1(new_n16493_), .A2(new_n16508_), .ZN(new_n16509_));
  XOR2_X1    g16212(.A1(new_n16488_), .A2(new_n334_), .Z(new_n16510_));
  INV_X1     g16213(.I(new_n16510_), .ZN(new_n16511_));
  OAI21_X1   g16214(.A1(new_n16493_), .A2(new_n16508_), .B(new_n16511_), .ZN(new_n16512_));
  NAND2_X1   g16215(.A1(new_n16482_), .A2(new_n16478_), .ZN(new_n16513_));
  AND2_X2    g16216(.A1(new_n16513_), .A2(new_n16480_), .Z(new_n16514_));
  INV_X1     g16217(.I(new_n16444_), .ZN(new_n16515_));
  OAI21_X1   g16218(.A1(new_n16448_), .A2(new_n16450_), .B(new_n16187_), .ZN(new_n16516_));
  AOI21_X1   g16219(.A1(new_n16515_), .A2(new_n16516_), .B(new_n16456_), .ZN(new_n16517_));
  AOI21_X1   g16220(.A1(new_n16460_), .A2(new_n16463_), .B(new_n16517_), .ZN(new_n16518_));
  NOR2_X1    g16221(.A1(new_n16189_), .A2(new_n16432_), .ZN(new_n16519_));
  NOR2_X1    g16222(.A1(new_n16519_), .A2(new_n16430_), .ZN(new_n16520_));
  NOR2_X1    g16223(.A1(new_n16192_), .A2(new_n16417_), .ZN(new_n16521_));
  NOR2_X1    g16224(.A1(new_n16521_), .A2(new_n16414_), .ZN(new_n16522_));
  INV_X1     g16225(.I(new_n16522_), .ZN(new_n16523_));
  NOR2_X1    g16226(.A1(new_n16405_), .A2(new_n16403_), .ZN(new_n16524_));
  INV_X1     g16227(.I(new_n16381_), .ZN(new_n16525_));
  NOR3_X1    g16228(.A1(new_n16369_), .A2(new_n16375_), .A3(new_n16380_), .ZN(new_n16526_));
  NOR2_X1    g16229(.A1(new_n16387_), .A2(new_n16526_), .ZN(new_n16527_));
  INV_X1     g16230(.I(new_n16363_), .ZN(new_n16528_));
  OAI21_X1   g16231(.A1(new_n16196_), .A2(new_n16367_), .B(new_n16528_), .ZN(new_n16529_));
  INV_X1     g16232(.I(new_n16529_), .ZN(new_n16530_));
  NAND2_X1   g16233(.A1(new_n16198_), .A2(new_n16352_), .ZN(new_n16531_));
  NAND2_X1   g16234(.A1(new_n16531_), .A2(new_n16351_), .ZN(new_n16532_));
  INV_X1     g16235(.I(new_n16532_), .ZN(new_n16533_));
  OAI22_X1   g16236(.A1(new_n4072_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n4067_), .ZN(new_n16534_));
  OAI21_X1   g16237(.A1(new_n4253_), .A2(new_n4318_), .B(new_n16534_), .ZN(new_n16535_));
  AOI21_X1   g16238(.A1(new_n16535_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n16536_));
  XNOR2_X1   g16239(.A1(new_n4778_), .A2(new_n16536_), .ZN(new_n16537_));
  INV_X1     g16240(.I(new_n16537_), .ZN(new_n16538_));
  AOI21_X1   g16241(.A1(new_n16203_), .A2(new_n16326_), .B(new_n16324_), .ZN(new_n16539_));
  INV_X1     g16242(.I(new_n16332_), .ZN(new_n16540_));
  NOR2_X1    g16243(.A1(new_n16327_), .A2(new_n16323_), .ZN(new_n16541_));
  OAI21_X1   g16244(.A1(new_n16541_), .A2(new_n16338_), .B(new_n16201_), .ZN(new_n16542_));
  OAI21_X1   g16245(.A1(new_n16205_), .A2(new_n16305_), .B(new_n16318_), .ZN(new_n16543_));
  INV_X1     g16246(.I(new_n16543_), .ZN(new_n16544_));
  NOR2_X1    g16247(.A1(new_n16286_), .A2(new_n16287_), .ZN(new_n16545_));
  NAND2_X1   g16248(.A1(new_n16286_), .A2(new_n16287_), .ZN(new_n16546_));
  XOR2_X1    g16249(.A1(new_n16290_), .A2(\a[44] ), .Z(new_n16547_));
  AOI21_X1   g16250(.A1(new_n16546_), .A2(new_n16547_), .B(new_n16545_), .ZN(new_n16548_));
  INV_X1     g16251(.I(new_n16548_), .ZN(new_n16549_));
  NAND2_X1   g16252(.A1(new_n16281_), .A2(new_n16283_), .ZN(new_n16550_));
  NAND2_X1   g16253(.A1(new_n16550_), .A2(new_n16279_), .ZN(new_n16551_));
  OAI21_X1   g16254(.A1(new_n16209_), .A2(new_n16272_), .B(new_n16270_), .ZN(new_n16552_));
  OAI21_X1   g16255(.A1(new_n16259_), .A2(new_n16257_), .B(new_n16255_), .ZN(new_n16553_));
  INV_X1     g16256(.I(new_n16553_), .ZN(new_n16554_));
  NOR2_X1    g16257(.A1(new_n16246_), .A2(new_n16214_), .ZN(new_n16555_));
  NOR2_X1    g16258(.A1(new_n16555_), .A2(new_n16245_), .ZN(new_n16556_));
  INV_X1     g16259(.I(new_n16556_), .ZN(new_n16557_));
  NOR2_X1    g16260(.A1(new_n16240_), .A2(new_n16230_), .ZN(new_n16558_));
  NOR2_X1    g16261(.A1(new_n16558_), .A2(new_n16239_), .ZN(new_n16559_));
  AOI22_X1   g16262(.A1(new_n13078_), .A2(\b[10] ), .B1(new_n14320_), .B2(new_n12218_), .ZN(new_n16560_));
  OAI21_X1   g16263(.A1(new_n16560_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n16561_));
  XOR2_X1    g16264(.A1(new_n785_), .A2(new_n16561_), .Z(new_n16562_));
  INV_X1     g16265(.I(new_n16562_), .ZN(new_n16563_));
  INV_X1     g16266(.I(new_n16224_), .ZN(new_n16564_));
  AOI21_X1   g16267(.A1(new_n16218_), .A2(new_n16564_), .B(new_n16225_), .ZN(new_n16565_));
  INV_X1     g16268(.I(new_n16565_), .ZN(new_n16566_));
  OAI22_X1   g16269(.A1(new_n13880_), .A2(new_n649_), .B1(new_n472_), .B2(new_n13885_), .ZN(new_n16567_));
  AOI21_X1   g16270(.A1(new_n16567_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n16568_));
  XOR2_X1    g16271(.A1(new_n569_), .A2(new_n16568_), .Z(new_n16569_));
  NOR2_X1    g16272(.A1(new_n13476_), .A2(new_n419_), .ZN(new_n16570_));
  XOR2_X1    g16273(.A1(new_n14736_), .A2(new_n419_), .Z(new_n16571_));
  NAND2_X1   g16274(.A1(new_n16571_), .A2(\b[6] ), .ZN(new_n16572_));
  XOR2_X1    g16275(.A1(new_n16572_), .A2(new_n16570_), .Z(new_n16573_));
  NOR2_X1    g16276(.A1(new_n16573_), .A2(new_n364_), .ZN(new_n16574_));
  NOR2_X1    g16277(.A1(new_n260_), .A2(new_n334_), .ZN(new_n16575_));
  NOR2_X1    g16278(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n16576_));
  NOR2_X1    g16279(.A1(new_n16575_), .A2(new_n16576_), .ZN(new_n16577_));
  INV_X1     g16280(.I(new_n16577_), .ZN(new_n16578_));
  AOI21_X1   g16281(.A1(new_n16573_), .A2(new_n16578_), .B(new_n16574_), .ZN(new_n16579_));
  XOR2_X1    g16282(.A1(new_n16569_), .A2(new_n16579_), .Z(new_n16580_));
  NAND2_X1   g16283(.A1(new_n16580_), .A2(new_n16566_), .ZN(new_n16581_));
  XOR2_X1    g16284(.A1(new_n759_), .A2(new_n16568_), .Z(new_n16582_));
  INV_X1     g16285(.I(new_n16579_), .ZN(new_n16583_));
  NAND2_X1   g16286(.A1(new_n16582_), .A2(new_n16583_), .ZN(new_n16584_));
  NAND2_X1   g16287(.A1(new_n16569_), .A2(new_n16579_), .ZN(new_n16585_));
  NAND2_X1   g16288(.A1(new_n16584_), .A2(new_n16585_), .ZN(new_n16586_));
  NAND2_X1   g16289(.A1(new_n16586_), .A2(new_n16565_), .ZN(new_n16587_));
  NAND2_X1   g16290(.A1(new_n16581_), .A2(new_n16587_), .ZN(new_n16588_));
  NAND2_X1   g16291(.A1(new_n16563_), .A2(new_n16588_), .ZN(new_n16589_));
  NAND3_X1   g16292(.A1(new_n16562_), .A2(new_n16581_), .A3(new_n16587_), .ZN(new_n16590_));
  AOI21_X1   g16293(.A1(new_n16590_), .A2(new_n16589_), .B(new_n16559_), .ZN(new_n16591_));
  INV_X1     g16294(.I(new_n16559_), .ZN(new_n16592_));
  XOR2_X1    g16295(.A1(new_n16588_), .A2(new_n16562_), .Z(new_n16593_));
  NOR2_X1    g16296(.A1(new_n16593_), .A2(new_n16592_), .ZN(new_n16594_));
  NOR2_X1    g16297(.A1(new_n16594_), .A2(new_n16591_), .ZN(new_n16595_));
  AOI22_X1   g16298(.A1(new_n10969_), .A2(new_n1105_), .B1(new_n11394_), .B2(\b[13] ), .ZN(new_n16596_));
  OAI21_X1   g16299(.A1(new_n16596_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n16597_));
  XNOR2_X1   g16300(.A1(new_n1024_), .A2(new_n16597_), .ZN(new_n16598_));
  XOR2_X1    g16301(.A1(new_n16595_), .A2(new_n16598_), .Z(new_n16599_));
  NAND2_X1   g16302(.A1(new_n16599_), .A2(new_n16557_), .ZN(new_n16600_));
  NOR2_X1    g16303(.A1(new_n16595_), .A2(new_n16598_), .ZN(new_n16601_));
  INV_X1     g16304(.I(new_n16595_), .ZN(new_n16602_));
  INV_X1     g16305(.I(new_n16598_), .ZN(new_n16603_));
  NOR2_X1    g16306(.A1(new_n16602_), .A2(new_n16603_), .ZN(new_n16604_));
  OAI21_X1   g16307(.A1(new_n16604_), .A2(new_n16601_), .B(new_n16556_), .ZN(new_n16605_));
  NAND2_X1   g16308(.A1(new_n16600_), .A2(new_n16605_), .ZN(new_n16606_));
  AOI22_X1   g16309(.A1(new_n11415_), .A2(new_n1296_), .B1(\b[16] ), .B2(new_n10145_), .ZN(new_n16607_));
  OAI21_X1   g16310(.A1(new_n16607_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n16608_));
  XOR2_X1    g16311(.A1(new_n1299_), .A2(new_n16608_), .Z(new_n16609_));
  XOR2_X1    g16312(.A1(new_n16606_), .A2(new_n16609_), .Z(new_n16610_));
  NOR2_X1    g16313(.A1(new_n16610_), .A2(new_n16554_), .ZN(new_n16611_));
  NAND3_X1   g16314(.A1(new_n16600_), .A2(new_n16605_), .A3(new_n16609_), .ZN(new_n16612_));
  INV_X1     g16315(.I(new_n16609_), .ZN(new_n16613_));
  NAND2_X1   g16316(.A1(new_n16606_), .A2(new_n16613_), .ZN(new_n16614_));
  AOI21_X1   g16317(.A1(new_n16614_), .A2(new_n16612_), .B(new_n16553_), .ZN(new_n16615_));
  OAI22_X1   g16318(.A1(new_n8644_), .A2(new_n1525_), .B1(new_n1634_), .B2(new_n9388_), .ZN(new_n16616_));
  OAI21_X1   g16319(.A1(new_n1518_), .A2(new_n10154_), .B(new_n16616_), .ZN(new_n16617_));
  AOI21_X1   g16320(.A1(new_n16617_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n16618_));
  XNOR2_X1   g16321(.A1(new_n1638_), .A2(new_n16618_), .ZN(new_n16619_));
  NOR3_X1    g16322(.A1(new_n16611_), .A2(new_n16615_), .A3(new_n16619_), .ZN(new_n16620_));
  NOR2_X1    g16323(.A1(new_n16611_), .A2(new_n16615_), .ZN(new_n16621_));
  INV_X1     g16324(.I(new_n16619_), .ZN(new_n16622_));
  NOR2_X1    g16325(.A1(new_n16621_), .A2(new_n16622_), .ZN(new_n16623_));
  OAI21_X1   g16326(.A1(new_n16623_), .A2(new_n16620_), .B(new_n16552_), .ZN(new_n16624_));
  INV_X1     g16327(.I(new_n16552_), .ZN(new_n16625_));
  XOR2_X1    g16328(.A1(new_n16621_), .A2(new_n16622_), .Z(new_n16626_));
  NAND2_X1   g16329(.A1(new_n16626_), .A2(new_n16625_), .ZN(new_n16627_));
  NAND2_X1   g16330(.A1(new_n16627_), .A2(new_n16624_), .ZN(new_n16628_));
  OAI22_X1   g16331(.A1(new_n7619_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n8309_), .ZN(new_n16629_));
  OAI21_X1   g16332(.A1(new_n1803_), .A2(new_n7947_), .B(new_n16629_), .ZN(new_n16630_));
  AOI21_X1   g16333(.A1(new_n16630_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n16631_));
  XOR2_X1    g16334(.A1(new_n2106_), .A2(new_n16631_), .Z(new_n16632_));
  INV_X1     g16335(.I(new_n16632_), .ZN(new_n16633_));
  XOR2_X1    g16336(.A1(new_n16628_), .A2(new_n16633_), .Z(new_n16634_));
  NAND2_X1   g16337(.A1(new_n16634_), .A2(new_n16551_), .ZN(new_n16635_));
  INV_X1     g16338(.I(new_n16551_), .ZN(new_n16636_));
  NAND2_X1   g16339(.A1(new_n16628_), .A2(new_n16633_), .ZN(new_n16637_));
  INV_X1     g16340(.I(new_n16637_), .ZN(new_n16638_));
  NOR2_X1    g16341(.A1(new_n16628_), .A2(new_n16633_), .ZN(new_n16639_));
  OAI21_X1   g16342(.A1(new_n16638_), .A2(new_n16639_), .B(new_n16636_), .ZN(new_n16640_));
  NAND2_X1   g16343(.A1(new_n16635_), .A2(new_n16640_), .ZN(new_n16641_));
  OAI22_X1   g16344(.A1(new_n6644_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n6647_), .ZN(new_n16642_));
  OAI21_X1   g16345(.A1(new_n2281_), .A2(new_n7284_), .B(new_n16642_), .ZN(new_n16643_));
  AOI21_X1   g16346(.A1(new_n16643_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n16644_));
  XNOR2_X1   g16347(.A1(new_n2647_), .A2(new_n16644_), .ZN(new_n16645_));
  XOR2_X1    g16348(.A1(new_n16641_), .A2(new_n16645_), .Z(new_n16646_));
  NAND2_X1   g16349(.A1(new_n16646_), .A2(new_n16549_), .ZN(new_n16647_));
  NOR2_X1    g16350(.A1(new_n16641_), .A2(new_n16645_), .ZN(new_n16648_));
  AND2_X2    g16351(.A1(new_n16641_), .A2(new_n16645_), .Z(new_n16649_));
  OAI21_X1   g16352(.A1(new_n16649_), .A2(new_n16648_), .B(new_n16548_), .ZN(new_n16650_));
  OAI22_X1   g16353(.A1(new_n5993_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n5991_), .ZN(new_n16651_));
  OAI21_X1   g16354(.A1(new_n2842_), .A2(new_n5997_), .B(new_n16651_), .ZN(new_n16652_));
  AOI21_X1   g16355(.A1(new_n16652_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n16653_));
  XNOR2_X1   g16356(.A1(new_n3264_), .A2(new_n16653_), .ZN(new_n16654_));
  INV_X1     g16357(.I(new_n16654_), .ZN(new_n16655_));
  NAND3_X1   g16358(.A1(new_n16647_), .A2(new_n16650_), .A3(new_n16655_), .ZN(new_n16656_));
  NAND2_X1   g16359(.A1(new_n16647_), .A2(new_n16650_), .ZN(new_n16657_));
  NAND2_X1   g16360(.A1(new_n16657_), .A2(new_n16654_), .ZN(new_n16658_));
  AOI21_X1   g16361(.A1(new_n16656_), .A2(new_n16658_), .B(new_n16544_), .ZN(new_n16659_));
  XOR2_X1    g16362(.A1(new_n16657_), .A2(new_n16655_), .Z(new_n16660_));
  NOR2_X1    g16363(.A1(new_n16660_), .A2(new_n16543_), .ZN(new_n16661_));
  NOR2_X1    g16364(.A1(new_n16661_), .A2(new_n16659_), .ZN(new_n16662_));
  OAI22_X1   g16365(.A1(new_n5420_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n5107_), .ZN(new_n16663_));
  OAI21_X1   g16366(.A1(new_n3709_), .A2(new_n5112_), .B(new_n16663_), .ZN(new_n16664_));
  AOI21_X1   g16367(.A1(new_n16664_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n16665_));
  XNOR2_X1   g16368(.A1(new_n3993_), .A2(new_n16665_), .ZN(new_n16666_));
  NOR2_X1    g16369(.A1(new_n16662_), .A2(new_n16666_), .ZN(new_n16667_));
  INV_X1     g16370(.I(new_n16667_), .ZN(new_n16668_));
  NAND2_X1   g16371(.A1(new_n16662_), .A2(new_n16666_), .ZN(new_n16669_));
  NAND2_X1   g16372(.A1(new_n16668_), .A2(new_n16669_), .ZN(new_n16670_));
  NAND3_X1   g16373(.A1(new_n16670_), .A2(new_n16540_), .A3(new_n16542_), .ZN(new_n16671_));
  NAND2_X1   g16374(.A1(new_n16542_), .A2(new_n16540_), .ZN(new_n16672_));
  INV_X1     g16375(.I(new_n16669_), .ZN(new_n16673_));
  NOR2_X1    g16376(.A1(new_n16673_), .A2(new_n16667_), .ZN(new_n16674_));
  NAND2_X1   g16377(.A1(new_n16672_), .A2(new_n16674_), .ZN(new_n16675_));
  NAND2_X1   g16378(.A1(new_n16675_), .A2(new_n16671_), .ZN(new_n16676_));
  NAND2_X1   g16379(.A1(new_n16676_), .A2(new_n16539_), .ZN(new_n16677_));
  INV_X1     g16380(.I(new_n16539_), .ZN(new_n16678_));
  NAND3_X1   g16381(.A1(new_n16675_), .A2(new_n16671_), .A3(new_n16678_), .ZN(new_n16679_));
  AOI21_X1   g16382(.A1(new_n16677_), .A2(new_n16679_), .B(new_n16538_), .ZN(new_n16680_));
  AOI21_X1   g16383(.A1(new_n16675_), .A2(new_n16671_), .B(new_n16678_), .ZN(new_n16681_));
  INV_X1     g16384(.I(new_n16679_), .ZN(new_n16682_));
  NOR3_X1    g16385(.A1(new_n16682_), .A2(new_n16681_), .A3(new_n16537_), .ZN(new_n16683_));
  OAI22_X1   g16386(.A1(new_n5353_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n5913_), .ZN(new_n16684_));
  OAI21_X1   g16387(.A1(new_n5068_), .A2(new_n3569_), .B(new_n16684_), .ZN(new_n16685_));
  AOI21_X1   g16388(.A1(new_n16685_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n16686_));
  XNOR2_X1   g16389(.A1(new_n5600_), .A2(new_n16686_), .ZN(new_n16687_));
  INV_X1     g16390(.I(new_n16687_), .ZN(new_n16688_));
  OAI21_X1   g16391(.A1(new_n16683_), .A2(new_n16680_), .B(new_n16688_), .ZN(new_n16689_));
  OAI21_X1   g16392(.A1(new_n16682_), .A2(new_n16681_), .B(new_n16537_), .ZN(new_n16690_));
  NAND3_X1   g16393(.A1(new_n16677_), .A2(new_n16679_), .A3(new_n16538_), .ZN(new_n16691_));
  NAND3_X1   g16394(.A1(new_n16690_), .A2(new_n16691_), .A3(new_n16687_), .ZN(new_n16692_));
  AOI21_X1   g16395(.A1(new_n16689_), .A2(new_n16692_), .B(new_n16533_), .ZN(new_n16693_));
  NAND3_X1   g16396(.A1(new_n16690_), .A2(new_n16691_), .A3(new_n16688_), .ZN(new_n16694_));
  OAI21_X1   g16397(.A1(new_n16683_), .A2(new_n16680_), .B(new_n16687_), .ZN(new_n16695_));
  AOI21_X1   g16398(.A1(new_n16695_), .A2(new_n16694_), .B(new_n16532_), .ZN(new_n16696_));
  OAI22_X1   g16399(.A1(new_n6229_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n6538_), .ZN(new_n16697_));
  OAI21_X1   g16400(.A1(new_n5921_), .A2(new_n2884_), .B(new_n16697_), .ZN(new_n16698_));
  AOI21_X1   g16401(.A1(new_n16698_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n16699_));
  XOR2_X1    g16402(.A1(new_n6543_), .A2(new_n16699_), .Z(new_n16700_));
  INV_X1     g16403(.I(new_n16700_), .ZN(new_n16701_));
  OAI21_X1   g16404(.A1(new_n16693_), .A2(new_n16696_), .B(new_n16701_), .ZN(new_n16702_));
  NOR3_X1    g16405(.A1(new_n16693_), .A2(new_n16696_), .A3(new_n16701_), .ZN(new_n16703_));
  INV_X1     g16406(.I(new_n16703_), .ZN(new_n16704_));
  AOI21_X1   g16407(.A1(new_n16704_), .A2(new_n16702_), .B(new_n16530_), .ZN(new_n16705_));
  AOI21_X1   g16408(.A1(new_n16690_), .A2(new_n16691_), .B(new_n16687_), .ZN(new_n16706_));
  NOR3_X1    g16409(.A1(new_n16683_), .A2(new_n16680_), .A3(new_n16688_), .ZN(new_n16707_));
  OAI21_X1   g16410(.A1(new_n16707_), .A2(new_n16706_), .B(new_n16532_), .ZN(new_n16708_));
  NOR3_X1    g16411(.A1(new_n16683_), .A2(new_n16680_), .A3(new_n16687_), .ZN(new_n16709_));
  AOI21_X1   g16412(.A1(new_n16690_), .A2(new_n16691_), .B(new_n16688_), .ZN(new_n16710_));
  OAI21_X1   g16413(.A1(new_n16709_), .A2(new_n16710_), .B(new_n16533_), .ZN(new_n16711_));
  NAND3_X1   g16414(.A1(new_n16711_), .A2(new_n16708_), .A3(new_n16701_), .ZN(new_n16712_));
  OAI21_X1   g16415(.A1(new_n16693_), .A2(new_n16696_), .B(new_n16700_), .ZN(new_n16713_));
  AOI21_X1   g16416(.A1(new_n16712_), .A2(new_n16713_), .B(new_n16529_), .ZN(new_n16714_));
  OAI22_X1   g16417(.A1(new_n2171_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n2166_), .ZN(new_n16715_));
  OAI21_X1   g16418(.A1(new_n6847_), .A2(new_n2322_), .B(new_n16715_), .ZN(new_n16716_));
  AOI21_X1   g16419(.A1(new_n16716_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n16717_));
  XOR2_X1    g16420(.A1(new_n7516_), .A2(new_n16717_), .Z(new_n16718_));
  NOR3_X1    g16421(.A1(new_n16705_), .A2(new_n16714_), .A3(new_n16718_), .ZN(new_n16719_));
  INV_X1     g16422(.I(new_n16702_), .ZN(new_n16720_));
  OAI21_X1   g16423(.A1(new_n16720_), .A2(new_n16703_), .B(new_n16529_), .ZN(new_n16721_));
  INV_X1     g16424(.I(new_n16714_), .ZN(new_n16722_));
  INV_X1     g16425(.I(new_n16718_), .ZN(new_n16723_));
  AOI21_X1   g16426(.A1(new_n16722_), .A2(new_n16721_), .B(new_n16723_), .ZN(new_n16724_));
  OAI22_X1   g16427(.A1(new_n16724_), .A2(new_n16719_), .B1(new_n16527_), .B2(new_n16525_), .ZN(new_n16725_));
  NOR2_X1    g16428(.A1(new_n16527_), .A2(new_n16525_), .ZN(new_n16726_));
  AOI21_X1   g16429(.A1(new_n16722_), .A2(new_n16721_), .B(new_n16718_), .ZN(new_n16727_));
  NOR3_X1    g16430(.A1(new_n16705_), .A2(new_n16714_), .A3(new_n16723_), .ZN(new_n16728_));
  OAI21_X1   g16431(.A1(new_n16727_), .A2(new_n16728_), .B(new_n16726_), .ZN(new_n16729_));
  OAI22_X1   g16432(.A1(new_n1712_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n1707_), .ZN(new_n16730_));
  OAI21_X1   g16433(.A1(new_n7870_), .A2(new_n1850_), .B(new_n16730_), .ZN(new_n16731_));
  AOI21_X1   g16434(.A1(new_n16731_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n16732_));
  XOR2_X1    g16435(.A1(new_n8568_), .A2(new_n16732_), .Z(new_n16733_));
  AOI21_X1   g16436(.A1(new_n16729_), .A2(new_n16725_), .B(new_n16733_), .ZN(new_n16734_));
  NAND2_X1   g16437(.A1(new_n16729_), .A2(new_n16725_), .ZN(new_n16735_));
  INV_X1     g16438(.I(new_n16733_), .ZN(new_n16736_));
  NOR2_X1    g16439(.A1(new_n16735_), .A2(new_n16736_), .ZN(new_n16737_));
  OAI22_X1   g16440(.A1(new_n16737_), .A2(new_n16734_), .B1(new_n16524_), .B2(new_n16396_), .ZN(new_n16738_));
  INV_X1     g16441(.I(new_n16738_), .ZN(new_n16739_));
  NOR2_X1    g16442(.A1(new_n16524_), .A2(new_n16396_), .ZN(new_n16740_));
  NOR2_X1    g16443(.A1(new_n16735_), .A2(new_n16733_), .ZN(new_n16741_));
  AOI21_X1   g16444(.A1(new_n16729_), .A2(new_n16725_), .B(new_n16736_), .ZN(new_n16742_));
  OAI21_X1   g16445(.A1(new_n16741_), .A2(new_n16742_), .B(new_n16740_), .ZN(new_n16743_));
  INV_X1     g16446(.I(new_n16743_), .ZN(new_n16744_));
  OAI22_X1   g16447(.A1(new_n1347_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n1344_), .ZN(new_n16745_));
  OAI21_X1   g16448(.A1(new_n8948_), .A2(new_n1457_), .B(new_n16745_), .ZN(new_n16746_));
  AOI21_X1   g16449(.A1(new_n16746_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n16747_));
  XNOR2_X1   g16450(.A1(new_n9642_), .A2(new_n16747_), .ZN(new_n16748_));
  INV_X1     g16451(.I(new_n16748_), .ZN(new_n16749_));
  OAI21_X1   g16452(.A1(new_n16739_), .A2(new_n16744_), .B(new_n16749_), .ZN(new_n16750_));
  NAND3_X1   g16453(.A1(new_n16738_), .A2(new_n16743_), .A3(new_n16748_), .ZN(new_n16751_));
  NAND2_X1   g16454(.A1(new_n16750_), .A2(new_n16751_), .ZN(new_n16752_));
  NAND2_X1   g16455(.A1(new_n16752_), .A2(new_n16523_), .ZN(new_n16753_));
  NOR3_X1    g16456(.A1(new_n16739_), .A2(new_n16744_), .A3(new_n16748_), .ZN(new_n16754_));
  AOI21_X1   g16457(.A1(new_n16738_), .A2(new_n16743_), .B(new_n16749_), .ZN(new_n16755_));
  OAI21_X1   g16458(.A1(new_n16754_), .A2(new_n16755_), .B(new_n16522_), .ZN(new_n16756_));
  OAI22_X1   g16459(.A1(new_n1055_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n1061_), .ZN(new_n16757_));
  OAI21_X1   g16460(.A1(new_n10031_), .A2(new_n1332_), .B(new_n16757_), .ZN(new_n16758_));
  AOI21_X1   g16461(.A1(new_n16758_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n16759_));
  XNOR2_X1   g16462(.A1(new_n10866_), .A2(new_n16759_), .ZN(new_n16760_));
  AOI21_X1   g16463(.A1(new_n16753_), .A2(new_n16756_), .B(new_n16760_), .ZN(new_n16761_));
  NAND2_X1   g16464(.A1(new_n16753_), .A2(new_n16756_), .ZN(new_n16762_));
  INV_X1     g16465(.I(new_n16760_), .ZN(new_n16763_));
  NOR2_X1    g16466(.A1(new_n16762_), .A2(new_n16763_), .ZN(new_n16764_));
  NOR2_X1    g16467(.A1(new_n16764_), .A2(new_n16761_), .ZN(new_n16765_));
  NOR2_X1    g16468(.A1(new_n16765_), .A2(new_n16520_), .ZN(new_n16766_));
  XOR2_X1    g16469(.A1(new_n16762_), .A2(new_n16763_), .Z(new_n16767_));
  AOI21_X1   g16470(.A1(new_n16520_), .A2(new_n16767_), .B(new_n16766_), .ZN(new_n16768_));
  OAI21_X1   g16471(.A1(new_n16186_), .A2(new_n16103_), .B(new_n16443_), .ZN(new_n16769_));
  OAI22_X1   g16472(.A1(new_n970_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n820_), .ZN(new_n16770_));
  OAI21_X1   g16473(.A1(new_n11738_), .A2(new_n894_), .B(new_n16770_), .ZN(new_n16771_));
  AOI21_X1   g16474(.A1(new_n16771_), .A2(new_n827_), .B(new_n970_), .ZN(new_n16772_));
  XNOR2_X1   g16475(.A1(new_n12128_), .A2(new_n16772_), .ZN(new_n16773_));
  AOI21_X1   g16476(.A1(new_n16769_), .A2(new_n16442_), .B(new_n16773_), .ZN(new_n16774_));
  INV_X1     g16477(.I(new_n16774_), .ZN(new_n16775_));
  NAND3_X1   g16478(.A1(new_n16769_), .A2(new_n16442_), .A3(new_n16773_), .ZN(new_n16776_));
  AOI21_X1   g16479(.A1(new_n16775_), .A2(new_n16776_), .B(new_n16768_), .ZN(new_n16777_));
  NAND2_X1   g16480(.A1(new_n16767_), .A2(new_n16520_), .ZN(new_n16778_));
  OAI21_X1   g16481(.A1(new_n16520_), .A2(new_n16765_), .B(new_n16778_), .ZN(new_n16779_));
  INV_X1     g16482(.I(new_n16773_), .ZN(new_n16780_));
  NAND3_X1   g16483(.A1(new_n16769_), .A2(new_n16442_), .A3(new_n16780_), .ZN(new_n16781_));
  AOI21_X1   g16484(.A1(new_n16769_), .A2(new_n16442_), .B(new_n16780_), .ZN(new_n16782_));
  INV_X1     g16485(.I(new_n16782_), .ZN(new_n16783_));
  AOI21_X1   g16486(.A1(new_n16783_), .A2(new_n16781_), .B(new_n16779_), .ZN(new_n16784_));
  OAI22_X1   g16487(.A1(new_n607_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n610_), .ZN(new_n16785_));
  OAI21_X1   g16488(.A1(new_n12542_), .A2(new_n684_), .B(new_n16785_), .ZN(new_n16786_));
  AOI21_X1   g16489(.A1(new_n16786_), .A2(new_n612_), .B(new_n607_), .ZN(new_n16787_));
  XNOR2_X1   g16490(.A1(new_n13371_), .A2(new_n16787_), .ZN(new_n16788_));
  INV_X1     g16491(.I(new_n16788_), .ZN(new_n16789_));
  OAI21_X1   g16492(.A1(new_n16784_), .A2(new_n16777_), .B(new_n16789_), .ZN(new_n16790_));
  INV_X1     g16493(.I(new_n16776_), .ZN(new_n16791_));
  OAI21_X1   g16494(.A1(new_n16791_), .A2(new_n16774_), .B(new_n16779_), .ZN(new_n16792_));
  INV_X1     g16495(.I(new_n16781_), .ZN(new_n16793_));
  OAI21_X1   g16496(.A1(new_n16793_), .A2(new_n16782_), .B(new_n16768_), .ZN(new_n16794_));
  NAND3_X1   g16497(.A1(new_n16792_), .A2(new_n16794_), .A3(new_n16788_), .ZN(new_n16795_));
  AOI21_X1   g16498(.A1(new_n16790_), .A2(new_n16795_), .B(new_n16518_), .ZN(new_n16796_));
  OAI21_X1   g16499(.A1(new_n16185_), .A2(new_n16459_), .B(new_n16458_), .ZN(new_n16797_));
  NAND3_X1   g16500(.A1(new_n16792_), .A2(new_n16794_), .A3(new_n16789_), .ZN(new_n16798_));
  OAI21_X1   g16501(.A1(new_n16784_), .A2(new_n16777_), .B(new_n16788_), .ZN(new_n16799_));
  AOI21_X1   g16502(.A1(new_n16799_), .A2(new_n16798_), .B(new_n16797_), .ZN(new_n16800_));
  OAI22_X1   g16503(.A1(new_n448_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n450_), .ZN(new_n16801_));
  OAI21_X1   g16504(.A1(new_n13785_), .A2(new_n496_), .B(new_n16801_), .ZN(new_n16802_));
  AOI21_X1   g16505(.A1(new_n16802_), .A2(new_n452_), .B(new_n448_), .ZN(new_n16803_));
  XNOR2_X1   g16506(.A1(new_n14599_), .A2(new_n16803_), .ZN(new_n16804_));
  INV_X1     g16507(.I(new_n16804_), .ZN(new_n16805_));
  OAI21_X1   g16508(.A1(new_n16796_), .A2(new_n16800_), .B(new_n16805_), .ZN(new_n16806_));
  AOI21_X1   g16509(.A1(new_n16792_), .A2(new_n16794_), .B(new_n16788_), .ZN(new_n16807_));
  NOR3_X1    g16510(.A1(new_n16784_), .A2(new_n16777_), .A3(new_n16789_), .ZN(new_n16808_));
  OAI21_X1   g16511(.A1(new_n16808_), .A2(new_n16807_), .B(new_n16797_), .ZN(new_n16809_));
  NOR3_X1    g16512(.A1(new_n16784_), .A2(new_n16777_), .A3(new_n16788_), .ZN(new_n16810_));
  AOI21_X1   g16513(.A1(new_n16792_), .A2(new_n16794_), .B(new_n16789_), .ZN(new_n16811_));
  OAI21_X1   g16514(.A1(new_n16811_), .A2(new_n16810_), .B(new_n16518_), .ZN(new_n16812_));
  NAND3_X1   g16515(.A1(new_n16812_), .A2(new_n16809_), .A3(new_n16804_), .ZN(new_n16813_));
  AND2_X2    g16516(.A1(new_n16806_), .A2(new_n16813_), .Z(new_n16814_));
  NAND3_X1   g16517(.A1(new_n16812_), .A2(new_n16809_), .A3(new_n16805_), .ZN(new_n16815_));
  OAI21_X1   g16518(.A1(new_n16796_), .A2(new_n16800_), .B(new_n16804_), .ZN(new_n16816_));
  NAND2_X1   g16519(.A1(new_n16816_), .A2(new_n16815_), .ZN(new_n16817_));
  NAND3_X1   g16520(.A1(new_n16817_), .A2(new_n16480_), .A3(new_n16513_), .ZN(new_n16818_));
  OAI21_X1   g16521(.A1(new_n16514_), .A2(new_n16814_), .B(new_n16818_), .ZN(new_n16819_));
  NAND3_X1   g16522(.A1(new_n16512_), .A2(new_n16819_), .A3(new_n16509_), .ZN(new_n16820_));
  NOR2_X1    g16523(.A1(new_n16484_), .A2(new_n16485_), .ZN(new_n16821_));
  AOI21_X1   g16524(.A1(new_n16484_), .A2(new_n16485_), .B(new_n16510_), .ZN(new_n16822_));
  AOI22_X1   g16525(.A1(new_n16513_), .A2(new_n16480_), .B1(new_n16806_), .B2(new_n16813_), .ZN(new_n16823_));
  AOI21_X1   g16526(.A1(new_n16514_), .A2(new_n16817_), .B(new_n16823_), .ZN(new_n16824_));
  OAI21_X1   g16527(.A1(new_n16821_), .A2(new_n16822_), .B(new_n16824_), .ZN(new_n16825_));
  NAND2_X1   g16528(.A1(new_n16820_), .A2(new_n16825_), .ZN(new_n16826_));
  NAND2_X1   g16529(.A1(new_n16505_), .A2(new_n16826_), .ZN(new_n16827_));
  XOR2_X1    g16530(.A1(new_n16827_), .A2(new_n16500_), .Z(new_n16828_));
  XOR2_X1    g16531(.A1(new_n16828_), .A2(new_n16181_), .Z(\f[69] ));
  AOI21_X1   g16532(.A1(new_n16797_), .A2(new_n16795_), .B(new_n16807_), .ZN(new_n16830_));
  INV_X1     g16533(.I(new_n16830_), .ZN(new_n16831_));
  AOI21_X1   g16534(.A1(new_n16779_), .A2(new_n16776_), .B(new_n16774_), .ZN(new_n16832_));
  INV_X1     g16535(.I(new_n16832_), .ZN(new_n16833_));
  NOR2_X1    g16536(.A1(new_n16764_), .A2(new_n16520_), .ZN(new_n16834_));
  NOR2_X1    g16537(.A1(new_n16834_), .A2(new_n16761_), .ZN(new_n16835_));
  INV_X1     g16538(.I(new_n16835_), .ZN(new_n16836_));
  NAND2_X1   g16539(.A1(new_n16523_), .A2(new_n16751_), .ZN(new_n16837_));
  NAND2_X1   g16540(.A1(new_n16837_), .A2(new_n16750_), .ZN(new_n16838_));
  INV_X1     g16541(.I(new_n16838_), .ZN(new_n16839_));
  NOR2_X1    g16542(.A1(new_n16737_), .A2(new_n16740_), .ZN(new_n16840_));
  NOR2_X1    g16543(.A1(new_n16840_), .A2(new_n16734_), .ZN(new_n16841_));
  INV_X1     g16544(.I(new_n16841_), .ZN(new_n16842_));
  NOR2_X1    g16545(.A1(new_n16726_), .A2(new_n16724_), .ZN(new_n16843_));
  NOR2_X1    g16546(.A1(new_n16843_), .A2(new_n16719_), .ZN(new_n16844_));
  INV_X1     g16547(.I(new_n16844_), .ZN(new_n16845_));
  AND2_X2    g16548(.A1(new_n16713_), .A2(new_n16529_), .Z(new_n16846_));
  INV_X1     g16549(.I(new_n16846_), .ZN(new_n16847_));
  NAND2_X1   g16550(.A1(new_n16847_), .A2(new_n16712_), .ZN(new_n16848_));
  INV_X1     g16551(.I(new_n16848_), .ZN(new_n16849_));
  AOI21_X1   g16552(.A1(new_n16532_), .A2(new_n16695_), .B(new_n16709_), .ZN(new_n16850_));
  AOI21_X1   g16553(.A1(new_n16542_), .A2(new_n16540_), .B(new_n16537_), .ZN(new_n16851_));
  NOR2_X1    g16554(.A1(new_n16672_), .A2(new_n16538_), .ZN(new_n16852_));
  XOR2_X1    g16555(.A1(new_n16670_), .A2(new_n16539_), .Z(new_n16853_));
  NOR2_X1    g16556(.A1(new_n16853_), .A2(new_n16852_), .ZN(new_n16854_));
  NOR2_X1    g16557(.A1(new_n16854_), .A2(new_n16851_), .ZN(new_n16855_));
  AOI21_X1   g16558(.A1(new_n16678_), .A2(new_n16669_), .B(new_n16667_), .ZN(new_n16856_));
  NOR2_X1    g16559(.A1(new_n16649_), .A2(new_n16548_), .ZN(new_n16857_));
  NOR2_X1    g16560(.A1(new_n16857_), .A2(new_n16648_), .ZN(new_n16858_));
  NOR2_X1    g16561(.A1(new_n16623_), .A2(new_n16625_), .ZN(new_n16859_));
  NOR2_X1    g16562(.A1(new_n16859_), .A2(new_n16620_), .ZN(new_n16860_));
  NAND2_X1   g16563(.A1(new_n16614_), .A2(new_n16553_), .ZN(new_n16861_));
  AND2_X2    g16564(.A1(new_n16861_), .A2(new_n16612_), .Z(new_n16862_));
  INV_X1     g16565(.I(new_n16862_), .ZN(new_n16863_));
  AOI22_X1   g16566(.A1(new_n8631_), .A2(\b[21] ), .B1(\b[22] ), .B2(new_n9382_), .ZN(new_n16864_));
  AOI21_X1   g16567(.A1(\b[20] ), .A2(new_n9731_), .B(new_n16864_), .ZN(new_n16865_));
  OAI21_X1   g16568(.A1(new_n16865_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n16866_));
  XNOR2_X1   g16569(.A1(new_n1808_), .A2(new_n16866_), .ZN(new_n16867_));
  AOI22_X1   g16570(.A1(new_n10969_), .A2(new_n1111_), .B1(new_n11394_), .B2(\b[14] ), .ZN(new_n16868_));
  OAI21_X1   g16571(.A1(new_n16868_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n16869_));
  XNOR2_X1   g16572(.A1(new_n1114_), .A2(new_n16869_), .ZN(new_n16870_));
  INV_X1     g16573(.I(new_n16585_), .ZN(new_n16871_));
  AOI21_X1   g16574(.A1(new_n16566_), .A2(new_n16584_), .B(new_n16871_), .ZN(new_n16872_));
  INV_X1     g16575(.I(new_n16872_), .ZN(new_n16873_));
  OAI22_X1   g16576(.A1(new_n13880_), .A2(new_n657_), .B1(new_n515_), .B2(new_n13885_), .ZN(new_n16874_));
  AOI21_X1   g16577(.A1(new_n16874_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n16875_));
  XOR2_X1    g16578(.A1(new_n660_), .A2(new_n16875_), .Z(new_n16876_));
  INV_X1     g16579(.I(new_n16876_), .ZN(new_n16877_));
  NOR2_X1    g16580(.A1(new_n16573_), .A2(new_n16576_), .ZN(new_n16878_));
  NOR2_X1    g16581(.A1(new_n16878_), .A2(new_n16575_), .ZN(new_n16879_));
  NOR2_X1    g16582(.A1(new_n13476_), .A2(new_n420_), .ZN(new_n16880_));
  XOR2_X1    g16583(.A1(new_n14736_), .A2(new_n420_), .Z(new_n16881_));
  NAND2_X1   g16584(.A1(new_n16881_), .A2(\b[7] ), .ZN(new_n16882_));
  XOR2_X1    g16585(.A1(new_n16882_), .A2(new_n16880_), .Z(new_n16883_));
  XOR2_X1    g16586(.A1(new_n16879_), .A2(new_n16883_), .Z(new_n16884_));
  NOR2_X1    g16587(.A1(new_n16877_), .A2(new_n16884_), .ZN(new_n16885_));
  INV_X1     g16588(.I(new_n16879_), .ZN(new_n16886_));
  NOR2_X1    g16589(.A1(new_n16886_), .A2(new_n16883_), .ZN(new_n16887_));
  INV_X1     g16590(.I(new_n16883_), .ZN(new_n16888_));
  NOR2_X1    g16591(.A1(new_n16879_), .A2(new_n16888_), .ZN(new_n16889_));
  NOR2_X1    g16592(.A1(new_n16887_), .A2(new_n16889_), .ZN(new_n16890_));
  NOR2_X1    g16593(.A1(new_n16876_), .A2(new_n16890_), .ZN(new_n16891_));
  NOR2_X1    g16594(.A1(new_n16885_), .A2(new_n16891_), .ZN(new_n16892_));
  AOI22_X1   g16595(.A1(new_n13078_), .A2(\b[11] ), .B1(new_n927_), .B2(new_n12218_), .ZN(new_n16893_));
  OAI21_X1   g16596(.A1(new_n16893_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n16894_));
  XOR2_X1    g16597(.A1(new_n860_), .A2(new_n16894_), .Z(new_n16895_));
  INV_X1     g16598(.I(new_n16895_), .ZN(new_n16896_));
  NAND2_X1   g16599(.A1(new_n16892_), .A2(new_n16896_), .ZN(new_n16897_));
  INV_X1     g16600(.I(new_n16897_), .ZN(new_n16898_));
  NOR2_X1    g16601(.A1(new_n16892_), .A2(new_n16896_), .ZN(new_n16899_));
  OAI21_X1   g16602(.A1(new_n16898_), .A2(new_n16899_), .B(new_n16873_), .ZN(new_n16900_));
  XOR2_X1    g16603(.A1(new_n16892_), .A2(new_n16895_), .Z(new_n16901_));
  OAI21_X1   g16604(.A1(new_n16873_), .A2(new_n16901_), .B(new_n16900_), .ZN(new_n16902_));
  NAND2_X1   g16605(.A1(new_n16592_), .A2(new_n16589_), .ZN(new_n16903_));
  NAND2_X1   g16606(.A1(new_n16903_), .A2(new_n16590_), .ZN(new_n16904_));
  AND2_X2    g16607(.A1(new_n16902_), .A2(new_n16904_), .Z(new_n16905_));
  NOR2_X1    g16608(.A1(new_n16902_), .A2(new_n16904_), .ZN(new_n16906_));
  NOR2_X1    g16609(.A1(new_n16905_), .A2(new_n16906_), .ZN(new_n16907_));
  XOR2_X1    g16610(.A1(new_n16902_), .A2(new_n16904_), .Z(new_n16908_));
  NAND2_X1   g16611(.A1(new_n16908_), .A2(new_n16870_), .ZN(new_n16909_));
  OAI21_X1   g16612(.A1(new_n16870_), .A2(new_n16907_), .B(new_n16909_), .ZN(new_n16910_));
  INV_X1     g16613(.I(new_n16601_), .ZN(new_n16911_));
  OAI21_X1   g16614(.A1(new_n16602_), .A2(new_n16603_), .B(new_n16557_), .ZN(new_n16912_));
  AOI22_X1   g16615(.A1(new_n11415_), .A2(new_n1520_), .B1(\b[17] ), .B2(new_n10145_), .ZN(new_n16913_));
  OAI21_X1   g16616(.A1(new_n16913_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n16914_));
  XOR2_X1    g16617(.A1(new_n1421_), .A2(new_n16914_), .Z(new_n16915_));
  AOI21_X1   g16618(.A1(new_n16912_), .A2(new_n16911_), .B(new_n16915_), .ZN(new_n16916_));
  NAND2_X1   g16619(.A1(new_n16912_), .A2(new_n16911_), .ZN(new_n16917_));
  INV_X1     g16620(.I(new_n16915_), .ZN(new_n16918_));
  NOR2_X1    g16621(.A1(new_n16917_), .A2(new_n16918_), .ZN(new_n16919_));
  OAI21_X1   g16622(.A1(new_n16919_), .A2(new_n16916_), .B(new_n16910_), .ZN(new_n16920_));
  XOR2_X1    g16623(.A1(new_n16917_), .A2(new_n16915_), .Z(new_n16921_));
  OAI21_X1   g16624(.A1(new_n16921_), .A2(new_n16910_), .B(new_n16920_), .ZN(new_n16922_));
  INV_X1     g16625(.I(new_n16922_), .ZN(new_n16923_));
  NOR2_X1    g16626(.A1(new_n16923_), .A2(new_n16867_), .ZN(new_n16924_));
  INV_X1     g16627(.I(new_n16867_), .ZN(new_n16925_));
  NOR2_X1    g16628(.A1(new_n16925_), .A2(new_n16922_), .ZN(new_n16926_));
  OAI21_X1   g16629(.A1(new_n16924_), .A2(new_n16926_), .B(new_n16863_), .ZN(new_n16927_));
  XOR2_X1    g16630(.A1(new_n16922_), .A2(new_n16867_), .Z(new_n16928_));
  OAI21_X1   g16631(.A1(new_n16928_), .A2(new_n16863_), .B(new_n16927_), .ZN(new_n16929_));
  OAI22_X1   g16632(.A1(new_n7619_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n8309_), .ZN(new_n16930_));
  OAI21_X1   g16633(.A1(new_n1936_), .A2(new_n7947_), .B(new_n16930_), .ZN(new_n16931_));
  AOI21_X1   g16634(.A1(new_n16931_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n16932_));
  XNOR2_X1   g16635(.A1(new_n2280_), .A2(new_n16932_), .ZN(new_n16933_));
  INV_X1     g16636(.I(new_n16933_), .ZN(new_n16934_));
  NAND2_X1   g16637(.A1(new_n16929_), .A2(new_n16934_), .ZN(new_n16935_));
  NOR2_X1    g16638(.A1(new_n16929_), .A2(new_n16934_), .ZN(new_n16936_));
  INV_X1     g16639(.I(new_n16936_), .ZN(new_n16937_));
  AOI21_X1   g16640(.A1(new_n16937_), .A2(new_n16935_), .B(new_n16860_), .ZN(new_n16938_));
  XOR2_X1    g16641(.A1(new_n16929_), .A2(new_n16933_), .Z(new_n16939_));
  INV_X1     g16642(.I(new_n16939_), .ZN(new_n16940_));
  AOI21_X1   g16643(.A1(new_n16940_), .A2(new_n16860_), .B(new_n16938_), .ZN(new_n16941_));
  OAI21_X1   g16644(.A1(new_n16636_), .A2(new_n16639_), .B(new_n16637_), .ZN(new_n16942_));
  OAI22_X1   g16645(.A1(new_n6644_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n6647_), .ZN(new_n16943_));
  OAI21_X1   g16646(.A1(new_n2439_), .A2(new_n7284_), .B(new_n16943_), .ZN(new_n16944_));
  AOI21_X1   g16647(.A1(new_n2846_), .A2(new_n6631_), .B(new_n16944_), .ZN(new_n16945_));
  XOR2_X1    g16648(.A1(new_n16942_), .A2(new_n16945_), .Z(new_n16946_));
  XOR2_X1    g16649(.A1(new_n16946_), .A2(new_n16941_), .Z(new_n16947_));
  XOR2_X1    g16650(.A1(new_n16947_), .A2(new_n6632_), .Z(new_n16948_));
  OAI22_X1   g16651(.A1(new_n5993_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n5991_), .ZN(new_n16949_));
  OAI21_X1   g16652(.A1(new_n3018_), .A2(new_n5997_), .B(new_n16949_), .ZN(new_n16950_));
  AOI21_X1   g16653(.A1(new_n16950_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n16951_));
  XNOR2_X1   g16654(.A1(new_n3514_), .A2(new_n16951_), .ZN(new_n16952_));
  XOR2_X1    g16655(.A1(new_n16948_), .A2(new_n16952_), .Z(new_n16953_));
  XOR2_X1    g16656(.A1(new_n16947_), .A2(\a[44] ), .Z(new_n16954_));
  NOR2_X1    g16657(.A1(new_n16954_), .A2(new_n16952_), .ZN(new_n16955_));
  INV_X1     g16658(.I(new_n16952_), .ZN(new_n16956_));
  NOR2_X1    g16659(.A1(new_n16948_), .A2(new_n16956_), .ZN(new_n16957_));
  OAI21_X1   g16660(.A1(new_n16955_), .A2(new_n16957_), .B(new_n16858_), .ZN(new_n16958_));
  OAI21_X1   g16661(.A1(new_n16953_), .A2(new_n16858_), .B(new_n16958_), .ZN(new_n16959_));
  NAND2_X1   g16662(.A1(new_n16658_), .A2(new_n16543_), .ZN(new_n16960_));
  NAND2_X1   g16663(.A1(new_n16960_), .A2(new_n16656_), .ZN(new_n16961_));
  INV_X1     g16664(.I(new_n4257_), .ZN(new_n16962_));
  AOI22_X1   g16665(.A1(new_n4859_), .A2(\b[33] ), .B1(new_n4865_), .B2(\b[34] ), .ZN(new_n16963_));
  AOI21_X1   g16666(.A1(\b[32] ), .A2(new_n6005_), .B(new_n16963_), .ZN(new_n16964_));
  OAI21_X1   g16667(.A1(new_n16962_), .A2(new_n5420_), .B(new_n16964_), .ZN(new_n16965_));
  XOR2_X1    g16668(.A1(new_n16961_), .A2(new_n16965_), .Z(new_n16966_));
  XOR2_X1    g16669(.A1(new_n16966_), .A2(new_n16959_), .Z(new_n16967_));
  NOR2_X1    g16670(.A1(new_n16967_), .A2(\a[38] ), .ZN(new_n16968_));
  XNOR2_X1   g16671(.A1(new_n16966_), .A2(new_n16959_), .ZN(new_n16969_));
  NOR2_X1    g16672(.A1(new_n16969_), .A2(new_n4860_), .ZN(new_n16970_));
  NOR2_X1    g16673(.A1(new_n16970_), .A2(new_n16968_), .ZN(new_n16971_));
  OAI22_X1   g16674(.A1(new_n4072_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n4067_), .ZN(new_n16972_));
  OAI21_X1   g16675(.A1(new_n4500_), .A2(new_n4318_), .B(new_n16972_), .ZN(new_n16973_));
  AOI21_X1   g16676(.A1(new_n16973_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n16974_));
  XOR2_X1    g16677(.A1(new_n5067_), .A2(new_n16974_), .Z(new_n16975_));
  INV_X1     g16678(.I(new_n16975_), .ZN(new_n16976_));
  NAND2_X1   g16679(.A1(new_n16971_), .A2(new_n16976_), .ZN(new_n16977_));
  NAND2_X1   g16680(.A1(new_n16969_), .A2(new_n4860_), .ZN(new_n16978_));
  NAND2_X1   g16681(.A1(new_n16967_), .A2(\a[38] ), .ZN(new_n16979_));
  NAND2_X1   g16682(.A1(new_n16978_), .A2(new_n16979_), .ZN(new_n16980_));
  NAND2_X1   g16683(.A1(new_n16980_), .A2(new_n16975_), .ZN(new_n16981_));
  AOI21_X1   g16684(.A1(new_n16977_), .A2(new_n16981_), .B(new_n16856_), .ZN(new_n16982_));
  INV_X1     g16685(.I(new_n16856_), .ZN(new_n16983_));
  NAND2_X1   g16686(.A1(new_n16980_), .A2(new_n16976_), .ZN(new_n16984_));
  NAND2_X1   g16687(.A1(new_n16971_), .A2(new_n16975_), .ZN(new_n16985_));
  AOI21_X1   g16688(.A1(new_n16985_), .A2(new_n16984_), .B(new_n16983_), .ZN(new_n16986_));
  OAI22_X1   g16689(.A1(new_n5913_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n5921_), .ZN(new_n16987_));
  OAI21_X1   g16690(.A1(new_n5353_), .A2(new_n3569_), .B(new_n16987_), .ZN(new_n16988_));
  AOI21_X1   g16691(.A1(new_n16988_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n16989_));
  XOR2_X1    g16692(.A1(new_n5926_), .A2(new_n16989_), .Z(new_n16990_));
  INV_X1     g16693(.I(new_n16990_), .ZN(new_n16991_));
  OAI21_X1   g16694(.A1(new_n16982_), .A2(new_n16986_), .B(new_n16991_), .ZN(new_n16992_));
  NOR2_X1    g16695(.A1(new_n16982_), .A2(new_n16986_), .ZN(new_n16993_));
  NAND2_X1   g16696(.A1(new_n16993_), .A2(new_n16990_), .ZN(new_n16994_));
  AOI21_X1   g16697(.A1(new_n16994_), .A2(new_n16992_), .B(new_n16855_), .ZN(new_n16995_));
  INV_X1     g16698(.I(new_n16855_), .ZN(new_n16996_));
  NAND2_X1   g16699(.A1(new_n16993_), .A2(new_n16991_), .ZN(new_n16997_));
  OAI21_X1   g16700(.A1(new_n16982_), .A2(new_n16986_), .B(new_n16990_), .ZN(new_n16998_));
  AOI21_X1   g16701(.A1(new_n16997_), .A2(new_n16998_), .B(new_n16996_), .ZN(new_n16999_));
  OAI22_X1   g16702(.A1(new_n6538_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n6847_), .ZN(new_n17000_));
  OAI21_X1   g16703(.A1(new_n6229_), .A2(new_n2884_), .B(new_n17000_), .ZN(new_n17001_));
  AOI21_X1   g16704(.A1(new_n17001_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n17002_));
  XOR2_X1    g16705(.A1(new_n6851_), .A2(new_n17002_), .Z(new_n17003_));
  INV_X1     g16706(.I(new_n17003_), .ZN(new_n17004_));
  OAI21_X1   g16707(.A1(new_n16995_), .A2(new_n16999_), .B(new_n17004_), .ZN(new_n17005_));
  NOR2_X1    g16708(.A1(new_n16995_), .A2(new_n16999_), .ZN(new_n17006_));
  NAND2_X1   g16709(.A1(new_n17006_), .A2(new_n17003_), .ZN(new_n17007_));
  AOI21_X1   g16710(.A1(new_n17007_), .A2(new_n17005_), .B(new_n16850_), .ZN(new_n17008_));
  INV_X1     g16711(.I(new_n16850_), .ZN(new_n17009_));
  NAND2_X1   g16712(.A1(new_n17006_), .A2(new_n17004_), .ZN(new_n17010_));
  OAI21_X1   g16713(.A1(new_n16995_), .A2(new_n16999_), .B(new_n17003_), .ZN(new_n17011_));
  AOI21_X1   g16714(.A1(new_n17010_), .A2(new_n17011_), .B(new_n17009_), .ZN(new_n17012_));
  OAI22_X1   g16715(.A1(new_n2171_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n2166_), .ZN(new_n17013_));
  OAI21_X1   g16716(.A1(new_n7198_), .A2(new_n2322_), .B(new_n17013_), .ZN(new_n17014_));
  AOI21_X1   g16717(.A1(new_n17014_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n17015_));
  XNOR2_X1   g16718(.A1(new_n7874_), .A2(new_n17015_), .ZN(new_n17016_));
  INV_X1     g16719(.I(new_n17016_), .ZN(new_n17017_));
  OAI21_X1   g16720(.A1(new_n17012_), .A2(new_n17008_), .B(new_n17017_), .ZN(new_n17018_));
  NOR3_X1    g16721(.A1(new_n17008_), .A2(new_n17012_), .A3(new_n17017_), .ZN(new_n17019_));
  INV_X1     g16722(.I(new_n17019_), .ZN(new_n17020_));
  AOI21_X1   g16723(.A1(new_n17020_), .A2(new_n17018_), .B(new_n16849_), .ZN(new_n17021_));
  OR3_X2     g16724(.A1(new_n17008_), .A2(new_n17012_), .A3(new_n17016_), .Z(new_n17022_));
  OAI21_X1   g16725(.A1(new_n17012_), .A2(new_n17008_), .B(new_n17016_), .ZN(new_n17023_));
  AOI21_X1   g16726(.A1(new_n17022_), .A2(new_n17023_), .B(new_n16848_), .ZN(new_n17024_));
  OAI22_X1   g16727(.A1(new_n1712_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n1707_), .ZN(new_n17025_));
  OAI21_X1   g16728(.A1(new_n8218_), .A2(new_n1850_), .B(new_n17025_), .ZN(new_n17026_));
  AOI21_X1   g16729(.A1(new_n17026_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n17027_));
  XOR2_X1    g16730(.A1(new_n8952_), .A2(new_n17027_), .Z(new_n17028_));
  INV_X1     g16731(.I(new_n17028_), .ZN(new_n17029_));
  OAI21_X1   g16732(.A1(new_n17021_), .A2(new_n17024_), .B(new_n17029_), .ZN(new_n17030_));
  NOR2_X1    g16733(.A1(new_n17021_), .A2(new_n17024_), .ZN(new_n17031_));
  NAND2_X1   g16734(.A1(new_n17031_), .A2(new_n17028_), .ZN(new_n17032_));
  NAND2_X1   g16735(.A1(new_n17032_), .A2(new_n17030_), .ZN(new_n17033_));
  NAND2_X1   g16736(.A1(new_n17033_), .A2(new_n16845_), .ZN(new_n17034_));
  XOR2_X1    g16737(.A1(new_n17031_), .A2(new_n17028_), .Z(new_n17035_));
  NAND2_X1   g16738(.A1(new_n17035_), .A2(new_n16844_), .ZN(new_n17036_));
  OAI22_X1   g16739(.A1(new_n1347_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n1344_), .ZN(new_n17037_));
  OAI21_X1   g16740(.A1(new_n9295_), .A2(new_n1457_), .B(new_n17037_), .ZN(new_n17038_));
  AOI21_X1   g16741(.A1(new_n17038_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n17039_));
  XNOR2_X1   g16742(.A1(new_n10035_), .A2(new_n17039_), .ZN(new_n17040_));
  AOI21_X1   g16743(.A1(new_n17036_), .A2(new_n17034_), .B(new_n17040_), .ZN(new_n17041_));
  NAND2_X1   g16744(.A1(new_n17036_), .A2(new_n17034_), .ZN(new_n17042_));
  INV_X1     g16745(.I(new_n17040_), .ZN(new_n17043_));
  NOR2_X1    g16746(.A1(new_n17042_), .A2(new_n17043_), .ZN(new_n17044_));
  OAI21_X1   g16747(.A1(new_n17044_), .A2(new_n17041_), .B(new_n16842_), .ZN(new_n17045_));
  NOR2_X1    g16748(.A1(new_n17042_), .A2(new_n17040_), .ZN(new_n17046_));
  AOI21_X1   g16749(.A1(new_n17036_), .A2(new_n17034_), .B(new_n17043_), .ZN(new_n17047_));
  OAI21_X1   g16750(.A1(new_n17046_), .A2(new_n17047_), .B(new_n16841_), .ZN(new_n17048_));
  NAND2_X1   g16751(.A1(new_n17045_), .A2(new_n17048_), .ZN(new_n17049_));
  OAI22_X1   g16752(.A1(new_n1055_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n1061_), .ZN(new_n17050_));
  OAI21_X1   g16753(.A1(new_n10477_), .A2(new_n1332_), .B(new_n17050_), .ZN(new_n17051_));
  AOI21_X1   g16754(.A1(new_n17051_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n17052_));
  XOR2_X1    g16755(.A1(new_n11298_), .A2(new_n17052_), .Z(new_n17053_));
  XOR2_X1    g16756(.A1(new_n17049_), .A2(new_n17053_), .Z(new_n17054_));
  NOR2_X1    g16757(.A1(new_n17054_), .A2(new_n16839_), .ZN(new_n17055_));
  INV_X1     g16758(.I(new_n17053_), .ZN(new_n17056_));
  NAND2_X1   g16759(.A1(new_n17049_), .A2(new_n17056_), .ZN(new_n17057_));
  NAND3_X1   g16760(.A1(new_n17045_), .A2(new_n17048_), .A3(new_n17053_), .ZN(new_n17058_));
  AOI21_X1   g16761(.A1(new_n17057_), .A2(new_n17058_), .B(new_n16838_), .ZN(new_n17059_));
  NOR2_X1    g16762(.A1(new_n17055_), .A2(new_n17059_), .ZN(new_n17060_));
  OAI22_X1   g16763(.A1(new_n970_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n820_), .ZN(new_n17061_));
  OAI21_X1   g16764(.A1(new_n11744_), .A2(new_n894_), .B(new_n17061_), .ZN(new_n17062_));
  AOI21_X1   g16765(.A1(new_n17062_), .A2(new_n827_), .B(new_n970_), .ZN(new_n17063_));
  XNOR2_X1   g16766(.A1(new_n12546_), .A2(new_n17063_), .ZN(new_n17064_));
  INV_X1     g16767(.I(new_n17064_), .ZN(new_n17065_));
  NAND2_X1   g16768(.A1(new_n17060_), .A2(new_n17065_), .ZN(new_n17066_));
  INV_X1     g16769(.I(new_n17059_), .ZN(new_n17067_));
  OAI21_X1   g16770(.A1(new_n16839_), .A2(new_n17054_), .B(new_n17067_), .ZN(new_n17068_));
  NAND2_X1   g16771(.A1(new_n17068_), .A2(new_n17064_), .ZN(new_n17069_));
  NAND2_X1   g16772(.A1(new_n17066_), .A2(new_n17069_), .ZN(new_n17070_));
  NAND2_X1   g16773(.A1(new_n17070_), .A2(new_n16836_), .ZN(new_n17071_));
  NOR2_X1    g16774(.A1(new_n17060_), .A2(new_n17064_), .ZN(new_n17072_));
  NOR2_X1    g16775(.A1(new_n17068_), .A2(new_n17065_), .ZN(new_n17073_));
  OAI21_X1   g16776(.A1(new_n17072_), .A2(new_n17073_), .B(new_n16835_), .ZN(new_n17074_));
  NAND2_X1   g16777(.A1(new_n17071_), .A2(new_n17074_), .ZN(new_n17075_));
  OAI22_X1   g16778(.A1(new_n607_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n610_), .ZN(new_n17076_));
  OAI21_X1   g16779(.A1(new_n12970_), .A2(new_n684_), .B(new_n17076_), .ZN(new_n17077_));
  AOI21_X1   g16780(.A1(new_n17077_), .A2(new_n612_), .B(new_n607_), .ZN(new_n17078_));
  XOR2_X1    g16781(.A1(new_n13784_), .A2(new_n17078_), .Z(new_n17079_));
  NOR2_X1    g16782(.A1(new_n17075_), .A2(new_n17079_), .ZN(new_n17080_));
  INV_X1     g16783(.I(new_n17079_), .ZN(new_n17081_));
  AOI21_X1   g16784(.A1(new_n17071_), .A2(new_n17074_), .B(new_n17081_), .ZN(new_n17082_));
  OAI21_X1   g16785(.A1(new_n17080_), .A2(new_n17082_), .B(new_n16833_), .ZN(new_n17083_));
  AOI21_X1   g16786(.A1(new_n17071_), .A2(new_n17074_), .B(new_n17079_), .ZN(new_n17084_));
  NOR2_X1    g16787(.A1(new_n17075_), .A2(new_n17081_), .ZN(new_n17085_));
  OAI21_X1   g16788(.A1(new_n17085_), .A2(new_n17084_), .B(new_n16832_), .ZN(new_n17086_));
  NAND2_X1   g16789(.A1(new_n17083_), .A2(new_n17086_), .ZN(new_n17087_));
  NOR2_X1    g16790(.A1(new_n496_), .A2(new_n450_), .ZN(new_n17088_));
  NAND2_X1   g16791(.A1(new_n16148_), .A2(new_n452_), .ZN(new_n17089_));
  OAI21_X1   g16792(.A1(new_n17088_), .A2(new_n17089_), .B(new_n447_), .ZN(new_n17090_));
  XNOR2_X1   g16793(.A1(new_n14978_), .A2(new_n17090_), .ZN(new_n17091_));
  NOR2_X1    g16794(.A1(new_n17087_), .A2(new_n17091_), .ZN(new_n17092_));
  INV_X1     g16795(.I(new_n17091_), .ZN(new_n17093_));
  AOI21_X1   g16796(.A1(new_n17083_), .A2(new_n17086_), .B(new_n17093_), .ZN(new_n17094_));
  OAI21_X1   g16797(.A1(new_n17092_), .A2(new_n17094_), .B(new_n16831_), .ZN(new_n17095_));
  XOR2_X1    g16798(.A1(new_n17087_), .A2(new_n17093_), .Z(new_n17096_));
  OAI21_X1   g16799(.A1(new_n17096_), .A2(new_n16831_), .B(new_n17095_), .ZN(new_n17097_));
  NOR3_X1    g16800(.A1(new_n16796_), .A2(new_n16800_), .A3(new_n16805_), .ZN(new_n17098_));
  NOR2_X1    g16801(.A1(new_n16514_), .A2(new_n17098_), .ZN(new_n17099_));
  INV_X1     g16802(.I(new_n17099_), .ZN(new_n17100_));
  NAND2_X1   g16803(.A1(new_n17100_), .A2(new_n16806_), .ZN(new_n17101_));
  XOR2_X1    g16804(.A1(new_n17097_), .A2(new_n17101_), .Z(new_n17102_));
  INV_X1     g16805(.I(new_n16166_), .ZN(new_n17103_));
  AOI21_X1   g16806(.A1(new_n15830_), .A2(new_n16165_), .B(new_n15814_), .ZN(new_n17104_));
  NAND4_X1   g16807(.A1(new_n15825_), .A2(new_n15817_), .A3(new_n15826_), .A4(new_n17104_), .ZN(new_n17105_));
  OAI21_X1   g16808(.A1(new_n16497_), .A2(new_n16498_), .B(new_n334_), .ZN(new_n17106_));
  NAND3_X1   g16809(.A1(new_n16492_), .A2(new_n16495_), .A3(\a[5] ), .ZN(new_n17107_));
  NOR3_X1    g16810(.A1(new_n16824_), .A2(new_n16822_), .A3(new_n16821_), .ZN(new_n17108_));
  AOI21_X1   g16811(.A1(new_n16512_), .A2(new_n16509_), .B(new_n16819_), .ZN(new_n17109_));
  NOR2_X1    g16812(.A1(new_n17109_), .A2(new_n17108_), .ZN(new_n17110_));
  NAND3_X1   g16813(.A1(new_n17110_), .A2(new_n17106_), .A3(new_n17107_), .ZN(new_n17111_));
  AOI21_X1   g16814(.A1(new_n17106_), .A2(new_n17107_), .B(new_n17110_), .ZN(new_n17112_));
  OAI21_X1   g16815(.A1(new_n17112_), .A2(new_n16183_), .B(new_n17111_), .ZN(new_n17113_));
  AOI21_X1   g16816(.A1(new_n17105_), .A2(new_n17103_), .B(new_n17113_), .ZN(new_n17114_));
  NOR3_X1    g16817(.A1(new_n16819_), .A2(new_n16821_), .A3(new_n16822_), .ZN(new_n17115_));
  NOR2_X1    g16818(.A1(new_n17114_), .A2(new_n17115_), .ZN(new_n17116_));
  INV_X1     g16819(.I(new_n17115_), .ZN(new_n17117_));
  NAND2_X1   g16820(.A1(new_n17102_), .A2(new_n17117_), .ZN(new_n17118_));
  OAI22_X1   g16821(.A1(new_n17116_), .A2(new_n17102_), .B1(new_n17114_), .B2(new_n17118_), .ZN(\f[70] ));
  NOR3_X1    g16822(.A1(new_n16826_), .A2(new_n16496_), .A3(new_n16499_), .ZN(new_n17120_));
  OAI21_X1   g16823(.A1(new_n16496_), .A2(new_n16499_), .B(new_n16826_), .ZN(new_n17121_));
  AOI21_X1   g16824(.A1(new_n17121_), .A2(new_n16182_), .B(new_n17120_), .ZN(new_n17122_));
  OAI21_X1   g16825(.A1(new_n16179_), .A2(new_n16166_), .B(new_n17122_), .ZN(new_n17123_));
  INV_X1     g16826(.I(new_n17097_), .ZN(new_n17124_));
  NOR2_X1    g16827(.A1(new_n17124_), .A2(new_n17117_), .ZN(new_n17125_));
  INV_X1     g16828(.I(new_n17125_), .ZN(new_n17126_));
  OAI21_X1   g16829(.A1(new_n17097_), .A2(new_n17115_), .B(new_n17101_), .ZN(new_n17127_));
  OAI21_X1   g16830(.A1(new_n17123_), .A2(new_n17127_), .B(new_n17126_), .ZN(new_n17128_));
  INV_X1     g16831(.I(new_n17094_), .ZN(new_n17129_));
  AOI21_X1   g16832(.A1(new_n16831_), .A2(new_n17129_), .B(new_n17092_), .ZN(new_n17130_));
  INV_X1     g16833(.I(new_n17130_), .ZN(new_n17131_));
  NAND2_X1   g16834(.A1(new_n17058_), .A2(new_n16838_), .ZN(new_n17132_));
  NAND2_X1   g16835(.A1(new_n17132_), .A2(new_n17057_), .ZN(new_n17133_));
  OAI21_X1   g16836(.A1(new_n17042_), .A2(new_n17043_), .B(new_n16842_), .ZN(new_n17134_));
  INV_X1     g16837(.I(new_n17134_), .ZN(new_n17135_));
  NAND2_X1   g16838(.A1(new_n17032_), .A2(new_n16845_), .ZN(new_n17136_));
  OAI21_X1   g16839(.A1(new_n17019_), .A2(new_n16849_), .B(new_n17018_), .ZN(new_n17137_));
  NAND2_X1   g16840(.A1(new_n17007_), .A2(new_n17009_), .ZN(new_n17138_));
  NAND2_X1   g16841(.A1(new_n17138_), .A2(new_n17005_), .ZN(new_n17139_));
  INV_X1     g16842(.I(new_n17139_), .ZN(new_n17140_));
  NAND2_X1   g16843(.A1(new_n16994_), .A2(new_n16996_), .ZN(new_n17141_));
  NAND2_X1   g16844(.A1(new_n17141_), .A2(new_n16992_), .ZN(new_n17142_));
  NAND2_X1   g16845(.A1(new_n16981_), .A2(new_n16983_), .ZN(new_n17143_));
  INV_X1     g16846(.I(new_n16858_), .ZN(new_n17144_));
  INV_X1     g16847(.I(new_n16957_), .ZN(new_n17145_));
  AOI21_X1   g16848(.A1(new_n17145_), .A2(new_n17144_), .B(new_n16955_), .ZN(new_n17146_));
  INV_X1     g16849(.I(new_n17146_), .ZN(new_n17147_));
  INV_X1     g16850(.I(new_n16941_), .ZN(new_n17148_));
  INV_X1     g16851(.I(new_n16942_), .ZN(new_n17149_));
  XOR2_X1    g16852(.A1(new_n16945_), .A2(new_n6632_), .Z(new_n17150_));
  AOI21_X1   g16853(.A1(new_n17149_), .A2(new_n16941_), .B(new_n17150_), .ZN(new_n17151_));
  AOI21_X1   g16854(.A1(new_n17148_), .A2(new_n16942_), .B(new_n17151_), .ZN(new_n17152_));
  OAI21_X1   g16855(.A1(new_n16860_), .A2(new_n16936_), .B(new_n16935_), .ZN(new_n17153_));
  NOR2_X1    g16856(.A1(new_n16926_), .A2(new_n16862_), .ZN(new_n17154_));
  NOR2_X1    g16857(.A1(new_n17154_), .A2(new_n16924_), .ZN(new_n17155_));
  INV_X1     g16858(.I(new_n17155_), .ZN(new_n17156_));
  OAI22_X1   g16859(.A1(new_n7619_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n8309_), .ZN(new_n17157_));
  OAI21_X1   g16860(.A1(new_n2102_), .A2(new_n7947_), .B(new_n17157_), .ZN(new_n17158_));
  AOI21_X1   g16861(.A1(new_n17158_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n17159_));
  INV_X1     g16862(.I(new_n17159_), .ZN(new_n17160_));
  NOR2_X1    g16863(.A1(new_n2443_), .A2(new_n17160_), .ZN(new_n17161_));
  AND2_X2    g16864(.A1(new_n2443_), .A2(new_n17160_), .Z(new_n17162_));
  OAI22_X1   g16865(.A1(new_n8644_), .A2(new_n1803_), .B1(new_n1936_), .B2(new_n9388_), .ZN(new_n17163_));
  OAI21_X1   g16866(.A1(new_n1634_), .A2(new_n10154_), .B(new_n17163_), .ZN(new_n17164_));
  AOI21_X1   g16867(.A1(new_n17164_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n17165_));
  XNOR2_X1   g16868(.A1(new_n1940_), .A2(new_n17165_), .ZN(new_n17166_));
  AOI22_X1   g16869(.A1(new_n11415_), .A2(new_n1527_), .B1(\b[18] ), .B2(new_n10145_), .ZN(new_n17167_));
  OAI21_X1   g16870(.A1(new_n17167_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n17168_));
  XNOR2_X1   g16871(.A1(new_n1530_), .A2(new_n17168_), .ZN(new_n17169_));
  INV_X1     g16872(.I(new_n16889_), .ZN(new_n17170_));
  OAI21_X1   g16873(.A1(new_n16877_), .A2(new_n16887_), .B(new_n17170_), .ZN(new_n17171_));
  NOR2_X1    g16874(.A1(new_n13476_), .A2(new_n472_), .ZN(new_n17172_));
  XOR2_X1    g16875(.A1(new_n14736_), .A2(new_n472_), .Z(new_n17173_));
  NAND2_X1   g16876(.A1(new_n17173_), .A2(\b[8] ), .ZN(new_n17174_));
  XOR2_X1    g16877(.A1(new_n17174_), .A2(new_n17172_), .Z(new_n17175_));
  NOR2_X1    g16878(.A1(new_n16888_), .A2(new_n17175_), .ZN(new_n17176_));
  INV_X1     g16879(.I(new_n17175_), .ZN(new_n17177_));
  NOR2_X1    g16880(.A1(new_n17177_), .A2(new_n16883_), .ZN(new_n17178_));
  NOR2_X1    g16881(.A1(new_n17176_), .A2(new_n17178_), .ZN(new_n17179_));
  INV_X1     g16882(.I(new_n17179_), .ZN(new_n17180_));
  XOR2_X1    g16883(.A1(new_n16883_), .A2(new_n17175_), .Z(new_n17181_));
  NOR2_X1    g16884(.A1(new_n17171_), .A2(new_n17181_), .ZN(new_n17182_));
  AOI21_X1   g16885(.A1(new_n17171_), .A2(new_n17180_), .B(new_n17182_), .ZN(new_n17183_));
  INV_X1     g16886(.I(new_n17183_), .ZN(new_n17184_));
  AOI22_X1   g16887(.A1(new_n13078_), .A2(\b[12] ), .B1(new_n932_), .B2(new_n12218_), .ZN(new_n17185_));
  OAI21_X1   g16888(.A1(new_n17185_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n17186_));
  INV_X1     g16889(.I(new_n17186_), .ZN(new_n17187_));
  XOR2_X1    g16890(.A1(new_n937_), .A2(new_n17187_), .Z(new_n17188_));
  OAI22_X1   g16891(.A1(new_n13880_), .A2(new_n772_), .B1(new_n565_), .B2(new_n13885_), .ZN(new_n17189_));
  AOI21_X1   g16892(.A1(new_n17189_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n17190_));
  XNOR2_X1   g16893(.A1(new_n710_), .A2(new_n17190_), .ZN(new_n17191_));
  INV_X1     g16894(.I(new_n17191_), .ZN(new_n17192_));
  XOR2_X1    g16895(.A1(new_n17188_), .A2(new_n17192_), .Z(new_n17193_));
  NAND2_X1   g16896(.A1(new_n17188_), .A2(new_n17192_), .ZN(new_n17194_));
  OR2_X2     g16897(.A1(new_n17188_), .A2(new_n17192_), .Z(new_n17195_));
  AOI21_X1   g16898(.A1(new_n17195_), .A2(new_n17194_), .B(new_n17184_), .ZN(new_n17196_));
  AOI21_X1   g16899(.A1(new_n17184_), .A2(new_n17193_), .B(new_n17196_), .ZN(new_n17197_));
  AOI22_X1   g16900(.A1(new_n10969_), .A2(new_n1292_), .B1(new_n11394_), .B2(\b[15] ), .ZN(new_n17198_));
  OAI21_X1   g16901(.A1(new_n17198_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n17199_));
  XNOR2_X1   g16902(.A1(new_n1196_), .A2(new_n17199_), .ZN(new_n17200_));
  OAI21_X1   g16903(.A1(new_n16872_), .A2(new_n16899_), .B(new_n16897_), .ZN(new_n17201_));
  XNOR2_X1   g16904(.A1(new_n17200_), .A2(new_n17201_), .ZN(new_n17202_));
  NOR2_X1    g16905(.A1(new_n17202_), .A2(new_n17197_), .ZN(new_n17203_));
  NAND2_X1   g16906(.A1(new_n17200_), .A2(new_n17201_), .ZN(new_n17204_));
  OR2_X2     g16907(.A1(new_n17200_), .A2(new_n17201_), .Z(new_n17205_));
  NAND2_X1   g16908(.A1(new_n17205_), .A2(new_n17204_), .ZN(new_n17206_));
  AND2_X2    g16909(.A1(new_n17206_), .A2(new_n17197_), .Z(new_n17207_));
  NOR2_X1    g16910(.A1(new_n17207_), .A2(new_n17203_), .ZN(new_n17208_));
  NOR2_X1    g16911(.A1(new_n16906_), .A2(new_n16870_), .ZN(new_n17209_));
  NOR2_X1    g16912(.A1(new_n17209_), .A2(new_n16905_), .ZN(new_n17210_));
  INV_X1     g16913(.I(new_n17210_), .ZN(new_n17211_));
  XOR2_X1    g16914(.A1(new_n17208_), .A2(new_n17211_), .Z(new_n17212_));
  NOR2_X1    g16915(.A1(new_n17212_), .A2(new_n17169_), .ZN(new_n17213_));
  INV_X1     g16916(.I(new_n17169_), .ZN(new_n17214_));
  OAI21_X1   g16917(.A1(new_n17203_), .A2(new_n17207_), .B(new_n17211_), .ZN(new_n17215_));
  NAND2_X1   g16918(.A1(new_n17208_), .A2(new_n17210_), .ZN(new_n17216_));
  AOI21_X1   g16919(.A1(new_n17216_), .A2(new_n17215_), .B(new_n17214_), .ZN(new_n17217_));
  NOR2_X1    g16920(.A1(new_n17213_), .A2(new_n17217_), .ZN(new_n17218_));
  INV_X1     g16921(.I(new_n16919_), .ZN(new_n17219_));
  AOI21_X1   g16922(.A1(new_n17219_), .A2(new_n16910_), .B(new_n16916_), .ZN(new_n17220_));
  XOR2_X1    g16923(.A1(new_n17218_), .A2(new_n17220_), .Z(new_n17221_));
  NOR2_X1    g16924(.A1(new_n17221_), .A2(new_n17166_), .ZN(new_n17222_));
  INV_X1     g16925(.I(new_n17166_), .ZN(new_n17223_));
  INV_X1     g16926(.I(new_n17220_), .ZN(new_n17224_));
  NAND2_X1   g16927(.A1(new_n17218_), .A2(new_n17224_), .ZN(new_n17225_));
  OAI21_X1   g16928(.A1(new_n17213_), .A2(new_n17217_), .B(new_n17220_), .ZN(new_n17226_));
  AOI21_X1   g16929(.A1(new_n17225_), .A2(new_n17226_), .B(new_n17223_), .ZN(new_n17227_));
  NOR2_X1    g16930(.A1(new_n17222_), .A2(new_n17227_), .ZN(new_n17228_));
  NOR3_X1    g16931(.A1(new_n17228_), .A2(new_n17161_), .A3(new_n17162_), .ZN(new_n17229_));
  NOR2_X1    g16932(.A1(new_n17162_), .A2(new_n17161_), .ZN(new_n17230_));
  NOR3_X1    g16933(.A1(new_n17222_), .A2(new_n17230_), .A3(new_n17227_), .ZN(new_n17231_));
  OAI21_X1   g16934(.A1(new_n17229_), .A2(new_n17231_), .B(new_n17156_), .ZN(new_n17232_));
  XOR2_X1    g16935(.A1(new_n17228_), .A2(new_n17230_), .Z(new_n17233_));
  OAI21_X1   g16936(.A1(new_n17233_), .A2(new_n17156_), .B(new_n17232_), .ZN(new_n17234_));
  OAI22_X1   g16937(.A1(new_n6644_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n6647_), .ZN(new_n17235_));
  OAI21_X1   g16938(.A1(new_n2643_), .A2(new_n7284_), .B(new_n17235_), .ZN(new_n17236_));
  AOI21_X1   g16939(.A1(new_n17236_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n17237_));
  XNOR2_X1   g16940(.A1(new_n3022_), .A2(new_n17237_), .ZN(new_n17238_));
  INV_X1     g16941(.I(new_n17238_), .ZN(new_n17239_));
  NAND2_X1   g16942(.A1(new_n17234_), .A2(new_n17239_), .ZN(new_n17240_));
  INV_X1     g16943(.I(new_n17240_), .ZN(new_n17241_));
  NOR2_X1    g16944(.A1(new_n17234_), .A2(new_n17239_), .ZN(new_n17242_));
  OAI21_X1   g16945(.A1(new_n17241_), .A2(new_n17242_), .B(new_n17153_), .ZN(new_n17243_));
  INV_X1     g16946(.I(new_n17153_), .ZN(new_n17244_));
  XOR2_X1    g16947(.A1(new_n17234_), .A2(new_n17239_), .Z(new_n17245_));
  NAND2_X1   g16948(.A1(new_n17245_), .A2(new_n17244_), .ZN(new_n17246_));
  NAND2_X1   g16949(.A1(new_n17246_), .A2(new_n17243_), .ZN(new_n17247_));
  OAI22_X1   g16950(.A1(new_n5993_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n5991_), .ZN(new_n17248_));
  OAI21_X1   g16951(.A1(new_n3260_), .A2(new_n5997_), .B(new_n17248_), .ZN(new_n17249_));
  AOI21_X1   g16952(.A1(new_n17249_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n17250_));
  XOR2_X1    g16953(.A1(new_n3722_), .A2(new_n17250_), .Z(new_n17251_));
  XOR2_X1    g16954(.A1(new_n17247_), .A2(new_n17251_), .Z(new_n17252_));
  INV_X1     g16955(.I(new_n17251_), .ZN(new_n17253_));
  NAND2_X1   g16956(.A1(new_n17247_), .A2(new_n17253_), .ZN(new_n17254_));
  INV_X1     g16957(.I(new_n17254_), .ZN(new_n17255_));
  NOR2_X1    g16958(.A1(new_n17247_), .A2(new_n17253_), .ZN(new_n17256_));
  OAI21_X1   g16959(.A1(new_n17255_), .A2(new_n17256_), .B(new_n17152_), .ZN(new_n17257_));
  OAI21_X1   g16960(.A1(new_n17152_), .A2(new_n17252_), .B(new_n17257_), .ZN(new_n17258_));
  OAI22_X1   g16961(.A1(new_n5420_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n5107_), .ZN(new_n17259_));
  OAI21_X1   g16962(.A1(new_n3989_), .A2(new_n5112_), .B(new_n17259_), .ZN(new_n17260_));
  AOI21_X1   g16963(.A1(new_n17260_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n17261_));
  XOR2_X1    g16964(.A1(new_n4499_), .A2(new_n17261_), .Z(new_n17262_));
  OR2_X2     g16965(.A1(new_n17258_), .A2(new_n17262_), .Z(new_n17263_));
  NAND2_X1   g16966(.A1(new_n17258_), .A2(new_n17262_), .ZN(new_n17264_));
  NAND2_X1   g16967(.A1(new_n17263_), .A2(new_n17264_), .ZN(new_n17265_));
  NAND2_X1   g16968(.A1(new_n17265_), .A2(new_n17147_), .ZN(new_n17266_));
  XNOR2_X1   g16969(.A1(new_n17258_), .A2(new_n17262_), .ZN(new_n17267_));
  OAI21_X1   g16970(.A1(new_n17147_), .A2(new_n17267_), .B(new_n17266_), .ZN(new_n17268_));
  NAND2_X1   g16971(.A1(new_n16959_), .A2(new_n16961_), .ZN(new_n17269_));
  XOR2_X1    g16972(.A1(new_n16965_), .A2(new_n4860_), .Z(new_n17270_));
  OAI21_X1   g16973(.A1(new_n16959_), .A2(new_n16961_), .B(new_n17270_), .ZN(new_n17271_));
  NAND2_X1   g16974(.A1(new_n17271_), .A2(new_n17269_), .ZN(new_n17272_));
  INV_X1     g16975(.I(new_n5357_), .ZN(new_n17273_));
  AOI22_X1   g16976(.A1(new_n4062_), .A2(\b[37] ), .B1(new_n5438_), .B2(\b[38] ), .ZN(new_n17274_));
  AOI21_X1   g16977(.A1(\b[36] ), .A2(new_n4319_), .B(new_n17274_), .ZN(new_n17275_));
  OAI21_X1   g16978(.A1(new_n17273_), .A2(new_n4072_), .B(new_n17275_), .ZN(new_n17276_));
  XOR2_X1    g16979(.A1(new_n17272_), .A2(new_n17276_), .Z(new_n17277_));
  XOR2_X1    g16980(.A1(new_n17277_), .A2(new_n17268_), .Z(new_n17278_));
  XOR2_X1    g16981(.A1(new_n17278_), .A2(new_n4069_), .Z(new_n17279_));
  INV_X1     g16982(.I(new_n17279_), .ZN(new_n17280_));
  OAI22_X1   g16983(.A1(new_n5921_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n6229_), .ZN(new_n17281_));
  OAI21_X1   g16984(.A1(new_n5913_), .A2(new_n3569_), .B(new_n17281_), .ZN(new_n17282_));
  AOI21_X1   g16985(.A1(new_n17282_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n17283_));
  XOR2_X1    g16986(.A1(new_n6233_), .A2(new_n17283_), .Z(new_n17284_));
  INV_X1     g16987(.I(new_n17284_), .ZN(new_n17285_));
  NAND2_X1   g16988(.A1(new_n17280_), .A2(new_n17285_), .ZN(new_n17286_));
  NAND2_X1   g16989(.A1(new_n17279_), .A2(new_n17284_), .ZN(new_n17287_));
  AOI22_X1   g16990(.A1(new_n17286_), .A2(new_n17287_), .B1(new_n16977_), .B2(new_n17143_), .ZN(new_n17288_));
  NAND2_X1   g16991(.A1(new_n17143_), .A2(new_n16977_), .ZN(new_n17289_));
  NAND2_X1   g16992(.A1(new_n17279_), .A2(new_n17285_), .ZN(new_n17290_));
  NAND2_X1   g16993(.A1(new_n17280_), .A2(new_n17284_), .ZN(new_n17291_));
  AOI21_X1   g16994(.A1(new_n17291_), .A2(new_n17290_), .B(new_n17289_), .ZN(new_n17292_));
  NOR2_X1    g16995(.A1(new_n17288_), .A2(new_n17292_), .ZN(new_n17293_));
  OAI22_X1   g16996(.A1(new_n6847_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n7198_), .ZN(new_n17294_));
  OAI21_X1   g16997(.A1(new_n6538_), .A2(new_n2884_), .B(new_n17294_), .ZN(new_n17295_));
  AOI21_X1   g16998(.A1(new_n17295_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n17296_));
  XNOR2_X1   g16999(.A1(new_n7202_), .A2(new_n17296_), .ZN(new_n17297_));
  NOR2_X1    g17000(.A1(new_n17293_), .A2(new_n17297_), .ZN(new_n17298_));
  INV_X1     g17001(.I(new_n17293_), .ZN(new_n17299_));
  INV_X1     g17002(.I(new_n17297_), .ZN(new_n17300_));
  NOR2_X1    g17003(.A1(new_n17299_), .A2(new_n17300_), .ZN(new_n17301_));
  OAI21_X1   g17004(.A1(new_n17301_), .A2(new_n17298_), .B(new_n17142_), .ZN(new_n17302_));
  INV_X1     g17005(.I(new_n17142_), .ZN(new_n17303_));
  NAND2_X1   g17006(.A1(new_n17293_), .A2(new_n17300_), .ZN(new_n17304_));
  INV_X1     g17007(.I(new_n17304_), .ZN(new_n17305_));
  NOR2_X1    g17008(.A1(new_n17293_), .A2(new_n17300_), .ZN(new_n17306_));
  OAI21_X1   g17009(.A1(new_n17305_), .A2(new_n17306_), .B(new_n17303_), .ZN(new_n17307_));
  OAI22_X1   g17010(.A1(new_n2171_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n2166_), .ZN(new_n17308_));
  OAI21_X1   g17011(.A1(new_n7864_), .A2(new_n2322_), .B(new_n17308_), .ZN(new_n17309_));
  AOI21_X1   g17012(.A1(new_n17309_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n17310_));
  XOR2_X1    g17013(.A1(new_n8217_), .A2(new_n17310_), .Z(new_n17311_));
  AOI21_X1   g17014(.A1(new_n17302_), .A2(new_n17307_), .B(new_n17311_), .ZN(new_n17312_));
  INV_X1     g17015(.I(new_n17312_), .ZN(new_n17313_));
  NAND3_X1   g17016(.A1(new_n17302_), .A2(new_n17307_), .A3(new_n17311_), .ZN(new_n17314_));
  AOI21_X1   g17017(.A1(new_n17313_), .A2(new_n17314_), .B(new_n17140_), .ZN(new_n17315_));
  INV_X1     g17018(.I(new_n17311_), .ZN(new_n17316_));
  NAND3_X1   g17019(.A1(new_n17302_), .A2(new_n17307_), .A3(new_n17316_), .ZN(new_n17317_));
  INV_X1     g17020(.I(new_n17302_), .ZN(new_n17318_));
  INV_X1     g17021(.I(new_n17306_), .ZN(new_n17319_));
  AOI21_X1   g17022(.A1(new_n17319_), .A2(new_n17304_), .B(new_n17142_), .ZN(new_n17320_));
  OAI21_X1   g17023(.A1(new_n17318_), .A2(new_n17320_), .B(new_n17311_), .ZN(new_n17321_));
  AOI21_X1   g17024(.A1(new_n17321_), .A2(new_n17317_), .B(new_n17139_), .ZN(new_n17322_));
  OAI22_X1   g17025(.A1(new_n1712_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n1707_), .ZN(new_n17323_));
  OAI21_X1   g17026(.A1(new_n8563_), .A2(new_n1850_), .B(new_n17323_), .ZN(new_n17324_));
  AOI21_X1   g17027(.A1(new_n17324_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n17325_));
  XNOR2_X1   g17028(.A1(new_n9299_), .A2(new_n17325_), .ZN(new_n17326_));
  NOR3_X1    g17029(.A1(new_n17315_), .A2(new_n17322_), .A3(new_n17326_), .ZN(new_n17327_));
  INV_X1     g17030(.I(new_n17314_), .ZN(new_n17328_));
  OAI21_X1   g17031(.A1(new_n17328_), .A2(new_n17312_), .B(new_n17139_), .ZN(new_n17329_));
  INV_X1     g17032(.I(new_n17317_), .ZN(new_n17330_));
  AOI21_X1   g17033(.A1(new_n17302_), .A2(new_n17307_), .B(new_n17316_), .ZN(new_n17331_));
  OAI21_X1   g17034(.A1(new_n17330_), .A2(new_n17331_), .B(new_n17140_), .ZN(new_n17332_));
  INV_X1     g17035(.I(new_n17326_), .ZN(new_n17333_));
  AOI21_X1   g17036(.A1(new_n17329_), .A2(new_n17332_), .B(new_n17333_), .ZN(new_n17334_));
  OAI21_X1   g17037(.A1(new_n17334_), .A2(new_n17327_), .B(new_n17137_), .ZN(new_n17335_));
  OAI21_X1   g17038(.A1(new_n17315_), .A2(new_n17322_), .B(new_n17333_), .ZN(new_n17336_));
  NAND3_X1   g17039(.A1(new_n17329_), .A2(new_n17332_), .A3(new_n17326_), .ZN(new_n17337_));
  AOI21_X1   g17040(.A1(new_n17337_), .A2(new_n17336_), .B(new_n17137_), .ZN(new_n17338_));
  INV_X1     g17041(.I(new_n17338_), .ZN(new_n17339_));
  OAI22_X1   g17042(.A1(new_n1347_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n1344_), .ZN(new_n17340_));
  OAI21_X1   g17043(.A1(new_n10025_), .A2(new_n1457_), .B(new_n17340_), .ZN(new_n17341_));
  AOI21_X1   g17044(.A1(new_n17341_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n17342_));
  XOR2_X1    g17045(.A1(new_n10476_), .A2(new_n17342_), .Z(new_n17343_));
  INV_X1     g17046(.I(new_n17343_), .ZN(new_n17344_));
  NAND3_X1   g17047(.A1(new_n17339_), .A2(new_n17335_), .A3(new_n17344_), .ZN(new_n17345_));
  INV_X1     g17048(.I(new_n17335_), .ZN(new_n17346_));
  OAI21_X1   g17049(.A1(new_n17346_), .A2(new_n17338_), .B(new_n17343_), .ZN(new_n17347_));
  AOI22_X1   g17050(.A1(new_n17347_), .A2(new_n17345_), .B1(new_n17030_), .B2(new_n17136_), .ZN(new_n17348_));
  NAND2_X1   g17051(.A1(new_n17136_), .A2(new_n17030_), .ZN(new_n17349_));
  NAND2_X1   g17052(.A1(new_n17339_), .A2(new_n17335_), .ZN(new_n17350_));
  NAND2_X1   g17053(.A1(new_n17350_), .A2(new_n17344_), .ZN(new_n17351_));
  NAND3_X1   g17054(.A1(new_n17339_), .A2(new_n17335_), .A3(new_n17343_), .ZN(new_n17352_));
  AOI21_X1   g17055(.A1(new_n17351_), .A2(new_n17352_), .B(new_n17349_), .ZN(new_n17353_));
  NOR2_X1    g17056(.A1(new_n17353_), .A2(new_n17348_), .ZN(new_n17354_));
  OAI22_X1   g17057(.A1(new_n1055_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n1061_), .ZN(new_n17355_));
  OAI21_X1   g17058(.A1(new_n10862_), .A2(new_n1332_), .B(new_n17355_), .ZN(new_n17356_));
  AOI21_X1   g17059(.A1(new_n17356_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n17357_));
  XNOR2_X1   g17060(.A1(new_n11748_), .A2(new_n17357_), .ZN(new_n17358_));
  NOR2_X1    g17061(.A1(new_n17354_), .A2(new_n17358_), .ZN(new_n17359_));
  INV_X1     g17062(.I(new_n17354_), .ZN(new_n17360_));
  INV_X1     g17063(.I(new_n17358_), .ZN(new_n17361_));
  NOR2_X1    g17064(.A1(new_n17360_), .A2(new_n17361_), .ZN(new_n17362_));
  OAI22_X1   g17065(.A1(new_n17362_), .A2(new_n17359_), .B1(new_n17041_), .B2(new_n17135_), .ZN(new_n17363_));
  NOR2_X1    g17066(.A1(new_n17135_), .A2(new_n17041_), .ZN(new_n17364_));
  XOR2_X1    g17067(.A1(new_n17354_), .A2(new_n17358_), .Z(new_n17365_));
  NAND2_X1   g17068(.A1(new_n17365_), .A2(new_n17364_), .ZN(new_n17366_));
  NAND2_X1   g17069(.A1(new_n17366_), .A2(new_n17363_), .ZN(new_n17367_));
  OAI22_X1   g17070(.A1(new_n970_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n820_), .ZN(new_n17368_));
  OAI21_X1   g17071(.A1(new_n12536_), .A2(new_n894_), .B(new_n17368_), .ZN(new_n17369_));
  AOI21_X1   g17072(.A1(new_n17369_), .A2(new_n827_), .B(new_n970_), .ZN(new_n17370_));
  XOR2_X1    g17073(.A1(new_n12969_), .A2(new_n17370_), .Z(new_n17371_));
  INV_X1     g17074(.I(new_n17371_), .ZN(new_n17372_));
  XOR2_X1    g17075(.A1(new_n17367_), .A2(new_n17372_), .Z(new_n17373_));
  XOR2_X1    g17076(.A1(new_n17367_), .A2(new_n17371_), .Z(new_n17374_));
  MUX2_X1    g17077(.I0(new_n17374_), .I1(new_n17373_), .S(new_n17133_), .Z(new_n17375_));
  NAND2_X1   g17078(.A1(new_n17069_), .A2(new_n16836_), .ZN(new_n17376_));
  NAND2_X1   g17079(.A1(new_n17376_), .A2(new_n17066_), .ZN(new_n17377_));
  OAI22_X1   g17080(.A1(new_n607_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n610_), .ZN(new_n17378_));
  OAI21_X1   g17081(.A1(new_n13367_), .A2(new_n684_), .B(new_n17378_), .ZN(new_n17379_));
  AOI21_X1   g17082(.A1(new_n17379_), .A2(new_n612_), .B(new_n607_), .ZN(new_n17380_));
  XOR2_X1    g17083(.A1(new_n14213_), .A2(new_n17380_), .Z(new_n17381_));
  XOR2_X1    g17084(.A1(new_n17377_), .A2(new_n17381_), .Z(new_n17382_));
  INV_X1     g17085(.I(new_n17381_), .ZN(new_n17383_));
  NAND2_X1   g17086(.A1(new_n17377_), .A2(new_n17383_), .ZN(new_n17384_));
  NOR2_X1    g17087(.A1(new_n17377_), .A2(new_n17383_), .ZN(new_n17385_));
  INV_X1     g17088(.I(new_n17385_), .ZN(new_n17386_));
  NAND2_X1   g17089(.A1(new_n17386_), .A2(new_n17384_), .ZN(new_n17387_));
  NAND2_X1   g17090(.A1(new_n17375_), .A2(new_n17387_), .ZN(new_n17388_));
  OAI21_X1   g17091(.A1(new_n17375_), .A2(new_n17382_), .B(new_n17388_), .ZN(new_n17389_));
  INV_X1     g17092(.I(new_n17084_), .ZN(new_n17390_));
  OAI21_X1   g17093(.A1(new_n17075_), .A2(new_n17081_), .B(new_n16833_), .ZN(new_n17391_));
  AOI21_X1   g17094(.A1(new_n447_), .A2(new_n749_), .B(new_n16486_), .ZN(new_n17392_));
  INV_X1     g17095(.I(new_n17392_), .ZN(new_n17393_));
  NAND3_X1   g17096(.A1(new_n17391_), .A2(new_n17390_), .A3(new_n17393_), .ZN(new_n17394_));
  NAND2_X1   g17097(.A1(new_n17391_), .A2(new_n17390_), .ZN(new_n17395_));
  NAND2_X1   g17098(.A1(new_n17395_), .A2(new_n17392_), .ZN(new_n17396_));
  AOI21_X1   g17099(.A1(new_n17394_), .A2(new_n17396_), .B(new_n17389_), .ZN(new_n17397_));
  OR2_X2     g17100(.A1(new_n17375_), .A2(new_n17382_), .Z(new_n17398_));
  NAND2_X1   g17101(.A1(new_n17396_), .A2(new_n17394_), .ZN(new_n17399_));
  AOI21_X1   g17102(.A1(new_n17398_), .A2(new_n17388_), .B(new_n17399_), .ZN(new_n17400_));
  OAI21_X1   g17103(.A1(new_n17397_), .A2(new_n17400_), .B(new_n452_), .ZN(new_n17401_));
  INV_X1     g17104(.I(new_n17401_), .ZN(new_n17402_));
  NOR3_X1    g17105(.A1(new_n17397_), .A2(new_n17400_), .A3(new_n452_), .ZN(new_n17403_));
  OAI21_X1   g17106(.A1(new_n17402_), .A2(new_n17403_), .B(new_n17131_), .ZN(new_n17404_));
  NOR2_X1    g17107(.A1(new_n17402_), .A2(new_n17403_), .ZN(new_n17405_));
  NAND2_X1   g17108(.A1(new_n17405_), .A2(new_n17130_), .ZN(new_n17406_));
  NAND2_X1   g17109(.A1(new_n17406_), .A2(new_n17404_), .ZN(new_n17407_));
  NAND2_X1   g17110(.A1(new_n17128_), .A2(new_n17407_), .ZN(new_n17408_));
  INV_X1     g17111(.I(new_n17127_), .ZN(new_n17409_));
  AOI21_X1   g17112(.A1(new_n17114_), .A2(new_n17409_), .B(new_n17125_), .ZN(new_n17410_));
  XOR2_X1    g17113(.A1(new_n17405_), .A2(new_n17130_), .Z(new_n17411_));
  NAND2_X1   g17114(.A1(new_n17410_), .A2(new_n17411_), .ZN(new_n17412_));
  NAND2_X1   g17115(.A1(new_n17408_), .A2(new_n17412_), .ZN(\f[71] ));
  NAND2_X1   g17116(.A1(new_n17389_), .A2(new_n17395_), .ZN(new_n17414_));
  XOR2_X1    g17117(.A1(new_n17392_), .A2(new_n452_), .Z(new_n17415_));
  OAI21_X1   g17118(.A1(new_n17389_), .A2(new_n17395_), .B(new_n17415_), .ZN(new_n17416_));
  NAND2_X1   g17119(.A1(new_n17416_), .A2(new_n17414_), .ZN(new_n17417_));
  INV_X1     g17120(.I(new_n17384_), .ZN(new_n17418_));
  NOR2_X1    g17121(.A1(new_n17375_), .A2(new_n17385_), .ZN(new_n17419_));
  NOR2_X1    g17122(.A1(new_n17419_), .A2(new_n17418_), .ZN(new_n17420_));
  NAND2_X1   g17123(.A1(new_n17367_), .A2(new_n17372_), .ZN(new_n17421_));
  OAI21_X1   g17124(.A1(new_n17367_), .A2(new_n17372_), .B(new_n17133_), .ZN(new_n17422_));
  NAND2_X1   g17125(.A1(new_n17422_), .A2(new_n17421_), .ZN(new_n17423_));
  NOR2_X1    g17126(.A1(new_n17362_), .A2(new_n17364_), .ZN(new_n17424_));
  INV_X1     g17127(.I(new_n17345_), .ZN(new_n17425_));
  AOI22_X1   g17128(.A1(new_n17350_), .A2(new_n17343_), .B1(new_n17030_), .B2(new_n17136_), .ZN(new_n17426_));
  NOR2_X1    g17129(.A1(new_n17426_), .A2(new_n17425_), .ZN(new_n17427_));
  NAND2_X1   g17130(.A1(new_n17337_), .A2(new_n17137_), .ZN(new_n17428_));
  NAND2_X1   g17131(.A1(new_n17428_), .A2(new_n17336_), .ZN(new_n17429_));
  AOI21_X1   g17132(.A1(new_n17139_), .A2(new_n17314_), .B(new_n17312_), .ZN(new_n17430_));
  INV_X1     g17133(.I(new_n17430_), .ZN(new_n17431_));
  XOR2_X1    g17134(.A1(new_n17142_), .A2(new_n17297_), .Z(new_n17432_));
  NOR2_X1    g17135(.A1(new_n17299_), .A2(new_n17432_), .ZN(new_n17433_));
  INV_X1     g17136(.I(new_n17433_), .ZN(new_n17434_));
  NOR2_X1    g17137(.A1(new_n17142_), .A2(new_n17300_), .ZN(new_n17435_));
  INV_X1     g17138(.I(new_n17435_), .ZN(new_n17436_));
  NAND2_X1   g17139(.A1(new_n17287_), .A2(new_n17289_), .ZN(new_n17437_));
  NAND2_X1   g17140(.A1(new_n17437_), .A2(new_n17286_), .ZN(new_n17438_));
  NAND2_X1   g17141(.A1(new_n17268_), .A2(new_n17272_), .ZN(new_n17439_));
  XOR2_X1    g17142(.A1(new_n17276_), .A2(new_n4069_), .Z(new_n17440_));
  OAI21_X1   g17143(.A1(new_n17268_), .A2(new_n17272_), .B(new_n17440_), .ZN(new_n17441_));
  NAND2_X1   g17144(.A1(new_n17441_), .A2(new_n17439_), .ZN(new_n17442_));
  NAND2_X1   g17145(.A1(new_n17264_), .A2(new_n17147_), .ZN(new_n17443_));
  NAND2_X1   g17146(.A1(new_n17443_), .A2(new_n17263_), .ZN(new_n17444_));
  OAI21_X1   g17147(.A1(new_n17152_), .A2(new_n17256_), .B(new_n17254_), .ZN(new_n17445_));
  OAI21_X1   g17148(.A1(new_n17244_), .A2(new_n17242_), .B(new_n17240_), .ZN(new_n17446_));
  NOR2_X1    g17149(.A1(new_n17229_), .A2(new_n17155_), .ZN(new_n17447_));
  NAND2_X1   g17150(.A1(new_n17226_), .A2(new_n17223_), .ZN(new_n17448_));
  NAND2_X1   g17151(.A1(new_n17448_), .A2(new_n17225_), .ZN(new_n17449_));
  OAI22_X1   g17152(.A1(new_n8644_), .A2(new_n1936_), .B1(new_n2102_), .B2(new_n9388_), .ZN(new_n17450_));
  OAI21_X1   g17153(.A1(new_n1803_), .A2(new_n10154_), .B(new_n17450_), .ZN(new_n17451_));
  AOI21_X1   g17154(.A1(new_n17451_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n17452_));
  XOR2_X1    g17155(.A1(new_n2106_), .A2(new_n17452_), .Z(new_n17453_));
  INV_X1     g17156(.I(new_n17453_), .ZN(new_n17454_));
  NAND2_X1   g17157(.A1(new_n17216_), .A2(new_n17214_), .ZN(new_n17455_));
  NAND2_X1   g17158(.A1(new_n17195_), .A2(new_n17184_), .ZN(new_n17456_));
  NAND2_X1   g17159(.A1(new_n17456_), .A2(new_n17194_), .ZN(new_n17457_));
  INV_X1     g17160(.I(new_n17176_), .ZN(new_n17458_));
  AOI21_X1   g17161(.A1(new_n17171_), .A2(new_n17458_), .B(new_n17178_), .ZN(new_n17459_));
  OAI22_X1   g17162(.A1(new_n13880_), .A2(new_n781_), .B1(new_n656_), .B2(new_n13885_), .ZN(new_n17460_));
  AOI21_X1   g17163(.A1(new_n17460_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n17461_));
  XOR2_X1    g17164(.A1(new_n785_), .A2(new_n17461_), .Z(new_n17462_));
  NOR2_X1    g17165(.A1(new_n13476_), .A2(new_n515_), .ZN(new_n17463_));
  XOR2_X1    g17166(.A1(new_n14736_), .A2(new_n515_), .Z(new_n17464_));
  NAND2_X1   g17167(.A1(new_n17464_), .A2(\b[9] ), .ZN(new_n17465_));
  XOR2_X1    g17168(.A1(new_n17465_), .A2(new_n17463_), .Z(new_n17466_));
  XOR2_X1    g17169(.A1(new_n17466_), .A2(\a[8] ), .Z(new_n17467_));
  NOR2_X1    g17170(.A1(new_n17467_), .A2(new_n17175_), .ZN(new_n17468_));
  NOR2_X1    g17171(.A1(new_n17466_), .A2(new_n452_), .ZN(new_n17469_));
  INV_X1     g17172(.I(new_n17469_), .ZN(new_n17470_));
  NAND2_X1   g17173(.A1(new_n17466_), .A2(new_n452_), .ZN(new_n17471_));
  AOI21_X1   g17174(.A1(new_n17470_), .A2(new_n17471_), .B(new_n17177_), .ZN(new_n17472_));
  OAI21_X1   g17175(.A1(new_n17468_), .A2(new_n17472_), .B(new_n17462_), .ZN(new_n17473_));
  INV_X1     g17176(.I(new_n17462_), .ZN(new_n17474_));
  NOR2_X1    g17177(.A1(new_n17468_), .A2(new_n17472_), .ZN(new_n17475_));
  NAND2_X1   g17178(.A1(new_n17474_), .A2(new_n17475_), .ZN(new_n17476_));
  AOI21_X1   g17179(.A1(new_n17476_), .A2(new_n17473_), .B(new_n17459_), .ZN(new_n17477_));
  INV_X1     g17180(.I(new_n17459_), .ZN(new_n17478_));
  XOR2_X1    g17181(.A1(new_n17462_), .A2(new_n17475_), .Z(new_n17479_));
  NOR2_X1    g17182(.A1(new_n17479_), .A2(new_n17478_), .ZN(new_n17480_));
  NOR2_X1    g17183(.A1(new_n17480_), .A2(new_n17477_), .ZN(new_n17481_));
  AOI22_X1   g17184(.A1(new_n13078_), .A2(\b[13] ), .B1(new_n1105_), .B2(new_n12218_), .ZN(new_n17482_));
  OAI21_X1   g17185(.A1(new_n17482_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n17483_));
  XOR2_X1    g17186(.A1(new_n1024_), .A2(new_n17483_), .Z(new_n17484_));
  INV_X1     g17187(.I(new_n17484_), .ZN(new_n17485_));
  XOR2_X1    g17188(.A1(new_n17481_), .A2(new_n17485_), .Z(new_n17486_));
  OAI21_X1   g17189(.A1(new_n17480_), .A2(new_n17477_), .B(new_n17484_), .ZN(new_n17487_));
  NAND2_X1   g17190(.A1(new_n17481_), .A2(new_n17485_), .ZN(new_n17488_));
  AOI21_X1   g17191(.A1(new_n17487_), .A2(new_n17488_), .B(new_n17457_), .ZN(new_n17489_));
  AOI21_X1   g17192(.A1(new_n17486_), .A2(new_n17457_), .B(new_n17489_), .ZN(new_n17490_));
  INV_X1     g17193(.I(new_n17490_), .ZN(new_n17491_));
  AOI22_X1   g17194(.A1(new_n10969_), .A2(new_n1296_), .B1(new_n11394_), .B2(\b[16] ), .ZN(new_n17492_));
  OAI21_X1   g17195(.A1(new_n17492_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n17493_));
  XNOR2_X1   g17196(.A1(new_n1299_), .A2(new_n17493_), .ZN(new_n17494_));
  NAND2_X1   g17197(.A1(new_n17197_), .A2(new_n17205_), .ZN(new_n17495_));
  AOI21_X1   g17198(.A1(new_n17495_), .A2(new_n17204_), .B(new_n17494_), .ZN(new_n17496_));
  INV_X1     g17199(.I(new_n17494_), .ZN(new_n17497_));
  NAND2_X1   g17200(.A1(new_n17495_), .A2(new_n17204_), .ZN(new_n17498_));
  NOR2_X1    g17201(.A1(new_n17498_), .A2(new_n17497_), .ZN(new_n17499_));
  OAI21_X1   g17202(.A1(new_n17496_), .A2(new_n17499_), .B(new_n17491_), .ZN(new_n17500_));
  XOR2_X1    g17203(.A1(new_n17498_), .A2(new_n17497_), .Z(new_n17501_));
  NAND2_X1   g17204(.A1(new_n17501_), .A2(new_n17490_), .ZN(new_n17502_));
  NAND2_X1   g17205(.A1(new_n17502_), .A2(new_n17500_), .ZN(new_n17503_));
  AOI22_X1   g17206(.A1(new_n11415_), .A2(new_n1797_), .B1(\b[19] ), .B2(new_n10145_), .ZN(new_n17504_));
  OAI21_X1   g17207(.A1(new_n17504_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n17505_));
  XOR2_X1    g17208(.A1(new_n1638_), .A2(new_n17505_), .Z(new_n17506_));
  INV_X1     g17209(.I(new_n17506_), .ZN(new_n17507_));
  NAND2_X1   g17210(.A1(new_n17503_), .A2(new_n17507_), .ZN(new_n17508_));
  INV_X1     g17211(.I(new_n17503_), .ZN(new_n17509_));
  NAND2_X1   g17212(.A1(new_n17509_), .A2(new_n17506_), .ZN(new_n17510_));
  AOI22_X1   g17213(.A1(new_n17510_), .A2(new_n17508_), .B1(new_n17215_), .B2(new_n17455_), .ZN(new_n17511_));
  NAND2_X1   g17214(.A1(new_n17455_), .A2(new_n17215_), .ZN(new_n17512_));
  NAND2_X1   g17215(.A1(new_n17509_), .A2(new_n17507_), .ZN(new_n17513_));
  NAND2_X1   g17216(.A1(new_n17503_), .A2(new_n17506_), .ZN(new_n17514_));
  AOI21_X1   g17217(.A1(new_n17513_), .A2(new_n17514_), .B(new_n17512_), .ZN(new_n17515_));
  NOR2_X1    g17218(.A1(new_n17511_), .A2(new_n17515_), .ZN(new_n17516_));
  NOR2_X1    g17219(.A1(new_n17516_), .A2(new_n17454_), .ZN(new_n17517_));
  INV_X1     g17220(.I(new_n17516_), .ZN(new_n17518_));
  NOR2_X1    g17221(.A1(new_n17518_), .A2(new_n17453_), .ZN(new_n17519_));
  OAI21_X1   g17222(.A1(new_n17519_), .A2(new_n17517_), .B(new_n17449_), .ZN(new_n17520_));
  XOR2_X1    g17223(.A1(new_n17516_), .A2(new_n17454_), .Z(new_n17521_));
  NAND3_X1   g17224(.A1(new_n17521_), .A2(new_n17225_), .A3(new_n17448_), .ZN(new_n17522_));
  NAND2_X1   g17225(.A1(new_n17522_), .A2(new_n17520_), .ZN(new_n17523_));
  OAI22_X1   g17226(.A1(new_n7619_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n8309_), .ZN(new_n17524_));
  OAI21_X1   g17227(.A1(new_n2281_), .A2(new_n7947_), .B(new_n17524_), .ZN(new_n17525_));
  AOI21_X1   g17228(.A1(new_n17525_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n17526_));
  XNOR2_X1   g17229(.A1(new_n2647_), .A2(new_n17526_), .ZN(new_n17527_));
  INV_X1     g17230(.I(new_n17527_), .ZN(new_n17528_));
  XOR2_X1    g17231(.A1(new_n17523_), .A2(new_n17528_), .Z(new_n17529_));
  OAI21_X1   g17232(.A1(new_n17231_), .A2(new_n17447_), .B(new_n17529_), .ZN(new_n17530_));
  NOR2_X1    g17233(.A1(new_n17447_), .A2(new_n17231_), .ZN(new_n17531_));
  AOI21_X1   g17234(.A1(new_n17522_), .A2(new_n17520_), .B(new_n17527_), .ZN(new_n17532_));
  NOR2_X1    g17235(.A1(new_n17523_), .A2(new_n17528_), .ZN(new_n17533_));
  OAI21_X1   g17236(.A1(new_n17533_), .A2(new_n17532_), .B(new_n17531_), .ZN(new_n17534_));
  NAND2_X1   g17237(.A1(new_n17530_), .A2(new_n17534_), .ZN(new_n17535_));
  OAI22_X1   g17238(.A1(new_n6644_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n6647_), .ZN(new_n17536_));
  OAI21_X1   g17239(.A1(new_n2842_), .A2(new_n7284_), .B(new_n17536_), .ZN(new_n17537_));
  AOI21_X1   g17240(.A1(new_n17537_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n17538_));
  XNOR2_X1   g17241(.A1(new_n3264_), .A2(new_n17538_), .ZN(new_n17539_));
  NOR2_X1    g17242(.A1(new_n17535_), .A2(new_n17539_), .ZN(new_n17540_));
  AND2_X2    g17243(.A1(new_n17535_), .A2(new_n17539_), .Z(new_n17541_));
  OAI21_X1   g17244(.A1(new_n17541_), .A2(new_n17540_), .B(new_n17446_), .ZN(new_n17542_));
  INV_X1     g17245(.I(new_n17446_), .ZN(new_n17543_));
  XOR2_X1    g17246(.A1(new_n17535_), .A2(new_n17539_), .Z(new_n17544_));
  NAND2_X1   g17247(.A1(new_n17544_), .A2(new_n17543_), .ZN(new_n17545_));
  NAND2_X1   g17248(.A1(new_n17545_), .A2(new_n17542_), .ZN(new_n17546_));
  OAI22_X1   g17249(.A1(new_n5993_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n5991_), .ZN(new_n17547_));
  OAI21_X1   g17250(.A1(new_n3709_), .A2(new_n5997_), .B(new_n17547_), .ZN(new_n17548_));
  AOI21_X1   g17251(.A1(new_n17548_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n17549_));
  XNOR2_X1   g17252(.A1(new_n3993_), .A2(new_n17549_), .ZN(new_n17550_));
  INV_X1     g17253(.I(new_n17550_), .ZN(new_n17551_));
  NAND2_X1   g17254(.A1(new_n17546_), .A2(new_n17551_), .ZN(new_n17552_));
  INV_X1     g17255(.I(new_n17552_), .ZN(new_n17553_));
  NOR2_X1    g17256(.A1(new_n17546_), .A2(new_n17551_), .ZN(new_n17554_));
  OAI21_X1   g17257(.A1(new_n17553_), .A2(new_n17554_), .B(new_n17445_), .ZN(new_n17555_));
  INV_X1     g17258(.I(new_n17445_), .ZN(new_n17556_));
  XOR2_X1    g17259(.A1(new_n17546_), .A2(new_n17551_), .Z(new_n17557_));
  NAND2_X1   g17260(.A1(new_n17557_), .A2(new_n17556_), .ZN(new_n17558_));
  NAND2_X1   g17261(.A1(new_n17558_), .A2(new_n17555_), .ZN(new_n17559_));
  OAI22_X1   g17262(.A1(new_n5420_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n5107_), .ZN(new_n17560_));
  OAI21_X1   g17263(.A1(new_n4253_), .A2(new_n5112_), .B(new_n17560_), .ZN(new_n17561_));
  AOI21_X1   g17264(.A1(new_n17561_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n17562_));
  XNOR2_X1   g17265(.A1(new_n4778_), .A2(new_n17562_), .ZN(new_n17563_));
  INV_X1     g17266(.I(new_n17563_), .ZN(new_n17564_));
  XOR2_X1    g17267(.A1(new_n17559_), .A2(new_n17564_), .Z(new_n17565_));
  NAND2_X1   g17268(.A1(new_n17565_), .A2(new_n17444_), .ZN(new_n17566_));
  INV_X1     g17269(.I(new_n17444_), .ZN(new_n17567_));
  NAND2_X1   g17270(.A1(new_n17559_), .A2(new_n17564_), .ZN(new_n17568_));
  INV_X1     g17271(.I(new_n17568_), .ZN(new_n17569_));
  NOR2_X1    g17272(.A1(new_n17559_), .A2(new_n17564_), .ZN(new_n17570_));
  OAI21_X1   g17273(.A1(new_n17569_), .A2(new_n17570_), .B(new_n17567_), .ZN(new_n17571_));
  NAND2_X1   g17274(.A1(new_n17566_), .A2(new_n17571_), .ZN(new_n17572_));
  OAI22_X1   g17275(.A1(new_n4072_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n4067_), .ZN(new_n17573_));
  OAI21_X1   g17276(.A1(new_n5068_), .A2(new_n4318_), .B(new_n17573_), .ZN(new_n17574_));
  AOI21_X1   g17277(.A1(new_n17574_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n17575_));
  XNOR2_X1   g17278(.A1(new_n5600_), .A2(new_n17575_), .ZN(new_n17576_));
  NOR2_X1    g17279(.A1(new_n17572_), .A2(new_n17576_), .ZN(new_n17577_));
  AND2_X2    g17280(.A1(new_n17572_), .A2(new_n17576_), .Z(new_n17578_));
  OAI21_X1   g17281(.A1(new_n17578_), .A2(new_n17577_), .B(new_n17442_), .ZN(new_n17579_));
  INV_X1     g17282(.I(new_n17442_), .ZN(new_n17580_));
  XOR2_X1    g17283(.A1(new_n17572_), .A2(new_n17576_), .Z(new_n17581_));
  NAND2_X1   g17284(.A1(new_n17581_), .A2(new_n17580_), .ZN(new_n17582_));
  NAND2_X1   g17285(.A1(new_n17582_), .A2(new_n17579_), .ZN(new_n17583_));
  OAI22_X1   g17286(.A1(new_n6229_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n6538_), .ZN(new_n17584_));
  OAI21_X1   g17287(.A1(new_n5921_), .A2(new_n3569_), .B(new_n17584_), .ZN(new_n17585_));
  AOI21_X1   g17288(.A1(new_n17585_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n17586_));
  XOR2_X1    g17289(.A1(new_n6543_), .A2(new_n17586_), .Z(new_n17587_));
  INV_X1     g17290(.I(new_n17587_), .ZN(new_n17588_));
  NAND2_X1   g17291(.A1(new_n17583_), .A2(new_n17588_), .ZN(new_n17589_));
  INV_X1     g17292(.I(new_n17589_), .ZN(new_n17590_));
  NOR2_X1    g17293(.A1(new_n17583_), .A2(new_n17588_), .ZN(new_n17591_));
  OAI21_X1   g17294(.A1(new_n17590_), .A2(new_n17591_), .B(new_n17438_), .ZN(new_n17592_));
  INV_X1     g17295(.I(new_n17438_), .ZN(new_n17593_));
  XOR2_X1    g17296(.A1(new_n17583_), .A2(new_n17588_), .Z(new_n17594_));
  NAND2_X1   g17297(.A1(new_n17594_), .A2(new_n17593_), .ZN(new_n17595_));
  NAND2_X1   g17298(.A1(new_n17595_), .A2(new_n17592_), .ZN(new_n17596_));
  OAI22_X1   g17299(.A1(new_n7864_), .A2(new_n2700_), .B1(new_n2705_), .B2(new_n7198_), .ZN(new_n17597_));
  OAI21_X1   g17300(.A1(new_n6847_), .A2(new_n2884_), .B(new_n17597_), .ZN(new_n17598_));
  AOI21_X1   g17301(.A1(new_n17598_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n17599_));
  XNOR2_X1   g17302(.A1(new_n7516_), .A2(new_n17599_), .ZN(new_n17600_));
  NAND3_X1   g17303(.A1(new_n17596_), .A2(new_n17436_), .A3(new_n17600_), .ZN(new_n17601_));
  INV_X1     g17304(.I(new_n17601_), .ZN(new_n17602_));
  AOI21_X1   g17305(.A1(new_n17596_), .A2(new_n17600_), .B(new_n17436_), .ZN(new_n17603_));
  OAI21_X1   g17306(.A1(new_n17602_), .A2(new_n17603_), .B(new_n17434_), .ZN(new_n17604_));
  INV_X1     g17307(.I(new_n17603_), .ZN(new_n17605_));
  NAND3_X1   g17308(.A1(new_n17605_), .A2(new_n17433_), .A3(new_n17601_), .ZN(new_n17606_));
  OAI22_X1   g17309(.A1(new_n2171_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n2166_), .ZN(new_n17607_));
  OAI21_X1   g17310(.A1(new_n7870_), .A2(new_n2322_), .B(new_n17607_), .ZN(new_n17608_));
  AOI21_X1   g17311(.A1(new_n17608_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n17609_));
  XOR2_X1    g17312(.A1(new_n8568_), .A2(new_n17609_), .Z(new_n17610_));
  AOI21_X1   g17313(.A1(new_n17606_), .A2(new_n17604_), .B(new_n17610_), .ZN(new_n17611_));
  NAND3_X1   g17314(.A1(new_n17606_), .A2(new_n17604_), .A3(new_n17610_), .ZN(new_n17612_));
  INV_X1     g17315(.I(new_n17612_), .ZN(new_n17613_));
  OAI21_X1   g17316(.A1(new_n17613_), .A2(new_n17611_), .B(new_n17431_), .ZN(new_n17614_));
  INV_X1     g17317(.I(new_n17610_), .ZN(new_n17615_));
  NAND3_X1   g17318(.A1(new_n17606_), .A2(new_n17604_), .A3(new_n17615_), .ZN(new_n17616_));
  INV_X1     g17319(.I(new_n17616_), .ZN(new_n17617_));
  AOI21_X1   g17320(.A1(new_n17606_), .A2(new_n17604_), .B(new_n17615_), .ZN(new_n17618_));
  OAI21_X1   g17321(.A1(new_n17617_), .A2(new_n17618_), .B(new_n17430_), .ZN(new_n17619_));
  OAI22_X1   g17322(.A1(new_n1712_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n1707_), .ZN(new_n17620_));
  OAI21_X1   g17323(.A1(new_n8948_), .A2(new_n1850_), .B(new_n17620_), .ZN(new_n17621_));
  AOI21_X1   g17324(.A1(new_n17621_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n17622_));
  XNOR2_X1   g17325(.A1(new_n9642_), .A2(new_n17622_), .ZN(new_n17623_));
  AOI21_X1   g17326(.A1(new_n17614_), .A2(new_n17619_), .B(new_n17623_), .ZN(new_n17624_));
  INV_X1     g17327(.I(new_n17611_), .ZN(new_n17625_));
  AOI21_X1   g17328(.A1(new_n17625_), .A2(new_n17612_), .B(new_n17430_), .ZN(new_n17626_));
  INV_X1     g17329(.I(new_n17618_), .ZN(new_n17627_));
  AOI21_X1   g17330(.A1(new_n17627_), .A2(new_n17616_), .B(new_n17431_), .ZN(new_n17628_));
  INV_X1     g17331(.I(new_n17623_), .ZN(new_n17629_));
  NOR3_X1    g17332(.A1(new_n17626_), .A2(new_n17628_), .A3(new_n17629_), .ZN(new_n17630_));
  OAI21_X1   g17333(.A1(new_n17630_), .A2(new_n17624_), .B(new_n17429_), .ZN(new_n17631_));
  INV_X1     g17334(.I(new_n17429_), .ZN(new_n17632_));
  NOR3_X1    g17335(.A1(new_n17626_), .A2(new_n17628_), .A3(new_n17623_), .ZN(new_n17633_));
  AOI21_X1   g17336(.A1(new_n17614_), .A2(new_n17619_), .B(new_n17629_), .ZN(new_n17634_));
  OAI21_X1   g17337(.A1(new_n17633_), .A2(new_n17634_), .B(new_n17632_), .ZN(new_n17635_));
  OAI22_X1   g17338(.A1(new_n1347_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n1344_), .ZN(new_n17636_));
  OAI21_X1   g17339(.A1(new_n10031_), .A2(new_n1457_), .B(new_n17636_), .ZN(new_n17637_));
  AOI21_X1   g17340(.A1(new_n17637_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n17638_));
  XNOR2_X1   g17341(.A1(new_n10866_), .A2(new_n17638_), .ZN(new_n17639_));
  AOI21_X1   g17342(.A1(new_n17631_), .A2(new_n17635_), .B(new_n17639_), .ZN(new_n17640_));
  INV_X1     g17343(.I(new_n17640_), .ZN(new_n17641_));
  NAND3_X1   g17344(.A1(new_n17631_), .A2(new_n17635_), .A3(new_n17639_), .ZN(new_n17642_));
  AOI21_X1   g17345(.A1(new_n17641_), .A2(new_n17642_), .B(new_n17427_), .ZN(new_n17643_));
  OAI21_X1   g17346(.A1(new_n17626_), .A2(new_n17628_), .B(new_n17629_), .ZN(new_n17644_));
  NAND3_X1   g17347(.A1(new_n17614_), .A2(new_n17619_), .A3(new_n17623_), .ZN(new_n17645_));
  AOI21_X1   g17348(.A1(new_n17644_), .A2(new_n17645_), .B(new_n17632_), .ZN(new_n17646_));
  NAND3_X1   g17349(.A1(new_n17614_), .A2(new_n17619_), .A3(new_n17629_), .ZN(new_n17647_));
  OAI21_X1   g17350(.A1(new_n17626_), .A2(new_n17628_), .B(new_n17623_), .ZN(new_n17648_));
  AOI21_X1   g17351(.A1(new_n17648_), .A2(new_n17647_), .B(new_n17429_), .ZN(new_n17649_));
  NOR3_X1    g17352(.A1(new_n17646_), .A2(new_n17649_), .A3(new_n17639_), .ZN(new_n17650_));
  INV_X1     g17353(.I(new_n17639_), .ZN(new_n17651_));
  AOI21_X1   g17354(.A1(new_n17631_), .A2(new_n17635_), .B(new_n17651_), .ZN(new_n17652_));
  OAI21_X1   g17355(.A1(new_n17652_), .A2(new_n17650_), .B(new_n17427_), .ZN(new_n17653_));
  INV_X1     g17356(.I(new_n17653_), .ZN(new_n17654_));
  OAI22_X1   g17357(.A1(new_n1055_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n1061_), .ZN(new_n17655_));
  OAI21_X1   g17358(.A1(new_n11738_), .A2(new_n1332_), .B(new_n17655_), .ZN(new_n17656_));
  AOI21_X1   g17359(.A1(new_n17656_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n17657_));
  XNOR2_X1   g17360(.A1(new_n12128_), .A2(new_n17657_), .ZN(new_n17658_));
  NOR3_X1    g17361(.A1(new_n17654_), .A2(new_n17643_), .A3(new_n17658_), .ZN(new_n17659_));
  INV_X1     g17362(.I(new_n17427_), .ZN(new_n17660_));
  NOR3_X1    g17363(.A1(new_n17646_), .A2(new_n17649_), .A3(new_n17651_), .ZN(new_n17661_));
  OAI21_X1   g17364(.A1(new_n17640_), .A2(new_n17661_), .B(new_n17660_), .ZN(new_n17662_));
  INV_X1     g17365(.I(new_n17658_), .ZN(new_n17663_));
  AOI21_X1   g17366(.A1(new_n17662_), .A2(new_n17653_), .B(new_n17663_), .ZN(new_n17664_));
  OAI22_X1   g17367(.A1(new_n17424_), .A2(new_n17359_), .B1(new_n17659_), .B2(new_n17664_), .ZN(new_n17665_));
  NOR2_X1    g17368(.A1(new_n17424_), .A2(new_n17359_), .ZN(new_n17666_));
  OAI21_X1   g17369(.A1(new_n17654_), .A2(new_n17643_), .B(new_n17663_), .ZN(new_n17667_));
  NAND3_X1   g17370(.A1(new_n17662_), .A2(new_n17653_), .A3(new_n17658_), .ZN(new_n17668_));
  NAND2_X1   g17371(.A1(new_n17667_), .A2(new_n17668_), .ZN(new_n17669_));
  NAND2_X1   g17372(.A1(new_n17669_), .A2(new_n17666_), .ZN(new_n17670_));
  OAI22_X1   g17373(.A1(new_n970_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n820_), .ZN(new_n17671_));
  OAI21_X1   g17374(.A1(new_n12542_), .A2(new_n894_), .B(new_n17671_), .ZN(new_n17672_));
  AOI21_X1   g17375(.A1(new_n17672_), .A2(new_n827_), .B(new_n970_), .ZN(new_n17673_));
  XNOR2_X1   g17376(.A1(new_n13371_), .A2(new_n17673_), .ZN(new_n17674_));
  INV_X1     g17377(.I(new_n17674_), .ZN(new_n17675_));
  NAND3_X1   g17378(.A1(new_n17670_), .A2(new_n17665_), .A3(new_n17675_), .ZN(new_n17676_));
  NAND2_X1   g17379(.A1(new_n17670_), .A2(new_n17665_), .ZN(new_n17677_));
  NAND2_X1   g17380(.A1(new_n17677_), .A2(new_n17674_), .ZN(new_n17678_));
  NAND2_X1   g17381(.A1(new_n17678_), .A2(new_n17676_), .ZN(new_n17679_));
  NAND2_X1   g17382(.A1(new_n17679_), .A2(new_n17423_), .ZN(new_n17680_));
  INV_X1     g17383(.I(new_n17423_), .ZN(new_n17681_));
  AOI21_X1   g17384(.A1(new_n17670_), .A2(new_n17665_), .B(new_n17674_), .ZN(new_n17682_));
  NOR2_X1    g17385(.A1(new_n17677_), .A2(new_n17675_), .ZN(new_n17683_));
  OAI21_X1   g17386(.A1(new_n17682_), .A2(new_n17683_), .B(new_n17681_), .ZN(new_n17684_));
  OAI22_X1   g17387(.A1(new_n607_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n610_), .ZN(new_n17685_));
  OAI21_X1   g17388(.A1(new_n13785_), .A2(new_n684_), .B(new_n17685_), .ZN(new_n17686_));
  AOI21_X1   g17389(.A1(new_n17686_), .A2(new_n612_), .B(new_n607_), .ZN(new_n17687_));
  XNOR2_X1   g17390(.A1(new_n14599_), .A2(new_n17687_), .ZN(new_n17688_));
  AOI21_X1   g17391(.A1(new_n17684_), .A2(new_n17680_), .B(new_n17688_), .ZN(new_n17689_));
  AOI21_X1   g17392(.A1(new_n17676_), .A2(new_n17678_), .B(new_n17681_), .ZN(new_n17690_));
  NOR2_X1    g17393(.A1(new_n17683_), .A2(new_n17682_), .ZN(new_n17691_));
  NOR2_X1    g17394(.A1(new_n17691_), .A2(new_n17423_), .ZN(new_n17692_));
  INV_X1     g17395(.I(new_n17688_), .ZN(new_n17693_));
  NOR3_X1    g17396(.A1(new_n17692_), .A2(new_n17690_), .A3(new_n17693_), .ZN(new_n17694_));
  NOR2_X1    g17397(.A1(new_n17689_), .A2(new_n17694_), .ZN(new_n17695_));
  NOR3_X1    g17398(.A1(new_n17692_), .A2(new_n17690_), .A3(new_n17688_), .ZN(new_n17696_));
  AOI21_X1   g17399(.A1(new_n17684_), .A2(new_n17680_), .B(new_n17693_), .ZN(new_n17697_));
  OAI21_X1   g17400(.A1(new_n17696_), .A2(new_n17697_), .B(new_n17420_), .ZN(new_n17698_));
  OAI21_X1   g17401(.A1(new_n17420_), .A2(new_n17695_), .B(new_n17698_), .ZN(new_n17699_));
  NAND2_X1   g17402(.A1(new_n17699_), .A2(new_n17417_), .ZN(new_n17700_));
  INV_X1     g17403(.I(new_n17420_), .ZN(new_n17701_));
  OAI21_X1   g17404(.A1(new_n17689_), .A2(new_n17694_), .B(new_n17701_), .ZN(new_n17702_));
  NAND4_X1   g17405(.A1(new_n17702_), .A2(new_n17416_), .A3(new_n17414_), .A4(new_n17698_), .ZN(new_n17703_));
  NAND2_X1   g17406(.A1(new_n17700_), .A2(new_n17703_), .ZN(new_n17704_));
  NAND2_X1   g17407(.A1(new_n17411_), .A2(new_n17704_), .ZN(new_n17705_));
  XOR2_X1    g17408(.A1(new_n17705_), .A2(new_n17404_), .Z(new_n17706_));
  XOR2_X1    g17409(.A1(new_n17706_), .A2(new_n17128_), .Z(\f[72] ));
  INV_X1     g17410(.I(new_n17703_), .ZN(new_n17708_));
  NAND3_X1   g17411(.A1(new_n17405_), .A2(new_n17700_), .A3(new_n17703_), .ZN(new_n17709_));
  INV_X1     g17412(.I(new_n17403_), .ZN(new_n17710_));
  AOI22_X1   g17413(.A1(new_n17710_), .A2(new_n17401_), .B1(new_n17700_), .B2(new_n17703_), .ZN(new_n17711_));
  OAI21_X1   g17414(.A1(new_n17711_), .A2(new_n17131_), .B(new_n17709_), .ZN(new_n17712_));
  NOR2_X1    g17415(.A1(new_n17410_), .A2(new_n17712_), .ZN(new_n17713_));
  NOR2_X1    g17416(.A1(new_n17420_), .A2(new_n17694_), .ZN(new_n17714_));
  NOR2_X1    g17417(.A1(new_n17714_), .A2(new_n17689_), .ZN(new_n17715_));
  NAND2_X1   g17418(.A1(new_n17678_), .A2(new_n17423_), .ZN(new_n17716_));
  NAND2_X1   g17419(.A1(new_n17716_), .A2(new_n17676_), .ZN(new_n17717_));
  INV_X1     g17420(.I(new_n17717_), .ZN(new_n17718_));
  OAI21_X1   g17421(.A1(new_n17424_), .A2(new_n17359_), .B(new_n17668_), .ZN(new_n17719_));
  NAND2_X1   g17422(.A1(new_n17719_), .A2(new_n17667_), .ZN(new_n17720_));
  INV_X1     g17423(.I(new_n17720_), .ZN(new_n17721_));
  AOI21_X1   g17424(.A1(new_n17660_), .A2(new_n17642_), .B(new_n17640_), .ZN(new_n17722_));
  AOI21_X1   g17425(.A1(new_n17429_), .A2(new_n17645_), .B(new_n17624_), .ZN(new_n17723_));
  NAND2_X1   g17426(.A1(new_n17596_), .A2(new_n17433_), .ZN(new_n17724_));
  NAND3_X1   g17427(.A1(new_n17434_), .A2(new_n17592_), .A3(new_n17595_), .ZN(new_n17725_));
  NAND3_X1   g17428(.A1(new_n17725_), .A2(new_n17435_), .A3(new_n17600_), .ZN(new_n17726_));
  NAND2_X1   g17429(.A1(new_n17726_), .A2(new_n17724_), .ZN(new_n17727_));
  INV_X1     g17430(.I(new_n17577_), .ZN(new_n17728_));
  OAI21_X1   g17431(.A1(new_n17580_), .A2(new_n17578_), .B(new_n17728_), .ZN(new_n17729_));
  OAI21_X1   g17432(.A1(new_n17567_), .A2(new_n17570_), .B(new_n17568_), .ZN(new_n17730_));
  INV_X1     g17433(.I(new_n17730_), .ZN(new_n17731_));
  OAI21_X1   g17434(.A1(new_n17556_), .A2(new_n17554_), .B(new_n17552_), .ZN(new_n17732_));
  INV_X1     g17435(.I(new_n17732_), .ZN(new_n17733_));
  NOR2_X1    g17436(.A1(new_n17541_), .A2(new_n17543_), .ZN(new_n17734_));
  NOR2_X1    g17437(.A1(new_n17734_), .A2(new_n17540_), .ZN(new_n17735_));
  OAI22_X1   g17438(.A1(new_n5993_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n5991_), .ZN(new_n17736_));
  OAI21_X1   g17439(.A1(new_n3717_), .A2(new_n5997_), .B(new_n17736_), .ZN(new_n17737_));
  AOI21_X1   g17440(.A1(new_n17737_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n17738_));
  INV_X1     g17441(.I(new_n17738_), .ZN(new_n17739_));
  NOR2_X1    g17442(.A1(new_n4257_), .A2(new_n17739_), .ZN(new_n17740_));
  NOR2_X1    g17443(.A1(new_n16962_), .A2(new_n17738_), .ZN(new_n17741_));
  NOR2_X1    g17444(.A1(new_n17741_), .A2(new_n17740_), .ZN(new_n17742_));
  OAI22_X1   g17445(.A1(new_n7619_), .A2(new_n2643_), .B1(new_n2842_), .B2(new_n8309_), .ZN(new_n17743_));
  OAI21_X1   g17446(.A1(new_n2439_), .A2(new_n7947_), .B(new_n17743_), .ZN(new_n17744_));
  AOI21_X1   g17447(.A1(new_n17744_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n17745_));
  XNOR2_X1   g17448(.A1(new_n2846_), .A2(new_n17745_), .ZN(new_n17746_));
  AOI22_X1   g17449(.A1(new_n11415_), .A2(new_n1805_), .B1(\b[20] ), .B2(new_n10145_), .ZN(new_n17747_));
  OAI21_X1   g17450(.A1(new_n17747_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n17748_));
  XNOR2_X1   g17451(.A1(new_n1808_), .A2(new_n17748_), .ZN(new_n17749_));
  INV_X1     g17452(.I(new_n17749_), .ZN(new_n17750_));
  NAND2_X1   g17453(.A1(new_n17478_), .A2(new_n17473_), .ZN(new_n17751_));
  AND2_X2    g17454(.A1(new_n17751_), .A2(new_n17476_), .Z(new_n17752_));
  INV_X1     g17455(.I(new_n17752_), .ZN(new_n17753_));
  AOI22_X1   g17456(.A1(new_n13078_), .A2(\b[14] ), .B1(new_n1111_), .B2(new_n12218_), .ZN(new_n17754_));
  OAI21_X1   g17457(.A1(new_n17754_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n17755_));
  XOR2_X1    g17458(.A1(new_n1114_), .A2(new_n17755_), .Z(new_n17756_));
  OAI22_X1   g17459(.A1(new_n13880_), .A2(new_n921_), .B1(new_n706_), .B2(new_n13885_), .ZN(new_n17757_));
  AOI21_X1   g17460(.A1(new_n17757_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n17758_));
  XOR2_X1    g17461(.A1(new_n860_), .A2(new_n17758_), .Z(new_n17759_));
  NAND2_X1   g17462(.A1(new_n17471_), .A2(new_n17177_), .ZN(new_n17760_));
  NAND2_X1   g17463(.A1(new_n17760_), .A2(new_n17470_), .ZN(new_n17761_));
  NOR2_X1    g17464(.A1(new_n13476_), .A2(new_n565_), .ZN(new_n17762_));
  XOR2_X1    g17465(.A1(new_n14736_), .A2(new_n565_), .Z(new_n17763_));
  NAND2_X1   g17466(.A1(new_n17763_), .A2(\b[10] ), .ZN(new_n17764_));
  XOR2_X1    g17467(.A1(new_n17764_), .A2(new_n17762_), .Z(new_n17765_));
  NOR2_X1    g17468(.A1(new_n17761_), .A2(new_n17765_), .ZN(new_n17766_));
  INV_X1     g17469(.I(new_n17766_), .ZN(new_n17767_));
  NAND2_X1   g17470(.A1(new_n17761_), .A2(new_n17765_), .ZN(new_n17768_));
  NAND2_X1   g17471(.A1(new_n17767_), .A2(new_n17768_), .ZN(new_n17769_));
  INV_X1     g17472(.I(new_n17765_), .ZN(new_n17770_));
  XOR2_X1    g17473(.A1(new_n17761_), .A2(new_n17770_), .Z(new_n17771_));
  NOR2_X1    g17474(.A1(new_n17759_), .A2(new_n17771_), .ZN(new_n17772_));
  AOI21_X1   g17475(.A1(new_n17759_), .A2(new_n17769_), .B(new_n17772_), .ZN(new_n17773_));
  INV_X1     g17476(.I(new_n17773_), .ZN(new_n17774_));
  NAND2_X1   g17477(.A1(new_n17756_), .A2(new_n17774_), .ZN(new_n17775_));
  INV_X1     g17478(.I(new_n17775_), .ZN(new_n17776_));
  NOR2_X1    g17479(.A1(new_n17756_), .A2(new_n17774_), .ZN(new_n17777_));
  OAI21_X1   g17480(.A1(new_n17776_), .A2(new_n17777_), .B(new_n17753_), .ZN(new_n17778_));
  XOR2_X1    g17481(.A1(new_n17756_), .A2(new_n17773_), .Z(new_n17779_));
  OAI21_X1   g17482(.A1(new_n17753_), .A2(new_n17779_), .B(new_n17778_), .ZN(new_n17780_));
  INV_X1     g17483(.I(new_n17780_), .ZN(new_n17781_));
  NAND2_X1   g17484(.A1(new_n17457_), .A2(new_n17488_), .ZN(new_n17782_));
  AND2_X2    g17485(.A1(new_n17782_), .A2(new_n17487_), .Z(new_n17783_));
  AOI22_X1   g17486(.A1(new_n10969_), .A2(new_n1520_), .B1(new_n11394_), .B2(\b[17] ), .ZN(new_n17784_));
  OAI21_X1   g17487(.A1(new_n17784_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n17785_));
  XOR2_X1    g17488(.A1(new_n1421_), .A2(new_n17785_), .Z(new_n17786_));
  NOR2_X1    g17489(.A1(new_n17783_), .A2(new_n17786_), .ZN(new_n17787_));
  AND2_X2    g17490(.A1(new_n17783_), .A2(new_n17786_), .Z(new_n17788_));
  NOR2_X1    g17491(.A1(new_n17788_), .A2(new_n17787_), .ZN(new_n17789_));
  NOR2_X1    g17492(.A1(new_n17789_), .A2(new_n17781_), .ZN(new_n17790_));
  XNOR2_X1   g17493(.A1(new_n17783_), .A2(new_n17786_), .ZN(new_n17791_));
  NOR2_X1    g17494(.A1(new_n17791_), .A2(new_n17780_), .ZN(new_n17792_));
  NOR2_X1    g17495(.A1(new_n17790_), .A2(new_n17792_), .ZN(new_n17793_));
  NOR2_X1    g17496(.A1(new_n17491_), .A2(new_n17499_), .ZN(new_n17794_));
  NOR2_X1    g17497(.A1(new_n17794_), .A2(new_n17496_), .ZN(new_n17795_));
  NOR2_X1    g17498(.A1(new_n17793_), .A2(new_n17795_), .ZN(new_n17796_));
  INV_X1     g17499(.I(new_n17795_), .ZN(new_n17797_));
  NOR3_X1    g17500(.A1(new_n17797_), .A2(new_n17790_), .A3(new_n17792_), .ZN(new_n17798_));
  OAI21_X1   g17501(.A1(new_n17796_), .A2(new_n17798_), .B(new_n17750_), .ZN(new_n17799_));
  XOR2_X1    g17502(.A1(new_n17793_), .A2(new_n17797_), .Z(new_n17800_));
  OAI21_X1   g17503(.A1(new_n17800_), .A2(new_n17750_), .B(new_n17799_), .ZN(new_n17801_));
  NAND2_X1   g17504(.A1(new_n17514_), .A2(new_n17512_), .ZN(new_n17802_));
  OAI22_X1   g17505(.A1(new_n8644_), .A2(new_n2102_), .B1(new_n2281_), .B2(new_n9388_), .ZN(new_n17803_));
  OAI21_X1   g17506(.A1(new_n1936_), .A2(new_n10154_), .B(new_n17803_), .ZN(new_n17804_));
  AOI21_X1   g17507(.A1(new_n17804_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n17805_));
  XNOR2_X1   g17508(.A1(new_n2280_), .A2(new_n17805_), .ZN(new_n17806_));
  AOI21_X1   g17509(.A1(new_n17802_), .A2(new_n17513_), .B(new_n17806_), .ZN(new_n17807_));
  NAND2_X1   g17510(.A1(new_n17802_), .A2(new_n17513_), .ZN(new_n17808_));
  INV_X1     g17511(.I(new_n17806_), .ZN(new_n17809_));
  NOR2_X1    g17512(.A1(new_n17808_), .A2(new_n17809_), .ZN(new_n17810_));
  OAI21_X1   g17513(.A1(new_n17807_), .A2(new_n17810_), .B(new_n17801_), .ZN(new_n17811_));
  XOR2_X1    g17514(.A1(new_n17808_), .A2(new_n17806_), .Z(new_n17812_));
  OAI21_X1   g17515(.A1(new_n17801_), .A2(new_n17812_), .B(new_n17811_), .ZN(new_n17813_));
  OAI21_X1   g17516(.A1(new_n17516_), .A2(new_n17454_), .B(new_n17449_), .ZN(new_n17814_));
  OAI21_X1   g17517(.A1(new_n17453_), .A2(new_n17518_), .B(new_n17814_), .ZN(new_n17815_));
  NAND2_X1   g17518(.A1(new_n17813_), .A2(new_n17815_), .ZN(new_n17816_));
  OR2_X2     g17519(.A1(new_n17813_), .A2(new_n17815_), .Z(new_n17817_));
  AOI21_X1   g17520(.A1(new_n17817_), .A2(new_n17816_), .B(new_n17746_), .ZN(new_n17818_));
  XOR2_X1    g17521(.A1(new_n17813_), .A2(new_n17815_), .Z(new_n17819_));
  AOI21_X1   g17522(.A1(new_n17819_), .A2(new_n17746_), .B(new_n17818_), .ZN(new_n17820_));
  NOR2_X1    g17523(.A1(new_n17533_), .A2(new_n17531_), .ZN(new_n17821_));
  NOR2_X1    g17524(.A1(new_n17821_), .A2(new_n17532_), .ZN(new_n17822_));
  OAI22_X1   g17525(.A1(new_n6644_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n6647_), .ZN(new_n17823_));
  OAI21_X1   g17526(.A1(new_n3018_), .A2(new_n7284_), .B(new_n17823_), .ZN(new_n17824_));
  AOI21_X1   g17527(.A1(new_n17824_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n17825_));
  XNOR2_X1   g17528(.A1(new_n3514_), .A2(new_n17825_), .ZN(new_n17826_));
  INV_X1     g17529(.I(new_n17826_), .ZN(new_n17827_));
  XOR2_X1    g17530(.A1(new_n17822_), .A2(new_n17827_), .Z(new_n17828_));
  NOR2_X1    g17531(.A1(new_n17828_), .A2(new_n17820_), .ZN(new_n17829_));
  INV_X1     g17532(.I(new_n17820_), .ZN(new_n17830_));
  OAI21_X1   g17533(.A1(new_n17821_), .A2(new_n17532_), .B(new_n17827_), .ZN(new_n17831_));
  NAND2_X1   g17534(.A1(new_n17822_), .A2(new_n17826_), .ZN(new_n17832_));
  AOI21_X1   g17535(.A1(new_n17832_), .A2(new_n17831_), .B(new_n17830_), .ZN(new_n17833_));
  NOR2_X1    g17536(.A1(new_n17829_), .A2(new_n17833_), .ZN(new_n17834_));
  XOR2_X1    g17537(.A1(new_n17834_), .A2(new_n17742_), .Z(new_n17835_));
  NOR3_X1    g17538(.A1(new_n17834_), .A2(new_n17740_), .A3(new_n17741_), .ZN(new_n17836_));
  NOR3_X1    g17539(.A1(new_n17829_), .A2(new_n17742_), .A3(new_n17833_), .ZN(new_n17837_));
  OAI21_X1   g17540(.A1(new_n17837_), .A2(new_n17836_), .B(new_n17735_), .ZN(new_n17838_));
  OAI21_X1   g17541(.A1(new_n17735_), .A2(new_n17835_), .B(new_n17838_), .ZN(new_n17839_));
  OAI22_X1   g17542(.A1(new_n5420_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n5107_), .ZN(new_n17840_));
  OAI21_X1   g17543(.A1(new_n4500_), .A2(new_n5112_), .B(new_n17840_), .ZN(new_n17841_));
  AOI21_X1   g17544(.A1(new_n17841_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n17842_));
  XOR2_X1    g17545(.A1(new_n5067_), .A2(new_n17842_), .Z(new_n17843_));
  XNOR2_X1   g17546(.A1(new_n17839_), .A2(new_n17843_), .ZN(new_n17844_));
  NOR2_X1    g17547(.A1(new_n17844_), .A2(new_n17733_), .ZN(new_n17845_));
  NOR2_X1    g17548(.A1(new_n17839_), .A2(new_n17843_), .ZN(new_n17846_));
  INV_X1     g17549(.I(new_n17846_), .ZN(new_n17847_));
  NAND2_X1   g17550(.A1(new_n17839_), .A2(new_n17843_), .ZN(new_n17848_));
  AOI21_X1   g17551(.A1(new_n17847_), .A2(new_n17848_), .B(new_n17732_), .ZN(new_n17849_));
  NOR2_X1    g17552(.A1(new_n17845_), .A2(new_n17849_), .ZN(new_n17850_));
  INV_X1     g17553(.I(new_n17850_), .ZN(new_n17851_));
  OAI22_X1   g17554(.A1(new_n4072_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n4067_), .ZN(new_n17852_));
  OAI21_X1   g17555(.A1(new_n5353_), .A2(new_n4318_), .B(new_n17852_), .ZN(new_n17853_));
  AOI21_X1   g17556(.A1(new_n17853_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n17854_));
  XOR2_X1    g17557(.A1(new_n5926_), .A2(new_n17854_), .Z(new_n17855_));
  NOR2_X1    g17558(.A1(new_n17851_), .A2(new_n17855_), .ZN(new_n17856_));
  INV_X1     g17559(.I(new_n17856_), .ZN(new_n17857_));
  NAND2_X1   g17560(.A1(new_n17851_), .A2(new_n17855_), .ZN(new_n17858_));
  AOI21_X1   g17561(.A1(new_n17857_), .A2(new_n17858_), .B(new_n17731_), .ZN(new_n17859_));
  XOR2_X1    g17562(.A1(new_n17850_), .A2(new_n17855_), .Z(new_n17860_));
  NOR2_X1    g17563(.A1(new_n17860_), .A2(new_n17730_), .ZN(new_n17861_));
  NOR2_X1    g17564(.A1(new_n17859_), .A2(new_n17861_), .ZN(new_n17862_));
  OAI22_X1   g17565(.A1(new_n6538_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n6847_), .ZN(new_n17863_));
  OAI21_X1   g17566(.A1(new_n6229_), .A2(new_n3569_), .B(new_n17863_), .ZN(new_n17864_));
  AOI21_X1   g17567(.A1(new_n17864_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n17865_));
  XOR2_X1    g17568(.A1(new_n6851_), .A2(new_n17865_), .Z(new_n17866_));
  NOR2_X1    g17569(.A1(new_n17862_), .A2(new_n17866_), .ZN(new_n17867_));
  AND2_X2    g17570(.A1(new_n17862_), .A2(new_n17866_), .Z(new_n17868_));
  OAI21_X1   g17571(.A1(new_n17868_), .A2(new_n17867_), .B(new_n17729_), .ZN(new_n17869_));
  INV_X1     g17572(.I(new_n17729_), .ZN(new_n17870_));
  XOR2_X1    g17573(.A1(new_n17862_), .A2(new_n17866_), .Z(new_n17871_));
  NAND2_X1   g17574(.A1(new_n17871_), .A2(new_n17870_), .ZN(new_n17872_));
  NAND2_X1   g17575(.A1(new_n17872_), .A2(new_n17869_), .ZN(new_n17873_));
  OAI21_X1   g17576(.A1(new_n17593_), .A2(new_n17591_), .B(new_n17589_), .ZN(new_n17874_));
  OAI22_X1   g17577(.A1(new_n7864_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n7870_), .ZN(new_n17875_));
  OAI21_X1   g17578(.A1(new_n7198_), .A2(new_n2884_), .B(new_n17875_), .ZN(new_n17876_));
  AOI21_X1   g17579(.A1(new_n7874_), .A2(new_n2694_), .B(new_n17876_), .ZN(new_n17877_));
  XOR2_X1    g17580(.A1(new_n17874_), .A2(new_n17877_), .Z(new_n17878_));
  XOR2_X1    g17581(.A1(new_n17878_), .A2(new_n17873_), .Z(new_n17879_));
  OR2_X2     g17582(.A1(new_n17879_), .A2(\a[29] ), .Z(new_n17880_));
  NAND2_X1   g17583(.A1(new_n17879_), .A2(\a[29] ), .ZN(new_n17881_));
  NAND2_X1   g17584(.A1(new_n17880_), .A2(new_n17881_), .ZN(new_n17882_));
  OAI22_X1   g17585(.A1(new_n2171_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n2166_), .ZN(new_n17883_));
  OAI21_X1   g17586(.A1(new_n8218_), .A2(new_n2322_), .B(new_n17883_), .ZN(new_n17884_));
  AOI21_X1   g17587(.A1(new_n17884_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n17885_));
  XOR2_X1    g17588(.A1(new_n8952_), .A2(new_n17885_), .Z(new_n17886_));
  INV_X1     g17589(.I(new_n17886_), .ZN(new_n17887_));
  NAND2_X1   g17590(.A1(new_n17882_), .A2(new_n17887_), .ZN(new_n17888_));
  INV_X1     g17591(.I(new_n17888_), .ZN(new_n17889_));
  NOR2_X1    g17592(.A1(new_n17882_), .A2(new_n17887_), .ZN(new_n17890_));
  OAI21_X1   g17593(.A1(new_n17889_), .A2(new_n17890_), .B(new_n17727_), .ZN(new_n17891_));
  INV_X1     g17594(.I(new_n17727_), .ZN(new_n17892_));
  NOR2_X1    g17595(.A1(new_n17882_), .A2(new_n17886_), .ZN(new_n17893_));
  NAND2_X1   g17596(.A1(new_n17882_), .A2(new_n17886_), .ZN(new_n17894_));
  INV_X1     g17597(.I(new_n17894_), .ZN(new_n17895_));
  OAI21_X1   g17598(.A1(new_n17895_), .A2(new_n17893_), .B(new_n17892_), .ZN(new_n17896_));
  NAND2_X1   g17599(.A1(new_n17891_), .A2(new_n17896_), .ZN(new_n17897_));
  OAI21_X1   g17600(.A1(new_n17430_), .A2(new_n17613_), .B(new_n17625_), .ZN(new_n17898_));
  OAI22_X1   g17601(.A1(new_n1712_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n1707_), .ZN(new_n17899_));
  OAI21_X1   g17602(.A1(new_n9295_), .A2(new_n1850_), .B(new_n17899_), .ZN(new_n17900_));
  AOI21_X1   g17603(.A1(new_n10035_), .A2(new_n1702_), .B(new_n17900_), .ZN(new_n17901_));
  INV_X1     g17604(.I(new_n17901_), .ZN(new_n17902_));
  NOR2_X1    g17605(.A1(new_n17898_), .A2(new_n17902_), .ZN(new_n17903_));
  NAND2_X1   g17606(.A1(new_n17898_), .A2(new_n17902_), .ZN(new_n17904_));
  INV_X1     g17607(.I(new_n17904_), .ZN(new_n17905_));
  NOR2_X1    g17608(.A1(new_n17905_), .A2(new_n17903_), .ZN(new_n17906_));
  NOR2_X1    g17609(.A1(new_n17897_), .A2(new_n17906_), .ZN(new_n17907_));
  NAND2_X1   g17610(.A1(new_n17897_), .A2(new_n17906_), .ZN(new_n17908_));
  INV_X1     g17611(.I(new_n17908_), .ZN(new_n17909_));
  OAI21_X1   g17612(.A1(new_n17909_), .A2(new_n17907_), .B(new_n1709_), .ZN(new_n17910_));
  INV_X1     g17613(.I(new_n17907_), .ZN(new_n17911_));
  NAND3_X1   g17614(.A1(new_n17911_), .A2(new_n17908_), .A3(\a[23] ), .ZN(new_n17912_));
  OAI22_X1   g17615(.A1(new_n1347_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n1344_), .ZN(new_n17913_));
  OAI21_X1   g17616(.A1(new_n10477_), .A2(new_n1457_), .B(new_n17913_), .ZN(new_n17914_));
  AOI21_X1   g17617(.A1(new_n17914_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n17915_));
  XOR2_X1    g17618(.A1(new_n11298_), .A2(new_n17915_), .Z(new_n17916_));
  INV_X1     g17619(.I(new_n17916_), .ZN(new_n17917_));
  NAND3_X1   g17620(.A1(new_n17910_), .A2(new_n17912_), .A3(new_n17917_), .ZN(new_n17918_));
  AOI21_X1   g17621(.A1(new_n17911_), .A2(new_n17908_), .B(\a[23] ), .ZN(new_n17919_));
  NOR3_X1    g17622(.A1(new_n17909_), .A2(new_n17907_), .A3(new_n1709_), .ZN(new_n17920_));
  OAI21_X1   g17623(.A1(new_n17919_), .A2(new_n17920_), .B(new_n17916_), .ZN(new_n17921_));
  AOI21_X1   g17624(.A1(new_n17921_), .A2(new_n17918_), .B(new_n17723_), .ZN(new_n17922_));
  INV_X1     g17625(.I(new_n17723_), .ZN(new_n17923_));
  OAI21_X1   g17626(.A1(new_n17919_), .A2(new_n17920_), .B(new_n17917_), .ZN(new_n17924_));
  NAND3_X1   g17627(.A1(new_n17910_), .A2(new_n17912_), .A3(new_n17916_), .ZN(new_n17925_));
  AOI21_X1   g17628(.A1(new_n17924_), .A2(new_n17925_), .B(new_n17923_), .ZN(new_n17926_));
  OAI22_X1   g17629(.A1(new_n1055_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n1061_), .ZN(new_n17927_));
  OAI21_X1   g17630(.A1(new_n11744_), .A2(new_n1332_), .B(new_n17927_), .ZN(new_n17928_));
  AOI21_X1   g17631(.A1(new_n17928_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n17929_));
  XNOR2_X1   g17632(.A1(new_n12546_), .A2(new_n17929_), .ZN(new_n17930_));
  INV_X1     g17633(.I(new_n17930_), .ZN(new_n17931_));
  OAI21_X1   g17634(.A1(new_n17922_), .A2(new_n17926_), .B(new_n17931_), .ZN(new_n17932_));
  NOR3_X1    g17635(.A1(new_n17919_), .A2(new_n17920_), .A3(new_n17916_), .ZN(new_n17933_));
  AOI21_X1   g17636(.A1(new_n17910_), .A2(new_n17912_), .B(new_n17917_), .ZN(new_n17934_));
  OAI21_X1   g17637(.A1(new_n17934_), .A2(new_n17933_), .B(new_n17923_), .ZN(new_n17935_));
  AOI21_X1   g17638(.A1(new_n17910_), .A2(new_n17912_), .B(new_n17916_), .ZN(new_n17936_));
  NOR3_X1    g17639(.A1(new_n17919_), .A2(new_n17920_), .A3(new_n17917_), .ZN(new_n17937_));
  OAI21_X1   g17640(.A1(new_n17936_), .A2(new_n17937_), .B(new_n17723_), .ZN(new_n17938_));
  NAND3_X1   g17641(.A1(new_n17938_), .A2(new_n17935_), .A3(new_n17930_), .ZN(new_n17939_));
  AOI21_X1   g17642(.A1(new_n17932_), .A2(new_n17939_), .B(new_n17722_), .ZN(new_n17940_));
  INV_X1     g17643(.I(new_n17722_), .ZN(new_n17941_));
  NAND3_X1   g17644(.A1(new_n17938_), .A2(new_n17935_), .A3(new_n17931_), .ZN(new_n17942_));
  OAI21_X1   g17645(.A1(new_n17922_), .A2(new_n17926_), .B(new_n17930_), .ZN(new_n17943_));
  AOI21_X1   g17646(.A1(new_n17943_), .A2(new_n17942_), .B(new_n17941_), .ZN(new_n17944_));
  OAI22_X1   g17647(.A1(new_n970_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n820_), .ZN(new_n17945_));
  OAI21_X1   g17648(.A1(new_n12970_), .A2(new_n894_), .B(new_n17945_), .ZN(new_n17946_));
  AOI21_X1   g17649(.A1(new_n17946_), .A2(new_n827_), .B(new_n970_), .ZN(new_n17947_));
  XOR2_X1    g17650(.A1(new_n13784_), .A2(new_n17947_), .Z(new_n17948_));
  INV_X1     g17651(.I(new_n17948_), .ZN(new_n17949_));
  OAI21_X1   g17652(.A1(new_n17940_), .A2(new_n17944_), .B(new_n17949_), .ZN(new_n17950_));
  NOR3_X1    g17653(.A1(new_n17940_), .A2(new_n17944_), .A3(new_n17949_), .ZN(new_n17951_));
  INV_X1     g17654(.I(new_n17951_), .ZN(new_n17952_));
  AOI21_X1   g17655(.A1(new_n17952_), .A2(new_n17950_), .B(new_n17721_), .ZN(new_n17953_));
  INV_X1     g17656(.I(new_n17953_), .ZN(new_n17954_));
  OR3_X2     g17657(.A1(new_n17940_), .A2(new_n17944_), .A3(new_n17948_), .Z(new_n17955_));
  OAI21_X1   g17658(.A1(new_n17940_), .A2(new_n17944_), .B(new_n17948_), .ZN(new_n17956_));
  AOI21_X1   g17659(.A1(new_n17955_), .A2(new_n17956_), .B(new_n17720_), .ZN(new_n17957_));
  INV_X1     g17660(.I(new_n17957_), .ZN(new_n17958_));
  NOR2_X1    g17661(.A1(new_n684_), .A2(new_n610_), .ZN(new_n17959_));
  NAND2_X1   g17662(.A1(new_n16148_), .A2(new_n612_), .ZN(new_n17960_));
  OAI21_X1   g17663(.A1(new_n17959_), .A2(new_n17960_), .B(new_n606_), .ZN(new_n17961_));
  XNOR2_X1   g17664(.A1(new_n14978_), .A2(new_n17961_), .ZN(new_n17962_));
  INV_X1     g17665(.I(new_n17962_), .ZN(new_n17963_));
  NAND3_X1   g17666(.A1(new_n17954_), .A2(new_n17958_), .A3(new_n17963_), .ZN(new_n17964_));
  OAI21_X1   g17667(.A1(new_n17953_), .A2(new_n17957_), .B(new_n17962_), .ZN(new_n17965_));
  AOI21_X1   g17668(.A1(new_n17964_), .A2(new_n17965_), .B(new_n17718_), .ZN(new_n17966_));
  OAI21_X1   g17669(.A1(new_n17953_), .A2(new_n17957_), .B(new_n17963_), .ZN(new_n17967_));
  NAND3_X1   g17670(.A1(new_n17954_), .A2(new_n17958_), .A3(new_n17962_), .ZN(new_n17968_));
  AOI21_X1   g17671(.A1(new_n17968_), .A2(new_n17967_), .B(new_n17717_), .ZN(new_n17969_));
  NOR2_X1    g17672(.A1(new_n17966_), .A2(new_n17969_), .ZN(new_n17970_));
  NOR2_X1    g17673(.A1(new_n17970_), .A2(new_n17715_), .ZN(new_n17971_));
  XOR2_X1    g17674(.A1(new_n17713_), .A2(new_n17971_), .Z(new_n17972_));
  XOR2_X1    g17675(.A1(new_n17972_), .A2(new_n17708_), .Z(\f[73] ));
  AOI21_X1   g17676(.A1(new_n17970_), .A2(new_n17715_), .B(new_n17703_), .ZN(new_n17974_));
  INV_X1     g17677(.I(new_n17974_), .ZN(new_n17975_));
  NOR3_X1    g17678(.A1(new_n17410_), .A2(new_n17712_), .A3(new_n17975_), .ZN(new_n17976_));
  NOR2_X1    g17679(.A1(new_n17976_), .A2(new_n17971_), .ZN(new_n17977_));
  NAND2_X1   g17680(.A1(new_n17968_), .A2(new_n17717_), .ZN(new_n17978_));
  AND2_X2    g17681(.A1(new_n17978_), .A2(new_n17967_), .Z(new_n17979_));
  AOI21_X1   g17682(.A1(new_n17923_), .A2(new_n17921_), .B(new_n17933_), .ZN(new_n17980_));
  INV_X1     g17683(.I(new_n17980_), .ZN(new_n17981_));
  OAI21_X1   g17684(.A1(new_n17892_), .A2(new_n17890_), .B(new_n17888_), .ZN(new_n17982_));
  NOR2_X1    g17685(.A1(new_n17868_), .A2(new_n17870_), .ZN(new_n17983_));
  NOR2_X1    g17686(.A1(new_n17983_), .A2(new_n17867_), .ZN(new_n17984_));
  AOI21_X1   g17687(.A1(new_n17732_), .A2(new_n17848_), .B(new_n17846_), .ZN(new_n17985_));
  OAI22_X1   g17688(.A1(new_n4072_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n4067_), .ZN(new_n17986_));
  OAI21_X1   g17689(.A1(new_n5913_), .A2(new_n4318_), .B(new_n17986_), .ZN(new_n17987_));
  AOI21_X1   g17690(.A1(new_n17987_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n17988_));
  XOR2_X1    g17691(.A1(new_n6233_), .A2(new_n17988_), .Z(new_n17989_));
  NOR2_X1    g17692(.A1(new_n17836_), .A2(new_n17735_), .ZN(new_n17990_));
  NOR2_X1    g17693(.A1(new_n17990_), .A2(new_n17837_), .ZN(new_n17991_));
  OAI22_X1   g17694(.A1(new_n5420_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n5107_), .ZN(new_n17992_));
  OAI21_X1   g17695(.A1(new_n4774_), .A2(new_n5112_), .B(new_n17992_), .ZN(new_n17993_));
  AOI21_X1   g17696(.A1(new_n17993_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n17994_));
  XOR2_X1    g17697(.A1(new_n5357_), .A2(new_n17994_), .Z(new_n17995_));
  OAI22_X1   g17698(.A1(new_n6644_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n6647_), .ZN(new_n17996_));
  OAI21_X1   g17699(.A1(new_n3260_), .A2(new_n7284_), .B(new_n17996_), .ZN(new_n17997_));
  AOI21_X1   g17700(.A1(new_n17997_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n17998_));
  XOR2_X1    g17701(.A1(new_n3722_), .A2(new_n17998_), .Z(new_n17999_));
  INV_X1     g17702(.I(new_n17999_), .ZN(new_n18000_));
  OAI22_X1   g17703(.A1(new_n8644_), .A2(new_n2281_), .B1(new_n2439_), .B2(new_n9388_), .ZN(new_n18001_));
  OAI21_X1   g17704(.A1(new_n2102_), .A2(new_n10154_), .B(new_n18001_), .ZN(new_n18002_));
  AOI21_X1   g17705(.A1(new_n18002_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n18003_));
  XNOR2_X1   g17706(.A1(new_n2443_), .A2(new_n18003_), .ZN(new_n18004_));
  INV_X1     g17707(.I(new_n18004_), .ZN(new_n18005_));
  NOR2_X1    g17708(.A1(new_n17798_), .A2(new_n17749_), .ZN(new_n18006_));
  NOR2_X1    g17709(.A1(new_n18006_), .A2(new_n17796_), .ZN(new_n18007_));
  AOI22_X1   g17710(.A1(new_n11415_), .A2(new_n2097_), .B1(\b[21] ), .B2(new_n10145_), .ZN(new_n18008_));
  OAI21_X1   g17711(.A1(new_n18008_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n18009_));
  XOR2_X1    g17712(.A1(new_n1940_), .A2(new_n18009_), .Z(new_n18010_));
  AOI22_X1   g17713(.A1(new_n10969_), .A2(new_n1527_), .B1(new_n11394_), .B2(\b[18] ), .ZN(new_n18011_));
  OAI21_X1   g17714(.A1(new_n18011_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n18012_));
  XNOR2_X1   g17715(.A1(new_n1530_), .A2(new_n18012_), .ZN(new_n18013_));
  NAND2_X1   g17716(.A1(new_n17759_), .A2(new_n17767_), .ZN(new_n18014_));
  NAND2_X1   g17717(.A1(new_n18014_), .A2(new_n17768_), .ZN(new_n18015_));
  NOR2_X1    g17718(.A1(new_n13476_), .A2(new_n656_), .ZN(new_n18016_));
  XOR2_X1    g17719(.A1(new_n14736_), .A2(new_n656_), .Z(new_n18017_));
  NAND2_X1   g17720(.A1(new_n18017_), .A2(\b[11] ), .ZN(new_n18018_));
  XOR2_X1    g17721(.A1(new_n18018_), .A2(new_n18016_), .Z(new_n18019_));
  NOR2_X1    g17722(.A1(new_n17770_), .A2(new_n18019_), .ZN(new_n18020_));
  INV_X1     g17723(.I(new_n18019_), .ZN(new_n18021_));
  NOR2_X1    g17724(.A1(new_n18021_), .A2(new_n17765_), .ZN(new_n18022_));
  NOR2_X1    g17725(.A1(new_n18020_), .A2(new_n18022_), .ZN(new_n18023_));
  INV_X1     g17726(.I(new_n18023_), .ZN(new_n18024_));
  NAND2_X1   g17727(.A1(new_n18015_), .A2(new_n18024_), .ZN(new_n18025_));
  XOR2_X1    g17728(.A1(new_n17765_), .A2(new_n18019_), .Z(new_n18026_));
  OAI21_X1   g17729(.A1(new_n18015_), .A2(new_n18026_), .B(new_n18025_), .ZN(new_n18027_));
  INV_X1     g17730(.I(new_n18027_), .ZN(new_n18028_));
  AOI22_X1   g17731(.A1(new_n13078_), .A2(\b[15] ), .B1(new_n1292_), .B2(new_n12218_), .ZN(new_n18029_));
  OAI21_X1   g17732(.A1(new_n18029_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n18030_));
  XOR2_X1    g17733(.A1(new_n1196_), .A2(new_n18030_), .Z(new_n18031_));
  OAI22_X1   g17734(.A1(new_n13880_), .A2(new_n931_), .B1(new_n780_), .B2(new_n13885_), .ZN(new_n18032_));
  AOI21_X1   g17735(.A1(new_n18032_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n18033_));
  XNOR2_X1   g17736(.A1(new_n937_), .A2(new_n18033_), .ZN(new_n18034_));
  OR2_X2     g17737(.A1(new_n18031_), .A2(new_n18034_), .Z(new_n18035_));
  NAND2_X1   g17738(.A1(new_n18031_), .A2(new_n18034_), .ZN(new_n18036_));
  AOI21_X1   g17739(.A1(new_n18035_), .A2(new_n18036_), .B(new_n18028_), .ZN(new_n18037_));
  XNOR2_X1   g17740(.A1(new_n18031_), .A2(new_n18034_), .ZN(new_n18038_));
  NOR2_X1    g17741(.A1(new_n18038_), .A2(new_n18027_), .ZN(new_n18039_));
  NOR2_X1    g17742(.A1(new_n18039_), .A2(new_n18037_), .ZN(new_n18040_));
  OAI21_X1   g17743(.A1(new_n17752_), .A2(new_n17777_), .B(new_n17775_), .ZN(new_n18041_));
  XOR2_X1    g17744(.A1(new_n18040_), .A2(new_n18041_), .Z(new_n18042_));
  NOR2_X1    g17745(.A1(new_n18042_), .A2(new_n18013_), .ZN(new_n18043_));
  INV_X1     g17746(.I(new_n18013_), .ZN(new_n18044_));
  INV_X1     g17747(.I(new_n18041_), .ZN(new_n18045_));
  NOR2_X1    g17748(.A1(new_n18040_), .A2(new_n18045_), .ZN(new_n18046_));
  INV_X1     g17749(.I(new_n18046_), .ZN(new_n18047_));
  NAND2_X1   g17750(.A1(new_n18040_), .A2(new_n18045_), .ZN(new_n18048_));
  AOI21_X1   g17751(.A1(new_n18047_), .A2(new_n18048_), .B(new_n18044_), .ZN(new_n18049_));
  NOR2_X1    g17752(.A1(new_n18043_), .A2(new_n18049_), .ZN(new_n18050_));
  INV_X1     g17753(.I(new_n17788_), .ZN(new_n18051_));
  AOI21_X1   g17754(.A1(new_n18051_), .A2(new_n17780_), .B(new_n17787_), .ZN(new_n18052_));
  XOR2_X1    g17755(.A1(new_n18050_), .A2(new_n18052_), .Z(new_n18053_));
  INV_X1     g17756(.I(new_n18052_), .ZN(new_n18054_));
  NAND2_X1   g17757(.A1(new_n18050_), .A2(new_n18054_), .ZN(new_n18055_));
  INV_X1     g17758(.I(new_n18055_), .ZN(new_n18056_));
  NOR2_X1    g17759(.A1(new_n18050_), .A2(new_n18054_), .ZN(new_n18057_));
  OAI21_X1   g17760(.A1(new_n18056_), .A2(new_n18057_), .B(new_n18010_), .ZN(new_n18058_));
  OAI21_X1   g17761(.A1(new_n18010_), .A2(new_n18053_), .B(new_n18058_), .ZN(new_n18059_));
  XOR2_X1    g17762(.A1(new_n18059_), .A2(new_n18007_), .Z(new_n18060_));
  NAND2_X1   g17763(.A1(new_n18059_), .A2(new_n18007_), .ZN(new_n18061_));
  OR2_X2     g17764(.A1(new_n18059_), .A2(new_n18007_), .Z(new_n18062_));
  AOI21_X1   g17765(.A1(new_n18062_), .A2(new_n18061_), .B(new_n18005_), .ZN(new_n18063_));
  AOI21_X1   g17766(.A1(new_n18005_), .A2(new_n18060_), .B(new_n18063_), .ZN(new_n18064_));
  OAI22_X1   g17767(.A1(new_n7619_), .A2(new_n2842_), .B1(new_n3018_), .B2(new_n8309_), .ZN(new_n18065_));
  OAI21_X1   g17768(.A1(new_n2643_), .A2(new_n7947_), .B(new_n18065_), .ZN(new_n18066_));
  AOI21_X1   g17769(.A1(new_n18066_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n18067_));
  XNOR2_X1   g17770(.A1(new_n3022_), .A2(new_n18067_), .ZN(new_n18068_));
  INV_X1     g17771(.I(new_n17810_), .ZN(new_n18069_));
  AOI21_X1   g17772(.A1(new_n18069_), .A2(new_n17801_), .B(new_n17807_), .ZN(new_n18070_));
  XNOR2_X1   g17773(.A1(new_n18070_), .A2(new_n18068_), .ZN(new_n18071_));
  NOR2_X1    g17774(.A1(new_n18070_), .A2(new_n18068_), .ZN(new_n18072_));
  NAND2_X1   g17775(.A1(new_n18070_), .A2(new_n18068_), .ZN(new_n18073_));
  INV_X1     g17776(.I(new_n18073_), .ZN(new_n18074_));
  OAI21_X1   g17777(.A1(new_n18072_), .A2(new_n18074_), .B(new_n18064_), .ZN(new_n18075_));
  OAI21_X1   g17778(.A1(new_n18064_), .A2(new_n18071_), .B(new_n18075_), .ZN(new_n18076_));
  INV_X1     g17779(.I(new_n17746_), .ZN(new_n18077_));
  NAND2_X1   g17780(.A1(new_n17817_), .A2(new_n18077_), .ZN(new_n18078_));
  AND2_X2    g17781(.A1(new_n18078_), .A2(new_n17816_), .Z(new_n18079_));
  XNOR2_X1   g17782(.A1(new_n18076_), .A2(new_n18079_), .ZN(new_n18080_));
  INV_X1     g17783(.I(new_n18079_), .ZN(new_n18081_));
  NAND2_X1   g17784(.A1(new_n18076_), .A2(new_n18081_), .ZN(new_n18082_));
  INV_X1     g17785(.I(new_n18076_), .ZN(new_n18083_));
  NAND2_X1   g17786(.A1(new_n18083_), .A2(new_n18079_), .ZN(new_n18084_));
  AOI21_X1   g17787(.A1(new_n18084_), .A2(new_n18082_), .B(new_n18000_), .ZN(new_n18085_));
  AOI21_X1   g17788(.A1(new_n18000_), .A2(new_n18080_), .B(new_n18085_), .ZN(new_n18086_));
  OAI22_X1   g17789(.A1(new_n5993_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n5991_), .ZN(new_n18087_));
  OAI21_X1   g17790(.A1(new_n3989_), .A2(new_n5997_), .B(new_n18087_), .ZN(new_n18088_));
  AOI21_X1   g17791(.A1(new_n18088_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n18089_));
  XOR2_X1    g17792(.A1(new_n4499_), .A2(new_n18089_), .Z(new_n18090_));
  NAND2_X1   g17793(.A1(new_n17832_), .A2(new_n17830_), .ZN(new_n18091_));
  NAND2_X1   g17794(.A1(new_n18091_), .A2(new_n17831_), .ZN(new_n18092_));
  XOR2_X1    g17795(.A1(new_n18092_), .A2(new_n18090_), .Z(new_n18093_));
  AOI21_X1   g17796(.A1(new_n18091_), .A2(new_n17831_), .B(new_n18090_), .ZN(new_n18094_));
  INV_X1     g17797(.I(new_n18090_), .ZN(new_n18095_));
  NOR2_X1    g17798(.A1(new_n18092_), .A2(new_n18095_), .ZN(new_n18096_));
  OAI21_X1   g17799(.A1(new_n18094_), .A2(new_n18096_), .B(new_n18086_), .ZN(new_n18097_));
  OAI21_X1   g17800(.A1(new_n18086_), .A2(new_n18093_), .B(new_n18097_), .ZN(new_n18098_));
  XNOR2_X1   g17801(.A1(new_n18098_), .A2(new_n17995_), .ZN(new_n18099_));
  NOR2_X1    g17802(.A1(new_n18099_), .A2(new_n17991_), .ZN(new_n18100_));
  INV_X1     g17803(.I(new_n17991_), .ZN(new_n18101_));
  NAND2_X1   g17804(.A1(new_n18098_), .A2(new_n17995_), .ZN(new_n18102_));
  NOR2_X1    g17805(.A1(new_n18098_), .A2(new_n17995_), .ZN(new_n18103_));
  INV_X1     g17806(.I(new_n18103_), .ZN(new_n18104_));
  AOI21_X1   g17807(.A1(new_n18104_), .A2(new_n18102_), .B(new_n18101_), .ZN(new_n18105_));
  OAI21_X1   g17808(.A1(new_n18100_), .A2(new_n18105_), .B(new_n17989_), .ZN(new_n18106_));
  INV_X1     g17809(.I(new_n17989_), .ZN(new_n18107_));
  NOR2_X1    g17810(.A1(new_n18100_), .A2(new_n18105_), .ZN(new_n18108_));
  NAND2_X1   g17811(.A1(new_n18108_), .A2(new_n18107_), .ZN(new_n18109_));
  AOI21_X1   g17812(.A1(new_n18109_), .A2(new_n18106_), .B(new_n17985_), .ZN(new_n18110_));
  XOR2_X1    g17813(.A1(new_n18108_), .A2(new_n18107_), .Z(new_n18111_));
  AOI21_X1   g17814(.A1(new_n18111_), .A2(new_n17985_), .B(new_n18110_), .ZN(new_n18112_));
  AOI21_X1   g17815(.A1(new_n17730_), .A2(new_n17858_), .B(new_n17856_), .ZN(new_n18113_));
  OAI22_X1   g17816(.A1(new_n6847_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n7198_), .ZN(new_n18114_));
  OAI21_X1   g17817(.A1(new_n6538_), .A2(new_n3569_), .B(new_n18114_), .ZN(new_n18115_));
  AOI21_X1   g17818(.A1(new_n7202_), .A2(new_n3346_), .B(new_n18115_), .ZN(new_n18116_));
  XOR2_X1    g17819(.A1(new_n18113_), .A2(new_n18116_), .Z(new_n18117_));
  XOR2_X1    g17820(.A1(new_n18117_), .A2(new_n18112_), .Z(new_n18118_));
  XOR2_X1    g17821(.A1(new_n18118_), .A2(\a[32] ), .Z(new_n18119_));
  OAI22_X1   g17822(.A1(new_n7870_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n8218_), .ZN(new_n18120_));
  OAI21_X1   g17823(.A1(new_n7864_), .A2(new_n2884_), .B(new_n18120_), .ZN(new_n18121_));
  AOI21_X1   g17824(.A1(new_n18121_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n18122_));
  XOR2_X1    g17825(.A1(new_n8217_), .A2(new_n18122_), .Z(new_n18123_));
  XNOR2_X1   g17826(.A1(new_n18119_), .A2(new_n18123_), .ZN(new_n18124_));
  NOR2_X1    g17827(.A1(new_n18119_), .A2(new_n18123_), .ZN(new_n18125_));
  AND2_X2    g17828(.A1(new_n18119_), .A2(new_n18123_), .Z(new_n18126_));
  OAI21_X1   g17829(.A1(new_n18126_), .A2(new_n18125_), .B(new_n17984_), .ZN(new_n18127_));
  OAI21_X1   g17830(.A1(new_n17984_), .A2(new_n18124_), .B(new_n18127_), .ZN(new_n18128_));
  NAND2_X1   g17831(.A1(new_n17873_), .A2(new_n17874_), .ZN(new_n18129_));
  NOR2_X1    g17832(.A1(new_n17873_), .A2(new_n17874_), .ZN(new_n18130_));
  XOR2_X1    g17833(.A1(new_n17877_), .A2(\a[29] ), .Z(new_n18131_));
  OAI21_X1   g17834(.A1(new_n18130_), .A2(new_n18131_), .B(new_n18129_), .ZN(new_n18132_));
  OAI22_X1   g17835(.A1(new_n2171_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n2166_), .ZN(new_n18133_));
  OAI21_X1   g17836(.A1(new_n8563_), .A2(new_n2322_), .B(new_n18133_), .ZN(new_n18134_));
  AOI21_X1   g17837(.A1(new_n9299_), .A2(new_n2161_), .B(new_n18134_), .ZN(new_n18135_));
  XOR2_X1    g17838(.A1(new_n18132_), .A2(new_n18135_), .Z(new_n18136_));
  XOR2_X1    g17839(.A1(new_n18128_), .A2(new_n18136_), .Z(new_n18137_));
  XOR2_X1    g17840(.A1(new_n18137_), .A2(\a[26] ), .Z(new_n18138_));
  OAI22_X1   g17841(.A1(new_n1712_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n1707_), .ZN(new_n18139_));
  OAI21_X1   g17842(.A1(new_n10025_), .A2(new_n1850_), .B(new_n18139_), .ZN(new_n18140_));
  AOI21_X1   g17843(.A1(new_n18140_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n18141_));
  XOR2_X1    g17844(.A1(new_n10476_), .A2(new_n18141_), .Z(new_n18142_));
  NOR2_X1    g17845(.A1(new_n18138_), .A2(new_n18142_), .ZN(new_n18143_));
  AND2_X2    g17846(.A1(new_n18138_), .A2(new_n18142_), .Z(new_n18144_));
  OAI21_X1   g17847(.A1(new_n18144_), .A2(new_n18143_), .B(new_n17982_), .ZN(new_n18145_));
  INV_X1     g17848(.I(new_n17982_), .ZN(new_n18146_));
  XOR2_X1    g17849(.A1(new_n18138_), .A2(new_n18142_), .Z(new_n18147_));
  NAND2_X1   g17850(.A1(new_n18147_), .A2(new_n18146_), .ZN(new_n18148_));
  NAND2_X1   g17851(.A1(new_n18148_), .A2(new_n18145_), .ZN(new_n18149_));
  INV_X1     g17852(.I(new_n18149_), .ZN(new_n18150_));
  NAND2_X1   g17853(.A1(new_n17897_), .A2(new_n17898_), .ZN(new_n18151_));
  XOR2_X1    g17854(.A1(new_n17901_), .A2(\a[23] ), .Z(new_n18152_));
  OAI21_X1   g17855(.A1(new_n17897_), .A2(new_n17898_), .B(new_n18152_), .ZN(new_n18153_));
  NAND2_X1   g17856(.A1(new_n18153_), .A2(new_n18151_), .ZN(new_n18154_));
  OAI22_X1   g17857(.A1(new_n1347_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n1344_), .ZN(new_n18155_));
  OAI21_X1   g17858(.A1(new_n10862_), .A2(new_n1457_), .B(new_n18155_), .ZN(new_n18156_));
  AOI21_X1   g17859(.A1(new_n11748_), .A2(new_n1340_), .B(new_n18156_), .ZN(new_n18157_));
  XOR2_X1    g17860(.A1(new_n18154_), .A2(new_n18157_), .Z(new_n18158_));
  NAND2_X1   g17861(.A1(new_n18158_), .A2(new_n18150_), .ZN(new_n18159_));
  XNOR2_X1   g17862(.A1(new_n18154_), .A2(new_n18157_), .ZN(new_n18160_));
  NAND2_X1   g17863(.A1(new_n18160_), .A2(new_n18149_), .ZN(new_n18161_));
  AOI21_X1   g17864(.A1(new_n18161_), .A2(new_n18159_), .B(\a[20] ), .ZN(new_n18162_));
  NOR2_X1    g17865(.A1(new_n18160_), .A2(new_n18149_), .ZN(new_n18163_));
  NOR2_X1    g17866(.A1(new_n18158_), .A2(new_n18150_), .ZN(new_n18164_));
  NOR3_X1    g17867(.A1(new_n18163_), .A2(new_n18164_), .A3(new_n1346_), .ZN(new_n18165_));
  OAI22_X1   g17868(.A1(new_n1055_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n1061_), .ZN(new_n18166_));
  OAI21_X1   g17869(.A1(new_n12536_), .A2(new_n1332_), .B(new_n18166_), .ZN(new_n18167_));
  AOI21_X1   g17870(.A1(new_n18167_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n18168_));
  XOR2_X1    g17871(.A1(new_n12969_), .A2(new_n18168_), .Z(new_n18169_));
  NOR3_X1    g17872(.A1(new_n18162_), .A2(new_n18165_), .A3(new_n18169_), .ZN(new_n18170_));
  OAI21_X1   g17873(.A1(new_n18163_), .A2(new_n18164_), .B(new_n1346_), .ZN(new_n18171_));
  NAND3_X1   g17874(.A1(new_n18161_), .A2(new_n18159_), .A3(\a[20] ), .ZN(new_n18172_));
  INV_X1     g17875(.I(new_n18169_), .ZN(new_n18173_));
  AOI21_X1   g17876(.A1(new_n18171_), .A2(new_n18172_), .B(new_n18173_), .ZN(new_n18174_));
  OAI21_X1   g17877(.A1(new_n18170_), .A2(new_n18174_), .B(new_n17981_), .ZN(new_n18175_));
  AOI21_X1   g17878(.A1(new_n18171_), .A2(new_n18172_), .B(new_n18169_), .ZN(new_n18176_));
  NAND3_X1   g17879(.A1(new_n18171_), .A2(new_n18172_), .A3(new_n18169_), .ZN(new_n18177_));
  INV_X1     g17880(.I(new_n18177_), .ZN(new_n18178_));
  OAI21_X1   g17881(.A1(new_n18178_), .A2(new_n18176_), .B(new_n17980_), .ZN(new_n18179_));
  NAND2_X1   g17882(.A1(new_n18179_), .A2(new_n18175_), .ZN(new_n18180_));
  NOR3_X1    g17883(.A1(new_n17922_), .A2(new_n17926_), .A3(new_n17931_), .ZN(new_n18181_));
  OAI21_X1   g17884(.A1(new_n17722_), .A2(new_n18181_), .B(new_n17932_), .ZN(new_n18182_));
  INV_X1     g17885(.I(new_n14213_), .ZN(new_n18183_));
  OAI22_X1   g17886(.A1(new_n970_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n820_), .ZN(new_n18184_));
  OAI21_X1   g17887(.A1(new_n13367_), .A2(new_n894_), .B(new_n18184_), .ZN(new_n18185_));
  AOI21_X1   g17888(.A1(new_n18183_), .A2(new_n817_), .B(new_n18185_), .ZN(new_n18186_));
  XOR2_X1    g17889(.A1(new_n18182_), .A2(new_n18186_), .Z(new_n18187_));
  NOR2_X1    g17890(.A1(new_n18180_), .A2(new_n18187_), .ZN(new_n18188_));
  NAND3_X1   g17891(.A1(new_n18171_), .A2(new_n18172_), .A3(new_n18173_), .ZN(new_n18189_));
  OAI21_X1   g17892(.A1(new_n18162_), .A2(new_n18165_), .B(new_n18169_), .ZN(new_n18190_));
  AOI21_X1   g17893(.A1(new_n18190_), .A2(new_n18189_), .B(new_n17980_), .ZN(new_n18191_));
  OAI21_X1   g17894(.A1(new_n18162_), .A2(new_n18165_), .B(new_n18173_), .ZN(new_n18192_));
  AOI21_X1   g17895(.A1(new_n18192_), .A2(new_n18177_), .B(new_n17981_), .ZN(new_n18193_));
  NOR2_X1    g17896(.A1(new_n18191_), .A2(new_n18193_), .ZN(new_n18194_));
  INV_X1     g17897(.I(new_n18186_), .ZN(new_n18195_));
  XOR2_X1    g17898(.A1(new_n18182_), .A2(new_n18195_), .Z(new_n18196_));
  NOR2_X1    g17899(.A1(new_n18196_), .A2(new_n18194_), .ZN(new_n18197_));
  OAI21_X1   g17900(.A1(new_n18188_), .A2(new_n18197_), .B(new_n827_), .ZN(new_n18198_));
  NAND2_X1   g17901(.A1(new_n18196_), .A2(new_n18194_), .ZN(new_n18199_));
  NAND2_X1   g17902(.A1(new_n18180_), .A2(new_n18187_), .ZN(new_n18200_));
  NAND3_X1   g17903(.A1(new_n18200_), .A2(new_n18199_), .A3(\a[14] ), .ZN(new_n18201_));
  NAND2_X1   g17904(.A1(new_n18198_), .A2(new_n18201_), .ZN(new_n18202_));
  OAI21_X1   g17905(.A1(new_n17721_), .A2(new_n17951_), .B(new_n17950_), .ZN(new_n18203_));
  OAI21_X1   g17906(.A1(new_n607_), .A2(new_n684_), .B(new_n16487_), .ZN(new_n18204_));
  XOR2_X1    g17907(.A1(new_n18203_), .A2(new_n18204_), .Z(new_n18205_));
  INV_X1     g17908(.I(new_n18205_), .ZN(new_n18206_));
  NOR2_X1    g17909(.A1(new_n18202_), .A2(new_n18206_), .ZN(new_n18207_));
  AOI21_X1   g17910(.A1(new_n18198_), .A2(new_n18201_), .B(new_n18205_), .ZN(new_n18208_));
  OAI21_X1   g17911(.A1(new_n18207_), .A2(new_n18208_), .B(new_n612_), .ZN(new_n18209_));
  INV_X1     g17912(.I(new_n18209_), .ZN(new_n18210_));
  NOR3_X1    g17913(.A1(new_n18207_), .A2(new_n612_), .A3(new_n18208_), .ZN(new_n18211_));
  NOR2_X1    g17914(.A1(new_n18210_), .A2(new_n18211_), .ZN(new_n18212_));
  XOR2_X1    g17915(.A1(new_n18212_), .A2(new_n17979_), .Z(new_n18213_));
  INV_X1     g17916(.I(new_n17979_), .ZN(new_n18214_));
  OAI21_X1   g17917(.A1(new_n18210_), .A2(new_n18211_), .B(new_n18214_), .ZN(new_n18215_));
  NAND2_X1   g17918(.A1(new_n18212_), .A2(new_n17979_), .ZN(new_n18216_));
  NAND2_X1   g17919(.A1(new_n18216_), .A2(new_n18215_), .ZN(new_n18217_));
  MUX2_X1    g17920(.I0(new_n18213_), .I1(new_n18217_), .S(new_n17977_), .Z(\f[74] ));
  NAND2_X1   g17921(.A1(new_n18202_), .A2(new_n18203_), .ZN(new_n18219_));
  XOR2_X1    g17922(.A1(new_n18204_), .A2(new_n612_), .Z(new_n18220_));
  INV_X1     g17923(.I(new_n18220_), .ZN(new_n18221_));
  OAI21_X1   g17924(.A1(new_n18202_), .A2(new_n18203_), .B(new_n18221_), .ZN(new_n18222_));
  NAND2_X1   g17925(.A1(new_n18180_), .A2(new_n18182_), .ZN(new_n18223_));
  XOR2_X1    g17926(.A1(new_n18186_), .A2(\a[14] ), .Z(new_n18224_));
  INV_X1     g17927(.I(new_n18224_), .ZN(new_n18225_));
  OAI21_X1   g17928(.A1(new_n18180_), .A2(new_n18182_), .B(new_n18225_), .ZN(new_n18226_));
  NAND2_X1   g17929(.A1(new_n18226_), .A2(new_n18223_), .ZN(new_n18227_));
  AOI21_X1   g17930(.A1(new_n17981_), .A2(new_n18177_), .B(new_n18176_), .ZN(new_n18228_));
  NAND2_X1   g17931(.A1(new_n18149_), .A2(new_n18154_), .ZN(new_n18229_));
  NOR2_X1    g17932(.A1(new_n18149_), .A2(new_n18154_), .ZN(new_n18230_));
  XOR2_X1    g17933(.A1(new_n18157_), .A2(new_n1346_), .Z(new_n18231_));
  OAI21_X1   g17934(.A1(new_n18230_), .A2(new_n18231_), .B(new_n18229_), .ZN(new_n18232_));
  INV_X1     g17935(.I(new_n18232_), .ZN(new_n18233_));
  NOR2_X1    g17936(.A1(new_n18144_), .A2(new_n18146_), .ZN(new_n18234_));
  OR2_X2     g17937(.A1(new_n18234_), .A2(new_n18143_), .Z(new_n18235_));
  NAND2_X1   g17938(.A1(new_n18128_), .A2(new_n18132_), .ZN(new_n18236_));
  XOR2_X1    g17939(.A1(new_n18135_), .A2(new_n2168_), .Z(new_n18237_));
  OAI21_X1   g17940(.A1(new_n18128_), .A2(new_n18132_), .B(new_n18237_), .ZN(new_n18238_));
  NAND2_X1   g17941(.A1(new_n18238_), .A2(new_n18236_), .ZN(new_n18239_));
  NOR2_X1    g17942(.A1(new_n18126_), .A2(new_n17984_), .ZN(new_n18240_));
  NOR2_X1    g17943(.A1(new_n18240_), .A2(new_n18125_), .ZN(new_n18241_));
  NOR2_X1    g17944(.A1(new_n18113_), .A2(new_n18112_), .ZN(new_n18242_));
  NAND2_X1   g17945(.A1(new_n18113_), .A2(new_n18112_), .ZN(new_n18243_));
  XOR2_X1    g17946(.A1(new_n18116_), .A2(new_n3354_), .Z(new_n18244_));
  AOI21_X1   g17947(.A1(new_n18243_), .A2(new_n18244_), .B(new_n18242_), .ZN(new_n18245_));
  INV_X1     g17948(.I(new_n17985_), .ZN(new_n18246_));
  NAND2_X1   g17949(.A1(new_n18106_), .A2(new_n18246_), .ZN(new_n18247_));
  NAND2_X1   g17950(.A1(new_n18247_), .A2(new_n18109_), .ZN(new_n18248_));
  OAI21_X1   g17951(.A1(new_n17991_), .A2(new_n18103_), .B(new_n18102_), .ZN(new_n18249_));
  INV_X1     g17952(.I(new_n18249_), .ZN(new_n18250_));
  INV_X1     g17953(.I(new_n18096_), .ZN(new_n18251_));
  AOI21_X1   g17954(.A1(new_n18086_), .A2(new_n18251_), .B(new_n18094_), .ZN(new_n18252_));
  NAND2_X1   g17955(.A1(new_n18084_), .A2(new_n18000_), .ZN(new_n18253_));
  AOI21_X1   g17956(.A1(new_n18064_), .A2(new_n18073_), .B(new_n18072_), .ZN(new_n18254_));
  INV_X1     g17957(.I(new_n18254_), .ZN(new_n18255_));
  NAND2_X1   g17958(.A1(new_n18061_), .A2(new_n18005_), .ZN(new_n18256_));
  NAND2_X1   g17959(.A1(new_n18256_), .A2(new_n18062_), .ZN(new_n18257_));
  INV_X1     g17960(.I(new_n18257_), .ZN(new_n18258_));
  OAI21_X1   g17961(.A1(new_n18010_), .A2(new_n18057_), .B(new_n18055_), .ZN(new_n18259_));
  INV_X1     g17962(.I(new_n2103_), .ZN(new_n18260_));
  AOI22_X1   g17963(.A1(new_n11415_), .A2(new_n18260_), .B1(\b[22] ), .B2(new_n10145_), .ZN(new_n18261_));
  OAI21_X1   g17964(.A1(new_n18261_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n18262_));
  XOR2_X1    g17965(.A1(new_n2106_), .A2(new_n18262_), .Z(new_n18263_));
  AOI21_X1   g17966(.A1(new_n18044_), .A2(new_n18048_), .B(new_n18046_), .ZN(new_n18264_));
  INV_X1     g17967(.I(new_n18022_), .ZN(new_n18265_));
  AOI21_X1   g17968(.A1(new_n18015_), .A2(new_n18265_), .B(new_n18020_), .ZN(new_n18266_));
  OAI22_X1   g17969(.A1(new_n13880_), .A2(new_n1104_), .B1(new_n861_), .B2(new_n13885_), .ZN(new_n18267_));
  AOI21_X1   g17970(.A1(new_n18267_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n18268_));
  XOR2_X1    g17971(.A1(new_n1024_), .A2(new_n18268_), .Z(new_n18269_));
  NOR2_X1    g17972(.A1(new_n13476_), .A2(new_n706_), .ZN(new_n18270_));
  XOR2_X1    g17973(.A1(new_n14736_), .A2(new_n706_), .Z(new_n18271_));
  NAND2_X1   g17974(.A1(new_n18271_), .A2(\b[12] ), .ZN(new_n18272_));
  XOR2_X1    g17975(.A1(new_n18272_), .A2(new_n18270_), .Z(new_n18273_));
  XOR2_X1    g17976(.A1(new_n18273_), .A2(\a[11] ), .Z(new_n18274_));
  NOR2_X1    g17977(.A1(new_n18274_), .A2(new_n17765_), .ZN(new_n18275_));
  NOR2_X1    g17978(.A1(new_n18273_), .A2(new_n612_), .ZN(new_n18276_));
  INV_X1     g17979(.I(new_n18276_), .ZN(new_n18277_));
  NAND2_X1   g17980(.A1(new_n18273_), .A2(new_n612_), .ZN(new_n18278_));
  AOI21_X1   g17981(.A1(new_n18277_), .A2(new_n18278_), .B(new_n17770_), .ZN(new_n18279_));
  OAI21_X1   g17982(.A1(new_n18275_), .A2(new_n18279_), .B(new_n18269_), .ZN(new_n18280_));
  INV_X1     g17983(.I(new_n18269_), .ZN(new_n18281_));
  NOR2_X1    g17984(.A1(new_n18275_), .A2(new_n18279_), .ZN(new_n18282_));
  NAND2_X1   g17985(.A1(new_n18281_), .A2(new_n18282_), .ZN(new_n18283_));
  AOI21_X1   g17986(.A1(new_n18283_), .A2(new_n18280_), .B(new_n18266_), .ZN(new_n18284_));
  XNOR2_X1   g17987(.A1(new_n18269_), .A2(new_n18282_), .ZN(new_n18285_));
  AOI21_X1   g17988(.A1(new_n18285_), .A2(new_n18266_), .B(new_n18284_), .ZN(new_n18286_));
  INV_X1     g17989(.I(new_n18286_), .ZN(new_n18287_));
  AOI22_X1   g17990(.A1(new_n13078_), .A2(\b[16] ), .B1(new_n1296_), .B2(new_n12218_), .ZN(new_n18288_));
  OAI21_X1   g17991(.A1(new_n18288_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n18289_));
  XOR2_X1    g17992(.A1(new_n1299_), .A2(new_n18289_), .Z(new_n18290_));
  NAND2_X1   g17993(.A1(new_n18036_), .A2(new_n18027_), .ZN(new_n18291_));
  NAND2_X1   g17994(.A1(new_n18291_), .A2(new_n18035_), .ZN(new_n18292_));
  XOR2_X1    g17995(.A1(new_n18292_), .A2(new_n18290_), .Z(new_n18293_));
  NAND2_X1   g17996(.A1(new_n18293_), .A2(new_n18287_), .ZN(new_n18294_));
  NAND2_X1   g17997(.A1(new_n18292_), .A2(new_n18290_), .ZN(new_n18295_));
  INV_X1     g17998(.I(new_n18295_), .ZN(new_n18296_));
  NOR2_X1    g17999(.A1(new_n18292_), .A2(new_n18290_), .ZN(new_n18297_));
  OAI21_X1   g18000(.A1(new_n18296_), .A2(new_n18297_), .B(new_n18286_), .ZN(new_n18298_));
  NAND2_X1   g18001(.A1(new_n18294_), .A2(new_n18298_), .ZN(new_n18299_));
  AOI22_X1   g18002(.A1(new_n10969_), .A2(new_n1797_), .B1(new_n11394_), .B2(\b[19] ), .ZN(new_n18300_));
  OAI21_X1   g18003(.A1(new_n18300_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n18301_));
  XOR2_X1    g18004(.A1(new_n1638_), .A2(new_n18301_), .Z(new_n18302_));
  INV_X1     g18005(.I(new_n18302_), .ZN(new_n18303_));
  XOR2_X1    g18006(.A1(new_n18299_), .A2(new_n18303_), .Z(new_n18304_));
  NOR2_X1    g18007(.A1(new_n18304_), .A2(new_n18264_), .ZN(new_n18305_));
  INV_X1     g18008(.I(new_n18264_), .ZN(new_n18306_));
  NAND3_X1   g18009(.A1(new_n18294_), .A2(new_n18298_), .A3(new_n18303_), .ZN(new_n18307_));
  NAND2_X1   g18010(.A1(new_n18299_), .A2(new_n18302_), .ZN(new_n18308_));
  AOI21_X1   g18011(.A1(new_n18308_), .A2(new_n18307_), .B(new_n18306_), .ZN(new_n18309_));
  NOR2_X1    g18012(.A1(new_n18305_), .A2(new_n18309_), .ZN(new_n18310_));
  NOR2_X1    g18013(.A1(new_n18310_), .A2(new_n18263_), .ZN(new_n18311_));
  AND2_X2    g18014(.A1(new_n18310_), .A2(new_n18263_), .Z(new_n18312_));
  OAI21_X1   g18015(.A1(new_n18312_), .A2(new_n18311_), .B(new_n18259_), .ZN(new_n18313_));
  INV_X1     g18016(.I(new_n18259_), .ZN(new_n18314_));
  XOR2_X1    g18017(.A1(new_n18310_), .A2(new_n18263_), .Z(new_n18315_));
  NAND2_X1   g18018(.A1(new_n18315_), .A2(new_n18314_), .ZN(new_n18316_));
  NAND2_X1   g18019(.A1(new_n18316_), .A2(new_n18313_), .ZN(new_n18317_));
  OAI22_X1   g18020(.A1(new_n8644_), .A2(new_n2439_), .B1(new_n2643_), .B2(new_n9388_), .ZN(new_n18318_));
  OAI21_X1   g18021(.A1(new_n2281_), .A2(new_n10154_), .B(new_n18318_), .ZN(new_n18319_));
  AOI21_X1   g18022(.A1(new_n18319_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n18320_));
  XNOR2_X1   g18023(.A1(new_n2647_), .A2(new_n18320_), .ZN(new_n18321_));
  XOR2_X1    g18024(.A1(new_n18317_), .A2(new_n18321_), .Z(new_n18322_));
  INV_X1     g18025(.I(new_n18321_), .ZN(new_n18323_));
  NAND2_X1   g18026(.A1(new_n18317_), .A2(new_n18323_), .ZN(new_n18324_));
  INV_X1     g18027(.I(new_n18324_), .ZN(new_n18325_));
  NOR2_X1    g18028(.A1(new_n18317_), .A2(new_n18323_), .ZN(new_n18326_));
  OAI21_X1   g18029(.A1(new_n18325_), .A2(new_n18326_), .B(new_n18258_), .ZN(new_n18327_));
  OAI21_X1   g18030(.A1(new_n18258_), .A2(new_n18322_), .B(new_n18327_), .ZN(new_n18328_));
  OAI22_X1   g18031(.A1(new_n7619_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n8309_), .ZN(new_n18329_));
  OAI21_X1   g18032(.A1(new_n2842_), .A2(new_n7947_), .B(new_n18329_), .ZN(new_n18330_));
  AOI21_X1   g18033(.A1(new_n18330_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n18331_));
  XNOR2_X1   g18034(.A1(new_n3264_), .A2(new_n18331_), .ZN(new_n18332_));
  NOR2_X1    g18035(.A1(new_n18328_), .A2(new_n18332_), .ZN(new_n18333_));
  OR2_X2     g18036(.A1(new_n18322_), .A2(new_n18258_), .Z(new_n18334_));
  INV_X1     g18037(.I(new_n18332_), .ZN(new_n18335_));
  AOI21_X1   g18038(.A1(new_n18334_), .A2(new_n18327_), .B(new_n18335_), .ZN(new_n18336_));
  OAI21_X1   g18039(.A1(new_n18336_), .A2(new_n18333_), .B(new_n18255_), .ZN(new_n18337_));
  XOR2_X1    g18040(.A1(new_n18328_), .A2(new_n18335_), .Z(new_n18338_));
  OAI21_X1   g18041(.A1(new_n18338_), .A2(new_n18255_), .B(new_n18337_), .ZN(new_n18339_));
  OAI22_X1   g18042(.A1(new_n6644_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n6647_), .ZN(new_n18340_));
  OAI21_X1   g18043(.A1(new_n3709_), .A2(new_n7284_), .B(new_n18340_), .ZN(new_n18341_));
  AOI21_X1   g18044(.A1(new_n18341_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n18342_));
  XNOR2_X1   g18045(.A1(new_n3993_), .A2(new_n18342_), .ZN(new_n18343_));
  INV_X1     g18046(.I(new_n18343_), .ZN(new_n18344_));
  NAND2_X1   g18047(.A1(new_n18339_), .A2(new_n18344_), .ZN(new_n18345_));
  OR2_X2     g18048(.A1(new_n18339_), .A2(new_n18344_), .Z(new_n18346_));
  AOI22_X1   g18049(.A1(new_n18346_), .A2(new_n18345_), .B1(new_n18082_), .B2(new_n18253_), .ZN(new_n18347_));
  NAND2_X1   g18050(.A1(new_n18253_), .A2(new_n18082_), .ZN(new_n18348_));
  XOR2_X1    g18051(.A1(new_n18339_), .A2(new_n18343_), .Z(new_n18349_));
  NOR2_X1    g18052(.A1(new_n18349_), .A2(new_n18348_), .ZN(new_n18350_));
  NOR2_X1    g18053(.A1(new_n18350_), .A2(new_n18347_), .ZN(new_n18351_));
  OAI22_X1   g18054(.A1(new_n5993_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n5991_), .ZN(new_n18352_));
  OAI21_X1   g18055(.A1(new_n4253_), .A2(new_n5997_), .B(new_n18352_), .ZN(new_n18353_));
  AOI21_X1   g18056(.A1(new_n18353_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n18354_));
  XNOR2_X1   g18057(.A1(new_n4778_), .A2(new_n18354_), .ZN(new_n18355_));
  INV_X1     g18058(.I(new_n18355_), .ZN(new_n18356_));
  XOR2_X1    g18059(.A1(new_n18351_), .A2(new_n18356_), .Z(new_n18357_));
  NOR2_X1    g18060(.A1(new_n18357_), .A2(new_n18252_), .ZN(new_n18358_));
  INV_X1     g18061(.I(new_n18252_), .ZN(new_n18359_));
  OAI21_X1   g18062(.A1(new_n18350_), .A2(new_n18347_), .B(new_n18356_), .ZN(new_n18360_));
  NAND2_X1   g18063(.A1(new_n18351_), .A2(new_n18355_), .ZN(new_n18361_));
  AOI21_X1   g18064(.A1(new_n18361_), .A2(new_n18360_), .B(new_n18359_), .ZN(new_n18362_));
  NOR2_X1    g18065(.A1(new_n18358_), .A2(new_n18362_), .ZN(new_n18363_));
  OAI22_X1   g18066(.A1(new_n5420_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n5107_), .ZN(new_n18364_));
  OAI21_X1   g18067(.A1(new_n5068_), .A2(new_n5112_), .B(new_n18364_), .ZN(new_n18365_));
  AOI21_X1   g18068(.A1(new_n18365_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n18366_));
  XNOR2_X1   g18069(.A1(new_n5600_), .A2(new_n18366_), .ZN(new_n18367_));
  INV_X1     g18070(.I(new_n18367_), .ZN(new_n18368_));
  NAND2_X1   g18071(.A1(new_n18363_), .A2(new_n18368_), .ZN(new_n18369_));
  OAI21_X1   g18072(.A1(new_n18358_), .A2(new_n18362_), .B(new_n18367_), .ZN(new_n18370_));
  AOI21_X1   g18073(.A1(new_n18369_), .A2(new_n18370_), .B(new_n18250_), .ZN(new_n18371_));
  XOR2_X1    g18074(.A1(new_n18363_), .A2(new_n18367_), .Z(new_n18372_));
  NOR2_X1    g18075(.A1(new_n18372_), .A2(new_n18249_), .ZN(new_n18373_));
  NOR2_X1    g18076(.A1(new_n18373_), .A2(new_n18371_), .ZN(new_n18374_));
  OAI22_X1   g18077(.A1(new_n4072_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n4067_), .ZN(new_n18375_));
  OAI21_X1   g18078(.A1(new_n5921_), .A2(new_n4318_), .B(new_n18375_), .ZN(new_n18376_));
  AOI21_X1   g18079(.A1(new_n18376_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n18377_));
  XOR2_X1    g18080(.A1(new_n6543_), .A2(new_n18377_), .Z(new_n18378_));
  XOR2_X1    g18081(.A1(new_n18374_), .A2(new_n18378_), .Z(new_n18379_));
  INV_X1     g18082(.I(new_n18374_), .ZN(new_n18380_));
  INV_X1     g18083(.I(new_n18378_), .ZN(new_n18381_));
  NAND2_X1   g18084(.A1(new_n18380_), .A2(new_n18381_), .ZN(new_n18382_));
  NAND2_X1   g18085(.A1(new_n18374_), .A2(new_n18378_), .ZN(new_n18383_));
  AOI21_X1   g18086(.A1(new_n18382_), .A2(new_n18383_), .B(new_n18248_), .ZN(new_n18384_));
  AOI21_X1   g18087(.A1(new_n18248_), .A2(new_n18379_), .B(new_n18384_), .ZN(new_n18385_));
  OAI22_X1   g18088(.A1(new_n7198_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n7864_), .ZN(new_n18386_));
  OAI21_X1   g18089(.A1(new_n6847_), .A2(new_n3569_), .B(new_n18386_), .ZN(new_n18387_));
  AOI21_X1   g18090(.A1(new_n18387_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n18388_));
  XOR2_X1    g18091(.A1(new_n7516_), .A2(new_n18388_), .Z(new_n18389_));
  XOR2_X1    g18092(.A1(new_n18385_), .A2(new_n18389_), .Z(new_n18390_));
  NOR2_X1    g18093(.A1(new_n18390_), .A2(new_n18245_), .ZN(new_n18391_));
  INV_X1     g18094(.I(new_n18245_), .ZN(new_n18392_));
  INV_X1     g18095(.I(new_n18389_), .ZN(new_n18393_));
  NAND2_X1   g18096(.A1(new_n18385_), .A2(new_n18393_), .ZN(new_n18394_));
  NOR2_X1    g18097(.A1(new_n18385_), .A2(new_n18393_), .ZN(new_n18395_));
  INV_X1     g18098(.I(new_n18395_), .ZN(new_n18396_));
  AOI21_X1   g18099(.A1(new_n18396_), .A2(new_n18394_), .B(new_n18392_), .ZN(new_n18397_));
  NOR2_X1    g18100(.A1(new_n18391_), .A2(new_n18397_), .ZN(new_n18398_));
  OAI22_X1   g18101(.A1(new_n8218_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n8563_), .ZN(new_n18399_));
  OAI21_X1   g18102(.A1(new_n7870_), .A2(new_n2884_), .B(new_n18399_), .ZN(new_n18400_));
  AOI21_X1   g18103(.A1(new_n18400_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n18401_));
  XOR2_X1    g18104(.A1(new_n8568_), .A2(new_n18401_), .Z(new_n18402_));
  INV_X1     g18105(.I(new_n18402_), .ZN(new_n18403_));
  NAND2_X1   g18106(.A1(new_n18398_), .A2(new_n18403_), .ZN(new_n18404_));
  OAI21_X1   g18107(.A1(new_n18391_), .A2(new_n18397_), .B(new_n18402_), .ZN(new_n18405_));
  AOI21_X1   g18108(.A1(new_n18405_), .A2(new_n18404_), .B(new_n18241_), .ZN(new_n18406_));
  XOR2_X1    g18109(.A1(new_n18398_), .A2(new_n18403_), .Z(new_n18407_));
  AOI21_X1   g18110(.A1(new_n18241_), .A2(new_n18407_), .B(new_n18406_), .ZN(new_n18408_));
  OAI22_X1   g18111(.A1(new_n2171_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n2166_), .ZN(new_n18409_));
  OAI21_X1   g18112(.A1(new_n8948_), .A2(new_n2322_), .B(new_n18409_), .ZN(new_n18410_));
  AOI21_X1   g18113(.A1(new_n18410_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n18411_));
  XNOR2_X1   g18114(.A1(new_n9642_), .A2(new_n18411_), .ZN(new_n18412_));
  XOR2_X1    g18115(.A1(new_n18408_), .A2(new_n18412_), .Z(new_n18413_));
  NAND2_X1   g18116(.A1(new_n18413_), .A2(new_n18239_), .ZN(new_n18414_));
  INV_X1     g18117(.I(new_n18239_), .ZN(new_n18415_));
  NOR2_X1    g18118(.A1(new_n18408_), .A2(new_n18412_), .ZN(new_n18416_));
  AND2_X2    g18119(.A1(new_n18408_), .A2(new_n18412_), .Z(new_n18417_));
  OAI21_X1   g18120(.A1(new_n18417_), .A2(new_n18416_), .B(new_n18415_), .ZN(new_n18418_));
  OAI22_X1   g18121(.A1(new_n1712_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n1707_), .ZN(new_n18419_));
  OAI21_X1   g18122(.A1(new_n10031_), .A2(new_n1850_), .B(new_n18419_), .ZN(new_n18420_));
  AOI21_X1   g18123(.A1(new_n18420_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n18421_));
  XNOR2_X1   g18124(.A1(new_n10866_), .A2(new_n18421_), .ZN(new_n18422_));
  INV_X1     g18125(.I(new_n18422_), .ZN(new_n18423_));
  NAND3_X1   g18126(.A1(new_n18414_), .A2(new_n18418_), .A3(new_n18423_), .ZN(new_n18424_));
  NAND2_X1   g18127(.A1(new_n18414_), .A2(new_n18418_), .ZN(new_n18425_));
  NAND2_X1   g18128(.A1(new_n18425_), .A2(new_n18422_), .ZN(new_n18426_));
  NAND2_X1   g18129(.A1(new_n18426_), .A2(new_n18424_), .ZN(new_n18427_));
  NAND2_X1   g18130(.A1(new_n18235_), .A2(new_n18427_), .ZN(new_n18428_));
  NOR2_X1    g18131(.A1(new_n18234_), .A2(new_n18143_), .ZN(new_n18429_));
  XOR2_X1    g18132(.A1(new_n18425_), .A2(new_n18422_), .Z(new_n18430_));
  NAND2_X1   g18133(.A1(new_n18430_), .A2(new_n18429_), .ZN(new_n18431_));
  NAND2_X1   g18134(.A1(new_n18428_), .A2(new_n18431_), .ZN(new_n18432_));
  OAI22_X1   g18135(.A1(new_n1347_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n1344_), .ZN(new_n18433_));
  OAI21_X1   g18136(.A1(new_n11738_), .A2(new_n1457_), .B(new_n18433_), .ZN(new_n18434_));
  AOI21_X1   g18137(.A1(new_n18434_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n18435_));
  XNOR2_X1   g18138(.A1(new_n12128_), .A2(new_n18435_), .ZN(new_n18436_));
  NOR2_X1    g18139(.A1(new_n18432_), .A2(new_n18436_), .ZN(new_n18437_));
  INV_X1     g18140(.I(new_n18437_), .ZN(new_n18438_));
  NAND2_X1   g18141(.A1(new_n18432_), .A2(new_n18436_), .ZN(new_n18439_));
  AOI21_X1   g18142(.A1(new_n18438_), .A2(new_n18439_), .B(new_n18233_), .ZN(new_n18440_));
  INV_X1     g18143(.I(new_n18436_), .ZN(new_n18441_));
  NAND2_X1   g18144(.A1(new_n18432_), .A2(new_n18441_), .ZN(new_n18442_));
  NAND3_X1   g18145(.A1(new_n18428_), .A2(new_n18431_), .A3(new_n18436_), .ZN(new_n18443_));
  AOI21_X1   g18146(.A1(new_n18442_), .A2(new_n18443_), .B(new_n18232_), .ZN(new_n18444_));
  OAI22_X1   g18147(.A1(new_n1055_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n1061_), .ZN(new_n18445_));
  OAI21_X1   g18148(.A1(new_n12542_), .A2(new_n1332_), .B(new_n18445_), .ZN(new_n18446_));
  AOI21_X1   g18149(.A1(new_n18446_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n18447_));
  XNOR2_X1   g18150(.A1(new_n13371_), .A2(new_n18447_), .ZN(new_n18448_));
  NOR3_X1    g18151(.A1(new_n18440_), .A2(new_n18444_), .A3(new_n18448_), .ZN(new_n18449_));
  INV_X1     g18152(.I(new_n18449_), .ZN(new_n18450_));
  OAI21_X1   g18153(.A1(new_n18440_), .A2(new_n18444_), .B(new_n18448_), .ZN(new_n18451_));
  AOI21_X1   g18154(.A1(new_n18450_), .A2(new_n18451_), .B(new_n18228_), .ZN(new_n18452_));
  INV_X1     g18155(.I(new_n18228_), .ZN(new_n18453_));
  INV_X1     g18156(.I(new_n18448_), .ZN(new_n18454_));
  OAI21_X1   g18157(.A1(new_n18440_), .A2(new_n18444_), .B(new_n18454_), .ZN(new_n18455_));
  INV_X1     g18158(.I(new_n18439_), .ZN(new_n18456_));
  OAI21_X1   g18159(.A1(new_n18456_), .A2(new_n18437_), .B(new_n18232_), .ZN(new_n18457_));
  INV_X1     g18160(.I(new_n18444_), .ZN(new_n18458_));
  NAND3_X1   g18161(.A1(new_n18458_), .A2(new_n18457_), .A3(new_n18448_), .ZN(new_n18459_));
  AOI21_X1   g18162(.A1(new_n18455_), .A2(new_n18459_), .B(new_n18453_), .ZN(new_n18460_));
  OAI22_X1   g18163(.A1(new_n970_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n820_), .ZN(new_n18461_));
  OAI21_X1   g18164(.A1(new_n13785_), .A2(new_n894_), .B(new_n18461_), .ZN(new_n18462_));
  AOI21_X1   g18165(.A1(new_n18462_), .A2(new_n827_), .B(new_n970_), .ZN(new_n18463_));
  XNOR2_X1   g18166(.A1(new_n14599_), .A2(new_n18463_), .ZN(new_n18464_));
  INV_X1     g18167(.I(new_n18464_), .ZN(new_n18465_));
  OAI21_X1   g18168(.A1(new_n18460_), .A2(new_n18452_), .B(new_n18465_), .ZN(new_n18466_));
  INV_X1     g18169(.I(new_n18451_), .ZN(new_n18467_));
  OAI21_X1   g18170(.A1(new_n18467_), .A2(new_n18449_), .B(new_n18453_), .ZN(new_n18468_));
  NAND2_X1   g18171(.A1(new_n18459_), .A2(new_n18455_), .ZN(new_n18469_));
  NAND2_X1   g18172(.A1(new_n18469_), .A2(new_n18228_), .ZN(new_n18470_));
  NAND3_X1   g18173(.A1(new_n18468_), .A2(new_n18470_), .A3(new_n18464_), .ZN(new_n18471_));
  NAND2_X1   g18174(.A1(new_n18471_), .A2(new_n18466_), .ZN(new_n18472_));
  NAND3_X1   g18175(.A1(new_n18468_), .A2(new_n18470_), .A3(new_n18465_), .ZN(new_n18473_));
  OAI21_X1   g18176(.A1(new_n18460_), .A2(new_n18452_), .B(new_n18464_), .ZN(new_n18474_));
  AOI21_X1   g18177(.A1(new_n18473_), .A2(new_n18474_), .B(new_n18227_), .ZN(new_n18475_));
  AOI21_X1   g18178(.A1(new_n18227_), .A2(new_n18472_), .B(new_n18475_), .ZN(new_n18476_));
  AOI21_X1   g18179(.A1(new_n18219_), .A2(new_n18222_), .B(new_n18476_), .ZN(new_n18477_));
  NAND2_X1   g18180(.A1(new_n18222_), .A2(new_n18219_), .ZN(new_n18478_));
  NAND2_X1   g18181(.A1(new_n18473_), .A2(new_n18474_), .ZN(new_n18479_));
  MUX2_X1    g18182(.I0(new_n18479_), .I1(new_n18472_), .S(new_n18227_), .Z(new_n18480_));
  NOR2_X1    g18183(.A1(new_n18478_), .A2(new_n18480_), .ZN(new_n18481_));
  OAI21_X1   g18184(.A1(new_n18477_), .A2(new_n18481_), .B(new_n18213_), .ZN(new_n18482_));
  XNOR2_X1   g18185(.A1(new_n18482_), .A2(new_n18215_), .ZN(new_n18483_));
  XOR2_X1    g18186(.A1(new_n18483_), .A2(new_n17977_), .Z(\f[75] ));
  NAND3_X1   g18187(.A1(new_n18476_), .A2(new_n18222_), .A3(new_n18219_), .ZN(new_n18485_));
  NOR4_X1    g18188(.A1(new_n18477_), .A2(new_n18481_), .A3(new_n18210_), .A4(new_n18211_), .ZN(new_n18486_));
  OAI22_X1   g18189(.A1(new_n18477_), .A2(new_n18481_), .B1(new_n18210_), .B2(new_n18211_), .ZN(new_n18487_));
  AOI21_X1   g18190(.A1(new_n17979_), .A2(new_n18487_), .B(new_n18486_), .ZN(new_n18488_));
  OAI21_X1   g18191(.A1(new_n17976_), .A2(new_n17971_), .B(new_n18488_), .ZN(new_n18489_));
  NAND2_X1   g18192(.A1(new_n18227_), .A2(new_n18471_), .ZN(new_n18490_));
  AND2_X2    g18193(.A1(new_n18490_), .A2(new_n18466_), .Z(new_n18491_));
  AOI21_X1   g18194(.A1(new_n18453_), .A2(new_n18451_), .B(new_n18449_), .ZN(new_n18492_));
  INV_X1     g18195(.I(new_n18442_), .ZN(new_n18493_));
  AOI21_X1   g18196(.A1(new_n18232_), .A2(new_n18443_), .B(new_n18493_), .ZN(new_n18494_));
  NOR2_X1    g18197(.A1(new_n18417_), .A2(new_n18415_), .ZN(new_n18495_));
  NOR2_X1    g18198(.A1(new_n18495_), .A2(new_n18416_), .ZN(new_n18496_));
  OAI21_X1   g18199(.A1(new_n18125_), .A2(new_n18240_), .B(new_n18405_), .ZN(new_n18497_));
  AND2_X2    g18200(.A1(new_n18497_), .A2(new_n18404_), .Z(new_n18498_));
  OAI21_X1   g18201(.A1(new_n18245_), .A2(new_n18395_), .B(new_n18394_), .ZN(new_n18499_));
  OAI22_X1   g18202(.A1(new_n7864_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n7870_), .ZN(new_n18500_));
  OAI21_X1   g18203(.A1(new_n7198_), .A2(new_n3569_), .B(new_n18500_), .ZN(new_n18501_));
  AOI21_X1   g18204(.A1(new_n7874_), .A2(new_n3346_), .B(new_n18501_), .ZN(new_n18502_));
  NAND2_X1   g18205(.A1(new_n18383_), .A2(new_n18248_), .ZN(new_n18503_));
  NAND2_X1   g18206(.A1(new_n18503_), .A2(new_n18382_), .ZN(new_n18504_));
  NAND2_X1   g18207(.A1(new_n18370_), .A2(new_n18249_), .ZN(new_n18505_));
  NAND2_X1   g18208(.A1(new_n18505_), .A2(new_n18369_), .ZN(new_n18506_));
  OAI22_X1   g18209(.A1(new_n5420_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n5107_), .ZN(new_n18507_));
  OAI21_X1   g18210(.A1(new_n5353_), .A2(new_n5112_), .B(new_n18507_), .ZN(new_n18508_));
  AOI21_X1   g18211(.A1(new_n18508_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n18509_));
  XOR2_X1    g18212(.A1(new_n5926_), .A2(new_n18509_), .Z(new_n18510_));
  NAND2_X1   g18213(.A1(new_n18361_), .A2(new_n18359_), .ZN(new_n18511_));
  NAND2_X1   g18214(.A1(new_n18511_), .A2(new_n18360_), .ZN(new_n18512_));
  INV_X1     g18215(.I(new_n18512_), .ZN(new_n18513_));
  OAI22_X1   g18216(.A1(new_n5993_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n5991_), .ZN(new_n18514_));
  OAI21_X1   g18217(.A1(new_n4500_), .A2(new_n5997_), .B(new_n18514_), .ZN(new_n18515_));
  AOI21_X1   g18218(.A1(new_n18515_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n18516_));
  XOR2_X1    g18219(.A1(new_n5067_), .A2(new_n18516_), .Z(new_n18517_));
  NAND2_X1   g18220(.A1(new_n18346_), .A2(new_n18348_), .ZN(new_n18518_));
  NAND2_X1   g18221(.A1(new_n18518_), .A2(new_n18345_), .ZN(new_n18519_));
  OAI22_X1   g18222(.A1(new_n6644_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n6647_), .ZN(new_n18520_));
  OAI21_X1   g18223(.A1(new_n3717_), .A2(new_n7284_), .B(new_n18520_), .ZN(new_n18521_));
  AOI21_X1   g18224(.A1(new_n18521_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n18522_));
  XNOR2_X1   g18225(.A1(new_n4257_), .A2(new_n18522_), .ZN(new_n18523_));
  INV_X1     g18226(.I(new_n18523_), .ZN(new_n18524_));
  NOR2_X1    g18227(.A1(new_n18336_), .A2(new_n18254_), .ZN(new_n18525_));
  NOR2_X1    g18228(.A1(new_n18525_), .A2(new_n18333_), .ZN(new_n18526_));
  OAI22_X1   g18229(.A1(new_n7619_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n8309_), .ZN(new_n18527_));
  OAI21_X1   g18230(.A1(new_n3018_), .A2(new_n7947_), .B(new_n18527_), .ZN(new_n18528_));
  AOI21_X1   g18231(.A1(new_n18528_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n18529_));
  XNOR2_X1   g18232(.A1(new_n3514_), .A2(new_n18529_), .ZN(new_n18530_));
  INV_X1     g18233(.I(new_n18530_), .ZN(new_n18531_));
  OAI21_X1   g18234(.A1(new_n18258_), .A2(new_n18326_), .B(new_n18324_), .ZN(new_n18532_));
  AOI22_X1   g18235(.A1(new_n8631_), .A2(\b[27] ), .B1(\b[28] ), .B2(new_n9382_), .ZN(new_n18533_));
  AOI21_X1   g18236(.A1(\b[26] ), .A2(new_n9731_), .B(new_n18533_), .ZN(new_n18534_));
  OAI21_X1   g18237(.A1(new_n18534_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n18535_));
  XNOR2_X1   g18238(.A1(new_n2846_), .A2(new_n18535_), .ZN(new_n18536_));
  INV_X1     g18239(.I(new_n18536_), .ZN(new_n18537_));
  AOI22_X1   g18240(.A1(new_n10969_), .A2(new_n1805_), .B1(new_n11394_), .B2(\b[20] ), .ZN(new_n18538_));
  OAI21_X1   g18241(.A1(new_n18538_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n18539_));
  XOR2_X1    g18242(.A1(new_n1808_), .A2(new_n18539_), .Z(new_n18540_));
  OAI22_X1   g18243(.A1(new_n13880_), .A2(new_n1110_), .B1(new_n930_), .B2(new_n13885_), .ZN(new_n18541_));
  AOI21_X1   g18244(.A1(new_n18541_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n18542_));
  XNOR2_X1   g18245(.A1(new_n1114_), .A2(new_n18542_), .ZN(new_n18543_));
  NAND2_X1   g18246(.A1(new_n18278_), .A2(new_n17770_), .ZN(new_n18544_));
  NAND2_X1   g18247(.A1(new_n18544_), .A2(new_n18277_), .ZN(new_n18545_));
  NOR2_X1    g18248(.A1(new_n13476_), .A2(new_n780_), .ZN(new_n18546_));
  XOR2_X1    g18249(.A1(new_n14736_), .A2(new_n780_), .Z(new_n18547_));
  NAND2_X1   g18250(.A1(new_n18547_), .A2(\b[13] ), .ZN(new_n18548_));
  XOR2_X1    g18251(.A1(new_n18548_), .A2(new_n18546_), .Z(new_n18549_));
  NOR2_X1    g18252(.A1(new_n18545_), .A2(new_n18549_), .ZN(new_n18550_));
  NAND2_X1   g18253(.A1(new_n18545_), .A2(new_n18549_), .ZN(new_n18551_));
  INV_X1     g18254(.I(new_n18551_), .ZN(new_n18552_));
  NOR2_X1    g18255(.A1(new_n18552_), .A2(new_n18550_), .ZN(new_n18553_));
  INV_X1     g18256(.I(new_n18553_), .ZN(new_n18554_));
  NAND2_X1   g18257(.A1(new_n18543_), .A2(new_n18554_), .ZN(new_n18555_));
  INV_X1     g18258(.I(new_n18549_), .ZN(new_n18556_));
  XOR2_X1    g18259(.A1(new_n18545_), .A2(new_n18556_), .Z(new_n18557_));
  OAI21_X1   g18260(.A1(new_n18543_), .A2(new_n18557_), .B(new_n18555_), .ZN(new_n18558_));
  INV_X1     g18261(.I(new_n18558_), .ZN(new_n18559_));
  INV_X1     g18262(.I(new_n18266_), .ZN(new_n18560_));
  NAND2_X1   g18263(.A1(new_n18560_), .A2(new_n18280_), .ZN(new_n18561_));
  NAND2_X1   g18264(.A1(new_n18561_), .A2(new_n18283_), .ZN(new_n18562_));
  INV_X1     g18265(.I(new_n18562_), .ZN(new_n18563_));
  AOI22_X1   g18266(.A1(new_n13078_), .A2(\b[17] ), .B1(new_n1520_), .B2(new_n12218_), .ZN(new_n18564_));
  OAI21_X1   g18267(.A1(new_n18564_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n18565_));
  XOR2_X1    g18268(.A1(new_n1421_), .A2(new_n18565_), .Z(new_n18566_));
  OR2_X2     g18269(.A1(new_n18566_), .A2(new_n18563_), .Z(new_n18567_));
  NAND2_X1   g18270(.A1(new_n18566_), .A2(new_n18563_), .ZN(new_n18568_));
  AOI21_X1   g18271(.A1(new_n18567_), .A2(new_n18568_), .B(new_n18559_), .ZN(new_n18569_));
  XOR2_X1    g18272(.A1(new_n18566_), .A2(new_n18562_), .Z(new_n18570_));
  NOR2_X1    g18273(.A1(new_n18570_), .A2(new_n18558_), .ZN(new_n18571_));
  NOR2_X1    g18274(.A1(new_n18571_), .A2(new_n18569_), .ZN(new_n18572_));
  OAI21_X1   g18275(.A1(new_n18292_), .A2(new_n18290_), .B(new_n18287_), .ZN(new_n18573_));
  NAND2_X1   g18276(.A1(new_n18573_), .A2(new_n18295_), .ZN(new_n18574_));
  INV_X1     g18277(.I(new_n18574_), .ZN(new_n18575_));
  NOR2_X1    g18278(.A1(new_n18572_), .A2(new_n18575_), .ZN(new_n18576_));
  NAND2_X1   g18279(.A1(new_n18572_), .A2(new_n18575_), .ZN(new_n18577_));
  INV_X1     g18280(.I(new_n18577_), .ZN(new_n18578_));
  OAI21_X1   g18281(.A1(new_n18578_), .A2(new_n18576_), .B(new_n18540_), .ZN(new_n18579_));
  INV_X1     g18282(.I(new_n18540_), .ZN(new_n18580_));
  XOR2_X1    g18283(.A1(new_n18572_), .A2(new_n18575_), .Z(new_n18581_));
  NAND2_X1   g18284(.A1(new_n18581_), .A2(new_n18580_), .ZN(new_n18582_));
  NAND2_X1   g18285(.A1(new_n18582_), .A2(new_n18579_), .ZN(new_n18583_));
  NAND2_X1   g18286(.A1(new_n18308_), .A2(new_n18306_), .ZN(new_n18584_));
  NAND2_X1   g18287(.A1(new_n18584_), .A2(new_n18307_), .ZN(new_n18585_));
  AOI22_X1   g18288(.A1(new_n11415_), .A2(new_n2435_), .B1(\b[23] ), .B2(new_n10145_), .ZN(new_n18586_));
  OAI21_X1   g18289(.A1(new_n18586_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n18587_));
  XOR2_X1    g18290(.A1(new_n2280_), .A2(new_n18587_), .Z(new_n18588_));
  INV_X1     g18291(.I(new_n18588_), .ZN(new_n18589_));
  NAND2_X1   g18292(.A1(new_n18585_), .A2(new_n18589_), .ZN(new_n18590_));
  INV_X1     g18293(.I(new_n18590_), .ZN(new_n18591_));
  NOR2_X1    g18294(.A1(new_n18585_), .A2(new_n18589_), .ZN(new_n18592_));
  OAI21_X1   g18295(.A1(new_n18591_), .A2(new_n18592_), .B(new_n18583_), .ZN(new_n18593_));
  INV_X1     g18296(.I(new_n18583_), .ZN(new_n18594_));
  XOR2_X1    g18297(.A1(new_n18585_), .A2(new_n18589_), .Z(new_n18595_));
  NAND2_X1   g18298(.A1(new_n18595_), .A2(new_n18594_), .ZN(new_n18596_));
  NAND2_X1   g18299(.A1(new_n18596_), .A2(new_n18593_), .ZN(new_n18597_));
  NOR2_X1    g18300(.A1(new_n18311_), .A2(new_n18314_), .ZN(new_n18598_));
  NOR2_X1    g18301(.A1(new_n18598_), .A2(new_n18312_), .ZN(new_n18599_));
  XOR2_X1    g18302(.A1(new_n18599_), .A2(new_n18597_), .Z(new_n18600_));
  NOR2_X1    g18303(.A1(new_n18600_), .A2(new_n18537_), .ZN(new_n18601_));
  OAI21_X1   g18304(.A1(new_n18312_), .A2(new_n18598_), .B(new_n18597_), .ZN(new_n18602_));
  NAND3_X1   g18305(.A1(new_n18599_), .A2(new_n18593_), .A3(new_n18596_), .ZN(new_n18603_));
  AOI21_X1   g18306(.A1(new_n18602_), .A2(new_n18603_), .B(new_n18536_), .ZN(new_n18604_));
  NOR2_X1    g18307(.A1(new_n18601_), .A2(new_n18604_), .ZN(new_n18605_));
  XOR2_X1    g18308(.A1(new_n18605_), .A2(new_n18532_), .Z(new_n18606_));
  NAND2_X1   g18309(.A1(new_n18606_), .A2(new_n18531_), .ZN(new_n18607_));
  NOR2_X1    g18310(.A1(new_n18605_), .A2(new_n18532_), .ZN(new_n18608_));
  NAND2_X1   g18311(.A1(new_n18605_), .A2(new_n18532_), .ZN(new_n18609_));
  INV_X1     g18312(.I(new_n18609_), .ZN(new_n18610_));
  OAI21_X1   g18313(.A1(new_n18610_), .A2(new_n18608_), .B(new_n18530_), .ZN(new_n18611_));
  NAND2_X1   g18314(.A1(new_n18607_), .A2(new_n18611_), .ZN(new_n18612_));
  XOR2_X1    g18315(.A1(new_n18612_), .A2(new_n18526_), .Z(new_n18613_));
  NAND2_X1   g18316(.A1(new_n18613_), .A2(new_n18524_), .ZN(new_n18614_));
  INV_X1     g18317(.I(new_n18526_), .ZN(new_n18615_));
  INV_X1     g18318(.I(new_n18612_), .ZN(new_n18616_));
  NOR2_X1    g18319(.A1(new_n18616_), .A2(new_n18615_), .ZN(new_n18617_));
  NOR2_X1    g18320(.A1(new_n18612_), .A2(new_n18526_), .ZN(new_n18618_));
  OAI21_X1   g18321(.A1(new_n18617_), .A2(new_n18618_), .B(new_n18523_), .ZN(new_n18619_));
  NAND2_X1   g18322(.A1(new_n18614_), .A2(new_n18619_), .ZN(new_n18620_));
  XOR2_X1    g18323(.A1(new_n18620_), .A2(new_n18519_), .Z(new_n18621_));
  NOR2_X1    g18324(.A1(new_n18621_), .A2(new_n18517_), .ZN(new_n18622_));
  INV_X1     g18325(.I(new_n18517_), .ZN(new_n18623_));
  NAND3_X1   g18326(.A1(new_n18620_), .A2(new_n18345_), .A3(new_n18518_), .ZN(new_n18624_));
  NAND3_X1   g18327(.A1(new_n18519_), .A2(new_n18614_), .A3(new_n18619_), .ZN(new_n18625_));
  AOI21_X1   g18328(.A1(new_n18624_), .A2(new_n18625_), .B(new_n18623_), .ZN(new_n18626_));
  NOR2_X1    g18329(.A1(new_n18622_), .A2(new_n18626_), .ZN(new_n18627_));
  XOR2_X1    g18330(.A1(new_n18627_), .A2(new_n18513_), .Z(new_n18628_));
  NOR2_X1    g18331(.A1(new_n18628_), .A2(new_n18510_), .ZN(new_n18629_));
  INV_X1     g18332(.I(new_n18510_), .ZN(new_n18630_));
  OAI21_X1   g18333(.A1(new_n18622_), .A2(new_n18626_), .B(new_n18513_), .ZN(new_n18631_));
  NAND2_X1   g18334(.A1(new_n18627_), .A2(new_n18512_), .ZN(new_n18632_));
  AOI21_X1   g18335(.A1(new_n18631_), .A2(new_n18632_), .B(new_n18630_), .ZN(new_n18633_));
  NOR2_X1    g18336(.A1(new_n18629_), .A2(new_n18633_), .ZN(new_n18634_));
  OAI22_X1   g18337(.A1(new_n4072_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n4067_), .ZN(new_n18635_));
  OAI21_X1   g18338(.A1(new_n6229_), .A2(new_n4318_), .B(new_n18635_), .ZN(new_n18636_));
  AOI21_X1   g18339(.A1(new_n18636_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n18637_));
  XOR2_X1    g18340(.A1(new_n6851_), .A2(new_n18637_), .Z(new_n18638_));
  INV_X1     g18341(.I(new_n18638_), .ZN(new_n18639_));
  NAND2_X1   g18342(.A1(new_n18634_), .A2(new_n18639_), .ZN(new_n18640_));
  INV_X1     g18343(.I(new_n18640_), .ZN(new_n18641_));
  NOR2_X1    g18344(.A1(new_n18634_), .A2(new_n18639_), .ZN(new_n18642_));
  OAI21_X1   g18345(.A1(new_n18641_), .A2(new_n18642_), .B(new_n18506_), .ZN(new_n18643_));
  INV_X1     g18346(.I(new_n18506_), .ZN(new_n18644_));
  XOR2_X1    g18347(.A1(new_n18634_), .A2(new_n18639_), .Z(new_n18645_));
  NAND2_X1   g18348(.A1(new_n18645_), .A2(new_n18644_), .ZN(new_n18646_));
  NAND2_X1   g18349(.A1(new_n18646_), .A2(new_n18643_), .ZN(new_n18647_));
  XOR2_X1    g18350(.A1(new_n18647_), .A2(new_n18504_), .Z(new_n18648_));
  XOR2_X1    g18351(.A1(new_n18648_), .A2(new_n18502_), .Z(new_n18649_));
  XOR2_X1    g18352(.A1(new_n18649_), .A2(\a[32] ), .Z(new_n18650_));
  OAI22_X1   g18353(.A1(new_n8563_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n8948_), .ZN(new_n18651_));
  OAI21_X1   g18354(.A1(new_n8218_), .A2(new_n2884_), .B(new_n18651_), .ZN(new_n18652_));
  AOI21_X1   g18355(.A1(new_n18652_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n18653_));
  XOR2_X1    g18356(.A1(new_n8952_), .A2(new_n18653_), .Z(new_n18654_));
  NOR2_X1    g18357(.A1(new_n18650_), .A2(new_n18654_), .ZN(new_n18655_));
  XOR2_X1    g18358(.A1(new_n18649_), .A2(new_n3354_), .Z(new_n18656_));
  INV_X1     g18359(.I(new_n18654_), .ZN(new_n18657_));
  NOR2_X1    g18360(.A1(new_n18656_), .A2(new_n18657_), .ZN(new_n18658_));
  OAI21_X1   g18361(.A1(new_n18655_), .A2(new_n18658_), .B(new_n18499_), .ZN(new_n18659_));
  XOR2_X1    g18362(.A1(new_n18656_), .A2(new_n18654_), .Z(new_n18660_));
  OAI21_X1   g18363(.A1(new_n18660_), .A2(new_n18499_), .B(new_n18659_), .ZN(new_n18661_));
  OAI22_X1   g18364(.A1(new_n2171_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n2166_), .ZN(new_n18662_));
  OAI21_X1   g18365(.A1(new_n9295_), .A2(new_n2322_), .B(new_n18662_), .ZN(new_n18663_));
  AOI21_X1   g18366(.A1(new_n18663_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n18664_));
  XNOR2_X1   g18367(.A1(new_n10035_), .A2(new_n18664_), .ZN(new_n18665_));
  INV_X1     g18368(.I(new_n18665_), .ZN(new_n18666_));
  NAND2_X1   g18369(.A1(new_n18661_), .A2(new_n18666_), .ZN(new_n18667_));
  INV_X1     g18370(.I(new_n18661_), .ZN(new_n18668_));
  NAND2_X1   g18371(.A1(new_n18668_), .A2(new_n18665_), .ZN(new_n18669_));
  AOI21_X1   g18372(.A1(new_n18669_), .A2(new_n18667_), .B(new_n18498_), .ZN(new_n18670_));
  INV_X1     g18373(.I(new_n18498_), .ZN(new_n18671_));
  XOR2_X1    g18374(.A1(new_n18661_), .A2(new_n18665_), .Z(new_n18672_));
  NOR2_X1    g18375(.A1(new_n18672_), .A2(new_n18671_), .ZN(new_n18673_));
  OAI22_X1   g18376(.A1(new_n1712_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n1707_), .ZN(new_n18674_));
  OAI21_X1   g18377(.A1(new_n10477_), .A2(new_n1850_), .B(new_n18674_), .ZN(new_n18675_));
  AOI21_X1   g18378(.A1(new_n18675_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n18676_));
  XOR2_X1    g18379(.A1(new_n11298_), .A2(new_n18676_), .Z(new_n18677_));
  INV_X1     g18380(.I(new_n18677_), .ZN(new_n18678_));
  OAI21_X1   g18381(.A1(new_n18673_), .A2(new_n18670_), .B(new_n18678_), .ZN(new_n18679_));
  NOR2_X1    g18382(.A1(new_n18673_), .A2(new_n18670_), .ZN(new_n18680_));
  NAND2_X1   g18383(.A1(new_n18680_), .A2(new_n18677_), .ZN(new_n18681_));
  AOI21_X1   g18384(.A1(new_n18681_), .A2(new_n18679_), .B(new_n18496_), .ZN(new_n18682_));
  XOR2_X1    g18385(.A1(new_n18680_), .A2(new_n18677_), .Z(new_n18683_));
  AOI21_X1   g18386(.A1(new_n18496_), .A2(new_n18683_), .B(new_n18682_), .ZN(new_n18684_));
  INV_X1     g18387(.I(new_n18424_), .ZN(new_n18685_));
  AOI21_X1   g18388(.A1(new_n18235_), .A2(new_n18426_), .B(new_n18685_), .ZN(new_n18686_));
  NAND2_X1   g18389(.A1(new_n12546_), .A2(new_n1340_), .ZN(new_n18687_));
  AOI22_X1   g18390(.A1(\b[58] ), .A2(new_n1999_), .B1(new_n1340_), .B2(\b[57] ), .ZN(new_n18688_));
  AOI21_X1   g18391(.A1(\b[56] ), .A2(new_n1458_), .B(new_n18688_), .ZN(new_n18689_));
  NAND2_X1   g18392(.A1(new_n18687_), .A2(new_n18689_), .ZN(new_n18690_));
  XOR2_X1    g18393(.A1(new_n18686_), .A2(new_n18690_), .Z(new_n18691_));
  XOR2_X1    g18394(.A1(new_n18691_), .A2(new_n18684_), .Z(new_n18692_));
  XOR2_X1    g18395(.A1(new_n18692_), .A2(\a[20] ), .Z(new_n18693_));
  OAI22_X1   g18396(.A1(new_n1055_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n1061_), .ZN(new_n18694_));
  OAI21_X1   g18397(.A1(new_n12970_), .A2(new_n1332_), .B(new_n18694_), .ZN(new_n18695_));
  AOI21_X1   g18398(.A1(new_n18695_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n18696_));
  XOR2_X1    g18399(.A1(new_n13784_), .A2(new_n18696_), .Z(new_n18697_));
  INV_X1     g18400(.I(new_n18697_), .ZN(new_n18698_));
  NAND2_X1   g18401(.A1(new_n18693_), .A2(new_n18698_), .ZN(new_n18699_));
  XOR2_X1    g18402(.A1(new_n18692_), .A2(new_n1346_), .Z(new_n18700_));
  NAND2_X1   g18403(.A1(new_n18700_), .A2(new_n18697_), .ZN(new_n18701_));
  AOI21_X1   g18404(.A1(new_n18701_), .A2(new_n18699_), .B(new_n18494_), .ZN(new_n18702_));
  INV_X1     g18405(.I(new_n18494_), .ZN(new_n18703_));
  NAND2_X1   g18406(.A1(new_n18700_), .A2(new_n18698_), .ZN(new_n18704_));
  NAND2_X1   g18407(.A1(new_n18693_), .A2(new_n18697_), .ZN(new_n18705_));
  AOI21_X1   g18408(.A1(new_n18704_), .A2(new_n18705_), .B(new_n18703_), .ZN(new_n18706_));
  NOR2_X1    g18409(.A1(new_n18706_), .A2(new_n18702_), .ZN(new_n18707_));
  NOR2_X1    g18410(.A1(new_n894_), .A2(new_n820_), .ZN(new_n18708_));
  NAND2_X1   g18411(.A1(new_n16148_), .A2(new_n827_), .ZN(new_n18709_));
  OAI21_X1   g18412(.A1(new_n18708_), .A2(new_n18709_), .B(new_n817_), .ZN(new_n18710_));
  XNOR2_X1   g18413(.A1(new_n14978_), .A2(new_n18710_), .ZN(new_n18711_));
  INV_X1     g18414(.I(new_n18711_), .ZN(new_n18712_));
  NAND2_X1   g18415(.A1(new_n18707_), .A2(new_n18712_), .ZN(new_n18713_));
  INV_X1     g18416(.I(new_n18707_), .ZN(new_n18714_));
  NAND2_X1   g18417(.A1(new_n18714_), .A2(new_n18711_), .ZN(new_n18715_));
  AOI21_X1   g18418(.A1(new_n18715_), .A2(new_n18713_), .B(new_n18492_), .ZN(new_n18716_));
  INV_X1     g18419(.I(new_n18716_), .ZN(new_n18717_));
  NOR2_X1    g18420(.A1(new_n18707_), .A2(new_n18711_), .ZN(new_n18718_));
  NAND2_X1   g18421(.A1(new_n18707_), .A2(new_n18711_), .ZN(new_n18719_));
  INV_X1     g18422(.I(new_n18719_), .ZN(new_n18720_));
  OAI21_X1   g18423(.A1(new_n18720_), .A2(new_n18718_), .B(new_n18492_), .ZN(new_n18721_));
  AOI21_X1   g18424(.A1(new_n18717_), .A2(new_n18721_), .B(new_n18491_), .ZN(new_n18722_));
  XOR2_X1    g18425(.A1(new_n18489_), .A2(new_n18722_), .Z(new_n18723_));
  XOR2_X1    g18426(.A1(new_n18723_), .A2(new_n18485_), .Z(\f[76] ));
  INV_X1     g18427(.I(new_n18722_), .ZN(new_n18725_));
  NAND3_X1   g18428(.A1(new_n18717_), .A2(new_n18491_), .A3(new_n18721_), .ZN(new_n18726_));
  NAND2_X1   g18429(.A1(new_n18726_), .A2(new_n18481_), .ZN(new_n18727_));
  OAI21_X1   g18430(.A1(new_n18489_), .A2(new_n18727_), .B(new_n18725_), .ZN(new_n18728_));
  INV_X1     g18431(.I(new_n18492_), .ZN(new_n18729_));
  AOI21_X1   g18432(.A1(new_n18729_), .A2(new_n18719_), .B(new_n18718_), .ZN(new_n18730_));
  INV_X1     g18433(.I(new_n18730_), .ZN(new_n18731_));
  OAI21_X1   g18434(.A1(new_n18416_), .A2(new_n18495_), .B(new_n18681_), .ZN(new_n18732_));
  AND2_X2    g18435(.A1(new_n18732_), .A2(new_n18679_), .Z(new_n18733_));
  INV_X1     g18436(.I(new_n18658_), .ZN(new_n18734_));
  AOI21_X1   g18437(.A1(new_n18734_), .A2(new_n18499_), .B(new_n18655_), .ZN(new_n18735_));
  OAI22_X1   g18438(.A1(new_n2171_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n2166_), .ZN(new_n18736_));
  OAI21_X1   g18439(.A1(new_n10025_), .A2(new_n2322_), .B(new_n18736_), .ZN(new_n18737_));
  AOI21_X1   g18440(.A1(new_n18737_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n18738_));
  XOR2_X1    g18441(.A1(new_n10476_), .A2(new_n18738_), .Z(new_n18739_));
  OAI22_X1   g18442(.A1(new_n8948_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n9295_), .ZN(new_n18740_));
  OAI21_X1   g18443(.A1(new_n8563_), .A2(new_n2884_), .B(new_n18740_), .ZN(new_n18741_));
  AOI21_X1   g18444(.A1(new_n9299_), .A2(new_n2694_), .B(new_n18741_), .ZN(new_n18742_));
  NAND2_X1   g18445(.A1(new_n18647_), .A2(new_n18504_), .ZN(new_n18743_));
  XOR2_X1    g18446(.A1(new_n18502_), .A2(\a[32] ), .Z(new_n18744_));
  INV_X1     g18447(.I(new_n18744_), .ZN(new_n18745_));
  OAI21_X1   g18448(.A1(new_n18647_), .A2(new_n18504_), .B(new_n18745_), .ZN(new_n18746_));
  NAND2_X1   g18449(.A1(new_n18746_), .A2(new_n18743_), .ZN(new_n18747_));
  INV_X1     g18450(.I(new_n18747_), .ZN(new_n18748_));
  OAI22_X1   g18451(.A1(new_n7870_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n8218_), .ZN(new_n18749_));
  OAI21_X1   g18452(.A1(new_n7864_), .A2(new_n3569_), .B(new_n18749_), .ZN(new_n18750_));
  AOI21_X1   g18453(.A1(new_n18750_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n18751_));
  XOR2_X1    g18454(.A1(new_n8217_), .A2(new_n18751_), .Z(new_n18752_));
  OAI22_X1   g18455(.A1(new_n4072_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n4067_), .ZN(new_n18753_));
  OAI21_X1   g18456(.A1(new_n6538_), .A2(new_n4318_), .B(new_n18753_), .ZN(new_n18754_));
  AOI21_X1   g18457(.A1(new_n18754_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n18755_));
  XNOR2_X1   g18458(.A1(new_n7202_), .A2(new_n18755_), .ZN(new_n18756_));
  NAND2_X1   g18459(.A1(new_n18631_), .A2(new_n18630_), .ZN(new_n18757_));
  NAND2_X1   g18460(.A1(new_n18757_), .A2(new_n18632_), .ZN(new_n18758_));
  OAI22_X1   g18461(.A1(new_n5420_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n5107_), .ZN(new_n18759_));
  OAI21_X1   g18462(.A1(new_n5913_), .A2(new_n5112_), .B(new_n18759_), .ZN(new_n18760_));
  AOI21_X1   g18463(.A1(new_n18760_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n18761_));
  XOR2_X1    g18464(.A1(new_n6233_), .A2(new_n18761_), .Z(new_n18762_));
  OAI22_X1   g18465(.A1(new_n5993_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n5991_), .ZN(new_n18763_));
  OAI21_X1   g18466(.A1(new_n4774_), .A2(new_n5997_), .B(new_n18763_), .ZN(new_n18764_));
  AOI21_X1   g18467(.A1(new_n18764_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n18765_));
  XNOR2_X1   g18468(.A1(new_n5357_), .A2(new_n18765_), .ZN(new_n18766_));
  INV_X1     g18469(.I(new_n18766_), .ZN(new_n18767_));
  OAI22_X1   g18470(.A1(new_n7619_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n8309_), .ZN(new_n18768_));
  OAI21_X1   g18471(.A1(new_n3260_), .A2(new_n7947_), .B(new_n18768_), .ZN(new_n18769_));
  AOI21_X1   g18472(.A1(new_n18769_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n18770_));
  XOR2_X1    g18473(.A1(new_n3722_), .A2(new_n18770_), .Z(new_n18771_));
  INV_X1     g18474(.I(new_n18771_), .ZN(new_n18772_));
  INV_X1     g18475(.I(new_n2440_), .ZN(new_n18773_));
  AOI22_X1   g18476(.A1(new_n11415_), .A2(new_n18773_), .B1(\b[24] ), .B2(new_n10145_), .ZN(new_n18774_));
  OAI21_X1   g18477(.A1(new_n18774_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n18775_));
  XOR2_X1    g18478(.A1(new_n2443_), .A2(new_n18775_), .Z(new_n18776_));
  AOI21_X1   g18479(.A1(new_n18540_), .A2(new_n18577_), .B(new_n18576_), .ZN(new_n18777_));
  AOI22_X1   g18480(.A1(new_n13078_), .A2(\b[18] ), .B1(new_n1527_), .B2(new_n12218_), .ZN(new_n18778_));
  OAI21_X1   g18481(.A1(new_n18778_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n18779_));
  XNOR2_X1   g18482(.A1(new_n1530_), .A2(new_n18779_), .ZN(new_n18780_));
  INV_X1     g18483(.I(new_n18550_), .ZN(new_n18781_));
  AOI21_X1   g18484(.A1(new_n18543_), .A2(new_n18781_), .B(new_n18552_), .ZN(new_n18782_));
  OAI22_X1   g18485(.A1(new_n13880_), .A2(new_n1287_), .B1(new_n1017_), .B2(new_n13885_), .ZN(new_n18783_));
  AOI21_X1   g18486(.A1(new_n18783_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n18784_));
  XOR2_X1    g18487(.A1(new_n1196_), .A2(new_n18784_), .Z(new_n18785_));
  NOR2_X1    g18488(.A1(new_n13476_), .A2(new_n861_), .ZN(new_n18786_));
  XOR2_X1    g18489(.A1(new_n14736_), .A2(new_n861_), .Z(new_n18787_));
  NAND2_X1   g18490(.A1(new_n18787_), .A2(\b[14] ), .ZN(new_n18788_));
  XOR2_X1    g18491(.A1(new_n18788_), .A2(new_n18786_), .Z(new_n18789_));
  XNOR2_X1   g18492(.A1(new_n18549_), .A2(new_n18789_), .ZN(new_n18790_));
  NAND2_X1   g18493(.A1(new_n18785_), .A2(new_n18790_), .ZN(new_n18791_));
  NOR2_X1    g18494(.A1(new_n18556_), .A2(new_n18789_), .ZN(new_n18792_));
  NAND2_X1   g18495(.A1(new_n18556_), .A2(new_n18789_), .ZN(new_n18793_));
  INV_X1     g18496(.I(new_n18793_), .ZN(new_n18794_));
  NOR2_X1    g18497(.A1(new_n18794_), .A2(new_n18792_), .ZN(new_n18795_));
  OAI21_X1   g18498(.A1(new_n18785_), .A2(new_n18795_), .B(new_n18791_), .ZN(new_n18796_));
  NAND2_X1   g18499(.A1(new_n18796_), .A2(new_n18782_), .ZN(new_n18797_));
  NOR2_X1    g18500(.A1(new_n18796_), .A2(new_n18782_), .ZN(new_n18798_));
  INV_X1     g18501(.I(new_n18798_), .ZN(new_n18799_));
  AOI21_X1   g18502(.A1(new_n18797_), .A2(new_n18799_), .B(new_n18780_), .ZN(new_n18800_));
  INV_X1     g18503(.I(new_n18780_), .ZN(new_n18801_));
  XNOR2_X1   g18504(.A1(new_n18796_), .A2(new_n18782_), .ZN(new_n18802_));
  NOR2_X1    g18505(.A1(new_n18801_), .A2(new_n18802_), .ZN(new_n18803_));
  NOR2_X1    g18506(.A1(new_n18803_), .A2(new_n18800_), .ZN(new_n18804_));
  AOI22_X1   g18507(.A1(new_n10969_), .A2(new_n2097_), .B1(new_n11394_), .B2(\b[21] ), .ZN(new_n18805_));
  OAI21_X1   g18508(.A1(new_n18805_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n18806_));
  XOR2_X1    g18509(.A1(new_n1940_), .A2(new_n18806_), .Z(new_n18807_));
  NAND2_X1   g18510(.A1(new_n18568_), .A2(new_n18558_), .ZN(new_n18808_));
  AND2_X2    g18511(.A1(new_n18808_), .A2(new_n18567_), .Z(new_n18809_));
  INV_X1     g18512(.I(new_n18809_), .ZN(new_n18810_));
  XOR2_X1    g18513(.A1(new_n18807_), .A2(new_n18810_), .Z(new_n18811_));
  NOR2_X1    g18514(.A1(new_n18811_), .A2(new_n18804_), .ZN(new_n18812_));
  INV_X1     g18515(.I(new_n18804_), .ZN(new_n18813_));
  OR2_X2     g18516(.A1(new_n18807_), .A2(new_n18809_), .Z(new_n18814_));
  NAND2_X1   g18517(.A1(new_n18807_), .A2(new_n18809_), .ZN(new_n18815_));
  AOI21_X1   g18518(.A1(new_n18814_), .A2(new_n18815_), .B(new_n18813_), .ZN(new_n18816_));
  NOR2_X1    g18519(.A1(new_n18812_), .A2(new_n18816_), .ZN(new_n18817_));
  XOR2_X1    g18520(.A1(new_n18817_), .A2(new_n18777_), .Z(new_n18818_));
  INV_X1     g18521(.I(new_n18777_), .ZN(new_n18819_));
  NOR2_X1    g18522(.A1(new_n18817_), .A2(new_n18819_), .ZN(new_n18820_));
  NAND2_X1   g18523(.A1(new_n18817_), .A2(new_n18819_), .ZN(new_n18821_));
  INV_X1     g18524(.I(new_n18821_), .ZN(new_n18822_));
  OAI21_X1   g18525(.A1(new_n18822_), .A2(new_n18820_), .B(new_n18776_), .ZN(new_n18823_));
  OAI21_X1   g18526(.A1(new_n18818_), .A2(new_n18776_), .B(new_n18823_), .ZN(new_n18824_));
  AOI22_X1   g18527(.A1(new_n8631_), .A2(\b[28] ), .B1(\b[29] ), .B2(new_n9382_), .ZN(new_n18825_));
  AOI21_X1   g18528(.A1(\b[27] ), .A2(new_n9731_), .B(new_n18825_), .ZN(new_n18826_));
  OAI21_X1   g18529(.A1(new_n18826_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n18827_));
  XNOR2_X1   g18530(.A1(new_n3022_), .A2(new_n18827_), .ZN(new_n18828_));
  OAI21_X1   g18531(.A1(new_n18594_), .A2(new_n18592_), .B(new_n18590_), .ZN(new_n18829_));
  XOR2_X1    g18532(.A1(new_n18828_), .A2(new_n18829_), .Z(new_n18830_));
  AND2_X2    g18533(.A1(new_n18828_), .A2(new_n18829_), .Z(new_n18831_));
  NOR2_X1    g18534(.A1(new_n18828_), .A2(new_n18829_), .ZN(new_n18832_));
  NOR2_X1    g18535(.A1(new_n18831_), .A2(new_n18832_), .ZN(new_n18833_));
  NOR2_X1    g18536(.A1(new_n18833_), .A2(new_n18824_), .ZN(new_n18834_));
  AOI21_X1   g18537(.A1(new_n18824_), .A2(new_n18830_), .B(new_n18834_), .ZN(new_n18835_));
  NAND2_X1   g18538(.A1(new_n18603_), .A2(new_n18536_), .ZN(new_n18836_));
  NAND2_X1   g18539(.A1(new_n18836_), .A2(new_n18602_), .ZN(new_n18837_));
  INV_X1     g18540(.I(new_n18837_), .ZN(new_n18838_));
  NOR2_X1    g18541(.A1(new_n18835_), .A2(new_n18838_), .ZN(new_n18839_));
  NAND2_X1   g18542(.A1(new_n18835_), .A2(new_n18838_), .ZN(new_n18840_));
  INV_X1     g18543(.I(new_n18840_), .ZN(new_n18841_));
  OAI21_X1   g18544(.A1(new_n18841_), .A2(new_n18839_), .B(new_n18772_), .ZN(new_n18842_));
  XOR2_X1    g18545(.A1(new_n18835_), .A2(new_n18837_), .Z(new_n18843_));
  OAI21_X1   g18546(.A1(new_n18772_), .A2(new_n18843_), .B(new_n18842_), .ZN(new_n18844_));
  OAI22_X1   g18547(.A1(new_n6644_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n6647_), .ZN(new_n18845_));
  OAI21_X1   g18548(.A1(new_n3989_), .A2(new_n7284_), .B(new_n18845_), .ZN(new_n18846_));
  AOI21_X1   g18549(.A1(new_n18846_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n18847_));
  XOR2_X1    g18550(.A1(new_n4499_), .A2(new_n18847_), .Z(new_n18848_));
  INV_X1     g18551(.I(new_n18848_), .ZN(new_n18849_));
  OAI21_X1   g18552(.A1(new_n18530_), .A2(new_n18608_), .B(new_n18609_), .ZN(new_n18850_));
  AND2_X2    g18553(.A1(new_n18850_), .A2(new_n18849_), .Z(new_n18851_));
  NOR2_X1    g18554(.A1(new_n18850_), .A2(new_n18849_), .ZN(new_n18852_));
  OAI21_X1   g18555(.A1(new_n18851_), .A2(new_n18852_), .B(new_n18844_), .ZN(new_n18853_));
  XOR2_X1    g18556(.A1(new_n18850_), .A2(new_n18848_), .Z(new_n18854_));
  OAI21_X1   g18557(.A1(new_n18844_), .A2(new_n18854_), .B(new_n18853_), .ZN(new_n18855_));
  INV_X1     g18558(.I(new_n18618_), .ZN(new_n18856_));
  OAI21_X1   g18559(.A1(new_n18523_), .A2(new_n18617_), .B(new_n18856_), .ZN(new_n18857_));
  XOR2_X1    g18560(.A1(new_n18857_), .A2(new_n18855_), .Z(new_n18858_));
  NAND2_X1   g18561(.A1(new_n18857_), .A2(new_n18855_), .ZN(new_n18859_));
  OR2_X2     g18562(.A1(new_n18857_), .A2(new_n18855_), .Z(new_n18860_));
  AOI21_X1   g18563(.A1(new_n18860_), .A2(new_n18859_), .B(new_n18767_), .ZN(new_n18861_));
  AOI21_X1   g18564(.A1(new_n18767_), .A2(new_n18858_), .B(new_n18861_), .ZN(new_n18862_));
  NAND2_X1   g18565(.A1(new_n18624_), .A2(new_n18623_), .ZN(new_n18863_));
  NAND2_X1   g18566(.A1(new_n18863_), .A2(new_n18625_), .ZN(new_n18864_));
  XNOR2_X1   g18567(.A1(new_n18862_), .A2(new_n18864_), .ZN(new_n18865_));
  NOR2_X1    g18568(.A1(new_n18865_), .A2(new_n18762_), .ZN(new_n18866_));
  INV_X1     g18569(.I(new_n18762_), .ZN(new_n18867_));
  NAND2_X1   g18570(.A1(new_n18862_), .A2(new_n18864_), .ZN(new_n18868_));
  NOR2_X1    g18571(.A1(new_n18862_), .A2(new_n18864_), .ZN(new_n18869_));
  INV_X1     g18572(.I(new_n18869_), .ZN(new_n18870_));
  AOI21_X1   g18573(.A1(new_n18870_), .A2(new_n18868_), .B(new_n18867_), .ZN(new_n18871_));
  NOR2_X1    g18574(.A1(new_n18866_), .A2(new_n18871_), .ZN(new_n18872_));
  OR2_X2     g18575(.A1(new_n18872_), .A2(new_n18758_), .Z(new_n18873_));
  NAND2_X1   g18576(.A1(new_n18872_), .A2(new_n18758_), .ZN(new_n18874_));
  AOI21_X1   g18577(.A1(new_n18873_), .A2(new_n18874_), .B(new_n18756_), .ZN(new_n18875_));
  INV_X1     g18578(.I(new_n18756_), .ZN(new_n18876_));
  XNOR2_X1   g18579(.A1(new_n18872_), .A2(new_n18758_), .ZN(new_n18877_));
  NOR2_X1    g18580(.A1(new_n18877_), .A2(new_n18876_), .ZN(new_n18878_));
  NOR2_X1    g18581(.A1(new_n18878_), .A2(new_n18875_), .ZN(new_n18879_));
  OAI21_X1   g18582(.A1(new_n18644_), .A2(new_n18642_), .B(new_n18640_), .ZN(new_n18880_));
  INV_X1     g18583(.I(new_n18880_), .ZN(new_n18881_));
  NOR2_X1    g18584(.A1(new_n18879_), .A2(new_n18881_), .ZN(new_n18882_));
  INV_X1     g18585(.I(new_n18882_), .ZN(new_n18883_));
  NAND2_X1   g18586(.A1(new_n18879_), .A2(new_n18881_), .ZN(new_n18884_));
  AOI21_X1   g18587(.A1(new_n18883_), .A2(new_n18884_), .B(new_n18752_), .ZN(new_n18885_));
  INV_X1     g18588(.I(new_n18752_), .ZN(new_n18886_));
  XOR2_X1    g18589(.A1(new_n18879_), .A2(new_n18880_), .Z(new_n18887_));
  NOR2_X1    g18590(.A1(new_n18887_), .A2(new_n18886_), .ZN(new_n18888_));
  NOR2_X1    g18591(.A1(new_n18888_), .A2(new_n18885_), .ZN(new_n18889_));
  XOR2_X1    g18592(.A1(new_n18889_), .A2(new_n18748_), .Z(new_n18890_));
  XOR2_X1    g18593(.A1(new_n18890_), .A2(new_n18742_), .Z(new_n18891_));
  XOR2_X1    g18594(.A1(new_n18891_), .A2(\a[29] ), .Z(new_n18892_));
  OR2_X2     g18595(.A1(new_n18892_), .A2(new_n18739_), .Z(new_n18893_));
  NAND2_X1   g18596(.A1(new_n18892_), .A2(new_n18739_), .ZN(new_n18894_));
  AOI21_X1   g18597(.A1(new_n18893_), .A2(new_n18894_), .B(new_n18735_), .ZN(new_n18895_));
  INV_X1     g18598(.I(new_n18735_), .ZN(new_n18896_));
  XNOR2_X1   g18599(.A1(new_n18892_), .A2(new_n18739_), .ZN(new_n18897_));
  NOR2_X1    g18600(.A1(new_n18897_), .A2(new_n18896_), .ZN(new_n18898_));
  NOR2_X1    g18601(.A1(new_n18898_), .A2(new_n18895_), .ZN(new_n18899_));
  INV_X1     g18602(.I(new_n18667_), .ZN(new_n18900_));
  AOI21_X1   g18603(.A1(new_n18668_), .A2(new_n18665_), .B(new_n18498_), .ZN(new_n18901_));
  NOR2_X1    g18604(.A1(new_n18901_), .A2(new_n18900_), .ZN(new_n18902_));
  NAND2_X1   g18605(.A1(new_n11748_), .A2(new_n1702_), .ZN(new_n18903_));
  AOI22_X1   g18606(.A1(\b[56] ), .A2(new_n2725_), .B1(new_n1702_), .B2(\b[55] ), .ZN(new_n18904_));
  AOI21_X1   g18607(.A1(\b[54] ), .A2(new_n1851_), .B(new_n18904_), .ZN(new_n18905_));
  NAND2_X1   g18608(.A1(new_n18903_), .A2(new_n18905_), .ZN(new_n18906_));
  XOR2_X1    g18609(.A1(new_n18902_), .A2(new_n18906_), .Z(new_n18907_));
  XOR2_X1    g18610(.A1(new_n18907_), .A2(new_n18899_), .Z(new_n18908_));
  XOR2_X1    g18611(.A1(new_n18908_), .A2(\a[23] ), .Z(new_n18909_));
  OAI22_X1   g18612(.A1(new_n1347_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n1344_), .ZN(new_n18910_));
  OAI21_X1   g18613(.A1(new_n12536_), .A2(new_n1457_), .B(new_n18910_), .ZN(new_n18911_));
  AOI21_X1   g18614(.A1(new_n18911_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n18912_));
  XOR2_X1    g18615(.A1(new_n12969_), .A2(new_n18912_), .Z(new_n18913_));
  INV_X1     g18616(.I(new_n18913_), .ZN(new_n18914_));
  NAND2_X1   g18617(.A1(new_n18909_), .A2(new_n18914_), .ZN(new_n18915_));
  XOR2_X1    g18618(.A1(new_n18908_), .A2(new_n1709_), .Z(new_n18916_));
  NAND2_X1   g18619(.A1(new_n18916_), .A2(new_n18913_), .ZN(new_n18917_));
  AOI21_X1   g18620(.A1(new_n18915_), .A2(new_n18917_), .B(new_n18733_), .ZN(new_n18918_));
  INV_X1     g18621(.I(new_n18733_), .ZN(new_n18919_));
  NAND2_X1   g18622(.A1(new_n18916_), .A2(new_n18914_), .ZN(new_n18920_));
  NAND2_X1   g18623(.A1(new_n18909_), .A2(new_n18913_), .ZN(new_n18921_));
  AOI21_X1   g18624(.A1(new_n18921_), .A2(new_n18920_), .B(new_n18919_), .ZN(new_n18922_));
  NOR2_X1    g18625(.A1(new_n18684_), .A2(new_n18686_), .ZN(new_n18923_));
  NAND2_X1   g18626(.A1(new_n18684_), .A2(new_n18686_), .ZN(new_n18924_));
  XOR2_X1    g18627(.A1(new_n18690_), .A2(new_n1346_), .Z(new_n18925_));
  INV_X1     g18628(.I(new_n18925_), .ZN(new_n18926_));
  AOI21_X1   g18629(.A1(new_n18924_), .A2(new_n18926_), .B(new_n18923_), .ZN(new_n18927_));
  OAI22_X1   g18630(.A1(new_n1055_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n1061_), .ZN(new_n18928_));
  OAI21_X1   g18631(.A1(new_n13367_), .A2(new_n1332_), .B(new_n18928_), .ZN(new_n18929_));
  AOI21_X1   g18632(.A1(new_n18183_), .A2(new_n1056_), .B(new_n18929_), .ZN(new_n18930_));
  XNOR2_X1   g18633(.A1(new_n18927_), .A2(new_n18930_), .ZN(new_n18931_));
  NOR3_X1    g18634(.A1(new_n18931_), .A2(new_n18918_), .A3(new_n18922_), .ZN(new_n18932_));
  NOR2_X1    g18635(.A1(new_n18918_), .A2(new_n18922_), .ZN(new_n18933_));
  INV_X1     g18636(.I(new_n18931_), .ZN(new_n18934_));
  NOR2_X1    g18637(.A1(new_n18934_), .A2(new_n18933_), .ZN(new_n18935_));
  OAI21_X1   g18638(.A1(new_n18935_), .A2(new_n18932_), .B(new_n1057_), .ZN(new_n18936_));
  NOR3_X1    g18639(.A1(new_n18935_), .A2(new_n1057_), .A3(new_n18932_), .ZN(new_n18937_));
  INV_X1     g18640(.I(new_n18937_), .ZN(new_n18938_));
  NAND2_X1   g18641(.A1(new_n18938_), .A2(new_n18936_), .ZN(new_n18939_));
  INV_X1     g18642(.I(new_n18939_), .ZN(new_n18940_));
  NOR2_X1    g18643(.A1(new_n18700_), .A2(new_n18697_), .ZN(new_n18941_));
  AOI21_X1   g18644(.A1(new_n18700_), .A2(new_n18697_), .B(new_n18494_), .ZN(new_n18942_));
  NOR2_X1    g18645(.A1(new_n18942_), .A2(new_n18941_), .ZN(new_n18943_));
  AOI21_X1   g18646(.A1(new_n817_), .A2(new_n895_), .B(new_n16486_), .ZN(new_n18944_));
  XOR2_X1    g18647(.A1(new_n18943_), .A2(new_n18944_), .Z(new_n18945_));
  NAND2_X1   g18648(.A1(new_n18940_), .A2(new_n18945_), .ZN(new_n18946_));
  XNOR2_X1   g18649(.A1(new_n18943_), .A2(new_n18944_), .ZN(new_n18947_));
  NAND2_X1   g18650(.A1(new_n18947_), .A2(new_n18939_), .ZN(new_n18948_));
  AOI21_X1   g18651(.A1(new_n18946_), .A2(new_n18948_), .B(\a[14] ), .ZN(new_n18949_));
  NOR2_X1    g18652(.A1(new_n18947_), .A2(new_n18939_), .ZN(new_n18950_));
  NOR2_X1    g18653(.A1(new_n18940_), .A2(new_n18945_), .ZN(new_n18951_));
  NOR3_X1    g18654(.A1(new_n18951_), .A2(new_n18950_), .A3(new_n827_), .ZN(new_n18952_));
  OAI21_X1   g18655(.A1(new_n18952_), .A2(new_n18949_), .B(new_n18731_), .ZN(new_n18953_));
  NOR2_X1    g18656(.A1(new_n18952_), .A2(new_n18949_), .ZN(new_n18954_));
  NAND2_X1   g18657(.A1(new_n18954_), .A2(new_n18730_), .ZN(new_n18955_));
  NAND2_X1   g18658(.A1(new_n18955_), .A2(new_n18953_), .ZN(new_n18956_));
  NAND2_X1   g18659(.A1(new_n18728_), .A2(new_n18956_), .ZN(new_n18957_));
  INV_X1     g18660(.I(new_n17971_), .ZN(new_n18958_));
  NOR3_X1    g18661(.A1(new_n17704_), .A2(new_n17402_), .A3(new_n17403_), .ZN(new_n18959_));
  NOR2_X1    g18662(.A1(new_n17711_), .A2(new_n17131_), .ZN(new_n18960_));
  NOR2_X1    g18663(.A1(new_n18960_), .A2(new_n18959_), .ZN(new_n18961_));
  NAND3_X1   g18664(.A1(new_n17128_), .A2(new_n18961_), .A3(new_n17974_), .ZN(new_n18962_));
  INV_X1     g18665(.I(new_n18211_), .ZN(new_n18963_));
  NAND2_X1   g18666(.A1(new_n18478_), .A2(new_n18480_), .ZN(new_n18964_));
  NAND4_X1   g18667(.A1(new_n18964_), .A2(new_n18963_), .A3(new_n18485_), .A4(new_n18209_), .ZN(new_n18965_));
  AOI22_X1   g18668(.A1(new_n18964_), .A2(new_n18485_), .B1(new_n18963_), .B2(new_n18209_), .ZN(new_n18966_));
  OAI21_X1   g18669(.A1(new_n18966_), .A2(new_n18214_), .B(new_n18965_), .ZN(new_n18967_));
  AOI21_X1   g18670(.A1(new_n18962_), .A2(new_n18958_), .B(new_n18967_), .ZN(new_n18968_));
  INV_X1     g18671(.I(new_n18721_), .ZN(new_n18969_));
  NOR2_X1    g18672(.A1(new_n18969_), .A2(new_n18716_), .ZN(new_n18970_));
  AOI21_X1   g18673(.A1(new_n18970_), .A2(new_n18491_), .B(new_n18485_), .ZN(new_n18971_));
  AOI21_X1   g18674(.A1(new_n18968_), .A2(new_n18971_), .B(new_n18722_), .ZN(new_n18972_));
  XOR2_X1    g18675(.A1(new_n18954_), .A2(new_n18730_), .Z(new_n18973_));
  NAND2_X1   g18676(.A1(new_n18973_), .A2(new_n18972_), .ZN(new_n18974_));
  NAND2_X1   g18677(.A1(new_n18974_), .A2(new_n18957_), .ZN(\f[77] ));
  INV_X1     g18678(.I(new_n18943_), .ZN(new_n18976_));
  NAND2_X1   g18679(.A1(new_n18939_), .A2(new_n18976_), .ZN(new_n18977_));
  XOR2_X1    g18680(.A1(new_n18944_), .A2(\a[14] ), .Z(new_n18978_));
  INV_X1     g18681(.I(new_n18978_), .ZN(new_n18979_));
  OAI21_X1   g18682(.A1(new_n18939_), .A2(new_n18976_), .B(new_n18979_), .ZN(new_n18980_));
  NOR2_X1    g18683(.A1(new_n18933_), .A2(new_n18927_), .ZN(new_n18981_));
  NAND2_X1   g18684(.A1(new_n18933_), .A2(new_n18927_), .ZN(new_n18982_));
  XOR2_X1    g18685(.A1(new_n18930_), .A2(\a[17] ), .Z(new_n18983_));
  INV_X1     g18686(.I(new_n18983_), .ZN(new_n18984_));
  AOI21_X1   g18687(.A1(new_n18982_), .A2(new_n18984_), .B(new_n18981_), .ZN(new_n18985_));
  NOR2_X1    g18688(.A1(new_n18916_), .A2(new_n18913_), .ZN(new_n18986_));
  AOI21_X1   g18689(.A1(new_n18919_), .A2(new_n18917_), .B(new_n18986_), .ZN(new_n18987_));
  NAND2_X1   g18690(.A1(new_n18899_), .A2(new_n18902_), .ZN(new_n18988_));
  XOR2_X1    g18691(.A1(new_n18906_), .A2(new_n1709_), .Z(new_n18989_));
  NAND2_X1   g18692(.A1(new_n18988_), .A2(new_n18989_), .ZN(new_n18990_));
  OAI21_X1   g18693(.A1(new_n18899_), .A2(new_n18902_), .B(new_n18990_), .ZN(new_n18991_));
  NAND2_X1   g18694(.A1(new_n18894_), .A2(new_n18896_), .ZN(new_n18992_));
  OAI22_X1   g18695(.A1(new_n2171_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n2166_), .ZN(new_n18993_));
  OAI21_X1   g18696(.A1(new_n10031_), .A2(new_n2322_), .B(new_n18993_), .ZN(new_n18994_));
  AOI21_X1   g18697(.A1(new_n18994_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n18995_));
  XNOR2_X1   g18698(.A1(new_n10866_), .A2(new_n18995_), .ZN(new_n18996_));
  OAI21_X1   g18699(.A1(new_n18888_), .A2(new_n18885_), .B(new_n18747_), .ZN(new_n18997_));
  NAND2_X1   g18700(.A1(new_n18889_), .A2(new_n18748_), .ZN(new_n18998_));
  XOR2_X1    g18701(.A1(new_n18742_), .A2(new_n2702_), .Z(new_n18999_));
  NAND2_X1   g18702(.A1(new_n18998_), .A2(new_n18999_), .ZN(new_n19000_));
  NAND2_X1   g18703(.A1(new_n19000_), .A2(new_n18997_), .ZN(new_n19001_));
  OAI22_X1   g18704(.A1(new_n9295_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n10025_), .ZN(new_n19002_));
  OAI21_X1   g18705(.A1(new_n8948_), .A2(new_n2884_), .B(new_n19002_), .ZN(new_n19003_));
  AOI21_X1   g18706(.A1(new_n19003_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n19004_));
  XNOR2_X1   g18707(.A1(new_n9642_), .A2(new_n19004_), .ZN(new_n19005_));
  NAND2_X1   g18708(.A1(new_n18873_), .A2(new_n18876_), .ZN(new_n19006_));
  NAND2_X1   g18709(.A1(new_n19006_), .A2(new_n18874_), .ZN(new_n19007_));
  OAI21_X1   g18710(.A1(new_n18762_), .A2(new_n18869_), .B(new_n18868_), .ZN(new_n19008_));
  INV_X1     g18711(.I(new_n19008_), .ZN(new_n19009_));
  NAND2_X1   g18712(.A1(new_n18860_), .A2(new_n18767_), .ZN(new_n19010_));
  AND2_X2    g18713(.A1(new_n19010_), .A2(new_n18859_), .Z(new_n19011_));
  INV_X1     g18714(.I(new_n19011_), .ZN(new_n19012_));
  INV_X1     g18715(.I(new_n18852_), .ZN(new_n19013_));
  AOI21_X1   g18716(.A1(new_n18844_), .A2(new_n19013_), .B(new_n18851_), .ZN(new_n19014_));
  AOI21_X1   g18717(.A1(new_n18772_), .A2(new_n18840_), .B(new_n18839_), .ZN(new_n19015_));
  OAI21_X1   g18718(.A1(new_n18776_), .A2(new_n18820_), .B(new_n18821_), .ZN(new_n19016_));
  NAND2_X1   g18719(.A1(new_n18813_), .A2(new_n18815_), .ZN(new_n19017_));
  AOI21_X1   g18720(.A1(new_n18801_), .A2(new_n18797_), .B(new_n18798_), .ZN(new_n19018_));
  INV_X1     g18721(.I(new_n19018_), .ZN(new_n19019_));
  OAI22_X1   g18722(.A1(new_n13880_), .A2(new_n1295_), .B1(new_n1109_), .B2(new_n13885_), .ZN(new_n19020_));
  AOI21_X1   g18723(.A1(new_n19020_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n19021_));
  XOR2_X1    g18724(.A1(new_n1299_), .A2(new_n19021_), .Z(new_n19022_));
  AOI21_X1   g18725(.A1(new_n18785_), .A2(new_n18793_), .B(new_n18792_), .ZN(new_n19023_));
  NOR2_X1    g18726(.A1(new_n13476_), .A2(new_n930_), .ZN(new_n19024_));
  XOR2_X1    g18727(.A1(new_n14736_), .A2(new_n930_), .Z(new_n19025_));
  NAND2_X1   g18728(.A1(new_n19025_), .A2(\b[15] ), .ZN(new_n19026_));
  XOR2_X1    g18729(.A1(new_n19026_), .A2(new_n19024_), .Z(new_n19027_));
  NOR2_X1    g18730(.A1(new_n19027_), .A2(new_n827_), .ZN(new_n19028_));
  INV_X1     g18731(.I(new_n19028_), .ZN(new_n19029_));
  NAND2_X1   g18732(.A1(new_n19027_), .A2(new_n827_), .ZN(new_n19030_));
  AOI21_X1   g18733(.A1(new_n19029_), .A2(new_n19030_), .B(new_n18549_), .ZN(new_n19031_));
  XOR2_X1    g18734(.A1(new_n19027_), .A2(\a[14] ), .Z(new_n19032_));
  NOR2_X1    g18735(.A1(new_n19032_), .A2(new_n18556_), .ZN(new_n19033_));
  NOR2_X1    g18736(.A1(new_n19033_), .A2(new_n19031_), .ZN(new_n19034_));
  INV_X1     g18737(.I(new_n19034_), .ZN(new_n19035_));
  XOR2_X1    g18738(.A1(new_n19023_), .A2(new_n19035_), .Z(new_n19036_));
  NOR2_X1    g18739(.A1(new_n19036_), .A2(new_n19022_), .ZN(new_n19037_));
  XNOR2_X1   g18740(.A1(new_n1299_), .A2(new_n19021_), .ZN(new_n19038_));
  OR2_X2     g18741(.A1(new_n19023_), .A2(new_n19034_), .Z(new_n19039_));
  NAND2_X1   g18742(.A1(new_n19023_), .A2(new_n19034_), .ZN(new_n19040_));
  AOI21_X1   g18743(.A1(new_n19040_), .A2(new_n19039_), .B(new_n19038_), .ZN(new_n19041_));
  NOR2_X1    g18744(.A1(new_n19037_), .A2(new_n19041_), .ZN(new_n19042_));
  AOI22_X1   g18745(.A1(new_n13078_), .A2(\b[19] ), .B1(new_n1797_), .B2(new_n12218_), .ZN(new_n19043_));
  OAI21_X1   g18746(.A1(new_n19043_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n19044_));
  XNOR2_X1   g18747(.A1(new_n1638_), .A2(new_n19044_), .ZN(new_n19045_));
  XOR2_X1    g18748(.A1(new_n19042_), .A2(new_n19045_), .Z(new_n19046_));
  NAND2_X1   g18749(.A1(new_n19046_), .A2(new_n19019_), .ZN(new_n19047_));
  NAND2_X1   g18750(.A1(new_n19042_), .A2(new_n19045_), .ZN(new_n19048_));
  INV_X1     g18751(.I(new_n19048_), .ZN(new_n19049_));
  NOR2_X1    g18752(.A1(new_n19042_), .A2(new_n19045_), .ZN(new_n19050_));
  OAI21_X1   g18753(.A1(new_n19049_), .A2(new_n19050_), .B(new_n19018_), .ZN(new_n19051_));
  AOI22_X1   g18754(.A1(new_n10969_), .A2(new_n18260_), .B1(new_n11394_), .B2(\b[22] ), .ZN(new_n19052_));
  OAI21_X1   g18755(.A1(new_n19052_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n19053_));
  XOR2_X1    g18756(.A1(new_n2106_), .A2(new_n19053_), .Z(new_n19054_));
  NAND3_X1   g18757(.A1(new_n19054_), .A2(new_n19047_), .A3(new_n19051_), .ZN(new_n19055_));
  NAND2_X1   g18758(.A1(new_n19047_), .A2(new_n19051_), .ZN(new_n19056_));
  INV_X1     g18759(.I(new_n19054_), .ZN(new_n19057_));
  NAND2_X1   g18760(.A1(new_n19057_), .A2(new_n19056_), .ZN(new_n19058_));
  AOI22_X1   g18761(.A1(new_n19058_), .A2(new_n19055_), .B1(new_n18814_), .B2(new_n19017_), .ZN(new_n19059_));
  NAND2_X1   g18762(.A1(new_n19017_), .A2(new_n18814_), .ZN(new_n19060_));
  XOR2_X1    g18763(.A1(new_n19056_), .A2(new_n19054_), .Z(new_n19061_));
  NOR2_X1    g18764(.A1(new_n19061_), .A2(new_n19060_), .ZN(new_n19062_));
  NOR2_X1    g18765(.A1(new_n19062_), .A2(new_n19059_), .ZN(new_n19063_));
  AOI22_X1   g18766(.A1(new_n11415_), .A2(new_n2838_), .B1(\b[25] ), .B2(new_n10145_), .ZN(new_n19064_));
  OAI21_X1   g18767(.A1(new_n19064_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n19065_));
  XOR2_X1    g18768(.A1(new_n2647_), .A2(new_n19065_), .Z(new_n19066_));
  XOR2_X1    g18769(.A1(new_n19063_), .A2(new_n19066_), .Z(new_n19067_));
  AND2_X2    g18770(.A1(new_n19067_), .A2(new_n19016_), .Z(new_n19068_));
  OR2_X2     g18771(.A1(new_n19063_), .A2(new_n19066_), .Z(new_n19069_));
  NAND2_X1   g18772(.A1(new_n19063_), .A2(new_n19066_), .ZN(new_n19070_));
  AOI21_X1   g18773(.A1(new_n19069_), .A2(new_n19070_), .B(new_n19016_), .ZN(new_n19071_));
  NOR2_X1    g18774(.A1(new_n19068_), .A2(new_n19071_), .ZN(new_n19072_));
  OAI22_X1   g18775(.A1(new_n8644_), .A2(new_n3018_), .B1(new_n3260_), .B2(new_n9388_), .ZN(new_n19073_));
  OAI21_X1   g18776(.A1(new_n2842_), .A2(new_n10154_), .B(new_n19073_), .ZN(new_n19074_));
  AOI21_X1   g18777(.A1(new_n19074_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n19075_));
  XOR2_X1    g18778(.A1(new_n3264_), .A2(new_n19075_), .Z(new_n19076_));
  INV_X1     g18779(.I(new_n19076_), .ZN(new_n19077_));
  NOR2_X1    g18780(.A1(new_n18824_), .A2(new_n18832_), .ZN(new_n19078_));
  NOR2_X1    g18781(.A1(new_n19078_), .A2(new_n18831_), .ZN(new_n19079_));
  NOR2_X1    g18782(.A1(new_n19079_), .A2(new_n19077_), .ZN(new_n19080_));
  INV_X1     g18783(.I(new_n19080_), .ZN(new_n19081_));
  NAND2_X1   g18784(.A1(new_n19079_), .A2(new_n19077_), .ZN(new_n19082_));
  AOI21_X1   g18785(.A1(new_n19081_), .A2(new_n19082_), .B(new_n19072_), .ZN(new_n19083_));
  XOR2_X1    g18786(.A1(new_n19079_), .A2(new_n19076_), .Z(new_n19084_));
  NOR3_X1    g18787(.A1(new_n19084_), .A2(new_n19068_), .A3(new_n19071_), .ZN(new_n19085_));
  NOR2_X1    g18788(.A1(new_n19085_), .A2(new_n19083_), .ZN(new_n19086_));
  OAI22_X1   g18789(.A1(new_n7619_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n8309_), .ZN(new_n19087_));
  OAI21_X1   g18790(.A1(new_n3709_), .A2(new_n7947_), .B(new_n19087_), .ZN(new_n19088_));
  AOI21_X1   g18791(.A1(new_n19088_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n19089_));
  XNOR2_X1   g18792(.A1(new_n3993_), .A2(new_n19089_), .ZN(new_n19090_));
  INV_X1     g18793(.I(new_n19090_), .ZN(new_n19091_));
  NAND2_X1   g18794(.A1(new_n19086_), .A2(new_n19091_), .ZN(new_n19092_));
  OAI21_X1   g18795(.A1(new_n19085_), .A2(new_n19083_), .B(new_n19090_), .ZN(new_n19093_));
  AOI21_X1   g18796(.A1(new_n19092_), .A2(new_n19093_), .B(new_n19015_), .ZN(new_n19094_));
  INV_X1     g18797(.I(new_n19015_), .ZN(new_n19095_));
  XOR2_X1    g18798(.A1(new_n19086_), .A2(new_n19090_), .Z(new_n19096_));
  NOR2_X1    g18799(.A1(new_n19096_), .A2(new_n19095_), .ZN(new_n19097_));
  NOR2_X1    g18800(.A1(new_n19097_), .A2(new_n19094_), .ZN(new_n19098_));
  OAI22_X1   g18801(.A1(new_n6644_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n6647_), .ZN(new_n19099_));
  OAI21_X1   g18802(.A1(new_n4253_), .A2(new_n7284_), .B(new_n19099_), .ZN(new_n19100_));
  AOI21_X1   g18803(.A1(new_n19100_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n19101_));
  XNOR2_X1   g18804(.A1(new_n4778_), .A2(new_n19101_), .ZN(new_n19102_));
  INV_X1     g18805(.I(new_n19102_), .ZN(new_n19103_));
  XOR2_X1    g18806(.A1(new_n19098_), .A2(new_n19103_), .Z(new_n19104_));
  NOR2_X1    g18807(.A1(new_n19104_), .A2(new_n19014_), .ZN(new_n19105_));
  INV_X1     g18808(.I(new_n19014_), .ZN(new_n19106_));
  OAI21_X1   g18809(.A1(new_n19097_), .A2(new_n19094_), .B(new_n19103_), .ZN(new_n19107_));
  NAND2_X1   g18810(.A1(new_n19098_), .A2(new_n19102_), .ZN(new_n19108_));
  AOI21_X1   g18811(.A1(new_n19108_), .A2(new_n19107_), .B(new_n19106_), .ZN(new_n19109_));
  NOR2_X1    g18812(.A1(new_n19105_), .A2(new_n19109_), .ZN(new_n19110_));
  OAI22_X1   g18813(.A1(new_n5993_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n5991_), .ZN(new_n19111_));
  OAI21_X1   g18814(.A1(new_n5068_), .A2(new_n5997_), .B(new_n19111_), .ZN(new_n19112_));
  AOI21_X1   g18815(.A1(new_n19112_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n19113_));
  XNOR2_X1   g18816(.A1(new_n5600_), .A2(new_n19113_), .ZN(new_n19114_));
  INV_X1     g18817(.I(new_n19114_), .ZN(new_n19115_));
  NAND2_X1   g18818(.A1(new_n19110_), .A2(new_n19115_), .ZN(new_n19116_));
  INV_X1     g18819(.I(new_n19116_), .ZN(new_n19117_));
  NOR2_X1    g18820(.A1(new_n19110_), .A2(new_n19115_), .ZN(new_n19118_));
  OAI21_X1   g18821(.A1(new_n19117_), .A2(new_n19118_), .B(new_n19012_), .ZN(new_n19119_));
  XOR2_X1    g18822(.A1(new_n19110_), .A2(new_n19115_), .Z(new_n19120_));
  NAND2_X1   g18823(.A1(new_n19120_), .A2(new_n19011_), .ZN(new_n19121_));
  NAND2_X1   g18824(.A1(new_n19121_), .A2(new_n19119_), .ZN(new_n19122_));
  OAI22_X1   g18825(.A1(new_n5420_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n5107_), .ZN(new_n19123_));
  OAI21_X1   g18826(.A1(new_n5921_), .A2(new_n5112_), .B(new_n19123_), .ZN(new_n19124_));
  AOI21_X1   g18827(.A1(new_n19124_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n19125_));
  XOR2_X1    g18828(.A1(new_n6543_), .A2(new_n19125_), .Z(new_n19126_));
  XOR2_X1    g18829(.A1(new_n19122_), .A2(new_n19126_), .Z(new_n19127_));
  NOR2_X1    g18830(.A1(new_n19127_), .A2(new_n19009_), .ZN(new_n19128_));
  INV_X1     g18831(.I(new_n19126_), .ZN(new_n19129_));
  NAND2_X1   g18832(.A1(new_n19122_), .A2(new_n19129_), .ZN(new_n19130_));
  NAND3_X1   g18833(.A1(new_n19121_), .A2(new_n19119_), .A3(new_n19126_), .ZN(new_n19131_));
  AOI21_X1   g18834(.A1(new_n19130_), .A2(new_n19131_), .B(new_n19008_), .ZN(new_n19132_));
  NOR2_X1    g18835(.A1(new_n19128_), .A2(new_n19132_), .ZN(new_n19133_));
  OAI22_X1   g18836(.A1(new_n4072_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n4067_), .ZN(new_n19134_));
  OAI21_X1   g18837(.A1(new_n6847_), .A2(new_n4318_), .B(new_n19134_), .ZN(new_n19135_));
  AOI21_X1   g18838(.A1(new_n19135_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n19136_));
  XOR2_X1    g18839(.A1(new_n7516_), .A2(new_n19136_), .Z(new_n19137_));
  INV_X1     g18840(.I(new_n19137_), .ZN(new_n19138_));
  XOR2_X1    g18841(.A1(new_n19133_), .A2(new_n19138_), .Z(new_n19139_));
  INV_X1     g18842(.I(new_n19133_), .ZN(new_n19140_));
  NOR2_X1    g18843(.A1(new_n19140_), .A2(new_n19137_), .ZN(new_n19141_));
  INV_X1     g18844(.I(new_n19141_), .ZN(new_n19142_));
  NAND2_X1   g18845(.A1(new_n19140_), .A2(new_n19137_), .ZN(new_n19143_));
  AOI21_X1   g18846(.A1(new_n19143_), .A2(new_n19142_), .B(new_n19007_), .ZN(new_n19144_));
  AOI21_X1   g18847(.A1(new_n19007_), .A2(new_n19139_), .B(new_n19144_), .ZN(new_n19145_));
  AOI21_X1   g18848(.A1(new_n18879_), .A2(new_n18881_), .B(new_n18752_), .ZN(new_n19146_));
  NOR2_X1    g18849(.A1(new_n19146_), .A2(new_n18882_), .ZN(new_n19147_));
  OAI22_X1   g18850(.A1(new_n8218_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n8563_), .ZN(new_n19148_));
  OAI21_X1   g18851(.A1(new_n7870_), .A2(new_n3569_), .B(new_n19148_), .ZN(new_n19149_));
  AOI21_X1   g18852(.A1(new_n19149_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n19150_));
  XOR2_X1    g18853(.A1(new_n8568_), .A2(new_n19150_), .Z(new_n19151_));
  NOR2_X1    g18854(.A1(new_n19147_), .A2(new_n19151_), .ZN(new_n19152_));
  INV_X1     g18855(.I(new_n19147_), .ZN(new_n19153_));
  INV_X1     g18856(.I(new_n19151_), .ZN(new_n19154_));
  NOR2_X1    g18857(.A1(new_n19153_), .A2(new_n19154_), .ZN(new_n19155_));
  NOR2_X1    g18858(.A1(new_n19155_), .A2(new_n19152_), .ZN(new_n19156_));
  XOR2_X1    g18859(.A1(new_n19147_), .A2(new_n19151_), .Z(new_n19157_));
  NAND2_X1   g18860(.A1(new_n19145_), .A2(new_n19157_), .ZN(new_n19158_));
  OAI21_X1   g18861(.A1(new_n19145_), .A2(new_n19156_), .B(new_n19158_), .ZN(new_n19159_));
  NAND2_X1   g18862(.A1(new_n19159_), .A2(new_n19005_), .ZN(new_n19160_));
  OR2_X2     g18863(.A1(new_n19159_), .A2(new_n19005_), .Z(new_n19161_));
  NAND2_X1   g18864(.A1(new_n19161_), .A2(new_n19160_), .ZN(new_n19162_));
  XNOR2_X1   g18865(.A1(new_n19159_), .A2(new_n19005_), .ZN(new_n19163_));
  NOR2_X1    g18866(.A1(new_n19163_), .A2(new_n19001_), .ZN(new_n19164_));
  AOI21_X1   g18867(.A1(new_n19001_), .A2(new_n19162_), .B(new_n19164_), .ZN(new_n19165_));
  XNOR2_X1   g18868(.A1(new_n19165_), .A2(new_n18996_), .ZN(new_n19166_));
  AOI21_X1   g18869(.A1(new_n18893_), .A2(new_n18992_), .B(new_n19166_), .ZN(new_n19167_));
  NAND2_X1   g18870(.A1(new_n18992_), .A2(new_n18893_), .ZN(new_n19168_));
  NOR2_X1    g18871(.A1(new_n19165_), .A2(new_n18996_), .ZN(new_n19169_));
  INV_X1     g18872(.I(new_n19169_), .ZN(new_n19170_));
  NAND2_X1   g18873(.A1(new_n19165_), .A2(new_n18996_), .ZN(new_n19171_));
  AOI21_X1   g18874(.A1(new_n19170_), .A2(new_n19171_), .B(new_n19168_), .ZN(new_n19172_));
  OAI22_X1   g18875(.A1(new_n1712_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n1707_), .ZN(new_n19173_));
  OAI21_X1   g18876(.A1(new_n11738_), .A2(new_n1850_), .B(new_n19173_), .ZN(new_n19174_));
  AOI21_X1   g18877(.A1(new_n19174_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n19175_));
  XNOR2_X1   g18878(.A1(new_n12128_), .A2(new_n19175_), .ZN(new_n19176_));
  NOR3_X1    g18879(.A1(new_n19167_), .A2(new_n19172_), .A3(new_n19176_), .ZN(new_n19177_));
  NOR2_X1    g18880(.A1(new_n19167_), .A2(new_n19172_), .ZN(new_n19178_));
  INV_X1     g18881(.I(new_n19176_), .ZN(new_n19179_));
  NOR2_X1    g18882(.A1(new_n19178_), .A2(new_n19179_), .ZN(new_n19180_));
  OAI21_X1   g18883(.A1(new_n19177_), .A2(new_n19180_), .B(new_n18991_), .ZN(new_n19181_));
  XOR2_X1    g18884(.A1(new_n19178_), .A2(new_n19176_), .Z(new_n19182_));
  OAI21_X1   g18885(.A1(new_n18991_), .A2(new_n19182_), .B(new_n19181_), .ZN(new_n19183_));
  OAI22_X1   g18886(.A1(new_n1347_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n1344_), .ZN(new_n19184_));
  OAI21_X1   g18887(.A1(new_n12542_), .A2(new_n1457_), .B(new_n19184_), .ZN(new_n19185_));
  AOI21_X1   g18888(.A1(new_n19185_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n19186_));
  XNOR2_X1   g18889(.A1(new_n13371_), .A2(new_n19186_), .ZN(new_n19187_));
  XOR2_X1    g18890(.A1(new_n19183_), .A2(new_n19187_), .Z(new_n19188_));
  INV_X1     g18891(.I(new_n19183_), .ZN(new_n19189_));
  NOR2_X1    g18892(.A1(new_n19189_), .A2(new_n19187_), .ZN(new_n19190_));
  NAND2_X1   g18893(.A1(new_n19189_), .A2(new_n19187_), .ZN(new_n19191_));
  INV_X1     g18894(.I(new_n19191_), .ZN(new_n19192_));
  OAI21_X1   g18895(.A1(new_n19192_), .A2(new_n19190_), .B(new_n18987_), .ZN(new_n19193_));
  OAI21_X1   g18896(.A1(new_n18987_), .A2(new_n19188_), .B(new_n19193_), .ZN(new_n19194_));
  OAI22_X1   g18897(.A1(new_n1055_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n1061_), .ZN(new_n19195_));
  OAI21_X1   g18898(.A1(new_n13785_), .A2(new_n1332_), .B(new_n19195_), .ZN(new_n19196_));
  AOI21_X1   g18899(.A1(new_n19196_), .A2(new_n1057_), .B(new_n1055_), .ZN(new_n19197_));
  XNOR2_X1   g18900(.A1(new_n14599_), .A2(new_n19197_), .ZN(new_n19198_));
  NOR2_X1    g18901(.A1(new_n19194_), .A2(new_n19198_), .ZN(new_n19199_));
  NOR2_X1    g18902(.A1(new_n19188_), .A2(new_n18987_), .ZN(new_n19200_));
  INV_X1     g18903(.I(new_n19190_), .ZN(new_n19201_));
  NAND2_X1   g18904(.A1(new_n19201_), .A2(new_n19191_), .ZN(new_n19202_));
  AOI21_X1   g18905(.A1(new_n18987_), .A2(new_n19202_), .B(new_n19200_), .ZN(new_n19203_));
  INV_X1     g18906(.I(new_n19198_), .ZN(new_n19204_));
  NOR2_X1    g18907(.A1(new_n19203_), .A2(new_n19204_), .ZN(new_n19205_));
  NOR2_X1    g18908(.A1(new_n19199_), .A2(new_n19205_), .ZN(new_n19206_));
  NOR2_X1    g18909(.A1(new_n19203_), .A2(new_n19198_), .ZN(new_n19207_));
  NOR2_X1    g18910(.A1(new_n19194_), .A2(new_n19204_), .ZN(new_n19208_));
  OAI21_X1   g18911(.A1(new_n19208_), .A2(new_n19207_), .B(new_n18985_), .ZN(new_n19209_));
  OAI21_X1   g18912(.A1(new_n18985_), .A2(new_n19206_), .B(new_n19209_), .ZN(new_n19210_));
  NAND3_X1   g18913(.A1(new_n19210_), .A2(new_n18980_), .A3(new_n18977_), .ZN(new_n19211_));
  INV_X1     g18914(.I(new_n19211_), .ZN(new_n19212_));
  AOI21_X1   g18915(.A1(new_n18980_), .A2(new_n18977_), .B(new_n19210_), .ZN(new_n19213_));
  OAI21_X1   g18916(.A1(new_n19212_), .A2(new_n19213_), .B(new_n18973_), .ZN(new_n19214_));
  XOR2_X1    g18917(.A1(new_n19214_), .A2(new_n18953_), .Z(new_n19215_));
  XOR2_X1    g18918(.A1(new_n19215_), .A2(new_n18728_), .Z(\f[78] ));
  NAND2_X1   g18919(.A1(new_n18980_), .A2(new_n18977_), .ZN(new_n19217_));
  OR2_X2     g18920(.A1(new_n19217_), .A2(new_n19210_), .Z(new_n19218_));
  NOR4_X1    g18921(.A1(new_n19212_), .A2(new_n18949_), .A3(new_n18952_), .A4(new_n19213_), .ZN(new_n19219_));
  OAI22_X1   g18922(.A1(new_n19212_), .A2(new_n19213_), .B1(new_n18952_), .B2(new_n18949_), .ZN(new_n19220_));
  AOI21_X1   g18923(.A1(new_n18730_), .A2(new_n19220_), .B(new_n19219_), .ZN(new_n19221_));
  NAND2_X1   g18924(.A1(new_n18728_), .A2(new_n19221_), .ZN(new_n19222_));
  NOR2_X1    g18925(.A1(new_n19205_), .A2(new_n18985_), .ZN(new_n19223_));
  NOR2_X1    g18926(.A1(new_n19223_), .A2(new_n19199_), .ZN(new_n19224_));
  OAI21_X1   g18927(.A1(new_n18987_), .A2(new_n19192_), .B(new_n19201_), .ZN(new_n19225_));
  INV_X1     g18928(.I(new_n19180_), .ZN(new_n19226_));
  AOI21_X1   g18929(.A1(new_n18991_), .A2(new_n19226_), .B(new_n19177_), .ZN(new_n19227_));
  INV_X1     g18930(.I(new_n19227_), .ZN(new_n19228_));
  OAI22_X1   g18931(.A1(new_n1712_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n1707_), .ZN(new_n19229_));
  OAI21_X1   g18932(.A1(new_n11744_), .A2(new_n1850_), .B(new_n19229_), .ZN(new_n19230_));
  AOI21_X1   g18933(.A1(new_n12546_), .A2(new_n1702_), .B(new_n19230_), .ZN(new_n19231_));
  AOI21_X1   g18934(.A1(new_n19168_), .A2(new_n19171_), .B(new_n19169_), .ZN(new_n19232_));
  INV_X1     g18935(.I(new_n19232_), .ZN(new_n19233_));
  OAI22_X1   g18936(.A1(new_n2171_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n2166_), .ZN(new_n19234_));
  OAI21_X1   g18937(.A1(new_n10477_), .A2(new_n2322_), .B(new_n19234_), .ZN(new_n19235_));
  AOI21_X1   g18938(.A1(new_n19235_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n19236_));
  XOR2_X1    g18939(.A1(new_n11298_), .A2(new_n19236_), .Z(new_n19237_));
  INV_X1     g18940(.I(new_n19237_), .ZN(new_n19238_));
  NAND2_X1   g18941(.A1(new_n19160_), .A2(new_n19001_), .ZN(new_n19239_));
  AND2_X2    g18942(.A1(new_n19239_), .A2(new_n19161_), .Z(new_n19240_));
  INV_X1     g18943(.I(new_n19155_), .ZN(new_n19241_));
  AOI21_X1   g18944(.A1(new_n19145_), .A2(new_n19241_), .B(new_n19152_), .ZN(new_n19242_));
  NAND2_X1   g18945(.A1(new_n10035_), .A2(new_n2694_), .ZN(new_n19243_));
  AOI22_X1   g18946(.A1(new_n2694_), .A2(\b[51] ), .B1(\b[52] ), .B2(new_n2699_), .ZN(new_n19244_));
  AOI21_X1   g18947(.A1(\b[50] ), .A2(new_n4094_), .B(new_n19244_), .ZN(new_n19245_));
  NAND2_X1   g18948(.A1(new_n19243_), .A2(new_n19245_), .ZN(new_n19246_));
  OAI22_X1   g18949(.A1(new_n8563_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n8948_), .ZN(new_n19247_));
  OAI21_X1   g18950(.A1(new_n8218_), .A2(new_n3569_), .B(new_n19247_), .ZN(new_n19248_));
  AOI21_X1   g18951(.A1(new_n19248_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n19249_));
  XOR2_X1    g18952(.A1(new_n8952_), .A2(new_n19249_), .Z(new_n19250_));
  INV_X1     g18953(.I(new_n19250_), .ZN(new_n19251_));
  AOI21_X1   g18954(.A1(new_n19007_), .A2(new_n19143_), .B(new_n19141_), .ZN(new_n19252_));
  OAI22_X1   g18955(.A1(new_n4072_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n4067_), .ZN(new_n19253_));
  OAI21_X1   g18956(.A1(new_n7198_), .A2(new_n4318_), .B(new_n19253_), .ZN(new_n19254_));
  AOI21_X1   g18957(.A1(new_n19254_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n19255_));
  XNOR2_X1   g18958(.A1(new_n7874_), .A2(new_n19255_), .ZN(new_n19256_));
  INV_X1     g18959(.I(new_n19256_), .ZN(new_n19257_));
  OAI21_X1   g18960(.A1(new_n19011_), .A2(new_n19118_), .B(new_n19116_), .ZN(new_n19258_));
  INV_X1     g18961(.I(new_n19258_), .ZN(new_n19259_));
  OAI22_X1   g18962(.A1(new_n5993_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n5991_), .ZN(new_n19260_));
  OAI21_X1   g18963(.A1(new_n5353_), .A2(new_n5997_), .B(new_n19260_), .ZN(new_n19261_));
  AOI21_X1   g18964(.A1(new_n19261_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n19262_));
  XOR2_X1    g18965(.A1(new_n5926_), .A2(new_n19262_), .Z(new_n19263_));
  INV_X1     g18966(.I(new_n19263_), .ZN(new_n19264_));
  NAND2_X1   g18967(.A1(new_n19108_), .A2(new_n19106_), .ZN(new_n19265_));
  NAND2_X1   g18968(.A1(new_n19265_), .A2(new_n19107_), .ZN(new_n19266_));
  OAI22_X1   g18969(.A1(new_n6644_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n6647_), .ZN(new_n19267_));
  OAI21_X1   g18970(.A1(new_n4500_), .A2(new_n7284_), .B(new_n19267_), .ZN(new_n19268_));
  AOI21_X1   g18971(.A1(new_n19268_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n19269_));
  XOR2_X1    g18972(.A1(new_n5067_), .A2(new_n19269_), .Z(new_n19270_));
  INV_X1     g18973(.I(new_n19270_), .ZN(new_n19271_));
  NAND2_X1   g18974(.A1(new_n19093_), .A2(new_n19095_), .ZN(new_n19272_));
  AND2_X2    g18975(.A1(new_n19272_), .A2(new_n19092_), .Z(new_n19273_));
  OAI22_X1   g18976(.A1(new_n7619_), .A2(new_n3989_), .B1(new_n4253_), .B2(new_n8309_), .ZN(new_n19274_));
  OAI21_X1   g18977(.A1(new_n3717_), .A2(new_n7947_), .B(new_n19274_), .ZN(new_n19275_));
  AOI21_X1   g18978(.A1(new_n19275_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n19276_));
  XNOR2_X1   g18979(.A1(new_n4257_), .A2(new_n19276_), .ZN(new_n19277_));
  INV_X1     g18980(.I(new_n2843_), .ZN(new_n19278_));
  AOI22_X1   g18981(.A1(new_n11415_), .A2(new_n19278_), .B1(\b[26] ), .B2(new_n10145_), .ZN(new_n19279_));
  OAI21_X1   g18982(.A1(new_n19279_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n19280_));
  XNOR2_X1   g18983(.A1(new_n2846_), .A2(new_n19280_), .ZN(new_n19281_));
  INV_X1     g18984(.I(new_n19281_), .ZN(new_n19282_));
  INV_X1     g18985(.I(new_n19055_), .ZN(new_n19283_));
  AOI22_X1   g18986(.A1(new_n19057_), .A2(new_n19056_), .B1(new_n18814_), .B2(new_n19017_), .ZN(new_n19284_));
  NOR2_X1    g18987(.A1(new_n19284_), .A2(new_n19283_), .ZN(new_n19285_));
  INV_X1     g18988(.I(new_n19285_), .ZN(new_n19286_));
  AOI22_X1   g18989(.A1(new_n13078_), .A2(\b[20] ), .B1(new_n1805_), .B2(new_n12218_), .ZN(new_n19287_));
  OAI21_X1   g18990(.A1(new_n19287_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n19288_));
  XNOR2_X1   g18991(.A1(new_n1808_), .A2(new_n19288_), .ZN(new_n19289_));
  NAND2_X1   g18992(.A1(new_n19038_), .A2(new_n19040_), .ZN(new_n19290_));
  NAND2_X1   g18993(.A1(new_n19290_), .A2(new_n19039_), .ZN(new_n19291_));
  OAI22_X1   g18994(.A1(new_n13880_), .A2(new_n1519_), .B1(new_n1189_), .B2(new_n13885_), .ZN(new_n19292_));
  AOI21_X1   g18995(.A1(new_n19292_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n19293_));
  XNOR2_X1   g18996(.A1(new_n1421_), .A2(new_n19293_), .ZN(new_n19294_));
  NAND2_X1   g18997(.A1(new_n19030_), .A2(new_n18556_), .ZN(new_n19295_));
  NAND2_X1   g18998(.A1(new_n19295_), .A2(new_n19029_), .ZN(new_n19296_));
  NOR2_X1    g18999(.A1(new_n13476_), .A2(new_n1017_), .ZN(new_n19297_));
  XOR2_X1    g19000(.A1(new_n14736_), .A2(new_n1017_), .Z(new_n19298_));
  NAND2_X1   g19001(.A1(new_n19298_), .A2(\b[16] ), .ZN(new_n19299_));
  XOR2_X1    g19002(.A1(new_n19299_), .A2(new_n19297_), .Z(new_n19300_));
  INV_X1     g19003(.I(new_n19300_), .ZN(new_n19301_));
  XOR2_X1    g19004(.A1(new_n19296_), .A2(new_n19301_), .Z(new_n19302_));
  OR2_X2     g19005(.A1(new_n19294_), .A2(new_n19302_), .Z(new_n19303_));
  NOR2_X1    g19006(.A1(new_n19296_), .A2(new_n19300_), .ZN(new_n19304_));
  NAND2_X1   g19007(.A1(new_n19296_), .A2(new_n19300_), .ZN(new_n19305_));
  INV_X1     g19008(.I(new_n19305_), .ZN(new_n19306_));
  OAI21_X1   g19009(.A1(new_n19304_), .A2(new_n19306_), .B(new_n19294_), .ZN(new_n19307_));
  AOI21_X1   g19010(.A1(new_n19303_), .A2(new_n19307_), .B(new_n19291_), .ZN(new_n19308_));
  NAND2_X1   g19011(.A1(new_n19303_), .A2(new_n19307_), .ZN(new_n19309_));
  AOI21_X1   g19012(.A1(new_n19039_), .A2(new_n19290_), .B(new_n19309_), .ZN(new_n19310_));
  NOR2_X1    g19013(.A1(new_n19310_), .A2(new_n19308_), .ZN(new_n19311_));
  NOR2_X1    g19014(.A1(new_n19289_), .A2(new_n19311_), .ZN(new_n19312_));
  XOR2_X1    g19015(.A1(new_n19309_), .A2(new_n19291_), .Z(new_n19313_));
  INV_X1     g19016(.I(new_n19313_), .ZN(new_n19314_));
  AOI21_X1   g19017(.A1(new_n19289_), .A2(new_n19314_), .B(new_n19312_), .ZN(new_n19315_));
  OAI21_X1   g19018(.A1(new_n19018_), .A2(new_n19050_), .B(new_n19048_), .ZN(new_n19316_));
  INV_X1     g19019(.I(new_n19316_), .ZN(new_n19317_));
  AOI22_X1   g19020(.A1(new_n10969_), .A2(new_n2435_), .B1(new_n11394_), .B2(\b[23] ), .ZN(new_n19318_));
  OAI21_X1   g19021(.A1(new_n19318_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n19319_));
  XOR2_X1    g19022(.A1(new_n2280_), .A2(new_n19319_), .Z(new_n19320_));
  NOR2_X1    g19023(.A1(new_n19317_), .A2(new_n19320_), .ZN(new_n19321_));
  INV_X1     g19024(.I(new_n19320_), .ZN(new_n19322_));
  NOR2_X1    g19025(.A1(new_n19322_), .A2(new_n19316_), .ZN(new_n19323_));
  NOR2_X1    g19026(.A1(new_n19323_), .A2(new_n19321_), .ZN(new_n19324_));
  NOR2_X1    g19027(.A1(new_n19324_), .A2(new_n19315_), .ZN(new_n19325_));
  NAND2_X1   g19028(.A1(new_n19314_), .A2(new_n19289_), .ZN(new_n19326_));
  OAI21_X1   g19029(.A1(new_n19289_), .A2(new_n19311_), .B(new_n19326_), .ZN(new_n19327_));
  XOR2_X1    g19030(.A1(new_n19320_), .A2(new_n19316_), .Z(new_n19328_));
  NOR2_X1    g19031(.A1(new_n19328_), .A2(new_n19327_), .ZN(new_n19329_));
  NOR2_X1    g19032(.A1(new_n19325_), .A2(new_n19329_), .ZN(new_n19330_));
  XOR2_X1    g19033(.A1(new_n19330_), .A2(new_n19286_), .Z(new_n19331_));
  NOR2_X1    g19034(.A1(new_n19331_), .A2(new_n19282_), .ZN(new_n19332_));
  OAI21_X1   g19035(.A1(new_n19325_), .A2(new_n19329_), .B(new_n19286_), .ZN(new_n19333_));
  NAND2_X1   g19036(.A1(new_n19330_), .A2(new_n19285_), .ZN(new_n19334_));
  AOI21_X1   g19037(.A1(new_n19333_), .A2(new_n19334_), .B(new_n19281_), .ZN(new_n19335_));
  NOR2_X1    g19038(.A1(new_n19332_), .A2(new_n19335_), .ZN(new_n19336_));
  INV_X1     g19039(.I(new_n19336_), .ZN(new_n19337_));
  NAND2_X1   g19040(.A1(new_n19070_), .A2(new_n19016_), .ZN(new_n19338_));
  NAND2_X1   g19041(.A1(new_n19338_), .A2(new_n19069_), .ZN(new_n19339_));
  OAI22_X1   g19042(.A1(new_n8644_), .A2(new_n3260_), .B1(new_n3709_), .B2(new_n9388_), .ZN(new_n19340_));
  OAI21_X1   g19043(.A1(new_n3018_), .A2(new_n10154_), .B(new_n19340_), .ZN(new_n19341_));
  AOI21_X1   g19044(.A1(new_n19341_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n19342_));
  XNOR2_X1   g19045(.A1(new_n3514_), .A2(new_n19342_), .ZN(new_n19343_));
  INV_X1     g19046(.I(new_n19343_), .ZN(new_n19344_));
  XOR2_X1    g19047(.A1(new_n19339_), .A2(new_n19344_), .Z(new_n19345_));
  NAND2_X1   g19048(.A1(new_n19345_), .A2(new_n19337_), .ZN(new_n19346_));
  NAND2_X1   g19049(.A1(new_n19339_), .A2(new_n19344_), .ZN(new_n19347_));
  INV_X1     g19050(.I(new_n19347_), .ZN(new_n19348_));
  NOR2_X1    g19051(.A1(new_n19339_), .A2(new_n19344_), .ZN(new_n19349_));
  OAI21_X1   g19052(.A1(new_n19348_), .A2(new_n19349_), .B(new_n19336_), .ZN(new_n19350_));
  NAND2_X1   g19053(.A1(new_n19346_), .A2(new_n19350_), .ZN(new_n19351_));
  AOI21_X1   g19054(.A1(new_n19072_), .A2(new_n19082_), .B(new_n19080_), .ZN(new_n19352_));
  XOR2_X1    g19055(.A1(new_n19351_), .A2(new_n19352_), .Z(new_n19353_));
  NOR2_X1    g19056(.A1(new_n19353_), .A2(new_n19277_), .ZN(new_n19354_));
  INV_X1     g19057(.I(new_n19277_), .ZN(new_n19355_));
  INV_X1     g19058(.I(new_n19352_), .ZN(new_n19356_));
  NAND2_X1   g19059(.A1(new_n19351_), .A2(new_n19356_), .ZN(new_n19357_));
  NAND3_X1   g19060(.A1(new_n19352_), .A2(new_n19346_), .A3(new_n19350_), .ZN(new_n19358_));
  AOI21_X1   g19061(.A1(new_n19357_), .A2(new_n19358_), .B(new_n19355_), .ZN(new_n19359_));
  NOR2_X1    g19062(.A1(new_n19354_), .A2(new_n19359_), .ZN(new_n19360_));
  XNOR2_X1   g19063(.A1(new_n19360_), .A2(new_n19273_), .ZN(new_n19361_));
  OAI21_X1   g19064(.A1(new_n19354_), .A2(new_n19359_), .B(new_n19273_), .ZN(new_n19362_));
  INV_X1     g19065(.I(new_n19273_), .ZN(new_n19363_));
  NAND2_X1   g19066(.A1(new_n19363_), .A2(new_n19360_), .ZN(new_n19364_));
  AOI21_X1   g19067(.A1(new_n19364_), .A2(new_n19362_), .B(new_n19271_), .ZN(new_n19365_));
  AOI21_X1   g19068(.A1(new_n19271_), .A2(new_n19361_), .B(new_n19365_), .ZN(new_n19366_));
  XOR2_X1    g19069(.A1(new_n19366_), .A2(new_n19266_), .Z(new_n19367_));
  NAND2_X1   g19070(.A1(new_n19367_), .A2(new_n19264_), .ZN(new_n19368_));
  NOR2_X1    g19071(.A1(new_n19366_), .A2(new_n19266_), .ZN(new_n19369_));
  AND2_X2    g19072(.A1(new_n19366_), .A2(new_n19266_), .Z(new_n19370_));
  OAI21_X1   g19073(.A1(new_n19370_), .A2(new_n19369_), .B(new_n19263_), .ZN(new_n19371_));
  NAND2_X1   g19074(.A1(new_n19368_), .A2(new_n19371_), .ZN(new_n19372_));
  OAI22_X1   g19075(.A1(new_n5420_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n5107_), .ZN(new_n19373_));
  OAI21_X1   g19076(.A1(new_n6229_), .A2(new_n5112_), .B(new_n19373_), .ZN(new_n19374_));
  AOI21_X1   g19077(.A1(new_n19374_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n19375_));
  XOR2_X1    g19078(.A1(new_n6851_), .A2(new_n19375_), .Z(new_n19376_));
  NOR2_X1    g19079(.A1(new_n19372_), .A2(new_n19376_), .ZN(new_n19377_));
  AND2_X2    g19080(.A1(new_n19372_), .A2(new_n19376_), .Z(new_n19378_));
  NOR2_X1    g19081(.A1(new_n19378_), .A2(new_n19377_), .ZN(new_n19379_));
  XOR2_X1    g19082(.A1(new_n19372_), .A2(new_n19376_), .Z(new_n19380_));
  NAND2_X1   g19083(.A1(new_n19380_), .A2(new_n19259_), .ZN(new_n19381_));
  OAI21_X1   g19084(.A1(new_n19259_), .A2(new_n19379_), .B(new_n19381_), .ZN(new_n19382_));
  NAND2_X1   g19085(.A1(new_n19131_), .A2(new_n19008_), .ZN(new_n19383_));
  NAND2_X1   g19086(.A1(new_n19383_), .A2(new_n19130_), .ZN(new_n19384_));
  AND2_X2    g19087(.A1(new_n19382_), .A2(new_n19384_), .Z(new_n19385_));
  NOR2_X1    g19088(.A1(new_n19382_), .A2(new_n19384_), .ZN(new_n19386_));
  OAI21_X1   g19089(.A1(new_n19385_), .A2(new_n19386_), .B(new_n19257_), .ZN(new_n19387_));
  XOR2_X1    g19090(.A1(new_n19382_), .A2(new_n19384_), .Z(new_n19388_));
  NAND2_X1   g19091(.A1(new_n19388_), .A2(new_n19256_), .ZN(new_n19389_));
  NAND2_X1   g19092(.A1(new_n19389_), .A2(new_n19387_), .ZN(new_n19390_));
  XNOR2_X1   g19093(.A1(new_n19390_), .A2(new_n19252_), .ZN(new_n19391_));
  INV_X1     g19094(.I(new_n19252_), .ZN(new_n19392_));
  NAND2_X1   g19095(.A1(new_n19392_), .A2(new_n19390_), .ZN(new_n19393_));
  NAND3_X1   g19096(.A1(new_n19252_), .A2(new_n19387_), .A3(new_n19389_), .ZN(new_n19394_));
  AOI21_X1   g19097(.A1(new_n19393_), .A2(new_n19394_), .B(new_n19251_), .ZN(new_n19395_));
  AOI21_X1   g19098(.A1(new_n19251_), .A2(new_n19391_), .B(new_n19395_), .ZN(new_n19396_));
  XOR2_X1    g19099(.A1(new_n19396_), .A2(new_n19246_), .Z(new_n19397_));
  XOR2_X1    g19100(.A1(new_n19397_), .A2(new_n19242_), .Z(new_n19398_));
  XOR2_X1    g19101(.A1(new_n19398_), .A2(\a[29] ), .Z(new_n19399_));
  XOR2_X1    g19102(.A1(new_n19399_), .A2(new_n19240_), .Z(new_n19400_));
  NAND2_X1   g19103(.A1(new_n19400_), .A2(new_n19238_), .ZN(new_n19401_));
  NOR2_X1    g19104(.A1(new_n19399_), .A2(new_n19240_), .ZN(new_n19402_));
  AND2_X2    g19105(.A1(new_n19399_), .A2(new_n19240_), .Z(new_n19403_));
  OAI21_X1   g19106(.A1(new_n19403_), .A2(new_n19402_), .B(new_n19237_), .ZN(new_n19404_));
  NAND2_X1   g19107(.A1(new_n19401_), .A2(new_n19404_), .ZN(new_n19405_));
  XOR2_X1    g19108(.A1(new_n19405_), .A2(new_n19233_), .Z(new_n19406_));
  XOR2_X1    g19109(.A1(new_n19406_), .A2(new_n19231_), .Z(new_n19407_));
  XOR2_X1    g19110(.A1(new_n19407_), .A2(\a[23] ), .Z(new_n19408_));
  INV_X1     g19111(.I(new_n19408_), .ZN(new_n19409_));
  OAI22_X1   g19112(.A1(new_n1347_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n1344_), .ZN(new_n19410_));
  OAI21_X1   g19113(.A1(new_n12970_), .A2(new_n1457_), .B(new_n19410_), .ZN(new_n19411_));
  AOI21_X1   g19114(.A1(new_n19411_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n19412_));
  XOR2_X1    g19115(.A1(new_n13784_), .A2(new_n19412_), .Z(new_n19413_));
  NOR2_X1    g19116(.A1(new_n19409_), .A2(new_n19413_), .ZN(new_n19414_));
  INV_X1     g19117(.I(new_n19413_), .ZN(new_n19415_));
  NOR2_X1    g19118(.A1(new_n19408_), .A2(new_n19415_), .ZN(new_n19416_));
  OAI21_X1   g19119(.A1(new_n19414_), .A2(new_n19416_), .B(new_n19228_), .ZN(new_n19417_));
  NOR2_X1    g19120(.A1(new_n19408_), .A2(new_n19413_), .ZN(new_n19418_));
  INV_X1     g19121(.I(new_n19418_), .ZN(new_n19419_));
  NAND2_X1   g19122(.A1(new_n19408_), .A2(new_n19413_), .ZN(new_n19420_));
  AOI21_X1   g19123(.A1(new_n19419_), .A2(new_n19420_), .B(new_n19228_), .ZN(new_n19421_));
  INV_X1     g19124(.I(new_n19421_), .ZN(new_n19422_));
  NAND2_X1   g19125(.A1(new_n19422_), .A2(new_n19417_), .ZN(new_n19423_));
  NOR2_X1    g19126(.A1(new_n1332_), .A2(new_n1061_), .ZN(new_n19424_));
  NAND2_X1   g19127(.A1(new_n16148_), .A2(new_n1057_), .ZN(new_n19425_));
  OAI21_X1   g19128(.A1(new_n19424_), .A2(new_n19425_), .B(new_n1056_), .ZN(new_n19426_));
  XNOR2_X1   g19129(.A1(new_n14978_), .A2(new_n19426_), .ZN(new_n19427_));
  NOR2_X1    g19130(.A1(new_n19423_), .A2(new_n19427_), .ZN(new_n19428_));
  INV_X1     g19131(.I(new_n19417_), .ZN(new_n19429_));
  NOR2_X1    g19132(.A1(new_n19429_), .A2(new_n19421_), .ZN(new_n19430_));
  INV_X1     g19133(.I(new_n19427_), .ZN(new_n19431_));
  NOR2_X1    g19134(.A1(new_n19430_), .A2(new_n19431_), .ZN(new_n19432_));
  OAI21_X1   g19135(.A1(new_n19432_), .A2(new_n19428_), .B(new_n19225_), .ZN(new_n19433_));
  INV_X1     g19136(.I(new_n19225_), .ZN(new_n19434_));
  NOR2_X1    g19137(.A1(new_n19430_), .A2(new_n19427_), .ZN(new_n19435_));
  NOR2_X1    g19138(.A1(new_n19423_), .A2(new_n19431_), .ZN(new_n19436_));
  OAI21_X1   g19139(.A1(new_n19435_), .A2(new_n19436_), .B(new_n19434_), .ZN(new_n19437_));
  AOI21_X1   g19140(.A1(new_n19433_), .A2(new_n19437_), .B(new_n19224_), .ZN(new_n19438_));
  XOR2_X1    g19141(.A1(new_n19222_), .A2(new_n19438_), .Z(new_n19439_));
  XOR2_X1    g19142(.A1(new_n19439_), .A2(new_n19218_), .Z(\f[79] ));
  NOR2_X1    g19143(.A1(new_n19218_), .A2(new_n19224_), .ZN(new_n19441_));
  OAI21_X1   g19144(.A1(new_n18951_), .A2(new_n18950_), .B(new_n827_), .ZN(new_n19442_));
  NAND3_X1   g19145(.A1(new_n18946_), .A2(new_n18948_), .A3(\a[14] ), .ZN(new_n19443_));
  INV_X1     g19146(.I(new_n19213_), .ZN(new_n19444_));
  NAND4_X1   g19147(.A1(new_n19444_), .A2(new_n19442_), .A3(new_n19211_), .A4(new_n19443_), .ZN(new_n19445_));
  AOI22_X1   g19148(.A1(new_n19444_), .A2(new_n19211_), .B1(new_n19442_), .B2(new_n19443_), .ZN(new_n19446_));
  OAI21_X1   g19149(.A1(new_n18731_), .A2(new_n19446_), .B(new_n19445_), .ZN(new_n19447_));
  NAND2_X1   g19150(.A1(new_n19433_), .A2(new_n19437_), .ZN(new_n19448_));
  NAND2_X1   g19151(.A1(new_n19218_), .A2(new_n19224_), .ZN(new_n19449_));
  NAND2_X1   g19152(.A1(new_n19448_), .A2(new_n19449_), .ZN(new_n19450_));
  NOR3_X1    g19153(.A1(new_n18972_), .A2(new_n19447_), .A3(new_n19450_), .ZN(new_n19451_));
  NOR2_X1    g19154(.A1(new_n19451_), .A2(new_n19441_), .ZN(new_n19452_));
  NAND2_X1   g19155(.A1(new_n19430_), .A2(new_n19431_), .ZN(new_n19453_));
  OAI21_X1   g19156(.A1(new_n19434_), .A2(new_n19432_), .B(new_n19453_), .ZN(new_n19454_));
  AOI21_X1   g19157(.A1(new_n1056_), .A2(new_n1142_), .B(new_n16486_), .ZN(new_n19455_));
  INV_X1     g19158(.I(new_n19455_), .ZN(new_n19456_));
  AOI21_X1   g19159(.A1(new_n19228_), .A2(new_n19420_), .B(new_n19418_), .ZN(new_n19457_));
  AOI21_X1   g19160(.A1(new_n19401_), .A2(new_n19404_), .B(new_n19232_), .ZN(new_n19458_));
  NOR2_X1    g19161(.A1(new_n19405_), .A2(new_n19233_), .ZN(new_n19459_));
  XOR2_X1    g19162(.A1(new_n19231_), .A2(\a[23] ), .Z(new_n19460_));
  NOR2_X1    g19163(.A1(new_n19459_), .A2(new_n19460_), .ZN(new_n19461_));
  NOR2_X1    g19164(.A1(new_n19461_), .A2(new_n19458_), .ZN(new_n19462_));
  OAI22_X1   g19165(.A1(new_n1347_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n1344_), .ZN(new_n19463_));
  OAI21_X1   g19166(.A1(new_n13367_), .A2(new_n1457_), .B(new_n19463_), .ZN(new_n19464_));
  AOI21_X1   g19167(.A1(new_n18183_), .A2(new_n1340_), .B(new_n19464_), .ZN(new_n19465_));
  OAI22_X1   g19168(.A1(new_n1712_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n1707_), .ZN(new_n19466_));
  OAI21_X1   g19169(.A1(new_n12536_), .A2(new_n1850_), .B(new_n19466_), .ZN(new_n19467_));
  AOI21_X1   g19170(.A1(new_n19467_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n19468_));
  XOR2_X1    g19171(.A1(new_n12969_), .A2(new_n19468_), .Z(new_n19469_));
  NOR2_X1    g19172(.A1(new_n19396_), .A2(new_n19242_), .ZN(new_n19470_));
  XOR2_X1    g19173(.A1(new_n19246_), .A2(\a[29] ), .Z(new_n19471_));
  AOI21_X1   g19174(.A1(new_n19396_), .A2(new_n19242_), .B(new_n19471_), .ZN(new_n19472_));
  NOR2_X1    g19175(.A1(new_n19472_), .A2(new_n19470_), .ZN(new_n19473_));
  OAI22_X1   g19176(.A1(new_n2171_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n2166_), .ZN(new_n19474_));
  OAI21_X1   g19177(.A1(new_n10862_), .A2(new_n2322_), .B(new_n19474_), .ZN(new_n19475_));
  AOI21_X1   g19178(.A1(new_n11748_), .A2(new_n2161_), .B(new_n19475_), .ZN(new_n19476_));
  OAI22_X1   g19179(.A1(new_n10031_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n10477_), .ZN(new_n19477_));
  OAI21_X1   g19180(.A1(new_n10025_), .A2(new_n2884_), .B(new_n19477_), .ZN(new_n19478_));
  AOI21_X1   g19181(.A1(new_n19478_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n19479_));
  XOR2_X1    g19182(.A1(new_n10476_), .A2(new_n19479_), .Z(new_n19480_));
  INV_X1     g19183(.I(new_n19480_), .ZN(new_n19481_));
  OAI22_X1   g19184(.A1(new_n8948_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n9295_), .ZN(new_n19482_));
  OAI21_X1   g19185(.A1(new_n8563_), .A2(new_n3569_), .B(new_n19482_), .ZN(new_n19483_));
  AOI21_X1   g19186(.A1(new_n19483_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n19484_));
  XNOR2_X1   g19187(.A1(new_n9299_), .A2(new_n19484_), .ZN(new_n19485_));
  NOR2_X1    g19188(.A1(new_n19386_), .A2(new_n19256_), .ZN(new_n19486_));
  NOR2_X1    g19189(.A1(new_n19486_), .A2(new_n19385_), .ZN(new_n19487_));
  OAI22_X1   g19190(.A1(new_n5420_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n5107_), .ZN(new_n19488_));
  OAI21_X1   g19191(.A1(new_n6538_), .A2(new_n5112_), .B(new_n19488_), .ZN(new_n19489_));
  AOI21_X1   g19192(.A1(new_n19489_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n19490_));
  XNOR2_X1   g19193(.A1(new_n7202_), .A2(new_n19490_), .ZN(new_n19491_));
  NOR2_X1    g19194(.A1(new_n19369_), .A2(new_n19263_), .ZN(new_n19492_));
  NOR2_X1    g19195(.A1(new_n19492_), .A2(new_n19370_), .ZN(new_n19493_));
  INV_X1     g19196(.I(new_n19493_), .ZN(new_n19494_));
  OAI22_X1   g19197(.A1(new_n5993_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n5991_), .ZN(new_n19495_));
  OAI21_X1   g19198(.A1(new_n5913_), .A2(new_n5997_), .B(new_n19495_), .ZN(new_n19496_));
  AOI21_X1   g19199(.A1(new_n19496_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n19497_));
  XOR2_X1    g19200(.A1(new_n6233_), .A2(new_n19497_), .Z(new_n19498_));
  OAI22_X1   g19201(.A1(new_n6644_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n6647_), .ZN(new_n19499_));
  OAI21_X1   g19202(.A1(new_n4774_), .A2(new_n7284_), .B(new_n19499_), .ZN(new_n19500_));
  AOI21_X1   g19203(.A1(new_n19500_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n19501_));
  XNOR2_X1   g19204(.A1(new_n5357_), .A2(new_n19501_), .ZN(new_n19502_));
  OAI22_X1   g19205(.A1(new_n8644_), .A2(new_n3709_), .B1(new_n3717_), .B2(new_n9388_), .ZN(new_n19503_));
  OAI21_X1   g19206(.A1(new_n3260_), .A2(new_n10154_), .B(new_n19503_), .ZN(new_n19504_));
  AOI21_X1   g19207(.A1(new_n19504_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n19505_));
  XOR2_X1    g19208(.A1(new_n3722_), .A2(new_n19505_), .Z(new_n19506_));
  INV_X1     g19209(.I(new_n19506_), .ZN(new_n19507_));
  AOI22_X1   g19210(.A1(new_n10969_), .A2(new_n18773_), .B1(new_n11394_), .B2(\b[24] ), .ZN(new_n19508_));
  OAI21_X1   g19211(.A1(new_n19508_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n19509_));
  XOR2_X1    g19212(.A1(new_n2443_), .A2(new_n19509_), .Z(new_n19510_));
  NOR2_X1    g19213(.A1(new_n19289_), .A2(new_n19308_), .ZN(new_n19511_));
  NOR2_X1    g19214(.A1(new_n19511_), .A2(new_n19310_), .ZN(new_n19512_));
  OAI22_X1   g19215(.A1(new_n13880_), .A2(new_n1526_), .B1(new_n1294_), .B2(new_n13885_), .ZN(new_n19513_));
  AOI21_X1   g19216(.A1(new_n19513_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n19514_));
  XNOR2_X1   g19217(.A1(new_n1530_), .A2(new_n19514_), .ZN(new_n19515_));
  NOR2_X1    g19218(.A1(new_n13476_), .A2(new_n1109_), .ZN(new_n19516_));
  XOR2_X1    g19219(.A1(new_n14736_), .A2(new_n1109_), .Z(new_n19517_));
  NAND2_X1   g19220(.A1(new_n19517_), .A2(\b[17] ), .ZN(new_n19518_));
  XOR2_X1    g19221(.A1(new_n19518_), .A2(new_n19516_), .Z(new_n19519_));
  NOR2_X1    g19222(.A1(new_n19301_), .A2(new_n19519_), .ZN(new_n19520_));
  INV_X1     g19223(.I(new_n19519_), .ZN(new_n19521_));
  NOR2_X1    g19224(.A1(new_n19521_), .A2(new_n19300_), .ZN(new_n19522_));
  NOR2_X1    g19225(.A1(new_n19520_), .A2(new_n19522_), .ZN(new_n19523_));
  INV_X1     g19226(.I(new_n19523_), .ZN(new_n19524_));
  XOR2_X1    g19227(.A1(new_n19300_), .A2(new_n19519_), .Z(new_n19525_));
  NOR2_X1    g19228(.A1(new_n19515_), .A2(new_n19525_), .ZN(new_n19526_));
  AOI21_X1   g19229(.A1(new_n19515_), .A2(new_n19524_), .B(new_n19526_), .ZN(new_n19527_));
  AOI22_X1   g19230(.A1(new_n13078_), .A2(\b[21] ), .B1(new_n2097_), .B2(new_n12218_), .ZN(new_n19528_));
  OAI21_X1   g19231(.A1(new_n19528_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n19529_));
  XOR2_X1    g19232(.A1(new_n1940_), .A2(new_n19529_), .Z(new_n19530_));
  OAI21_X1   g19233(.A1(new_n19294_), .A2(new_n19304_), .B(new_n19305_), .ZN(new_n19531_));
  XOR2_X1    g19234(.A1(new_n19530_), .A2(new_n19531_), .Z(new_n19532_));
  INV_X1     g19235(.I(new_n19531_), .ZN(new_n19533_));
  NOR2_X1    g19236(.A1(new_n19530_), .A2(new_n19533_), .ZN(new_n19534_));
  AND2_X2    g19237(.A1(new_n19530_), .A2(new_n19533_), .Z(new_n19535_));
  OAI21_X1   g19238(.A1(new_n19535_), .A2(new_n19534_), .B(new_n19527_), .ZN(new_n19536_));
  OAI21_X1   g19239(.A1(new_n19527_), .A2(new_n19532_), .B(new_n19536_), .ZN(new_n19537_));
  XNOR2_X1   g19240(.A1(new_n19537_), .A2(new_n19512_), .ZN(new_n19538_));
  NAND2_X1   g19241(.A1(new_n19537_), .A2(new_n19512_), .ZN(new_n19539_));
  INV_X1     g19242(.I(new_n19539_), .ZN(new_n19540_));
  NOR2_X1    g19243(.A1(new_n19537_), .A2(new_n19512_), .ZN(new_n19541_));
  OAI21_X1   g19244(.A1(new_n19540_), .A2(new_n19541_), .B(new_n19510_), .ZN(new_n19542_));
  OAI21_X1   g19245(.A1(new_n19510_), .A2(new_n19538_), .B(new_n19542_), .ZN(new_n19543_));
  AOI22_X1   g19246(.A1(new_n11415_), .A2(new_n3256_), .B1(\b[27] ), .B2(new_n10145_), .ZN(new_n19544_));
  OAI21_X1   g19247(.A1(new_n19544_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n19545_));
  XNOR2_X1   g19248(.A1(new_n3022_), .A2(new_n19545_), .ZN(new_n19546_));
  NOR2_X1    g19249(.A1(new_n19315_), .A2(new_n19323_), .ZN(new_n19547_));
  NOR2_X1    g19250(.A1(new_n19547_), .A2(new_n19321_), .ZN(new_n19548_));
  INV_X1     g19251(.I(new_n19548_), .ZN(new_n19549_));
  XOR2_X1    g19252(.A1(new_n19546_), .A2(new_n19549_), .Z(new_n19550_));
  NAND2_X1   g19253(.A1(new_n19546_), .A2(new_n19549_), .ZN(new_n19551_));
  NOR2_X1    g19254(.A1(new_n19546_), .A2(new_n19549_), .ZN(new_n19552_));
  INV_X1     g19255(.I(new_n19552_), .ZN(new_n19553_));
  AOI21_X1   g19256(.A1(new_n19551_), .A2(new_n19553_), .B(new_n19543_), .ZN(new_n19554_));
  AOI21_X1   g19257(.A1(new_n19543_), .A2(new_n19550_), .B(new_n19554_), .ZN(new_n19555_));
  INV_X1     g19258(.I(new_n19333_), .ZN(new_n19556_));
  AOI21_X1   g19259(.A1(new_n19281_), .A2(new_n19334_), .B(new_n19556_), .ZN(new_n19557_));
  NOR2_X1    g19260(.A1(new_n19555_), .A2(new_n19557_), .ZN(new_n19558_));
  NAND2_X1   g19261(.A1(new_n19555_), .A2(new_n19557_), .ZN(new_n19559_));
  INV_X1     g19262(.I(new_n19559_), .ZN(new_n19560_));
  OAI21_X1   g19263(.A1(new_n19560_), .A2(new_n19558_), .B(new_n19507_), .ZN(new_n19561_));
  XNOR2_X1   g19264(.A1(new_n19555_), .A2(new_n19557_), .ZN(new_n19562_));
  OAI21_X1   g19265(.A1(new_n19507_), .A2(new_n19562_), .B(new_n19561_), .ZN(new_n19563_));
  OAI22_X1   g19266(.A1(new_n7619_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n8309_), .ZN(new_n19564_));
  OAI21_X1   g19267(.A1(new_n3989_), .A2(new_n7947_), .B(new_n19564_), .ZN(new_n19565_));
  AOI21_X1   g19268(.A1(new_n19565_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n19566_));
  XOR2_X1    g19269(.A1(new_n4499_), .A2(new_n19566_), .Z(new_n19567_));
  OAI21_X1   g19270(.A1(new_n19337_), .A2(new_n19349_), .B(new_n19347_), .ZN(new_n19568_));
  INV_X1     g19271(.I(new_n19568_), .ZN(new_n19569_));
  NOR2_X1    g19272(.A1(new_n19569_), .A2(new_n19567_), .ZN(new_n19570_));
  NAND2_X1   g19273(.A1(new_n19569_), .A2(new_n19567_), .ZN(new_n19571_));
  INV_X1     g19274(.I(new_n19571_), .ZN(new_n19572_));
  OAI21_X1   g19275(.A1(new_n19570_), .A2(new_n19572_), .B(new_n19563_), .ZN(new_n19573_));
  XOR2_X1    g19276(.A1(new_n19567_), .A2(new_n19568_), .Z(new_n19574_));
  OAI21_X1   g19277(.A1(new_n19563_), .A2(new_n19574_), .B(new_n19573_), .ZN(new_n19575_));
  NAND2_X1   g19278(.A1(new_n19358_), .A2(new_n19355_), .ZN(new_n19576_));
  NAND2_X1   g19279(.A1(new_n19576_), .A2(new_n19357_), .ZN(new_n19577_));
  NAND2_X1   g19280(.A1(new_n19575_), .A2(new_n19577_), .ZN(new_n19578_));
  OR2_X2     g19281(.A1(new_n19575_), .A2(new_n19577_), .Z(new_n19579_));
  AOI21_X1   g19282(.A1(new_n19579_), .A2(new_n19578_), .B(new_n19502_), .ZN(new_n19580_));
  INV_X1     g19283(.I(new_n19502_), .ZN(new_n19581_));
  XNOR2_X1   g19284(.A1(new_n19575_), .A2(new_n19577_), .ZN(new_n19582_));
  NOR2_X1    g19285(.A1(new_n19582_), .A2(new_n19581_), .ZN(new_n19583_));
  NOR2_X1    g19286(.A1(new_n19583_), .A2(new_n19580_), .ZN(new_n19584_));
  NAND2_X1   g19287(.A1(new_n19362_), .A2(new_n19271_), .ZN(new_n19585_));
  NAND2_X1   g19288(.A1(new_n19585_), .A2(new_n19364_), .ZN(new_n19586_));
  XOR2_X1    g19289(.A1(new_n19584_), .A2(new_n19586_), .Z(new_n19587_));
  AOI21_X1   g19290(.A1(new_n19364_), .A2(new_n19585_), .B(new_n19584_), .ZN(new_n19588_));
  NOR3_X1    g19291(.A1(new_n19583_), .A2(new_n19586_), .A3(new_n19580_), .ZN(new_n19589_));
  OAI21_X1   g19292(.A1(new_n19588_), .A2(new_n19589_), .B(new_n19498_), .ZN(new_n19590_));
  OAI21_X1   g19293(.A1(new_n19587_), .A2(new_n19498_), .B(new_n19590_), .ZN(new_n19591_));
  XOR2_X1    g19294(.A1(new_n19591_), .A2(new_n19494_), .Z(new_n19592_));
  AND2_X2    g19295(.A1(new_n19591_), .A2(new_n19493_), .Z(new_n19593_));
  NOR2_X1    g19296(.A1(new_n19591_), .A2(new_n19493_), .ZN(new_n19594_));
  OAI21_X1   g19297(.A1(new_n19593_), .A2(new_n19594_), .B(new_n19491_), .ZN(new_n19595_));
  OAI21_X1   g19298(.A1(new_n19491_), .A2(new_n19592_), .B(new_n19595_), .ZN(new_n19596_));
  OAI22_X1   g19299(.A1(new_n4072_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n4067_), .ZN(new_n19597_));
  OAI21_X1   g19300(.A1(new_n7864_), .A2(new_n4318_), .B(new_n19597_), .ZN(new_n19598_));
  AOI21_X1   g19301(.A1(new_n19598_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n19599_));
  XOR2_X1    g19302(.A1(new_n8217_), .A2(new_n19599_), .Z(new_n19600_));
  INV_X1     g19303(.I(new_n19600_), .ZN(new_n19601_));
  INV_X1     g19304(.I(new_n19377_), .ZN(new_n19602_));
  OAI21_X1   g19305(.A1(new_n19259_), .A2(new_n19378_), .B(new_n19602_), .ZN(new_n19603_));
  XOR2_X1    g19306(.A1(new_n19603_), .A2(new_n19601_), .Z(new_n19604_));
  AND2_X2    g19307(.A1(new_n19604_), .A2(new_n19596_), .Z(new_n19605_));
  NAND2_X1   g19308(.A1(new_n19603_), .A2(new_n19601_), .ZN(new_n19606_));
  OR2_X2     g19309(.A1(new_n19603_), .A2(new_n19601_), .Z(new_n19607_));
  AOI21_X1   g19310(.A1(new_n19607_), .A2(new_n19606_), .B(new_n19596_), .ZN(new_n19608_));
  NOR2_X1    g19311(.A1(new_n19605_), .A2(new_n19608_), .ZN(new_n19609_));
  XNOR2_X1   g19312(.A1(new_n19609_), .A2(new_n19487_), .ZN(new_n19610_));
  NOR2_X1    g19313(.A1(new_n19609_), .A2(new_n19487_), .ZN(new_n19611_));
  NOR4_X1    g19314(.A1(new_n19605_), .A2(new_n19385_), .A3(new_n19486_), .A4(new_n19608_), .ZN(new_n19612_));
  OAI21_X1   g19315(.A1(new_n19611_), .A2(new_n19612_), .B(new_n19485_), .ZN(new_n19613_));
  OAI21_X1   g19316(.A1(new_n19610_), .A2(new_n19485_), .B(new_n19613_), .ZN(new_n19614_));
  INV_X1     g19317(.I(new_n19393_), .ZN(new_n19615_));
  AOI21_X1   g19318(.A1(new_n19251_), .A2(new_n19394_), .B(new_n19615_), .ZN(new_n19616_));
  NOR2_X1    g19319(.A1(new_n19616_), .A2(new_n19614_), .ZN(new_n19617_));
  AND2_X2    g19320(.A1(new_n19616_), .A2(new_n19614_), .Z(new_n19618_));
  OAI21_X1   g19321(.A1(new_n19618_), .A2(new_n19617_), .B(new_n19481_), .ZN(new_n19619_));
  XOR2_X1    g19322(.A1(new_n19616_), .A2(new_n19614_), .Z(new_n19620_));
  NAND2_X1   g19323(.A1(new_n19620_), .A2(new_n19480_), .ZN(new_n19621_));
  NAND2_X1   g19324(.A1(new_n19621_), .A2(new_n19619_), .ZN(new_n19622_));
  XOR2_X1    g19325(.A1(new_n19622_), .A2(new_n19476_), .Z(new_n19623_));
  XOR2_X1    g19326(.A1(new_n19623_), .A2(new_n19473_), .Z(new_n19624_));
  XOR2_X1    g19327(.A1(new_n19624_), .A2(\a[26] ), .Z(new_n19625_));
  NOR2_X1    g19328(.A1(new_n19403_), .A2(new_n19237_), .ZN(new_n19626_));
  OAI21_X1   g19329(.A1(new_n19402_), .A2(new_n19626_), .B(new_n19625_), .ZN(new_n19627_));
  INV_X1     g19330(.I(new_n19625_), .ZN(new_n19628_));
  NOR2_X1    g19331(.A1(new_n19626_), .A2(new_n19402_), .ZN(new_n19629_));
  NAND2_X1   g19332(.A1(new_n19628_), .A2(new_n19629_), .ZN(new_n19630_));
  AOI21_X1   g19333(.A1(new_n19630_), .A2(new_n19627_), .B(new_n19469_), .ZN(new_n19631_));
  INV_X1     g19334(.I(new_n19469_), .ZN(new_n19632_));
  XOR2_X1    g19335(.A1(new_n19625_), .A2(new_n19629_), .Z(new_n19633_));
  NOR2_X1    g19336(.A1(new_n19633_), .A2(new_n19632_), .ZN(new_n19634_));
  NOR2_X1    g19337(.A1(new_n19634_), .A2(new_n19631_), .ZN(new_n19635_));
  XOR2_X1    g19338(.A1(new_n19635_), .A2(new_n19465_), .Z(new_n19636_));
  XNOR2_X1   g19339(.A1(new_n19636_), .A2(new_n19462_), .ZN(new_n19637_));
  NOR2_X1    g19340(.A1(new_n19637_), .A2(\a[20] ), .ZN(new_n19638_));
  XOR2_X1    g19341(.A1(new_n19636_), .A2(new_n19462_), .Z(new_n19639_));
  NOR2_X1    g19342(.A1(new_n19639_), .A2(new_n1346_), .ZN(new_n19640_));
  OAI21_X1   g19343(.A1(new_n19638_), .A2(new_n19640_), .B(new_n19457_), .ZN(new_n19641_));
  NOR3_X1    g19344(.A1(new_n19638_), .A2(new_n19640_), .A3(new_n19457_), .ZN(new_n19642_));
  INV_X1     g19345(.I(new_n19642_), .ZN(new_n19643_));
  AOI21_X1   g19346(.A1(new_n19643_), .A2(new_n19641_), .B(new_n19456_), .ZN(new_n19644_));
  INV_X1     g19347(.I(new_n19641_), .ZN(new_n19645_));
  NOR3_X1    g19348(.A1(new_n19645_), .A2(new_n19642_), .A3(new_n19455_), .ZN(new_n19646_));
  OAI21_X1   g19349(.A1(new_n19646_), .A2(new_n19644_), .B(new_n1057_), .ZN(new_n19647_));
  OAI21_X1   g19350(.A1(new_n19645_), .A2(new_n19642_), .B(new_n19455_), .ZN(new_n19648_));
  NAND3_X1   g19351(.A1(new_n19643_), .A2(new_n19456_), .A3(new_n19641_), .ZN(new_n19649_));
  NAND3_X1   g19352(.A1(new_n19648_), .A2(new_n19649_), .A3(\a[17] ), .ZN(new_n19650_));
  AOI21_X1   g19353(.A1(new_n19647_), .A2(new_n19650_), .B(new_n19454_), .ZN(new_n19651_));
  NAND3_X1   g19354(.A1(new_n19454_), .A2(new_n19647_), .A3(new_n19650_), .ZN(new_n19652_));
  INV_X1     g19355(.I(new_n19652_), .ZN(new_n19653_));
  NOR2_X1    g19356(.A1(new_n19653_), .A2(new_n19651_), .ZN(new_n19654_));
  XOR2_X1    g19357(.A1(new_n19452_), .A2(new_n19654_), .Z(\f[80] ));
  INV_X1     g19358(.I(new_n19651_), .ZN(new_n19656_));
  NOR2_X1    g19359(.A1(new_n19638_), .A2(new_n19640_), .ZN(new_n19657_));
  NOR2_X1    g19360(.A1(new_n19657_), .A2(new_n19457_), .ZN(new_n19658_));
  XOR2_X1    g19361(.A1(new_n19455_), .A2(\a[17] ), .Z(new_n19659_));
  AOI21_X1   g19362(.A1(new_n19657_), .A2(new_n19457_), .B(new_n19659_), .ZN(new_n19660_));
  NOR2_X1    g19363(.A1(new_n19660_), .A2(new_n19658_), .ZN(new_n19661_));
  NOR2_X1    g19364(.A1(new_n19635_), .A2(new_n19462_), .ZN(new_n19662_));
  NAND2_X1   g19365(.A1(new_n19635_), .A2(new_n19462_), .ZN(new_n19663_));
  XOR2_X1    g19366(.A1(new_n19465_), .A2(new_n1346_), .Z(new_n19664_));
  INV_X1     g19367(.I(new_n19664_), .ZN(new_n19665_));
  AOI21_X1   g19368(.A1(new_n19663_), .A2(new_n19665_), .B(new_n19662_), .ZN(new_n19666_));
  OAI22_X1   g19369(.A1(new_n1347_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n1344_), .ZN(new_n19667_));
  OAI21_X1   g19370(.A1(new_n13785_), .A2(new_n1457_), .B(new_n19667_), .ZN(new_n19668_));
  AOI21_X1   g19371(.A1(new_n19668_), .A2(new_n1346_), .B(new_n1347_), .ZN(new_n19669_));
  XNOR2_X1   g19372(.A1(new_n14599_), .A2(new_n19669_), .ZN(new_n19670_));
  OAI22_X1   g19373(.A1(new_n1712_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n1707_), .ZN(new_n19671_));
  OAI21_X1   g19374(.A1(new_n12542_), .A2(new_n1850_), .B(new_n19671_), .ZN(new_n19672_));
  AOI21_X1   g19375(.A1(new_n19672_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n19673_));
  XNOR2_X1   g19376(.A1(new_n13371_), .A2(new_n19673_), .ZN(new_n19674_));
  NAND2_X1   g19377(.A1(new_n19630_), .A2(new_n19632_), .ZN(new_n19675_));
  INV_X1     g19378(.I(new_n19622_), .ZN(new_n19676_));
  NOR2_X1    g19379(.A1(new_n19676_), .A2(new_n19473_), .ZN(new_n19677_));
  NAND2_X1   g19380(.A1(new_n19676_), .A2(new_n19473_), .ZN(new_n19678_));
  XOR2_X1    g19381(.A1(new_n19476_), .A2(\a[26] ), .Z(new_n19679_));
  AOI21_X1   g19382(.A1(new_n19678_), .A2(new_n19679_), .B(new_n19677_), .ZN(new_n19680_));
  OAI22_X1   g19383(.A1(new_n10477_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n10862_), .ZN(new_n19681_));
  OAI21_X1   g19384(.A1(new_n10031_), .A2(new_n2884_), .B(new_n19681_), .ZN(new_n19682_));
  AOI21_X1   g19385(.A1(new_n19682_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n19683_));
  XNOR2_X1   g19386(.A1(new_n10866_), .A2(new_n19683_), .ZN(new_n19684_));
  NOR2_X1    g19387(.A1(new_n19618_), .A2(new_n19480_), .ZN(new_n19685_));
  NOR2_X1    g19388(.A1(new_n19685_), .A2(new_n19617_), .ZN(new_n19686_));
  NOR2_X1    g19389(.A1(new_n19612_), .A2(new_n19485_), .ZN(new_n19687_));
  NOR2_X1    g19390(.A1(new_n19593_), .A2(new_n19491_), .ZN(new_n19688_));
  NOR2_X1    g19391(.A1(new_n19688_), .A2(new_n19594_), .ZN(new_n19689_));
  NOR2_X1    g19392(.A1(new_n19589_), .A2(new_n19498_), .ZN(new_n19690_));
  NOR2_X1    g19393(.A1(new_n19588_), .A2(new_n19690_), .ZN(new_n19691_));
  NAND2_X1   g19394(.A1(new_n19579_), .A2(new_n19581_), .ZN(new_n19692_));
  AND2_X2    g19395(.A1(new_n19692_), .A2(new_n19578_), .Z(new_n19693_));
  AOI21_X1   g19396(.A1(new_n19563_), .A2(new_n19571_), .B(new_n19570_), .ZN(new_n19694_));
  AOI21_X1   g19397(.A1(new_n19507_), .A2(new_n19559_), .B(new_n19558_), .ZN(new_n19695_));
  INV_X1     g19398(.I(new_n19695_), .ZN(new_n19696_));
  INV_X1     g19399(.I(new_n19510_), .ZN(new_n19697_));
  AOI21_X1   g19400(.A1(new_n19697_), .A2(new_n19539_), .B(new_n19541_), .ZN(new_n19698_));
  NOR2_X1    g19401(.A1(new_n19535_), .A2(new_n19527_), .ZN(new_n19699_));
  NOR2_X1    g19402(.A1(new_n19699_), .A2(new_n19534_), .ZN(new_n19700_));
  INV_X1     g19403(.I(new_n19700_), .ZN(new_n19701_));
  INV_X1     g19404(.I(new_n19520_), .ZN(new_n19702_));
  AOI21_X1   g19405(.A1(new_n19515_), .A2(new_n19702_), .B(new_n19522_), .ZN(new_n19703_));
  INV_X1     g19406(.I(new_n19703_), .ZN(new_n19704_));
  OAI22_X1   g19407(.A1(new_n13880_), .A2(new_n1796_), .B1(new_n1518_), .B2(new_n13885_), .ZN(new_n19705_));
  AOI21_X1   g19408(.A1(new_n19705_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n19706_));
  XNOR2_X1   g19409(.A1(new_n1638_), .A2(new_n19706_), .ZN(new_n19707_));
  INV_X1     g19410(.I(new_n19707_), .ZN(new_n19708_));
  NOR2_X1    g19411(.A1(new_n13476_), .A2(new_n1189_), .ZN(new_n19709_));
  XOR2_X1    g19412(.A1(new_n14736_), .A2(new_n1189_), .Z(new_n19710_));
  NAND2_X1   g19413(.A1(new_n19710_), .A2(\b[18] ), .ZN(new_n19711_));
  XOR2_X1    g19414(.A1(new_n19711_), .A2(new_n19709_), .Z(new_n19712_));
  XOR2_X1    g19415(.A1(new_n19712_), .A2(\a[17] ), .Z(new_n19713_));
  NOR2_X1    g19416(.A1(new_n19713_), .A2(new_n19519_), .ZN(new_n19714_));
  NOR2_X1    g19417(.A1(new_n19712_), .A2(new_n1057_), .ZN(new_n19715_));
  INV_X1     g19418(.I(new_n19715_), .ZN(new_n19716_));
  NAND2_X1   g19419(.A1(new_n19712_), .A2(new_n1057_), .ZN(new_n19717_));
  AOI21_X1   g19420(.A1(new_n19716_), .A2(new_n19717_), .B(new_n19521_), .ZN(new_n19718_));
  NOR2_X1    g19421(.A1(new_n19714_), .A2(new_n19718_), .ZN(new_n19719_));
  NOR2_X1    g19422(.A1(new_n19708_), .A2(new_n19719_), .ZN(new_n19720_));
  NAND2_X1   g19423(.A1(new_n19708_), .A2(new_n19719_), .ZN(new_n19721_));
  INV_X1     g19424(.I(new_n19721_), .ZN(new_n19722_));
  OAI21_X1   g19425(.A1(new_n19722_), .A2(new_n19720_), .B(new_n19704_), .ZN(new_n19723_));
  XNOR2_X1   g19426(.A1(new_n19707_), .A2(new_n19719_), .ZN(new_n19724_));
  NAND2_X1   g19427(.A1(new_n19724_), .A2(new_n19703_), .ZN(new_n19725_));
  NAND2_X1   g19428(.A1(new_n19723_), .A2(new_n19725_), .ZN(new_n19726_));
  AOI22_X1   g19429(.A1(new_n13078_), .A2(\b[22] ), .B1(new_n18260_), .B2(new_n12218_), .ZN(new_n19727_));
  OAI21_X1   g19430(.A1(new_n19727_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n19728_));
  XNOR2_X1   g19431(.A1(new_n2106_), .A2(new_n19728_), .ZN(new_n19729_));
  XNOR2_X1   g19432(.A1(new_n19726_), .A2(new_n19729_), .ZN(new_n19730_));
  INV_X1     g19433(.I(new_n19726_), .ZN(new_n19731_));
  NOR2_X1    g19434(.A1(new_n19731_), .A2(new_n19729_), .ZN(new_n19732_));
  INV_X1     g19435(.I(new_n19729_), .ZN(new_n19733_));
  NOR2_X1    g19436(.A1(new_n19733_), .A2(new_n19726_), .ZN(new_n19734_));
  NOR2_X1    g19437(.A1(new_n19732_), .A2(new_n19734_), .ZN(new_n19735_));
  NOR2_X1    g19438(.A1(new_n19735_), .A2(new_n19701_), .ZN(new_n19736_));
  AOI21_X1   g19439(.A1(new_n19701_), .A2(new_n19730_), .B(new_n19736_), .ZN(new_n19737_));
  AOI22_X1   g19440(.A1(new_n10969_), .A2(new_n2838_), .B1(new_n11394_), .B2(\b[25] ), .ZN(new_n19738_));
  OAI21_X1   g19441(.A1(new_n19738_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n19739_));
  XOR2_X1    g19442(.A1(new_n2647_), .A2(new_n19739_), .Z(new_n19740_));
  XOR2_X1    g19443(.A1(new_n19737_), .A2(new_n19740_), .Z(new_n19741_));
  NOR2_X1    g19444(.A1(new_n19741_), .A2(new_n19698_), .ZN(new_n19742_));
  INV_X1     g19445(.I(new_n19698_), .ZN(new_n19743_));
  INV_X1     g19446(.I(new_n19737_), .ZN(new_n19744_));
  NOR2_X1    g19447(.A1(new_n19744_), .A2(new_n19740_), .ZN(new_n19745_));
  INV_X1     g19448(.I(new_n19745_), .ZN(new_n19746_));
  NAND2_X1   g19449(.A1(new_n19744_), .A2(new_n19740_), .ZN(new_n19747_));
  AOI21_X1   g19450(.A1(new_n19746_), .A2(new_n19747_), .B(new_n19743_), .ZN(new_n19748_));
  NOR2_X1    g19451(.A1(new_n19748_), .A2(new_n19742_), .ZN(new_n19749_));
  INV_X1     g19452(.I(new_n19749_), .ZN(new_n19750_));
  INV_X1     g19453(.I(new_n3261_), .ZN(new_n19751_));
  AOI22_X1   g19454(.A1(new_n11415_), .A2(new_n19751_), .B1(\b[28] ), .B2(new_n10145_), .ZN(new_n19752_));
  OAI21_X1   g19455(.A1(new_n19752_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n19753_));
  XOR2_X1    g19456(.A1(new_n3264_), .A2(new_n19753_), .Z(new_n19754_));
  OAI21_X1   g19457(.A1(new_n19543_), .A2(new_n19552_), .B(new_n19551_), .ZN(new_n19755_));
  INV_X1     g19458(.I(new_n19755_), .ZN(new_n19756_));
  NOR2_X1    g19459(.A1(new_n19756_), .A2(new_n19754_), .ZN(new_n19757_));
  NAND2_X1   g19460(.A1(new_n19756_), .A2(new_n19754_), .ZN(new_n19758_));
  INV_X1     g19461(.I(new_n19758_), .ZN(new_n19759_));
  OAI21_X1   g19462(.A1(new_n19759_), .A2(new_n19757_), .B(new_n19750_), .ZN(new_n19760_));
  XNOR2_X1   g19463(.A1(new_n19755_), .A2(new_n19754_), .ZN(new_n19761_));
  NAND2_X1   g19464(.A1(new_n19749_), .A2(new_n19761_), .ZN(new_n19762_));
  NAND2_X1   g19465(.A1(new_n19760_), .A2(new_n19762_), .ZN(new_n19763_));
  OAI22_X1   g19466(.A1(new_n8644_), .A2(new_n3717_), .B1(new_n3989_), .B2(new_n9388_), .ZN(new_n19764_));
  OAI21_X1   g19467(.A1(new_n3709_), .A2(new_n10154_), .B(new_n19764_), .ZN(new_n19765_));
  AOI21_X1   g19468(.A1(new_n19765_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n19766_));
  XNOR2_X1   g19469(.A1(new_n3993_), .A2(new_n19766_), .ZN(new_n19767_));
  OR2_X2     g19470(.A1(new_n19763_), .A2(new_n19767_), .Z(new_n19768_));
  NAND2_X1   g19471(.A1(new_n19763_), .A2(new_n19767_), .ZN(new_n19769_));
  NAND2_X1   g19472(.A1(new_n19768_), .A2(new_n19769_), .ZN(new_n19770_));
  NAND2_X1   g19473(.A1(new_n19770_), .A2(new_n19696_), .ZN(new_n19771_));
  XOR2_X1    g19474(.A1(new_n19763_), .A2(new_n19767_), .Z(new_n19772_));
  NAND2_X1   g19475(.A1(new_n19772_), .A2(new_n19695_), .ZN(new_n19773_));
  NAND2_X1   g19476(.A1(new_n19771_), .A2(new_n19773_), .ZN(new_n19774_));
  OAI22_X1   g19477(.A1(new_n7619_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n8309_), .ZN(new_n19775_));
  OAI21_X1   g19478(.A1(new_n4253_), .A2(new_n7947_), .B(new_n19775_), .ZN(new_n19776_));
  AOI21_X1   g19479(.A1(new_n19776_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n19777_));
  XNOR2_X1   g19480(.A1(new_n4778_), .A2(new_n19777_), .ZN(new_n19778_));
  XOR2_X1    g19481(.A1(new_n19774_), .A2(new_n19778_), .Z(new_n19779_));
  NOR2_X1    g19482(.A1(new_n19779_), .A2(new_n19694_), .ZN(new_n19780_));
  INV_X1     g19483(.I(new_n19694_), .ZN(new_n19781_));
  INV_X1     g19484(.I(new_n19778_), .ZN(new_n19782_));
  NAND2_X1   g19485(.A1(new_n19774_), .A2(new_n19782_), .ZN(new_n19783_));
  NOR2_X1    g19486(.A1(new_n19774_), .A2(new_n19782_), .ZN(new_n19784_));
  INV_X1     g19487(.I(new_n19784_), .ZN(new_n19785_));
  AOI21_X1   g19488(.A1(new_n19785_), .A2(new_n19783_), .B(new_n19781_), .ZN(new_n19786_));
  OAI22_X1   g19489(.A1(new_n6644_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n6647_), .ZN(new_n19787_));
  OAI21_X1   g19490(.A1(new_n5068_), .A2(new_n7284_), .B(new_n19787_), .ZN(new_n19788_));
  AOI21_X1   g19491(.A1(new_n19788_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n19789_));
  XNOR2_X1   g19492(.A1(new_n5600_), .A2(new_n19789_), .ZN(new_n19790_));
  NOR3_X1    g19493(.A1(new_n19780_), .A2(new_n19786_), .A3(new_n19790_), .ZN(new_n19791_));
  NOR2_X1    g19494(.A1(new_n19780_), .A2(new_n19786_), .ZN(new_n19792_));
  INV_X1     g19495(.I(new_n19790_), .ZN(new_n19793_));
  NOR2_X1    g19496(.A1(new_n19792_), .A2(new_n19793_), .ZN(new_n19794_));
  NOR2_X1    g19497(.A1(new_n19794_), .A2(new_n19791_), .ZN(new_n19795_));
  XOR2_X1    g19498(.A1(new_n19792_), .A2(new_n19793_), .Z(new_n19796_));
  NAND2_X1   g19499(.A1(new_n19796_), .A2(new_n19693_), .ZN(new_n19797_));
  OAI21_X1   g19500(.A1(new_n19693_), .A2(new_n19795_), .B(new_n19797_), .ZN(new_n19798_));
  OAI22_X1   g19501(.A1(new_n5993_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n5991_), .ZN(new_n19799_));
  OAI21_X1   g19502(.A1(new_n5921_), .A2(new_n5997_), .B(new_n19799_), .ZN(new_n19800_));
  AOI21_X1   g19503(.A1(new_n19800_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n19801_));
  XOR2_X1    g19504(.A1(new_n6543_), .A2(new_n19801_), .Z(new_n19802_));
  XOR2_X1    g19505(.A1(new_n19798_), .A2(new_n19802_), .Z(new_n19803_));
  INV_X1     g19506(.I(new_n19802_), .ZN(new_n19804_));
  NAND2_X1   g19507(.A1(new_n19798_), .A2(new_n19804_), .ZN(new_n19805_));
  INV_X1     g19508(.I(new_n19805_), .ZN(new_n19806_));
  NOR2_X1    g19509(.A1(new_n19798_), .A2(new_n19804_), .ZN(new_n19807_));
  OAI21_X1   g19510(.A1(new_n19806_), .A2(new_n19807_), .B(new_n19691_), .ZN(new_n19808_));
  OAI21_X1   g19511(.A1(new_n19691_), .A2(new_n19803_), .B(new_n19808_), .ZN(new_n19809_));
  AOI22_X1   g19512(.A1(new_n4859_), .A2(\b[44] ), .B1(new_n4865_), .B2(\b[45] ), .ZN(new_n19810_));
  AOI21_X1   g19513(.A1(\b[43] ), .A2(new_n6005_), .B(new_n19810_), .ZN(new_n19811_));
  OAI21_X1   g19514(.A1(new_n19811_), .A2(\a[38] ), .B(new_n4859_), .ZN(new_n19812_));
  XNOR2_X1   g19515(.A1(new_n7516_), .A2(new_n19812_), .ZN(new_n19813_));
  XNOR2_X1   g19516(.A1(new_n19809_), .A2(new_n19813_), .ZN(new_n19814_));
  NOR2_X1    g19517(.A1(new_n19814_), .A2(new_n19689_), .ZN(new_n19815_));
  NOR2_X1    g19518(.A1(new_n19809_), .A2(new_n19813_), .ZN(new_n19816_));
  INV_X1     g19519(.I(new_n19816_), .ZN(new_n19817_));
  NAND2_X1   g19520(.A1(new_n19809_), .A2(new_n19813_), .ZN(new_n19818_));
  NAND2_X1   g19521(.A1(new_n19817_), .A2(new_n19818_), .ZN(new_n19819_));
  AOI21_X1   g19522(.A1(new_n19689_), .A2(new_n19819_), .B(new_n19815_), .ZN(new_n19820_));
  AOI22_X1   g19523(.A1(new_n4062_), .A2(\b[47] ), .B1(new_n5438_), .B2(\b[48] ), .ZN(new_n19821_));
  AOI21_X1   g19524(.A1(\b[46] ), .A2(new_n4319_), .B(new_n19821_), .ZN(new_n19822_));
  OAI21_X1   g19525(.A1(new_n19822_), .A2(\a[35] ), .B(new_n4062_), .ZN(new_n19823_));
  XOR2_X1    g19526(.A1(new_n8568_), .A2(new_n19823_), .Z(new_n19824_));
  INV_X1     g19527(.I(new_n19607_), .ZN(new_n19825_));
  OAI21_X1   g19528(.A1(new_n19825_), .A2(new_n19596_), .B(new_n19606_), .ZN(new_n19826_));
  NAND2_X1   g19529(.A1(new_n19826_), .A2(new_n19824_), .ZN(new_n19827_));
  NOR2_X1    g19530(.A1(new_n19826_), .A2(new_n19824_), .ZN(new_n19828_));
  INV_X1     g19531(.I(new_n19828_), .ZN(new_n19829_));
  AOI21_X1   g19532(.A1(new_n19829_), .A2(new_n19827_), .B(new_n19820_), .ZN(new_n19830_));
  INV_X1     g19533(.I(new_n19820_), .ZN(new_n19831_));
  XNOR2_X1   g19534(.A1(new_n19826_), .A2(new_n19824_), .ZN(new_n19832_));
  NOR2_X1    g19535(.A1(new_n19831_), .A2(new_n19832_), .ZN(new_n19833_));
  OAI22_X1   g19536(.A1(new_n9295_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n10025_), .ZN(new_n19834_));
  OAI21_X1   g19537(.A1(new_n8948_), .A2(new_n3569_), .B(new_n19834_), .ZN(new_n19835_));
  AOI21_X1   g19538(.A1(new_n19835_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n19836_));
  XNOR2_X1   g19539(.A1(new_n9642_), .A2(new_n19836_), .ZN(new_n19837_));
  NOR3_X1    g19540(.A1(new_n19833_), .A2(new_n19830_), .A3(new_n19837_), .ZN(new_n19838_));
  NOR2_X1    g19541(.A1(new_n19833_), .A2(new_n19830_), .ZN(new_n19839_));
  INV_X1     g19542(.I(new_n19837_), .ZN(new_n19840_));
  NOR2_X1    g19543(.A1(new_n19839_), .A2(new_n19840_), .ZN(new_n19841_));
  OAI22_X1   g19544(.A1(new_n19841_), .A2(new_n19838_), .B1(new_n19611_), .B2(new_n19687_), .ZN(new_n19842_));
  NOR2_X1    g19545(.A1(new_n19687_), .A2(new_n19611_), .ZN(new_n19843_));
  XOR2_X1    g19546(.A1(new_n19839_), .A2(new_n19840_), .Z(new_n19844_));
  NAND2_X1   g19547(.A1(new_n19844_), .A2(new_n19843_), .ZN(new_n19845_));
  NAND2_X1   g19548(.A1(new_n19845_), .A2(new_n19842_), .ZN(new_n19846_));
  INV_X1     g19549(.I(new_n19846_), .ZN(new_n19847_));
  NOR2_X1    g19550(.A1(new_n19847_), .A2(new_n19686_), .ZN(new_n19848_));
  NOR3_X1    g19551(.A1(new_n19846_), .A2(new_n19617_), .A3(new_n19685_), .ZN(new_n19849_));
  NOR2_X1    g19552(.A1(new_n19848_), .A2(new_n19849_), .ZN(new_n19850_));
  NOR2_X1    g19553(.A1(new_n19850_), .A2(new_n19684_), .ZN(new_n19851_));
  INV_X1     g19554(.I(new_n19684_), .ZN(new_n19852_));
  XOR2_X1    g19555(.A1(new_n19846_), .A2(new_n19686_), .Z(new_n19853_));
  NOR2_X1    g19556(.A1(new_n19853_), .A2(new_n19852_), .ZN(new_n19854_));
  NOR2_X1    g19557(.A1(new_n19851_), .A2(new_n19854_), .ZN(new_n19855_));
  OAI22_X1   g19558(.A1(new_n2171_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n2166_), .ZN(new_n19856_));
  OAI21_X1   g19559(.A1(new_n11738_), .A2(new_n2322_), .B(new_n19856_), .ZN(new_n19857_));
  AOI21_X1   g19560(.A1(new_n19857_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n19858_));
  XNOR2_X1   g19561(.A1(new_n12128_), .A2(new_n19858_), .ZN(new_n19859_));
  NOR2_X1    g19562(.A1(new_n19855_), .A2(new_n19859_), .ZN(new_n19860_));
  INV_X1     g19563(.I(new_n19859_), .ZN(new_n19861_));
  NOR3_X1    g19564(.A1(new_n19851_), .A2(new_n19854_), .A3(new_n19861_), .ZN(new_n19862_));
  NOR2_X1    g19565(.A1(new_n19860_), .A2(new_n19862_), .ZN(new_n19863_));
  NOR2_X1    g19566(.A1(new_n19863_), .A2(new_n19680_), .ZN(new_n19864_));
  XOR2_X1    g19567(.A1(new_n19855_), .A2(new_n19861_), .Z(new_n19865_));
  INV_X1     g19568(.I(new_n19865_), .ZN(new_n19866_));
  AOI21_X1   g19569(.A1(new_n19866_), .A2(new_n19680_), .B(new_n19864_), .ZN(new_n19867_));
  AOI21_X1   g19570(.A1(new_n19627_), .A2(new_n19675_), .B(new_n19867_), .ZN(new_n19868_));
  INV_X1     g19571(.I(new_n19868_), .ZN(new_n19869_));
  NAND2_X1   g19572(.A1(new_n19675_), .A2(new_n19627_), .ZN(new_n19870_));
  INV_X1     g19573(.I(new_n19867_), .ZN(new_n19871_));
  NOR2_X1    g19574(.A1(new_n19871_), .A2(new_n19870_), .ZN(new_n19872_));
  INV_X1     g19575(.I(new_n19872_), .ZN(new_n19873_));
  AOI21_X1   g19576(.A1(new_n19873_), .A2(new_n19869_), .B(new_n19674_), .ZN(new_n19874_));
  INV_X1     g19577(.I(new_n19674_), .ZN(new_n19875_));
  XOR2_X1    g19578(.A1(new_n19870_), .A2(new_n19867_), .Z(new_n19876_));
  NOR2_X1    g19579(.A1(new_n19876_), .A2(new_n19875_), .ZN(new_n19877_));
  NOR2_X1    g19580(.A1(new_n19877_), .A2(new_n19874_), .ZN(new_n19878_));
  NOR2_X1    g19581(.A1(new_n19878_), .A2(new_n19670_), .ZN(new_n19879_));
  INV_X1     g19582(.I(new_n19879_), .ZN(new_n19880_));
  NAND2_X1   g19583(.A1(new_n19878_), .A2(new_n19670_), .ZN(new_n19881_));
  AOI21_X1   g19584(.A1(new_n19880_), .A2(new_n19881_), .B(new_n19666_), .ZN(new_n19882_));
  XOR2_X1    g19585(.A1(new_n19878_), .A2(new_n19670_), .Z(new_n19883_));
  AOI21_X1   g19586(.A1(new_n19666_), .A2(new_n19883_), .B(new_n19882_), .ZN(new_n19884_));
  XOR2_X1    g19587(.A1(new_n19661_), .A2(new_n19884_), .Z(new_n19885_));
  OAI21_X1   g19588(.A1(new_n19652_), .A2(new_n19885_), .B(new_n19656_), .ZN(new_n19886_));
  XNOR2_X1   g19589(.A1(new_n19452_), .A2(new_n19886_), .ZN(\f[81] ));
  NAND2_X1   g19590(.A1(new_n19661_), .A2(new_n19884_), .ZN(new_n19888_));
  INV_X1     g19591(.I(new_n19441_), .ZN(new_n19889_));
  AOI22_X1   g19592(.A1(new_n19218_), .A2(new_n19224_), .B1(new_n19433_), .B2(new_n19437_), .ZN(new_n19890_));
  NAND3_X1   g19593(.A1(new_n18728_), .A2(new_n19221_), .A3(new_n19890_), .ZN(new_n19891_));
  NOR2_X1    g19594(.A1(new_n19653_), .A2(new_n19651_), .ZN(new_n19892_));
  AOI21_X1   g19595(.A1(new_n19891_), .A2(new_n19889_), .B(new_n19892_), .ZN(new_n19893_));
  INV_X1     g19596(.I(new_n19881_), .ZN(new_n19894_));
  OAI21_X1   g19597(.A1(new_n19666_), .A2(new_n19894_), .B(new_n19880_), .ZN(new_n19895_));
  INV_X1     g19598(.I(new_n19895_), .ZN(new_n19896_));
  NOR2_X1    g19599(.A1(new_n1457_), .A2(new_n1344_), .ZN(new_n19897_));
  NAND2_X1   g19600(.A1(new_n16148_), .A2(new_n1346_), .ZN(new_n19898_));
  OAI21_X1   g19601(.A1(new_n19897_), .A2(new_n19898_), .B(new_n1340_), .ZN(new_n19899_));
  XNOR2_X1   g19602(.A1(new_n14978_), .A2(new_n19899_), .ZN(new_n19900_));
  OAI22_X1   g19603(.A1(new_n1712_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n1707_), .ZN(new_n19901_));
  OAI21_X1   g19604(.A1(new_n12970_), .A2(new_n1850_), .B(new_n19901_), .ZN(new_n19902_));
  AOI21_X1   g19605(.A1(new_n19902_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n19903_));
  XOR2_X1    g19606(.A1(new_n13784_), .A2(new_n19903_), .Z(new_n19904_));
  INV_X1     g19607(.I(new_n19904_), .ZN(new_n19905_));
  NOR2_X1    g19608(.A1(new_n19862_), .A2(new_n19680_), .ZN(new_n19906_));
  OAI22_X1   g19609(.A1(new_n2171_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n2166_), .ZN(new_n19907_));
  OAI21_X1   g19610(.A1(new_n11744_), .A2(new_n2322_), .B(new_n19907_), .ZN(new_n19908_));
  AOI21_X1   g19611(.A1(new_n19908_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n19909_));
  XNOR2_X1   g19612(.A1(new_n12546_), .A2(new_n19909_), .ZN(new_n19910_));
  INV_X1     g19613(.I(new_n19849_), .ZN(new_n19911_));
  AOI21_X1   g19614(.A1(new_n19911_), .A2(new_n19852_), .B(new_n19848_), .ZN(new_n19912_));
  OAI22_X1   g19615(.A1(new_n10862_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n11738_), .ZN(new_n19913_));
  OAI21_X1   g19616(.A1(new_n10477_), .A2(new_n2884_), .B(new_n19913_), .ZN(new_n19914_));
  AOI21_X1   g19617(.A1(new_n19914_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n19915_));
  XOR2_X1    g19618(.A1(new_n11298_), .A2(new_n19915_), .Z(new_n19916_));
  NOR2_X1    g19619(.A1(new_n19841_), .A2(new_n19843_), .ZN(new_n19917_));
  NOR2_X1    g19620(.A1(new_n19917_), .A2(new_n19838_), .ZN(new_n19918_));
  INV_X1     g19621(.I(new_n19918_), .ZN(new_n19919_));
  OAI22_X1   g19622(.A1(new_n10025_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n10031_), .ZN(new_n19920_));
  OAI21_X1   g19623(.A1(new_n9295_), .A2(new_n3569_), .B(new_n19920_), .ZN(new_n19921_));
  AOI21_X1   g19624(.A1(new_n19921_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n19922_));
  XNOR2_X1   g19625(.A1(new_n10035_), .A2(new_n19922_), .ZN(new_n19923_));
  OAI21_X1   g19626(.A1(new_n19831_), .A2(new_n19828_), .B(new_n19827_), .ZN(new_n19924_));
  OAI22_X1   g19627(.A1(new_n5420_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n5107_), .ZN(new_n19925_));
  OAI21_X1   g19628(.A1(new_n7198_), .A2(new_n5112_), .B(new_n19925_), .ZN(new_n19926_));
  AOI21_X1   g19629(.A1(new_n19926_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n19927_));
  XNOR2_X1   g19630(.A1(new_n7874_), .A2(new_n19927_), .ZN(new_n19928_));
  NOR2_X1    g19631(.A1(new_n19794_), .A2(new_n19693_), .ZN(new_n19929_));
  NOR2_X1    g19632(.A1(new_n19929_), .A2(new_n19791_), .ZN(new_n19930_));
  INV_X1     g19633(.I(new_n19930_), .ZN(new_n19931_));
  OAI22_X1   g19634(.A1(new_n6644_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n6647_), .ZN(new_n19932_));
  OAI21_X1   g19635(.A1(new_n5353_), .A2(new_n7284_), .B(new_n19932_), .ZN(new_n19933_));
  AOI21_X1   g19636(.A1(new_n19933_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n19934_));
  XOR2_X1    g19637(.A1(new_n5926_), .A2(new_n19934_), .Z(new_n19935_));
  INV_X1     g19638(.I(new_n19935_), .ZN(new_n19936_));
  OAI21_X1   g19639(.A1(new_n19694_), .A2(new_n19784_), .B(new_n19783_), .ZN(new_n19937_));
  AOI22_X1   g19640(.A1(new_n8631_), .A2(\b[33] ), .B1(\b[34] ), .B2(new_n9382_), .ZN(new_n19938_));
  AOI21_X1   g19641(.A1(\b[32] ), .A2(new_n9731_), .B(new_n19938_), .ZN(new_n19939_));
  OAI21_X1   g19642(.A1(new_n19939_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n19940_));
  XOR2_X1    g19643(.A1(new_n4257_), .A2(new_n19940_), .Z(new_n19941_));
  INV_X1     g19644(.I(new_n19941_), .ZN(new_n19942_));
  AOI22_X1   g19645(.A1(new_n10969_), .A2(new_n19278_), .B1(new_n11394_), .B2(\b[26] ), .ZN(new_n19943_));
  OAI21_X1   g19646(.A1(new_n19943_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n19944_));
  XOR2_X1    g19647(.A1(new_n2846_), .A2(new_n19944_), .Z(new_n19945_));
  NOR2_X1    g19648(.A1(new_n19734_), .A2(new_n19700_), .ZN(new_n19946_));
  NOR2_X1    g19649(.A1(new_n19946_), .A2(new_n19732_), .ZN(new_n19947_));
  OAI22_X1   g19650(.A1(new_n13880_), .A2(new_n1804_), .B1(new_n1525_), .B2(new_n13885_), .ZN(new_n19948_));
  AOI21_X1   g19651(.A1(new_n19948_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n19949_));
  XNOR2_X1   g19652(.A1(new_n1808_), .A2(new_n19949_), .ZN(new_n19950_));
  NAND2_X1   g19653(.A1(new_n19717_), .A2(new_n19521_), .ZN(new_n19951_));
  NAND2_X1   g19654(.A1(new_n19951_), .A2(new_n19716_), .ZN(new_n19952_));
  NOR2_X1    g19655(.A1(new_n13476_), .A2(new_n1294_), .ZN(new_n19953_));
  XOR2_X1    g19656(.A1(new_n14736_), .A2(new_n1294_), .Z(new_n19954_));
  NAND2_X1   g19657(.A1(new_n19954_), .A2(\b[19] ), .ZN(new_n19955_));
  XOR2_X1    g19658(.A1(new_n19955_), .A2(new_n19953_), .Z(new_n19956_));
  INV_X1     g19659(.I(new_n19956_), .ZN(new_n19957_));
  XOR2_X1    g19660(.A1(new_n19952_), .A2(new_n19957_), .Z(new_n19958_));
  INV_X1     g19661(.I(new_n19958_), .ZN(new_n19959_));
  NOR2_X1    g19662(.A1(new_n19952_), .A2(new_n19956_), .ZN(new_n19960_));
  INV_X1     g19663(.I(new_n19960_), .ZN(new_n19961_));
  NAND2_X1   g19664(.A1(new_n19952_), .A2(new_n19956_), .ZN(new_n19962_));
  AOI21_X1   g19665(.A1(new_n19961_), .A2(new_n19962_), .B(new_n19950_), .ZN(new_n19963_));
  AOI21_X1   g19666(.A1(new_n19950_), .A2(new_n19959_), .B(new_n19963_), .ZN(new_n19964_));
  OAI21_X1   g19667(.A1(new_n19703_), .A2(new_n19720_), .B(new_n19721_), .ZN(new_n19965_));
  AOI22_X1   g19668(.A1(new_n13078_), .A2(\b[23] ), .B1(new_n2435_), .B2(new_n12218_), .ZN(new_n19966_));
  OAI21_X1   g19669(.A1(new_n19966_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n19967_));
  XOR2_X1    g19670(.A1(new_n2280_), .A2(new_n19967_), .Z(new_n19968_));
  XOR2_X1    g19671(.A1(new_n19968_), .A2(new_n19965_), .Z(new_n19969_));
  NOR2_X1    g19672(.A1(new_n19964_), .A2(new_n19969_), .ZN(new_n19970_));
  INV_X1     g19673(.I(new_n19965_), .ZN(new_n19971_));
  NOR2_X1    g19674(.A1(new_n19971_), .A2(new_n19968_), .ZN(new_n19972_));
  INV_X1     g19675(.I(new_n19972_), .ZN(new_n19973_));
  NAND2_X1   g19676(.A1(new_n19971_), .A2(new_n19968_), .ZN(new_n19974_));
  NAND2_X1   g19677(.A1(new_n19973_), .A2(new_n19974_), .ZN(new_n19975_));
  AOI21_X1   g19678(.A1(new_n19964_), .A2(new_n19975_), .B(new_n19970_), .ZN(new_n19976_));
  XNOR2_X1   g19679(.A1(new_n19976_), .A2(new_n19947_), .ZN(new_n19977_));
  NOR2_X1    g19680(.A1(new_n19977_), .A2(new_n19945_), .ZN(new_n19978_));
  INV_X1     g19681(.I(new_n19945_), .ZN(new_n19979_));
  NOR2_X1    g19682(.A1(new_n19976_), .A2(new_n19947_), .ZN(new_n19980_));
  INV_X1     g19683(.I(new_n19980_), .ZN(new_n19981_));
  NAND2_X1   g19684(.A1(new_n19976_), .A2(new_n19947_), .ZN(new_n19982_));
  AOI21_X1   g19685(.A1(new_n19981_), .A2(new_n19982_), .B(new_n19979_), .ZN(new_n19983_));
  NOR2_X1    g19686(.A1(new_n19978_), .A2(new_n19983_), .ZN(new_n19984_));
  AOI21_X1   g19687(.A1(new_n19743_), .A2(new_n19747_), .B(new_n19745_), .ZN(new_n19985_));
  AOI22_X1   g19688(.A1(new_n11415_), .A2(new_n3711_), .B1(\b[29] ), .B2(new_n10145_), .ZN(new_n19986_));
  OAI21_X1   g19689(.A1(new_n19986_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n19987_));
  XOR2_X1    g19690(.A1(new_n3514_), .A2(new_n19987_), .Z(new_n19988_));
  XNOR2_X1   g19691(.A1(new_n19985_), .A2(new_n19988_), .ZN(new_n19989_));
  NOR2_X1    g19692(.A1(new_n19989_), .A2(new_n19984_), .ZN(new_n19990_));
  INV_X1     g19693(.I(new_n19984_), .ZN(new_n19991_));
  NOR2_X1    g19694(.A1(new_n19985_), .A2(new_n19988_), .ZN(new_n19992_));
  INV_X1     g19695(.I(new_n19992_), .ZN(new_n19993_));
  NAND2_X1   g19696(.A1(new_n19985_), .A2(new_n19988_), .ZN(new_n19994_));
  AOI21_X1   g19697(.A1(new_n19993_), .A2(new_n19994_), .B(new_n19991_), .ZN(new_n19995_));
  NOR2_X1    g19698(.A1(new_n19990_), .A2(new_n19995_), .ZN(new_n19996_));
  NOR2_X1    g19699(.A1(new_n19750_), .A2(new_n19759_), .ZN(new_n19997_));
  NOR2_X1    g19700(.A1(new_n19997_), .A2(new_n19757_), .ZN(new_n19998_));
  NOR2_X1    g19701(.A1(new_n19996_), .A2(new_n19998_), .ZN(new_n19999_));
  NOR4_X1    g19702(.A1(new_n19990_), .A2(new_n19757_), .A3(new_n19997_), .A4(new_n19995_), .ZN(new_n20000_));
  OAI21_X1   g19703(.A1(new_n19999_), .A2(new_n20000_), .B(new_n19942_), .ZN(new_n20001_));
  XNOR2_X1   g19704(.A1(new_n19996_), .A2(new_n19998_), .ZN(new_n20002_));
  OAI21_X1   g19705(.A1(new_n20002_), .A2(new_n19942_), .B(new_n20001_), .ZN(new_n20003_));
  INV_X1     g19706(.I(new_n20003_), .ZN(new_n20004_));
  NAND2_X1   g19707(.A1(new_n19769_), .A2(new_n19696_), .ZN(new_n20005_));
  NAND2_X1   g19708(.A1(new_n20005_), .A2(new_n19768_), .ZN(new_n20006_));
  OAI22_X1   g19709(.A1(new_n7619_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n8309_), .ZN(new_n20007_));
  OAI21_X1   g19710(.A1(new_n4500_), .A2(new_n7947_), .B(new_n20007_), .ZN(new_n20008_));
  AOI21_X1   g19711(.A1(new_n20008_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n20009_));
  XOR2_X1    g19712(.A1(new_n5067_), .A2(new_n20009_), .Z(new_n20010_));
  XOR2_X1    g19713(.A1(new_n20006_), .A2(new_n20010_), .Z(new_n20011_));
  NOR2_X1    g19714(.A1(new_n20011_), .A2(new_n20004_), .ZN(new_n20012_));
  INV_X1     g19715(.I(new_n20010_), .ZN(new_n20013_));
  NAND2_X1   g19716(.A1(new_n20006_), .A2(new_n20013_), .ZN(new_n20014_));
  NOR2_X1    g19717(.A1(new_n20006_), .A2(new_n20013_), .ZN(new_n20015_));
  INV_X1     g19718(.I(new_n20015_), .ZN(new_n20016_));
  AOI21_X1   g19719(.A1(new_n20016_), .A2(new_n20014_), .B(new_n20003_), .ZN(new_n20017_));
  NOR2_X1    g19720(.A1(new_n20012_), .A2(new_n20017_), .ZN(new_n20018_));
  XOR2_X1    g19721(.A1(new_n20018_), .A2(new_n19937_), .Z(new_n20019_));
  NAND2_X1   g19722(.A1(new_n20019_), .A2(new_n19936_), .ZN(new_n20020_));
  NOR2_X1    g19723(.A1(new_n20018_), .A2(new_n19937_), .ZN(new_n20021_));
  NAND2_X1   g19724(.A1(new_n20018_), .A2(new_n19937_), .ZN(new_n20022_));
  INV_X1     g19725(.I(new_n20022_), .ZN(new_n20023_));
  OAI21_X1   g19726(.A1(new_n20023_), .A2(new_n20021_), .B(new_n19935_), .ZN(new_n20024_));
  NAND2_X1   g19727(.A1(new_n20020_), .A2(new_n20024_), .ZN(new_n20025_));
  INV_X1     g19728(.I(new_n20025_), .ZN(new_n20026_));
  OAI22_X1   g19729(.A1(new_n5993_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n5991_), .ZN(new_n20027_));
  OAI21_X1   g19730(.A1(new_n6229_), .A2(new_n5997_), .B(new_n20027_), .ZN(new_n20028_));
  AOI21_X1   g19731(.A1(new_n20028_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n20029_));
  XOR2_X1    g19732(.A1(new_n6851_), .A2(new_n20029_), .Z(new_n20030_));
  INV_X1     g19733(.I(new_n20030_), .ZN(new_n20031_));
  NAND2_X1   g19734(.A1(new_n20026_), .A2(new_n20031_), .ZN(new_n20032_));
  INV_X1     g19735(.I(new_n20032_), .ZN(new_n20033_));
  NOR2_X1    g19736(.A1(new_n20026_), .A2(new_n20031_), .ZN(new_n20034_));
  OAI21_X1   g19737(.A1(new_n20033_), .A2(new_n20034_), .B(new_n19931_), .ZN(new_n20035_));
  XOR2_X1    g19738(.A1(new_n20025_), .A2(new_n20031_), .Z(new_n20036_));
  OAI21_X1   g19739(.A1(new_n19931_), .A2(new_n20036_), .B(new_n20035_), .ZN(new_n20037_));
  OAI21_X1   g19740(.A1(new_n19691_), .A2(new_n19807_), .B(new_n19805_), .ZN(new_n20038_));
  NAND2_X1   g19741(.A1(new_n20037_), .A2(new_n20038_), .ZN(new_n20039_));
  NOR2_X1    g19742(.A1(new_n20037_), .A2(new_n20038_), .ZN(new_n20040_));
  INV_X1     g19743(.I(new_n20040_), .ZN(new_n20041_));
  AOI21_X1   g19744(.A1(new_n20041_), .A2(new_n20039_), .B(new_n19928_), .ZN(new_n20042_));
  INV_X1     g19745(.I(new_n19928_), .ZN(new_n20043_));
  XNOR2_X1   g19746(.A1(new_n20037_), .A2(new_n20038_), .ZN(new_n20044_));
  NOR2_X1    g19747(.A1(new_n20044_), .A2(new_n20043_), .ZN(new_n20045_));
  NOR2_X1    g19748(.A1(new_n20045_), .A2(new_n20042_), .ZN(new_n20046_));
  INV_X1     g19749(.I(new_n20046_), .ZN(new_n20047_));
  OAI21_X1   g19750(.A1(new_n19594_), .A2(new_n19688_), .B(new_n19818_), .ZN(new_n20048_));
  OAI22_X1   g19751(.A1(new_n4072_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n4067_), .ZN(new_n20049_));
  OAI21_X1   g19752(.A1(new_n8218_), .A2(new_n4318_), .B(new_n20049_), .ZN(new_n20050_));
  AOI21_X1   g19753(.A1(new_n20050_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n20051_));
  XOR2_X1    g19754(.A1(new_n8952_), .A2(new_n20051_), .Z(new_n20052_));
  AOI21_X1   g19755(.A1(new_n20048_), .A2(new_n19817_), .B(new_n20052_), .ZN(new_n20053_));
  NAND2_X1   g19756(.A1(new_n20048_), .A2(new_n19817_), .ZN(new_n20054_));
  INV_X1     g19757(.I(new_n20052_), .ZN(new_n20055_));
  NOR2_X1    g19758(.A1(new_n20054_), .A2(new_n20055_), .ZN(new_n20056_));
  OAI21_X1   g19759(.A1(new_n20056_), .A2(new_n20053_), .B(new_n20047_), .ZN(new_n20057_));
  XOR2_X1    g19760(.A1(new_n20054_), .A2(new_n20052_), .Z(new_n20058_));
  OAI21_X1   g19761(.A1(new_n20058_), .A2(new_n20047_), .B(new_n20057_), .ZN(new_n20059_));
  XNOR2_X1   g19762(.A1(new_n19924_), .A2(new_n20059_), .ZN(new_n20060_));
  NOR2_X1    g19763(.A1(new_n20060_), .A2(new_n19923_), .ZN(new_n20061_));
  NAND2_X1   g19764(.A1(new_n19924_), .A2(new_n20059_), .ZN(new_n20062_));
  NOR2_X1    g19765(.A1(new_n19924_), .A2(new_n20059_), .ZN(new_n20063_));
  INV_X1     g19766(.I(new_n20063_), .ZN(new_n20064_));
  NAND2_X1   g19767(.A1(new_n20064_), .A2(new_n20062_), .ZN(new_n20065_));
  AOI21_X1   g19768(.A1(new_n19923_), .A2(new_n20065_), .B(new_n20061_), .ZN(new_n20066_));
  NOR2_X1    g19769(.A1(new_n20066_), .A2(new_n19919_), .ZN(new_n20067_));
  INV_X1     g19770(.I(new_n20067_), .ZN(new_n20068_));
  NAND2_X1   g19771(.A1(new_n20066_), .A2(new_n19919_), .ZN(new_n20069_));
  AOI21_X1   g19772(.A1(new_n20068_), .A2(new_n20069_), .B(new_n19916_), .ZN(new_n20070_));
  XOR2_X1    g19773(.A1(new_n20066_), .A2(new_n19918_), .Z(new_n20071_));
  INV_X1     g19774(.I(new_n20071_), .ZN(new_n20072_));
  AOI21_X1   g19775(.A1(new_n20072_), .A2(new_n19916_), .B(new_n20070_), .ZN(new_n20073_));
  XNOR2_X1   g19776(.A1(new_n20073_), .A2(new_n19912_), .ZN(new_n20074_));
  NOR2_X1    g19777(.A1(new_n20074_), .A2(new_n19910_), .ZN(new_n20075_));
  INV_X1     g19778(.I(new_n19910_), .ZN(new_n20076_));
  NOR2_X1    g19779(.A1(new_n20073_), .A2(new_n19912_), .ZN(new_n20077_));
  INV_X1     g19780(.I(new_n20077_), .ZN(new_n20078_));
  NAND2_X1   g19781(.A1(new_n20073_), .A2(new_n19912_), .ZN(new_n20079_));
  AOI21_X1   g19782(.A1(new_n20078_), .A2(new_n20079_), .B(new_n20076_), .ZN(new_n20080_));
  NOR2_X1    g19783(.A1(new_n20075_), .A2(new_n20080_), .ZN(new_n20081_));
  NOR3_X1    g19784(.A1(new_n20081_), .A2(new_n19860_), .A3(new_n19906_), .ZN(new_n20082_));
  NOR2_X1    g19785(.A1(new_n19906_), .A2(new_n19860_), .ZN(new_n20083_));
  NOR3_X1    g19786(.A1(new_n20075_), .A2(new_n20083_), .A3(new_n20080_), .ZN(new_n20084_));
  OAI21_X1   g19787(.A1(new_n20082_), .A2(new_n20084_), .B(new_n19905_), .ZN(new_n20085_));
  XOR2_X1    g19788(.A1(new_n20081_), .A2(new_n20083_), .Z(new_n20086_));
  OAI21_X1   g19789(.A1(new_n20086_), .A2(new_n19905_), .B(new_n20085_), .ZN(new_n20087_));
  INV_X1     g19790(.I(new_n20087_), .ZN(new_n20088_));
  NAND2_X1   g19791(.A1(new_n19873_), .A2(new_n19875_), .ZN(new_n20089_));
  NAND2_X1   g19792(.A1(new_n20089_), .A2(new_n19869_), .ZN(new_n20090_));
  XOR2_X1    g19793(.A1(new_n20090_), .A2(new_n20088_), .Z(new_n20091_));
  NOR2_X1    g19794(.A1(new_n20091_), .A2(new_n19900_), .ZN(new_n20092_));
  INV_X1     g19795(.I(new_n19900_), .ZN(new_n20093_));
  INV_X1     g19796(.I(new_n20090_), .ZN(new_n20094_));
  NOR2_X1    g19797(.A1(new_n20094_), .A2(new_n20088_), .ZN(new_n20095_));
  NOR2_X1    g19798(.A1(new_n20090_), .A2(new_n20087_), .ZN(new_n20096_));
  NOR2_X1    g19799(.A1(new_n20095_), .A2(new_n20096_), .ZN(new_n20097_));
  NOR2_X1    g19800(.A1(new_n20097_), .A2(new_n20093_), .ZN(new_n20098_));
  NOR2_X1    g19801(.A1(new_n20098_), .A2(new_n20092_), .ZN(new_n20099_));
  NOR2_X1    g19802(.A1(new_n20099_), .A2(new_n19896_), .ZN(new_n20100_));
  INV_X1     g19803(.I(new_n20100_), .ZN(new_n20101_));
  XOR2_X1    g19804(.A1(new_n19893_), .A2(new_n20101_), .Z(new_n20102_));
  XOR2_X1    g19805(.A1(new_n20102_), .A2(new_n19888_), .Z(\f[82] ));
  NAND2_X1   g19806(.A1(new_n19656_), .A2(new_n19652_), .ZN(new_n20104_));
  OAI21_X1   g19807(.A1(new_n19451_), .A2(new_n19441_), .B(new_n20104_), .ZN(new_n20105_));
  AOI21_X1   g19808(.A1(new_n19896_), .A2(new_n20099_), .B(new_n19888_), .ZN(new_n20106_));
  INV_X1     g19809(.I(new_n20106_), .ZN(new_n20107_));
  OAI21_X1   g19810(.A1(new_n20105_), .A2(new_n20107_), .B(new_n20101_), .ZN(new_n20108_));
  INV_X1     g19811(.I(new_n20096_), .ZN(new_n20109_));
  AOI21_X1   g19812(.A1(new_n20093_), .A2(new_n20109_), .B(new_n20095_), .ZN(new_n20110_));
  INV_X1     g19813(.I(new_n20110_), .ZN(new_n20111_));
  AOI21_X1   g19814(.A1(new_n20076_), .A2(new_n20079_), .B(new_n20077_), .ZN(new_n20112_));
  INV_X1     g19815(.I(new_n20112_), .ZN(new_n20113_));
  OAI22_X1   g19816(.A1(new_n1712_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n1707_), .ZN(new_n20114_));
  OAI21_X1   g19817(.A1(new_n13367_), .A2(new_n1850_), .B(new_n20114_), .ZN(new_n20115_));
  AOI21_X1   g19818(.A1(new_n18183_), .A2(new_n1702_), .B(new_n20115_), .ZN(new_n20116_));
  OAI22_X1   g19819(.A1(new_n2171_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n2166_), .ZN(new_n20117_));
  OAI21_X1   g19820(.A1(new_n12536_), .A2(new_n2322_), .B(new_n20117_), .ZN(new_n20118_));
  AOI21_X1   g19821(.A1(new_n20118_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n20119_));
  XOR2_X1    g19822(.A1(new_n12969_), .A2(new_n20119_), .Z(new_n20120_));
  OAI22_X1   g19823(.A1(new_n11738_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n11744_), .ZN(new_n20121_));
  OAI21_X1   g19824(.A1(new_n10862_), .A2(new_n2884_), .B(new_n20121_), .ZN(new_n20122_));
  AOI21_X1   g19825(.A1(new_n20122_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n20123_));
  XNOR2_X1   g19826(.A1(new_n11748_), .A2(new_n20123_), .ZN(new_n20124_));
  OAI21_X1   g19827(.A1(new_n19923_), .A2(new_n20063_), .B(new_n20062_), .ZN(new_n20125_));
  INV_X1     g19828(.I(new_n20125_), .ZN(new_n20126_));
  OAI22_X1   g19829(.A1(new_n10031_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n10477_), .ZN(new_n20127_));
  OAI21_X1   g19830(.A1(new_n10025_), .A2(new_n3569_), .B(new_n20127_), .ZN(new_n20128_));
  AOI21_X1   g19831(.A1(new_n20128_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n20129_));
  XOR2_X1    g19832(.A1(new_n10476_), .A2(new_n20129_), .Z(new_n20130_));
  OAI22_X1   g19833(.A1(new_n4072_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n4067_), .ZN(new_n20131_));
  OAI21_X1   g19834(.A1(new_n8563_), .A2(new_n4318_), .B(new_n20131_), .ZN(new_n20132_));
  AOI21_X1   g19835(.A1(new_n20132_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n20133_));
  XNOR2_X1   g19836(.A1(new_n9299_), .A2(new_n20133_), .ZN(new_n20134_));
  OAI22_X1   g19837(.A1(new_n5993_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n5991_), .ZN(new_n20135_));
  OAI21_X1   g19838(.A1(new_n6538_), .A2(new_n5997_), .B(new_n20135_), .ZN(new_n20136_));
  AOI21_X1   g19839(.A1(new_n20136_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n20137_));
  XNOR2_X1   g19840(.A1(new_n7202_), .A2(new_n20137_), .ZN(new_n20138_));
  OAI21_X1   g19841(.A1(new_n19935_), .A2(new_n20021_), .B(new_n20022_), .ZN(new_n20139_));
  OAI22_X1   g19842(.A1(new_n6644_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n6647_), .ZN(new_n20140_));
  OAI21_X1   g19843(.A1(new_n5913_), .A2(new_n7284_), .B(new_n20140_), .ZN(new_n20141_));
  AOI21_X1   g19844(.A1(new_n20141_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n20142_));
  XOR2_X1    g19845(.A1(new_n6233_), .A2(new_n20142_), .Z(new_n20143_));
  OAI22_X1   g19846(.A1(new_n7619_), .A2(new_n5068_), .B1(new_n5353_), .B2(new_n8309_), .ZN(new_n20144_));
  OAI21_X1   g19847(.A1(new_n4774_), .A2(new_n7947_), .B(new_n20144_), .ZN(new_n20145_));
  AOI21_X1   g19848(.A1(new_n20145_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n20146_));
  XNOR2_X1   g19849(.A1(new_n5357_), .A2(new_n20146_), .ZN(new_n20147_));
  INV_X1     g19850(.I(new_n20147_), .ZN(new_n20148_));
  INV_X1     g19851(.I(new_n19999_), .ZN(new_n20149_));
  OAI21_X1   g19852(.A1(new_n19941_), .A2(new_n20000_), .B(new_n20149_), .ZN(new_n20150_));
  INV_X1     g19853(.I(new_n20150_), .ZN(new_n20151_));
  OAI22_X1   g19854(.A1(new_n8644_), .A2(new_n4253_), .B1(new_n4500_), .B2(new_n9388_), .ZN(new_n20152_));
  OAI21_X1   g19855(.A1(new_n3989_), .A2(new_n10154_), .B(new_n20152_), .ZN(new_n20153_));
  AOI21_X1   g19856(.A1(new_n20153_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n20154_));
  XOR2_X1    g19857(.A1(new_n4499_), .A2(new_n20154_), .Z(new_n20155_));
  AOI22_X1   g19858(.A1(new_n11415_), .A2(new_n3719_), .B1(\b[30] ), .B2(new_n10145_), .ZN(new_n20156_));
  OAI21_X1   g19859(.A1(new_n20156_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n20157_));
  XNOR2_X1   g19860(.A1(new_n3722_), .A2(new_n20157_), .ZN(new_n20158_));
  AOI22_X1   g19861(.A1(new_n13078_), .A2(\b[24] ), .B1(new_n18773_), .B2(new_n12218_), .ZN(new_n20159_));
  OAI21_X1   g19862(.A1(new_n20159_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n20160_));
  XOR2_X1    g19863(.A1(new_n2443_), .A2(new_n20160_), .Z(new_n20161_));
  NAND2_X1   g19864(.A1(new_n19950_), .A2(new_n19961_), .ZN(new_n20162_));
  NAND2_X1   g19865(.A1(new_n20162_), .A2(new_n19962_), .ZN(new_n20163_));
  OAI22_X1   g19866(.A1(new_n13880_), .A2(new_n2096_), .B1(new_n1634_), .B2(new_n13885_), .ZN(new_n20164_));
  AOI21_X1   g19867(.A1(new_n20164_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n20165_));
  XNOR2_X1   g19868(.A1(new_n1940_), .A2(new_n20165_), .ZN(new_n20166_));
  NOR2_X1    g19869(.A1(new_n13476_), .A2(new_n1518_), .ZN(new_n20167_));
  XOR2_X1    g19870(.A1(new_n14736_), .A2(new_n1518_), .Z(new_n20168_));
  NAND2_X1   g19871(.A1(new_n20168_), .A2(\b[20] ), .ZN(new_n20169_));
  XOR2_X1    g19872(.A1(new_n20169_), .A2(new_n20167_), .Z(new_n20170_));
  XOR2_X1    g19873(.A1(new_n19956_), .A2(new_n20170_), .Z(new_n20171_));
  OR2_X2     g19874(.A1(new_n20166_), .A2(new_n20171_), .Z(new_n20172_));
  NOR2_X1    g19875(.A1(new_n19957_), .A2(new_n20170_), .ZN(new_n20173_));
  INV_X1     g19876(.I(new_n20170_), .ZN(new_n20174_));
  NOR2_X1    g19877(.A1(new_n20174_), .A2(new_n19956_), .ZN(new_n20175_));
  OAI21_X1   g19878(.A1(new_n20173_), .A2(new_n20175_), .B(new_n20166_), .ZN(new_n20176_));
  NAND2_X1   g19879(.A1(new_n20172_), .A2(new_n20176_), .ZN(new_n20177_));
  XOR2_X1    g19880(.A1(new_n20163_), .A2(new_n20177_), .Z(new_n20178_));
  NAND3_X1   g19881(.A1(new_n20177_), .A2(new_n19962_), .A3(new_n20162_), .ZN(new_n20179_));
  NAND3_X1   g19882(.A1(new_n20163_), .A2(new_n20172_), .A3(new_n20176_), .ZN(new_n20180_));
  NAND2_X1   g19883(.A1(new_n20180_), .A2(new_n20179_), .ZN(new_n20181_));
  NAND2_X1   g19884(.A1(new_n20181_), .A2(new_n20161_), .ZN(new_n20182_));
  OAI21_X1   g19885(.A1(new_n20161_), .A2(new_n20178_), .B(new_n20182_), .ZN(new_n20183_));
  AOI22_X1   g19886(.A1(new_n10969_), .A2(new_n3256_), .B1(new_n11394_), .B2(\b[27] ), .ZN(new_n20184_));
  OAI21_X1   g19887(.A1(new_n20184_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n20185_));
  XNOR2_X1   g19888(.A1(new_n3022_), .A2(new_n20185_), .ZN(new_n20186_));
  AOI21_X1   g19889(.A1(new_n19964_), .A2(new_n19974_), .B(new_n19972_), .ZN(new_n20187_));
  INV_X1     g19890(.I(new_n20187_), .ZN(new_n20188_));
  XOR2_X1    g19891(.A1(new_n20186_), .A2(new_n20188_), .Z(new_n20189_));
  AND2_X2    g19892(.A1(new_n20186_), .A2(new_n20188_), .Z(new_n20190_));
  NOR2_X1    g19893(.A1(new_n20186_), .A2(new_n20188_), .ZN(new_n20191_));
  NOR2_X1    g19894(.A1(new_n20190_), .A2(new_n20191_), .ZN(new_n20192_));
  NOR2_X1    g19895(.A1(new_n20192_), .A2(new_n20183_), .ZN(new_n20193_));
  AOI21_X1   g19896(.A1(new_n20183_), .A2(new_n20189_), .B(new_n20193_), .ZN(new_n20194_));
  AOI21_X1   g19897(.A1(new_n19979_), .A2(new_n19982_), .B(new_n19980_), .ZN(new_n20195_));
  NOR2_X1    g19898(.A1(new_n20194_), .A2(new_n20195_), .ZN(new_n20196_));
  INV_X1     g19899(.I(new_n20196_), .ZN(new_n20197_));
  NAND2_X1   g19900(.A1(new_n20194_), .A2(new_n20195_), .ZN(new_n20198_));
  AOI21_X1   g19901(.A1(new_n20197_), .A2(new_n20198_), .B(new_n20158_), .ZN(new_n20199_));
  INV_X1     g19902(.I(new_n20158_), .ZN(new_n20200_));
  XNOR2_X1   g19903(.A1(new_n20194_), .A2(new_n20195_), .ZN(new_n20201_));
  NOR2_X1    g19904(.A1(new_n20201_), .A2(new_n20200_), .ZN(new_n20202_));
  NOR2_X1    g19905(.A1(new_n20202_), .A2(new_n20199_), .ZN(new_n20203_));
  AOI21_X1   g19906(.A1(new_n19984_), .A2(new_n19994_), .B(new_n19992_), .ZN(new_n20204_));
  INV_X1     g19907(.I(new_n20204_), .ZN(new_n20205_));
  XOR2_X1    g19908(.A1(new_n20203_), .A2(new_n20205_), .Z(new_n20206_));
  NOR2_X1    g19909(.A1(new_n20203_), .A2(new_n20204_), .ZN(new_n20207_));
  NOR3_X1    g19910(.A1(new_n20202_), .A2(new_n20199_), .A3(new_n20205_), .ZN(new_n20208_));
  OAI21_X1   g19911(.A1(new_n20207_), .A2(new_n20208_), .B(new_n20155_), .ZN(new_n20209_));
  OAI21_X1   g19912(.A1(new_n20206_), .A2(new_n20155_), .B(new_n20209_), .ZN(new_n20210_));
  XOR2_X1    g19913(.A1(new_n20210_), .A2(new_n20151_), .Z(new_n20211_));
  NAND2_X1   g19914(.A1(new_n20211_), .A2(new_n20148_), .ZN(new_n20212_));
  NAND2_X1   g19915(.A1(new_n20210_), .A2(new_n20151_), .ZN(new_n20213_));
  OR2_X2     g19916(.A1(new_n20210_), .A2(new_n20151_), .Z(new_n20214_));
  NAND2_X1   g19917(.A1(new_n20214_), .A2(new_n20213_), .ZN(new_n20215_));
  NAND2_X1   g19918(.A1(new_n20215_), .A2(new_n20147_), .ZN(new_n20216_));
  NAND2_X1   g19919(.A1(new_n20216_), .A2(new_n20212_), .ZN(new_n20217_));
  OAI21_X1   g19920(.A1(new_n20004_), .A2(new_n20015_), .B(new_n20014_), .ZN(new_n20218_));
  XOR2_X1    g19921(.A1(new_n20217_), .A2(new_n20218_), .Z(new_n20219_));
  NOR2_X1    g19922(.A1(new_n20219_), .A2(new_n20143_), .ZN(new_n20220_));
  INV_X1     g19923(.I(new_n20143_), .ZN(new_n20221_));
  INV_X1     g19924(.I(new_n20218_), .ZN(new_n20222_));
  NOR2_X1    g19925(.A1(new_n20217_), .A2(new_n20222_), .ZN(new_n20223_));
  INV_X1     g19926(.I(new_n20223_), .ZN(new_n20224_));
  NAND2_X1   g19927(.A1(new_n20217_), .A2(new_n20222_), .ZN(new_n20225_));
  AOI21_X1   g19928(.A1(new_n20224_), .A2(new_n20225_), .B(new_n20221_), .ZN(new_n20226_));
  NOR2_X1    g19929(.A1(new_n20220_), .A2(new_n20226_), .ZN(new_n20227_));
  XNOR2_X1   g19930(.A1(new_n20227_), .A2(new_n20139_), .ZN(new_n20228_));
  NOR2_X1    g19931(.A1(new_n20227_), .A2(new_n20139_), .ZN(new_n20229_));
  NAND2_X1   g19932(.A1(new_n20227_), .A2(new_n20139_), .ZN(new_n20230_));
  INV_X1     g19933(.I(new_n20230_), .ZN(new_n20231_));
  OAI21_X1   g19934(.A1(new_n20231_), .A2(new_n20229_), .B(new_n20138_), .ZN(new_n20232_));
  OAI21_X1   g19935(.A1(new_n20138_), .A2(new_n20228_), .B(new_n20232_), .ZN(new_n20233_));
  OAI22_X1   g19936(.A1(new_n5420_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n5107_), .ZN(new_n20234_));
  OAI21_X1   g19937(.A1(new_n7864_), .A2(new_n5112_), .B(new_n20234_), .ZN(new_n20235_));
  AOI21_X1   g19938(.A1(new_n20235_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n20236_));
  XOR2_X1    g19939(.A1(new_n8217_), .A2(new_n20236_), .Z(new_n20237_));
  INV_X1     g19940(.I(new_n20237_), .ZN(new_n20238_));
  OAI21_X1   g19941(.A1(new_n19930_), .A2(new_n20034_), .B(new_n20032_), .ZN(new_n20239_));
  XOR2_X1    g19942(.A1(new_n20239_), .A2(new_n20238_), .Z(new_n20240_));
  NAND2_X1   g19943(.A1(new_n20239_), .A2(new_n20238_), .ZN(new_n20241_));
  NOR2_X1    g19944(.A1(new_n20239_), .A2(new_n20238_), .ZN(new_n20242_));
  INV_X1     g19945(.I(new_n20242_), .ZN(new_n20243_));
  AOI21_X1   g19946(.A1(new_n20241_), .A2(new_n20243_), .B(new_n20233_), .ZN(new_n20244_));
  AOI21_X1   g19947(.A1(new_n20233_), .A2(new_n20240_), .B(new_n20244_), .ZN(new_n20245_));
  OAI21_X1   g19948(.A1(new_n19928_), .A2(new_n20040_), .B(new_n20039_), .ZN(new_n20246_));
  XOR2_X1    g19949(.A1(new_n20245_), .A2(new_n20246_), .Z(new_n20247_));
  INV_X1     g19950(.I(new_n20246_), .ZN(new_n20248_));
  NOR2_X1    g19951(.A1(new_n20245_), .A2(new_n20248_), .ZN(new_n20249_));
  NAND2_X1   g19952(.A1(new_n20245_), .A2(new_n20248_), .ZN(new_n20250_));
  INV_X1     g19953(.I(new_n20250_), .ZN(new_n20251_));
  OAI21_X1   g19954(.A1(new_n20251_), .A2(new_n20249_), .B(new_n20134_), .ZN(new_n20252_));
  OAI21_X1   g19955(.A1(new_n20134_), .A2(new_n20247_), .B(new_n20252_), .ZN(new_n20253_));
  NOR2_X1    g19956(.A1(new_n20056_), .A2(new_n20046_), .ZN(new_n20254_));
  NOR2_X1    g19957(.A1(new_n20254_), .A2(new_n20053_), .ZN(new_n20255_));
  NOR2_X1    g19958(.A1(new_n20253_), .A2(new_n20255_), .ZN(new_n20256_));
  INV_X1     g19959(.I(new_n20256_), .ZN(new_n20257_));
  NAND2_X1   g19960(.A1(new_n20253_), .A2(new_n20255_), .ZN(new_n20258_));
  AOI21_X1   g19961(.A1(new_n20257_), .A2(new_n20258_), .B(new_n20130_), .ZN(new_n20259_));
  INV_X1     g19962(.I(new_n20130_), .ZN(new_n20260_));
  XNOR2_X1   g19963(.A1(new_n20253_), .A2(new_n20255_), .ZN(new_n20261_));
  NOR2_X1    g19964(.A1(new_n20261_), .A2(new_n20260_), .ZN(new_n20262_));
  NOR2_X1    g19965(.A1(new_n20262_), .A2(new_n20259_), .ZN(new_n20263_));
  NOR2_X1    g19966(.A1(new_n20263_), .A2(new_n20126_), .ZN(new_n20264_));
  INV_X1     g19967(.I(new_n20264_), .ZN(new_n20265_));
  NAND2_X1   g19968(.A1(new_n20263_), .A2(new_n20126_), .ZN(new_n20266_));
  AOI21_X1   g19969(.A1(new_n20265_), .A2(new_n20266_), .B(new_n20124_), .ZN(new_n20267_));
  INV_X1     g19970(.I(new_n20124_), .ZN(new_n20268_));
  XOR2_X1    g19971(.A1(new_n20263_), .A2(new_n20125_), .Z(new_n20269_));
  NOR2_X1    g19972(.A1(new_n20269_), .A2(new_n20268_), .ZN(new_n20270_));
  NOR2_X1    g19973(.A1(new_n20270_), .A2(new_n20267_), .ZN(new_n20271_));
  OAI21_X1   g19974(.A1(new_n19916_), .A2(new_n20067_), .B(new_n20069_), .ZN(new_n20272_));
  INV_X1     g19975(.I(new_n20272_), .ZN(new_n20273_));
  NOR2_X1    g19976(.A1(new_n20271_), .A2(new_n20273_), .ZN(new_n20274_));
  INV_X1     g19977(.I(new_n20274_), .ZN(new_n20275_));
  NAND2_X1   g19978(.A1(new_n20271_), .A2(new_n20273_), .ZN(new_n20276_));
  AOI21_X1   g19979(.A1(new_n20275_), .A2(new_n20276_), .B(new_n20120_), .ZN(new_n20277_));
  INV_X1     g19980(.I(new_n20120_), .ZN(new_n20278_));
  XOR2_X1    g19981(.A1(new_n20271_), .A2(new_n20272_), .Z(new_n20279_));
  NOR2_X1    g19982(.A1(new_n20279_), .A2(new_n20278_), .ZN(new_n20280_));
  NOR2_X1    g19983(.A1(new_n20280_), .A2(new_n20277_), .ZN(new_n20281_));
  XOR2_X1    g19984(.A1(new_n20281_), .A2(new_n20116_), .Z(new_n20282_));
  XOR2_X1    g19985(.A1(new_n20282_), .A2(new_n20113_), .Z(new_n20283_));
  XOR2_X1    g19986(.A1(new_n20283_), .A2(\a[23] ), .Z(new_n20284_));
  OAI21_X1   g19987(.A1(new_n1347_), .A2(new_n1457_), .B(new_n16487_), .ZN(new_n20285_));
  NOR2_X1    g19988(.A1(new_n20082_), .A2(new_n19904_), .ZN(new_n20286_));
  NOR2_X1    g19989(.A1(new_n20286_), .A2(new_n20084_), .ZN(new_n20287_));
  XNOR2_X1   g19990(.A1(new_n20287_), .A2(new_n20285_), .ZN(new_n20288_));
  XOR2_X1    g19991(.A1(new_n20284_), .A2(new_n20288_), .Z(new_n20289_));
  NOR2_X1    g19992(.A1(new_n20289_), .A2(\a[20] ), .ZN(new_n20290_));
  NAND2_X1   g19993(.A1(new_n20289_), .A2(\a[20] ), .ZN(new_n20291_));
  INV_X1     g19994(.I(new_n20291_), .ZN(new_n20292_));
  OAI21_X1   g19995(.A1(new_n20292_), .A2(new_n20290_), .B(new_n20111_), .ZN(new_n20293_));
  NOR2_X1    g19996(.A1(new_n20292_), .A2(new_n20290_), .ZN(new_n20294_));
  NAND2_X1   g19997(.A1(new_n20294_), .A2(new_n20110_), .ZN(new_n20295_));
  NAND2_X1   g19998(.A1(new_n20295_), .A2(new_n20293_), .ZN(new_n20296_));
  NAND2_X1   g19999(.A1(new_n20108_), .A2(new_n20296_), .ZN(new_n20297_));
  AOI21_X1   g20000(.A1(new_n19893_), .A2(new_n20106_), .B(new_n20100_), .ZN(new_n20298_));
  XOR2_X1    g20001(.A1(new_n20294_), .A2(new_n20110_), .Z(new_n20299_));
  NAND2_X1   g20002(.A1(new_n20298_), .A2(new_n20299_), .ZN(new_n20300_));
  NAND2_X1   g20003(.A1(new_n20297_), .A2(new_n20300_), .ZN(\f[83] ));
  NAND2_X1   g20004(.A1(new_n20281_), .A2(new_n20112_), .ZN(new_n20302_));
  XOR2_X1    g20005(.A1(new_n20116_), .A2(\a[23] ), .Z(new_n20303_));
  NAND2_X1   g20006(.A1(new_n20302_), .A2(new_n20303_), .ZN(new_n20304_));
  OAI21_X1   g20007(.A1(new_n20112_), .A2(new_n20281_), .B(new_n20304_), .ZN(new_n20305_));
  OAI22_X1   g20008(.A1(new_n1712_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n1707_), .ZN(new_n20306_));
  OAI21_X1   g20009(.A1(new_n13785_), .A2(new_n1850_), .B(new_n20306_), .ZN(new_n20307_));
  AOI21_X1   g20010(.A1(new_n20307_), .A2(new_n1709_), .B(new_n1712_), .ZN(new_n20308_));
  XNOR2_X1   g20011(.A1(new_n14599_), .A2(new_n20308_), .ZN(new_n20309_));
  INV_X1     g20012(.I(new_n20309_), .ZN(new_n20310_));
  OAI22_X1   g20013(.A1(new_n2171_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n2166_), .ZN(new_n20311_));
  OAI21_X1   g20014(.A1(new_n12542_), .A2(new_n2322_), .B(new_n20311_), .ZN(new_n20312_));
  AOI21_X1   g20015(.A1(new_n20312_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n20313_));
  XNOR2_X1   g20016(.A1(new_n13371_), .A2(new_n20313_), .ZN(new_n20314_));
  NAND2_X1   g20017(.A1(new_n20276_), .A2(new_n20278_), .ZN(new_n20315_));
  NAND2_X1   g20018(.A1(new_n20315_), .A2(new_n20275_), .ZN(new_n20316_));
  AOI21_X1   g20019(.A1(new_n20268_), .A2(new_n20266_), .B(new_n20264_), .ZN(new_n20317_));
  OAI22_X1   g20020(.A1(new_n11744_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n12536_), .ZN(new_n20318_));
  OAI21_X1   g20021(.A1(new_n11738_), .A2(new_n2884_), .B(new_n20318_), .ZN(new_n20319_));
  AOI21_X1   g20022(.A1(new_n20319_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n20320_));
  XNOR2_X1   g20023(.A1(new_n12128_), .A2(new_n20320_), .ZN(new_n20321_));
  INV_X1     g20024(.I(new_n20321_), .ZN(new_n20322_));
  OAI22_X1   g20025(.A1(new_n10477_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n10862_), .ZN(new_n20323_));
  OAI21_X1   g20026(.A1(new_n10031_), .A2(new_n3569_), .B(new_n20323_), .ZN(new_n20324_));
  AOI21_X1   g20027(.A1(new_n20324_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n20325_));
  XNOR2_X1   g20028(.A1(new_n10866_), .A2(new_n20325_), .ZN(new_n20326_));
  INV_X1     g20029(.I(new_n20326_), .ZN(new_n20327_));
  NAND2_X1   g20030(.A1(new_n20258_), .A2(new_n20260_), .ZN(new_n20328_));
  NAND2_X1   g20031(.A1(new_n20328_), .A2(new_n20257_), .ZN(new_n20329_));
  NOR2_X1    g20032(.A1(new_n20251_), .A2(new_n20134_), .ZN(new_n20330_));
  OAI21_X1   g20033(.A1(new_n20138_), .A2(new_n20229_), .B(new_n20230_), .ZN(new_n20331_));
  INV_X1     g20034(.I(new_n20214_), .ZN(new_n20332_));
  AOI21_X1   g20035(.A1(new_n20148_), .A2(new_n20213_), .B(new_n20332_), .ZN(new_n20333_));
  NOR2_X1    g20036(.A1(new_n20208_), .A2(new_n20155_), .ZN(new_n20334_));
  NOR2_X1    g20037(.A1(new_n20334_), .A2(new_n20207_), .ZN(new_n20335_));
  AOI21_X1   g20038(.A1(new_n20200_), .A2(new_n20198_), .B(new_n20196_), .ZN(new_n20336_));
  INV_X1     g20039(.I(new_n20161_), .ZN(new_n20337_));
  NAND2_X1   g20040(.A1(new_n20337_), .A2(new_n20179_), .ZN(new_n20338_));
  AND2_X2    g20041(.A1(new_n20338_), .A2(new_n20180_), .Z(new_n20339_));
  OAI22_X1   g20042(.A1(new_n13880_), .A2(new_n2103_), .B1(new_n1803_), .B2(new_n13885_), .ZN(new_n20340_));
  AOI21_X1   g20043(.A1(new_n20340_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n20341_));
  XOR2_X1    g20044(.A1(new_n2106_), .A2(new_n20341_), .Z(new_n20342_));
  NOR2_X1    g20045(.A1(new_n20166_), .A2(new_n20173_), .ZN(new_n20343_));
  NOR2_X1    g20046(.A1(new_n20343_), .A2(new_n20175_), .ZN(new_n20344_));
  INV_X1     g20047(.I(new_n20344_), .ZN(new_n20345_));
  NOR2_X1    g20048(.A1(new_n13476_), .A2(new_n1525_), .ZN(new_n20346_));
  XOR2_X1    g20049(.A1(new_n14736_), .A2(new_n1525_), .Z(new_n20347_));
  NAND2_X1   g20050(.A1(new_n20347_), .A2(\b[21] ), .ZN(new_n20348_));
  XOR2_X1    g20051(.A1(new_n20348_), .A2(new_n20346_), .Z(new_n20349_));
  XOR2_X1    g20052(.A1(new_n20349_), .A2(\a[20] ), .Z(new_n20350_));
  NOR2_X1    g20053(.A1(new_n20350_), .A2(new_n20170_), .ZN(new_n20351_));
  NOR2_X1    g20054(.A1(new_n20349_), .A2(new_n1346_), .ZN(new_n20352_));
  INV_X1     g20055(.I(new_n20352_), .ZN(new_n20353_));
  NAND2_X1   g20056(.A1(new_n20349_), .A2(new_n1346_), .ZN(new_n20354_));
  AOI21_X1   g20057(.A1(new_n20353_), .A2(new_n20354_), .B(new_n20174_), .ZN(new_n20355_));
  NOR2_X1    g20058(.A1(new_n20351_), .A2(new_n20355_), .ZN(new_n20356_));
  NOR2_X1    g20059(.A1(new_n20345_), .A2(new_n20356_), .ZN(new_n20357_));
  INV_X1     g20060(.I(new_n20357_), .ZN(new_n20358_));
  NAND2_X1   g20061(.A1(new_n20345_), .A2(new_n20356_), .ZN(new_n20359_));
  AOI21_X1   g20062(.A1(new_n20358_), .A2(new_n20359_), .B(new_n20342_), .ZN(new_n20360_));
  XOR2_X1    g20063(.A1(new_n20344_), .A2(new_n20356_), .Z(new_n20361_));
  INV_X1     g20064(.I(new_n20361_), .ZN(new_n20362_));
  AOI21_X1   g20065(.A1(new_n20342_), .A2(new_n20362_), .B(new_n20360_), .ZN(new_n20363_));
  AOI22_X1   g20066(.A1(new_n13078_), .A2(\b[25] ), .B1(new_n2838_), .B2(new_n12218_), .ZN(new_n20364_));
  OAI21_X1   g20067(.A1(new_n20364_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n20365_));
  XOR2_X1    g20068(.A1(new_n2647_), .A2(new_n20365_), .Z(new_n20366_));
  XNOR2_X1   g20069(.A1(new_n20363_), .A2(new_n20366_), .ZN(new_n20367_));
  NOR2_X1    g20070(.A1(new_n20367_), .A2(new_n20339_), .ZN(new_n20368_));
  INV_X1     g20071(.I(new_n20339_), .ZN(new_n20369_));
  NOR2_X1    g20072(.A1(new_n20363_), .A2(new_n20366_), .ZN(new_n20370_));
  INV_X1     g20073(.I(new_n20370_), .ZN(new_n20371_));
  NAND2_X1   g20074(.A1(new_n20363_), .A2(new_n20366_), .ZN(new_n20372_));
  AOI21_X1   g20075(.A1(new_n20371_), .A2(new_n20372_), .B(new_n20369_), .ZN(new_n20373_));
  NOR2_X1    g20076(.A1(new_n20368_), .A2(new_n20373_), .ZN(new_n20374_));
  AOI22_X1   g20077(.A1(new_n10969_), .A2(new_n19751_), .B1(new_n11394_), .B2(\b[28] ), .ZN(new_n20375_));
  OAI21_X1   g20078(.A1(new_n20375_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n20376_));
  XOR2_X1    g20079(.A1(new_n3264_), .A2(new_n20376_), .Z(new_n20377_));
  INV_X1     g20080(.I(new_n20190_), .ZN(new_n20378_));
  OAI21_X1   g20081(.A1(new_n20183_), .A2(new_n20191_), .B(new_n20378_), .ZN(new_n20379_));
  INV_X1     g20082(.I(new_n20379_), .ZN(new_n20380_));
  NOR2_X1    g20083(.A1(new_n20380_), .A2(new_n20377_), .ZN(new_n20381_));
  NAND2_X1   g20084(.A1(new_n20380_), .A2(new_n20377_), .ZN(new_n20382_));
  INV_X1     g20085(.I(new_n20382_), .ZN(new_n20383_));
  NOR2_X1    g20086(.A1(new_n20383_), .A2(new_n20381_), .ZN(new_n20384_));
  XNOR2_X1   g20087(.A1(new_n20379_), .A2(new_n20377_), .ZN(new_n20385_));
  NAND2_X1   g20088(.A1(new_n20385_), .A2(new_n20374_), .ZN(new_n20386_));
  OAI21_X1   g20089(.A1(new_n20374_), .A2(new_n20384_), .B(new_n20386_), .ZN(new_n20387_));
  AOI22_X1   g20090(.A1(new_n11415_), .A2(new_n4249_), .B1(\b[31] ), .B2(new_n10145_), .ZN(new_n20388_));
  OAI21_X1   g20091(.A1(new_n20388_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n20389_));
  XOR2_X1    g20092(.A1(new_n3993_), .A2(new_n20389_), .Z(new_n20390_));
  NOR2_X1    g20093(.A1(new_n20387_), .A2(new_n20390_), .ZN(new_n20391_));
  INV_X1     g20094(.I(new_n20391_), .ZN(new_n20392_));
  NAND2_X1   g20095(.A1(new_n20387_), .A2(new_n20390_), .ZN(new_n20393_));
  AOI21_X1   g20096(.A1(new_n20392_), .A2(new_n20393_), .B(new_n20336_), .ZN(new_n20394_));
  INV_X1     g20097(.I(new_n20336_), .ZN(new_n20395_));
  XNOR2_X1   g20098(.A1(new_n20387_), .A2(new_n20390_), .ZN(new_n20396_));
  NOR2_X1    g20099(.A1(new_n20396_), .A2(new_n20395_), .ZN(new_n20397_));
  NOR2_X1    g20100(.A1(new_n20397_), .A2(new_n20394_), .ZN(new_n20398_));
  OAI22_X1   g20101(.A1(new_n8644_), .A2(new_n4500_), .B1(new_n4774_), .B2(new_n9388_), .ZN(new_n20399_));
  OAI21_X1   g20102(.A1(new_n4253_), .A2(new_n10154_), .B(new_n20399_), .ZN(new_n20400_));
  AOI21_X1   g20103(.A1(new_n20400_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n20401_));
  XNOR2_X1   g20104(.A1(new_n4778_), .A2(new_n20401_), .ZN(new_n20402_));
  XNOR2_X1   g20105(.A1(new_n20398_), .A2(new_n20402_), .ZN(new_n20403_));
  NOR2_X1    g20106(.A1(new_n20403_), .A2(new_n20335_), .ZN(new_n20404_));
  INV_X1     g20107(.I(new_n20335_), .ZN(new_n20405_));
  NOR2_X1    g20108(.A1(new_n20398_), .A2(new_n20402_), .ZN(new_n20406_));
  INV_X1     g20109(.I(new_n20406_), .ZN(new_n20407_));
  NAND2_X1   g20110(.A1(new_n20398_), .A2(new_n20402_), .ZN(new_n20408_));
  AOI21_X1   g20111(.A1(new_n20407_), .A2(new_n20408_), .B(new_n20405_), .ZN(new_n20409_));
  NOR2_X1    g20112(.A1(new_n20404_), .A2(new_n20409_), .ZN(new_n20410_));
  OAI22_X1   g20113(.A1(new_n7619_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n8309_), .ZN(new_n20411_));
  OAI21_X1   g20114(.A1(new_n5068_), .A2(new_n7947_), .B(new_n20411_), .ZN(new_n20412_));
  AOI21_X1   g20115(.A1(new_n20412_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n20413_));
  XNOR2_X1   g20116(.A1(new_n5600_), .A2(new_n20413_), .ZN(new_n20414_));
  XOR2_X1    g20117(.A1(new_n20410_), .A2(new_n20414_), .Z(new_n20415_));
  NOR2_X1    g20118(.A1(new_n20415_), .A2(new_n20333_), .ZN(new_n20416_));
  INV_X1     g20119(.I(new_n20333_), .ZN(new_n20417_));
  INV_X1     g20120(.I(new_n20410_), .ZN(new_n20418_));
  NOR2_X1    g20121(.A1(new_n20418_), .A2(new_n20414_), .ZN(new_n20419_));
  INV_X1     g20122(.I(new_n20419_), .ZN(new_n20420_));
  NAND2_X1   g20123(.A1(new_n20418_), .A2(new_n20414_), .ZN(new_n20421_));
  AOI21_X1   g20124(.A1(new_n20420_), .A2(new_n20421_), .B(new_n20417_), .ZN(new_n20422_));
  NOR2_X1    g20125(.A1(new_n20422_), .A2(new_n20416_), .ZN(new_n20423_));
  INV_X1     g20126(.I(new_n20423_), .ZN(new_n20424_));
  OAI22_X1   g20127(.A1(new_n6644_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n6647_), .ZN(new_n20425_));
  OAI21_X1   g20128(.A1(new_n5921_), .A2(new_n7284_), .B(new_n20425_), .ZN(new_n20426_));
  AOI21_X1   g20129(.A1(new_n20426_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n20427_));
  XOR2_X1    g20130(.A1(new_n6543_), .A2(new_n20427_), .Z(new_n20428_));
  NAND2_X1   g20131(.A1(new_n20225_), .A2(new_n20221_), .ZN(new_n20429_));
  AOI21_X1   g20132(.A1(new_n20429_), .A2(new_n20224_), .B(new_n20428_), .ZN(new_n20430_));
  INV_X1     g20133(.I(new_n20428_), .ZN(new_n20431_));
  NAND2_X1   g20134(.A1(new_n20429_), .A2(new_n20224_), .ZN(new_n20432_));
  NOR2_X1    g20135(.A1(new_n20432_), .A2(new_n20431_), .ZN(new_n20433_));
  OAI21_X1   g20136(.A1(new_n20430_), .A2(new_n20433_), .B(new_n20424_), .ZN(new_n20434_));
  XOR2_X1    g20137(.A1(new_n20432_), .A2(new_n20428_), .Z(new_n20435_));
  OAI21_X1   g20138(.A1(new_n20424_), .A2(new_n20435_), .B(new_n20434_), .ZN(new_n20436_));
  AOI22_X1   g20139(.A1(new_n5680_), .A2(\b[44] ), .B1(\b[45] ), .B2(new_n5686_), .ZN(new_n20437_));
  AOI21_X1   g20140(.A1(\b[43] ), .A2(new_n6923_), .B(new_n20437_), .ZN(new_n20438_));
  OAI21_X1   g20141(.A1(new_n20438_), .A2(\a[41] ), .B(new_n5680_), .ZN(new_n20439_));
  XNOR2_X1   g20142(.A1(new_n7516_), .A2(new_n20439_), .ZN(new_n20440_));
  XOR2_X1    g20143(.A1(new_n20436_), .A2(new_n20440_), .Z(new_n20441_));
  AND2_X2    g20144(.A1(new_n20441_), .A2(new_n20331_), .Z(new_n20442_));
  NOR2_X1    g20145(.A1(new_n20436_), .A2(new_n20440_), .ZN(new_n20443_));
  INV_X1     g20146(.I(new_n20443_), .ZN(new_n20444_));
  NAND2_X1   g20147(.A1(new_n20436_), .A2(new_n20440_), .ZN(new_n20445_));
  AOI21_X1   g20148(.A1(new_n20444_), .A2(new_n20445_), .B(new_n20331_), .ZN(new_n20446_));
  NOR2_X1    g20149(.A1(new_n20442_), .A2(new_n20446_), .ZN(new_n20447_));
  AOI22_X1   g20150(.A1(new_n4859_), .A2(\b[47] ), .B1(new_n4865_), .B2(\b[48] ), .ZN(new_n20448_));
  AOI21_X1   g20151(.A1(\b[46] ), .A2(new_n6005_), .B(new_n20448_), .ZN(new_n20449_));
  OAI21_X1   g20152(.A1(new_n20449_), .A2(\a[38] ), .B(new_n4859_), .ZN(new_n20450_));
  XOR2_X1    g20153(.A1(new_n8568_), .A2(new_n20450_), .Z(new_n20451_));
  OAI21_X1   g20154(.A1(new_n20233_), .A2(new_n20242_), .B(new_n20241_), .ZN(new_n20452_));
  NAND2_X1   g20155(.A1(new_n20452_), .A2(new_n20451_), .ZN(new_n20453_));
  NOR2_X1    g20156(.A1(new_n20452_), .A2(new_n20451_), .ZN(new_n20454_));
  INV_X1     g20157(.I(new_n20454_), .ZN(new_n20455_));
  AOI21_X1   g20158(.A1(new_n20455_), .A2(new_n20453_), .B(new_n20447_), .ZN(new_n20456_));
  XNOR2_X1   g20159(.A1(new_n20452_), .A2(new_n20451_), .ZN(new_n20457_));
  NOR3_X1    g20160(.A1(new_n20442_), .A2(new_n20457_), .A3(new_n20446_), .ZN(new_n20458_));
  OAI22_X1   g20161(.A1(new_n4072_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n4067_), .ZN(new_n20459_));
  OAI21_X1   g20162(.A1(new_n8948_), .A2(new_n4318_), .B(new_n20459_), .ZN(new_n20460_));
  AOI21_X1   g20163(.A1(new_n20460_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n20461_));
  XNOR2_X1   g20164(.A1(new_n9642_), .A2(new_n20461_), .ZN(new_n20462_));
  NOR3_X1    g20165(.A1(new_n20456_), .A2(new_n20458_), .A3(new_n20462_), .ZN(new_n20463_));
  NOR2_X1    g20166(.A1(new_n20456_), .A2(new_n20458_), .ZN(new_n20464_));
  INV_X1     g20167(.I(new_n20462_), .ZN(new_n20465_));
  NOR2_X1    g20168(.A1(new_n20464_), .A2(new_n20465_), .ZN(new_n20466_));
  OAI22_X1   g20169(.A1(new_n20466_), .A2(new_n20463_), .B1(new_n20249_), .B2(new_n20330_), .ZN(new_n20467_));
  NOR2_X1    g20170(.A1(new_n20330_), .A2(new_n20249_), .ZN(new_n20468_));
  XOR2_X1    g20171(.A1(new_n20464_), .A2(new_n20465_), .Z(new_n20469_));
  NAND2_X1   g20172(.A1(new_n20469_), .A2(new_n20468_), .ZN(new_n20470_));
  NAND2_X1   g20173(.A1(new_n20470_), .A2(new_n20467_), .ZN(new_n20471_));
  XOR2_X1    g20174(.A1(new_n20471_), .A2(new_n20329_), .Z(new_n20472_));
  NAND2_X1   g20175(.A1(new_n20472_), .A2(new_n20327_), .ZN(new_n20473_));
  AOI22_X1   g20176(.A1(new_n20470_), .A2(new_n20467_), .B1(new_n20257_), .B2(new_n20328_), .ZN(new_n20474_));
  NOR2_X1    g20177(.A1(new_n20471_), .A2(new_n20329_), .ZN(new_n20475_));
  OAI21_X1   g20178(.A1(new_n20475_), .A2(new_n20474_), .B(new_n20326_), .ZN(new_n20476_));
  AOI21_X1   g20179(.A1(new_n20473_), .A2(new_n20476_), .B(new_n20322_), .ZN(new_n20477_));
  NAND2_X1   g20180(.A1(new_n20473_), .A2(new_n20476_), .ZN(new_n20478_));
  NOR2_X1    g20181(.A1(new_n20478_), .A2(new_n20321_), .ZN(new_n20479_));
  NOR2_X1    g20182(.A1(new_n20479_), .A2(new_n20477_), .ZN(new_n20480_));
  NOR2_X1    g20183(.A1(new_n20480_), .A2(new_n20317_), .ZN(new_n20481_));
  INV_X1     g20184(.I(new_n20317_), .ZN(new_n20482_));
  XOR2_X1    g20185(.A1(new_n20478_), .A2(new_n20322_), .Z(new_n20483_));
  NOR2_X1    g20186(.A1(new_n20483_), .A2(new_n20482_), .ZN(new_n20484_));
  NOR2_X1    g20187(.A1(new_n20484_), .A2(new_n20481_), .ZN(new_n20485_));
  XOR2_X1    g20188(.A1(new_n20485_), .A2(new_n20316_), .Z(new_n20486_));
  NOR2_X1    g20189(.A1(new_n20486_), .A2(new_n20314_), .ZN(new_n20487_));
  INV_X1     g20190(.I(new_n20314_), .ZN(new_n20488_));
  INV_X1     g20191(.I(new_n20316_), .ZN(new_n20489_));
  NOR2_X1    g20192(.A1(new_n20485_), .A2(new_n20489_), .ZN(new_n20490_));
  INV_X1     g20193(.I(new_n20490_), .ZN(new_n20491_));
  NAND2_X1   g20194(.A1(new_n20485_), .A2(new_n20489_), .ZN(new_n20492_));
  AOI21_X1   g20195(.A1(new_n20491_), .A2(new_n20492_), .B(new_n20488_), .ZN(new_n20493_));
  NOR2_X1    g20196(.A1(new_n20487_), .A2(new_n20493_), .ZN(new_n20494_));
  NOR2_X1    g20197(.A1(new_n20494_), .A2(new_n20310_), .ZN(new_n20495_));
  INV_X1     g20198(.I(new_n20495_), .ZN(new_n20496_));
  NAND2_X1   g20199(.A1(new_n20494_), .A2(new_n20310_), .ZN(new_n20497_));
  NAND2_X1   g20200(.A1(new_n20496_), .A2(new_n20497_), .ZN(new_n20498_));
  XOR2_X1    g20201(.A1(new_n20494_), .A2(new_n20309_), .Z(new_n20499_));
  NOR2_X1    g20202(.A1(new_n20499_), .A2(new_n20305_), .ZN(new_n20500_));
  AOI21_X1   g20203(.A1(new_n20305_), .A2(new_n20498_), .B(new_n20500_), .ZN(new_n20501_));
  NOR2_X1    g20204(.A1(new_n20284_), .A2(new_n20287_), .ZN(new_n20502_));
  XOR2_X1    g20205(.A1(new_n20285_), .A2(new_n1346_), .Z(new_n20503_));
  AOI21_X1   g20206(.A1(new_n20284_), .A2(new_n20287_), .B(new_n20503_), .ZN(new_n20504_));
  NOR2_X1    g20207(.A1(new_n20504_), .A2(new_n20502_), .ZN(new_n20505_));
  XNOR2_X1   g20208(.A1(new_n20505_), .A2(new_n20501_), .ZN(new_n20506_));
  INV_X1     g20209(.I(new_n20506_), .ZN(new_n20507_));
  NAND2_X1   g20210(.A1(new_n20299_), .A2(new_n20507_), .ZN(new_n20508_));
  XNOR2_X1   g20211(.A1(new_n20508_), .A2(new_n20293_), .ZN(new_n20509_));
  XOR2_X1    g20212(.A1(new_n20298_), .A2(new_n20509_), .Z(\f[84] ));
  NAND2_X1   g20213(.A1(new_n20505_), .A2(new_n20501_), .ZN(new_n20511_));
  NAND2_X1   g20214(.A1(new_n20294_), .A2(new_n20506_), .ZN(new_n20512_));
  NOR2_X1    g20215(.A1(new_n20294_), .A2(new_n20506_), .ZN(new_n20513_));
  OAI21_X1   g20216(.A1(new_n20111_), .A2(new_n20513_), .B(new_n20512_), .ZN(new_n20514_));
  INV_X1     g20217(.I(new_n20514_), .ZN(new_n20515_));
  NAND2_X1   g20218(.A1(new_n20108_), .A2(new_n20515_), .ZN(new_n20516_));
  NOR2_X1    g20219(.A1(new_n1850_), .A2(new_n1707_), .ZN(new_n20517_));
  NAND2_X1   g20220(.A1(new_n16148_), .A2(new_n1709_), .ZN(new_n20518_));
  OAI21_X1   g20221(.A1(new_n20517_), .A2(new_n20518_), .B(new_n1702_), .ZN(new_n20519_));
  XNOR2_X1   g20222(.A1(new_n14978_), .A2(new_n20519_), .ZN(new_n20520_));
  NAND2_X1   g20223(.A1(new_n20492_), .A2(new_n20488_), .ZN(new_n20521_));
  NAND2_X1   g20224(.A1(new_n20521_), .A2(new_n20491_), .ZN(new_n20522_));
  INV_X1     g20225(.I(new_n20522_), .ZN(new_n20523_));
  OAI22_X1   g20226(.A1(new_n2171_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n2166_), .ZN(new_n20524_));
  OAI21_X1   g20227(.A1(new_n12970_), .A2(new_n2322_), .B(new_n20524_), .ZN(new_n20525_));
  AOI21_X1   g20228(.A1(new_n20525_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n20526_));
  XOR2_X1    g20229(.A1(new_n13784_), .A2(new_n20526_), .Z(new_n20527_));
  INV_X1     g20230(.I(new_n20477_), .ZN(new_n20528_));
  AOI21_X1   g20231(.A1(new_n20528_), .A2(new_n20482_), .B(new_n20479_), .ZN(new_n20529_));
  OAI22_X1   g20232(.A1(new_n12536_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n12542_), .ZN(new_n20530_));
  OAI21_X1   g20233(.A1(new_n11744_), .A2(new_n2884_), .B(new_n20530_), .ZN(new_n20531_));
  AOI21_X1   g20234(.A1(new_n20531_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n20532_));
  XNOR2_X1   g20235(.A1(new_n12546_), .A2(new_n20532_), .ZN(new_n20533_));
  NOR2_X1    g20236(.A1(new_n20475_), .A2(new_n20326_), .ZN(new_n20534_));
  NOR2_X1    g20237(.A1(new_n20466_), .A2(new_n20468_), .ZN(new_n20535_));
  NOR2_X1    g20238(.A1(new_n20535_), .A2(new_n20463_), .ZN(new_n20536_));
  OAI22_X1   g20239(.A1(new_n10862_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n11738_), .ZN(new_n20537_));
  OAI21_X1   g20240(.A1(new_n10477_), .A2(new_n3569_), .B(new_n20537_), .ZN(new_n20538_));
  AOI21_X1   g20241(.A1(new_n20538_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n20539_));
  XOR2_X1    g20242(.A1(new_n11298_), .A2(new_n20539_), .Z(new_n20540_));
  OAI22_X1   g20243(.A1(new_n4072_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n4067_), .ZN(new_n20541_));
  OAI21_X1   g20244(.A1(new_n9295_), .A2(new_n4318_), .B(new_n20541_), .ZN(new_n20542_));
  AOI21_X1   g20245(.A1(new_n20542_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n20543_));
  XNOR2_X1   g20246(.A1(new_n10035_), .A2(new_n20543_), .ZN(new_n20544_));
  INV_X1     g20247(.I(new_n20544_), .ZN(new_n20545_));
  OAI22_X1   g20248(.A1(new_n5993_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n5991_), .ZN(new_n20546_));
  OAI21_X1   g20249(.A1(new_n7198_), .A2(new_n5997_), .B(new_n20546_), .ZN(new_n20547_));
  AOI21_X1   g20250(.A1(new_n20547_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n20548_));
  XNOR2_X1   g20251(.A1(new_n7874_), .A2(new_n20548_), .ZN(new_n20549_));
  AOI21_X1   g20252(.A1(new_n20417_), .A2(new_n20421_), .B(new_n20419_), .ZN(new_n20550_));
  OAI22_X1   g20253(.A1(new_n7619_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n8309_), .ZN(new_n20551_));
  OAI21_X1   g20254(.A1(new_n5353_), .A2(new_n7947_), .B(new_n20551_), .ZN(new_n20552_));
  AOI21_X1   g20255(.A1(new_n20552_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n20553_));
  XOR2_X1    g20256(.A1(new_n5926_), .A2(new_n20553_), .Z(new_n20554_));
  AOI21_X1   g20257(.A1(new_n20405_), .A2(new_n20408_), .B(new_n20406_), .ZN(new_n20555_));
  INV_X1     g20258(.I(new_n4254_), .ZN(new_n20556_));
  AOI22_X1   g20259(.A1(new_n11415_), .A2(new_n20556_), .B1(\b[32] ), .B2(new_n10145_), .ZN(new_n20557_));
  OAI21_X1   g20260(.A1(new_n20557_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n20558_));
  XOR2_X1    g20261(.A1(new_n4257_), .A2(new_n20558_), .Z(new_n20559_));
  INV_X1     g20262(.I(new_n20559_), .ZN(new_n20560_));
  AOI21_X1   g20263(.A1(new_n20369_), .A2(new_n20372_), .B(new_n20370_), .ZN(new_n20561_));
  AOI22_X1   g20264(.A1(new_n13078_), .A2(\b[26] ), .B1(new_n19278_), .B2(new_n12218_), .ZN(new_n20562_));
  OAI21_X1   g20265(.A1(new_n20562_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n20563_));
  XOR2_X1    g20266(.A1(new_n2846_), .A2(new_n20563_), .Z(new_n20564_));
  OAI21_X1   g20267(.A1(new_n20342_), .A2(new_n20357_), .B(new_n20359_), .ZN(new_n20565_));
  OAI22_X1   g20268(.A1(new_n13880_), .A2(new_n2434_), .B1(new_n1936_), .B2(new_n13885_), .ZN(new_n20566_));
  AOI21_X1   g20269(.A1(new_n20566_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n20567_));
  XNOR2_X1   g20270(.A1(new_n2280_), .A2(new_n20567_), .ZN(new_n20568_));
  NAND2_X1   g20271(.A1(new_n20354_), .A2(new_n20174_), .ZN(new_n20569_));
  NAND2_X1   g20272(.A1(new_n20569_), .A2(new_n20353_), .ZN(new_n20570_));
  NOR2_X1    g20273(.A1(new_n13476_), .A2(new_n1634_), .ZN(new_n20571_));
  XOR2_X1    g20274(.A1(new_n14736_), .A2(new_n1634_), .Z(new_n20572_));
  NAND2_X1   g20275(.A1(new_n20572_), .A2(\b[22] ), .ZN(new_n20573_));
  XOR2_X1    g20276(.A1(new_n20573_), .A2(new_n20571_), .Z(new_n20574_));
  INV_X1     g20277(.I(new_n20574_), .ZN(new_n20575_));
  XOR2_X1    g20278(.A1(new_n20570_), .A2(new_n20575_), .Z(new_n20576_));
  OR2_X2     g20279(.A1(new_n20568_), .A2(new_n20576_), .Z(new_n20577_));
  NOR2_X1    g20280(.A1(new_n20570_), .A2(new_n20574_), .ZN(new_n20578_));
  NAND2_X1   g20281(.A1(new_n20570_), .A2(new_n20574_), .ZN(new_n20579_));
  INV_X1     g20282(.I(new_n20579_), .ZN(new_n20580_));
  OAI21_X1   g20283(.A1(new_n20578_), .A2(new_n20580_), .B(new_n20568_), .ZN(new_n20581_));
  NAND2_X1   g20284(.A1(new_n20577_), .A2(new_n20581_), .ZN(new_n20582_));
  XOR2_X1    g20285(.A1(new_n20565_), .A2(new_n20582_), .Z(new_n20583_));
  INV_X1     g20286(.I(new_n20565_), .ZN(new_n20584_));
  NAND2_X1   g20287(.A1(new_n20584_), .A2(new_n20582_), .ZN(new_n20585_));
  NOR2_X1    g20288(.A1(new_n20584_), .A2(new_n20582_), .ZN(new_n20586_));
  INV_X1     g20289(.I(new_n20586_), .ZN(new_n20587_));
  NAND2_X1   g20290(.A1(new_n20587_), .A2(new_n20585_), .ZN(new_n20588_));
  NAND2_X1   g20291(.A1(new_n20588_), .A2(new_n20564_), .ZN(new_n20589_));
  OAI21_X1   g20292(.A1(new_n20564_), .A2(new_n20583_), .B(new_n20589_), .ZN(new_n20590_));
  AOI22_X1   g20293(.A1(new_n10969_), .A2(new_n3711_), .B1(new_n11394_), .B2(\b[29] ), .ZN(new_n20591_));
  OAI21_X1   g20294(.A1(new_n20591_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n20592_));
  XOR2_X1    g20295(.A1(new_n3514_), .A2(new_n20592_), .Z(new_n20593_));
  NOR2_X1    g20296(.A1(new_n20590_), .A2(new_n20593_), .ZN(new_n20594_));
  INV_X1     g20297(.I(new_n20594_), .ZN(new_n20595_));
  NAND2_X1   g20298(.A1(new_n20590_), .A2(new_n20593_), .ZN(new_n20596_));
  AOI21_X1   g20299(.A1(new_n20595_), .A2(new_n20596_), .B(new_n20561_), .ZN(new_n20597_));
  INV_X1     g20300(.I(new_n20561_), .ZN(new_n20598_));
  XNOR2_X1   g20301(.A1(new_n20590_), .A2(new_n20593_), .ZN(new_n20599_));
  NOR2_X1    g20302(.A1(new_n20599_), .A2(new_n20598_), .ZN(new_n20600_));
  NOR2_X1    g20303(.A1(new_n20600_), .A2(new_n20597_), .ZN(new_n20601_));
  AOI21_X1   g20304(.A1(new_n20374_), .A2(new_n20382_), .B(new_n20381_), .ZN(new_n20602_));
  NOR2_X1    g20305(.A1(new_n20601_), .A2(new_n20602_), .ZN(new_n20603_));
  NAND2_X1   g20306(.A1(new_n20601_), .A2(new_n20602_), .ZN(new_n20604_));
  INV_X1     g20307(.I(new_n20604_), .ZN(new_n20605_));
  OAI21_X1   g20308(.A1(new_n20605_), .A2(new_n20603_), .B(new_n20560_), .ZN(new_n20606_));
  XNOR2_X1   g20309(.A1(new_n20601_), .A2(new_n20602_), .ZN(new_n20607_));
  OAI21_X1   g20310(.A1(new_n20560_), .A2(new_n20607_), .B(new_n20606_), .ZN(new_n20608_));
  NAND2_X1   g20311(.A1(new_n20393_), .A2(new_n20395_), .ZN(new_n20609_));
  NAND2_X1   g20312(.A1(new_n20609_), .A2(new_n20392_), .ZN(new_n20610_));
  OAI22_X1   g20313(.A1(new_n8644_), .A2(new_n4774_), .B1(new_n5068_), .B2(new_n9388_), .ZN(new_n20611_));
  OAI21_X1   g20314(.A1(new_n4500_), .A2(new_n10154_), .B(new_n20611_), .ZN(new_n20612_));
  AOI21_X1   g20315(.A1(new_n20612_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n20613_));
  XOR2_X1    g20316(.A1(new_n5067_), .A2(new_n20613_), .Z(new_n20614_));
  INV_X1     g20317(.I(new_n20614_), .ZN(new_n20615_));
  XOR2_X1    g20318(.A1(new_n20610_), .A2(new_n20615_), .Z(new_n20616_));
  INV_X1     g20319(.I(new_n20610_), .ZN(new_n20617_));
  NOR2_X1    g20320(.A1(new_n20617_), .A2(new_n20614_), .ZN(new_n20618_));
  NOR2_X1    g20321(.A1(new_n20610_), .A2(new_n20615_), .ZN(new_n20619_));
  NOR2_X1    g20322(.A1(new_n20618_), .A2(new_n20619_), .ZN(new_n20620_));
  NOR2_X1    g20323(.A1(new_n20620_), .A2(new_n20608_), .ZN(new_n20621_));
  AOI21_X1   g20324(.A1(new_n20608_), .A2(new_n20616_), .B(new_n20621_), .ZN(new_n20622_));
  XOR2_X1    g20325(.A1(new_n20622_), .A2(new_n20555_), .Z(new_n20623_));
  INV_X1     g20326(.I(new_n20555_), .ZN(new_n20624_));
  NOR2_X1    g20327(.A1(new_n20622_), .A2(new_n20624_), .ZN(new_n20625_));
  NAND2_X1   g20328(.A1(new_n20622_), .A2(new_n20624_), .ZN(new_n20626_));
  INV_X1     g20329(.I(new_n20626_), .ZN(new_n20627_));
  OAI21_X1   g20330(.A1(new_n20627_), .A2(new_n20625_), .B(new_n20554_), .ZN(new_n20628_));
  OAI21_X1   g20331(.A1(new_n20554_), .A2(new_n20623_), .B(new_n20628_), .ZN(new_n20629_));
  OAI22_X1   g20332(.A1(new_n6644_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n6647_), .ZN(new_n20630_));
  OAI21_X1   g20333(.A1(new_n6229_), .A2(new_n7284_), .B(new_n20630_), .ZN(new_n20631_));
  AOI21_X1   g20334(.A1(new_n20631_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n20632_));
  XOR2_X1    g20335(.A1(new_n6851_), .A2(new_n20632_), .Z(new_n20633_));
  NOR2_X1    g20336(.A1(new_n20629_), .A2(new_n20633_), .ZN(new_n20634_));
  INV_X1     g20337(.I(new_n20634_), .ZN(new_n20635_));
  NAND2_X1   g20338(.A1(new_n20629_), .A2(new_n20633_), .ZN(new_n20636_));
  AOI21_X1   g20339(.A1(new_n20635_), .A2(new_n20636_), .B(new_n20550_), .ZN(new_n20637_));
  INV_X1     g20340(.I(new_n20550_), .ZN(new_n20638_));
  XNOR2_X1   g20341(.A1(new_n20629_), .A2(new_n20633_), .ZN(new_n20639_));
  NOR2_X1    g20342(.A1(new_n20639_), .A2(new_n20638_), .ZN(new_n20640_));
  NOR2_X1    g20343(.A1(new_n20640_), .A2(new_n20637_), .ZN(new_n20641_));
  NOR2_X1    g20344(.A1(new_n20424_), .A2(new_n20433_), .ZN(new_n20642_));
  NOR2_X1    g20345(.A1(new_n20642_), .A2(new_n20430_), .ZN(new_n20643_));
  NOR2_X1    g20346(.A1(new_n20641_), .A2(new_n20643_), .ZN(new_n20644_));
  NOR4_X1    g20347(.A1(new_n20640_), .A2(new_n20430_), .A3(new_n20637_), .A4(new_n20642_), .ZN(new_n20645_));
  NOR2_X1    g20348(.A1(new_n20644_), .A2(new_n20645_), .ZN(new_n20646_));
  NOR2_X1    g20349(.A1(new_n20646_), .A2(new_n20549_), .ZN(new_n20647_));
  INV_X1     g20350(.I(new_n20549_), .ZN(new_n20648_));
  XNOR2_X1   g20351(.A1(new_n20641_), .A2(new_n20643_), .ZN(new_n20649_));
  NOR2_X1    g20352(.A1(new_n20649_), .A2(new_n20648_), .ZN(new_n20650_));
  NOR2_X1    g20353(.A1(new_n20650_), .A2(new_n20647_), .ZN(new_n20651_));
  NAND2_X1   g20354(.A1(new_n20445_), .A2(new_n20331_), .ZN(new_n20652_));
  NAND2_X1   g20355(.A1(new_n20652_), .A2(new_n20444_), .ZN(new_n20653_));
  INV_X1     g20356(.I(new_n20653_), .ZN(new_n20654_));
  OAI22_X1   g20357(.A1(new_n5420_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n5107_), .ZN(new_n20655_));
  OAI21_X1   g20358(.A1(new_n8218_), .A2(new_n5112_), .B(new_n20655_), .ZN(new_n20656_));
  AOI21_X1   g20359(.A1(new_n20656_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n20657_));
  XOR2_X1    g20360(.A1(new_n8952_), .A2(new_n20657_), .Z(new_n20658_));
  NOR2_X1    g20361(.A1(new_n20654_), .A2(new_n20658_), .ZN(new_n20659_));
  INV_X1     g20362(.I(new_n20658_), .ZN(new_n20660_));
  NOR2_X1    g20363(.A1(new_n20653_), .A2(new_n20660_), .ZN(new_n20661_));
  NOR2_X1    g20364(.A1(new_n20659_), .A2(new_n20661_), .ZN(new_n20662_));
  NOR2_X1    g20365(.A1(new_n20662_), .A2(new_n20651_), .ZN(new_n20663_));
  INV_X1     g20366(.I(new_n20651_), .ZN(new_n20664_));
  XOR2_X1    g20367(.A1(new_n20653_), .A2(new_n20658_), .Z(new_n20665_));
  NOR2_X1    g20368(.A1(new_n20665_), .A2(new_n20664_), .ZN(new_n20666_));
  NOR2_X1    g20369(.A1(new_n20663_), .A2(new_n20666_), .ZN(new_n20667_));
  NAND2_X1   g20370(.A1(new_n20447_), .A2(new_n20455_), .ZN(new_n20668_));
  AOI21_X1   g20371(.A1(new_n20453_), .A2(new_n20668_), .B(new_n20667_), .ZN(new_n20669_));
  NAND2_X1   g20372(.A1(new_n20668_), .A2(new_n20453_), .ZN(new_n20670_));
  NOR3_X1    g20373(.A1(new_n20670_), .A2(new_n20663_), .A3(new_n20666_), .ZN(new_n20671_));
  OAI21_X1   g20374(.A1(new_n20669_), .A2(new_n20671_), .B(new_n20545_), .ZN(new_n20672_));
  XNOR2_X1   g20375(.A1(new_n20667_), .A2(new_n20670_), .ZN(new_n20673_));
  NAND2_X1   g20376(.A1(new_n20673_), .A2(new_n20544_), .ZN(new_n20674_));
  NAND2_X1   g20377(.A1(new_n20674_), .A2(new_n20672_), .ZN(new_n20675_));
  XOR2_X1    g20378(.A1(new_n20675_), .A2(new_n20540_), .Z(new_n20676_));
  NOR2_X1    g20379(.A1(new_n20676_), .A2(new_n20536_), .ZN(new_n20677_));
  INV_X1     g20380(.I(new_n20536_), .ZN(new_n20678_));
  INV_X1     g20381(.I(new_n20675_), .ZN(new_n20679_));
  NOR2_X1    g20382(.A1(new_n20679_), .A2(new_n20540_), .ZN(new_n20680_));
  INV_X1     g20383(.I(new_n20680_), .ZN(new_n20681_));
  NAND2_X1   g20384(.A1(new_n20679_), .A2(new_n20540_), .ZN(new_n20682_));
  AOI21_X1   g20385(.A1(new_n20681_), .A2(new_n20682_), .B(new_n20678_), .ZN(new_n20683_));
  NOR2_X1    g20386(.A1(new_n20683_), .A2(new_n20677_), .ZN(new_n20684_));
  NOR3_X1    g20387(.A1(new_n20684_), .A2(new_n20474_), .A3(new_n20534_), .ZN(new_n20685_));
  NOR2_X1    g20388(.A1(new_n20534_), .A2(new_n20474_), .ZN(new_n20686_));
  INV_X1     g20389(.I(new_n20684_), .ZN(new_n20687_));
  NOR2_X1    g20390(.A1(new_n20687_), .A2(new_n20686_), .ZN(new_n20688_));
  NOR2_X1    g20391(.A1(new_n20688_), .A2(new_n20685_), .ZN(new_n20689_));
  NOR2_X1    g20392(.A1(new_n20689_), .A2(new_n20533_), .ZN(new_n20690_));
  INV_X1     g20393(.I(new_n20533_), .ZN(new_n20691_));
  XOR2_X1    g20394(.A1(new_n20684_), .A2(new_n20686_), .Z(new_n20692_));
  NOR2_X1    g20395(.A1(new_n20692_), .A2(new_n20691_), .ZN(new_n20693_));
  NOR2_X1    g20396(.A1(new_n20690_), .A2(new_n20693_), .ZN(new_n20694_));
  XNOR2_X1   g20397(.A1(new_n20694_), .A2(new_n20529_), .ZN(new_n20695_));
  NOR2_X1    g20398(.A1(new_n20694_), .A2(new_n20529_), .ZN(new_n20696_));
  NAND2_X1   g20399(.A1(new_n20694_), .A2(new_n20529_), .ZN(new_n20697_));
  INV_X1     g20400(.I(new_n20697_), .ZN(new_n20698_));
  OAI21_X1   g20401(.A1(new_n20698_), .A2(new_n20696_), .B(new_n20527_), .ZN(new_n20699_));
  OAI21_X1   g20402(.A1(new_n20527_), .A2(new_n20695_), .B(new_n20699_), .ZN(new_n20700_));
  AND2_X2    g20403(.A1(new_n20700_), .A2(new_n20523_), .Z(new_n20701_));
  NOR2_X1    g20404(.A1(new_n20700_), .A2(new_n20523_), .ZN(new_n20702_));
  NOR2_X1    g20405(.A1(new_n20701_), .A2(new_n20702_), .ZN(new_n20703_));
  NOR2_X1    g20406(.A1(new_n20703_), .A2(new_n20520_), .ZN(new_n20704_));
  INV_X1     g20407(.I(new_n20520_), .ZN(new_n20705_));
  XOR2_X1    g20408(.A1(new_n20700_), .A2(new_n20522_), .Z(new_n20706_));
  NOR2_X1    g20409(.A1(new_n20706_), .A2(new_n20705_), .ZN(new_n20707_));
  NOR2_X1    g20410(.A1(new_n20704_), .A2(new_n20707_), .ZN(new_n20708_));
  NAND2_X1   g20411(.A1(new_n20496_), .A2(new_n20305_), .ZN(new_n20709_));
  AND2_X2    g20412(.A1(new_n20709_), .A2(new_n20497_), .Z(new_n20710_));
  NOR2_X1    g20413(.A1(new_n20708_), .A2(new_n20710_), .ZN(new_n20711_));
  XOR2_X1    g20414(.A1(new_n20516_), .A2(new_n20711_), .Z(new_n20712_));
  XOR2_X1    g20415(.A1(new_n20712_), .A2(new_n20511_), .Z(\f[85] ));
  NOR2_X1    g20416(.A1(new_n20511_), .A2(new_n20708_), .ZN(new_n20714_));
  INV_X1     g20417(.I(new_n20714_), .ZN(new_n20715_));
  AOI21_X1   g20418(.A1(new_n20511_), .A2(new_n20708_), .B(new_n20710_), .ZN(new_n20716_));
  INV_X1     g20419(.I(new_n20716_), .ZN(new_n20717_));
  OAI21_X1   g20420(.A1(new_n20516_), .A2(new_n20717_), .B(new_n20715_), .ZN(new_n20718_));
  NOR2_X1    g20421(.A1(new_n20701_), .A2(new_n20520_), .ZN(new_n20719_));
  NOR2_X1    g20422(.A1(new_n20719_), .A2(new_n20702_), .ZN(new_n20720_));
  INV_X1     g20423(.I(new_n20685_), .ZN(new_n20721_));
  AOI21_X1   g20424(.A1(new_n20721_), .A2(new_n20691_), .B(new_n20688_), .ZN(new_n20722_));
  OAI22_X1   g20425(.A1(new_n2171_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n2166_), .ZN(new_n20723_));
  OAI21_X1   g20426(.A1(new_n13367_), .A2(new_n2322_), .B(new_n20723_), .ZN(new_n20724_));
  AOI21_X1   g20427(.A1(new_n18183_), .A2(new_n2161_), .B(new_n20724_), .ZN(new_n20725_));
  OAI22_X1   g20428(.A1(new_n12542_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n12970_), .ZN(new_n20726_));
  OAI21_X1   g20429(.A1(new_n12536_), .A2(new_n2884_), .B(new_n20726_), .ZN(new_n20727_));
  AOI21_X1   g20430(.A1(new_n20727_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n20728_));
  XOR2_X1    g20431(.A1(new_n12969_), .A2(new_n20728_), .Z(new_n20729_));
  INV_X1     g20432(.I(new_n20729_), .ZN(new_n20730_));
  OAI22_X1   g20433(.A1(new_n11738_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n11744_), .ZN(new_n20731_));
  OAI21_X1   g20434(.A1(new_n10862_), .A2(new_n3569_), .B(new_n20731_), .ZN(new_n20732_));
  AOI21_X1   g20435(.A1(new_n20732_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n20733_));
  XNOR2_X1   g20436(.A1(new_n11748_), .A2(new_n20733_), .ZN(new_n20734_));
  INV_X1     g20437(.I(new_n20734_), .ZN(new_n20735_));
  NOR2_X1    g20438(.A1(new_n20671_), .A2(new_n20544_), .ZN(new_n20736_));
  NOR2_X1    g20439(.A1(new_n20736_), .A2(new_n20669_), .ZN(new_n20737_));
  OAI22_X1   g20440(.A1(new_n4072_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n4067_), .ZN(new_n20738_));
  OAI21_X1   g20441(.A1(new_n10025_), .A2(new_n4318_), .B(new_n20738_), .ZN(new_n20739_));
  AOI21_X1   g20442(.A1(new_n20739_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n20740_));
  XOR2_X1    g20443(.A1(new_n10476_), .A2(new_n20740_), .Z(new_n20741_));
  INV_X1     g20444(.I(new_n20741_), .ZN(new_n20742_));
  OAI22_X1   g20445(.A1(new_n5420_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n5107_), .ZN(new_n20743_));
  OAI21_X1   g20446(.A1(new_n8563_), .A2(new_n5112_), .B(new_n20743_), .ZN(new_n20744_));
  AOI21_X1   g20447(.A1(new_n20744_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n20745_));
  XNOR2_X1   g20448(.A1(new_n9299_), .A2(new_n20745_), .ZN(new_n20746_));
  OAI22_X1   g20449(.A1(new_n6644_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n6647_), .ZN(new_n20747_));
  OAI21_X1   g20450(.A1(new_n6538_), .A2(new_n7284_), .B(new_n20747_), .ZN(new_n20748_));
  AOI21_X1   g20451(.A1(new_n20748_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n20749_));
  XNOR2_X1   g20452(.A1(new_n7202_), .A2(new_n20749_), .ZN(new_n20750_));
  INV_X1     g20453(.I(new_n20750_), .ZN(new_n20751_));
  OAI21_X1   g20454(.A1(new_n20554_), .A2(new_n20625_), .B(new_n20626_), .ZN(new_n20752_));
  INV_X1     g20455(.I(new_n20752_), .ZN(new_n20753_));
  AOI22_X1   g20456(.A1(new_n8631_), .A2(\b[37] ), .B1(\b[38] ), .B2(new_n9382_), .ZN(new_n20754_));
  AOI21_X1   g20457(.A1(\b[36] ), .A2(new_n9731_), .B(new_n20754_), .ZN(new_n20755_));
  OAI21_X1   g20458(.A1(new_n20755_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n20756_));
  XOR2_X1    g20459(.A1(new_n5357_), .A2(new_n20756_), .Z(new_n20757_));
  AOI21_X1   g20460(.A1(new_n20560_), .A2(new_n20604_), .B(new_n20603_), .ZN(new_n20758_));
  INV_X1     g20461(.I(new_n20758_), .ZN(new_n20759_));
  AOI22_X1   g20462(.A1(new_n11415_), .A2(new_n4770_), .B1(\b[33] ), .B2(new_n10145_), .ZN(new_n20760_));
  OAI21_X1   g20463(.A1(new_n20760_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n20761_));
  XNOR2_X1   g20464(.A1(new_n4499_), .A2(new_n20761_), .ZN(new_n20762_));
  AOI22_X1   g20465(.A1(new_n10969_), .A2(new_n3719_), .B1(new_n11394_), .B2(\b[30] ), .ZN(new_n20763_));
  OAI21_X1   g20466(.A1(new_n20763_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n20764_));
  XNOR2_X1   g20467(.A1(new_n3722_), .A2(new_n20764_), .ZN(new_n20765_));
  OAI22_X1   g20468(.A1(new_n13880_), .A2(new_n2440_), .B1(new_n2102_), .B2(new_n13885_), .ZN(new_n20766_));
  AOI21_X1   g20469(.A1(new_n20766_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n20767_));
  XOR2_X1    g20470(.A1(new_n2443_), .A2(new_n20767_), .Z(new_n20768_));
  NOR2_X1    g20471(.A1(new_n13476_), .A2(new_n1803_), .ZN(new_n20769_));
  XOR2_X1    g20472(.A1(new_n14736_), .A2(new_n1803_), .Z(new_n20770_));
  NAND2_X1   g20473(.A1(new_n20770_), .A2(\b[23] ), .ZN(new_n20771_));
  XOR2_X1    g20474(.A1(new_n20771_), .A2(new_n20769_), .Z(new_n20772_));
  XOR2_X1    g20475(.A1(new_n20574_), .A2(new_n20772_), .Z(new_n20773_));
  INV_X1     g20476(.I(new_n20773_), .ZN(new_n20774_));
  NOR2_X1    g20477(.A1(new_n20575_), .A2(new_n20772_), .ZN(new_n20775_));
  INV_X1     g20478(.I(new_n20772_), .ZN(new_n20776_));
  NOR2_X1    g20479(.A1(new_n20776_), .A2(new_n20574_), .ZN(new_n20777_));
  NOR2_X1    g20480(.A1(new_n20775_), .A2(new_n20777_), .ZN(new_n20778_));
  NOR2_X1    g20481(.A1(new_n20768_), .A2(new_n20778_), .ZN(new_n20779_));
  AOI21_X1   g20482(.A1(new_n20768_), .A2(new_n20774_), .B(new_n20779_), .ZN(new_n20780_));
  AOI22_X1   g20483(.A1(new_n13078_), .A2(\b[27] ), .B1(new_n3256_), .B2(new_n12218_), .ZN(new_n20781_));
  OAI21_X1   g20484(.A1(new_n20781_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n20782_));
  XOR2_X1    g20485(.A1(new_n3022_), .A2(new_n20782_), .Z(new_n20783_));
  OAI21_X1   g20486(.A1(new_n20568_), .A2(new_n20578_), .B(new_n20579_), .ZN(new_n20784_));
  XOR2_X1    g20487(.A1(new_n20783_), .A2(new_n20784_), .Z(new_n20785_));
  NOR2_X1    g20488(.A1(new_n20785_), .A2(new_n20780_), .ZN(new_n20786_));
  INV_X1     g20489(.I(new_n20784_), .ZN(new_n20787_));
  NOR2_X1    g20490(.A1(new_n20783_), .A2(new_n20787_), .ZN(new_n20788_));
  INV_X1     g20491(.I(new_n20788_), .ZN(new_n20789_));
  NAND2_X1   g20492(.A1(new_n20783_), .A2(new_n20787_), .ZN(new_n20790_));
  NAND2_X1   g20493(.A1(new_n20789_), .A2(new_n20790_), .ZN(new_n20791_));
  AOI21_X1   g20494(.A1(new_n20780_), .A2(new_n20791_), .B(new_n20786_), .ZN(new_n20792_));
  INV_X1     g20495(.I(new_n20564_), .ZN(new_n20793_));
  AOI21_X1   g20496(.A1(new_n20793_), .A2(new_n20585_), .B(new_n20586_), .ZN(new_n20794_));
  XNOR2_X1   g20497(.A1(new_n20792_), .A2(new_n20794_), .ZN(new_n20795_));
  NOR2_X1    g20498(.A1(new_n20795_), .A2(new_n20765_), .ZN(new_n20796_));
  INV_X1     g20499(.I(new_n20765_), .ZN(new_n20797_));
  NOR2_X1    g20500(.A1(new_n20792_), .A2(new_n20794_), .ZN(new_n20798_));
  INV_X1     g20501(.I(new_n20798_), .ZN(new_n20799_));
  NAND2_X1   g20502(.A1(new_n20792_), .A2(new_n20794_), .ZN(new_n20800_));
  AOI21_X1   g20503(.A1(new_n20799_), .A2(new_n20800_), .B(new_n20797_), .ZN(new_n20801_));
  NOR2_X1    g20504(.A1(new_n20796_), .A2(new_n20801_), .ZN(new_n20802_));
  AOI21_X1   g20505(.A1(new_n20598_), .A2(new_n20596_), .B(new_n20594_), .ZN(new_n20803_));
  XOR2_X1    g20506(.A1(new_n20802_), .A2(new_n20803_), .Z(new_n20804_));
  NOR2_X1    g20507(.A1(new_n20804_), .A2(new_n20762_), .ZN(new_n20805_));
  INV_X1     g20508(.I(new_n20762_), .ZN(new_n20806_));
  INV_X1     g20509(.I(new_n20802_), .ZN(new_n20807_));
  NOR2_X1    g20510(.A1(new_n20807_), .A2(new_n20803_), .ZN(new_n20808_));
  INV_X1     g20511(.I(new_n20808_), .ZN(new_n20809_));
  NAND2_X1   g20512(.A1(new_n20807_), .A2(new_n20803_), .ZN(new_n20810_));
  AOI21_X1   g20513(.A1(new_n20809_), .A2(new_n20810_), .B(new_n20806_), .ZN(new_n20811_));
  NOR2_X1    g20514(.A1(new_n20811_), .A2(new_n20805_), .ZN(new_n20812_));
  NOR2_X1    g20515(.A1(new_n20812_), .A2(new_n20759_), .ZN(new_n20813_));
  INV_X1     g20516(.I(new_n20813_), .ZN(new_n20814_));
  NAND2_X1   g20517(.A1(new_n20812_), .A2(new_n20759_), .ZN(new_n20815_));
  AOI21_X1   g20518(.A1(new_n20814_), .A2(new_n20815_), .B(new_n20757_), .ZN(new_n20816_));
  INV_X1     g20519(.I(new_n20757_), .ZN(new_n20817_));
  XOR2_X1    g20520(.A1(new_n20812_), .A2(new_n20758_), .Z(new_n20818_));
  NOR2_X1    g20521(.A1(new_n20818_), .A2(new_n20817_), .ZN(new_n20819_));
  NOR2_X1    g20522(.A1(new_n20819_), .A2(new_n20816_), .ZN(new_n20820_));
  OAI22_X1   g20523(.A1(new_n7619_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n8309_), .ZN(new_n20821_));
  OAI21_X1   g20524(.A1(new_n5913_), .A2(new_n7947_), .B(new_n20821_), .ZN(new_n20822_));
  AOI21_X1   g20525(.A1(new_n20822_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n20823_));
  XOR2_X1    g20526(.A1(new_n6233_), .A2(new_n20823_), .Z(new_n20824_));
  INV_X1     g20527(.I(new_n20619_), .ZN(new_n20825_));
  AOI21_X1   g20528(.A1(new_n20608_), .A2(new_n20825_), .B(new_n20618_), .ZN(new_n20826_));
  NOR2_X1    g20529(.A1(new_n20826_), .A2(new_n20824_), .ZN(new_n20827_));
  INV_X1     g20530(.I(new_n20827_), .ZN(new_n20828_));
  NAND2_X1   g20531(.A1(new_n20826_), .A2(new_n20824_), .ZN(new_n20829_));
  AOI21_X1   g20532(.A1(new_n20828_), .A2(new_n20829_), .B(new_n20820_), .ZN(new_n20830_));
  INV_X1     g20533(.I(new_n20820_), .ZN(new_n20831_));
  XNOR2_X1   g20534(.A1(new_n20826_), .A2(new_n20824_), .ZN(new_n20832_));
  NOR2_X1    g20535(.A1(new_n20831_), .A2(new_n20832_), .ZN(new_n20833_));
  NOR2_X1    g20536(.A1(new_n20833_), .A2(new_n20830_), .ZN(new_n20834_));
  XOR2_X1    g20537(.A1(new_n20834_), .A2(new_n20753_), .Z(new_n20835_));
  NAND2_X1   g20538(.A1(new_n20835_), .A2(new_n20751_), .ZN(new_n20836_));
  NOR2_X1    g20539(.A1(new_n20834_), .A2(new_n20753_), .ZN(new_n20837_));
  NAND2_X1   g20540(.A1(new_n20834_), .A2(new_n20753_), .ZN(new_n20838_));
  INV_X1     g20541(.I(new_n20838_), .ZN(new_n20839_));
  OAI21_X1   g20542(.A1(new_n20839_), .A2(new_n20837_), .B(new_n20750_), .ZN(new_n20840_));
  NAND2_X1   g20543(.A1(new_n20836_), .A2(new_n20840_), .ZN(new_n20841_));
  INV_X1     g20544(.I(new_n20841_), .ZN(new_n20842_));
  OAI22_X1   g20545(.A1(new_n5993_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n5991_), .ZN(new_n20843_));
  OAI21_X1   g20546(.A1(new_n7864_), .A2(new_n5997_), .B(new_n20843_), .ZN(new_n20844_));
  AOI21_X1   g20547(.A1(new_n20844_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n20845_));
  XOR2_X1    g20548(.A1(new_n8217_), .A2(new_n20845_), .Z(new_n20846_));
  AOI21_X1   g20549(.A1(new_n20638_), .A2(new_n20636_), .B(new_n20634_), .ZN(new_n20847_));
  XNOR2_X1   g20550(.A1(new_n20847_), .A2(new_n20846_), .ZN(new_n20848_));
  NOR2_X1    g20551(.A1(new_n20848_), .A2(new_n20842_), .ZN(new_n20849_));
  NOR2_X1    g20552(.A1(new_n20847_), .A2(new_n20846_), .ZN(new_n20850_));
  INV_X1     g20553(.I(new_n20850_), .ZN(new_n20851_));
  NAND2_X1   g20554(.A1(new_n20847_), .A2(new_n20846_), .ZN(new_n20852_));
  AOI21_X1   g20555(.A1(new_n20851_), .A2(new_n20852_), .B(new_n20841_), .ZN(new_n20853_));
  NOR2_X1    g20556(.A1(new_n20849_), .A2(new_n20853_), .ZN(new_n20854_));
  NOR2_X1    g20557(.A1(new_n20645_), .A2(new_n20549_), .ZN(new_n20855_));
  NOR2_X1    g20558(.A1(new_n20855_), .A2(new_n20644_), .ZN(new_n20856_));
  XNOR2_X1   g20559(.A1(new_n20854_), .A2(new_n20856_), .ZN(new_n20857_));
  NOR2_X1    g20560(.A1(new_n20857_), .A2(new_n20746_), .ZN(new_n20858_));
  INV_X1     g20561(.I(new_n20746_), .ZN(new_n20859_));
  NOR2_X1    g20562(.A1(new_n20854_), .A2(new_n20856_), .ZN(new_n20860_));
  INV_X1     g20563(.I(new_n20860_), .ZN(new_n20861_));
  NAND2_X1   g20564(.A1(new_n20854_), .A2(new_n20856_), .ZN(new_n20862_));
  AOI21_X1   g20565(.A1(new_n20861_), .A2(new_n20862_), .B(new_n20859_), .ZN(new_n20863_));
  INV_X1     g20566(.I(new_n20661_), .ZN(new_n20864_));
  AOI21_X1   g20567(.A1(new_n20664_), .A2(new_n20864_), .B(new_n20659_), .ZN(new_n20865_));
  NOR3_X1    g20568(.A1(new_n20865_), .A2(new_n20858_), .A3(new_n20863_), .ZN(new_n20866_));
  NOR2_X1    g20569(.A1(new_n20858_), .A2(new_n20863_), .ZN(new_n20867_));
  INV_X1     g20570(.I(new_n20865_), .ZN(new_n20868_));
  NOR2_X1    g20571(.A1(new_n20868_), .A2(new_n20867_), .ZN(new_n20869_));
  OAI21_X1   g20572(.A1(new_n20869_), .A2(new_n20866_), .B(new_n20742_), .ZN(new_n20870_));
  XOR2_X1    g20573(.A1(new_n20867_), .A2(new_n20865_), .Z(new_n20871_));
  OAI21_X1   g20574(.A1(new_n20742_), .A2(new_n20871_), .B(new_n20870_), .ZN(new_n20872_));
  INV_X1     g20575(.I(new_n20872_), .ZN(new_n20873_));
  NOR2_X1    g20576(.A1(new_n20873_), .A2(new_n20737_), .ZN(new_n20874_));
  NOR3_X1    g20577(.A1(new_n20872_), .A2(new_n20669_), .A3(new_n20736_), .ZN(new_n20875_));
  OAI21_X1   g20578(.A1(new_n20874_), .A2(new_n20875_), .B(new_n20735_), .ZN(new_n20876_));
  XOR2_X1    g20579(.A1(new_n20872_), .A2(new_n20737_), .Z(new_n20877_));
  OAI21_X1   g20580(.A1(new_n20735_), .A2(new_n20877_), .B(new_n20876_), .ZN(new_n20878_));
  INV_X1     g20581(.I(new_n20878_), .ZN(new_n20879_));
  AOI21_X1   g20582(.A1(new_n20678_), .A2(new_n20682_), .B(new_n20680_), .ZN(new_n20880_));
  NOR2_X1    g20583(.A1(new_n20879_), .A2(new_n20880_), .ZN(new_n20881_));
  INV_X1     g20584(.I(new_n20880_), .ZN(new_n20882_));
  NOR2_X1    g20585(.A1(new_n20882_), .A2(new_n20878_), .ZN(new_n20883_));
  OAI21_X1   g20586(.A1(new_n20883_), .A2(new_n20881_), .B(new_n20730_), .ZN(new_n20884_));
  XOR2_X1    g20587(.A1(new_n20880_), .A2(new_n20878_), .Z(new_n20885_));
  OAI21_X1   g20588(.A1(new_n20730_), .A2(new_n20885_), .B(new_n20884_), .ZN(new_n20886_));
  XOR2_X1    g20589(.A1(new_n20886_), .A2(new_n20725_), .Z(new_n20887_));
  XOR2_X1    g20590(.A1(new_n20887_), .A2(new_n20722_), .Z(new_n20888_));
  XOR2_X1    g20591(.A1(new_n20888_), .A2(\a[26] ), .Z(new_n20889_));
  OAI21_X1   g20592(.A1(new_n1712_), .A2(new_n1850_), .B(new_n16487_), .ZN(new_n20890_));
  NOR2_X1    g20593(.A1(new_n20698_), .A2(new_n20527_), .ZN(new_n20891_));
  NOR2_X1    g20594(.A1(new_n20891_), .A2(new_n20696_), .ZN(new_n20892_));
  XNOR2_X1   g20595(.A1(new_n20892_), .A2(new_n20890_), .ZN(new_n20893_));
  XOR2_X1    g20596(.A1(new_n20893_), .A2(new_n20889_), .Z(new_n20894_));
  XOR2_X1    g20597(.A1(new_n20894_), .A2(\a[23] ), .Z(new_n20895_));
  NOR2_X1    g20598(.A1(new_n20895_), .A2(new_n20720_), .ZN(new_n20896_));
  NAND2_X1   g20599(.A1(new_n20895_), .A2(new_n20720_), .ZN(new_n20897_));
  INV_X1     g20600(.I(new_n20897_), .ZN(new_n20898_));
  NOR2_X1    g20601(.A1(new_n20898_), .A2(new_n20896_), .ZN(new_n20899_));
  XNOR2_X1   g20602(.A1(new_n20718_), .A2(new_n20899_), .ZN(\f[86] ));
  NOR2_X1    g20603(.A1(new_n20889_), .A2(new_n20892_), .ZN(new_n20901_));
  XOR2_X1    g20604(.A1(new_n20890_), .A2(new_n1709_), .Z(new_n20902_));
  AOI21_X1   g20605(.A1(new_n20889_), .A2(new_n20892_), .B(new_n20902_), .ZN(new_n20903_));
  NOR2_X1    g20606(.A1(new_n20903_), .A2(new_n20901_), .ZN(new_n20904_));
  INV_X1     g20607(.I(new_n20722_), .ZN(new_n20905_));
  NAND2_X1   g20608(.A1(new_n20905_), .A2(new_n20886_), .ZN(new_n20906_));
  XOR2_X1    g20609(.A1(new_n20725_), .A2(\a[26] ), .Z(new_n20907_));
  OAI21_X1   g20610(.A1(new_n20905_), .A2(new_n20886_), .B(new_n20907_), .ZN(new_n20908_));
  NAND2_X1   g20611(.A1(new_n20908_), .A2(new_n20906_), .ZN(new_n20909_));
  OAI22_X1   g20612(.A1(new_n2171_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n2166_), .ZN(new_n20910_));
  OAI21_X1   g20613(.A1(new_n13785_), .A2(new_n2322_), .B(new_n20910_), .ZN(new_n20911_));
  AOI21_X1   g20614(.A1(new_n20911_), .A2(new_n2168_), .B(new_n2171_), .ZN(new_n20912_));
  XNOR2_X1   g20615(.A1(new_n14599_), .A2(new_n20912_), .ZN(new_n20913_));
  NOR2_X1    g20616(.A1(new_n20883_), .A2(new_n20729_), .ZN(new_n20914_));
  AOI22_X1   g20617(.A1(new_n2694_), .A2(\b[59] ), .B1(\b[60] ), .B2(new_n2699_), .ZN(new_n20915_));
  AOI21_X1   g20618(.A1(\b[58] ), .A2(new_n4094_), .B(new_n20915_), .ZN(new_n20916_));
  OAI21_X1   g20619(.A1(new_n20916_), .A2(\a[29] ), .B(new_n2694_), .ZN(new_n20917_));
  XNOR2_X1   g20620(.A1(new_n13371_), .A2(new_n20917_), .ZN(new_n20918_));
  NOR2_X1    g20621(.A1(new_n20875_), .A2(new_n20734_), .ZN(new_n20919_));
  NOR2_X1    g20622(.A1(new_n20919_), .A2(new_n20874_), .ZN(new_n20920_));
  INV_X1     g20623(.I(new_n20920_), .ZN(new_n20921_));
  OAI22_X1   g20624(.A1(new_n11744_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n12536_), .ZN(new_n20922_));
  OAI21_X1   g20625(.A1(new_n11738_), .A2(new_n3569_), .B(new_n20922_), .ZN(new_n20923_));
  AOI21_X1   g20626(.A1(new_n20923_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n20924_));
  XNOR2_X1   g20627(.A1(new_n12128_), .A2(new_n20924_), .ZN(new_n20925_));
  INV_X1     g20628(.I(new_n20925_), .ZN(new_n20926_));
  NOR2_X1    g20629(.A1(new_n20869_), .A2(new_n20741_), .ZN(new_n20927_));
  NOR2_X1    g20630(.A1(new_n20927_), .A2(new_n20866_), .ZN(new_n20928_));
  AOI21_X1   g20631(.A1(new_n20859_), .A2(new_n20862_), .B(new_n20860_), .ZN(new_n20929_));
  INV_X1     g20632(.I(new_n20929_), .ZN(new_n20930_));
  AOI21_X1   g20633(.A1(new_n20751_), .A2(new_n20838_), .B(new_n20837_), .ZN(new_n20931_));
  AOI21_X1   g20634(.A1(new_n20831_), .A2(new_n20829_), .B(new_n20827_), .ZN(new_n20932_));
  OAI21_X1   g20635(.A1(new_n20757_), .A2(new_n20813_), .B(new_n20815_), .ZN(new_n20933_));
  INV_X1     g20636(.I(new_n20933_), .ZN(new_n20934_));
  AOI21_X1   g20637(.A1(new_n20797_), .A2(new_n20800_), .B(new_n20798_), .ZN(new_n20935_));
  AOI21_X1   g20638(.A1(new_n20780_), .A2(new_n20790_), .B(new_n20788_), .ZN(new_n20936_));
  INV_X1     g20639(.I(new_n20775_), .ZN(new_n20937_));
  AOI21_X1   g20640(.A1(new_n20768_), .A2(new_n20937_), .B(new_n20777_), .ZN(new_n20938_));
  INV_X1     g20641(.I(new_n20938_), .ZN(new_n20939_));
  OAI22_X1   g20642(.A1(new_n13880_), .A2(new_n2837_), .B1(new_n2281_), .B2(new_n13885_), .ZN(new_n20940_));
  AOI21_X1   g20643(.A1(new_n20940_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n20941_));
  XNOR2_X1   g20644(.A1(new_n2647_), .A2(new_n20941_), .ZN(new_n20942_));
  INV_X1     g20645(.I(new_n20942_), .ZN(new_n20943_));
  NOR2_X1    g20646(.A1(new_n13476_), .A2(new_n1936_), .ZN(new_n20944_));
  XOR2_X1    g20647(.A1(new_n14736_), .A2(new_n1936_), .Z(new_n20945_));
  NAND2_X1   g20648(.A1(new_n20945_), .A2(\b[24] ), .ZN(new_n20946_));
  XOR2_X1    g20649(.A1(new_n20946_), .A2(new_n20944_), .Z(new_n20947_));
  XOR2_X1    g20650(.A1(new_n20947_), .A2(\a[23] ), .Z(new_n20948_));
  NOR2_X1    g20651(.A1(new_n20948_), .A2(new_n20772_), .ZN(new_n20949_));
  NOR2_X1    g20652(.A1(new_n20947_), .A2(new_n1709_), .ZN(new_n20950_));
  INV_X1     g20653(.I(new_n20950_), .ZN(new_n20951_));
  NAND2_X1   g20654(.A1(new_n20947_), .A2(new_n1709_), .ZN(new_n20952_));
  AOI21_X1   g20655(.A1(new_n20951_), .A2(new_n20952_), .B(new_n20776_), .ZN(new_n20953_));
  NOR2_X1    g20656(.A1(new_n20949_), .A2(new_n20953_), .ZN(new_n20954_));
  NOR2_X1    g20657(.A1(new_n20943_), .A2(new_n20954_), .ZN(new_n20955_));
  NAND2_X1   g20658(.A1(new_n20943_), .A2(new_n20954_), .ZN(new_n20956_));
  INV_X1     g20659(.I(new_n20956_), .ZN(new_n20957_));
  OAI21_X1   g20660(.A1(new_n20957_), .A2(new_n20955_), .B(new_n20939_), .ZN(new_n20958_));
  XNOR2_X1   g20661(.A1(new_n20942_), .A2(new_n20954_), .ZN(new_n20959_));
  NAND2_X1   g20662(.A1(new_n20959_), .A2(new_n20938_), .ZN(new_n20960_));
  NAND2_X1   g20663(.A1(new_n20958_), .A2(new_n20960_), .ZN(new_n20961_));
  AOI22_X1   g20664(.A1(new_n13078_), .A2(\b[28] ), .B1(new_n19751_), .B2(new_n12218_), .ZN(new_n20962_));
  OAI21_X1   g20665(.A1(new_n20962_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n20963_));
  XOR2_X1    g20666(.A1(new_n3264_), .A2(new_n20963_), .Z(new_n20964_));
  XOR2_X1    g20667(.A1(new_n20961_), .A2(new_n20964_), .Z(new_n20965_));
  AOI21_X1   g20668(.A1(new_n20958_), .A2(new_n20960_), .B(new_n20964_), .ZN(new_n20966_));
  INV_X1     g20669(.I(new_n20964_), .ZN(new_n20967_));
  NOR2_X1    g20670(.A1(new_n20967_), .A2(new_n20961_), .ZN(new_n20968_));
  OAI21_X1   g20671(.A1(new_n20968_), .A2(new_n20966_), .B(new_n20936_), .ZN(new_n20969_));
  OAI21_X1   g20672(.A1(new_n20936_), .A2(new_n20965_), .B(new_n20969_), .ZN(new_n20970_));
  AOI22_X1   g20673(.A1(new_n10969_), .A2(new_n4249_), .B1(new_n11394_), .B2(\b[31] ), .ZN(new_n20971_));
  OAI21_X1   g20674(.A1(new_n20971_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n20972_));
  XOR2_X1    g20675(.A1(new_n3993_), .A2(new_n20972_), .Z(new_n20973_));
  XNOR2_X1   g20676(.A1(new_n20970_), .A2(new_n20973_), .ZN(new_n20974_));
  NOR2_X1    g20677(.A1(new_n20974_), .A2(new_n20935_), .ZN(new_n20975_));
  INV_X1     g20678(.I(new_n20935_), .ZN(new_n20976_));
  OR2_X2     g20679(.A1(new_n20970_), .A2(new_n20973_), .Z(new_n20977_));
  NAND2_X1   g20680(.A1(new_n20970_), .A2(new_n20973_), .ZN(new_n20978_));
  AOI21_X1   g20681(.A1(new_n20977_), .A2(new_n20978_), .B(new_n20976_), .ZN(new_n20979_));
  NOR2_X1    g20682(.A1(new_n20975_), .A2(new_n20979_), .ZN(new_n20980_));
  INV_X1     g20683(.I(new_n4775_), .ZN(new_n20981_));
  AOI22_X1   g20684(.A1(new_n11415_), .A2(new_n20981_), .B1(\b[34] ), .B2(new_n10145_), .ZN(new_n20982_));
  OAI21_X1   g20685(.A1(new_n20982_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n20983_));
  XOR2_X1    g20686(.A1(new_n4778_), .A2(new_n20983_), .Z(new_n20984_));
  NAND2_X1   g20687(.A1(new_n20810_), .A2(new_n20806_), .ZN(new_n20985_));
  AOI21_X1   g20688(.A1(new_n20985_), .A2(new_n20809_), .B(new_n20984_), .ZN(new_n20986_));
  INV_X1     g20689(.I(new_n20986_), .ZN(new_n20987_));
  INV_X1     g20690(.I(new_n20984_), .ZN(new_n20988_));
  NAND2_X1   g20691(.A1(new_n20985_), .A2(new_n20809_), .ZN(new_n20989_));
  NOR2_X1    g20692(.A1(new_n20989_), .A2(new_n20988_), .ZN(new_n20990_));
  INV_X1     g20693(.I(new_n20990_), .ZN(new_n20991_));
  AOI21_X1   g20694(.A1(new_n20991_), .A2(new_n20987_), .B(new_n20980_), .ZN(new_n20992_));
  XOR2_X1    g20695(.A1(new_n20989_), .A2(new_n20984_), .Z(new_n20993_));
  NOR3_X1    g20696(.A1(new_n20993_), .A2(new_n20975_), .A3(new_n20979_), .ZN(new_n20994_));
  NOR2_X1    g20697(.A1(new_n20994_), .A2(new_n20992_), .ZN(new_n20995_));
  OAI22_X1   g20698(.A1(new_n8644_), .A2(new_n5353_), .B1(new_n5913_), .B2(new_n9388_), .ZN(new_n20996_));
  OAI21_X1   g20699(.A1(new_n5068_), .A2(new_n10154_), .B(new_n20996_), .ZN(new_n20997_));
  AOI21_X1   g20700(.A1(new_n20997_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n20998_));
  XNOR2_X1   g20701(.A1(new_n5600_), .A2(new_n20998_), .ZN(new_n20999_));
  XOR2_X1    g20702(.A1(new_n20995_), .A2(new_n20999_), .Z(new_n21000_));
  NOR2_X1    g20703(.A1(new_n21000_), .A2(new_n20934_), .ZN(new_n21001_));
  INV_X1     g20704(.I(new_n20995_), .ZN(new_n21002_));
  NOR2_X1    g20705(.A1(new_n21002_), .A2(new_n20999_), .ZN(new_n21003_));
  INV_X1     g20706(.I(new_n21003_), .ZN(new_n21004_));
  NAND2_X1   g20707(.A1(new_n21002_), .A2(new_n20999_), .ZN(new_n21005_));
  AOI21_X1   g20708(.A1(new_n21004_), .A2(new_n21005_), .B(new_n20933_), .ZN(new_n21006_));
  NOR2_X1    g20709(.A1(new_n21006_), .A2(new_n21001_), .ZN(new_n21007_));
  INV_X1     g20710(.I(new_n21007_), .ZN(new_n21008_));
  OAI22_X1   g20711(.A1(new_n7619_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n8309_), .ZN(new_n21009_));
  OAI21_X1   g20712(.A1(new_n5921_), .A2(new_n7947_), .B(new_n21009_), .ZN(new_n21010_));
  AOI21_X1   g20713(.A1(new_n21010_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n21011_));
  XOR2_X1    g20714(.A1(new_n6543_), .A2(new_n21011_), .Z(new_n21012_));
  NOR2_X1    g20715(.A1(new_n21008_), .A2(new_n21012_), .ZN(new_n21013_));
  INV_X1     g20716(.I(new_n21013_), .ZN(new_n21014_));
  NAND2_X1   g20717(.A1(new_n21008_), .A2(new_n21012_), .ZN(new_n21015_));
  AOI21_X1   g20718(.A1(new_n21014_), .A2(new_n21015_), .B(new_n20932_), .ZN(new_n21016_));
  XNOR2_X1   g20719(.A1(new_n21007_), .A2(new_n21012_), .ZN(new_n21017_));
  AOI21_X1   g20720(.A1(new_n20932_), .A2(new_n21017_), .B(new_n21016_), .ZN(new_n21018_));
  OAI22_X1   g20721(.A1(new_n6644_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n6647_), .ZN(new_n21019_));
  OAI21_X1   g20722(.A1(new_n6847_), .A2(new_n7284_), .B(new_n21019_), .ZN(new_n21020_));
  AOI21_X1   g20723(.A1(new_n21020_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n21021_));
  XOR2_X1    g20724(.A1(new_n7516_), .A2(new_n21021_), .Z(new_n21022_));
  XNOR2_X1   g20725(.A1(new_n21018_), .A2(new_n21022_), .ZN(new_n21023_));
  NOR2_X1    g20726(.A1(new_n21023_), .A2(new_n20931_), .ZN(new_n21024_));
  INV_X1     g20727(.I(new_n20931_), .ZN(new_n21025_));
  NOR2_X1    g20728(.A1(new_n21018_), .A2(new_n21022_), .ZN(new_n21026_));
  INV_X1     g20729(.I(new_n21026_), .ZN(new_n21027_));
  NAND2_X1   g20730(.A1(new_n21018_), .A2(new_n21022_), .ZN(new_n21028_));
  AOI21_X1   g20731(.A1(new_n21027_), .A2(new_n21028_), .B(new_n21025_), .ZN(new_n21029_));
  NOR2_X1    g20732(.A1(new_n21024_), .A2(new_n21029_), .ZN(new_n21030_));
  AOI22_X1   g20733(.A1(new_n5680_), .A2(\b[47] ), .B1(\b[48] ), .B2(new_n5686_), .ZN(new_n21031_));
  AOI21_X1   g20734(.A1(\b[46] ), .A2(new_n6923_), .B(new_n21031_), .ZN(new_n21032_));
  OAI21_X1   g20735(.A1(new_n21032_), .A2(\a[41] ), .B(new_n5680_), .ZN(new_n21033_));
  XOR2_X1    g20736(.A1(new_n8568_), .A2(new_n21033_), .Z(new_n21034_));
  NAND2_X1   g20737(.A1(new_n20842_), .A2(new_n20852_), .ZN(new_n21035_));
  NAND2_X1   g20738(.A1(new_n21035_), .A2(new_n20851_), .ZN(new_n21036_));
  NAND2_X1   g20739(.A1(new_n21036_), .A2(new_n21034_), .ZN(new_n21037_));
  NOR2_X1    g20740(.A1(new_n21036_), .A2(new_n21034_), .ZN(new_n21038_));
  INV_X1     g20741(.I(new_n21038_), .ZN(new_n21039_));
  AOI21_X1   g20742(.A1(new_n21037_), .A2(new_n21039_), .B(new_n21030_), .ZN(new_n21040_));
  XNOR2_X1   g20743(.A1(new_n21036_), .A2(new_n21034_), .ZN(new_n21041_));
  NOR3_X1    g20744(.A1(new_n21024_), .A2(new_n21041_), .A3(new_n21029_), .ZN(new_n21042_));
  OAI22_X1   g20745(.A1(new_n5420_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n5107_), .ZN(new_n21043_));
  OAI21_X1   g20746(.A1(new_n8948_), .A2(new_n5112_), .B(new_n21043_), .ZN(new_n21044_));
  AOI21_X1   g20747(.A1(new_n21044_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n21045_));
  XNOR2_X1   g20748(.A1(new_n9642_), .A2(new_n21045_), .ZN(new_n21046_));
  NOR3_X1    g20749(.A1(new_n21040_), .A2(new_n21042_), .A3(new_n21046_), .ZN(new_n21047_));
  NOR2_X1    g20750(.A1(new_n21040_), .A2(new_n21042_), .ZN(new_n21048_));
  INV_X1     g20751(.I(new_n21046_), .ZN(new_n21049_));
  NOR2_X1    g20752(.A1(new_n21048_), .A2(new_n21049_), .ZN(new_n21050_));
  OAI21_X1   g20753(.A1(new_n21050_), .A2(new_n21047_), .B(new_n20930_), .ZN(new_n21051_));
  XOR2_X1    g20754(.A1(new_n21048_), .A2(new_n21049_), .Z(new_n21052_));
  NAND2_X1   g20755(.A1(new_n21052_), .A2(new_n20929_), .ZN(new_n21053_));
  NAND2_X1   g20756(.A1(new_n21053_), .A2(new_n21051_), .ZN(new_n21054_));
  OAI22_X1   g20757(.A1(new_n4072_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n4067_), .ZN(new_n21055_));
  OAI21_X1   g20758(.A1(new_n10031_), .A2(new_n4318_), .B(new_n21055_), .ZN(new_n21056_));
  AOI21_X1   g20759(.A1(new_n21056_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n21057_));
  XNOR2_X1   g20760(.A1(new_n10866_), .A2(new_n21057_), .ZN(new_n21058_));
  XOR2_X1    g20761(.A1(new_n21054_), .A2(new_n21058_), .Z(new_n21059_));
  NOR2_X1    g20762(.A1(new_n21059_), .A2(new_n20928_), .ZN(new_n21060_));
  INV_X1     g20763(.I(new_n20928_), .ZN(new_n21061_));
  INV_X1     g20764(.I(new_n21054_), .ZN(new_n21062_));
  NOR2_X1    g20765(.A1(new_n21062_), .A2(new_n21058_), .ZN(new_n21063_));
  INV_X1     g20766(.I(new_n21063_), .ZN(new_n21064_));
  NAND2_X1   g20767(.A1(new_n21062_), .A2(new_n21058_), .ZN(new_n21065_));
  AOI21_X1   g20768(.A1(new_n21064_), .A2(new_n21065_), .B(new_n21061_), .ZN(new_n21066_));
  NOR2_X1    g20769(.A1(new_n21066_), .A2(new_n21060_), .ZN(new_n21067_));
  XOR2_X1    g20770(.A1(new_n21067_), .A2(new_n20926_), .Z(new_n21068_));
  NOR2_X1    g20771(.A1(new_n21067_), .A2(new_n20926_), .ZN(new_n21069_));
  INV_X1     g20772(.I(new_n21069_), .ZN(new_n21070_));
  NAND2_X1   g20773(.A1(new_n21067_), .A2(new_n20926_), .ZN(new_n21071_));
  AOI21_X1   g20774(.A1(new_n21070_), .A2(new_n21071_), .B(new_n20921_), .ZN(new_n21072_));
  AOI21_X1   g20775(.A1(new_n20921_), .A2(new_n21068_), .B(new_n21072_), .ZN(new_n21073_));
  NOR2_X1    g20776(.A1(new_n21073_), .A2(new_n20918_), .ZN(new_n21074_));
  NAND2_X1   g20777(.A1(new_n21073_), .A2(new_n20918_), .ZN(new_n21075_));
  INV_X1     g20778(.I(new_n21075_), .ZN(new_n21076_));
  OAI22_X1   g20779(.A1(new_n21076_), .A2(new_n21074_), .B1(new_n20881_), .B2(new_n20914_), .ZN(new_n21077_));
  NOR2_X1    g20780(.A1(new_n20914_), .A2(new_n20881_), .ZN(new_n21078_));
  XOR2_X1    g20781(.A1(new_n21073_), .A2(new_n20918_), .Z(new_n21079_));
  NAND2_X1   g20782(.A1(new_n21079_), .A2(new_n21078_), .ZN(new_n21080_));
  NAND2_X1   g20783(.A1(new_n21080_), .A2(new_n21077_), .ZN(new_n21081_));
  INV_X1     g20784(.I(new_n21081_), .ZN(new_n21082_));
  NOR2_X1    g20785(.A1(new_n21082_), .A2(new_n20913_), .ZN(new_n21083_));
  INV_X1     g20786(.I(new_n21083_), .ZN(new_n21084_));
  NAND2_X1   g20787(.A1(new_n21082_), .A2(new_n20913_), .ZN(new_n21085_));
  NAND2_X1   g20788(.A1(new_n21084_), .A2(new_n21085_), .ZN(new_n21086_));
  XOR2_X1    g20789(.A1(new_n21081_), .A2(new_n20913_), .Z(new_n21087_));
  NOR2_X1    g20790(.A1(new_n21087_), .A2(new_n20909_), .ZN(new_n21088_));
  AOI21_X1   g20791(.A1(new_n20909_), .A2(new_n21086_), .B(new_n21088_), .ZN(new_n21089_));
  XOR2_X1    g20792(.A1(new_n21089_), .A2(new_n20904_), .Z(new_n21090_));
  AOI21_X1   g20793(.A1(new_n20897_), .A2(new_n21090_), .B(new_n20899_), .ZN(new_n21091_));
  XOR2_X1    g20794(.A1(new_n20718_), .A2(new_n21091_), .Z(\f[87] ));
  NAND2_X1   g20795(.A1(new_n21089_), .A2(new_n20904_), .ZN(new_n21093_));
  NOR3_X1    g20796(.A1(new_n20298_), .A2(new_n20514_), .A3(new_n20717_), .ZN(new_n21094_));
  NOR2_X1    g20797(.A1(new_n20898_), .A2(new_n20896_), .ZN(new_n21095_));
  INV_X1     g20798(.I(new_n21095_), .ZN(new_n21096_));
  OAI21_X1   g20799(.A1(new_n21094_), .A2(new_n20714_), .B(new_n21096_), .ZN(new_n21097_));
  AOI21_X1   g20800(.A1(new_n20909_), .A2(new_n21085_), .B(new_n21083_), .ZN(new_n21098_));
  NOR2_X1    g20801(.A1(new_n2322_), .A2(new_n2166_), .ZN(new_n21099_));
  NAND2_X1   g20802(.A1(new_n16148_), .A2(new_n2168_), .ZN(new_n21100_));
  OAI21_X1   g20803(.A1(new_n21099_), .A2(new_n21100_), .B(new_n2161_), .ZN(new_n21101_));
  XNOR2_X1   g20804(.A1(new_n14978_), .A2(new_n21101_), .ZN(new_n21102_));
  OAI22_X1   g20805(.A1(new_n13367_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n13785_), .ZN(new_n21103_));
  OAI21_X1   g20806(.A1(new_n12970_), .A2(new_n2884_), .B(new_n21103_), .ZN(new_n21104_));
  AOI21_X1   g20807(.A1(new_n21104_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n21105_));
  XOR2_X1    g20808(.A1(new_n13784_), .A2(new_n21105_), .Z(new_n21106_));
  OAI21_X1   g20809(.A1(new_n20920_), .A2(new_n21069_), .B(new_n21071_), .ZN(new_n21107_));
  OAI22_X1   g20810(.A1(new_n12536_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n12542_), .ZN(new_n21108_));
  OAI21_X1   g20811(.A1(new_n11744_), .A2(new_n3569_), .B(new_n21108_), .ZN(new_n21109_));
  AOI21_X1   g20812(.A1(new_n21109_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n21110_));
  XNOR2_X1   g20813(.A1(new_n12546_), .A2(new_n21110_), .ZN(new_n21111_));
  AOI21_X1   g20814(.A1(new_n21061_), .A2(new_n21065_), .B(new_n21063_), .ZN(new_n21112_));
  NOR2_X1    g20815(.A1(new_n21050_), .A2(new_n20929_), .ZN(new_n21113_));
  NOR2_X1    g20816(.A1(new_n21113_), .A2(new_n21047_), .ZN(new_n21114_));
  OAI22_X1   g20817(.A1(new_n5420_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n5107_), .ZN(new_n21115_));
  OAI21_X1   g20818(.A1(new_n9295_), .A2(new_n5112_), .B(new_n21115_), .ZN(new_n21116_));
  AOI21_X1   g20819(.A1(new_n21116_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n21117_));
  XNOR2_X1   g20820(.A1(new_n10035_), .A2(new_n21117_), .ZN(new_n21118_));
  INV_X1     g20821(.I(new_n21118_), .ZN(new_n21119_));
  OAI22_X1   g20822(.A1(new_n6644_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n6647_), .ZN(new_n21120_));
  OAI21_X1   g20823(.A1(new_n7198_), .A2(new_n7284_), .B(new_n21120_), .ZN(new_n21121_));
  AOI21_X1   g20824(.A1(new_n21121_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n21122_));
  XNOR2_X1   g20825(.A1(new_n7874_), .A2(new_n21122_), .ZN(new_n21123_));
  AOI21_X1   g20826(.A1(new_n20933_), .A2(new_n21005_), .B(new_n21003_), .ZN(new_n21124_));
  OAI22_X1   g20827(.A1(new_n8644_), .A2(new_n5913_), .B1(new_n5921_), .B2(new_n9388_), .ZN(new_n21125_));
  OAI21_X1   g20828(.A1(new_n5353_), .A2(new_n10154_), .B(new_n21125_), .ZN(new_n21126_));
  AOI21_X1   g20829(.A1(new_n21126_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n21127_));
  XOR2_X1    g20830(.A1(new_n5926_), .A2(new_n21127_), .Z(new_n21128_));
  NAND2_X1   g20831(.A1(new_n20991_), .A2(new_n20980_), .ZN(new_n21129_));
  NAND2_X1   g20832(.A1(new_n21129_), .A2(new_n20987_), .ZN(new_n21130_));
  AOI22_X1   g20833(.A1(new_n10969_), .A2(new_n20556_), .B1(new_n11394_), .B2(\b[32] ), .ZN(new_n21131_));
  OAI21_X1   g20834(.A1(new_n21131_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n21132_));
  XOR2_X1    g20835(.A1(new_n4257_), .A2(new_n21132_), .Z(new_n21133_));
  OAI21_X1   g20836(.A1(new_n20938_), .A2(new_n20955_), .B(new_n20956_), .ZN(new_n21134_));
  OAI22_X1   g20837(.A1(new_n13880_), .A2(new_n2843_), .B1(new_n2439_), .B2(new_n13885_), .ZN(new_n21135_));
  AOI21_X1   g20838(.A1(new_n21135_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n21136_));
  XNOR2_X1   g20839(.A1(new_n2846_), .A2(new_n21136_), .ZN(new_n21137_));
  NAND2_X1   g20840(.A1(new_n20952_), .A2(new_n20776_), .ZN(new_n21138_));
  NAND2_X1   g20841(.A1(new_n21138_), .A2(new_n20951_), .ZN(new_n21139_));
  NOR2_X1    g20842(.A1(new_n13476_), .A2(new_n2102_), .ZN(new_n21140_));
  XOR2_X1    g20843(.A1(new_n14736_), .A2(new_n2102_), .Z(new_n21141_));
  NAND2_X1   g20844(.A1(new_n21141_), .A2(\b[25] ), .ZN(new_n21142_));
  XOR2_X1    g20845(.A1(new_n21142_), .A2(new_n21140_), .Z(new_n21143_));
  INV_X1     g20846(.I(new_n21143_), .ZN(new_n21144_));
  XOR2_X1    g20847(.A1(new_n21139_), .A2(new_n21144_), .Z(new_n21145_));
  NOR2_X1    g20848(.A1(new_n21139_), .A2(new_n21143_), .ZN(new_n21146_));
  INV_X1     g20849(.I(new_n21146_), .ZN(new_n21147_));
  NAND2_X1   g20850(.A1(new_n21139_), .A2(new_n21143_), .ZN(new_n21148_));
  NAND2_X1   g20851(.A1(new_n21147_), .A2(new_n21148_), .ZN(new_n21149_));
  NAND2_X1   g20852(.A1(new_n21137_), .A2(new_n21149_), .ZN(new_n21150_));
  OAI21_X1   g20853(.A1(new_n21137_), .A2(new_n21145_), .B(new_n21150_), .ZN(new_n21151_));
  AOI22_X1   g20854(.A1(new_n13078_), .A2(\b[29] ), .B1(new_n3711_), .B2(new_n12218_), .ZN(new_n21152_));
  OAI21_X1   g20855(.A1(new_n21152_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n21153_));
  XOR2_X1    g20856(.A1(new_n3514_), .A2(new_n21153_), .Z(new_n21154_));
  NOR2_X1    g20857(.A1(new_n21151_), .A2(new_n21154_), .ZN(new_n21155_));
  INV_X1     g20858(.I(new_n21155_), .ZN(new_n21156_));
  NAND2_X1   g20859(.A1(new_n21151_), .A2(new_n21154_), .ZN(new_n21157_));
  NAND2_X1   g20860(.A1(new_n21156_), .A2(new_n21157_), .ZN(new_n21158_));
  XNOR2_X1   g20861(.A1(new_n21151_), .A2(new_n21154_), .ZN(new_n21159_));
  NOR2_X1    g20862(.A1(new_n21159_), .A2(new_n21134_), .ZN(new_n21160_));
  AOI21_X1   g20863(.A1(new_n21134_), .A2(new_n21158_), .B(new_n21160_), .ZN(new_n21161_));
  NOR2_X1    g20864(.A1(new_n20968_), .A2(new_n20936_), .ZN(new_n21162_));
  NOR2_X1    g20865(.A1(new_n21162_), .A2(new_n20966_), .ZN(new_n21163_));
  NOR2_X1    g20866(.A1(new_n21161_), .A2(new_n21163_), .ZN(new_n21164_));
  INV_X1     g20867(.I(new_n21164_), .ZN(new_n21165_));
  NAND2_X1   g20868(.A1(new_n21161_), .A2(new_n21163_), .ZN(new_n21166_));
  AOI21_X1   g20869(.A1(new_n21165_), .A2(new_n21166_), .B(new_n21133_), .ZN(new_n21167_));
  INV_X1     g20870(.I(new_n21133_), .ZN(new_n21168_));
  XNOR2_X1   g20871(.A1(new_n21161_), .A2(new_n21163_), .ZN(new_n21169_));
  NOR2_X1    g20872(.A1(new_n21169_), .A2(new_n21168_), .ZN(new_n21170_));
  NOR2_X1    g20873(.A1(new_n21170_), .A2(new_n21167_), .ZN(new_n21171_));
  INV_X1     g20874(.I(new_n21171_), .ZN(new_n21172_));
  NAND2_X1   g20875(.A1(new_n20976_), .A2(new_n20978_), .ZN(new_n21173_));
  NAND2_X1   g20876(.A1(new_n21173_), .A2(new_n20977_), .ZN(new_n21174_));
  AOI22_X1   g20877(.A1(new_n11415_), .A2(new_n5349_), .B1(\b[35] ), .B2(new_n10145_), .ZN(new_n21175_));
  OAI21_X1   g20878(.A1(new_n21175_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n21176_));
  XNOR2_X1   g20879(.A1(new_n5067_), .A2(new_n21176_), .ZN(new_n21177_));
  XNOR2_X1   g20880(.A1(new_n21174_), .A2(new_n21177_), .ZN(new_n21178_));
  INV_X1     g20881(.I(new_n21174_), .ZN(new_n21179_));
  NOR2_X1    g20882(.A1(new_n21179_), .A2(new_n21177_), .ZN(new_n21180_));
  INV_X1     g20883(.I(new_n21180_), .ZN(new_n21181_));
  NAND2_X1   g20884(.A1(new_n21179_), .A2(new_n21177_), .ZN(new_n21182_));
  AOI21_X1   g20885(.A1(new_n21181_), .A2(new_n21182_), .B(new_n21172_), .ZN(new_n21183_));
  AOI21_X1   g20886(.A1(new_n21172_), .A2(new_n21178_), .B(new_n21183_), .ZN(new_n21184_));
  XNOR2_X1   g20887(.A1(new_n21130_), .A2(new_n21184_), .ZN(new_n21185_));
  NOR2_X1    g20888(.A1(new_n21130_), .A2(new_n21184_), .ZN(new_n21186_));
  NAND2_X1   g20889(.A1(new_n21130_), .A2(new_n21184_), .ZN(new_n21187_));
  INV_X1     g20890(.I(new_n21187_), .ZN(new_n21188_));
  OAI21_X1   g20891(.A1(new_n21188_), .A2(new_n21186_), .B(new_n21128_), .ZN(new_n21189_));
  OAI21_X1   g20892(.A1(new_n21128_), .A2(new_n21185_), .B(new_n21189_), .ZN(new_n21190_));
  OAI22_X1   g20893(.A1(new_n7619_), .A2(new_n6538_), .B1(new_n6847_), .B2(new_n8309_), .ZN(new_n21191_));
  OAI21_X1   g20894(.A1(new_n6229_), .A2(new_n7947_), .B(new_n21191_), .ZN(new_n21192_));
  AOI21_X1   g20895(.A1(new_n21192_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n21193_));
  XOR2_X1    g20896(.A1(new_n6851_), .A2(new_n21193_), .Z(new_n21194_));
  NOR2_X1    g20897(.A1(new_n21190_), .A2(new_n21194_), .ZN(new_n21195_));
  INV_X1     g20898(.I(new_n21195_), .ZN(new_n21196_));
  NAND2_X1   g20899(.A1(new_n21190_), .A2(new_n21194_), .ZN(new_n21197_));
  AOI21_X1   g20900(.A1(new_n21196_), .A2(new_n21197_), .B(new_n21124_), .ZN(new_n21198_));
  INV_X1     g20901(.I(new_n21124_), .ZN(new_n21199_));
  XNOR2_X1   g20902(.A1(new_n21190_), .A2(new_n21194_), .ZN(new_n21200_));
  NOR2_X1    g20903(.A1(new_n21200_), .A2(new_n21199_), .ZN(new_n21201_));
  NOR2_X1    g20904(.A1(new_n21201_), .A2(new_n21198_), .ZN(new_n21202_));
  INV_X1     g20905(.I(new_n20932_), .ZN(new_n21203_));
  AOI21_X1   g20906(.A1(new_n21203_), .A2(new_n21015_), .B(new_n21013_), .ZN(new_n21204_));
  NOR2_X1    g20907(.A1(new_n21202_), .A2(new_n21204_), .ZN(new_n21205_));
  INV_X1     g20908(.I(new_n21205_), .ZN(new_n21206_));
  NAND2_X1   g20909(.A1(new_n21202_), .A2(new_n21204_), .ZN(new_n21207_));
  AOI21_X1   g20910(.A1(new_n21206_), .A2(new_n21207_), .B(new_n21123_), .ZN(new_n21208_));
  INV_X1     g20911(.I(new_n21123_), .ZN(new_n21209_));
  XNOR2_X1   g20912(.A1(new_n21202_), .A2(new_n21204_), .ZN(new_n21210_));
  NOR2_X1    g20913(.A1(new_n21210_), .A2(new_n21209_), .ZN(new_n21211_));
  NOR2_X1    g20914(.A1(new_n21211_), .A2(new_n21208_), .ZN(new_n21212_));
  NAND2_X1   g20915(.A1(new_n21028_), .A2(new_n21025_), .ZN(new_n21213_));
  NAND2_X1   g20916(.A1(new_n21213_), .A2(new_n21027_), .ZN(new_n21214_));
  INV_X1     g20917(.I(new_n21214_), .ZN(new_n21215_));
  OAI22_X1   g20918(.A1(new_n5993_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n5991_), .ZN(new_n21216_));
  OAI21_X1   g20919(.A1(new_n8218_), .A2(new_n5997_), .B(new_n21216_), .ZN(new_n21217_));
  AOI21_X1   g20920(.A1(new_n21217_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n21218_));
  XOR2_X1    g20921(.A1(new_n8952_), .A2(new_n21218_), .Z(new_n21219_));
  NOR2_X1    g20922(.A1(new_n21215_), .A2(new_n21219_), .ZN(new_n21220_));
  INV_X1     g20923(.I(new_n21219_), .ZN(new_n21221_));
  NOR2_X1    g20924(.A1(new_n21214_), .A2(new_n21221_), .ZN(new_n21222_));
  NOR2_X1    g20925(.A1(new_n21220_), .A2(new_n21222_), .ZN(new_n21223_));
  NOR2_X1    g20926(.A1(new_n21223_), .A2(new_n21212_), .ZN(new_n21224_));
  INV_X1     g20927(.I(new_n21212_), .ZN(new_n21225_));
  XOR2_X1    g20928(.A1(new_n21214_), .A2(new_n21219_), .Z(new_n21226_));
  NOR2_X1    g20929(.A1(new_n21226_), .A2(new_n21225_), .ZN(new_n21227_));
  NOR2_X1    g20930(.A1(new_n21224_), .A2(new_n21227_), .ZN(new_n21228_));
  NAND2_X1   g20931(.A1(new_n21030_), .A2(new_n21039_), .ZN(new_n21229_));
  AOI21_X1   g20932(.A1(new_n21037_), .A2(new_n21229_), .B(new_n21228_), .ZN(new_n21230_));
  NAND2_X1   g20933(.A1(new_n21229_), .A2(new_n21037_), .ZN(new_n21231_));
  NOR3_X1    g20934(.A1(new_n21231_), .A2(new_n21224_), .A3(new_n21227_), .ZN(new_n21232_));
  OAI21_X1   g20935(.A1(new_n21230_), .A2(new_n21232_), .B(new_n21119_), .ZN(new_n21233_));
  XNOR2_X1   g20936(.A1(new_n21228_), .A2(new_n21231_), .ZN(new_n21234_));
  NAND2_X1   g20937(.A1(new_n21234_), .A2(new_n21118_), .ZN(new_n21235_));
  NAND2_X1   g20938(.A1(new_n21235_), .A2(new_n21233_), .ZN(new_n21236_));
  OAI22_X1   g20939(.A1(new_n4072_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n4067_), .ZN(new_n21237_));
  OAI21_X1   g20940(.A1(new_n10477_), .A2(new_n4318_), .B(new_n21237_), .ZN(new_n21238_));
  AOI21_X1   g20941(.A1(new_n21238_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n21239_));
  XOR2_X1    g20942(.A1(new_n11298_), .A2(new_n21239_), .Z(new_n21240_));
  XOR2_X1    g20943(.A1(new_n21236_), .A2(new_n21240_), .Z(new_n21241_));
  NOR2_X1    g20944(.A1(new_n21241_), .A2(new_n21114_), .ZN(new_n21242_));
  INV_X1     g20945(.I(new_n21114_), .ZN(new_n21243_));
  INV_X1     g20946(.I(new_n21236_), .ZN(new_n21244_));
  NOR2_X1    g20947(.A1(new_n21244_), .A2(new_n21240_), .ZN(new_n21245_));
  INV_X1     g20948(.I(new_n21245_), .ZN(new_n21246_));
  NAND2_X1   g20949(.A1(new_n21244_), .A2(new_n21240_), .ZN(new_n21247_));
  AOI21_X1   g20950(.A1(new_n21246_), .A2(new_n21247_), .B(new_n21243_), .ZN(new_n21248_));
  NOR2_X1    g20951(.A1(new_n21248_), .A2(new_n21242_), .ZN(new_n21249_));
  XOR2_X1    g20952(.A1(new_n21249_), .A2(new_n21112_), .Z(new_n21250_));
  NOR2_X1    g20953(.A1(new_n21250_), .A2(new_n21111_), .ZN(new_n21251_));
  INV_X1     g20954(.I(new_n21111_), .ZN(new_n21252_));
  INV_X1     g20955(.I(new_n21112_), .ZN(new_n21253_));
  NOR2_X1    g20956(.A1(new_n21249_), .A2(new_n21253_), .ZN(new_n21254_));
  INV_X1     g20957(.I(new_n21254_), .ZN(new_n21255_));
  NAND2_X1   g20958(.A1(new_n21249_), .A2(new_n21253_), .ZN(new_n21256_));
  AOI21_X1   g20959(.A1(new_n21255_), .A2(new_n21256_), .B(new_n21252_), .ZN(new_n21257_));
  NOR2_X1    g20960(.A1(new_n21251_), .A2(new_n21257_), .ZN(new_n21258_));
  NOR2_X1    g20961(.A1(new_n21258_), .A2(new_n21107_), .ZN(new_n21259_));
  INV_X1     g20962(.I(new_n21107_), .ZN(new_n21260_));
  INV_X1     g20963(.I(new_n21258_), .ZN(new_n21261_));
  NOR2_X1    g20964(.A1(new_n21261_), .A2(new_n21260_), .ZN(new_n21262_));
  NOR2_X1    g20965(.A1(new_n21262_), .A2(new_n21259_), .ZN(new_n21263_));
  NOR2_X1    g20966(.A1(new_n21263_), .A2(new_n21106_), .ZN(new_n21264_));
  INV_X1     g20967(.I(new_n21106_), .ZN(new_n21265_));
  XOR2_X1    g20968(.A1(new_n21258_), .A2(new_n21260_), .Z(new_n21266_));
  NOR2_X1    g20969(.A1(new_n21266_), .A2(new_n21265_), .ZN(new_n21267_));
  NOR2_X1    g20970(.A1(new_n21264_), .A2(new_n21267_), .ZN(new_n21268_));
  OAI21_X1   g20971(.A1(new_n21078_), .A2(new_n21074_), .B(new_n21075_), .ZN(new_n21269_));
  XOR2_X1    g20972(.A1(new_n21268_), .A2(new_n21269_), .Z(new_n21270_));
  NOR2_X1    g20973(.A1(new_n21270_), .A2(new_n21102_), .ZN(new_n21271_));
  INV_X1     g20974(.I(new_n21102_), .ZN(new_n21272_));
  INV_X1     g20975(.I(new_n21269_), .ZN(new_n21273_));
  NOR2_X1    g20976(.A1(new_n21268_), .A2(new_n21273_), .ZN(new_n21274_));
  INV_X1     g20977(.I(new_n21274_), .ZN(new_n21275_));
  NAND2_X1   g20978(.A1(new_n21268_), .A2(new_n21273_), .ZN(new_n21276_));
  AOI21_X1   g20979(.A1(new_n21275_), .A2(new_n21276_), .B(new_n21272_), .ZN(new_n21277_));
  NOR2_X1    g20980(.A1(new_n21271_), .A2(new_n21277_), .ZN(new_n21278_));
  NOR2_X1    g20981(.A1(new_n21278_), .A2(new_n21098_), .ZN(new_n21279_));
  XOR2_X1    g20982(.A1(new_n21097_), .A2(new_n21279_), .Z(new_n21280_));
  XOR2_X1    g20983(.A1(new_n21280_), .A2(new_n21093_), .Z(\f[88] ));
  INV_X1     g20984(.I(new_n21279_), .ZN(new_n21282_));
  AOI21_X1   g20985(.A1(new_n21098_), .A2(new_n21278_), .B(new_n21093_), .ZN(new_n21283_));
  INV_X1     g20986(.I(new_n21283_), .ZN(new_n21284_));
  OAI21_X1   g20987(.A1(new_n21097_), .A2(new_n21284_), .B(new_n21282_), .ZN(new_n21285_));
  AOI21_X1   g20988(.A1(new_n21272_), .A2(new_n21276_), .B(new_n21274_), .ZN(new_n21286_));
  INV_X1     g20989(.I(new_n21286_), .ZN(new_n21287_));
  OAI22_X1   g20990(.A1(new_n13785_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n14208_), .ZN(new_n21288_));
  OAI21_X1   g20991(.A1(new_n13367_), .A2(new_n2884_), .B(new_n21288_), .ZN(new_n21289_));
  AOI21_X1   g20992(.A1(new_n21289_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n21290_));
  XOR2_X1    g20993(.A1(new_n14213_), .A2(new_n21290_), .Z(new_n21291_));
  INV_X1     g20994(.I(new_n21291_), .ZN(new_n21292_));
  OAI21_X1   g20995(.A1(new_n21111_), .A2(new_n21254_), .B(new_n21256_), .ZN(new_n21293_));
  OAI22_X1   g20996(.A1(new_n12542_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n12970_), .ZN(new_n21294_));
  OAI21_X1   g20997(.A1(new_n12536_), .A2(new_n3569_), .B(new_n21294_), .ZN(new_n21295_));
  AOI21_X1   g20998(.A1(new_n21295_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n21296_));
  XOR2_X1    g20999(.A1(new_n12969_), .A2(new_n21296_), .Z(new_n21297_));
  INV_X1     g21000(.I(new_n21297_), .ZN(new_n21298_));
  OAI22_X1   g21001(.A1(new_n4072_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n4067_), .ZN(new_n21299_));
  OAI21_X1   g21002(.A1(new_n10862_), .A2(new_n4318_), .B(new_n21299_), .ZN(new_n21300_));
  AOI21_X1   g21003(.A1(new_n21300_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n21301_));
  XNOR2_X1   g21004(.A1(new_n11748_), .A2(new_n21301_), .ZN(new_n21302_));
  NOR2_X1    g21005(.A1(new_n21232_), .A2(new_n21118_), .ZN(new_n21303_));
  OAI22_X1   g21006(.A1(new_n5420_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n5107_), .ZN(new_n21304_));
  OAI21_X1   g21007(.A1(new_n10025_), .A2(new_n5112_), .B(new_n21304_), .ZN(new_n21305_));
  AOI21_X1   g21008(.A1(new_n21305_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n21306_));
  XOR2_X1    g21009(.A1(new_n10476_), .A2(new_n21306_), .Z(new_n21307_));
  OAI22_X1   g21010(.A1(new_n5993_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n5991_), .ZN(new_n21308_));
  OAI21_X1   g21011(.A1(new_n8563_), .A2(new_n5997_), .B(new_n21308_), .ZN(new_n21309_));
  AOI21_X1   g21012(.A1(new_n21309_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n21310_));
  XNOR2_X1   g21013(.A1(new_n9299_), .A2(new_n21310_), .ZN(new_n21311_));
  OAI22_X1   g21014(.A1(new_n7619_), .A2(new_n6847_), .B1(new_n7198_), .B2(new_n8309_), .ZN(new_n21312_));
  OAI21_X1   g21015(.A1(new_n6538_), .A2(new_n7947_), .B(new_n21312_), .ZN(new_n21313_));
  AOI21_X1   g21016(.A1(new_n21313_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n21314_));
  XNOR2_X1   g21017(.A1(new_n7202_), .A2(new_n21314_), .ZN(new_n21315_));
  OAI21_X1   g21018(.A1(new_n21128_), .A2(new_n21186_), .B(new_n21187_), .ZN(new_n21316_));
  INV_X1     g21019(.I(new_n5354_), .ZN(new_n21317_));
  AOI22_X1   g21020(.A1(new_n11415_), .A2(new_n21317_), .B1(\b[36] ), .B2(new_n10145_), .ZN(new_n21318_));
  OAI21_X1   g21021(.A1(new_n21318_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n21319_));
  XOR2_X1    g21022(.A1(new_n5357_), .A2(new_n21319_), .Z(new_n21320_));
  AOI21_X1   g21023(.A1(new_n21168_), .A2(new_n21166_), .B(new_n21164_), .ZN(new_n21321_));
  INV_X1     g21024(.I(new_n21321_), .ZN(new_n21322_));
  AOI22_X1   g21025(.A1(new_n10969_), .A2(new_n4770_), .B1(new_n11394_), .B2(\b[33] ), .ZN(new_n21323_));
  OAI21_X1   g21026(.A1(new_n21323_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n21324_));
  XNOR2_X1   g21027(.A1(new_n4499_), .A2(new_n21324_), .ZN(new_n21325_));
  AOI22_X1   g21028(.A1(new_n13078_), .A2(\b[30] ), .B1(new_n3719_), .B2(new_n12218_), .ZN(new_n21326_));
  OAI21_X1   g21029(.A1(new_n21326_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n21327_));
  XNOR2_X1   g21030(.A1(new_n3722_), .A2(new_n21327_), .ZN(new_n21328_));
  OR2_X2     g21031(.A1(new_n21137_), .A2(new_n21146_), .Z(new_n21329_));
  NAND2_X1   g21032(.A1(new_n21329_), .A2(new_n21148_), .ZN(new_n21330_));
  OAI22_X1   g21033(.A1(new_n13880_), .A2(new_n3255_), .B1(new_n2643_), .B2(new_n13885_), .ZN(new_n21331_));
  AOI21_X1   g21034(.A1(new_n21331_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n21332_));
  XNOR2_X1   g21035(.A1(new_n3022_), .A2(new_n21332_), .ZN(new_n21333_));
  NOR2_X1    g21036(.A1(new_n13476_), .A2(new_n2281_), .ZN(new_n21334_));
  XOR2_X1    g21037(.A1(new_n14736_), .A2(new_n2281_), .Z(new_n21335_));
  NAND2_X1   g21038(.A1(new_n21335_), .A2(\b[26] ), .ZN(new_n21336_));
  XOR2_X1    g21039(.A1(new_n21336_), .A2(new_n21334_), .Z(new_n21337_));
  XOR2_X1    g21040(.A1(new_n21143_), .A2(new_n21337_), .Z(new_n21338_));
  NOR2_X1    g21041(.A1(new_n21144_), .A2(new_n21337_), .ZN(new_n21339_));
  INV_X1     g21042(.I(new_n21337_), .ZN(new_n21340_));
  NOR2_X1    g21043(.A1(new_n21340_), .A2(new_n21143_), .ZN(new_n21341_));
  OAI21_X1   g21044(.A1(new_n21339_), .A2(new_n21341_), .B(new_n21333_), .ZN(new_n21342_));
  OAI21_X1   g21045(.A1(new_n21333_), .A2(new_n21338_), .B(new_n21342_), .ZN(new_n21343_));
  XOR2_X1    g21046(.A1(new_n21330_), .A2(new_n21343_), .Z(new_n21344_));
  NOR2_X1    g21047(.A1(new_n21328_), .A2(new_n21344_), .ZN(new_n21345_));
  INV_X1     g21048(.I(new_n21328_), .ZN(new_n21346_));
  INV_X1     g21049(.I(new_n21330_), .ZN(new_n21347_));
  NAND2_X1   g21050(.A1(new_n21347_), .A2(new_n21343_), .ZN(new_n21348_));
  NOR2_X1    g21051(.A1(new_n21347_), .A2(new_n21343_), .ZN(new_n21349_));
  INV_X1     g21052(.I(new_n21349_), .ZN(new_n21350_));
  AOI21_X1   g21053(.A1(new_n21348_), .A2(new_n21350_), .B(new_n21346_), .ZN(new_n21351_));
  NOR2_X1    g21054(.A1(new_n21351_), .A2(new_n21345_), .ZN(new_n21352_));
  AOI21_X1   g21055(.A1(new_n21134_), .A2(new_n21157_), .B(new_n21155_), .ZN(new_n21353_));
  XOR2_X1    g21056(.A1(new_n21352_), .A2(new_n21353_), .Z(new_n21354_));
  NOR2_X1    g21057(.A1(new_n21354_), .A2(new_n21325_), .ZN(new_n21355_));
  INV_X1     g21058(.I(new_n21325_), .ZN(new_n21356_));
  INV_X1     g21059(.I(new_n21352_), .ZN(new_n21357_));
  NOR2_X1    g21060(.A1(new_n21357_), .A2(new_n21353_), .ZN(new_n21358_));
  INV_X1     g21061(.I(new_n21358_), .ZN(new_n21359_));
  NAND2_X1   g21062(.A1(new_n21357_), .A2(new_n21353_), .ZN(new_n21360_));
  AOI21_X1   g21063(.A1(new_n21359_), .A2(new_n21360_), .B(new_n21356_), .ZN(new_n21361_));
  NOR2_X1    g21064(.A1(new_n21361_), .A2(new_n21355_), .ZN(new_n21362_));
  NOR2_X1    g21065(.A1(new_n21362_), .A2(new_n21322_), .ZN(new_n21363_));
  INV_X1     g21066(.I(new_n21362_), .ZN(new_n21364_));
  NOR2_X1    g21067(.A1(new_n21364_), .A2(new_n21321_), .ZN(new_n21365_));
  NOR2_X1    g21068(.A1(new_n21365_), .A2(new_n21363_), .ZN(new_n21366_));
  NOR2_X1    g21069(.A1(new_n21366_), .A2(new_n21320_), .ZN(new_n21367_));
  INV_X1     g21070(.I(new_n21320_), .ZN(new_n21368_));
  XOR2_X1    g21071(.A1(new_n21362_), .A2(new_n21321_), .Z(new_n21369_));
  NOR2_X1    g21072(.A1(new_n21369_), .A2(new_n21368_), .ZN(new_n21370_));
  NOR2_X1    g21073(.A1(new_n21367_), .A2(new_n21370_), .ZN(new_n21371_));
  OAI22_X1   g21074(.A1(new_n8644_), .A2(new_n5921_), .B1(new_n6229_), .B2(new_n9388_), .ZN(new_n21372_));
  OAI21_X1   g21075(.A1(new_n5913_), .A2(new_n10154_), .B(new_n21372_), .ZN(new_n21373_));
  AOI21_X1   g21076(.A1(new_n21373_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n21374_));
  XOR2_X1    g21077(.A1(new_n6233_), .A2(new_n21374_), .Z(new_n21375_));
  AOI21_X1   g21078(.A1(new_n21172_), .A2(new_n21182_), .B(new_n21180_), .ZN(new_n21376_));
  NOR2_X1    g21079(.A1(new_n21376_), .A2(new_n21375_), .ZN(new_n21377_));
  AND2_X2    g21080(.A1(new_n21376_), .A2(new_n21375_), .Z(new_n21378_));
  NOR2_X1    g21081(.A1(new_n21378_), .A2(new_n21377_), .ZN(new_n21379_));
  NOR2_X1    g21082(.A1(new_n21371_), .A2(new_n21379_), .ZN(new_n21380_));
  INV_X1     g21083(.I(new_n21371_), .ZN(new_n21381_));
  XNOR2_X1   g21084(.A1(new_n21376_), .A2(new_n21375_), .ZN(new_n21382_));
  NOR2_X1    g21085(.A1(new_n21381_), .A2(new_n21382_), .ZN(new_n21383_));
  NOR2_X1    g21086(.A1(new_n21383_), .A2(new_n21380_), .ZN(new_n21384_));
  XOR2_X1    g21087(.A1(new_n21384_), .A2(new_n21316_), .Z(new_n21385_));
  INV_X1     g21088(.I(new_n21316_), .ZN(new_n21386_));
  NOR2_X1    g21089(.A1(new_n21384_), .A2(new_n21386_), .ZN(new_n21387_));
  NOR3_X1    g21090(.A1(new_n21383_), .A2(new_n21316_), .A3(new_n21380_), .ZN(new_n21388_));
  OAI21_X1   g21091(.A1(new_n21387_), .A2(new_n21388_), .B(new_n21315_), .ZN(new_n21389_));
  OAI21_X1   g21092(.A1(new_n21315_), .A2(new_n21385_), .B(new_n21389_), .ZN(new_n21390_));
  OAI22_X1   g21093(.A1(new_n6644_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n6647_), .ZN(new_n21391_));
  OAI21_X1   g21094(.A1(new_n7864_), .A2(new_n7284_), .B(new_n21391_), .ZN(new_n21392_));
  AOI21_X1   g21095(.A1(new_n21392_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n21393_));
  XOR2_X1    g21096(.A1(new_n8217_), .A2(new_n21393_), .Z(new_n21394_));
  AOI21_X1   g21097(.A1(new_n21199_), .A2(new_n21197_), .B(new_n21195_), .ZN(new_n21395_));
  XOR2_X1    g21098(.A1(new_n21395_), .A2(new_n21394_), .Z(new_n21396_));
  NOR2_X1    g21099(.A1(new_n21395_), .A2(new_n21394_), .ZN(new_n21397_));
  INV_X1     g21100(.I(new_n21397_), .ZN(new_n21398_));
  NAND2_X1   g21101(.A1(new_n21395_), .A2(new_n21394_), .ZN(new_n21399_));
  AOI21_X1   g21102(.A1(new_n21398_), .A2(new_n21399_), .B(new_n21390_), .ZN(new_n21400_));
  AOI21_X1   g21103(.A1(new_n21390_), .A2(new_n21396_), .B(new_n21400_), .ZN(new_n21401_));
  AOI21_X1   g21104(.A1(new_n21209_), .A2(new_n21207_), .B(new_n21205_), .ZN(new_n21402_));
  XNOR2_X1   g21105(.A1(new_n21402_), .A2(new_n21401_), .ZN(new_n21403_));
  NOR2_X1    g21106(.A1(new_n21403_), .A2(new_n21311_), .ZN(new_n21404_));
  INV_X1     g21107(.I(new_n21311_), .ZN(new_n21405_));
  NOR2_X1    g21108(.A1(new_n21402_), .A2(new_n21401_), .ZN(new_n21406_));
  INV_X1     g21109(.I(new_n21406_), .ZN(new_n21407_));
  NAND2_X1   g21110(.A1(new_n21402_), .A2(new_n21401_), .ZN(new_n21408_));
  AOI21_X1   g21111(.A1(new_n21407_), .A2(new_n21408_), .B(new_n21405_), .ZN(new_n21409_));
  NOR2_X1    g21112(.A1(new_n21404_), .A2(new_n21409_), .ZN(new_n21410_));
  NOR2_X1    g21113(.A1(new_n21222_), .A2(new_n21212_), .ZN(new_n21411_));
  NOR2_X1    g21114(.A1(new_n21411_), .A2(new_n21220_), .ZN(new_n21412_));
  XOR2_X1    g21115(.A1(new_n21412_), .A2(new_n21410_), .Z(new_n21413_));
  NOR2_X1    g21116(.A1(new_n21413_), .A2(new_n21307_), .ZN(new_n21414_));
  INV_X1     g21117(.I(new_n21307_), .ZN(new_n21415_));
  INV_X1     g21118(.I(new_n21410_), .ZN(new_n21416_));
  NOR2_X1    g21119(.A1(new_n21416_), .A2(new_n21412_), .ZN(new_n21417_));
  INV_X1     g21120(.I(new_n21417_), .ZN(new_n21418_));
  NAND2_X1   g21121(.A1(new_n21416_), .A2(new_n21412_), .ZN(new_n21419_));
  AOI21_X1   g21122(.A1(new_n21418_), .A2(new_n21419_), .B(new_n21415_), .ZN(new_n21420_));
  NOR2_X1    g21123(.A1(new_n21414_), .A2(new_n21420_), .ZN(new_n21421_));
  NOR3_X1    g21124(.A1(new_n21421_), .A2(new_n21230_), .A3(new_n21303_), .ZN(new_n21422_));
  NOR2_X1    g21125(.A1(new_n21230_), .A2(new_n21303_), .ZN(new_n21423_));
  INV_X1     g21126(.I(new_n21421_), .ZN(new_n21424_));
  NOR2_X1    g21127(.A1(new_n21424_), .A2(new_n21423_), .ZN(new_n21425_));
  NOR2_X1    g21128(.A1(new_n21425_), .A2(new_n21422_), .ZN(new_n21426_));
  NOR2_X1    g21129(.A1(new_n21426_), .A2(new_n21302_), .ZN(new_n21427_));
  INV_X1     g21130(.I(new_n21302_), .ZN(new_n21428_));
  XOR2_X1    g21131(.A1(new_n21421_), .A2(new_n21423_), .Z(new_n21429_));
  NOR2_X1    g21132(.A1(new_n21429_), .A2(new_n21428_), .ZN(new_n21430_));
  NOR2_X1    g21133(.A1(new_n21427_), .A2(new_n21430_), .ZN(new_n21431_));
  AOI21_X1   g21134(.A1(new_n21243_), .A2(new_n21247_), .B(new_n21245_), .ZN(new_n21432_));
  NOR2_X1    g21135(.A1(new_n21432_), .A2(new_n21431_), .ZN(new_n21433_));
  INV_X1     g21136(.I(new_n21431_), .ZN(new_n21434_));
  INV_X1     g21137(.I(new_n21432_), .ZN(new_n21435_));
  NOR2_X1    g21138(.A1(new_n21435_), .A2(new_n21434_), .ZN(new_n21436_));
  OAI21_X1   g21139(.A1(new_n21436_), .A2(new_n21433_), .B(new_n21298_), .ZN(new_n21437_));
  XNOR2_X1   g21140(.A1(new_n21432_), .A2(new_n21431_), .ZN(new_n21438_));
  OAI21_X1   g21141(.A1(new_n21298_), .A2(new_n21438_), .B(new_n21437_), .ZN(new_n21439_));
  XOR2_X1    g21142(.A1(new_n21439_), .A2(new_n21293_), .Z(new_n21440_));
  NAND2_X1   g21143(.A1(new_n21440_), .A2(new_n21292_), .ZN(new_n21441_));
  AND2_X2    g21144(.A1(new_n21439_), .A2(new_n21293_), .Z(new_n21442_));
  NOR2_X1    g21145(.A1(new_n21439_), .A2(new_n21293_), .ZN(new_n21443_));
  OAI21_X1   g21146(.A1(new_n21442_), .A2(new_n21443_), .B(new_n21291_), .ZN(new_n21444_));
  NAND2_X1   g21147(.A1(new_n21441_), .A2(new_n21444_), .ZN(new_n21445_));
  OAI21_X1   g21148(.A1(new_n2171_), .A2(new_n2322_), .B(new_n16487_), .ZN(new_n21446_));
  NOR2_X1    g21149(.A1(new_n21259_), .A2(new_n21106_), .ZN(new_n21447_));
  NOR2_X1    g21150(.A1(new_n21447_), .A2(new_n21262_), .ZN(new_n21448_));
  XOR2_X1    g21151(.A1(new_n21448_), .A2(new_n21446_), .Z(new_n21449_));
  XOR2_X1    g21152(.A1(new_n21449_), .A2(new_n21445_), .Z(new_n21450_));
  NOR2_X1    g21153(.A1(new_n21450_), .A2(\a[26] ), .ZN(new_n21451_));
  NAND2_X1   g21154(.A1(new_n21450_), .A2(\a[26] ), .ZN(new_n21452_));
  INV_X1     g21155(.I(new_n21452_), .ZN(new_n21453_));
  NOR2_X1    g21156(.A1(new_n21453_), .A2(new_n21451_), .ZN(new_n21454_));
  INV_X1     g21157(.I(new_n21454_), .ZN(new_n21455_));
  NAND2_X1   g21158(.A1(new_n21455_), .A2(new_n21287_), .ZN(new_n21456_));
  NAND2_X1   g21159(.A1(new_n21454_), .A2(new_n21286_), .ZN(new_n21457_));
  NAND2_X1   g21160(.A1(new_n21456_), .A2(new_n21457_), .ZN(new_n21458_));
  XOR2_X1    g21161(.A1(new_n21454_), .A2(new_n21286_), .Z(new_n21459_));
  MUX2_X1    g21162(.I0(new_n21459_), .I1(new_n21458_), .S(new_n21285_), .Z(\f[89] ));
  INV_X1     g21163(.I(new_n21445_), .ZN(new_n21461_));
  NAND2_X1   g21164(.A1(new_n21461_), .A2(new_n21448_), .ZN(new_n21462_));
  XOR2_X1    g21165(.A1(new_n21446_), .A2(\a[26] ), .Z(new_n21463_));
  NAND2_X1   g21166(.A1(new_n21462_), .A2(new_n21463_), .ZN(new_n21464_));
  OAI21_X1   g21167(.A1(new_n21461_), .A2(new_n21448_), .B(new_n21464_), .ZN(new_n21465_));
  NOR2_X1    g21168(.A1(new_n21443_), .A2(new_n21291_), .ZN(new_n21466_));
  NOR2_X1    g21169(.A1(new_n21466_), .A2(new_n21442_), .ZN(new_n21467_));
  OAI22_X1   g21170(.A1(new_n14208_), .A2(new_n2705_), .B1(new_n2700_), .B2(new_n14592_), .ZN(new_n21468_));
  OAI21_X1   g21171(.A1(new_n13785_), .A2(new_n2884_), .B(new_n21468_), .ZN(new_n21469_));
  AOI21_X1   g21172(.A1(new_n21469_), .A2(new_n2702_), .B(new_n2705_), .ZN(new_n21470_));
  XNOR2_X1   g21173(.A1(new_n14599_), .A2(new_n21470_), .ZN(new_n21471_));
  NOR2_X1    g21174(.A1(new_n21422_), .A2(new_n21302_), .ZN(new_n21472_));
  NOR2_X1    g21175(.A1(new_n21472_), .A2(new_n21425_), .ZN(new_n21473_));
  INV_X1     g21176(.I(new_n21473_), .ZN(new_n21474_));
  AOI21_X1   g21177(.A1(new_n21415_), .A2(new_n21419_), .B(new_n21417_), .ZN(new_n21475_));
  AOI21_X1   g21178(.A1(new_n21405_), .A2(new_n21408_), .B(new_n21406_), .ZN(new_n21476_));
  INV_X1     g21179(.I(new_n21476_), .ZN(new_n21477_));
  INV_X1     g21180(.I(new_n21387_), .ZN(new_n21478_));
  OAI21_X1   g21181(.A1(new_n21315_), .A2(new_n21388_), .B(new_n21478_), .ZN(new_n21479_));
  INV_X1     g21182(.I(new_n21378_), .ZN(new_n21480_));
  AOI21_X1   g21183(.A1(new_n21381_), .A2(new_n21480_), .B(new_n21377_), .ZN(new_n21481_));
  INV_X1     g21184(.I(new_n21363_), .ZN(new_n21482_));
  AOI21_X1   g21185(.A1(new_n21368_), .A2(new_n21482_), .B(new_n21365_), .ZN(new_n21483_));
  AOI21_X1   g21186(.A1(new_n21346_), .A2(new_n21348_), .B(new_n21349_), .ZN(new_n21484_));
  AOI22_X1   g21187(.A1(new_n13078_), .A2(\b[31] ), .B1(new_n4249_), .B2(new_n12218_), .ZN(new_n21485_));
  OAI21_X1   g21188(.A1(new_n21485_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n21486_));
  XOR2_X1    g21189(.A1(new_n3993_), .A2(new_n21486_), .Z(new_n21487_));
  NOR2_X1    g21190(.A1(new_n21333_), .A2(new_n21339_), .ZN(new_n21488_));
  NOR2_X1    g21191(.A1(new_n21488_), .A2(new_n21341_), .ZN(new_n21489_));
  OAI22_X1   g21192(.A1(new_n13880_), .A2(new_n3261_), .B1(new_n2842_), .B2(new_n13885_), .ZN(new_n21490_));
  AOI21_X1   g21193(.A1(new_n21490_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n21491_));
  XNOR2_X1   g21194(.A1(new_n3264_), .A2(new_n21491_), .ZN(new_n21492_));
  INV_X1     g21195(.I(new_n21492_), .ZN(new_n21493_));
  NOR2_X1    g21196(.A1(new_n13476_), .A2(new_n2439_), .ZN(new_n21494_));
  XOR2_X1    g21197(.A1(new_n14736_), .A2(new_n2439_), .Z(new_n21495_));
  NAND2_X1   g21198(.A1(new_n21495_), .A2(\b[27] ), .ZN(new_n21496_));
  XOR2_X1    g21199(.A1(new_n21496_), .A2(new_n21494_), .Z(new_n21497_));
  XOR2_X1    g21200(.A1(new_n21497_), .A2(\a[26] ), .Z(new_n21498_));
  NOR2_X1    g21201(.A1(new_n21498_), .A2(new_n21337_), .ZN(new_n21499_));
  NOR2_X1    g21202(.A1(new_n21497_), .A2(new_n2168_), .ZN(new_n21500_));
  INV_X1     g21203(.I(new_n21500_), .ZN(new_n21501_));
  NAND2_X1   g21204(.A1(new_n21497_), .A2(new_n2168_), .ZN(new_n21502_));
  AOI21_X1   g21205(.A1(new_n21501_), .A2(new_n21502_), .B(new_n21340_), .ZN(new_n21503_));
  NOR2_X1    g21206(.A1(new_n21499_), .A2(new_n21503_), .ZN(new_n21504_));
  NOR2_X1    g21207(.A1(new_n21493_), .A2(new_n21504_), .ZN(new_n21505_));
  INV_X1     g21208(.I(new_n21505_), .ZN(new_n21506_));
  NAND2_X1   g21209(.A1(new_n21493_), .A2(new_n21504_), .ZN(new_n21507_));
  AOI21_X1   g21210(.A1(new_n21506_), .A2(new_n21507_), .B(new_n21489_), .ZN(new_n21508_));
  XOR2_X1    g21211(.A1(new_n21492_), .A2(new_n21504_), .Z(new_n21509_));
  INV_X1     g21212(.I(new_n21509_), .ZN(new_n21510_));
  AOI21_X1   g21213(.A1(new_n21489_), .A2(new_n21510_), .B(new_n21508_), .ZN(new_n21511_));
  XNOR2_X1   g21214(.A1(new_n21511_), .A2(new_n21487_), .ZN(new_n21512_));
  NOR2_X1    g21215(.A1(new_n21512_), .A2(new_n21484_), .ZN(new_n21513_));
  INV_X1     g21216(.I(new_n21484_), .ZN(new_n21514_));
  NOR2_X1    g21217(.A1(new_n21511_), .A2(new_n21487_), .ZN(new_n21515_));
  INV_X1     g21218(.I(new_n21515_), .ZN(new_n21516_));
  NAND2_X1   g21219(.A1(new_n21511_), .A2(new_n21487_), .ZN(new_n21517_));
  AOI21_X1   g21220(.A1(new_n21516_), .A2(new_n21517_), .B(new_n21514_), .ZN(new_n21518_));
  NOR2_X1    g21221(.A1(new_n21513_), .A2(new_n21518_), .ZN(new_n21519_));
  AOI22_X1   g21222(.A1(new_n10969_), .A2(new_n20981_), .B1(new_n11394_), .B2(\b[34] ), .ZN(new_n21520_));
  OAI21_X1   g21223(.A1(new_n21520_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n21521_));
  XOR2_X1    g21224(.A1(new_n4778_), .A2(new_n21521_), .Z(new_n21522_));
  NAND2_X1   g21225(.A1(new_n21360_), .A2(new_n21356_), .ZN(new_n21523_));
  NAND2_X1   g21226(.A1(new_n21523_), .A2(new_n21359_), .ZN(new_n21524_));
  INV_X1     g21227(.I(new_n21524_), .ZN(new_n21525_));
  NOR2_X1    g21228(.A1(new_n21525_), .A2(new_n21522_), .ZN(new_n21526_));
  INV_X1     g21229(.I(new_n21522_), .ZN(new_n21527_));
  NOR2_X1    g21230(.A1(new_n21524_), .A2(new_n21527_), .ZN(new_n21528_));
  NOR2_X1    g21231(.A1(new_n21526_), .A2(new_n21528_), .ZN(new_n21529_));
  NOR2_X1    g21232(.A1(new_n21529_), .A2(new_n21519_), .ZN(new_n21530_));
  XOR2_X1    g21233(.A1(new_n21524_), .A2(new_n21522_), .Z(new_n21531_));
  NOR3_X1    g21234(.A1(new_n21531_), .A2(new_n21513_), .A3(new_n21518_), .ZN(new_n21532_));
  NOR2_X1    g21235(.A1(new_n21530_), .A2(new_n21532_), .ZN(new_n21533_));
  AOI22_X1   g21236(.A1(new_n11415_), .A2(new_n5915_), .B1(\b[37] ), .B2(new_n10145_), .ZN(new_n21534_));
  OAI21_X1   g21237(.A1(new_n21534_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n21535_));
  XOR2_X1    g21238(.A1(new_n5600_), .A2(new_n21535_), .Z(new_n21536_));
  XOR2_X1    g21239(.A1(new_n21533_), .A2(new_n21536_), .Z(new_n21537_));
  NOR3_X1    g21240(.A1(new_n21530_), .A2(new_n21532_), .A3(new_n21536_), .ZN(new_n21538_));
  INV_X1     g21241(.I(new_n21536_), .ZN(new_n21539_));
  NOR2_X1    g21242(.A1(new_n21533_), .A2(new_n21539_), .ZN(new_n21540_));
  OAI21_X1   g21243(.A1(new_n21540_), .A2(new_n21538_), .B(new_n21483_), .ZN(new_n21541_));
  OAI21_X1   g21244(.A1(new_n21483_), .A2(new_n21537_), .B(new_n21541_), .ZN(new_n21542_));
  OAI22_X1   g21245(.A1(new_n8644_), .A2(new_n6229_), .B1(new_n6538_), .B2(new_n9388_), .ZN(new_n21543_));
  OAI21_X1   g21246(.A1(new_n5921_), .A2(new_n10154_), .B(new_n21543_), .ZN(new_n21544_));
  AOI21_X1   g21247(.A1(new_n21544_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n21545_));
  XOR2_X1    g21248(.A1(new_n6543_), .A2(new_n21545_), .Z(new_n21546_));
  NOR2_X1    g21249(.A1(new_n21542_), .A2(new_n21546_), .ZN(new_n21547_));
  INV_X1     g21250(.I(new_n21547_), .ZN(new_n21548_));
  NAND2_X1   g21251(.A1(new_n21542_), .A2(new_n21546_), .ZN(new_n21549_));
  AOI21_X1   g21252(.A1(new_n21548_), .A2(new_n21549_), .B(new_n21481_), .ZN(new_n21550_));
  XOR2_X1    g21253(.A1(new_n21542_), .A2(new_n21546_), .Z(new_n21551_));
  AOI21_X1   g21254(.A1(new_n21481_), .A2(new_n21551_), .B(new_n21550_), .ZN(new_n21552_));
  OAI22_X1   g21255(.A1(new_n7619_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n8309_), .ZN(new_n21553_));
  OAI21_X1   g21256(.A1(new_n6847_), .A2(new_n7947_), .B(new_n21553_), .ZN(new_n21554_));
  AOI21_X1   g21257(.A1(new_n21554_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n21555_));
  XOR2_X1    g21258(.A1(new_n7516_), .A2(new_n21555_), .Z(new_n21556_));
  XOR2_X1    g21259(.A1(new_n21552_), .A2(new_n21556_), .Z(new_n21557_));
  AND2_X2    g21260(.A1(new_n21557_), .A2(new_n21479_), .Z(new_n21558_));
  NOR2_X1    g21261(.A1(new_n21552_), .A2(new_n21556_), .ZN(new_n21559_));
  INV_X1     g21262(.I(new_n21559_), .ZN(new_n21560_));
  NAND2_X1   g21263(.A1(new_n21552_), .A2(new_n21556_), .ZN(new_n21561_));
  AOI21_X1   g21264(.A1(new_n21560_), .A2(new_n21561_), .B(new_n21479_), .ZN(new_n21562_));
  NOR2_X1    g21265(.A1(new_n21558_), .A2(new_n21562_), .ZN(new_n21563_));
  OAI22_X1   g21266(.A1(new_n6644_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n6647_), .ZN(new_n21564_));
  OAI21_X1   g21267(.A1(new_n7870_), .A2(new_n7284_), .B(new_n21564_), .ZN(new_n21565_));
  AOI21_X1   g21268(.A1(new_n21565_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n21566_));
  XNOR2_X1   g21269(.A1(new_n8568_), .A2(new_n21566_), .ZN(new_n21567_));
  INV_X1     g21270(.I(new_n21399_), .ZN(new_n21568_));
  OAI21_X1   g21271(.A1(new_n21390_), .A2(new_n21568_), .B(new_n21398_), .ZN(new_n21569_));
  NAND2_X1   g21272(.A1(new_n21569_), .A2(new_n21567_), .ZN(new_n21570_));
  NOR2_X1    g21273(.A1(new_n21569_), .A2(new_n21567_), .ZN(new_n21571_));
  INV_X1     g21274(.I(new_n21571_), .ZN(new_n21572_));
  AOI21_X1   g21275(.A1(new_n21572_), .A2(new_n21570_), .B(new_n21563_), .ZN(new_n21573_));
  XNOR2_X1   g21276(.A1(new_n21569_), .A2(new_n21567_), .ZN(new_n21574_));
  NOR3_X1    g21277(.A1(new_n21558_), .A2(new_n21562_), .A3(new_n21574_), .ZN(new_n21575_));
  OAI22_X1   g21278(.A1(new_n5993_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n5991_), .ZN(new_n21576_));
  OAI21_X1   g21279(.A1(new_n8948_), .A2(new_n5997_), .B(new_n21576_), .ZN(new_n21577_));
  AOI21_X1   g21280(.A1(new_n21577_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n21578_));
  XNOR2_X1   g21281(.A1(new_n9642_), .A2(new_n21578_), .ZN(new_n21579_));
  NOR3_X1    g21282(.A1(new_n21573_), .A2(new_n21575_), .A3(new_n21579_), .ZN(new_n21580_));
  NOR2_X1    g21283(.A1(new_n21573_), .A2(new_n21575_), .ZN(new_n21581_));
  INV_X1     g21284(.I(new_n21579_), .ZN(new_n21582_));
  NOR2_X1    g21285(.A1(new_n21581_), .A2(new_n21582_), .ZN(new_n21583_));
  OAI21_X1   g21286(.A1(new_n21583_), .A2(new_n21580_), .B(new_n21477_), .ZN(new_n21584_));
  XOR2_X1    g21287(.A1(new_n21581_), .A2(new_n21582_), .Z(new_n21585_));
  NAND2_X1   g21288(.A1(new_n21585_), .A2(new_n21476_), .ZN(new_n21586_));
  NAND2_X1   g21289(.A1(new_n21586_), .A2(new_n21584_), .ZN(new_n21587_));
  OAI22_X1   g21290(.A1(new_n5420_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n5107_), .ZN(new_n21588_));
  OAI21_X1   g21291(.A1(new_n10031_), .A2(new_n5112_), .B(new_n21588_), .ZN(new_n21589_));
  AOI21_X1   g21292(.A1(new_n21589_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n21590_));
  XNOR2_X1   g21293(.A1(new_n10866_), .A2(new_n21590_), .ZN(new_n21591_));
  XOR2_X1    g21294(.A1(new_n21587_), .A2(new_n21591_), .Z(new_n21592_));
  NOR2_X1    g21295(.A1(new_n21592_), .A2(new_n21475_), .ZN(new_n21593_));
  INV_X1     g21296(.I(new_n21475_), .ZN(new_n21594_));
  INV_X1     g21297(.I(new_n21587_), .ZN(new_n21595_));
  NOR2_X1    g21298(.A1(new_n21595_), .A2(new_n21591_), .ZN(new_n21596_));
  INV_X1     g21299(.I(new_n21596_), .ZN(new_n21597_));
  NAND2_X1   g21300(.A1(new_n21595_), .A2(new_n21591_), .ZN(new_n21598_));
  AOI21_X1   g21301(.A1(new_n21597_), .A2(new_n21598_), .B(new_n21594_), .ZN(new_n21599_));
  NOR2_X1    g21302(.A1(new_n21599_), .A2(new_n21593_), .ZN(new_n21600_));
  OAI22_X1   g21303(.A1(new_n4072_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n4067_), .ZN(new_n21601_));
  OAI21_X1   g21304(.A1(new_n11738_), .A2(new_n4318_), .B(new_n21601_), .ZN(new_n21602_));
  AOI21_X1   g21305(.A1(new_n21602_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n21603_));
  XNOR2_X1   g21306(.A1(new_n12128_), .A2(new_n21603_), .ZN(new_n21604_));
  XOR2_X1    g21307(.A1(new_n21600_), .A2(new_n21604_), .Z(new_n21605_));
  INV_X1     g21308(.I(new_n21605_), .ZN(new_n21606_));
  INV_X1     g21309(.I(new_n21600_), .ZN(new_n21607_));
  NOR2_X1    g21310(.A1(new_n21607_), .A2(new_n21604_), .ZN(new_n21608_));
  INV_X1     g21311(.I(new_n21608_), .ZN(new_n21609_));
  NAND2_X1   g21312(.A1(new_n21607_), .A2(new_n21604_), .ZN(new_n21610_));
  AOI21_X1   g21313(.A1(new_n21609_), .A2(new_n21610_), .B(new_n21474_), .ZN(new_n21611_));
  AOI21_X1   g21314(.A1(new_n21474_), .A2(new_n21606_), .B(new_n21611_), .ZN(new_n21612_));
  OAI22_X1   g21315(.A1(new_n12970_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n13367_), .ZN(new_n21613_));
  OAI21_X1   g21316(.A1(new_n12542_), .A2(new_n3569_), .B(new_n21613_), .ZN(new_n21614_));
  AOI21_X1   g21317(.A1(new_n21614_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n21615_));
  XNOR2_X1   g21318(.A1(new_n13371_), .A2(new_n21615_), .ZN(new_n21616_));
  INV_X1     g21319(.I(new_n21433_), .ZN(new_n21617_));
  OAI21_X1   g21320(.A1(new_n21435_), .A2(new_n21434_), .B(new_n21298_), .ZN(new_n21618_));
  NAND2_X1   g21321(.A1(new_n21618_), .A2(new_n21617_), .ZN(new_n21619_));
  XOR2_X1    g21322(.A1(new_n21619_), .A2(new_n21616_), .Z(new_n21620_));
  NOR2_X1    g21323(.A1(new_n21620_), .A2(new_n21612_), .ZN(new_n21621_));
  INV_X1     g21324(.I(new_n21619_), .ZN(new_n21622_));
  NOR2_X1    g21325(.A1(new_n21622_), .A2(new_n21616_), .ZN(new_n21623_));
  INV_X1     g21326(.I(new_n21623_), .ZN(new_n21624_));
  NAND2_X1   g21327(.A1(new_n21622_), .A2(new_n21616_), .ZN(new_n21625_));
  NAND2_X1   g21328(.A1(new_n21624_), .A2(new_n21625_), .ZN(new_n21626_));
  AOI21_X1   g21329(.A1(new_n21612_), .A2(new_n21626_), .B(new_n21621_), .ZN(new_n21627_));
  XNOR2_X1   g21330(.A1(new_n21627_), .A2(new_n21471_), .ZN(new_n21628_));
  NOR2_X1    g21331(.A1(new_n21628_), .A2(new_n21467_), .ZN(new_n21629_));
  INV_X1     g21332(.I(new_n21467_), .ZN(new_n21630_));
  NOR2_X1    g21333(.A1(new_n21627_), .A2(new_n21471_), .ZN(new_n21631_));
  INV_X1     g21334(.I(new_n21631_), .ZN(new_n21632_));
  NAND2_X1   g21335(.A1(new_n21627_), .A2(new_n21471_), .ZN(new_n21633_));
  AOI21_X1   g21336(.A1(new_n21632_), .A2(new_n21633_), .B(new_n21630_), .ZN(new_n21634_));
  NOR2_X1    g21337(.A1(new_n21629_), .A2(new_n21634_), .ZN(new_n21635_));
  XNOR2_X1   g21338(.A1(new_n21465_), .A2(new_n21635_), .ZN(new_n21636_));
  INV_X1     g21339(.I(new_n21636_), .ZN(new_n21637_));
  NAND2_X1   g21340(.A1(new_n21459_), .A2(new_n21637_), .ZN(new_n21638_));
  XOR2_X1    g21341(.A1(new_n21638_), .A2(new_n21456_), .Z(new_n21639_));
  XOR2_X1    g21342(.A1(new_n21285_), .A2(new_n21639_), .Z(\f[90] ));
  NOR2_X1    g21343(.A1(new_n21465_), .A2(new_n21635_), .ZN(new_n21641_));
  NAND3_X1   g21344(.A1(new_n20718_), .A2(new_n21096_), .A3(new_n21283_), .ZN(new_n21642_));
  NOR2_X1    g21345(.A1(new_n21455_), .A2(new_n21637_), .ZN(new_n21643_));
  AOI21_X1   g21346(.A1(new_n21455_), .A2(new_n21637_), .B(new_n21287_), .ZN(new_n21644_));
  NOR2_X1    g21347(.A1(new_n21644_), .A2(new_n21643_), .ZN(new_n21645_));
  INV_X1     g21348(.I(new_n21645_), .ZN(new_n21646_));
  AOI21_X1   g21349(.A1(new_n21642_), .A2(new_n21282_), .B(new_n21646_), .ZN(new_n21647_));
  NOR2_X1    g21350(.A1(new_n2884_), .A2(new_n2700_), .ZN(new_n21648_));
  NAND2_X1   g21351(.A1(new_n16148_), .A2(new_n2702_), .ZN(new_n21649_));
  OAI21_X1   g21352(.A1(new_n21648_), .A2(new_n21649_), .B(new_n2694_), .ZN(new_n21650_));
  XNOR2_X1   g21353(.A1(new_n14978_), .A2(new_n21650_), .ZN(new_n21651_));
  AOI21_X1   g21354(.A1(new_n21612_), .A2(new_n21625_), .B(new_n21623_), .ZN(new_n21652_));
  INV_X1     g21355(.I(new_n21652_), .ZN(new_n21653_));
  OAI22_X1   g21356(.A1(new_n13367_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n13785_), .ZN(new_n21654_));
  OAI21_X1   g21357(.A1(new_n12970_), .A2(new_n3569_), .B(new_n21654_), .ZN(new_n21655_));
  AOI21_X1   g21358(.A1(new_n21655_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n21656_));
  XOR2_X1    g21359(.A1(new_n13784_), .A2(new_n21656_), .Z(new_n21657_));
  AOI21_X1   g21360(.A1(new_n21474_), .A2(new_n21610_), .B(new_n21608_), .ZN(new_n21658_));
  OAI22_X1   g21361(.A1(new_n4072_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n4067_), .ZN(new_n21659_));
  OAI21_X1   g21362(.A1(new_n11744_), .A2(new_n4318_), .B(new_n21659_), .ZN(new_n21660_));
  AOI21_X1   g21363(.A1(new_n21660_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n21661_));
  XNOR2_X1   g21364(.A1(new_n12546_), .A2(new_n21661_), .ZN(new_n21662_));
  AOI21_X1   g21365(.A1(new_n21594_), .A2(new_n21598_), .B(new_n21596_), .ZN(new_n21663_));
  INV_X1     g21366(.I(new_n21663_), .ZN(new_n21664_));
  NOR2_X1    g21367(.A1(new_n21583_), .A2(new_n21476_), .ZN(new_n21665_));
  NOR2_X1    g21368(.A1(new_n21665_), .A2(new_n21580_), .ZN(new_n21666_));
  OAI22_X1   g21369(.A1(new_n5993_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n5991_), .ZN(new_n21667_));
  OAI21_X1   g21370(.A1(new_n9295_), .A2(new_n5997_), .B(new_n21667_), .ZN(new_n21668_));
  AOI21_X1   g21371(.A1(new_n21668_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n21669_));
  XNOR2_X1   g21372(.A1(new_n10035_), .A2(new_n21669_), .ZN(new_n21670_));
  INV_X1     g21373(.I(new_n21670_), .ZN(new_n21671_));
  OAI22_X1   g21374(.A1(new_n7619_), .A2(new_n7864_), .B1(new_n7870_), .B2(new_n8309_), .ZN(new_n21672_));
  OAI21_X1   g21375(.A1(new_n7198_), .A2(new_n7947_), .B(new_n21672_), .ZN(new_n21673_));
  AOI21_X1   g21376(.A1(new_n21673_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n21674_));
  XNOR2_X1   g21377(.A1(new_n7874_), .A2(new_n21674_), .ZN(new_n21675_));
  NOR2_X1    g21378(.A1(new_n21540_), .A2(new_n21483_), .ZN(new_n21676_));
  NOR2_X1    g21379(.A1(new_n21676_), .A2(new_n21538_), .ZN(new_n21677_));
  AOI22_X1   g21380(.A1(new_n11415_), .A2(new_n5923_), .B1(\b[38] ), .B2(new_n10145_), .ZN(new_n21678_));
  OAI21_X1   g21381(.A1(new_n21678_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n21679_));
  XNOR2_X1   g21382(.A1(new_n5926_), .A2(new_n21679_), .ZN(new_n21680_));
  INV_X1     g21383(.I(new_n21528_), .ZN(new_n21681_));
  AOI21_X1   g21384(.A1(new_n21519_), .A2(new_n21681_), .B(new_n21526_), .ZN(new_n21682_));
  AOI22_X1   g21385(.A1(new_n13078_), .A2(\b[32] ), .B1(new_n20556_), .B2(new_n12218_), .ZN(new_n21683_));
  OAI21_X1   g21386(.A1(new_n21683_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n21684_));
  XOR2_X1    g21387(.A1(new_n4257_), .A2(new_n21684_), .Z(new_n21685_));
  OAI22_X1   g21388(.A1(new_n13880_), .A2(new_n3710_), .B1(new_n3018_), .B2(new_n13885_), .ZN(new_n21686_));
  AOI21_X1   g21389(.A1(new_n21686_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n21687_));
  XNOR2_X1   g21390(.A1(new_n3514_), .A2(new_n21687_), .ZN(new_n21688_));
  NAND2_X1   g21391(.A1(new_n21502_), .A2(new_n21340_), .ZN(new_n21689_));
  NAND2_X1   g21392(.A1(new_n21689_), .A2(new_n21501_), .ZN(new_n21690_));
  NOR2_X1    g21393(.A1(new_n13476_), .A2(new_n2643_), .ZN(new_n21691_));
  XOR2_X1    g21394(.A1(new_n14736_), .A2(new_n2643_), .Z(new_n21692_));
  NAND2_X1   g21395(.A1(new_n21692_), .A2(\b[28] ), .ZN(new_n21693_));
  XOR2_X1    g21396(.A1(new_n21693_), .A2(new_n21691_), .Z(new_n21694_));
  INV_X1     g21397(.I(new_n21694_), .ZN(new_n21695_));
  XOR2_X1    g21398(.A1(new_n21690_), .A2(new_n21695_), .Z(new_n21696_));
  NOR2_X1    g21399(.A1(new_n21688_), .A2(new_n21696_), .ZN(new_n21697_));
  INV_X1     g21400(.I(new_n21688_), .ZN(new_n21698_));
  NOR2_X1    g21401(.A1(new_n21690_), .A2(new_n21694_), .ZN(new_n21699_));
  INV_X1     g21402(.I(new_n21699_), .ZN(new_n21700_));
  NAND2_X1   g21403(.A1(new_n21690_), .A2(new_n21694_), .ZN(new_n21701_));
  AOI21_X1   g21404(.A1(new_n21700_), .A2(new_n21701_), .B(new_n21698_), .ZN(new_n21702_));
  NOR2_X1    g21405(.A1(new_n21702_), .A2(new_n21697_), .ZN(new_n21703_));
  OAI21_X1   g21406(.A1(new_n21489_), .A2(new_n21505_), .B(new_n21507_), .ZN(new_n21704_));
  AND2_X2    g21407(.A1(new_n21704_), .A2(new_n21703_), .Z(new_n21705_));
  NOR2_X1    g21408(.A1(new_n21704_), .A2(new_n21703_), .ZN(new_n21706_));
  NOR2_X1    g21409(.A1(new_n21705_), .A2(new_n21706_), .ZN(new_n21707_));
  NOR2_X1    g21410(.A1(new_n21707_), .A2(new_n21685_), .ZN(new_n21708_));
  XOR2_X1    g21411(.A1(new_n21704_), .A2(new_n21703_), .Z(new_n21709_));
  AOI21_X1   g21412(.A1(new_n21685_), .A2(new_n21709_), .B(new_n21708_), .ZN(new_n21710_));
  NAND2_X1   g21413(.A1(new_n21517_), .A2(new_n21514_), .ZN(new_n21711_));
  NAND2_X1   g21414(.A1(new_n21711_), .A2(new_n21516_), .ZN(new_n21712_));
  INV_X1     g21415(.I(new_n21712_), .ZN(new_n21713_));
  AOI22_X1   g21416(.A1(new_n10969_), .A2(new_n5349_), .B1(new_n11394_), .B2(\b[35] ), .ZN(new_n21714_));
  OAI21_X1   g21417(.A1(new_n21714_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n21715_));
  XNOR2_X1   g21418(.A1(new_n5067_), .A2(new_n21715_), .ZN(new_n21716_));
  NOR2_X1    g21419(.A1(new_n21713_), .A2(new_n21716_), .ZN(new_n21717_));
  INV_X1     g21420(.I(new_n21716_), .ZN(new_n21718_));
  NOR2_X1    g21421(.A1(new_n21712_), .A2(new_n21718_), .ZN(new_n21719_));
  NOR2_X1    g21422(.A1(new_n21717_), .A2(new_n21719_), .ZN(new_n21720_));
  NOR2_X1    g21423(.A1(new_n21720_), .A2(new_n21710_), .ZN(new_n21721_));
  INV_X1     g21424(.I(new_n21710_), .ZN(new_n21722_));
  XOR2_X1    g21425(.A1(new_n21712_), .A2(new_n21716_), .Z(new_n21723_));
  NOR2_X1    g21426(.A1(new_n21723_), .A2(new_n21722_), .ZN(new_n21724_));
  NOR2_X1    g21427(.A1(new_n21721_), .A2(new_n21724_), .ZN(new_n21725_));
  XNOR2_X1   g21428(.A1(new_n21682_), .A2(new_n21725_), .ZN(new_n21726_));
  NOR2_X1    g21429(.A1(new_n21682_), .A2(new_n21725_), .ZN(new_n21727_));
  NAND2_X1   g21430(.A1(new_n21682_), .A2(new_n21725_), .ZN(new_n21728_));
  INV_X1     g21431(.I(new_n21728_), .ZN(new_n21729_));
  OAI21_X1   g21432(.A1(new_n21729_), .A2(new_n21727_), .B(new_n21680_), .ZN(new_n21730_));
  OAI21_X1   g21433(.A1(new_n21680_), .A2(new_n21726_), .B(new_n21730_), .ZN(new_n21731_));
  AOI22_X1   g21434(.A1(new_n8631_), .A2(\b[42] ), .B1(\b[43] ), .B2(new_n9382_), .ZN(new_n21732_));
  AOI21_X1   g21435(.A1(\b[41] ), .A2(new_n9731_), .B(new_n21732_), .ZN(new_n21733_));
  OAI21_X1   g21436(.A1(new_n21733_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n21734_));
  XNOR2_X1   g21437(.A1(new_n6851_), .A2(new_n21734_), .ZN(new_n21735_));
  NOR2_X1    g21438(.A1(new_n21731_), .A2(new_n21735_), .ZN(new_n21736_));
  INV_X1     g21439(.I(new_n21736_), .ZN(new_n21737_));
  NAND2_X1   g21440(.A1(new_n21731_), .A2(new_n21735_), .ZN(new_n21738_));
  AOI21_X1   g21441(.A1(new_n21737_), .A2(new_n21738_), .B(new_n21677_), .ZN(new_n21739_));
  INV_X1     g21442(.I(new_n21677_), .ZN(new_n21740_));
  XNOR2_X1   g21443(.A1(new_n21731_), .A2(new_n21735_), .ZN(new_n21741_));
  NOR2_X1    g21444(.A1(new_n21741_), .A2(new_n21740_), .ZN(new_n21742_));
  NOR2_X1    g21445(.A1(new_n21742_), .A2(new_n21739_), .ZN(new_n21743_));
  INV_X1     g21446(.I(new_n21481_), .ZN(new_n21744_));
  AOI21_X1   g21447(.A1(new_n21744_), .A2(new_n21549_), .B(new_n21547_), .ZN(new_n21745_));
  NOR2_X1    g21448(.A1(new_n21743_), .A2(new_n21745_), .ZN(new_n21746_));
  INV_X1     g21449(.I(new_n21746_), .ZN(new_n21747_));
  NAND2_X1   g21450(.A1(new_n21743_), .A2(new_n21745_), .ZN(new_n21748_));
  AOI21_X1   g21451(.A1(new_n21747_), .A2(new_n21748_), .B(new_n21675_), .ZN(new_n21749_));
  INV_X1     g21452(.I(new_n21675_), .ZN(new_n21750_));
  XNOR2_X1   g21453(.A1(new_n21743_), .A2(new_n21745_), .ZN(new_n21751_));
  NOR2_X1    g21454(.A1(new_n21751_), .A2(new_n21750_), .ZN(new_n21752_));
  NOR2_X1    g21455(.A1(new_n21752_), .A2(new_n21749_), .ZN(new_n21753_));
  NAND2_X1   g21456(.A1(new_n21561_), .A2(new_n21479_), .ZN(new_n21754_));
  NAND2_X1   g21457(.A1(new_n21754_), .A2(new_n21560_), .ZN(new_n21755_));
  INV_X1     g21458(.I(new_n21755_), .ZN(new_n21756_));
  OAI22_X1   g21459(.A1(new_n6644_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n6647_), .ZN(new_n21757_));
  OAI21_X1   g21460(.A1(new_n8218_), .A2(new_n7284_), .B(new_n21757_), .ZN(new_n21758_));
  AOI21_X1   g21461(.A1(new_n21758_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n21759_));
  XOR2_X1    g21462(.A1(new_n8952_), .A2(new_n21759_), .Z(new_n21760_));
  NOR2_X1    g21463(.A1(new_n21756_), .A2(new_n21760_), .ZN(new_n21761_));
  INV_X1     g21464(.I(new_n21760_), .ZN(new_n21762_));
  NOR2_X1    g21465(.A1(new_n21755_), .A2(new_n21762_), .ZN(new_n21763_));
  NOR2_X1    g21466(.A1(new_n21761_), .A2(new_n21763_), .ZN(new_n21764_));
  NOR2_X1    g21467(.A1(new_n21764_), .A2(new_n21753_), .ZN(new_n21765_));
  INV_X1     g21468(.I(new_n21753_), .ZN(new_n21766_));
  XOR2_X1    g21469(.A1(new_n21755_), .A2(new_n21760_), .Z(new_n21767_));
  NOR2_X1    g21470(.A1(new_n21767_), .A2(new_n21766_), .ZN(new_n21768_));
  NOR2_X1    g21471(.A1(new_n21765_), .A2(new_n21768_), .ZN(new_n21769_));
  NAND2_X1   g21472(.A1(new_n21563_), .A2(new_n21572_), .ZN(new_n21770_));
  AOI21_X1   g21473(.A1(new_n21570_), .A2(new_n21770_), .B(new_n21769_), .ZN(new_n21771_));
  NAND2_X1   g21474(.A1(new_n21770_), .A2(new_n21570_), .ZN(new_n21772_));
  NOR3_X1    g21475(.A1(new_n21772_), .A2(new_n21765_), .A3(new_n21768_), .ZN(new_n21773_));
  OAI21_X1   g21476(.A1(new_n21771_), .A2(new_n21773_), .B(new_n21671_), .ZN(new_n21774_));
  XNOR2_X1   g21477(.A1(new_n21769_), .A2(new_n21772_), .ZN(new_n21775_));
  NAND2_X1   g21478(.A1(new_n21775_), .A2(new_n21670_), .ZN(new_n21776_));
  NAND2_X1   g21479(.A1(new_n21776_), .A2(new_n21774_), .ZN(new_n21777_));
  OAI22_X1   g21480(.A1(new_n5420_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n5107_), .ZN(new_n21778_));
  OAI21_X1   g21481(.A1(new_n10477_), .A2(new_n5112_), .B(new_n21778_), .ZN(new_n21779_));
  AOI21_X1   g21482(.A1(new_n21779_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n21780_));
  XOR2_X1    g21483(.A1(new_n11298_), .A2(new_n21780_), .Z(new_n21781_));
  XOR2_X1    g21484(.A1(new_n21777_), .A2(new_n21781_), .Z(new_n21782_));
  NOR2_X1    g21485(.A1(new_n21782_), .A2(new_n21666_), .ZN(new_n21783_));
  INV_X1     g21486(.I(new_n21666_), .ZN(new_n21784_));
  INV_X1     g21487(.I(new_n21777_), .ZN(new_n21785_));
  NOR2_X1    g21488(.A1(new_n21785_), .A2(new_n21781_), .ZN(new_n21786_));
  INV_X1     g21489(.I(new_n21786_), .ZN(new_n21787_));
  NAND2_X1   g21490(.A1(new_n21785_), .A2(new_n21781_), .ZN(new_n21788_));
  AOI21_X1   g21491(.A1(new_n21787_), .A2(new_n21788_), .B(new_n21784_), .ZN(new_n21789_));
  NOR2_X1    g21492(.A1(new_n21789_), .A2(new_n21783_), .ZN(new_n21790_));
  NOR2_X1    g21493(.A1(new_n21790_), .A2(new_n21664_), .ZN(new_n21791_));
  INV_X1     g21494(.I(new_n21790_), .ZN(new_n21792_));
  NOR2_X1    g21495(.A1(new_n21792_), .A2(new_n21663_), .ZN(new_n21793_));
  NOR2_X1    g21496(.A1(new_n21793_), .A2(new_n21791_), .ZN(new_n21794_));
  NOR2_X1    g21497(.A1(new_n21794_), .A2(new_n21662_), .ZN(new_n21795_));
  INV_X1     g21498(.I(new_n21662_), .ZN(new_n21796_));
  XOR2_X1    g21499(.A1(new_n21790_), .A2(new_n21663_), .Z(new_n21797_));
  NOR2_X1    g21500(.A1(new_n21797_), .A2(new_n21796_), .ZN(new_n21798_));
  NOR2_X1    g21501(.A1(new_n21795_), .A2(new_n21798_), .ZN(new_n21799_));
  XNOR2_X1   g21502(.A1(new_n21799_), .A2(new_n21658_), .ZN(new_n21800_));
  NOR2_X1    g21503(.A1(new_n21800_), .A2(new_n21657_), .ZN(new_n21801_));
  INV_X1     g21504(.I(new_n21657_), .ZN(new_n21802_));
  NOR2_X1    g21505(.A1(new_n21799_), .A2(new_n21658_), .ZN(new_n21803_));
  INV_X1     g21506(.I(new_n21803_), .ZN(new_n21804_));
  NAND2_X1   g21507(.A1(new_n21799_), .A2(new_n21658_), .ZN(new_n21805_));
  AOI21_X1   g21508(.A1(new_n21804_), .A2(new_n21805_), .B(new_n21802_), .ZN(new_n21806_));
  NOR2_X1    g21509(.A1(new_n21801_), .A2(new_n21806_), .ZN(new_n21807_));
  NOR2_X1    g21510(.A1(new_n21807_), .A2(new_n21653_), .ZN(new_n21808_));
  INV_X1     g21511(.I(new_n21807_), .ZN(new_n21809_));
  NOR2_X1    g21512(.A1(new_n21809_), .A2(new_n21652_), .ZN(new_n21810_));
  NOR2_X1    g21513(.A1(new_n21810_), .A2(new_n21808_), .ZN(new_n21811_));
  NOR2_X1    g21514(.A1(new_n21811_), .A2(new_n21651_), .ZN(new_n21812_));
  INV_X1     g21515(.I(new_n21651_), .ZN(new_n21813_));
  XOR2_X1    g21516(.A1(new_n21807_), .A2(new_n21652_), .Z(new_n21814_));
  NOR2_X1    g21517(.A1(new_n21814_), .A2(new_n21813_), .ZN(new_n21815_));
  NOR2_X1    g21518(.A1(new_n21812_), .A2(new_n21815_), .ZN(new_n21816_));
  AOI21_X1   g21519(.A1(new_n21630_), .A2(new_n21633_), .B(new_n21631_), .ZN(new_n21817_));
  NOR2_X1    g21520(.A1(new_n21816_), .A2(new_n21817_), .ZN(new_n21818_));
  XOR2_X1    g21521(.A1(new_n21647_), .A2(new_n21818_), .Z(new_n21819_));
  XOR2_X1    g21522(.A1(new_n21819_), .A2(new_n21641_), .Z(\f[91] ));
  INV_X1     g21523(.I(new_n21641_), .ZN(new_n21821_));
  NOR2_X1    g21524(.A1(new_n21821_), .A2(new_n21816_), .ZN(new_n21822_));
  INV_X1     g21525(.I(new_n21822_), .ZN(new_n21823_));
  AOI21_X1   g21526(.A1(new_n21821_), .A2(new_n21816_), .B(new_n21817_), .ZN(new_n21824_));
  NAND3_X1   g21527(.A1(new_n21285_), .A2(new_n21645_), .A3(new_n21824_), .ZN(new_n21825_));
  NAND2_X1   g21528(.A1(new_n21825_), .A2(new_n21823_), .ZN(new_n21826_));
  NOR2_X1    g21529(.A1(new_n21808_), .A2(new_n21651_), .ZN(new_n21827_));
  NOR2_X1    g21530(.A1(new_n21827_), .A2(new_n21810_), .ZN(new_n21828_));
  INV_X1     g21531(.I(new_n21828_), .ZN(new_n21829_));
  OAI22_X1   g21532(.A1(new_n13785_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n14208_), .ZN(new_n21830_));
  OAI21_X1   g21533(.A1(new_n13367_), .A2(new_n3569_), .B(new_n21830_), .ZN(new_n21831_));
  AOI21_X1   g21534(.A1(new_n21831_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n21832_));
  XOR2_X1    g21535(.A1(new_n14213_), .A2(new_n21832_), .Z(new_n21833_));
  NOR2_X1    g21536(.A1(new_n21791_), .A2(new_n21662_), .ZN(new_n21834_));
  NOR2_X1    g21537(.A1(new_n21834_), .A2(new_n21793_), .ZN(new_n21835_));
  OAI22_X1   g21538(.A1(new_n5420_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n5107_), .ZN(new_n21836_));
  OAI21_X1   g21539(.A1(new_n10862_), .A2(new_n5112_), .B(new_n21836_), .ZN(new_n21837_));
  AOI21_X1   g21540(.A1(new_n21837_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n21838_));
  XNOR2_X1   g21541(.A1(new_n11748_), .A2(new_n21838_), .ZN(new_n21839_));
  NOR2_X1    g21542(.A1(new_n21773_), .A2(new_n21670_), .ZN(new_n21840_));
  NOR2_X1    g21543(.A1(new_n21840_), .A2(new_n21771_), .ZN(new_n21841_));
  OAI22_X1   g21544(.A1(new_n5993_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n5991_), .ZN(new_n21842_));
  OAI21_X1   g21545(.A1(new_n10025_), .A2(new_n5997_), .B(new_n21842_), .ZN(new_n21843_));
  AOI21_X1   g21546(.A1(new_n21843_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n21844_));
  XOR2_X1    g21547(.A1(new_n10476_), .A2(new_n21844_), .Z(new_n21845_));
  OAI22_X1   g21548(.A1(new_n6644_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n6647_), .ZN(new_n21846_));
  OAI21_X1   g21549(.A1(new_n8563_), .A2(new_n7284_), .B(new_n21846_), .ZN(new_n21847_));
  AOI21_X1   g21550(.A1(new_n21847_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n21848_));
  XNOR2_X1   g21551(.A1(new_n9299_), .A2(new_n21848_), .ZN(new_n21849_));
  AOI22_X1   g21552(.A1(new_n8631_), .A2(\b[43] ), .B1(\b[44] ), .B2(new_n9382_), .ZN(new_n21850_));
  AOI21_X1   g21553(.A1(\b[42] ), .A2(new_n9731_), .B(new_n21850_), .ZN(new_n21851_));
  OAI21_X1   g21554(.A1(new_n21851_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n21852_));
  XOR2_X1    g21555(.A1(new_n7202_), .A2(new_n21852_), .Z(new_n21853_));
  NOR2_X1    g21556(.A1(new_n21729_), .A2(new_n21680_), .ZN(new_n21854_));
  NOR2_X1    g21557(.A1(new_n21854_), .A2(new_n21727_), .ZN(new_n21855_));
  AOI22_X1   g21558(.A1(new_n10969_), .A2(new_n21317_), .B1(new_n11394_), .B2(\b[36] ), .ZN(new_n21856_));
  OAI21_X1   g21559(.A1(new_n21856_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n21857_));
  XOR2_X1    g21560(.A1(new_n5357_), .A2(new_n21857_), .Z(new_n21858_));
  INV_X1     g21561(.I(new_n21858_), .ZN(new_n21859_));
  INV_X1     g21562(.I(new_n21705_), .ZN(new_n21860_));
  OAI21_X1   g21563(.A1(new_n21685_), .A2(new_n21706_), .B(new_n21860_), .ZN(new_n21861_));
  AOI22_X1   g21564(.A1(new_n13078_), .A2(\b[33] ), .B1(new_n4770_), .B2(new_n12218_), .ZN(new_n21862_));
  OAI21_X1   g21565(.A1(new_n21862_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n21863_));
  XNOR2_X1   g21566(.A1(new_n4499_), .A2(new_n21863_), .ZN(new_n21864_));
  OAI21_X1   g21567(.A1(new_n21688_), .A2(new_n21699_), .B(new_n21701_), .ZN(new_n21865_));
  NOR2_X1    g21568(.A1(new_n13476_), .A2(new_n2842_), .ZN(new_n21866_));
  XOR2_X1    g21569(.A1(new_n14736_), .A2(new_n2842_), .Z(new_n21867_));
  NAND2_X1   g21570(.A1(new_n21867_), .A2(\b[29] ), .ZN(new_n21868_));
  XOR2_X1    g21571(.A1(new_n21868_), .A2(new_n21866_), .Z(new_n21869_));
  NOR2_X1    g21572(.A1(new_n21695_), .A2(new_n21869_), .ZN(new_n21870_));
  INV_X1     g21573(.I(new_n21870_), .ZN(new_n21871_));
  INV_X1     g21574(.I(new_n21869_), .ZN(new_n21872_));
  NOR2_X1    g21575(.A1(new_n21872_), .A2(new_n21694_), .ZN(new_n21873_));
  INV_X1     g21576(.I(new_n21873_), .ZN(new_n21874_));
  NAND2_X1   g21577(.A1(new_n21871_), .A2(new_n21874_), .ZN(new_n21875_));
  XOR2_X1    g21578(.A1(new_n21694_), .A2(new_n21869_), .Z(new_n21876_));
  NOR2_X1    g21579(.A1(new_n21865_), .A2(new_n21876_), .ZN(new_n21877_));
  AOI21_X1   g21580(.A1(new_n21865_), .A2(new_n21875_), .B(new_n21877_), .ZN(new_n21878_));
  OAI22_X1   g21581(.A1(new_n13880_), .A2(new_n3718_), .B1(new_n3260_), .B2(new_n13885_), .ZN(new_n21879_));
  AOI21_X1   g21582(.A1(new_n21879_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n21880_));
  XOR2_X1    g21583(.A1(new_n3722_), .A2(new_n21880_), .Z(new_n21881_));
  XNOR2_X1   g21584(.A1(new_n21878_), .A2(new_n21881_), .ZN(new_n21882_));
  NOR2_X1    g21585(.A1(new_n21882_), .A2(new_n21864_), .ZN(new_n21883_));
  INV_X1     g21586(.I(new_n21864_), .ZN(new_n21884_));
  NOR2_X1    g21587(.A1(new_n21878_), .A2(new_n21881_), .ZN(new_n21885_));
  INV_X1     g21588(.I(new_n21885_), .ZN(new_n21886_));
  NAND2_X1   g21589(.A1(new_n21878_), .A2(new_n21881_), .ZN(new_n21887_));
  AOI21_X1   g21590(.A1(new_n21886_), .A2(new_n21887_), .B(new_n21884_), .ZN(new_n21888_));
  NOR2_X1    g21591(.A1(new_n21883_), .A2(new_n21888_), .ZN(new_n21889_));
  NOR2_X1    g21592(.A1(new_n21889_), .A2(new_n21861_), .ZN(new_n21890_));
  AND2_X2    g21593(.A1(new_n21889_), .A2(new_n21861_), .Z(new_n21891_));
  OAI21_X1   g21594(.A1(new_n21891_), .A2(new_n21890_), .B(new_n21859_), .ZN(new_n21892_));
  XOR2_X1    g21595(.A1(new_n21889_), .A2(new_n21861_), .Z(new_n21893_));
  NAND2_X1   g21596(.A1(new_n21893_), .A2(new_n21858_), .ZN(new_n21894_));
  NAND2_X1   g21597(.A1(new_n21894_), .A2(new_n21892_), .ZN(new_n21895_));
  AOI22_X1   g21598(.A1(new_n11415_), .A2(new_n6532_), .B1(\b[39] ), .B2(new_n10145_), .ZN(new_n21896_));
  OAI21_X1   g21599(.A1(new_n21896_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n21897_));
  XNOR2_X1   g21600(.A1(new_n6233_), .A2(new_n21897_), .ZN(new_n21898_));
  NOR2_X1    g21601(.A1(new_n21719_), .A2(new_n21710_), .ZN(new_n21899_));
  NOR2_X1    g21602(.A1(new_n21899_), .A2(new_n21717_), .ZN(new_n21900_));
  NOR2_X1    g21603(.A1(new_n21900_), .A2(new_n21898_), .ZN(new_n21901_));
  INV_X1     g21604(.I(new_n21901_), .ZN(new_n21902_));
  NAND2_X1   g21605(.A1(new_n21900_), .A2(new_n21898_), .ZN(new_n21903_));
  NAND2_X1   g21606(.A1(new_n21902_), .A2(new_n21903_), .ZN(new_n21904_));
  XNOR2_X1   g21607(.A1(new_n21900_), .A2(new_n21898_), .ZN(new_n21905_));
  NOR2_X1    g21608(.A1(new_n21905_), .A2(new_n21895_), .ZN(new_n21906_));
  AOI21_X1   g21609(.A1(new_n21895_), .A2(new_n21904_), .B(new_n21906_), .ZN(new_n21907_));
  XNOR2_X1   g21610(.A1(new_n21855_), .A2(new_n21907_), .ZN(new_n21908_));
  NOR2_X1    g21611(.A1(new_n21908_), .A2(new_n21853_), .ZN(new_n21909_));
  INV_X1     g21612(.I(new_n21853_), .ZN(new_n21910_));
  NOR2_X1    g21613(.A1(new_n21855_), .A2(new_n21907_), .ZN(new_n21911_));
  INV_X1     g21614(.I(new_n21911_), .ZN(new_n21912_));
  NAND2_X1   g21615(.A1(new_n21855_), .A2(new_n21907_), .ZN(new_n21913_));
  AOI21_X1   g21616(.A1(new_n21912_), .A2(new_n21913_), .B(new_n21910_), .ZN(new_n21914_));
  NOR2_X1    g21617(.A1(new_n21914_), .A2(new_n21909_), .ZN(new_n21915_));
  OAI22_X1   g21618(.A1(new_n7619_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n8309_), .ZN(new_n21916_));
  OAI21_X1   g21619(.A1(new_n7864_), .A2(new_n7947_), .B(new_n21916_), .ZN(new_n21917_));
  AOI21_X1   g21620(.A1(new_n21917_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n21918_));
  XOR2_X1    g21621(.A1(new_n8217_), .A2(new_n21918_), .Z(new_n21919_));
  AOI21_X1   g21622(.A1(new_n21740_), .A2(new_n21738_), .B(new_n21736_), .ZN(new_n21920_));
  XNOR2_X1   g21623(.A1(new_n21920_), .A2(new_n21919_), .ZN(new_n21921_));
  NOR2_X1    g21624(.A1(new_n21921_), .A2(new_n21915_), .ZN(new_n21922_));
  NOR2_X1    g21625(.A1(new_n21920_), .A2(new_n21919_), .ZN(new_n21923_));
  INV_X1     g21626(.I(new_n21923_), .ZN(new_n21924_));
  NAND2_X1   g21627(.A1(new_n21920_), .A2(new_n21919_), .ZN(new_n21925_));
  NAND2_X1   g21628(.A1(new_n21924_), .A2(new_n21925_), .ZN(new_n21926_));
  AOI21_X1   g21629(.A1(new_n21915_), .A2(new_n21926_), .B(new_n21922_), .ZN(new_n21927_));
  AOI21_X1   g21630(.A1(new_n21750_), .A2(new_n21748_), .B(new_n21746_), .ZN(new_n21928_));
  XNOR2_X1   g21631(.A1(new_n21927_), .A2(new_n21928_), .ZN(new_n21929_));
  NOR2_X1    g21632(.A1(new_n21929_), .A2(new_n21849_), .ZN(new_n21930_));
  INV_X1     g21633(.I(new_n21849_), .ZN(new_n21931_));
  NOR2_X1    g21634(.A1(new_n21927_), .A2(new_n21928_), .ZN(new_n21932_));
  INV_X1     g21635(.I(new_n21932_), .ZN(new_n21933_));
  NAND2_X1   g21636(.A1(new_n21927_), .A2(new_n21928_), .ZN(new_n21934_));
  AOI21_X1   g21637(.A1(new_n21933_), .A2(new_n21934_), .B(new_n21931_), .ZN(new_n21935_));
  NOR2_X1    g21638(.A1(new_n21930_), .A2(new_n21935_), .ZN(new_n21936_));
  NOR2_X1    g21639(.A1(new_n21763_), .A2(new_n21753_), .ZN(new_n21937_));
  NOR2_X1    g21640(.A1(new_n21937_), .A2(new_n21761_), .ZN(new_n21938_));
  XOR2_X1    g21641(.A1(new_n21936_), .A2(new_n21938_), .Z(new_n21939_));
  NOR2_X1    g21642(.A1(new_n21939_), .A2(new_n21845_), .ZN(new_n21940_));
  INV_X1     g21643(.I(new_n21845_), .ZN(new_n21941_));
  INV_X1     g21644(.I(new_n21936_), .ZN(new_n21942_));
  NOR2_X1    g21645(.A1(new_n21942_), .A2(new_n21938_), .ZN(new_n21943_));
  INV_X1     g21646(.I(new_n21943_), .ZN(new_n21944_));
  NAND2_X1   g21647(.A1(new_n21942_), .A2(new_n21938_), .ZN(new_n21945_));
  AOI21_X1   g21648(.A1(new_n21944_), .A2(new_n21945_), .B(new_n21941_), .ZN(new_n21946_));
  NOR2_X1    g21649(.A1(new_n21946_), .A2(new_n21940_), .ZN(new_n21947_));
  XOR2_X1    g21650(.A1(new_n21947_), .A2(new_n21841_), .Z(new_n21948_));
  NOR2_X1    g21651(.A1(new_n21948_), .A2(new_n21839_), .ZN(new_n21949_));
  INV_X1     g21652(.I(new_n21841_), .ZN(new_n21950_));
  NOR2_X1    g21653(.A1(new_n21947_), .A2(new_n21950_), .ZN(new_n21951_));
  INV_X1     g21654(.I(new_n21951_), .ZN(new_n21952_));
  NAND2_X1   g21655(.A1(new_n21947_), .A2(new_n21950_), .ZN(new_n21953_));
  NAND2_X1   g21656(.A1(new_n21952_), .A2(new_n21953_), .ZN(new_n21954_));
  AOI21_X1   g21657(.A1(new_n21839_), .A2(new_n21954_), .B(new_n21949_), .ZN(new_n21955_));
  OAI22_X1   g21658(.A1(new_n4072_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n4067_), .ZN(new_n21956_));
  OAI21_X1   g21659(.A1(new_n12536_), .A2(new_n4318_), .B(new_n21956_), .ZN(new_n21957_));
  AOI21_X1   g21660(.A1(new_n21957_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n21958_));
  XOR2_X1    g21661(.A1(new_n12969_), .A2(new_n21958_), .Z(new_n21959_));
  AOI21_X1   g21662(.A1(new_n21784_), .A2(new_n21788_), .B(new_n21786_), .ZN(new_n21960_));
  XNOR2_X1   g21663(.A1(new_n21960_), .A2(new_n21959_), .ZN(new_n21961_));
  NOR2_X1    g21664(.A1(new_n21961_), .A2(new_n21955_), .ZN(new_n21962_));
  NOR2_X1    g21665(.A1(new_n21960_), .A2(new_n21959_), .ZN(new_n21963_));
  INV_X1     g21666(.I(new_n21963_), .ZN(new_n21964_));
  NAND2_X1   g21667(.A1(new_n21960_), .A2(new_n21959_), .ZN(new_n21965_));
  NAND2_X1   g21668(.A1(new_n21964_), .A2(new_n21965_), .ZN(new_n21966_));
  AOI21_X1   g21669(.A1(new_n21955_), .A2(new_n21966_), .B(new_n21962_), .ZN(new_n21967_));
  XNOR2_X1   g21670(.A1(new_n21967_), .A2(new_n21835_), .ZN(new_n21968_));
  NOR2_X1    g21671(.A1(new_n21967_), .A2(new_n21835_), .ZN(new_n21969_));
  NAND2_X1   g21672(.A1(new_n21967_), .A2(new_n21835_), .ZN(new_n21970_));
  INV_X1     g21673(.I(new_n21970_), .ZN(new_n21971_));
  OAI21_X1   g21674(.A1(new_n21971_), .A2(new_n21969_), .B(new_n21833_), .ZN(new_n21972_));
  OAI21_X1   g21675(.A1(new_n21833_), .A2(new_n21968_), .B(new_n21972_), .ZN(new_n21973_));
  OAI21_X1   g21676(.A1(new_n2705_), .A2(new_n2884_), .B(new_n16487_), .ZN(new_n21974_));
  NAND2_X1   g21677(.A1(new_n21805_), .A2(new_n21802_), .ZN(new_n21975_));
  NAND2_X1   g21678(.A1(new_n21975_), .A2(new_n21804_), .ZN(new_n21976_));
  XOR2_X1    g21679(.A1(new_n21976_), .A2(new_n21974_), .Z(new_n21977_));
  XOR2_X1    g21680(.A1(new_n21977_), .A2(new_n21973_), .Z(new_n21978_));
  XOR2_X1    g21681(.A1(new_n21978_), .A2(new_n2702_), .Z(new_n21979_));
  NOR2_X1    g21682(.A1(new_n21979_), .A2(new_n21829_), .ZN(new_n21980_));
  INV_X1     g21683(.I(new_n21980_), .ZN(new_n21981_));
  NAND2_X1   g21684(.A1(new_n21979_), .A2(new_n21829_), .ZN(new_n21982_));
  NAND2_X1   g21685(.A1(new_n21981_), .A2(new_n21982_), .ZN(new_n21983_));
  XOR2_X1    g21686(.A1(new_n21826_), .A2(new_n21983_), .Z(\f[92] ));
  NAND2_X1   g21687(.A1(new_n21973_), .A2(new_n21976_), .ZN(new_n21985_));
  XOR2_X1    g21688(.A1(new_n21974_), .A2(\a[29] ), .Z(new_n21986_));
  OAI21_X1   g21689(.A1(new_n21973_), .A2(new_n21976_), .B(new_n21986_), .ZN(new_n21987_));
  NAND2_X1   g21690(.A1(new_n21987_), .A2(new_n21985_), .ZN(new_n21988_));
  NOR2_X1    g21691(.A1(new_n21971_), .A2(new_n21833_), .ZN(new_n21989_));
  OAI22_X1   g21692(.A1(new_n14208_), .A2(new_n3357_), .B1(new_n3352_), .B2(new_n14592_), .ZN(new_n21990_));
  OAI21_X1   g21693(.A1(new_n13785_), .A2(new_n3569_), .B(new_n21990_), .ZN(new_n21991_));
  AOI21_X1   g21694(.A1(new_n21991_), .A2(new_n3354_), .B(new_n3357_), .ZN(new_n21992_));
  XNOR2_X1   g21695(.A1(new_n14599_), .A2(new_n21992_), .ZN(new_n21993_));
  OAI21_X1   g21696(.A1(new_n21839_), .A2(new_n21951_), .B(new_n21953_), .ZN(new_n21994_));
  AOI21_X1   g21697(.A1(new_n21941_), .A2(new_n21945_), .B(new_n21943_), .ZN(new_n21995_));
  AOI21_X1   g21698(.A1(new_n21931_), .A2(new_n21934_), .B(new_n21932_), .ZN(new_n21996_));
  INV_X1     g21699(.I(new_n21996_), .ZN(new_n21997_));
  NAND2_X1   g21700(.A1(new_n21913_), .A2(new_n21910_), .ZN(new_n21998_));
  AOI21_X1   g21701(.A1(new_n21895_), .A2(new_n21903_), .B(new_n21901_), .ZN(new_n21999_));
  NOR2_X1    g21702(.A1(new_n21890_), .A2(new_n21858_), .ZN(new_n22000_));
  NOR2_X1    g21703(.A1(new_n22000_), .A2(new_n21891_), .ZN(new_n22001_));
  AOI21_X1   g21704(.A1(new_n21884_), .A2(new_n21887_), .B(new_n21885_), .ZN(new_n22002_));
  AOI21_X1   g21705(.A1(new_n21865_), .A2(new_n21871_), .B(new_n21873_), .ZN(new_n22003_));
  OAI22_X1   g21706(.A1(new_n13880_), .A2(new_n4248_), .B1(new_n3709_), .B2(new_n13885_), .ZN(new_n22004_));
  AOI21_X1   g21707(.A1(new_n22004_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n22005_));
  XNOR2_X1   g21708(.A1(new_n3993_), .A2(new_n22005_), .ZN(new_n22006_));
  NOR2_X1    g21709(.A1(new_n13476_), .A2(new_n3018_), .ZN(new_n22007_));
  XOR2_X1    g21710(.A1(new_n14736_), .A2(new_n3018_), .Z(new_n22008_));
  NAND2_X1   g21711(.A1(new_n22008_), .A2(\b[30] ), .ZN(new_n22009_));
  XOR2_X1    g21712(.A1(new_n22009_), .A2(new_n22007_), .Z(new_n22010_));
  NOR2_X1    g21713(.A1(new_n22010_), .A2(new_n2702_), .ZN(new_n22011_));
  INV_X1     g21714(.I(new_n22011_), .ZN(new_n22012_));
  NAND2_X1   g21715(.A1(new_n22010_), .A2(new_n2702_), .ZN(new_n22013_));
  AOI21_X1   g21716(.A1(new_n22012_), .A2(new_n22013_), .B(new_n21869_), .ZN(new_n22014_));
  XOR2_X1    g21717(.A1(new_n22010_), .A2(\a[29] ), .Z(new_n22015_));
  NOR2_X1    g21718(.A1(new_n22015_), .A2(new_n21872_), .ZN(new_n22016_));
  NOR2_X1    g21719(.A1(new_n22016_), .A2(new_n22014_), .ZN(new_n22017_));
  NOR2_X1    g21720(.A1(new_n22006_), .A2(new_n22017_), .ZN(new_n22018_));
  AND2_X2    g21721(.A1(new_n22006_), .A2(new_n22017_), .Z(new_n22019_));
  NOR2_X1    g21722(.A1(new_n22019_), .A2(new_n22018_), .ZN(new_n22020_));
  NOR2_X1    g21723(.A1(new_n22020_), .A2(new_n22003_), .ZN(new_n22021_));
  INV_X1     g21724(.I(new_n22003_), .ZN(new_n22022_));
  XNOR2_X1   g21725(.A1(new_n22006_), .A2(new_n22017_), .ZN(new_n22023_));
  NOR2_X1    g21726(.A1(new_n22023_), .A2(new_n22022_), .ZN(new_n22024_));
  NOR2_X1    g21727(.A1(new_n22021_), .A2(new_n22024_), .ZN(new_n22025_));
  AOI22_X1   g21728(.A1(new_n13078_), .A2(\b[34] ), .B1(new_n20981_), .B2(new_n12218_), .ZN(new_n22026_));
  OAI21_X1   g21729(.A1(new_n22026_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22027_));
  XOR2_X1    g21730(.A1(new_n4778_), .A2(new_n22027_), .Z(new_n22028_));
  XNOR2_X1   g21731(.A1(new_n22025_), .A2(new_n22028_), .ZN(new_n22029_));
  NOR2_X1    g21732(.A1(new_n22029_), .A2(new_n22002_), .ZN(new_n22030_));
  INV_X1     g21733(.I(new_n22002_), .ZN(new_n22031_));
  NOR2_X1    g21734(.A1(new_n22025_), .A2(new_n22028_), .ZN(new_n22032_));
  INV_X1     g21735(.I(new_n22032_), .ZN(new_n22033_));
  NAND2_X1   g21736(.A1(new_n22025_), .A2(new_n22028_), .ZN(new_n22034_));
  AOI21_X1   g21737(.A1(new_n22033_), .A2(new_n22034_), .B(new_n22031_), .ZN(new_n22035_));
  NOR2_X1    g21738(.A1(new_n22030_), .A2(new_n22035_), .ZN(new_n22036_));
  AOI22_X1   g21739(.A1(new_n10969_), .A2(new_n5915_), .B1(new_n11394_), .B2(\b[37] ), .ZN(new_n22037_));
  OAI21_X1   g21740(.A1(new_n22037_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22038_));
  XOR2_X1    g21741(.A1(new_n5600_), .A2(new_n22038_), .Z(new_n22039_));
  XOR2_X1    g21742(.A1(new_n22036_), .A2(new_n22039_), .Z(new_n22040_));
  NOR3_X1    g21743(.A1(new_n22030_), .A2(new_n22035_), .A3(new_n22039_), .ZN(new_n22041_));
  INV_X1     g21744(.I(new_n22039_), .ZN(new_n22042_));
  NOR2_X1    g21745(.A1(new_n22036_), .A2(new_n22042_), .ZN(new_n22043_));
  OAI21_X1   g21746(.A1(new_n22043_), .A2(new_n22041_), .B(new_n22001_), .ZN(new_n22044_));
  OAI21_X1   g21747(.A1(new_n22001_), .A2(new_n22040_), .B(new_n22044_), .ZN(new_n22045_));
  AOI22_X1   g21748(.A1(new_n11415_), .A2(new_n6540_), .B1(\b[40] ), .B2(new_n10145_), .ZN(new_n22046_));
  OAI21_X1   g21749(.A1(new_n22046_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22047_));
  XNOR2_X1   g21750(.A1(new_n6543_), .A2(new_n22047_), .ZN(new_n22048_));
  NOR2_X1    g21751(.A1(new_n22045_), .A2(new_n22048_), .ZN(new_n22049_));
  INV_X1     g21752(.I(new_n22049_), .ZN(new_n22050_));
  NAND2_X1   g21753(.A1(new_n22045_), .A2(new_n22048_), .ZN(new_n22051_));
  AOI21_X1   g21754(.A1(new_n22050_), .A2(new_n22051_), .B(new_n21999_), .ZN(new_n22052_));
  XOR2_X1    g21755(.A1(new_n22045_), .A2(new_n22048_), .Z(new_n22053_));
  AOI21_X1   g21756(.A1(new_n21999_), .A2(new_n22053_), .B(new_n22052_), .ZN(new_n22054_));
  OAI22_X1   g21757(.A1(new_n8644_), .A2(new_n7198_), .B1(new_n7864_), .B2(new_n9388_), .ZN(new_n22055_));
  OAI21_X1   g21758(.A1(new_n6847_), .A2(new_n10154_), .B(new_n22055_), .ZN(new_n22056_));
  AOI21_X1   g21759(.A1(new_n22056_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n22057_));
  XOR2_X1    g21760(.A1(new_n7516_), .A2(new_n22057_), .Z(new_n22058_));
  XNOR2_X1   g21761(.A1(new_n22054_), .A2(new_n22058_), .ZN(new_n22059_));
  AOI21_X1   g21762(.A1(new_n21912_), .A2(new_n21998_), .B(new_n22059_), .ZN(new_n22060_));
  NAND2_X1   g21763(.A1(new_n21998_), .A2(new_n21912_), .ZN(new_n22061_));
  NOR2_X1    g21764(.A1(new_n22054_), .A2(new_n22058_), .ZN(new_n22062_));
  INV_X1     g21765(.I(new_n22062_), .ZN(new_n22063_));
  NAND2_X1   g21766(.A1(new_n22054_), .A2(new_n22058_), .ZN(new_n22064_));
  AOI21_X1   g21767(.A1(new_n22063_), .A2(new_n22064_), .B(new_n22061_), .ZN(new_n22065_));
  NOR2_X1    g21768(.A1(new_n22060_), .A2(new_n22065_), .ZN(new_n22066_));
  OAI22_X1   g21769(.A1(new_n7619_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n8309_), .ZN(new_n22067_));
  OAI21_X1   g21770(.A1(new_n7870_), .A2(new_n7947_), .B(new_n22067_), .ZN(new_n22068_));
  AOI21_X1   g21771(.A1(new_n22068_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22069_));
  XOR2_X1    g21772(.A1(new_n8568_), .A2(new_n22069_), .Z(new_n22070_));
  NAND2_X1   g21773(.A1(new_n21915_), .A2(new_n21925_), .ZN(new_n22071_));
  AOI21_X1   g21774(.A1(new_n22071_), .A2(new_n21924_), .B(new_n22070_), .ZN(new_n22072_));
  INV_X1     g21775(.I(new_n22072_), .ZN(new_n22073_));
  INV_X1     g21776(.I(new_n22070_), .ZN(new_n22074_));
  NAND2_X1   g21777(.A1(new_n22071_), .A2(new_n21924_), .ZN(new_n22075_));
  NOR2_X1    g21778(.A1(new_n22075_), .A2(new_n22074_), .ZN(new_n22076_));
  INV_X1     g21779(.I(new_n22076_), .ZN(new_n22077_));
  AOI21_X1   g21780(.A1(new_n22077_), .A2(new_n22073_), .B(new_n22066_), .ZN(new_n22078_));
  XOR2_X1    g21781(.A1(new_n22075_), .A2(new_n22070_), .Z(new_n22079_));
  NOR3_X1    g21782(.A1(new_n22079_), .A2(new_n22060_), .A3(new_n22065_), .ZN(new_n22080_));
  OAI22_X1   g21783(.A1(new_n6644_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n6647_), .ZN(new_n22081_));
  OAI21_X1   g21784(.A1(new_n8948_), .A2(new_n7284_), .B(new_n22081_), .ZN(new_n22082_));
  AOI21_X1   g21785(.A1(new_n22082_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22083_));
  XNOR2_X1   g21786(.A1(new_n9642_), .A2(new_n22083_), .ZN(new_n22084_));
  NOR3_X1    g21787(.A1(new_n22080_), .A2(new_n22078_), .A3(new_n22084_), .ZN(new_n22085_));
  NOR2_X1    g21788(.A1(new_n22080_), .A2(new_n22078_), .ZN(new_n22086_));
  INV_X1     g21789(.I(new_n22084_), .ZN(new_n22087_));
  NOR2_X1    g21790(.A1(new_n22086_), .A2(new_n22087_), .ZN(new_n22088_));
  OAI21_X1   g21791(.A1(new_n22088_), .A2(new_n22085_), .B(new_n21997_), .ZN(new_n22089_));
  XOR2_X1    g21792(.A1(new_n22086_), .A2(new_n22087_), .Z(new_n22090_));
  NAND2_X1   g21793(.A1(new_n22090_), .A2(new_n21996_), .ZN(new_n22091_));
  NAND2_X1   g21794(.A1(new_n22091_), .A2(new_n22089_), .ZN(new_n22092_));
  OAI22_X1   g21795(.A1(new_n5993_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n5991_), .ZN(new_n22093_));
  OAI21_X1   g21796(.A1(new_n10031_), .A2(new_n5997_), .B(new_n22093_), .ZN(new_n22094_));
  AOI21_X1   g21797(.A1(new_n22094_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n22095_));
  XNOR2_X1   g21798(.A1(new_n10866_), .A2(new_n22095_), .ZN(new_n22096_));
  XOR2_X1    g21799(.A1(new_n22092_), .A2(new_n22096_), .Z(new_n22097_));
  AOI21_X1   g21800(.A1(new_n22091_), .A2(new_n22089_), .B(new_n22096_), .ZN(new_n22098_));
  INV_X1     g21801(.I(new_n22096_), .ZN(new_n22099_));
  NOR2_X1    g21802(.A1(new_n22092_), .A2(new_n22099_), .ZN(new_n22100_));
  OAI21_X1   g21803(.A1(new_n22100_), .A2(new_n22098_), .B(new_n21995_), .ZN(new_n22101_));
  OAI21_X1   g21804(.A1(new_n22097_), .A2(new_n21995_), .B(new_n22101_), .ZN(new_n22102_));
  AOI22_X1   g21805(.A1(new_n4859_), .A2(\b[56] ), .B1(new_n4865_), .B2(\b[57] ), .ZN(new_n22103_));
  AOI21_X1   g21806(.A1(\b[55] ), .A2(new_n6005_), .B(new_n22103_), .ZN(new_n22104_));
  OAI21_X1   g21807(.A1(new_n22104_), .A2(\a[38] ), .B(new_n4859_), .ZN(new_n22105_));
  XOR2_X1    g21808(.A1(new_n12128_), .A2(new_n22105_), .Z(new_n22106_));
  XOR2_X1    g21809(.A1(new_n22102_), .A2(new_n22106_), .Z(new_n22107_));
  NOR2_X1    g21810(.A1(new_n22102_), .A2(new_n22106_), .ZN(new_n22108_));
  INV_X1     g21811(.I(new_n22108_), .ZN(new_n22109_));
  NAND2_X1   g21812(.A1(new_n22102_), .A2(new_n22106_), .ZN(new_n22110_));
  NAND2_X1   g21813(.A1(new_n22109_), .A2(new_n22110_), .ZN(new_n22111_));
  MUX2_X1    g21814(.I0(new_n22111_), .I1(new_n22107_), .S(new_n21994_), .Z(new_n22112_));
  OAI22_X1   g21815(.A1(new_n4072_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n4067_), .ZN(new_n22113_));
  OAI21_X1   g21816(.A1(new_n12542_), .A2(new_n4318_), .B(new_n22113_), .ZN(new_n22114_));
  AOI21_X1   g21817(.A1(new_n22114_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n22115_));
  XNOR2_X1   g21818(.A1(new_n13371_), .A2(new_n22115_), .ZN(new_n22116_));
  INV_X1     g21819(.I(new_n22116_), .ZN(new_n22117_));
  NAND2_X1   g21820(.A1(new_n21965_), .A2(new_n21955_), .ZN(new_n22118_));
  NAND2_X1   g21821(.A1(new_n22118_), .A2(new_n21964_), .ZN(new_n22119_));
  NAND2_X1   g21822(.A1(new_n22119_), .A2(new_n22117_), .ZN(new_n22120_));
  INV_X1     g21823(.I(new_n22120_), .ZN(new_n22121_));
  NOR2_X1    g21824(.A1(new_n22119_), .A2(new_n22117_), .ZN(new_n22122_));
  OAI21_X1   g21825(.A1(new_n22121_), .A2(new_n22122_), .B(new_n22112_), .ZN(new_n22123_));
  XOR2_X1    g21826(.A1(new_n22119_), .A2(new_n22116_), .Z(new_n22124_));
  OR2_X2     g21827(.A1(new_n22124_), .A2(new_n22112_), .Z(new_n22125_));
  NAND2_X1   g21828(.A1(new_n22125_), .A2(new_n22123_), .ZN(new_n22126_));
  XOR2_X1    g21829(.A1(new_n22126_), .A2(new_n21993_), .Z(new_n22127_));
  OAI21_X1   g21830(.A1(new_n21969_), .A2(new_n21989_), .B(new_n22127_), .ZN(new_n22128_));
  NOR2_X1    g21831(.A1(new_n21989_), .A2(new_n21969_), .ZN(new_n22129_));
  AND2_X2    g21832(.A1(new_n22126_), .A2(new_n21993_), .Z(new_n22130_));
  NOR2_X1    g21833(.A1(new_n22126_), .A2(new_n21993_), .ZN(new_n22131_));
  OAI21_X1   g21834(.A1(new_n22130_), .A2(new_n22131_), .B(new_n22129_), .ZN(new_n22132_));
  NAND2_X1   g21835(.A1(new_n22128_), .A2(new_n22132_), .ZN(new_n22133_));
  XOR2_X1    g21836(.A1(new_n22133_), .A2(new_n21988_), .Z(new_n22134_));
  OAI21_X1   g21837(.A1(new_n21982_), .A2(new_n22134_), .B(new_n21981_), .ZN(new_n22135_));
  XOR2_X1    g21838(.A1(new_n21826_), .A2(new_n22135_), .Z(\f[93] ));
  AOI21_X1   g21839(.A1(new_n22128_), .A2(new_n22132_), .B(new_n21988_), .ZN(new_n22137_));
  AOI21_X1   g21840(.A1(new_n21647_), .A2(new_n21824_), .B(new_n21822_), .ZN(new_n22138_));
  NAND2_X1   g21841(.A1(new_n21981_), .A2(new_n21982_), .ZN(new_n22139_));
  INV_X1     g21842(.I(new_n22139_), .ZN(new_n22140_));
  NOR2_X1    g21843(.A1(new_n22138_), .A2(new_n22140_), .ZN(new_n22141_));
  NOR2_X1    g21844(.A1(new_n3569_), .A2(new_n3352_), .ZN(new_n22142_));
  NAND2_X1   g21845(.A1(new_n16148_), .A2(new_n3354_), .ZN(new_n22143_));
  OAI21_X1   g21846(.A1(new_n22142_), .A2(new_n22143_), .B(new_n3346_), .ZN(new_n22144_));
  XNOR2_X1   g21847(.A1(new_n14978_), .A2(new_n22144_), .ZN(new_n22145_));
  OAI21_X1   g21848(.A1(new_n22112_), .A2(new_n22122_), .B(new_n22120_), .ZN(new_n22146_));
  OAI22_X1   g21849(.A1(new_n5420_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n5107_), .ZN(new_n22147_));
  OAI21_X1   g21850(.A1(new_n11744_), .A2(new_n5112_), .B(new_n22147_), .ZN(new_n22148_));
  AOI21_X1   g21851(.A1(new_n22148_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n22149_));
  XNOR2_X1   g21852(.A1(new_n12546_), .A2(new_n22149_), .ZN(new_n22150_));
  NOR2_X1    g21853(.A1(new_n22100_), .A2(new_n21995_), .ZN(new_n22151_));
  NOR2_X1    g21854(.A1(new_n22088_), .A2(new_n21996_), .ZN(new_n22152_));
  NOR2_X1    g21855(.A1(new_n22152_), .A2(new_n22085_), .ZN(new_n22153_));
  OAI22_X1   g21856(.A1(new_n6644_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n6647_), .ZN(new_n22154_));
  OAI21_X1   g21857(.A1(new_n9295_), .A2(new_n7284_), .B(new_n22154_), .ZN(new_n22155_));
  AOI21_X1   g21858(.A1(new_n22155_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22156_));
  XNOR2_X1   g21859(.A1(new_n10035_), .A2(new_n22156_), .ZN(new_n22157_));
  INV_X1     g21860(.I(new_n22157_), .ZN(new_n22158_));
  AOI22_X1   g21861(.A1(new_n8631_), .A2(\b[45] ), .B1(\b[46] ), .B2(new_n9382_), .ZN(new_n22159_));
  AOI21_X1   g21862(.A1(\b[44] ), .A2(new_n9731_), .B(new_n22159_), .ZN(new_n22160_));
  OAI21_X1   g21863(.A1(new_n22160_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n22161_));
  XOR2_X1    g21864(.A1(new_n7874_), .A2(new_n22161_), .Z(new_n22162_));
  NOR2_X1    g21865(.A1(new_n22043_), .A2(new_n22001_), .ZN(new_n22163_));
  NOR2_X1    g21866(.A1(new_n22163_), .A2(new_n22041_), .ZN(new_n22164_));
  AOI22_X1   g21867(.A1(new_n10969_), .A2(new_n5923_), .B1(new_n11394_), .B2(\b[38] ), .ZN(new_n22165_));
  OAI21_X1   g21868(.A1(new_n22165_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22166_));
  XNOR2_X1   g21869(.A1(new_n5926_), .A2(new_n22166_), .ZN(new_n22167_));
  NAND2_X1   g21870(.A1(new_n22034_), .A2(new_n22031_), .ZN(new_n22168_));
  NAND2_X1   g21871(.A1(new_n22168_), .A2(new_n22033_), .ZN(new_n22169_));
  AOI22_X1   g21872(.A1(new_n13078_), .A2(\b[35] ), .B1(new_n5349_), .B2(new_n12218_), .ZN(new_n22170_));
  OAI21_X1   g21873(.A1(new_n22170_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22171_));
  XNOR2_X1   g21874(.A1(new_n5067_), .A2(new_n22171_), .ZN(new_n22172_));
  INV_X1     g21875(.I(new_n22019_), .ZN(new_n22173_));
  AOI21_X1   g21876(.A1(new_n22173_), .A2(new_n22022_), .B(new_n22018_), .ZN(new_n22174_));
  OAI22_X1   g21877(.A1(new_n13880_), .A2(new_n4254_), .B1(new_n3717_), .B2(new_n13885_), .ZN(new_n22175_));
  AOI21_X1   g21878(.A1(new_n22175_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n22176_));
  XNOR2_X1   g21879(.A1(new_n4257_), .A2(new_n22176_), .ZN(new_n22177_));
  NAND2_X1   g21880(.A1(new_n22013_), .A2(new_n21872_), .ZN(new_n22178_));
  NAND2_X1   g21881(.A1(new_n22178_), .A2(new_n22012_), .ZN(new_n22179_));
  NOR2_X1    g21882(.A1(new_n13476_), .A2(new_n3260_), .ZN(new_n22180_));
  XOR2_X1    g21883(.A1(new_n14736_), .A2(new_n3260_), .Z(new_n22181_));
  NAND2_X1   g21884(.A1(new_n22181_), .A2(\b[31] ), .ZN(new_n22182_));
  XOR2_X1    g21885(.A1(new_n22182_), .A2(new_n22180_), .Z(new_n22183_));
  INV_X1     g21886(.I(new_n22183_), .ZN(new_n22184_));
  XOR2_X1    g21887(.A1(new_n22179_), .A2(new_n22184_), .Z(new_n22185_));
  NOR2_X1    g21888(.A1(new_n22177_), .A2(new_n22185_), .ZN(new_n22186_));
  NOR2_X1    g21889(.A1(new_n22179_), .A2(new_n22183_), .ZN(new_n22187_));
  INV_X1     g21890(.I(new_n22187_), .ZN(new_n22188_));
  NAND2_X1   g21891(.A1(new_n22179_), .A2(new_n22183_), .ZN(new_n22189_));
  NAND2_X1   g21892(.A1(new_n22188_), .A2(new_n22189_), .ZN(new_n22190_));
  AOI21_X1   g21893(.A1(new_n22177_), .A2(new_n22190_), .B(new_n22186_), .ZN(new_n22191_));
  XOR2_X1    g21894(.A1(new_n22191_), .A2(new_n22174_), .Z(new_n22192_));
  NOR2_X1    g21895(.A1(new_n22192_), .A2(new_n22172_), .ZN(new_n22193_));
  INV_X1     g21896(.I(new_n22174_), .ZN(new_n22194_));
  NOR2_X1    g21897(.A1(new_n22191_), .A2(new_n22194_), .ZN(new_n22195_));
  INV_X1     g21898(.I(new_n22195_), .ZN(new_n22196_));
  NAND2_X1   g21899(.A1(new_n22191_), .A2(new_n22194_), .ZN(new_n22197_));
  NAND2_X1   g21900(.A1(new_n22196_), .A2(new_n22197_), .ZN(new_n22198_));
  AOI21_X1   g21901(.A1(new_n22172_), .A2(new_n22198_), .B(new_n22193_), .ZN(new_n22199_));
  XNOR2_X1   g21902(.A1(new_n22199_), .A2(new_n22169_), .ZN(new_n22200_));
  NOR2_X1    g21903(.A1(new_n22199_), .A2(new_n22169_), .ZN(new_n22201_));
  NAND2_X1   g21904(.A1(new_n22199_), .A2(new_n22169_), .ZN(new_n22202_));
  INV_X1     g21905(.I(new_n22202_), .ZN(new_n22203_));
  OAI21_X1   g21906(.A1(new_n22203_), .A2(new_n22201_), .B(new_n22167_), .ZN(new_n22204_));
  OAI21_X1   g21907(.A1(new_n22167_), .A2(new_n22200_), .B(new_n22204_), .ZN(new_n22205_));
  AOI22_X1   g21908(.A1(new_n11415_), .A2(new_n7194_), .B1(\b[41] ), .B2(new_n10145_), .ZN(new_n22206_));
  OAI21_X1   g21909(.A1(new_n22206_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22207_));
  XNOR2_X1   g21910(.A1(new_n6851_), .A2(new_n22207_), .ZN(new_n22208_));
  NOR2_X1    g21911(.A1(new_n22205_), .A2(new_n22208_), .ZN(new_n22209_));
  INV_X1     g21912(.I(new_n22209_), .ZN(new_n22210_));
  NAND2_X1   g21913(.A1(new_n22205_), .A2(new_n22208_), .ZN(new_n22211_));
  AOI21_X1   g21914(.A1(new_n22210_), .A2(new_n22211_), .B(new_n22164_), .ZN(new_n22212_));
  INV_X1     g21915(.I(new_n22164_), .ZN(new_n22213_));
  XNOR2_X1   g21916(.A1(new_n22205_), .A2(new_n22208_), .ZN(new_n22214_));
  NOR2_X1    g21917(.A1(new_n22214_), .A2(new_n22213_), .ZN(new_n22215_));
  NOR2_X1    g21918(.A1(new_n22215_), .A2(new_n22212_), .ZN(new_n22216_));
  INV_X1     g21919(.I(new_n21999_), .ZN(new_n22217_));
  AOI21_X1   g21920(.A1(new_n22217_), .A2(new_n22051_), .B(new_n22049_), .ZN(new_n22218_));
  NOR2_X1    g21921(.A1(new_n22216_), .A2(new_n22218_), .ZN(new_n22219_));
  INV_X1     g21922(.I(new_n22219_), .ZN(new_n22220_));
  NAND2_X1   g21923(.A1(new_n22216_), .A2(new_n22218_), .ZN(new_n22221_));
  AOI21_X1   g21924(.A1(new_n22220_), .A2(new_n22221_), .B(new_n22162_), .ZN(new_n22222_));
  INV_X1     g21925(.I(new_n22162_), .ZN(new_n22223_));
  XNOR2_X1   g21926(.A1(new_n22216_), .A2(new_n22218_), .ZN(new_n22224_));
  NOR2_X1    g21927(.A1(new_n22224_), .A2(new_n22223_), .ZN(new_n22225_));
  NOR2_X1    g21928(.A1(new_n22225_), .A2(new_n22222_), .ZN(new_n22226_));
  NAND2_X1   g21929(.A1(new_n22064_), .A2(new_n22061_), .ZN(new_n22227_));
  NAND2_X1   g21930(.A1(new_n22227_), .A2(new_n22063_), .ZN(new_n22228_));
  INV_X1     g21931(.I(new_n22228_), .ZN(new_n22229_));
  OAI22_X1   g21932(.A1(new_n7619_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n8309_), .ZN(new_n22230_));
  OAI21_X1   g21933(.A1(new_n8218_), .A2(new_n7947_), .B(new_n22230_), .ZN(new_n22231_));
  AOI21_X1   g21934(.A1(new_n22231_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22232_));
  XOR2_X1    g21935(.A1(new_n8952_), .A2(new_n22232_), .Z(new_n22233_));
  NOR2_X1    g21936(.A1(new_n22229_), .A2(new_n22233_), .ZN(new_n22234_));
  INV_X1     g21937(.I(new_n22233_), .ZN(new_n22235_));
  NOR2_X1    g21938(.A1(new_n22228_), .A2(new_n22235_), .ZN(new_n22236_));
  NOR2_X1    g21939(.A1(new_n22234_), .A2(new_n22236_), .ZN(new_n22237_));
  NOR2_X1    g21940(.A1(new_n22226_), .A2(new_n22237_), .ZN(new_n22238_));
  INV_X1     g21941(.I(new_n22226_), .ZN(new_n22239_));
  XOR2_X1    g21942(.A1(new_n22228_), .A2(new_n22233_), .Z(new_n22240_));
  NOR2_X1    g21943(.A1(new_n22239_), .A2(new_n22240_), .ZN(new_n22241_));
  NOR2_X1    g21944(.A1(new_n22241_), .A2(new_n22238_), .ZN(new_n22242_));
  NAND2_X1   g21945(.A1(new_n22077_), .A2(new_n22066_), .ZN(new_n22243_));
  AOI21_X1   g21946(.A1(new_n22073_), .A2(new_n22243_), .B(new_n22242_), .ZN(new_n22244_));
  NAND2_X1   g21947(.A1(new_n22243_), .A2(new_n22073_), .ZN(new_n22245_));
  NOR3_X1    g21948(.A1(new_n22245_), .A2(new_n22241_), .A3(new_n22238_), .ZN(new_n22246_));
  OAI21_X1   g21949(.A1(new_n22244_), .A2(new_n22246_), .B(new_n22158_), .ZN(new_n22247_));
  XNOR2_X1   g21950(.A1(new_n22242_), .A2(new_n22245_), .ZN(new_n22248_));
  NAND2_X1   g21951(.A1(new_n22248_), .A2(new_n22157_), .ZN(new_n22249_));
  NAND2_X1   g21952(.A1(new_n22249_), .A2(new_n22247_), .ZN(new_n22250_));
  OAI22_X1   g21953(.A1(new_n5993_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n5991_), .ZN(new_n22251_));
  OAI21_X1   g21954(.A1(new_n10477_), .A2(new_n5997_), .B(new_n22251_), .ZN(new_n22252_));
  AOI21_X1   g21955(.A1(new_n22252_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n22253_));
  XOR2_X1    g21956(.A1(new_n11298_), .A2(new_n22253_), .Z(new_n22254_));
  XOR2_X1    g21957(.A1(new_n22250_), .A2(new_n22254_), .Z(new_n22255_));
  NOR2_X1    g21958(.A1(new_n22255_), .A2(new_n22153_), .ZN(new_n22256_));
  INV_X1     g21959(.I(new_n22153_), .ZN(new_n22257_));
  INV_X1     g21960(.I(new_n22250_), .ZN(new_n22258_));
  NOR2_X1    g21961(.A1(new_n22258_), .A2(new_n22254_), .ZN(new_n22259_));
  INV_X1     g21962(.I(new_n22259_), .ZN(new_n22260_));
  NAND2_X1   g21963(.A1(new_n22258_), .A2(new_n22254_), .ZN(new_n22261_));
  AOI21_X1   g21964(.A1(new_n22260_), .A2(new_n22261_), .B(new_n22257_), .ZN(new_n22262_));
  NOR2_X1    g21965(.A1(new_n22262_), .A2(new_n22256_), .ZN(new_n22263_));
  NOR3_X1    g21966(.A1(new_n22263_), .A2(new_n22098_), .A3(new_n22151_), .ZN(new_n22264_));
  NOR2_X1    g21967(.A1(new_n22151_), .A2(new_n22098_), .ZN(new_n22265_));
  INV_X1     g21968(.I(new_n22263_), .ZN(new_n22266_));
  NOR2_X1    g21969(.A1(new_n22266_), .A2(new_n22265_), .ZN(new_n22267_));
  NOR2_X1    g21970(.A1(new_n22267_), .A2(new_n22264_), .ZN(new_n22268_));
  NOR2_X1    g21971(.A1(new_n22268_), .A2(new_n22150_), .ZN(new_n22269_));
  INV_X1     g21972(.I(new_n22150_), .ZN(new_n22270_));
  XOR2_X1    g21973(.A1(new_n22263_), .A2(new_n22265_), .Z(new_n22271_));
  NOR2_X1    g21974(.A1(new_n22271_), .A2(new_n22270_), .ZN(new_n22272_));
  NOR2_X1    g21975(.A1(new_n22269_), .A2(new_n22272_), .ZN(new_n22273_));
  NAND2_X1   g21976(.A1(new_n22110_), .A2(new_n21994_), .ZN(new_n22274_));
  NAND2_X1   g21977(.A1(new_n22274_), .A2(new_n22109_), .ZN(new_n22275_));
  OAI22_X1   g21978(.A1(new_n4072_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n4067_), .ZN(new_n22276_));
  OAI21_X1   g21979(.A1(new_n12970_), .A2(new_n4318_), .B(new_n22276_), .ZN(new_n22277_));
  AOI21_X1   g21980(.A1(new_n22277_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n22278_));
  XOR2_X1    g21981(.A1(new_n13784_), .A2(new_n22278_), .Z(new_n22279_));
  XOR2_X1    g21982(.A1(new_n22275_), .A2(new_n22279_), .Z(new_n22280_));
  NOR2_X1    g21983(.A1(new_n22273_), .A2(new_n22280_), .ZN(new_n22281_));
  INV_X1     g21984(.I(new_n22273_), .ZN(new_n22282_));
  INV_X1     g21985(.I(new_n22275_), .ZN(new_n22283_));
  NOR2_X1    g21986(.A1(new_n22283_), .A2(new_n22279_), .ZN(new_n22284_));
  INV_X1     g21987(.I(new_n22284_), .ZN(new_n22285_));
  NAND2_X1   g21988(.A1(new_n22283_), .A2(new_n22279_), .ZN(new_n22286_));
  AOI21_X1   g21989(.A1(new_n22286_), .A2(new_n22285_), .B(new_n22282_), .ZN(new_n22287_));
  NOR2_X1    g21990(.A1(new_n22287_), .A2(new_n22281_), .ZN(new_n22288_));
  NOR2_X1    g21991(.A1(new_n22288_), .A2(new_n22146_), .ZN(new_n22289_));
  INV_X1     g21992(.I(new_n22146_), .ZN(new_n22290_));
  INV_X1     g21993(.I(new_n22288_), .ZN(new_n22291_));
  NOR2_X1    g21994(.A1(new_n22291_), .A2(new_n22290_), .ZN(new_n22292_));
  NOR2_X1    g21995(.A1(new_n22292_), .A2(new_n22289_), .ZN(new_n22293_));
  NOR2_X1    g21996(.A1(new_n22293_), .A2(new_n22145_), .ZN(new_n22294_));
  INV_X1     g21997(.I(new_n22145_), .ZN(new_n22295_));
  XOR2_X1    g21998(.A1(new_n22288_), .A2(new_n22290_), .Z(new_n22296_));
  NOR2_X1    g21999(.A1(new_n22296_), .A2(new_n22295_), .ZN(new_n22297_));
  NOR2_X1    g22000(.A1(new_n22294_), .A2(new_n22297_), .ZN(new_n22298_));
  NOR2_X1    g22001(.A1(new_n22130_), .A2(new_n22129_), .ZN(new_n22299_));
  NOR2_X1    g22002(.A1(new_n22299_), .A2(new_n22131_), .ZN(new_n22300_));
  NOR2_X1    g22003(.A1(new_n22300_), .A2(new_n22298_), .ZN(new_n22301_));
  XOR2_X1    g22004(.A1(new_n22141_), .A2(new_n22301_), .Z(new_n22302_));
  XOR2_X1    g22005(.A1(new_n22302_), .A2(new_n22137_), .Z(\f[94] ));
  INV_X1     g22006(.I(new_n22137_), .ZN(new_n22304_));
  NOR2_X1    g22007(.A1(new_n22304_), .A2(new_n22298_), .ZN(new_n22305_));
  INV_X1     g22008(.I(new_n22305_), .ZN(new_n22306_));
  AOI21_X1   g22009(.A1(new_n22304_), .A2(new_n22298_), .B(new_n22300_), .ZN(new_n22307_));
  NAND3_X1   g22010(.A1(new_n21826_), .A2(new_n22139_), .A3(new_n22307_), .ZN(new_n22308_));
  NAND2_X1   g22011(.A1(new_n22308_), .A2(new_n22306_), .ZN(new_n22309_));
  NOR2_X1    g22012(.A1(new_n22289_), .A2(new_n22145_), .ZN(new_n22310_));
  NOR2_X1    g22013(.A1(new_n22310_), .A2(new_n22292_), .ZN(new_n22311_));
  OAI22_X1   g22014(.A1(new_n4072_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n4067_), .ZN(new_n22312_));
  OAI21_X1   g22015(.A1(new_n13367_), .A2(new_n4318_), .B(new_n22312_), .ZN(new_n22313_));
  AOI21_X1   g22016(.A1(new_n22313_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n22314_));
  XOR2_X1    g22017(.A1(new_n14213_), .A2(new_n22314_), .Z(new_n22315_));
  OAI22_X1   g22018(.A1(new_n5993_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n5991_), .ZN(new_n22316_));
  OAI21_X1   g22019(.A1(new_n10862_), .A2(new_n5997_), .B(new_n22316_), .ZN(new_n22317_));
  AOI21_X1   g22020(.A1(new_n22317_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n22318_));
  XNOR2_X1   g22021(.A1(new_n11748_), .A2(new_n22318_), .ZN(new_n22319_));
  NOR2_X1    g22022(.A1(new_n22246_), .A2(new_n22157_), .ZN(new_n22320_));
  NOR2_X1    g22023(.A1(new_n22244_), .A2(new_n22320_), .ZN(new_n22321_));
  OAI22_X1   g22024(.A1(new_n6644_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n6647_), .ZN(new_n22322_));
  OAI21_X1   g22025(.A1(new_n10025_), .A2(new_n7284_), .B(new_n22322_), .ZN(new_n22323_));
  AOI21_X1   g22026(.A1(new_n22323_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22324_));
  XOR2_X1    g22027(.A1(new_n10476_), .A2(new_n22324_), .Z(new_n22325_));
  OAI22_X1   g22028(.A1(new_n7619_), .A2(new_n8948_), .B1(new_n9295_), .B2(new_n8309_), .ZN(new_n22326_));
  OAI21_X1   g22029(.A1(new_n8563_), .A2(new_n7947_), .B(new_n22326_), .ZN(new_n22327_));
  AOI21_X1   g22030(.A1(new_n22327_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22328_));
  XNOR2_X1   g22031(.A1(new_n9299_), .A2(new_n22328_), .ZN(new_n22329_));
  INV_X1     g22032(.I(new_n7199_), .ZN(new_n22330_));
  AOI22_X1   g22033(.A1(new_n11415_), .A2(new_n22330_), .B1(\b[42] ), .B2(new_n10145_), .ZN(new_n22331_));
  OAI21_X1   g22034(.A1(new_n22331_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22332_));
  XOR2_X1    g22035(.A1(new_n7202_), .A2(new_n22332_), .Z(new_n22333_));
  OAI21_X1   g22036(.A1(new_n22167_), .A2(new_n22201_), .B(new_n22202_), .ZN(new_n22334_));
  AOI22_X1   g22037(.A1(new_n10969_), .A2(new_n6532_), .B1(new_n11394_), .B2(\b[39] ), .ZN(new_n22335_));
  OAI21_X1   g22038(.A1(new_n22335_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22336_));
  XNOR2_X1   g22039(.A1(new_n6233_), .A2(new_n22336_), .ZN(new_n22337_));
  OAI21_X1   g22040(.A1(new_n22177_), .A2(new_n22187_), .B(new_n22189_), .ZN(new_n22338_));
  NOR2_X1    g22041(.A1(new_n13476_), .A2(new_n3709_), .ZN(new_n22339_));
  XOR2_X1    g22042(.A1(new_n14736_), .A2(new_n3709_), .Z(new_n22340_));
  NAND2_X1   g22043(.A1(new_n22340_), .A2(\b[32] ), .ZN(new_n22341_));
  XOR2_X1    g22044(.A1(new_n22341_), .A2(new_n22339_), .Z(new_n22342_));
  NOR2_X1    g22045(.A1(new_n22184_), .A2(new_n22342_), .ZN(new_n22343_));
  INV_X1     g22046(.I(new_n22342_), .ZN(new_n22344_));
  NOR2_X1    g22047(.A1(new_n22344_), .A2(new_n22183_), .ZN(new_n22345_));
  NOR2_X1    g22048(.A1(new_n22343_), .A2(new_n22345_), .ZN(new_n22346_));
  INV_X1     g22049(.I(new_n22346_), .ZN(new_n22347_));
  XOR2_X1    g22050(.A1(new_n22183_), .A2(new_n22342_), .Z(new_n22348_));
  NOR2_X1    g22051(.A1(new_n22338_), .A2(new_n22348_), .ZN(new_n22349_));
  AOI21_X1   g22052(.A1(new_n22338_), .A2(new_n22347_), .B(new_n22349_), .ZN(new_n22350_));
  AOI22_X1   g22053(.A1(new_n13078_), .A2(\b[36] ), .B1(new_n21317_), .B2(new_n12218_), .ZN(new_n22351_));
  OAI21_X1   g22054(.A1(new_n22351_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22352_));
  XOR2_X1    g22055(.A1(new_n5357_), .A2(new_n22352_), .Z(new_n22353_));
  OAI22_X1   g22056(.A1(new_n13880_), .A2(new_n4769_), .B1(new_n3989_), .B2(new_n13885_), .ZN(new_n22354_));
  AOI21_X1   g22057(.A1(new_n22354_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n22355_));
  XOR2_X1    g22058(.A1(new_n4499_), .A2(new_n22355_), .Z(new_n22356_));
  NOR2_X1    g22059(.A1(new_n22353_), .A2(new_n22356_), .ZN(new_n22357_));
  INV_X1     g22060(.I(new_n22357_), .ZN(new_n22358_));
  NAND2_X1   g22061(.A1(new_n22353_), .A2(new_n22356_), .ZN(new_n22359_));
  AOI21_X1   g22062(.A1(new_n22358_), .A2(new_n22359_), .B(new_n22350_), .ZN(new_n22360_));
  INV_X1     g22063(.I(new_n22350_), .ZN(new_n22361_));
  XNOR2_X1   g22064(.A1(new_n22353_), .A2(new_n22356_), .ZN(new_n22362_));
  NOR2_X1    g22065(.A1(new_n22362_), .A2(new_n22361_), .ZN(new_n22363_));
  NOR2_X1    g22066(.A1(new_n22363_), .A2(new_n22360_), .ZN(new_n22364_));
  OAI21_X1   g22067(.A1(new_n22172_), .A2(new_n22195_), .B(new_n22197_), .ZN(new_n22365_));
  XOR2_X1    g22068(.A1(new_n22364_), .A2(new_n22365_), .Z(new_n22366_));
  NOR2_X1    g22069(.A1(new_n22366_), .A2(new_n22337_), .ZN(new_n22367_));
  INV_X1     g22070(.I(new_n22337_), .ZN(new_n22368_));
  INV_X1     g22071(.I(new_n22365_), .ZN(new_n22369_));
  NOR2_X1    g22072(.A1(new_n22364_), .A2(new_n22369_), .ZN(new_n22370_));
  INV_X1     g22073(.I(new_n22370_), .ZN(new_n22371_));
  NAND2_X1   g22074(.A1(new_n22364_), .A2(new_n22369_), .ZN(new_n22372_));
  AOI21_X1   g22075(.A1(new_n22371_), .A2(new_n22372_), .B(new_n22368_), .ZN(new_n22373_));
  NOR2_X1    g22076(.A1(new_n22367_), .A2(new_n22373_), .ZN(new_n22374_));
  XNOR2_X1   g22077(.A1(new_n22374_), .A2(new_n22334_), .ZN(new_n22375_));
  NOR2_X1    g22078(.A1(new_n22375_), .A2(new_n22333_), .ZN(new_n22376_));
  NOR2_X1    g22079(.A1(new_n22374_), .A2(new_n22334_), .ZN(new_n22377_));
  INV_X1     g22080(.I(new_n22377_), .ZN(new_n22378_));
  NAND2_X1   g22081(.A1(new_n22374_), .A2(new_n22334_), .ZN(new_n22379_));
  NAND2_X1   g22082(.A1(new_n22378_), .A2(new_n22379_), .ZN(new_n22380_));
  AOI21_X1   g22083(.A1(new_n22333_), .A2(new_n22380_), .B(new_n22376_), .ZN(new_n22381_));
  OAI22_X1   g22084(.A1(new_n8644_), .A2(new_n7870_), .B1(new_n8218_), .B2(new_n9388_), .ZN(new_n22382_));
  OAI21_X1   g22085(.A1(new_n7864_), .A2(new_n10154_), .B(new_n22382_), .ZN(new_n22383_));
  AOI21_X1   g22086(.A1(new_n22383_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n22384_));
  XOR2_X1    g22087(.A1(new_n8217_), .A2(new_n22384_), .Z(new_n22385_));
  AOI21_X1   g22088(.A1(new_n22213_), .A2(new_n22211_), .B(new_n22209_), .ZN(new_n22386_));
  XNOR2_X1   g22089(.A1(new_n22386_), .A2(new_n22385_), .ZN(new_n22387_));
  NOR2_X1    g22090(.A1(new_n22381_), .A2(new_n22387_), .ZN(new_n22388_));
  NOR2_X1    g22091(.A1(new_n22386_), .A2(new_n22385_), .ZN(new_n22389_));
  INV_X1     g22092(.I(new_n22389_), .ZN(new_n22390_));
  NAND2_X1   g22093(.A1(new_n22386_), .A2(new_n22385_), .ZN(new_n22391_));
  NAND2_X1   g22094(.A1(new_n22390_), .A2(new_n22391_), .ZN(new_n22392_));
  AOI21_X1   g22095(.A1(new_n22381_), .A2(new_n22392_), .B(new_n22388_), .ZN(new_n22393_));
  AOI21_X1   g22096(.A1(new_n22223_), .A2(new_n22221_), .B(new_n22219_), .ZN(new_n22394_));
  XNOR2_X1   g22097(.A1(new_n22393_), .A2(new_n22394_), .ZN(new_n22395_));
  NOR2_X1    g22098(.A1(new_n22395_), .A2(new_n22329_), .ZN(new_n22396_));
  INV_X1     g22099(.I(new_n22329_), .ZN(new_n22397_));
  NOR2_X1    g22100(.A1(new_n22393_), .A2(new_n22394_), .ZN(new_n22398_));
  INV_X1     g22101(.I(new_n22398_), .ZN(new_n22399_));
  NAND2_X1   g22102(.A1(new_n22393_), .A2(new_n22394_), .ZN(new_n22400_));
  AOI21_X1   g22103(.A1(new_n22399_), .A2(new_n22400_), .B(new_n22397_), .ZN(new_n22401_));
  NOR2_X1    g22104(.A1(new_n22396_), .A2(new_n22401_), .ZN(new_n22402_));
  NOR2_X1    g22105(.A1(new_n22226_), .A2(new_n22236_), .ZN(new_n22403_));
  NOR2_X1    g22106(.A1(new_n22403_), .A2(new_n22234_), .ZN(new_n22404_));
  XOR2_X1    g22107(.A1(new_n22402_), .A2(new_n22404_), .Z(new_n22405_));
  NOR2_X1    g22108(.A1(new_n22405_), .A2(new_n22325_), .ZN(new_n22406_));
  INV_X1     g22109(.I(new_n22325_), .ZN(new_n22407_));
  INV_X1     g22110(.I(new_n22402_), .ZN(new_n22408_));
  NOR2_X1    g22111(.A1(new_n22408_), .A2(new_n22404_), .ZN(new_n22409_));
  INV_X1     g22112(.I(new_n22409_), .ZN(new_n22410_));
  NAND2_X1   g22113(.A1(new_n22408_), .A2(new_n22404_), .ZN(new_n22411_));
  AOI21_X1   g22114(.A1(new_n22410_), .A2(new_n22411_), .B(new_n22407_), .ZN(new_n22412_));
  NOR2_X1    g22115(.A1(new_n22412_), .A2(new_n22406_), .ZN(new_n22413_));
  XOR2_X1    g22116(.A1(new_n22413_), .A2(new_n22321_), .Z(new_n22414_));
  NOR2_X1    g22117(.A1(new_n22414_), .A2(new_n22319_), .ZN(new_n22415_));
  INV_X1     g22118(.I(new_n22321_), .ZN(new_n22416_));
  NOR2_X1    g22119(.A1(new_n22413_), .A2(new_n22416_), .ZN(new_n22417_));
  INV_X1     g22120(.I(new_n22417_), .ZN(new_n22418_));
  NAND2_X1   g22121(.A1(new_n22413_), .A2(new_n22416_), .ZN(new_n22419_));
  NAND2_X1   g22122(.A1(new_n22418_), .A2(new_n22419_), .ZN(new_n22420_));
  AOI21_X1   g22123(.A1(new_n22319_), .A2(new_n22420_), .B(new_n22415_), .ZN(new_n22421_));
  OAI22_X1   g22124(.A1(new_n5420_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n5107_), .ZN(new_n22422_));
  OAI21_X1   g22125(.A1(new_n12536_), .A2(new_n5112_), .B(new_n22422_), .ZN(new_n22423_));
  AOI21_X1   g22126(.A1(new_n22423_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n22424_));
  XOR2_X1    g22127(.A1(new_n12969_), .A2(new_n22424_), .Z(new_n22425_));
  AOI21_X1   g22128(.A1(new_n22257_), .A2(new_n22261_), .B(new_n22259_), .ZN(new_n22426_));
  XNOR2_X1   g22129(.A1(new_n22426_), .A2(new_n22425_), .ZN(new_n22427_));
  NOR2_X1    g22130(.A1(new_n22421_), .A2(new_n22427_), .ZN(new_n22428_));
  NOR2_X1    g22131(.A1(new_n22426_), .A2(new_n22425_), .ZN(new_n22429_));
  INV_X1     g22132(.I(new_n22429_), .ZN(new_n22430_));
  NAND2_X1   g22133(.A1(new_n22426_), .A2(new_n22425_), .ZN(new_n22431_));
  NAND2_X1   g22134(.A1(new_n22430_), .A2(new_n22431_), .ZN(new_n22432_));
  AOI21_X1   g22135(.A1(new_n22421_), .A2(new_n22432_), .B(new_n22428_), .ZN(new_n22433_));
  NOR2_X1    g22136(.A1(new_n22264_), .A2(new_n22150_), .ZN(new_n22434_));
  NOR2_X1    g22137(.A1(new_n22434_), .A2(new_n22267_), .ZN(new_n22435_));
  NOR2_X1    g22138(.A1(new_n22433_), .A2(new_n22435_), .ZN(new_n22436_));
  INV_X1     g22139(.I(new_n22436_), .ZN(new_n22437_));
  NAND2_X1   g22140(.A1(new_n22433_), .A2(new_n22435_), .ZN(new_n22438_));
  AOI21_X1   g22141(.A1(new_n22437_), .A2(new_n22438_), .B(new_n22315_), .ZN(new_n22439_));
  XOR2_X1    g22142(.A1(new_n22433_), .A2(new_n22435_), .Z(new_n22440_));
  AOI21_X1   g22143(.A1(new_n22315_), .A2(new_n22440_), .B(new_n22439_), .ZN(new_n22441_));
  OAI21_X1   g22144(.A1(new_n3357_), .A2(new_n3569_), .B(new_n16487_), .ZN(new_n22442_));
  NAND2_X1   g22145(.A1(new_n22282_), .A2(new_n22286_), .ZN(new_n22443_));
  NAND2_X1   g22146(.A1(new_n22443_), .A2(new_n22285_), .ZN(new_n22444_));
  XOR2_X1    g22147(.A1(new_n22444_), .A2(new_n22442_), .Z(new_n22445_));
  XOR2_X1    g22148(.A1(new_n22445_), .A2(new_n22441_), .Z(new_n22446_));
  XOR2_X1    g22149(.A1(new_n22446_), .A2(\a[32] ), .Z(new_n22447_));
  NOR2_X1    g22150(.A1(new_n22447_), .A2(new_n22311_), .ZN(new_n22448_));
  NAND2_X1   g22151(.A1(new_n22447_), .A2(new_n22311_), .ZN(new_n22449_));
  INV_X1     g22152(.I(new_n22449_), .ZN(new_n22450_));
  NOR2_X1    g22153(.A1(new_n22450_), .A2(new_n22448_), .ZN(new_n22451_));
  XNOR2_X1   g22154(.A1(new_n22309_), .A2(new_n22451_), .ZN(\f[95] ));
  INV_X1     g22155(.I(new_n22444_), .ZN(new_n22453_));
  NOR2_X1    g22156(.A1(new_n22441_), .A2(new_n22453_), .ZN(new_n22454_));
  XOR2_X1    g22157(.A1(new_n22442_), .A2(new_n3354_), .Z(new_n22455_));
  AOI21_X1   g22158(.A1(new_n22441_), .A2(new_n22453_), .B(new_n22455_), .ZN(new_n22456_));
  NOR2_X1    g22159(.A1(new_n22456_), .A2(new_n22454_), .ZN(new_n22457_));
  INV_X1     g22160(.I(new_n22315_), .ZN(new_n22458_));
  AOI21_X1   g22161(.A1(new_n22458_), .A2(new_n22438_), .B(new_n22436_), .ZN(new_n22459_));
  OAI22_X1   g22162(.A1(new_n4072_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n4067_), .ZN(new_n22460_));
  OAI21_X1   g22163(.A1(new_n13785_), .A2(new_n4318_), .B(new_n22460_), .ZN(new_n22461_));
  AOI21_X1   g22164(.A1(new_n22461_), .A2(new_n4069_), .B(new_n4072_), .ZN(new_n22462_));
  XNOR2_X1   g22165(.A1(new_n14599_), .A2(new_n22462_), .ZN(new_n22463_));
  INV_X1     g22166(.I(new_n22463_), .ZN(new_n22464_));
  OAI21_X1   g22167(.A1(new_n22319_), .A2(new_n22417_), .B(new_n22419_), .ZN(new_n22465_));
  AOI21_X1   g22168(.A1(new_n22407_), .A2(new_n22411_), .B(new_n22409_), .ZN(new_n22466_));
  AOI21_X1   g22169(.A1(new_n22397_), .A2(new_n22400_), .B(new_n22398_), .ZN(new_n22467_));
  INV_X1     g22170(.I(new_n22467_), .ZN(new_n22468_));
  OAI21_X1   g22171(.A1(new_n22333_), .A2(new_n22377_), .B(new_n22379_), .ZN(new_n22469_));
  AOI21_X1   g22172(.A1(new_n22361_), .A2(new_n22359_), .B(new_n22357_), .ZN(new_n22470_));
  INV_X1     g22173(.I(new_n22343_), .ZN(new_n22471_));
  AOI21_X1   g22174(.A1(new_n22338_), .A2(new_n22471_), .B(new_n22345_), .ZN(new_n22472_));
  AOI22_X1   g22175(.A1(new_n13472_), .A2(new_n20981_), .B1(\b[34] ), .B2(new_n13884_), .ZN(new_n22473_));
  OAI21_X1   g22176(.A1(new_n22473_), .A2(\a[62] ), .B(new_n13466_), .ZN(new_n22474_));
  NOR2_X1    g22177(.A1(new_n4778_), .A2(new_n22474_), .ZN(new_n22475_));
  NAND2_X1   g22178(.A1(new_n4778_), .A2(new_n22474_), .ZN(new_n22476_));
  INV_X1     g22179(.I(new_n22476_), .ZN(new_n22477_));
  NOR2_X1    g22180(.A1(new_n22477_), .A2(new_n22475_), .ZN(new_n22478_));
  NOR2_X1    g22181(.A1(new_n13476_), .A2(new_n3717_), .ZN(new_n22479_));
  XOR2_X1    g22182(.A1(new_n14736_), .A2(new_n3717_), .Z(new_n22480_));
  NAND2_X1   g22183(.A1(new_n22480_), .A2(\b[33] ), .ZN(new_n22481_));
  XOR2_X1    g22184(.A1(new_n22481_), .A2(new_n22479_), .Z(new_n22482_));
  NOR2_X1    g22185(.A1(new_n22482_), .A2(new_n3354_), .ZN(new_n22483_));
  INV_X1     g22186(.I(new_n22483_), .ZN(new_n22484_));
  NAND2_X1   g22187(.A1(new_n22482_), .A2(new_n3354_), .ZN(new_n22485_));
  AOI21_X1   g22188(.A1(new_n22484_), .A2(new_n22485_), .B(new_n22342_), .ZN(new_n22486_));
  XOR2_X1    g22189(.A1(new_n22482_), .A2(\a[32] ), .Z(new_n22487_));
  NOR2_X1    g22190(.A1(new_n22487_), .A2(new_n22344_), .ZN(new_n22488_));
  NOR2_X1    g22191(.A1(new_n22488_), .A2(new_n22486_), .ZN(new_n22489_));
  NOR2_X1    g22192(.A1(new_n22478_), .A2(new_n22489_), .ZN(new_n22490_));
  INV_X1     g22193(.I(new_n22489_), .ZN(new_n22491_));
  NOR3_X1    g22194(.A1(new_n22477_), .A2(new_n22475_), .A3(new_n22491_), .ZN(new_n22492_));
  NOR2_X1    g22195(.A1(new_n22490_), .A2(new_n22492_), .ZN(new_n22493_));
  NOR2_X1    g22196(.A1(new_n22493_), .A2(new_n22472_), .ZN(new_n22494_));
  INV_X1     g22197(.I(new_n22472_), .ZN(new_n22495_));
  XOR2_X1    g22198(.A1(new_n22478_), .A2(new_n22491_), .Z(new_n22496_));
  NOR2_X1    g22199(.A1(new_n22496_), .A2(new_n22495_), .ZN(new_n22497_));
  NOR2_X1    g22200(.A1(new_n22497_), .A2(new_n22494_), .ZN(new_n22498_));
  AOI22_X1   g22201(.A1(new_n13078_), .A2(\b[37] ), .B1(new_n5915_), .B2(new_n12218_), .ZN(new_n22499_));
  OAI21_X1   g22202(.A1(new_n22499_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22500_));
  XOR2_X1    g22203(.A1(new_n5600_), .A2(new_n22500_), .Z(new_n22501_));
  XNOR2_X1   g22204(.A1(new_n22498_), .A2(new_n22501_), .ZN(new_n22502_));
  NOR2_X1    g22205(.A1(new_n22502_), .A2(new_n22470_), .ZN(new_n22503_));
  INV_X1     g22206(.I(new_n22470_), .ZN(new_n22504_));
  NOR2_X1    g22207(.A1(new_n22498_), .A2(new_n22501_), .ZN(new_n22505_));
  INV_X1     g22208(.I(new_n22505_), .ZN(new_n22506_));
  NAND2_X1   g22209(.A1(new_n22498_), .A2(new_n22501_), .ZN(new_n22507_));
  AOI21_X1   g22210(.A1(new_n22506_), .A2(new_n22507_), .B(new_n22504_), .ZN(new_n22508_));
  NOR2_X1    g22211(.A1(new_n22503_), .A2(new_n22508_), .ZN(new_n22509_));
  INV_X1     g22212(.I(new_n22509_), .ZN(new_n22510_));
  AOI22_X1   g22213(.A1(new_n10969_), .A2(new_n6540_), .B1(new_n11394_), .B2(\b[40] ), .ZN(new_n22511_));
  OAI21_X1   g22214(.A1(new_n22511_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22512_));
  XNOR2_X1   g22215(.A1(new_n6543_), .A2(new_n22512_), .ZN(new_n22513_));
  NAND2_X1   g22216(.A1(new_n22372_), .A2(new_n22368_), .ZN(new_n22514_));
  AOI21_X1   g22217(.A1(new_n22514_), .A2(new_n22371_), .B(new_n22513_), .ZN(new_n22515_));
  INV_X1     g22218(.I(new_n22513_), .ZN(new_n22516_));
  NAND2_X1   g22219(.A1(new_n22514_), .A2(new_n22371_), .ZN(new_n22517_));
  NOR2_X1    g22220(.A1(new_n22517_), .A2(new_n22516_), .ZN(new_n22518_));
  OAI21_X1   g22221(.A1(new_n22518_), .A2(new_n22515_), .B(new_n22510_), .ZN(new_n22519_));
  XOR2_X1    g22222(.A1(new_n22517_), .A2(new_n22513_), .Z(new_n22520_));
  OAI21_X1   g22223(.A1(new_n22510_), .A2(new_n22520_), .B(new_n22519_), .ZN(new_n22521_));
  AOI22_X1   g22224(.A1(new_n11415_), .A2(new_n7866_), .B1(\b[43] ), .B2(new_n10145_), .ZN(new_n22522_));
  OAI21_X1   g22225(.A1(new_n22522_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22523_));
  XNOR2_X1   g22226(.A1(new_n7516_), .A2(new_n22523_), .ZN(new_n22524_));
  XOR2_X1    g22227(.A1(new_n22521_), .A2(new_n22524_), .Z(new_n22525_));
  OR2_X2     g22228(.A1(new_n22521_), .A2(new_n22524_), .Z(new_n22526_));
  NAND2_X1   g22229(.A1(new_n22521_), .A2(new_n22524_), .ZN(new_n22527_));
  AOI21_X1   g22230(.A1(new_n22526_), .A2(new_n22527_), .B(new_n22469_), .ZN(new_n22528_));
  AOI21_X1   g22231(.A1(new_n22469_), .A2(new_n22525_), .B(new_n22528_), .ZN(new_n22529_));
  INV_X1     g22232(.I(new_n22529_), .ZN(new_n22530_));
  OAI22_X1   g22233(.A1(new_n8644_), .A2(new_n8218_), .B1(new_n8563_), .B2(new_n9388_), .ZN(new_n22531_));
  OAI21_X1   g22234(.A1(new_n7870_), .A2(new_n10154_), .B(new_n22531_), .ZN(new_n22532_));
  AOI21_X1   g22235(.A1(new_n22532_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n22533_));
  XOR2_X1    g22236(.A1(new_n8568_), .A2(new_n22533_), .Z(new_n22534_));
  NAND2_X1   g22237(.A1(new_n22381_), .A2(new_n22391_), .ZN(new_n22535_));
  AOI21_X1   g22238(.A1(new_n22535_), .A2(new_n22390_), .B(new_n22534_), .ZN(new_n22536_));
  INV_X1     g22239(.I(new_n22534_), .ZN(new_n22537_));
  NAND2_X1   g22240(.A1(new_n22535_), .A2(new_n22390_), .ZN(new_n22538_));
  NOR2_X1    g22241(.A1(new_n22538_), .A2(new_n22537_), .ZN(new_n22539_));
  OAI21_X1   g22242(.A1(new_n22539_), .A2(new_n22536_), .B(new_n22530_), .ZN(new_n22540_));
  XOR2_X1    g22243(.A1(new_n22538_), .A2(new_n22534_), .Z(new_n22541_));
  OAI21_X1   g22244(.A1(new_n22541_), .A2(new_n22530_), .B(new_n22540_), .ZN(new_n22542_));
  OAI22_X1   g22245(.A1(new_n7619_), .A2(new_n9295_), .B1(new_n10025_), .B2(new_n8309_), .ZN(new_n22543_));
  OAI21_X1   g22246(.A1(new_n8948_), .A2(new_n7947_), .B(new_n22543_), .ZN(new_n22544_));
  AOI21_X1   g22247(.A1(new_n22544_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22545_));
  XNOR2_X1   g22248(.A1(new_n9642_), .A2(new_n22545_), .ZN(new_n22546_));
  NOR2_X1    g22249(.A1(new_n22542_), .A2(new_n22546_), .ZN(new_n22547_));
  NAND2_X1   g22250(.A1(new_n22542_), .A2(new_n22546_), .ZN(new_n22548_));
  INV_X1     g22251(.I(new_n22548_), .ZN(new_n22549_));
  OAI21_X1   g22252(.A1(new_n22549_), .A2(new_n22547_), .B(new_n22468_), .ZN(new_n22550_));
  XOR2_X1    g22253(.A1(new_n22542_), .A2(new_n22546_), .Z(new_n22551_));
  NAND2_X1   g22254(.A1(new_n22551_), .A2(new_n22467_), .ZN(new_n22552_));
  NAND2_X1   g22255(.A1(new_n22552_), .A2(new_n22550_), .ZN(new_n22553_));
  OAI22_X1   g22256(.A1(new_n6644_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n6647_), .ZN(new_n22554_));
  OAI21_X1   g22257(.A1(new_n10031_), .A2(new_n7284_), .B(new_n22554_), .ZN(new_n22555_));
  AOI21_X1   g22258(.A1(new_n22555_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22556_));
  XNOR2_X1   g22259(.A1(new_n10866_), .A2(new_n22556_), .ZN(new_n22557_));
  XOR2_X1    g22260(.A1(new_n22553_), .A2(new_n22557_), .Z(new_n22558_));
  AOI21_X1   g22261(.A1(new_n22552_), .A2(new_n22550_), .B(new_n22557_), .ZN(new_n22559_));
  INV_X1     g22262(.I(new_n22557_), .ZN(new_n22560_));
  NOR2_X1    g22263(.A1(new_n22553_), .A2(new_n22560_), .ZN(new_n22561_));
  OAI21_X1   g22264(.A1(new_n22561_), .A2(new_n22559_), .B(new_n22466_), .ZN(new_n22562_));
  OAI21_X1   g22265(.A1(new_n22558_), .A2(new_n22466_), .B(new_n22562_), .ZN(new_n22563_));
  AOI22_X1   g22266(.A1(new_n5680_), .A2(\b[56] ), .B1(\b[57] ), .B2(new_n5686_), .ZN(new_n22564_));
  AOI21_X1   g22267(.A1(\b[55] ), .A2(new_n6923_), .B(new_n22564_), .ZN(new_n22565_));
  OAI21_X1   g22268(.A1(new_n22565_), .A2(\a[41] ), .B(new_n5680_), .ZN(new_n22566_));
  XOR2_X1    g22269(.A1(new_n12128_), .A2(new_n22566_), .Z(new_n22567_));
  XOR2_X1    g22270(.A1(new_n22563_), .A2(new_n22567_), .Z(new_n22568_));
  NOR2_X1    g22271(.A1(new_n22563_), .A2(new_n22567_), .ZN(new_n22569_));
  INV_X1     g22272(.I(new_n22569_), .ZN(new_n22570_));
  NAND2_X1   g22273(.A1(new_n22563_), .A2(new_n22567_), .ZN(new_n22571_));
  NAND2_X1   g22274(.A1(new_n22570_), .A2(new_n22571_), .ZN(new_n22572_));
  MUX2_X1    g22275(.I0(new_n22572_), .I1(new_n22568_), .S(new_n22465_), .Z(new_n22573_));
  OAI22_X1   g22276(.A1(new_n5420_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n5107_), .ZN(new_n22574_));
  OAI21_X1   g22277(.A1(new_n12542_), .A2(new_n5112_), .B(new_n22574_), .ZN(new_n22575_));
  AOI21_X1   g22278(.A1(new_n22575_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n22576_));
  XNOR2_X1   g22279(.A1(new_n13371_), .A2(new_n22576_), .ZN(new_n22577_));
  INV_X1     g22280(.I(new_n22577_), .ZN(new_n22578_));
  NAND2_X1   g22281(.A1(new_n22421_), .A2(new_n22431_), .ZN(new_n22579_));
  NAND2_X1   g22282(.A1(new_n22579_), .A2(new_n22430_), .ZN(new_n22580_));
  NAND2_X1   g22283(.A1(new_n22580_), .A2(new_n22578_), .ZN(new_n22581_));
  INV_X1     g22284(.I(new_n22581_), .ZN(new_n22582_));
  NOR2_X1    g22285(.A1(new_n22580_), .A2(new_n22578_), .ZN(new_n22583_));
  OAI21_X1   g22286(.A1(new_n22582_), .A2(new_n22583_), .B(new_n22573_), .ZN(new_n22584_));
  XOR2_X1    g22287(.A1(new_n22580_), .A2(new_n22577_), .Z(new_n22585_));
  OR2_X2     g22288(.A1(new_n22585_), .A2(new_n22573_), .Z(new_n22586_));
  NAND2_X1   g22289(.A1(new_n22586_), .A2(new_n22584_), .ZN(new_n22587_));
  XOR2_X1    g22290(.A1(new_n22587_), .A2(new_n22464_), .Z(new_n22588_));
  AND2_X2    g22291(.A1(new_n22587_), .A2(new_n22463_), .Z(new_n22589_));
  NOR2_X1    g22292(.A1(new_n22587_), .A2(new_n22463_), .ZN(new_n22590_));
  OAI21_X1   g22293(.A1(new_n22589_), .A2(new_n22590_), .B(new_n22459_), .ZN(new_n22591_));
  OAI21_X1   g22294(.A1(new_n22459_), .A2(new_n22588_), .B(new_n22591_), .ZN(new_n22592_));
  XNOR2_X1   g22295(.A1(new_n22592_), .A2(new_n22457_), .ZN(new_n22593_));
  AOI21_X1   g22296(.A1(new_n22593_), .A2(new_n22449_), .B(new_n22451_), .ZN(new_n22594_));
  XOR2_X1    g22297(.A1(new_n22309_), .A2(new_n22594_), .Z(\f[96] ));
  NAND2_X1   g22298(.A1(new_n22592_), .A2(new_n22457_), .ZN(new_n22596_));
  NOR2_X1    g22299(.A1(new_n22450_), .A2(new_n22448_), .ZN(new_n22597_));
  AOI21_X1   g22300(.A1(new_n22308_), .A2(new_n22306_), .B(new_n22597_), .ZN(new_n22598_));
  NOR2_X1    g22301(.A1(new_n4318_), .A2(new_n4067_), .ZN(new_n22599_));
  NAND2_X1   g22302(.A1(new_n16148_), .A2(new_n4069_), .ZN(new_n22600_));
  OAI21_X1   g22303(.A1(new_n22599_), .A2(new_n22600_), .B(new_n4062_), .ZN(new_n22601_));
  XNOR2_X1   g22304(.A1(new_n14978_), .A2(new_n22601_), .ZN(new_n22602_));
  OAI21_X1   g22305(.A1(new_n22573_), .A2(new_n22583_), .B(new_n22581_), .ZN(new_n22603_));
  OAI22_X1   g22306(.A1(new_n5993_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n5991_), .ZN(new_n22604_));
  OAI21_X1   g22307(.A1(new_n11744_), .A2(new_n5997_), .B(new_n22604_), .ZN(new_n22605_));
  AOI21_X1   g22308(.A1(new_n22605_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n22606_));
  XNOR2_X1   g22309(.A1(new_n12546_), .A2(new_n22606_), .ZN(new_n22607_));
  NOR2_X1    g22310(.A1(new_n22561_), .A2(new_n22466_), .ZN(new_n22608_));
  AOI21_X1   g22311(.A1(new_n22468_), .A2(new_n22548_), .B(new_n22547_), .ZN(new_n22609_));
  OAI22_X1   g22312(.A1(new_n7619_), .A2(new_n10025_), .B1(new_n10031_), .B2(new_n8309_), .ZN(new_n22610_));
  OAI21_X1   g22313(.A1(new_n9295_), .A2(new_n7947_), .B(new_n22610_), .ZN(new_n22611_));
  AOI21_X1   g22314(.A1(new_n22611_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22612_));
  XNOR2_X1   g22315(.A1(new_n10035_), .A2(new_n22612_), .ZN(new_n22613_));
  INV_X1     g22316(.I(new_n7871_), .ZN(new_n22614_));
  AOI22_X1   g22317(.A1(new_n11415_), .A2(new_n22614_), .B1(\b[44] ), .B2(new_n10145_), .ZN(new_n22615_));
  OAI21_X1   g22318(.A1(new_n22615_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22616_));
  XOR2_X1    g22319(.A1(new_n7874_), .A2(new_n22616_), .Z(new_n22617_));
  INV_X1     g22320(.I(new_n22617_), .ZN(new_n22618_));
  AOI21_X1   g22321(.A1(new_n22504_), .A2(new_n22507_), .B(new_n22505_), .ZN(new_n22619_));
  AOI22_X1   g22322(.A1(new_n13078_), .A2(\b[38] ), .B1(new_n5923_), .B2(new_n12218_), .ZN(new_n22620_));
  OAI21_X1   g22323(.A1(new_n22620_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22621_));
  XNOR2_X1   g22324(.A1(new_n5926_), .A2(new_n22621_), .ZN(new_n22622_));
  NOR2_X1    g22325(.A1(new_n22492_), .A2(new_n22472_), .ZN(new_n22623_));
  NOR2_X1    g22326(.A1(new_n22623_), .A2(new_n22490_), .ZN(new_n22624_));
  OAI22_X1   g22327(.A1(new_n13880_), .A2(new_n5348_), .B1(new_n4500_), .B2(new_n13885_), .ZN(new_n22625_));
  AOI21_X1   g22328(.A1(new_n22625_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n22626_));
  XNOR2_X1   g22329(.A1(new_n5067_), .A2(new_n22626_), .ZN(new_n22627_));
  NAND2_X1   g22330(.A1(new_n22485_), .A2(new_n22344_), .ZN(new_n22628_));
  NAND2_X1   g22331(.A1(new_n22628_), .A2(new_n22484_), .ZN(new_n22629_));
  NOR2_X1    g22332(.A1(new_n13476_), .A2(new_n3989_), .ZN(new_n22630_));
  XOR2_X1    g22333(.A1(new_n14736_), .A2(new_n3989_), .Z(new_n22631_));
  NAND2_X1   g22334(.A1(new_n22631_), .A2(\b[34] ), .ZN(new_n22632_));
  XOR2_X1    g22335(.A1(new_n22632_), .A2(new_n22630_), .Z(new_n22633_));
  INV_X1     g22336(.I(new_n22633_), .ZN(new_n22634_));
  XOR2_X1    g22337(.A1(new_n22629_), .A2(new_n22634_), .Z(new_n22635_));
  INV_X1     g22338(.I(new_n22635_), .ZN(new_n22636_));
  NOR2_X1    g22339(.A1(new_n22629_), .A2(new_n22633_), .ZN(new_n22637_));
  INV_X1     g22340(.I(new_n22637_), .ZN(new_n22638_));
  NAND2_X1   g22341(.A1(new_n22629_), .A2(new_n22633_), .ZN(new_n22639_));
  AOI21_X1   g22342(.A1(new_n22638_), .A2(new_n22639_), .B(new_n22627_), .ZN(new_n22640_));
  AOI21_X1   g22343(.A1(new_n22627_), .A2(new_n22636_), .B(new_n22640_), .ZN(new_n22641_));
  XOR2_X1    g22344(.A1(new_n22641_), .A2(new_n22624_), .Z(new_n22642_));
  INV_X1     g22345(.I(new_n22641_), .ZN(new_n22643_));
  NAND2_X1   g22346(.A1(new_n22643_), .A2(new_n22624_), .ZN(new_n22644_));
  NOR2_X1    g22347(.A1(new_n22643_), .A2(new_n22624_), .ZN(new_n22645_));
  INV_X1     g22348(.I(new_n22645_), .ZN(new_n22646_));
  NAND2_X1   g22349(.A1(new_n22646_), .A2(new_n22644_), .ZN(new_n22647_));
  NAND2_X1   g22350(.A1(new_n22647_), .A2(new_n22622_), .ZN(new_n22648_));
  OAI21_X1   g22351(.A1(new_n22622_), .A2(new_n22642_), .B(new_n22648_), .ZN(new_n22649_));
  AOI22_X1   g22352(.A1(new_n10969_), .A2(new_n7194_), .B1(new_n11394_), .B2(\b[41] ), .ZN(new_n22650_));
  OAI21_X1   g22353(.A1(new_n22650_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22651_));
  XNOR2_X1   g22354(.A1(new_n6851_), .A2(new_n22651_), .ZN(new_n22652_));
  NOR2_X1    g22355(.A1(new_n22649_), .A2(new_n22652_), .ZN(new_n22653_));
  INV_X1     g22356(.I(new_n22653_), .ZN(new_n22654_));
  NAND2_X1   g22357(.A1(new_n22649_), .A2(new_n22652_), .ZN(new_n22655_));
  AOI21_X1   g22358(.A1(new_n22654_), .A2(new_n22655_), .B(new_n22619_), .ZN(new_n22656_));
  INV_X1     g22359(.I(new_n22619_), .ZN(new_n22657_));
  XNOR2_X1   g22360(.A1(new_n22649_), .A2(new_n22652_), .ZN(new_n22658_));
  NOR2_X1    g22361(.A1(new_n22658_), .A2(new_n22657_), .ZN(new_n22659_));
  NOR2_X1    g22362(.A1(new_n22659_), .A2(new_n22656_), .ZN(new_n22660_));
  NOR2_X1    g22363(.A1(new_n22518_), .A2(new_n22510_), .ZN(new_n22661_));
  NOR2_X1    g22364(.A1(new_n22661_), .A2(new_n22515_), .ZN(new_n22662_));
  NOR2_X1    g22365(.A1(new_n22660_), .A2(new_n22662_), .ZN(new_n22663_));
  NAND2_X1   g22366(.A1(new_n22660_), .A2(new_n22662_), .ZN(new_n22664_));
  INV_X1     g22367(.I(new_n22664_), .ZN(new_n22665_));
  OAI21_X1   g22368(.A1(new_n22665_), .A2(new_n22663_), .B(new_n22618_), .ZN(new_n22666_));
  XOR2_X1    g22369(.A1(new_n22660_), .A2(new_n22662_), .Z(new_n22667_));
  NAND2_X1   g22370(.A1(new_n22667_), .A2(new_n22617_), .ZN(new_n22668_));
  NAND2_X1   g22371(.A1(new_n22668_), .A2(new_n22666_), .ZN(new_n22669_));
  NAND2_X1   g22372(.A1(new_n22527_), .A2(new_n22469_), .ZN(new_n22670_));
  NAND2_X1   g22373(.A1(new_n22670_), .A2(new_n22526_), .ZN(new_n22671_));
  INV_X1     g22374(.I(new_n22671_), .ZN(new_n22672_));
  OAI22_X1   g22375(.A1(new_n8644_), .A2(new_n8563_), .B1(new_n8948_), .B2(new_n9388_), .ZN(new_n22673_));
  OAI21_X1   g22376(.A1(new_n8218_), .A2(new_n10154_), .B(new_n22673_), .ZN(new_n22674_));
  AOI21_X1   g22377(.A1(new_n22674_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n22675_));
  XOR2_X1    g22378(.A1(new_n8952_), .A2(new_n22675_), .Z(new_n22676_));
  NOR2_X1    g22379(.A1(new_n22672_), .A2(new_n22676_), .ZN(new_n22677_));
  INV_X1     g22380(.I(new_n22676_), .ZN(new_n22678_));
  NOR2_X1    g22381(.A1(new_n22671_), .A2(new_n22678_), .ZN(new_n22679_));
  OAI21_X1   g22382(.A1(new_n22677_), .A2(new_n22679_), .B(new_n22669_), .ZN(new_n22680_));
  XOR2_X1    g22383(.A1(new_n22671_), .A2(new_n22676_), .Z(new_n22681_));
  OAI21_X1   g22384(.A1(new_n22669_), .A2(new_n22681_), .B(new_n22680_), .ZN(new_n22682_));
  INV_X1     g22385(.I(new_n22682_), .ZN(new_n22683_));
  NOR2_X1    g22386(.A1(new_n22539_), .A2(new_n22530_), .ZN(new_n22684_));
  NOR2_X1    g22387(.A1(new_n22684_), .A2(new_n22536_), .ZN(new_n22685_));
  NOR2_X1    g22388(.A1(new_n22683_), .A2(new_n22685_), .ZN(new_n22686_));
  INV_X1     g22389(.I(new_n22686_), .ZN(new_n22687_));
  NAND2_X1   g22390(.A1(new_n22683_), .A2(new_n22685_), .ZN(new_n22688_));
  AOI21_X1   g22391(.A1(new_n22687_), .A2(new_n22688_), .B(new_n22613_), .ZN(new_n22689_));
  INV_X1     g22392(.I(new_n22613_), .ZN(new_n22690_));
  XOR2_X1    g22393(.A1(new_n22685_), .A2(new_n22682_), .Z(new_n22691_));
  NOR2_X1    g22394(.A1(new_n22691_), .A2(new_n22690_), .ZN(new_n22692_));
  NOR2_X1    g22395(.A1(new_n22692_), .A2(new_n22689_), .ZN(new_n22693_));
  OAI22_X1   g22396(.A1(new_n6644_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n6647_), .ZN(new_n22694_));
  OAI21_X1   g22397(.A1(new_n10477_), .A2(new_n7284_), .B(new_n22694_), .ZN(new_n22695_));
  AOI21_X1   g22398(.A1(new_n22695_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22696_));
  XOR2_X1    g22399(.A1(new_n11298_), .A2(new_n22696_), .Z(new_n22697_));
  XNOR2_X1   g22400(.A1(new_n22693_), .A2(new_n22697_), .ZN(new_n22698_));
  NOR2_X1    g22401(.A1(new_n22698_), .A2(new_n22609_), .ZN(new_n22699_));
  INV_X1     g22402(.I(new_n22609_), .ZN(new_n22700_));
  NOR2_X1    g22403(.A1(new_n22693_), .A2(new_n22697_), .ZN(new_n22701_));
  INV_X1     g22404(.I(new_n22701_), .ZN(new_n22702_));
  NAND2_X1   g22405(.A1(new_n22693_), .A2(new_n22697_), .ZN(new_n22703_));
  AOI21_X1   g22406(.A1(new_n22702_), .A2(new_n22703_), .B(new_n22700_), .ZN(new_n22704_));
  NOR2_X1    g22407(.A1(new_n22699_), .A2(new_n22704_), .ZN(new_n22705_));
  NOR3_X1    g22408(.A1(new_n22705_), .A2(new_n22559_), .A3(new_n22608_), .ZN(new_n22706_));
  NOR2_X1    g22409(.A1(new_n22608_), .A2(new_n22559_), .ZN(new_n22707_));
  INV_X1     g22410(.I(new_n22705_), .ZN(new_n22708_));
  NOR2_X1    g22411(.A1(new_n22708_), .A2(new_n22707_), .ZN(new_n22709_));
  NOR2_X1    g22412(.A1(new_n22709_), .A2(new_n22706_), .ZN(new_n22710_));
  NOR2_X1    g22413(.A1(new_n22710_), .A2(new_n22607_), .ZN(new_n22711_));
  INV_X1     g22414(.I(new_n22607_), .ZN(new_n22712_));
  XOR2_X1    g22415(.A1(new_n22705_), .A2(new_n22707_), .Z(new_n22713_));
  NOR2_X1    g22416(.A1(new_n22713_), .A2(new_n22712_), .ZN(new_n22714_));
  NOR2_X1    g22417(.A1(new_n22711_), .A2(new_n22714_), .ZN(new_n22715_));
  NAND2_X1   g22418(.A1(new_n22571_), .A2(new_n22465_), .ZN(new_n22716_));
  NAND2_X1   g22419(.A1(new_n22716_), .A2(new_n22570_), .ZN(new_n22717_));
  OAI22_X1   g22420(.A1(new_n5420_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n5107_), .ZN(new_n22718_));
  OAI21_X1   g22421(.A1(new_n12970_), .A2(new_n5112_), .B(new_n22718_), .ZN(new_n22719_));
  AOI21_X1   g22422(.A1(new_n22719_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n22720_));
  XOR2_X1    g22423(.A1(new_n13784_), .A2(new_n22720_), .Z(new_n22721_));
  XOR2_X1    g22424(.A1(new_n22717_), .A2(new_n22721_), .Z(new_n22722_));
  NOR2_X1    g22425(.A1(new_n22722_), .A2(new_n22715_), .ZN(new_n22723_));
  INV_X1     g22426(.I(new_n22715_), .ZN(new_n22724_));
  INV_X1     g22427(.I(new_n22717_), .ZN(new_n22725_));
  NOR2_X1    g22428(.A1(new_n22725_), .A2(new_n22721_), .ZN(new_n22726_));
  INV_X1     g22429(.I(new_n22726_), .ZN(new_n22727_));
  NAND2_X1   g22430(.A1(new_n22725_), .A2(new_n22721_), .ZN(new_n22728_));
  AOI21_X1   g22431(.A1(new_n22727_), .A2(new_n22728_), .B(new_n22724_), .ZN(new_n22729_));
  NOR2_X1    g22432(.A1(new_n22729_), .A2(new_n22723_), .ZN(new_n22730_));
  NOR2_X1    g22433(.A1(new_n22730_), .A2(new_n22603_), .ZN(new_n22731_));
  INV_X1     g22434(.I(new_n22603_), .ZN(new_n22732_));
  INV_X1     g22435(.I(new_n22730_), .ZN(new_n22733_));
  NOR2_X1    g22436(.A1(new_n22733_), .A2(new_n22732_), .ZN(new_n22734_));
  NOR2_X1    g22437(.A1(new_n22734_), .A2(new_n22731_), .ZN(new_n22735_));
  NOR2_X1    g22438(.A1(new_n22735_), .A2(new_n22602_), .ZN(new_n22736_));
  INV_X1     g22439(.I(new_n22602_), .ZN(new_n22737_));
  XOR2_X1    g22440(.A1(new_n22730_), .A2(new_n22732_), .Z(new_n22738_));
  NOR2_X1    g22441(.A1(new_n22738_), .A2(new_n22737_), .ZN(new_n22739_));
  NOR2_X1    g22442(.A1(new_n22736_), .A2(new_n22739_), .ZN(new_n22740_));
  NOR2_X1    g22443(.A1(new_n22589_), .A2(new_n22459_), .ZN(new_n22741_));
  NOR2_X1    g22444(.A1(new_n22741_), .A2(new_n22590_), .ZN(new_n22742_));
  NOR2_X1    g22445(.A1(new_n22742_), .A2(new_n22740_), .ZN(new_n22743_));
  XNOR2_X1   g22446(.A1(new_n22598_), .A2(new_n22743_), .ZN(new_n22744_));
  XOR2_X1    g22447(.A1(new_n22744_), .A2(new_n22596_), .Z(\f[97] ));
  INV_X1     g22448(.I(new_n22307_), .ZN(new_n22746_));
  NOR3_X1    g22449(.A1(new_n22138_), .A2(new_n22140_), .A3(new_n22746_), .ZN(new_n22747_));
  INV_X1     g22450(.I(new_n22597_), .ZN(new_n22748_));
  OAI21_X1   g22451(.A1(new_n22747_), .A2(new_n22305_), .B(new_n22748_), .ZN(new_n22749_));
  NOR2_X1    g22452(.A1(new_n22596_), .A2(new_n22740_), .ZN(new_n22750_));
  INV_X1     g22453(.I(new_n22750_), .ZN(new_n22751_));
  AOI21_X1   g22454(.A1(new_n22596_), .A2(new_n22740_), .B(new_n22742_), .ZN(new_n22752_));
  INV_X1     g22455(.I(new_n22752_), .ZN(new_n22753_));
  OAI21_X1   g22456(.A1(new_n22749_), .A2(new_n22753_), .B(new_n22751_), .ZN(new_n22754_));
  INV_X1     g22457(.I(new_n22731_), .ZN(new_n22755_));
  AOI21_X1   g22458(.A1(new_n22737_), .A2(new_n22755_), .B(new_n22734_), .ZN(new_n22756_));
  OAI22_X1   g22459(.A1(new_n5420_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n5107_), .ZN(new_n22757_));
  OAI21_X1   g22460(.A1(new_n13367_), .A2(new_n5112_), .B(new_n22757_), .ZN(new_n22758_));
  AOI21_X1   g22461(.A1(new_n22758_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n22759_));
  XOR2_X1    g22462(.A1(new_n14213_), .A2(new_n22759_), .Z(new_n22760_));
  INV_X1     g22463(.I(new_n22760_), .ZN(new_n22761_));
  OAI22_X1   g22464(.A1(new_n6644_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n6647_), .ZN(new_n22762_));
  OAI21_X1   g22465(.A1(new_n10862_), .A2(new_n7284_), .B(new_n22762_), .ZN(new_n22763_));
  AOI21_X1   g22466(.A1(new_n22763_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22764_));
  XNOR2_X1   g22467(.A1(new_n11748_), .A2(new_n22764_), .ZN(new_n22765_));
  INV_X1     g22468(.I(new_n22765_), .ZN(new_n22766_));
  AOI21_X1   g22469(.A1(new_n22690_), .A2(new_n22688_), .B(new_n22686_), .ZN(new_n22767_));
  INV_X1     g22470(.I(new_n22767_), .ZN(new_n22768_));
  OAI22_X1   g22471(.A1(new_n7619_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n8309_), .ZN(new_n22769_));
  OAI21_X1   g22472(.A1(new_n10025_), .A2(new_n7947_), .B(new_n22769_), .ZN(new_n22770_));
  AOI21_X1   g22473(.A1(new_n22770_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22771_));
  XOR2_X1    g22474(.A1(new_n10476_), .A2(new_n22771_), .Z(new_n22772_));
  AOI22_X1   g22475(.A1(new_n8631_), .A2(\b[49] ), .B1(\b[50] ), .B2(new_n9382_), .ZN(new_n22773_));
  AOI21_X1   g22476(.A1(\b[48] ), .A2(new_n9731_), .B(new_n22773_), .ZN(new_n22774_));
  OAI21_X1   g22477(.A1(new_n22774_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n22775_));
  XOR2_X1    g22478(.A1(new_n9299_), .A2(new_n22775_), .Z(new_n22776_));
  INV_X1     g22479(.I(new_n22776_), .ZN(new_n22777_));
  AOI22_X1   g22480(.A1(new_n10969_), .A2(new_n22330_), .B1(new_n11394_), .B2(\b[42] ), .ZN(new_n22778_));
  OAI21_X1   g22481(.A1(new_n22778_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22779_));
  XOR2_X1    g22482(.A1(new_n7202_), .A2(new_n22779_), .Z(new_n22780_));
  INV_X1     g22483(.I(new_n22780_), .ZN(new_n22781_));
  INV_X1     g22484(.I(new_n22622_), .ZN(new_n22782_));
  AOI21_X1   g22485(.A1(new_n22782_), .A2(new_n22644_), .B(new_n22645_), .ZN(new_n22783_));
  NAND2_X1   g22486(.A1(new_n22627_), .A2(new_n22638_), .ZN(new_n22784_));
  NAND2_X1   g22487(.A1(new_n22784_), .A2(new_n22639_), .ZN(new_n22785_));
  NOR2_X1    g22488(.A1(new_n13476_), .A2(new_n4253_), .ZN(new_n22786_));
  XOR2_X1    g22489(.A1(new_n14736_), .A2(new_n4253_), .Z(new_n22787_));
  NAND2_X1   g22490(.A1(new_n22787_), .A2(\b[35] ), .ZN(new_n22788_));
  XOR2_X1    g22491(.A1(new_n22788_), .A2(new_n22786_), .Z(new_n22789_));
  NOR2_X1    g22492(.A1(new_n22634_), .A2(new_n22789_), .ZN(new_n22790_));
  INV_X1     g22493(.I(new_n22789_), .ZN(new_n22791_));
  NOR2_X1    g22494(.A1(new_n22791_), .A2(new_n22633_), .ZN(new_n22792_));
  NOR2_X1    g22495(.A1(new_n22790_), .A2(new_n22792_), .ZN(new_n22793_));
  INV_X1     g22496(.I(new_n22793_), .ZN(new_n22794_));
  XOR2_X1    g22497(.A1(new_n22633_), .A2(new_n22789_), .Z(new_n22795_));
  NOR2_X1    g22498(.A1(new_n22785_), .A2(new_n22795_), .ZN(new_n22796_));
  AOI21_X1   g22499(.A1(new_n22785_), .A2(new_n22794_), .B(new_n22796_), .ZN(new_n22797_));
  AOI22_X1   g22500(.A1(new_n13078_), .A2(\b[39] ), .B1(new_n6532_), .B2(new_n12218_), .ZN(new_n22798_));
  OAI21_X1   g22501(.A1(new_n22798_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22799_));
  XNOR2_X1   g22502(.A1(new_n6233_), .A2(new_n22799_), .ZN(new_n22800_));
  OAI22_X1   g22503(.A1(new_n13880_), .A2(new_n5354_), .B1(new_n4774_), .B2(new_n13885_), .ZN(new_n22801_));
  AOI21_X1   g22504(.A1(new_n22801_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n22802_));
  XNOR2_X1   g22505(.A1(new_n5357_), .A2(new_n22802_), .ZN(new_n22803_));
  NOR2_X1    g22506(.A1(new_n22800_), .A2(new_n22803_), .ZN(new_n22804_));
  INV_X1     g22507(.I(new_n22804_), .ZN(new_n22805_));
  NAND2_X1   g22508(.A1(new_n22800_), .A2(new_n22803_), .ZN(new_n22806_));
  AOI21_X1   g22509(.A1(new_n22805_), .A2(new_n22806_), .B(new_n22797_), .ZN(new_n22807_));
  INV_X1     g22510(.I(new_n22797_), .ZN(new_n22808_));
  XNOR2_X1   g22511(.A1(new_n22800_), .A2(new_n22803_), .ZN(new_n22809_));
  NOR2_X1    g22512(.A1(new_n22809_), .A2(new_n22808_), .ZN(new_n22810_));
  NOR2_X1    g22513(.A1(new_n22810_), .A2(new_n22807_), .ZN(new_n22811_));
  XNOR2_X1   g22514(.A1(new_n22811_), .A2(new_n22783_), .ZN(new_n22812_));
  INV_X1     g22515(.I(new_n22812_), .ZN(new_n22813_));
  NOR2_X1    g22516(.A1(new_n22811_), .A2(new_n22783_), .ZN(new_n22814_));
  INV_X1     g22517(.I(new_n22814_), .ZN(new_n22815_));
  NAND2_X1   g22518(.A1(new_n22811_), .A2(new_n22783_), .ZN(new_n22816_));
  AOI21_X1   g22519(.A1(new_n22815_), .A2(new_n22816_), .B(new_n22781_), .ZN(new_n22817_));
  AOI21_X1   g22520(.A1(new_n22813_), .A2(new_n22781_), .B(new_n22817_), .ZN(new_n22818_));
  AOI22_X1   g22521(.A1(new_n11415_), .A2(new_n8557_), .B1(\b[45] ), .B2(new_n10145_), .ZN(new_n22819_));
  OAI21_X1   g22522(.A1(new_n22819_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22820_));
  XNOR2_X1   g22523(.A1(new_n8217_), .A2(new_n22820_), .ZN(new_n22821_));
  AOI21_X1   g22524(.A1(new_n22657_), .A2(new_n22655_), .B(new_n22653_), .ZN(new_n22822_));
  XNOR2_X1   g22525(.A1(new_n22822_), .A2(new_n22821_), .ZN(new_n22823_));
  NOR2_X1    g22526(.A1(new_n22823_), .A2(new_n22818_), .ZN(new_n22824_));
  NOR2_X1    g22527(.A1(new_n22822_), .A2(new_n22821_), .ZN(new_n22825_));
  INV_X1     g22528(.I(new_n22825_), .ZN(new_n22826_));
  NAND2_X1   g22529(.A1(new_n22822_), .A2(new_n22821_), .ZN(new_n22827_));
  NAND2_X1   g22530(.A1(new_n22826_), .A2(new_n22827_), .ZN(new_n22828_));
  AOI21_X1   g22531(.A1(new_n22818_), .A2(new_n22828_), .B(new_n22824_), .ZN(new_n22829_));
  AOI21_X1   g22532(.A1(new_n22618_), .A2(new_n22664_), .B(new_n22663_), .ZN(new_n22830_));
  XOR2_X1    g22533(.A1(new_n22829_), .A2(new_n22830_), .Z(new_n22831_));
  NOR2_X1    g22534(.A1(new_n22829_), .A2(new_n22830_), .ZN(new_n22832_));
  INV_X1     g22535(.I(new_n22832_), .ZN(new_n22833_));
  NAND2_X1   g22536(.A1(new_n22829_), .A2(new_n22830_), .ZN(new_n22834_));
  AOI21_X1   g22537(.A1(new_n22833_), .A2(new_n22834_), .B(new_n22777_), .ZN(new_n22835_));
  AOI21_X1   g22538(.A1(new_n22777_), .A2(new_n22831_), .B(new_n22835_), .ZN(new_n22836_));
  INV_X1     g22539(.I(new_n22669_), .ZN(new_n22837_));
  INV_X1     g22540(.I(new_n22677_), .ZN(new_n22838_));
  OAI21_X1   g22541(.A1(new_n22837_), .A2(new_n22679_), .B(new_n22838_), .ZN(new_n22839_));
  XNOR2_X1   g22542(.A1(new_n22836_), .A2(new_n22839_), .ZN(new_n22840_));
  NOR2_X1    g22543(.A1(new_n22840_), .A2(new_n22772_), .ZN(new_n22841_));
  NAND2_X1   g22544(.A1(new_n22836_), .A2(new_n22839_), .ZN(new_n22842_));
  NOR2_X1    g22545(.A1(new_n22836_), .A2(new_n22839_), .ZN(new_n22843_));
  INV_X1     g22546(.I(new_n22843_), .ZN(new_n22844_));
  NAND2_X1   g22547(.A1(new_n22844_), .A2(new_n22842_), .ZN(new_n22845_));
  AOI21_X1   g22548(.A1(new_n22772_), .A2(new_n22845_), .B(new_n22841_), .ZN(new_n22846_));
  XOR2_X1    g22549(.A1(new_n22846_), .A2(new_n22768_), .Z(new_n22847_));
  NAND2_X1   g22550(.A1(new_n22847_), .A2(new_n22766_), .ZN(new_n22848_));
  NOR2_X1    g22551(.A1(new_n22846_), .A2(new_n22768_), .ZN(new_n22849_));
  NAND2_X1   g22552(.A1(new_n22846_), .A2(new_n22768_), .ZN(new_n22850_));
  INV_X1     g22553(.I(new_n22850_), .ZN(new_n22851_));
  OAI21_X1   g22554(.A1(new_n22851_), .A2(new_n22849_), .B(new_n22765_), .ZN(new_n22852_));
  NAND2_X1   g22555(.A1(new_n22848_), .A2(new_n22852_), .ZN(new_n22853_));
  OAI22_X1   g22556(.A1(new_n5993_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n5991_), .ZN(new_n22854_));
  OAI21_X1   g22557(.A1(new_n12536_), .A2(new_n5997_), .B(new_n22854_), .ZN(new_n22855_));
  AOI21_X1   g22558(.A1(new_n22855_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n22856_));
  XOR2_X1    g22559(.A1(new_n12969_), .A2(new_n22856_), .Z(new_n22857_));
  AOI21_X1   g22560(.A1(new_n22700_), .A2(new_n22703_), .B(new_n22701_), .ZN(new_n22858_));
  XOR2_X1    g22561(.A1(new_n22858_), .A2(new_n22857_), .Z(new_n22859_));
  NOR2_X1    g22562(.A1(new_n22858_), .A2(new_n22857_), .ZN(new_n22860_));
  INV_X1     g22563(.I(new_n22860_), .ZN(new_n22861_));
  NAND2_X1   g22564(.A1(new_n22858_), .A2(new_n22857_), .ZN(new_n22862_));
  AOI21_X1   g22565(.A1(new_n22861_), .A2(new_n22862_), .B(new_n22853_), .ZN(new_n22863_));
  AOI21_X1   g22566(.A1(new_n22853_), .A2(new_n22859_), .B(new_n22863_), .ZN(new_n22864_));
  NOR2_X1    g22567(.A1(new_n22706_), .A2(new_n22607_), .ZN(new_n22865_));
  NOR2_X1    g22568(.A1(new_n22865_), .A2(new_n22709_), .ZN(new_n22866_));
  NOR2_X1    g22569(.A1(new_n22866_), .A2(new_n22864_), .ZN(new_n22867_));
  NAND2_X1   g22570(.A1(new_n22866_), .A2(new_n22864_), .ZN(new_n22868_));
  INV_X1     g22571(.I(new_n22868_), .ZN(new_n22869_));
  OAI21_X1   g22572(.A1(new_n22869_), .A2(new_n22867_), .B(new_n22761_), .ZN(new_n22870_));
  XNOR2_X1   g22573(.A1(new_n22866_), .A2(new_n22864_), .ZN(new_n22871_));
  OAI21_X1   g22574(.A1(new_n22761_), .A2(new_n22871_), .B(new_n22870_), .ZN(new_n22872_));
  OAI21_X1   g22575(.A1(new_n4072_), .A2(new_n4318_), .B(new_n16487_), .ZN(new_n22873_));
  NAND2_X1   g22576(.A1(new_n22724_), .A2(new_n22728_), .ZN(new_n22874_));
  NAND2_X1   g22577(.A1(new_n22874_), .A2(new_n22727_), .ZN(new_n22875_));
  XNOR2_X1   g22578(.A1(new_n22875_), .A2(new_n22873_), .ZN(new_n22876_));
  XOR2_X1    g22579(.A1(new_n22876_), .A2(new_n22872_), .Z(new_n22877_));
  NOR2_X1    g22580(.A1(new_n22877_), .A2(\a[35] ), .ZN(new_n22878_));
  NAND2_X1   g22581(.A1(new_n22877_), .A2(\a[35] ), .ZN(new_n22879_));
  INV_X1     g22582(.I(new_n22879_), .ZN(new_n22880_));
  NOR2_X1    g22583(.A1(new_n22880_), .A2(new_n22878_), .ZN(new_n22881_));
  XOR2_X1    g22584(.A1(new_n22881_), .A2(new_n22756_), .Z(new_n22882_));
  NAND2_X1   g22585(.A1(new_n22754_), .A2(new_n22882_), .ZN(new_n22883_));
  AOI21_X1   g22586(.A1(new_n22598_), .A2(new_n22752_), .B(new_n22750_), .ZN(new_n22884_));
  INV_X1     g22587(.I(new_n22756_), .ZN(new_n22885_));
  INV_X1     g22588(.I(new_n22881_), .ZN(new_n22886_));
  NAND2_X1   g22589(.A1(new_n22886_), .A2(new_n22885_), .ZN(new_n22887_));
  NAND2_X1   g22590(.A1(new_n22881_), .A2(new_n22756_), .ZN(new_n22888_));
  NAND2_X1   g22591(.A1(new_n22887_), .A2(new_n22888_), .ZN(new_n22889_));
  NAND2_X1   g22592(.A1(new_n22884_), .A2(new_n22889_), .ZN(new_n22890_));
  NAND2_X1   g22593(.A1(new_n22883_), .A2(new_n22890_), .ZN(\f[98] ));
  OAI22_X1   g22594(.A1(new_n5420_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n5107_), .ZN(new_n22892_));
  OAI21_X1   g22595(.A1(new_n13785_), .A2(new_n5112_), .B(new_n22892_), .ZN(new_n22893_));
  AOI21_X1   g22596(.A1(new_n22893_), .A2(new_n4860_), .B(new_n5420_), .ZN(new_n22894_));
  XNOR2_X1   g22597(.A1(new_n14599_), .A2(new_n22894_), .ZN(new_n22895_));
  NOR2_X1    g22598(.A1(new_n22869_), .A2(new_n22760_), .ZN(new_n22896_));
  NOR2_X1    g22599(.A1(new_n22896_), .A2(new_n22867_), .ZN(new_n22897_));
  OAI21_X1   g22600(.A1(new_n22765_), .A2(new_n22849_), .B(new_n22850_), .ZN(new_n22898_));
  OAI21_X1   g22601(.A1(new_n22772_), .A2(new_n22843_), .B(new_n22842_), .ZN(new_n22899_));
  INV_X1     g22602(.I(new_n22899_), .ZN(new_n22900_));
  OAI22_X1   g22603(.A1(new_n7619_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n8309_), .ZN(new_n22901_));
  OAI21_X1   g22604(.A1(new_n10031_), .A2(new_n7947_), .B(new_n22901_), .ZN(new_n22902_));
  AOI21_X1   g22605(.A1(new_n22902_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n22903_));
  XNOR2_X1   g22606(.A1(new_n10866_), .A2(new_n22903_), .ZN(new_n22904_));
  AOI21_X1   g22607(.A1(new_n22777_), .A2(new_n22834_), .B(new_n22832_), .ZN(new_n22905_));
  AOI21_X1   g22608(.A1(new_n22781_), .A2(new_n22816_), .B(new_n22814_), .ZN(new_n22906_));
  INV_X1     g22609(.I(new_n22790_), .ZN(new_n22907_));
  AOI21_X1   g22610(.A1(new_n22785_), .A2(new_n22907_), .B(new_n22792_), .ZN(new_n22908_));
  OAI22_X1   g22611(.A1(new_n13880_), .A2(new_n5914_), .B1(new_n5068_), .B2(new_n13885_), .ZN(new_n22909_));
  AOI21_X1   g22612(.A1(new_n22909_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n22910_));
  XNOR2_X1   g22613(.A1(new_n5600_), .A2(new_n22910_), .ZN(new_n22911_));
  NOR2_X1    g22614(.A1(new_n13476_), .A2(new_n4500_), .ZN(new_n22912_));
  XOR2_X1    g22615(.A1(new_n14736_), .A2(new_n4500_), .Z(new_n22913_));
  NAND2_X1   g22616(.A1(new_n22913_), .A2(\b[36] ), .ZN(new_n22914_));
  XOR2_X1    g22617(.A1(new_n22914_), .A2(new_n22912_), .Z(new_n22915_));
  XOR2_X1    g22618(.A1(new_n22915_), .A2(\a[35] ), .Z(new_n22916_));
  NOR2_X1    g22619(.A1(new_n22916_), .A2(new_n22789_), .ZN(new_n22917_));
  NOR2_X1    g22620(.A1(new_n22915_), .A2(new_n4069_), .ZN(new_n22918_));
  INV_X1     g22621(.I(new_n22918_), .ZN(new_n22919_));
  NAND2_X1   g22622(.A1(new_n22915_), .A2(new_n4069_), .ZN(new_n22920_));
  AOI21_X1   g22623(.A1(new_n22919_), .A2(new_n22920_), .B(new_n22791_), .ZN(new_n22921_));
  NOR2_X1    g22624(.A1(new_n22917_), .A2(new_n22921_), .ZN(new_n22922_));
  XOR2_X1    g22625(.A1(new_n22911_), .A2(new_n22922_), .Z(new_n22923_));
  NOR2_X1    g22626(.A1(new_n22923_), .A2(new_n22908_), .ZN(new_n22924_));
  INV_X1     g22627(.I(new_n22911_), .ZN(new_n22925_));
  NOR2_X1    g22628(.A1(new_n22925_), .A2(new_n22922_), .ZN(new_n22926_));
  INV_X1     g22629(.I(new_n22926_), .ZN(new_n22927_));
  NAND2_X1   g22630(.A1(new_n22925_), .A2(new_n22922_), .ZN(new_n22928_));
  NAND2_X1   g22631(.A1(new_n22927_), .A2(new_n22928_), .ZN(new_n22929_));
  AOI21_X1   g22632(.A1(new_n22908_), .A2(new_n22929_), .B(new_n22924_), .ZN(new_n22930_));
  AOI22_X1   g22633(.A1(new_n13078_), .A2(\b[40] ), .B1(new_n6540_), .B2(new_n12218_), .ZN(new_n22931_));
  OAI21_X1   g22634(.A1(new_n22931_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n22932_));
  XNOR2_X1   g22635(.A1(new_n6543_), .A2(new_n22932_), .ZN(new_n22933_));
  NAND2_X1   g22636(.A1(new_n22806_), .A2(new_n22808_), .ZN(new_n22934_));
  NAND2_X1   g22637(.A1(new_n22934_), .A2(new_n22805_), .ZN(new_n22935_));
  XOR2_X1    g22638(.A1(new_n22933_), .A2(new_n22935_), .Z(new_n22936_));
  NOR2_X1    g22639(.A1(new_n22936_), .A2(new_n22930_), .ZN(new_n22937_));
  INV_X1     g22640(.I(new_n22935_), .ZN(new_n22938_));
  NOR2_X1    g22641(.A1(new_n22938_), .A2(new_n22933_), .ZN(new_n22939_));
  INV_X1     g22642(.I(new_n22939_), .ZN(new_n22940_));
  NAND2_X1   g22643(.A1(new_n22938_), .A2(new_n22933_), .ZN(new_n22941_));
  NAND2_X1   g22644(.A1(new_n22940_), .A2(new_n22941_), .ZN(new_n22942_));
  AOI21_X1   g22645(.A1(new_n22930_), .A2(new_n22942_), .B(new_n22937_), .ZN(new_n22943_));
  AOI22_X1   g22646(.A1(new_n10969_), .A2(new_n7866_), .B1(new_n11394_), .B2(\b[43] ), .ZN(new_n22944_));
  OAI21_X1   g22647(.A1(new_n22944_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n22945_));
  XNOR2_X1   g22648(.A1(new_n7516_), .A2(new_n22945_), .ZN(new_n22946_));
  XNOR2_X1   g22649(.A1(new_n22943_), .A2(new_n22946_), .ZN(new_n22947_));
  NOR2_X1    g22650(.A1(new_n22947_), .A2(new_n22906_), .ZN(new_n22948_));
  INV_X1     g22651(.I(new_n22906_), .ZN(new_n22949_));
  NOR2_X1    g22652(.A1(new_n22943_), .A2(new_n22946_), .ZN(new_n22950_));
  INV_X1     g22653(.I(new_n22950_), .ZN(new_n22951_));
  NAND2_X1   g22654(.A1(new_n22943_), .A2(new_n22946_), .ZN(new_n22952_));
  AOI21_X1   g22655(.A1(new_n22951_), .A2(new_n22952_), .B(new_n22949_), .ZN(new_n22953_));
  NOR2_X1    g22656(.A1(new_n22948_), .A2(new_n22953_), .ZN(new_n22954_));
  INV_X1     g22657(.I(new_n22954_), .ZN(new_n22955_));
  AOI22_X1   g22658(.A1(new_n11415_), .A2(new_n8565_), .B1(\b[46] ), .B2(new_n10145_), .ZN(new_n22956_));
  OAI21_X1   g22659(.A1(new_n22956_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n22957_));
  XNOR2_X1   g22660(.A1(new_n8568_), .A2(new_n22957_), .ZN(new_n22958_));
  NAND2_X1   g22661(.A1(new_n22818_), .A2(new_n22827_), .ZN(new_n22959_));
  NAND2_X1   g22662(.A1(new_n22959_), .A2(new_n22826_), .ZN(new_n22960_));
  INV_X1     g22663(.I(new_n22960_), .ZN(new_n22961_));
  NOR2_X1    g22664(.A1(new_n22961_), .A2(new_n22958_), .ZN(new_n22962_));
  NAND2_X1   g22665(.A1(new_n22961_), .A2(new_n22958_), .ZN(new_n22963_));
  INV_X1     g22666(.I(new_n22963_), .ZN(new_n22964_));
  OAI21_X1   g22667(.A1(new_n22962_), .A2(new_n22964_), .B(new_n22955_), .ZN(new_n22965_));
  XOR2_X1    g22668(.A1(new_n22960_), .A2(new_n22958_), .Z(new_n22966_));
  OAI21_X1   g22669(.A1(new_n22955_), .A2(new_n22966_), .B(new_n22965_), .ZN(new_n22967_));
  AOI22_X1   g22670(.A1(new_n8631_), .A2(\b[50] ), .B1(\b[51] ), .B2(new_n9382_), .ZN(new_n22968_));
  AOI21_X1   g22671(.A1(\b[49] ), .A2(new_n9731_), .B(new_n22968_), .ZN(new_n22969_));
  OAI21_X1   g22672(.A1(new_n22969_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n22970_));
  XOR2_X1    g22673(.A1(new_n9642_), .A2(new_n22970_), .Z(new_n22971_));
  XNOR2_X1   g22674(.A1(new_n22967_), .A2(new_n22971_), .ZN(new_n22972_));
  NOR2_X1    g22675(.A1(new_n22972_), .A2(new_n22905_), .ZN(new_n22973_));
  INV_X1     g22676(.I(new_n22905_), .ZN(new_n22974_));
  NOR2_X1    g22677(.A1(new_n22967_), .A2(new_n22971_), .ZN(new_n22975_));
  INV_X1     g22678(.I(new_n22975_), .ZN(new_n22976_));
  NAND2_X1   g22679(.A1(new_n22967_), .A2(new_n22971_), .ZN(new_n22977_));
  AOI21_X1   g22680(.A1(new_n22976_), .A2(new_n22977_), .B(new_n22974_), .ZN(new_n22978_));
  NOR2_X1    g22681(.A1(new_n22973_), .A2(new_n22978_), .ZN(new_n22979_));
  XOR2_X1    g22682(.A1(new_n22979_), .A2(new_n22904_), .Z(new_n22980_));
  INV_X1     g22683(.I(new_n22904_), .ZN(new_n22981_));
  NOR2_X1    g22684(.A1(new_n22979_), .A2(new_n22981_), .ZN(new_n22982_));
  NAND2_X1   g22685(.A1(new_n22979_), .A2(new_n22981_), .ZN(new_n22983_));
  INV_X1     g22686(.I(new_n22983_), .ZN(new_n22984_));
  OAI21_X1   g22687(.A1(new_n22984_), .A2(new_n22982_), .B(new_n22900_), .ZN(new_n22985_));
  OAI21_X1   g22688(.A1(new_n22900_), .A2(new_n22980_), .B(new_n22985_), .ZN(new_n22986_));
  OAI22_X1   g22689(.A1(new_n6644_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n6647_), .ZN(new_n22987_));
  OAI21_X1   g22690(.A1(new_n11738_), .A2(new_n7284_), .B(new_n22987_), .ZN(new_n22988_));
  AOI21_X1   g22691(.A1(new_n22988_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n22989_));
  XNOR2_X1   g22692(.A1(new_n12128_), .A2(new_n22989_), .ZN(new_n22990_));
  XNOR2_X1   g22693(.A1(new_n22986_), .A2(new_n22990_), .ZN(new_n22991_));
  INV_X1     g22694(.I(new_n22991_), .ZN(new_n22992_));
  NOR2_X1    g22695(.A1(new_n22986_), .A2(new_n22990_), .ZN(new_n22993_));
  INV_X1     g22696(.I(new_n22993_), .ZN(new_n22994_));
  NAND2_X1   g22697(.A1(new_n22986_), .A2(new_n22990_), .ZN(new_n22995_));
  AOI21_X1   g22698(.A1(new_n22994_), .A2(new_n22995_), .B(new_n22898_), .ZN(new_n22996_));
  AOI21_X1   g22699(.A1(new_n22992_), .A2(new_n22898_), .B(new_n22996_), .ZN(new_n22997_));
  OAI22_X1   g22700(.A1(new_n5993_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n5991_), .ZN(new_n22998_));
  OAI21_X1   g22701(.A1(new_n12542_), .A2(new_n5997_), .B(new_n22998_), .ZN(new_n22999_));
  AOI21_X1   g22702(.A1(new_n22999_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n23000_));
  XNOR2_X1   g22703(.A1(new_n13371_), .A2(new_n23000_), .ZN(new_n23001_));
  NAND3_X1   g22704(.A1(new_n22862_), .A2(new_n22848_), .A3(new_n22852_), .ZN(new_n23002_));
  AOI21_X1   g22705(.A1(new_n23002_), .A2(new_n22861_), .B(new_n23001_), .ZN(new_n23003_));
  INV_X1     g22706(.I(new_n23003_), .ZN(new_n23004_));
  INV_X1     g22707(.I(new_n23001_), .ZN(new_n23005_));
  NAND2_X1   g22708(.A1(new_n23002_), .A2(new_n22861_), .ZN(new_n23006_));
  NOR2_X1    g22709(.A1(new_n23006_), .A2(new_n23005_), .ZN(new_n23007_));
  INV_X1     g22710(.I(new_n23007_), .ZN(new_n23008_));
  AOI21_X1   g22711(.A1(new_n23008_), .A2(new_n23004_), .B(new_n22997_), .ZN(new_n23009_));
  XOR2_X1    g22712(.A1(new_n23006_), .A2(new_n23001_), .Z(new_n23010_));
  INV_X1     g22713(.I(new_n23010_), .ZN(new_n23011_));
  AOI21_X1   g22714(.A1(new_n22997_), .A2(new_n23011_), .B(new_n23009_), .ZN(new_n23012_));
  XOR2_X1    g22715(.A1(new_n22897_), .A2(new_n23012_), .Z(new_n23013_));
  NOR2_X1    g22716(.A1(new_n23013_), .A2(new_n22895_), .ZN(new_n23014_));
  INV_X1     g22717(.I(new_n22897_), .ZN(new_n23015_));
  NOR2_X1    g22718(.A1(new_n23015_), .A2(new_n23012_), .ZN(new_n23016_));
  INV_X1     g22719(.I(new_n23016_), .ZN(new_n23017_));
  NAND2_X1   g22720(.A1(new_n23015_), .A2(new_n23012_), .ZN(new_n23018_));
  NAND2_X1   g22721(.A1(new_n23017_), .A2(new_n23018_), .ZN(new_n23019_));
  AOI21_X1   g22722(.A1(new_n22895_), .A2(new_n23019_), .B(new_n23014_), .ZN(new_n23020_));
  NAND2_X1   g22723(.A1(new_n22872_), .A2(new_n22875_), .ZN(new_n23021_));
  XOR2_X1    g22724(.A1(new_n22873_), .A2(\a[35] ), .Z(new_n23022_));
  OAI21_X1   g22725(.A1(new_n22872_), .A2(new_n22875_), .B(new_n23022_), .ZN(new_n23023_));
  NAND2_X1   g22726(.A1(new_n23023_), .A2(new_n23021_), .ZN(new_n23024_));
  INV_X1     g22727(.I(new_n23024_), .ZN(new_n23025_));
  XOR2_X1    g22728(.A1(new_n23020_), .A2(new_n23025_), .Z(new_n23026_));
  INV_X1     g22729(.I(new_n23026_), .ZN(new_n23027_));
  NAND2_X1   g22730(.A1(new_n22882_), .A2(new_n23027_), .ZN(new_n23028_));
  XNOR2_X1   g22731(.A1(new_n23028_), .A2(new_n22887_), .ZN(new_n23029_));
  XOR2_X1    g22732(.A1(new_n22884_), .A2(new_n23029_), .Z(\f[99] ));
  NOR2_X1    g22733(.A1(new_n23020_), .A2(new_n23024_), .ZN(new_n23031_));
  NOR2_X1    g22734(.A1(new_n22886_), .A2(new_n23027_), .ZN(new_n23032_));
  AOI21_X1   g22735(.A1(new_n22886_), .A2(new_n23027_), .B(new_n22885_), .ZN(new_n23033_));
  NOR2_X1    g22736(.A1(new_n23033_), .A2(new_n23032_), .ZN(new_n23034_));
  NAND2_X1   g22737(.A1(new_n22754_), .A2(new_n23034_), .ZN(new_n23035_));
  NOR2_X1    g22738(.A1(new_n5112_), .A2(new_n5107_), .ZN(new_n23036_));
  NAND2_X1   g22739(.A1(new_n16148_), .A2(new_n4860_), .ZN(new_n23037_));
  OAI21_X1   g22740(.A1(new_n23036_), .A2(new_n23037_), .B(new_n4859_), .ZN(new_n23038_));
  XNOR2_X1   g22741(.A1(new_n14978_), .A2(new_n23038_), .ZN(new_n23039_));
  NAND2_X1   g22742(.A1(new_n22997_), .A2(new_n23008_), .ZN(new_n23040_));
  NAND2_X1   g22743(.A1(new_n23040_), .A2(new_n23004_), .ZN(new_n23041_));
  OAI22_X1   g22744(.A1(new_n6644_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n6647_), .ZN(new_n23042_));
  OAI21_X1   g22745(.A1(new_n11744_), .A2(new_n7284_), .B(new_n23042_), .ZN(new_n23043_));
  AOI21_X1   g22746(.A1(new_n23043_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n23044_));
  XNOR2_X1   g22747(.A1(new_n12546_), .A2(new_n23044_), .ZN(new_n23045_));
  AOI22_X1   g22748(.A1(new_n8631_), .A2(\b[51] ), .B1(\b[52] ), .B2(new_n9382_), .ZN(new_n23046_));
  AOI21_X1   g22749(.A1(\b[50] ), .A2(new_n9731_), .B(new_n23046_), .ZN(new_n23047_));
  OAI21_X1   g22750(.A1(new_n23047_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n23048_));
  XOR2_X1    g22751(.A1(new_n10035_), .A2(new_n23048_), .Z(new_n23049_));
  AOI22_X1   g22752(.A1(new_n10969_), .A2(new_n22614_), .B1(new_n11394_), .B2(\b[44] ), .ZN(new_n23050_));
  OAI21_X1   g22753(.A1(new_n23050_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n23051_));
  XOR2_X1    g22754(.A1(new_n7874_), .A2(new_n23051_), .Z(new_n23052_));
  INV_X1     g22755(.I(new_n23052_), .ZN(new_n23053_));
  OAI22_X1   g22756(.A1(new_n13880_), .A2(new_n5922_), .B1(new_n5353_), .B2(new_n13885_), .ZN(new_n23054_));
  AOI21_X1   g22757(.A1(new_n23054_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23055_));
  XOR2_X1    g22758(.A1(new_n5926_), .A2(new_n23055_), .Z(new_n23056_));
  INV_X1     g22759(.I(new_n23056_), .ZN(new_n23057_));
  NAND2_X1   g22760(.A1(new_n22920_), .A2(new_n22791_), .ZN(new_n23058_));
  NAND2_X1   g22761(.A1(new_n23058_), .A2(new_n22919_), .ZN(new_n23059_));
  NOR2_X1    g22762(.A1(new_n13476_), .A2(new_n4774_), .ZN(new_n23060_));
  XOR2_X1    g22763(.A1(new_n14736_), .A2(new_n4774_), .Z(new_n23061_));
  NAND2_X1   g22764(.A1(new_n23061_), .A2(\b[37] ), .ZN(new_n23062_));
  XOR2_X1    g22765(.A1(new_n23062_), .A2(new_n23060_), .Z(new_n23063_));
  NOR2_X1    g22766(.A1(new_n23059_), .A2(new_n23063_), .ZN(new_n23064_));
  INV_X1     g22767(.I(new_n23064_), .ZN(new_n23065_));
  NAND2_X1   g22768(.A1(new_n23059_), .A2(new_n23063_), .ZN(new_n23066_));
  NAND2_X1   g22769(.A1(new_n23065_), .A2(new_n23066_), .ZN(new_n23067_));
  INV_X1     g22770(.I(new_n23063_), .ZN(new_n23068_));
  XOR2_X1    g22771(.A1(new_n23059_), .A2(new_n23068_), .Z(new_n23069_));
  NOR2_X1    g22772(.A1(new_n23057_), .A2(new_n23069_), .ZN(new_n23070_));
  AOI21_X1   g22773(.A1(new_n23057_), .A2(new_n23067_), .B(new_n23070_), .ZN(new_n23071_));
  OAI21_X1   g22774(.A1(new_n22908_), .A2(new_n22926_), .B(new_n22928_), .ZN(new_n23072_));
  INV_X1     g22775(.I(new_n23072_), .ZN(new_n23073_));
  AOI22_X1   g22776(.A1(new_n13078_), .A2(\b[41] ), .B1(new_n7194_), .B2(new_n12218_), .ZN(new_n23074_));
  OAI21_X1   g22777(.A1(new_n23074_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23075_));
  XNOR2_X1   g22778(.A1(new_n6851_), .A2(new_n23075_), .ZN(new_n23076_));
  NOR2_X1    g22779(.A1(new_n23076_), .A2(new_n23073_), .ZN(new_n23077_));
  AND2_X2    g22780(.A1(new_n23076_), .A2(new_n23073_), .Z(new_n23078_));
  NOR2_X1    g22781(.A1(new_n23078_), .A2(new_n23077_), .ZN(new_n23079_));
  NOR2_X1    g22782(.A1(new_n23079_), .A2(new_n23071_), .ZN(new_n23080_));
  INV_X1     g22783(.I(new_n23071_), .ZN(new_n23081_));
  XOR2_X1    g22784(.A1(new_n23076_), .A2(new_n23072_), .Z(new_n23082_));
  NOR2_X1    g22785(.A1(new_n23081_), .A2(new_n23082_), .ZN(new_n23083_));
  NOR2_X1    g22786(.A1(new_n23083_), .A2(new_n23080_), .ZN(new_n23084_));
  NAND2_X1   g22787(.A1(new_n22941_), .A2(new_n22930_), .ZN(new_n23085_));
  AOI21_X1   g22788(.A1(new_n22940_), .A2(new_n23085_), .B(new_n23084_), .ZN(new_n23086_));
  NAND2_X1   g22789(.A1(new_n23085_), .A2(new_n22940_), .ZN(new_n23087_));
  NOR3_X1    g22790(.A1(new_n23087_), .A2(new_n23080_), .A3(new_n23083_), .ZN(new_n23088_));
  OAI21_X1   g22791(.A1(new_n23086_), .A2(new_n23088_), .B(new_n23053_), .ZN(new_n23089_));
  XOR2_X1    g22792(.A1(new_n23084_), .A2(new_n23087_), .Z(new_n23090_));
  OR2_X2     g22793(.A1(new_n23090_), .A2(new_n23053_), .Z(new_n23091_));
  NAND2_X1   g22794(.A1(new_n22952_), .A2(new_n22949_), .ZN(new_n23092_));
  NAND2_X1   g22795(.A1(new_n23092_), .A2(new_n22951_), .ZN(new_n23093_));
  INV_X1     g22796(.I(new_n23093_), .ZN(new_n23094_));
  AOI22_X1   g22797(.A1(new_n11415_), .A2(new_n9291_), .B1(\b[47] ), .B2(new_n10145_), .ZN(new_n23095_));
  OAI21_X1   g22798(.A1(new_n23095_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23096_));
  XNOR2_X1   g22799(.A1(new_n8952_), .A2(new_n23096_), .ZN(new_n23097_));
  NOR2_X1    g22800(.A1(new_n23094_), .A2(new_n23097_), .ZN(new_n23098_));
  INV_X1     g22801(.I(new_n23098_), .ZN(new_n23099_));
  NAND2_X1   g22802(.A1(new_n23094_), .A2(new_n23097_), .ZN(new_n23100_));
  AOI22_X1   g22803(.A1(new_n23099_), .A2(new_n23100_), .B1(new_n23089_), .B2(new_n23091_), .ZN(new_n23101_));
  NAND2_X1   g22804(.A1(new_n23091_), .A2(new_n23089_), .ZN(new_n23102_));
  XOR2_X1    g22805(.A1(new_n23093_), .A2(new_n23097_), .Z(new_n23103_));
  NOR2_X1    g22806(.A1(new_n23103_), .A2(new_n23102_), .ZN(new_n23104_));
  NOR2_X1    g22807(.A1(new_n23101_), .A2(new_n23104_), .ZN(new_n23105_));
  NOR2_X1    g22808(.A1(new_n22964_), .A2(new_n22955_), .ZN(new_n23106_));
  NOR2_X1    g22809(.A1(new_n23106_), .A2(new_n22962_), .ZN(new_n23107_));
  NOR2_X1    g22810(.A1(new_n23105_), .A2(new_n23107_), .ZN(new_n23108_));
  NOR4_X1    g22811(.A1(new_n23101_), .A2(new_n22962_), .A3(new_n23106_), .A4(new_n23104_), .ZN(new_n23109_));
  NOR2_X1    g22812(.A1(new_n23108_), .A2(new_n23109_), .ZN(new_n23110_));
  NOR2_X1    g22813(.A1(new_n23110_), .A2(new_n23049_), .ZN(new_n23111_));
  INV_X1     g22814(.I(new_n23049_), .ZN(new_n23112_));
  XNOR2_X1   g22815(.A1(new_n23105_), .A2(new_n23107_), .ZN(new_n23113_));
  NOR2_X1    g22816(.A1(new_n23113_), .A2(new_n23112_), .ZN(new_n23114_));
  NOR2_X1    g22817(.A1(new_n23114_), .A2(new_n23111_), .ZN(new_n23115_));
  NAND2_X1   g22818(.A1(new_n22977_), .A2(new_n22974_), .ZN(new_n23116_));
  NAND2_X1   g22819(.A1(new_n23116_), .A2(new_n22976_), .ZN(new_n23117_));
  INV_X1     g22820(.I(new_n23117_), .ZN(new_n23118_));
  OAI22_X1   g22821(.A1(new_n7619_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n8309_), .ZN(new_n23119_));
  OAI21_X1   g22822(.A1(new_n10477_), .A2(new_n7947_), .B(new_n23119_), .ZN(new_n23120_));
  AOI21_X1   g22823(.A1(new_n23120_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23121_));
  XOR2_X1    g22824(.A1(new_n11298_), .A2(new_n23121_), .Z(new_n23122_));
  NOR2_X1    g22825(.A1(new_n23118_), .A2(new_n23122_), .ZN(new_n23123_));
  INV_X1     g22826(.I(new_n23122_), .ZN(new_n23124_));
  NOR2_X1    g22827(.A1(new_n23117_), .A2(new_n23124_), .ZN(new_n23125_));
  NOR2_X1    g22828(.A1(new_n23123_), .A2(new_n23125_), .ZN(new_n23126_));
  NOR2_X1    g22829(.A1(new_n23126_), .A2(new_n23115_), .ZN(new_n23127_));
  INV_X1     g22830(.I(new_n23115_), .ZN(new_n23128_));
  XOR2_X1    g22831(.A1(new_n23117_), .A2(new_n23122_), .Z(new_n23129_));
  NOR2_X1    g22832(.A1(new_n23129_), .A2(new_n23128_), .ZN(new_n23130_));
  NOR2_X1    g22833(.A1(new_n23127_), .A2(new_n23130_), .ZN(new_n23131_));
  OAI21_X1   g22834(.A1(new_n22900_), .A2(new_n22982_), .B(new_n22983_), .ZN(new_n23132_));
  INV_X1     g22835(.I(new_n23132_), .ZN(new_n23133_));
  NOR2_X1    g22836(.A1(new_n23133_), .A2(new_n23131_), .ZN(new_n23134_));
  NOR3_X1    g22837(.A1(new_n23132_), .A2(new_n23127_), .A3(new_n23130_), .ZN(new_n23135_));
  NOR2_X1    g22838(.A1(new_n23134_), .A2(new_n23135_), .ZN(new_n23136_));
  NOR2_X1    g22839(.A1(new_n23136_), .A2(new_n23045_), .ZN(new_n23137_));
  INV_X1     g22840(.I(new_n23045_), .ZN(new_n23138_));
  XOR2_X1    g22841(.A1(new_n23131_), .A2(new_n23132_), .Z(new_n23139_));
  NOR2_X1    g22842(.A1(new_n23139_), .A2(new_n23138_), .ZN(new_n23140_));
  NOR2_X1    g22843(.A1(new_n23140_), .A2(new_n23137_), .ZN(new_n23141_));
  NAND2_X1   g22844(.A1(new_n22995_), .A2(new_n22898_), .ZN(new_n23142_));
  NAND2_X1   g22845(.A1(new_n23142_), .A2(new_n22994_), .ZN(new_n23143_));
  OAI22_X1   g22846(.A1(new_n5993_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n5991_), .ZN(new_n23144_));
  OAI21_X1   g22847(.A1(new_n12970_), .A2(new_n5997_), .B(new_n23144_), .ZN(new_n23145_));
  AOI21_X1   g22848(.A1(new_n23145_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n23146_));
  XOR2_X1    g22849(.A1(new_n13784_), .A2(new_n23146_), .Z(new_n23147_));
  XOR2_X1    g22850(.A1(new_n23143_), .A2(new_n23147_), .Z(new_n23148_));
  NOR2_X1    g22851(.A1(new_n23148_), .A2(new_n23141_), .ZN(new_n23149_));
  INV_X1     g22852(.I(new_n23141_), .ZN(new_n23150_));
  INV_X1     g22853(.I(new_n23143_), .ZN(new_n23151_));
  NOR2_X1    g22854(.A1(new_n23151_), .A2(new_n23147_), .ZN(new_n23152_));
  INV_X1     g22855(.I(new_n23152_), .ZN(new_n23153_));
  NAND2_X1   g22856(.A1(new_n23151_), .A2(new_n23147_), .ZN(new_n23154_));
  AOI21_X1   g22857(.A1(new_n23153_), .A2(new_n23154_), .B(new_n23150_), .ZN(new_n23155_));
  NOR2_X1    g22858(.A1(new_n23155_), .A2(new_n23149_), .ZN(new_n23156_));
  NOR2_X1    g22859(.A1(new_n23156_), .A2(new_n23041_), .ZN(new_n23157_));
  INV_X1     g22860(.I(new_n23157_), .ZN(new_n23158_));
  NAND2_X1   g22861(.A1(new_n23156_), .A2(new_n23041_), .ZN(new_n23159_));
  AOI21_X1   g22862(.A1(new_n23158_), .A2(new_n23159_), .B(new_n23039_), .ZN(new_n23160_));
  INV_X1     g22863(.I(new_n23039_), .ZN(new_n23161_));
  XNOR2_X1   g22864(.A1(new_n23156_), .A2(new_n23041_), .ZN(new_n23162_));
  NOR2_X1    g22865(.A1(new_n23162_), .A2(new_n23161_), .ZN(new_n23163_));
  NOR2_X1    g22866(.A1(new_n23163_), .A2(new_n23160_), .ZN(new_n23164_));
  INV_X1     g22867(.I(new_n23164_), .ZN(new_n23165_));
  OAI21_X1   g22868(.A1(new_n22895_), .A2(new_n23016_), .B(new_n23018_), .ZN(new_n23166_));
  NAND2_X1   g22869(.A1(new_n23165_), .A2(new_n23166_), .ZN(new_n23167_));
  XOR2_X1    g22870(.A1(new_n23035_), .A2(new_n23167_), .Z(new_n23168_));
  XOR2_X1    g22871(.A1(new_n23168_), .A2(new_n23031_), .Z(\f[100] ));
  INV_X1     g22872(.I(new_n23031_), .ZN(new_n23170_));
  NOR2_X1    g22873(.A1(new_n23170_), .A2(new_n23164_), .ZN(new_n23171_));
  INV_X1     g22874(.I(new_n23171_), .ZN(new_n23172_));
  OAI21_X1   g22875(.A1(new_n23031_), .A2(new_n23165_), .B(new_n23166_), .ZN(new_n23173_));
  INV_X1     g22876(.I(new_n23173_), .ZN(new_n23174_));
  NAND3_X1   g22877(.A1(new_n22754_), .A2(new_n23034_), .A3(new_n23174_), .ZN(new_n23175_));
  NAND2_X1   g22878(.A1(new_n23175_), .A2(new_n23172_), .ZN(new_n23176_));
  OAI21_X1   g22879(.A1(new_n23039_), .A2(new_n23157_), .B(new_n23159_), .ZN(new_n23177_));
  INV_X1     g22880(.I(new_n23177_), .ZN(new_n23178_));
  OAI22_X1   g22881(.A1(new_n5993_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n5991_), .ZN(new_n23179_));
  OAI21_X1   g22882(.A1(new_n13367_), .A2(new_n5997_), .B(new_n23179_), .ZN(new_n23180_));
  AOI21_X1   g22883(.A1(new_n23180_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n23181_));
  XOR2_X1    g22884(.A1(new_n14213_), .A2(new_n23181_), .Z(new_n23182_));
  OAI22_X1   g22885(.A1(new_n7619_), .A2(new_n11738_), .B1(new_n11744_), .B2(new_n8309_), .ZN(new_n23183_));
  OAI21_X1   g22886(.A1(new_n10862_), .A2(new_n7947_), .B(new_n23183_), .ZN(new_n23184_));
  AOI21_X1   g22887(.A1(new_n23184_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23185_));
  XNOR2_X1   g22888(.A1(new_n11748_), .A2(new_n23185_), .ZN(new_n23186_));
  INV_X1     g22889(.I(new_n23109_), .ZN(new_n23187_));
  AOI21_X1   g22890(.A1(new_n23187_), .A2(new_n23112_), .B(new_n23108_), .ZN(new_n23188_));
  OAI22_X1   g22891(.A1(new_n8644_), .A2(new_n10031_), .B1(new_n10477_), .B2(new_n9388_), .ZN(new_n23189_));
  OAI21_X1   g22892(.A1(new_n10025_), .A2(new_n10154_), .B(new_n23189_), .ZN(new_n23190_));
  AOI21_X1   g22893(.A1(new_n23190_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n23191_));
  XOR2_X1    g22894(.A1(new_n10476_), .A2(new_n23191_), .Z(new_n23192_));
  INV_X1     g22895(.I(new_n9296_), .ZN(new_n23193_));
  AOI22_X1   g22896(.A1(new_n11415_), .A2(new_n23193_), .B1(\b[48] ), .B2(new_n10145_), .ZN(new_n23194_));
  OAI21_X1   g22897(.A1(new_n23194_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23195_));
  XOR2_X1    g22898(.A1(new_n9299_), .A2(new_n23195_), .Z(new_n23196_));
  OAI21_X1   g22899(.A1(new_n23056_), .A2(new_n23064_), .B(new_n23066_), .ZN(new_n23197_));
  NOR2_X1    g22900(.A1(new_n13476_), .A2(new_n5068_), .ZN(new_n23198_));
  XOR2_X1    g22901(.A1(new_n14736_), .A2(new_n5068_), .Z(new_n23199_));
  NAND2_X1   g22902(.A1(new_n23199_), .A2(\b[38] ), .ZN(new_n23200_));
  XOR2_X1    g22903(.A1(new_n23200_), .A2(new_n23198_), .Z(new_n23201_));
  NOR2_X1    g22904(.A1(new_n23068_), .A2(new_n23201_), .ZN(new_n23202_));
  INV_X1     g22905(.I(new_n23201_), .ZN(new_n23203_));
  NOR2_X1    g22906(.A1(new_n23203_), .A2(new_n23063_), .ZN(new_n23204_));
  NOR2_X1    g22907(.A1(new_n23202_), .A2(new_n23204_), .ZN(new_n23205_));
  INV_X1     g22908(.I(new_n23205_), .ZN(new_n23206_));
  XOR2_X1    g22909(.A1(new_n23063_), .A2(new_n23201_), .Z(new_n23207_));
  NOR2_X1    g22910(.A1(new_n23197_), .A2(new_n23207_), .ZN(new_n23208_));
  AOI21_X1   g22911(.A1(new_n23197_), .A2(new_n23206_), .B(new_n23208_), .ZN(new_n23209_));
  AOI22_X1   g22912(.A1(new_n13078_), .A2(\b[42] ), .B1(new_n22330_), .B2(new_n12218_), .ZN(new_n23210_));
  OAI21_X1   g22913(.A1(new_n23210_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23211_));
  XOR2_X1    g22914(.A1(new_n7202_), .A2(new_n23211_), .Z(new_n23212_));
  OAI22_X1   g22915(.A1(new_n13880_), .A2(new_n6531_), .B1(new_n5913_), .B2(new_n13885_), .ZN(new_n23213_));
  AOI21_X1   g22916(.A1(new_n23213_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23214_));
  XOR2_X1    g22917(.A1(new_n6233_), .A2(new_n23214_), .Z(new_n23215_));
  NOR2_X1    g22918(.A1(new_n23212_), .A2(new_n23215_), .ZN(new_n23216_));
  INV_X1     g22919(.I(new_n23216_), .ZN(new_n23217_));
  NAND2_X1   g22920(.A1(new_n23212_), .A2(new_n23215_), .ZN(new_n23218_));
  AOI21_X1   g22921(.A1(new_n23217_), .A2(new_n23218_), .B(new_n23209_), .ZN(new_n23219_));
  INV_X1     g22922(.I(new_n23209_), .ZN(new_n23220_));
  XNOR2_X1   g22923(.A1(new_n23212_), .A2(new_n23215_), .ZN(new_n23221_));
  NOR2_X1    g22924(.A1(new_n23221_), .A2(new_n23220_), .ZN(new_n23222_));
  NOR2_X1    g22925(.A1(new_n23222_), .A2(new_n23219_), .ZN(new_n23223_));
  AOI22_X1   g22926(.A1(new_n10969_), .A2(new_n8557_), .B1(new_n11394_), .B2(\b[45] ), .ZN(new_n23224_));
  OAI21_X1   g22927(.A1(new_n23224_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n23225_));
  XNOR2_X1   g22928(.A1(new_n8217_), .A2(new_n23225_), .ZN(new_n23226_));
  INV_X1     g22929(.I(new_n23078_), .ZN(new_n23227_));
  AOI21_X1   g22930(.A1(new_n23081_), .A2(new_n23227_), .B(new_n23077_), .ZN(new_n23228_));
  NOR2_X1    g22931(.A1(new_n23226_), .A2(new_n23228_), .ZN(new_n23229_));
  INV_X1     g22932(.I(new_n23226_), .ZN(new_n23230_));
  INV_X1     g22933(.I(new_n23228_), .ZN(new_n23231_));
  NOR2_X1    g22934(.A1(new_n23230_), .A2(new_n23231_), .ZN(new_n23232_));
  NOR2_X1    g22935(.A1(new_n23232_), .A2(new_n23229_), .ZN(new_n23233_));
  XNOR2_X1   g22936(.A1(new_n23226_), .A2(new_n23228_), .ZN(new_n23234_));
  MUX2_X1    g22937(.I0(new_n23233_), .I1(new_n23234_), .S(new_n23223_), .Z(new_n23235_));
  NOR2_X1    g22938(.A1(new_n23088_), .A2(new_n23052_), .ZN(new_n23236_));
  NOR2_X1    g22939(.A1(new_n23236_), .A2(new_n23086_), .ZN(new_n23237_));
  XNOR2_X1   g22940(.A1(new_n23235_), .A2(new_n23237_), .ZN(new_n23238_));
  NOR2_X1    g22941(.A1(new_n23238_), .A2(new_n23196_), .ZN(new_n23239_));
  INV_X1     g22942(.I(new_n23196_), .ZN(new_n23240_));
  NOR2_X1    g22943(.A1(new_n23235_), .A2(new_n23237_), .ZN(new_n23241_));
  INV_X1     g22944(.I(new_n23241_), .ZN(new_n23242_));
  NAND2_X1   g22945(.A1(new_n23235_), .A2(new_n23237_), .ZN(new_n23243_));
  AOI21_X1   g22946(.A1(new_n23242_), .A2(new_n23243_), .B(new_n23240_), .ZN(new_n23244_));
  NOR2_X1    g22947(.A1(new_n23239_), .A2(new_n23244_), .ZN(new_n23245_));
  AOI21_X1   g22948(.A1(new_n23102_), .A2(new_n23100_), .B(new_n23098_), .ZN(new_n23246_));
  XOR2_X1    g22949(.A1(new_n23245_), .A2(new_n23246_), .Z(new_n23247_));
  NOR2_X1    g22950(.A1(new_n23247_), .A2(new_n23192_), .ZN(new_n23248_));
  INV_X1     g22951(.I(new_n23192_), .ZN(new_n23249_));
  INV_X1     g22952(.I(new_n23245_), .ZN(new_n23250_));
  NOR2_X1    g22953(.A1(new_n23250_), .A2(new_n23246_), .ZN(new_n23251_));
  INV_X1     g22954(.I(new_n23251_), .ZN(new_n23252_));
  NAND2_X1   g22955(.A1(new_n23250_), .A2(new_n23246_), .ZN(new_n23253_));
  AOI21_X1   g22956(.A1(new_n23252_), .A2(new_n23253_), .B(new_n23249_), .ZN(new_n23254_));
  NOR2_X1    g22957(.A1(new_n23254_), .A2(new_n23248_), .ZN(new_n23255_));
  XOR2_X1    g22958(.A1(new_n23255_), .A2(new_n23188_), .Z(new_n23256_));
  NOR2_X1    g22959(.A1(new_n23256_), .A2(new_n23186_), .ZN(new_n23257_));
  INV_X1     g22960(.I(new_n23188_), .ZN(new_n23258_));
  NOR2_X1    g22961(.A1(new_n23255_), .A2(new_n23258_), .ZN(new_n23259_));
  INV_X1     g22962(.I(new_n23259_), .ZN(new_n23260_));
  NAND2_X1   g22963(.A1(new_n23255_), .A2(new_n23258_), .ZN(new_n23261_));
  NAND2_X1   g22964(.A1(new_n23260_), .A2(new_n23261_), .ZN(new_n23262_));
  AOI21_X1   g22965(.A1(new_n23186_), .A2(new_n23262_), .B(new_n23257_), .ZN(new_n23263_));
  OAI22_X1   g22966(.A1(new_n6644_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n6647_), .ZN(new_n23264_));
  OAI21_X1   g22967(.A1(new_n12536_), .A2(new_n7284_), .B(new_n23264_), .ZN(new_n23265_));
  AOI21_X1   g22968(.A1(new_n23265_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n23266_));
  XOR2_X1    g22969(.A1(new_n12969_), .A2(new_n23266_), .Z(new_n23267_));
  NOR2_X1    g22970(.A1(new_n23115_), .A2(new_n23125_), .ZN(new_n23268_));
  NOR2_X1    g22971(.A1(new_n23268_), .A2(new_n23123_), .ZN(new_n23269_));
  XNOR2_X1   g22972(.A1(new_n23269_), .A2(new_n23267_), .ZN(new_n23270_));
  NOR2_X1    g22973(.A1(new_n23263_), .A2(new_n23270_), .ZN(new_n23271_));
  NOR2_X1    g22974(.A1(new_n23269_), .A2(new_n23267_), .ZN(new_n23272_));
  INV_X1     g22975(.I(new_n23272_), .ZN(new_n23273_));
  NAND2_X1   g22976(.A1(new_n23269_), .A2(new_n23267_), .ZN(new_n23274_));
  NAND2_X1   g22977(.A1(new_n23273_), .A2(new_n23274_), .ZN(new_n23275_));
  AOI21_X1   g22978(.A1(new_n23263_), .A2(new_n23275_), .B(new_n23271_), .ZN(new_n23276_));
  NOR2_X1    g22979(.A1(new_n23135_), .A2(new_n23045_), .ZN(new_n23277_));
  NOR2_X1    g22980(.A1(new_n23277_), .A2(new_n23134_), .ZN(new_n23278_));
  NOR2_X1    g22981(.A1(new_n23276_), .A2(new_n23278_), .ZN(new_n23279_));
  INV_X1     g22982(.I(new_n23279_), .ZN(new_n23280_));
  NAND2_X1   g22983(.A1(new_n23276_), .A2(new_n23278_), .ZN(new_n23281_));
  AOI21_X1   g22984(.A1(new_n23280_), .A2(new_n23281_), .B(new_n23182_), .ZN(new_n23282_));
  XOR2_X1    g22985(.A1(new_n23276_), .A2(new_n23278_), .Z(new_n23283_));
  AOI21_X1   g22986(.A1(new_n23182_), .A2(new_n23283_), .B(new_n23282_), .ZN(new_n23284_));
  OAI21_X1   g22987(.A1(new_n5420_), .A2(new_n5112_), .B(new_n16487_), .ZN(new_n23285_));
  NAND2_X1   g22988(.A1(new_n23154_), .A2(new_n23150_), .ZN(new_n23286_));
  NAND2_X1   g22989(.A1(new_n23286_), .A2(new_n23153_), .ZN(new_n23287_));
  XNOR2_X1   g22990(.A1(new_n23287_), .A2(new_n23285_), .ZN(new_n23288_));
  XNOR2_X1   g22991(.A1(new_n23288_), .A2(new_n23284_), .ZN(new_n23289_));
  NOR2_X1    g22992(.A1(new_n23289_), .A2(\a[38] ), .ZN(new_n23290_));
  NAND2_X1   g22993(.A1(new_n23289_), .A2(\a[38] ), .ZN(new_n23291_));
  INV_X1     g22994(.I(new_n23291_), .ZN(new_n23292_));
  NOR2_X1    g22995(.A1(new_n23292_), .A2(new_n23290_), .ZN(new_n23293_));
  XOR2_X1    g22996(.A1(new_n23293_), .A2(new_n23178_), .Z(new_n23294_));
  NAND2_X1   g22997(.A1(new_n23176_), .A2(new_n23294_), .ZN(new_n23295_));
  XOR2_X1    g22998(.A1(new_n23293_), .A2(new_n23178_), .Z(new_n23296_));
  OAI21_X1   g22999(.A1(new_n23176_), .A2(new_n23296_), .B(new_n23295_), .ZN(\f[101] ));
  INV_X1     g23000(.I(new_n23293_), .ZN(new_n23298_));
  NAND2_X1   g23001(.A1(new_n23298_), .A2(new_n23177_), .ZN(new_n23299_));
  OAI22_X1   g23002(.A1(new_n5993_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n5991_), .ZN(new_n23300_));
  OAI21_X1   g23003(.A1(new_n13785_), .A2(new_n5997_), .B(new_n23300_), .ZN(new_n23301_));
  AOI21_X1   g23004(.A1(new_n23301_), .A2(new_n5681_), .B(new_n5993_), .ZN(new_n23302_));
  XNOR2_X1   g23005(.A1(new_n14599_), .A2(new_n23302_), .ZN(new_n23303_));
  AOI21_X1   g23006(.A1(new_n23276_), .A2(new_n23278_), .B(new_n23182_), .ZN(new_n23304_));
  NOR2_X1    g23007(.A1(new_n23304_), .A2(new_n23279_), .ZN(new_n23305_));
  INV_X1     g23008(.I(new_n23305_), .ZN(new_n23306_));
  OAI21_X1   g23009(.A1(new_n23186_), .A2(new_n23259_), .B(new_n23261_), .ZN(new_n23307_));
  INV_X1     g23010(.I(new_n23307_), .ZN(new_n23308_));
  AOI21_X1   g23011(.A1(new_n23249_), .A2(new_n23253_), .B(new_n23251_), .ZN(new_n23309_));
  OAI22_X1   g23012(.A1(new_n8644_), .A2(new_n10477_), .B1(new_n10862_), .B2(new_n9388_), .ZN(new_n23310_));
  OAI21_X1   g23013(.A1(new_n10031_), .A2(new_n10154_), .B(new_n23310_), .ZN(new_n23311_));
  AOI21_X1   g23014(.A1(new_n23311_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n23312_));
  XNOR2_X1   g23015(.A1(new_n10866_), .A2(new_n23312_), .ZN(new_n23313_));
  INV_X1     g23016(.I(new_n23313_), .ZN(new_n23314_));
  AOI21_X1   g23017(.A1(new_n23240_), .A2(new_n23243_), .B(new_n23241_), .ZN(new_n23315_));
  INV_X1     g23018(.I(new_n23315_), .ZN(new_n23316_));
  INV_X1     g23019(.I(new_n23204_), .ZN(new_n23317_));
  AOI21_X1   g23020(.A1(new_n23197_), .A2(new_n23317_), .B(new_n23202_), .ZN(new_n23318_));
  OAI22_X1   g23021(.A1(new_n13880_), .A2(new_n6539_), .B1(new_n5921_), .B2(new_n13885_), .ZN(new_n23319_));
  AOI21_X1   g23022(.A1(new_n23319_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23320_));
  XOR2_X1    g23023(.A1(new_n6543_), .A2(new_n23320_), .Z(new_n23321_));
  INV_X1     g23024(.I(new_n23321_), .ZN(new_n23322_));
  NOR2_X1    g23025(.A1(new_n13476_), .A2(new_n5353_), .ZN(new_n23323_));
  XOR2_X1    g23026(.A1(new_n14736_), .A2(new_n5353_), .Z(new_n23324_));
  NAND2_X1   g23027(.A1(new_n23324_), .A2(\b[39] ), .ZN(new_n23325_));
  XOR2_X1    g23028(.A1(new_n23325_), .A2(new_n23323_), .Z(new_n23326_));
  XOR2_X1    g23029(.A1(new_n23326_), .A2(\a[38] ), .Z(new_n23327_));
  NOR2_X1    g23030(.A1(new_n23327_), .A2(new_n23063_), .ZN(new_n23328_));
  NOR2_X1    g23031(.A1(new_n23326_), .A2(new_n4860_), .ZN(new_n23329_));
  INV_X1     g23032(.I(new_n23329_), .ZN(new_n23330_));
  NAND2_X1   g23033(.A1(new_n23326_), .A2(new_n4860_), .ZN(new_n23331_));
  AOI21_X1   g23034(.A1(new_n23330_), .A2(new_n23331_), .B(new_n23068_), .ZN(new_n23332_));
  NOR2_X1    g23035(.A1(new_n23328_), .A2(new_n23332_), .ZN(new_n23333_));
  NOR2_X1    g23036(.A1(new_n23322_), .A2(new_n23333_), .ZN(new_n23334_));
  INV_X1     g23037(.I(new_n23334_), .ZN(new_n23335_));
  NAND2_X1   g23038(.A1(new_n23322_), .A2(new_n23333_), .ZN(new_n23336_));
  AOI21_X1   g23039(.A1(new_n23335_), .A2(new_n23336_), .B(new_n23318_), .ZN(new_n23337_));
  INV_X1     g23040(.I(new_n23318_), .ZN(new_n23338_));
  XOR2_X1    g23041(.A1(new_n23321_), .A2(new_n23333_), .Z(new_n23339_));
  NOR2_X1    g23042(.A1(new_n23339_), .A2(new_n23338_), .ZN(new_n23340_));
  NOR2_X1    g23043(.A1(new_n23337_), .A2(new_n23340_), .ZN(new_n23341_));
  NAND2_X1   g23044(.A1(new_n23218_), .A2(new_n23220_), .ZN(new_n23342_));
  AOI22_X1   g23045(.A1(new_n13078_), .A2(\b[43] ), .B1(new_n7866_), .B2(new_n12218_), .ZN(new_n23343_));
  OAI21_X1   g23046(.A1(new_n23343_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23344_));
  XNOR2_X1   g23047(.A1(new_n7516_), .A2(new_n23344_), .ZN(new_n23345_));
  AOI21_X1   g23048(.A1(new_n23342_), .A2(new_n23217_), .B(new_n23345_), .ZN(new_n23346_));
  INV_X1     g23049(.I(new_n23346_), .ZN(new_n23347_));
  NAND2_X1   g23050(.A1(new_n23342_), .A2(new_n23217_), .ZN(new_n23348_));
  INV_X1     g23051(.I(new_n23345_), .ZN(new_n23349_));
  NOR2_X1    g23052(.A1(new_n23348_), .A2(new_n23349_), .ZN(new_n23350_));
  INV_X1     g23053(.I(new_n23350_), .ZN(new_n23351_));
  AOI21_X1   g23054(.A1(new_n23351_), .A2(new_n23347_), .B(new_n23341_), .ZN(new_n23352_));
  INV_X1     g23055(.I(new_n23341_), .ZN(new_n23353_));
  XOR2_X1    g23056(.A1(new_n23348_), .A2(new_n23345_), .Z(new_n23354_));
  NOR2_X1    g23057(.A1(new_n23354_), .A2(new_n23353_), .ZN(new_n23355_));
  NOR2_X1    g23058(.A1(new_n23355_), .A2(new_n23352_), .ZN(new_n23356_));
  AOI22_X1   g23059(.A1(new_n10969_), .A2(new_n8565_), .B1(new_n11394_), .B2(\b[46] ), .ZN(new_n23357_));
  OAI21_X1   g23060(.A1(new_n23357_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n23358_));
  XOR2_X1    g23061(.A1(new_n8568_), .A2(new_n23358_), .Z(new_n23359_));
  INV_X1     g23062(.I(new_n23229_), .ZN(new_n23360_));
  OAI21_X1   g23063(.A1(new_n23223_), .A2(new_n23232_), .B(new_n23360_), .ZN(new_n23361_));
  XNOR2_X1   g23064(.A1(new_n23361_), .A2(new_n23359_), .ZN(new_n23362_));
  NAND2_X1   g23065(.A1(new_n23361_), .A2(new_n23359_), .ZN(new_n23363_));
  INV_X1     g23066(.I(new_n23363_), .ZN(new_n23364_));
  NOR2_X1    g23067(.A1(new_n23361_), .A2(new_n23359_), .ZN(new_n23365_));
  OAI21_X1   g23068(.A1(new_n23364_), .A2(new_n23365_), .B(new_n23356_), .ZN(new_n23366_));
  OAI21_X1   g23069(.A1(new_n23356_), .A2(new_n23362_), .B(new_n23366_), .ZN(new_n23367_));
  AOI22_X1   g23070(.A1(new_n11415_), .A2(new_n10027_), .B1(\b[49] ), .B2(new_n10145_), .ZN(new_n23368_));
  OAI21_X1   g23071(.A1(new_n23368_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23369_));
  XOR2_X1    g23072(.A1(new_n9642_), .A2(new_n23369_), .Z(new_n23370_));
  XOR2_X1    g23073(.A1(new_n23367_), .A2(new_n23370_), .Z(new_n23371_));
  NAND2_X1   g23074(.A1(new_n23371_), .A2(new_n23316_), .ZN(new_n23372_));
  NOR2_X1    g23075(.A1(new_n23367_), .A2(new_n23370_), .ZN(new_n23373_));
  NAND2_X1   g23076(.A1(new_n23367_), .A2(new_n23370_), .ZN(new_n23374_));
  INV_X1     g23077(.I(new_n23374_), .ZN(new_n23375_));
  OAI21_X1   g23078(.A1(new_n23375_), .A2(new_n23373_), .B(new_n23315_), .ZN(new_n23376_));
  NAND2_X1   g23079(.A1(new_n23372_), .A2(new_n23376_), .ZN(new_n23377_));
  XOR2_X1    g23080(.A1(new_n23377_), .A2(new_n23314_), .Z(new_n23378_));
  AND2_X2    g23081(.A1(new_n23377_), .A2(new_n23313_), .Z(new_n23379_));
  NOR2_X1    g23082(.A1(new_n23377_), .A2(new_n23313_), .ZN(new_n23380_));
  OAI21_X1   g23083(.A1(new_n23379_), .A2(new_n23380_), .B(new_n23309_), .ZN(new_n23381_));
  OAI21_X1   g23084(.A1(new_n23309_), .A2(new_n23378_), .B(new_n23381_), .ZN(new_n23382_));
  OAI22_X1   g23085(.A1(new_n7619_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n8309_), .ZN(new_n23383_));
  OAI21_X1   g23086(.A1(new_n11738_), .A2(new_n7947_), .B(new_n23383_), .ZN(new_n23384_));
  AOI21_X1   g23087(.A1(new_n23384_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23385_));
  XNOR2_X1   g23088(.A1(new_n12128_), .A2(new_n23385_), .ZN(new_n23386_));
  XNOR2_X1   g23089(.A1(new_n23382_), .A2(new_n23386_), .ZN(new_n23387_));
  NOR2_X1    g23090(.A1(new_n23382_), .A2(new_n23386_), .ZN(new_n23388_));
  NAND2_X1   g23091(.A1(new_n23382_), .A2(new_n23386_), .ZN(new_n23389_));
  INV_X1     g23092(.I(new_n23389_), .ZN(new_n23390_));
  OAI21_X1   g23093(.A1(new_n23390_), .A2(new_n23388_), .B(new_n23308_), .ZN(new_n23391_));
  OAI21_X1   g23094(.A1(new_n23308_), .A2(new_n23387_), .B(new_n23391_), .ZN(new_n23392_));
  OAI22_X1   g23095(.A1(new_n6644_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n6647_), .ZN(new_n23393_));
  OAI21_X1   g23096(.A1(new_n12542_), .A2(new_n7284_), .B(new_n23393_), .ZN(new_n23394_));
  AOI21_X1   g23097(.A1(new_n23394_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n23395_));
  XNOR2_X1   g23098(.A1(new_n13371_), .A2(new_n23395_), .ZN(new_n23396_));
  NAND2_X1   g23099(.A1(new_n23263_), .A2(new_n23274_), .ZN(new_n23397_));
  AOI21_X1   g23100(.A1(new_n23397_), .A2(new_n23273_), .B(new_n23396_), .ZN(new_n23398_));
  INV_X1     g23101(.I(new_n23396_), .ZN(new_n23399_));
  NAND2_X1   g23102(.A1(new_n23397_), .A2(new_n23273_), .ZN(new_n23400_));
  NOR2_X1    g23103(.A1(new_n23400_), .A2(new_n23399_), .ZN(new_n23401_));
  OAI21_X1   g23104(.A1(new_n23401_), .A2(new_n23398_), .B(new_n23392_), .ZN(new_n23402_));
  XOR2_X1    g23105(.A1(new_n23400_), .A2(new_n23396_), .Z(new_n23403_));
  OAI21_X1   g23106(.A1(new_n23403_), .A2(new_n23392_), .B(new_n23402_), .ZN(new_n23404_));
  XOR2_X1    g23107(.A1(new_n23404_), .A2(new_n23306_), .Z(new_n23405_));
  NOR2_X1    g23108(.A1(new_n23405_), .A2(new_n23303_), .ZN(new_n23406_));
  INV_X1     g23109(.I(new_n23303_), .ZN(new_n23407_));
  AND2_X2    g23110(.A1(new_n23404_), .A2(new_n23305_), .Z(new_n23408_));
  NOR2_X1    g23111(.A1(new_n23404_), .A2(new_n23305_), .ZN(new_n23409_));
  NOR2_X1    g23112(.A1(new_n23408_), .A2(new_n23409_), .ZN(new_n23410_));
  NOR2_X1    g23113(.A1(new_n23410_), .A2(new_n23407_), .ZN(new_n23411_));
  NOR2_X1    g23114(.A1(new_n23411_), .A2(new_n23406_), .ZN(new_n23412_));
  INV_X1     g23115(.I(new_n23287_), .ZN(new_n23413_));
  NOR2_X1    g23116(.A1(new_n23413_), .A2(new_n23284_), .ZN(new_n23414_));
  XOR2_X1    g23117(.A1(new_n23285_), .A2(new_n4860_), .Z(new_n23415_));
  AOI21_X1   g23118(.A1(new_n23413_), .A2(new_n23284_), .B(new_n23415_), .ZN(new_n23416_));
  NOR2_X1    g23119(.A1(new_n23416_), .A2(new_n23414_), .ZN(new_n23417_));
  XOR2_X1    g23120(.A1(new_n23412_), .A2(new_n23417_), .Z(new_n23418_));
  INV_X1     g23121(.I(new_n23418_), .ZN(new_n23419_));
  NAND2_X1   g23122(.A1(new_n23294_), .A2(new_n23419_), .ZN(new_n23420_));
  XOR2_X1    g23123(.A1(new_n23420_), .A2(new_n23299_), .Z(new_n23421_));
  XOR2_X1    g23124(.A1(new_n23176_), .A2(new_n23421_), .Z(\f[102] ));
  NOR3_X1    g23125(.A1(new_n23412_), .A2(new_n23414_), .A3(new_n23416_), .ZN(new_n23423_));
  INV_X1     g23126(.I(new_n23423_), .ZN(new_n23424_));
  INV_X1     g23127(.I(new_n23034_), .ZN(new_n23425_));
  NOR3_X1    g23128(.A1(new_n22884_), .A2(new_n23425_), .A3(new_n23173_), .ZN(new_n23426_));
  NOR2_X1    g23129(.A1(new_n23298_), .A2(new_n23419_), .ZN(new_n23427_));
  AOI21_X1   g23130(.A1(new_n23298_), .A2(new_n23419_), .B(new_n23177_), .ZN(new_n23428_));
  NOR2_X1    g23131(.A1(new_n23428_), .A2(new_n23427_), .ZN(new_n23429_));
  OAI21_X1   g23132(.A1(new_n23426_), .A2(new_n23171_), .B(new_n23429_), .ZN(new_n23430_));
  NOR2_X1    g23133(.A1(new_n5997_), .A2(new_n5991_), .ZN(new_n23431_));
  NAND2_X1   g23134(.A1(new_n16148_), .A2(new_n5681_), .ZN(new_n23432_));
  OAI21_X1   g23135(.A1(new_n23431_), .A2(new_n23432_), .B(new_n5680_), .ZN(new_n23433_));
  XNOR2_X1   g23136(.A1(new_n14978_), .A2(new_n23433_), .ZN(new_n23434_));
  NOR2_X1    g23137(.A1(new_n23401_), .A2(new_n23392_), .ZN(new_n23435_));
  OAI22_X1   g23138(.A1(new_n7619_), .A2(new_n12536_), .B1(new_n12542_), .B2(new_n8309_), .ZN(new_n23436_));
  OAI21_X1   g23139(.A1(new_n11744_), .A2(new_n7947_), .B(new_n23436_), .ZN(new_n23437_));
  AOI21_X1   g23140(.A1(new_n23437_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23438_));
  XNOR2_X1   g23141(.A1(new_n12546_), .A2(new_n23438_), .ZN(new_n23439_));
  INV_X1     g23142(.I(new_n10032_), .ZN(new_n23440_));
  AOI22_X1   g23143(.A1(new_n11415_), .A2(new_n23440_), .B1(\b[50] ), .B2(new_n10145_), .ZN(new_n23441_));
  OAI21_X1   g23144(.A1(new_n23441_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23442_));
  XOR2_X1    g23145(.A1(new_n10035_), .A2(new_n23442_), .Z(new_n23443_));
  OAI21_X1   g23146(.A1(new_n23318_), .A2(new_n23334_), .B(new_n23336_), .ZN(new_n23444_));
  AOI22_X1   g23147(.A1(new_n13078_), .A2(\b[44] ), .B1(new_n22614_), .B2(new_n12218_), .ZN(new_n23445_));
  OAI21_X1   g23148(.A1(new_n23445_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23446_));
  XOR2_X1    g23149(.A1(new_n7874_), .A2(new_n23446_), .Z(new_n23447_));
  OAI22_X1   g23150(.A1(new_n13880_), .A2(new_n7193_), .B1(new_n6229_), .B2(new_n13885_), .ZN(new_n23448_));
  AOI21_X1   g23151(.A1(new_n23448_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23449_));
  XNOR2_X1   g23152(.A1(new_n6851_), .A2(new_n23449_), .ZN(new_n23450_));
  NAND2_X1   g23153(.A1(new_n23331_), .A2(new_n23068_), .ZN(new_n23451_));
  NAND2_X1   g23154(.A1(new_n23451_), .A2(new_n23330_), .ZN(new_n23452_));
  NOR2_X1    g23155(.A1(new_n13476_), .A2(new_n5913_), .ZN(new_n23453_));
  XOR2_X1    g23156(.A1(new_n14736_), .A2(new_n5913_), .Z(new_n23454_));
  NAND2_X1   g23157(.A1(new_n23454_), .A2(\b[40] ), .ZN(new_n23455_));
  XOR2_X1    g23158(.A1(new_n23455_), .A2(new_n23453_), .Z(new_n23456_));
  INV_X1     g23159(.I(new_n23456_), .ZN(new_n23457_));
  XOR2_X1    g23160(.A1(new_n23452_), .A2(new_n23457_), .Z(new_n23458_));
  INV_X1     g23161(.I(new_n23458_), .ZN(new_n23459_));
  NOR2_X1    g23162(.A1(new_n23452_), .A2(new_n23456_), .ZN(new_n23460_));
  INV_X1     g23163(.I(new_n23460_), .ZN(new_n23461_));
  NAND2_X1   g23164(.A1(new_n23452_), .A2(new_n23456_), .ZN(new_n23462_));
  AOI21_X1   g23165(.A1(new_n23461_), .A2(new_n23462_), .B(new_n23450_), .ZN(new_n23463_));
  AOI21_X1   g23166(.A1(new_n23450_), .A2(new_n23459_), .B(new_n23463_), .ZN(new_n23464_));
  INV_X1     g23167(.I(new_n23464_), .ZN(new_n23465_));
  AND2_X2    g23168(.A1(new_n23447_), .A2(new_n23465_), .Z(new_n23466_));
  NOR2_X1    g23169(.A1(new_n23447_), .A2(new_n23465_), .ZN(new_n23467_));
  OAI21_X1   g23170(.A1(new_n23466_), .A2(new_n23467_), .B(new_n23444_), .ZN(new_n23468_));
  XOR2_X1    g23171(.A1(new_n23447_), .A2(new_n23464_), .Z(new_n23469_));
  OAI21_X1   g23172(.A1(new_n23444_), .A2(new_n23469_), .B(new_n23468_), .ZN(new_n23470_));
  INV_X1     g23173(.I(new_n23470_), .ZN(new_n23471_));
  NAND2_X1   g23174(.A1(new_n23351_), .A2(new_n23353_), .ZN(new_n23472_));
  NAND2_X1   g23175(.A1(new_n23472_), .A2(new_n23347_), .ZN(new_n23473_));
  INV_X1     g23176(.I(new_n23473_), .ZN(new_n23474_));
  AOI22_X1   g23177(.A1(new_n10969_), .A2(new_n9291_), .B1(new_n11394_), .B2(\b[47] ), .ZN(new_n23475_));
  OAI21_X1   g23178(.A1(new_n23475_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n23476_));
  XNOR2_X1   g23179(.A1(new_n8952_), .A2(new_n23476_), .ZN(new_n23477_));
  NOR2_X1    g23180(.A1(new_n23474_), .A2(new_n23477_), .ZN(new_n23478_));
  INV_X1     g23181(.I(new_n23477_), .ZN(new_n23479_));
  NOR2_X1    g23182(.A1(new_n23473_), .A2(new_n23479_), .ZN(new_n23480_));
  NOR2_X1    g23183(.A1(new_n23478_), .A2(new_n23480_), .ZN(new_n23481_));
  NOR2_X1    g23184(.A1(new_n23481_), .A2(new_n23471_), .ZN(new_n23482_));
  XOR2_X1    g23185(.A1(new_n23473_), .A2(new_n23477_), .Z(new_n23483_));
  NOR2_X1    g23186(.A1(new_n23483_), .A2(new_n23470_), .ZN(new_n23484_));
  NOR2_X1    g23187(.A1(new_n23482_), .A2(new_n23484_), .ZN(new_n23485_));
  OAI21_X1   g23188(.A1(new_n23356_), .A2(new_n23365_), .B(new_n23363_), .ZN(new_n23486_));
  INV_X1     g23189(.I(new_n23486_), .ZN(new_n23487_));
  NOR2_X1    g23190(.A1(new_n23485_), .A2(new_n23487_), .ZN(new_n23488_));
  NOR3_X1    g23191(.A1(new_n23482_), .A2(new_n23484_), .A3(new_n23486_), .ZN(new_n23489_));
  NOR2_X1    g23192(.A1(new_n23488_), .A2(new_n23489_), .ZN(new_n23490_));
  NOR2_X1    g23193(.A1(new_n23490_), .A2(new_n23443_), .ZN(new_n23491_));
  INV_X1     g23194(.I(new_n23443_), .ZN(new_n23492_));
  XOR2_X1    g23195(.A1(new_n23485_), .A2(new_n23486_), .Z(new_n23493_));
  NOR2_X1    g23196(.A1(new_n23493_), .A2(new_n23492_), .ZN(new_n23494_));
  NOR2_X1    g23197(.A1(new_n23375_), .A2(new_n23315_), .ZN(new_n23495_));
  NOR2_X1    g23198(.A1(new_n23495_), .A2(new_n23373_), .ZN(new_n23496_));
  OAI22_X1   g23199(.A1(new_n8644_), .A2(new_n10862_), .B1(new_n11738_), .B2(new_n9388_), .ZN(new_n23497_));
  OAI21_X1   g23200(.A1(new_n10477_), .A2(new_n10154_), .B(new_n23497_), .ZN(new_n23498_));
  AOI21_X1   g23201(.A1(new_n23498_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n23499_));
  XOR2_X1    g23202(.A1(new_n11298_), .A2(new_n23499_), .Z(new_n23500_));
  NOR2_X1    g23203(.A1(new_n23496_), .A2(new_n23500_), .ZN(new_n23501_));
  AND2_X2    g23204(.A1(new_n23496_), .A2(new_n23500_), .Z(new_n23502_));
  OAI22_X1   g23205(.A1(new_n23502_), .A2(new_n23501_), .B1(new_n23491_), .B2(new_n23494_), .ZN(new_n23503_));
  NOR2_X1    g23206(.A1(new_n23494_), .A2(new_n23491_), .ZN(new_n23504_));
  XOR2_X1    g23207(.A1(new_n23496_), .A2(new_n23500_), .Z(new_n23505_));
  NAND2_X1   g23208(.A1(new_n23505_), .A2(new_n23504_), .ZN(new_n23506_));
  NAND2_X1   g23209(.A1(new_n23506_), .A2(new_n23503_), .ZN(new_n23507_));
  INV_X1     g23210(.I(new_n23507_), .ZN(new_n23508_));
  NOR2_X1    g23211(.A1(new_n23379_), .A2(new_n23309_), .ZN(new_n23509_));
  NOR2_X1    g23212(.A1(new_n23509_), .A2(new_n23380_), .ZN(new_n23510_));
  NOR2_X1    g23213(.A1(new_n23508_), .A2(new_n23510_), .ZN(new_n23511_));
  INV_X1     g23214(.I(new_n23511_), .ZN(new_n23512_));
  NAND2_X1   g23215(.A1(new_n23508_), .A2(new_n23510_), .ZN(new_n23513_));
  AOI21_X1   g23216(.A1(new_n23512_), .A2(new_n23513_), .B(new_n23439_), .ZN(new_n23514_));
  INV_X1     g23217(.I(new_n23439_), .ZN(new_n23515_));
  XOR2_X1    g23218(.A1(new_n23507_), .A2(new_n23510_), .Z(new_n23516_));
  NOR2_X1    g23219(.A1(new_n23516_), .A2(new_n23515_), .ZN(new_n23517_));
  NOR2_X1    g23220(.A1(new_n23514_), .A2(new_n23517_), .ZN(new_n23518_));
  AOI21_X1   g23221(.A1(new_n23307_), .A2(new_n23389_), .B(new_n23388_), .ZN(new_n23519_));
  OAI22_X1   g23222(.A1(new_n6644_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n6647_), .ZN(new_n23520_));
  OAI21_X1   g23223(.A1(new_n12970_), .A2(new_n7284_), .B(new_n23520_), .ZN(new_n23521_));
  AOI21_X1   g23224(.A1(new_n23521_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n23522_));
  XOR2_X1    g23225(.A1(new_n13784_), .A2(new_n23522_), .Z(new_n23523_));
  XNOR2_X1   g23226(.A1(new_n23519_), .A2(new_n23523_), .ZN(new_n23524_));
  NOR2_X1    g23227(.A1(new_n23524_), .A2(new_n23518_), .ZN(new_n23525_));
  INV_X1     g23228(.I(new_n23518_), .ZN(new_n23526_));
  NOR2_X1    g23229(.A1(new_n23519_), .A2(new_n23523_), .ZN(new_n23527_));
  INV_X1     g23230(.I(new_n23527_), .ZN(new_n23528_));
  NAND2_X1   g23231(.A1(new_n23519_), .A2(new_n23523_), .ZN(new_n23529_));
  AOI21_X1   g23232(.A1(new_n23529_), .A2(new_n23528_), .B(new_n23526_), .ZN(new_n23530_));
  NOR2_X1    g23233(.A1(new_n23530_), .A2(new_n23525_), .ZN(new_n23531_));
  NOR3_X1    g23234(.A1(new_n23531_), .A2(new_n23398_), .A3(new_n23435_), .ZN(new_n23532_));
  NOR2_X1    g23235(.A1(new_n23435_), .A2(new_n23398_), .ZN(new_n23533_));
  INV_X1     g23236(.I(new_n23531_), .ZN(new_n23534_));
  NOR2_X1    g23237(.A1(new_n23534_), .A2(new_n23533_), .ZN(new_n23535_));
  NOR2_X1    g23238(.A1(new_n23535_), .A2(new_n23532_), .ZN(new_n23536_));
  NOR2_X1    g23239(.A1(new_n23536_), .A2(new_n23434_), .ZN(new_n23537_));
  INV_X1     g23240(.I(new_n23434_), .ZN(new_n23538_));
  XOR2_X1    g23241(.A1(new_n23531_), .A2(new_n23533_), .Z(new_n23539_));
  NOR2_X1    g23242(.A1(new_n23539_), .A2(new_n23538_), .ZN(new_n23540_));
  NOR2_X1    g23243(.A1(new_n23537_), .A2(new_n23540_), .ZN(new_n23541_));
  INV_X1     g23244(.I(new_n23408_), .ZN(new_n23542_));
  AOI21_X1   g23245(.A1(new_n23542_), .A2(new_n23407_), .B(new_n23409_), .ZN(new_n23543_));
  NOR2_X1    g23246(.A1(new_n23541_), .A2(new_n23543_), .ZN(new_n23544_));
  XOR2_X1    g23247(.A1(new_n23430_), .A2(new_n23544_), .Z(new_n23545_));
  XOR2_X1    g23248(.A1(new_n23545_), .A2(new_n23424_), .Z(\f[103] ));
  NOR2_X1    g23249(.A1(new_n23424_), .A2(new_n23541_), .ZN(new_n23547_));
  INV_X1     g23250(.I(new_n23547_), .ZN(new_n23548_));
  AOI21_X1   g23251(.A1(new_n23424_), .A2(new_n23541_), .B(new_n23543_), .ZN(new_n23549_));
  INV_X1     g23252(.I(new_n23549_), .ZN(new_n23550_));
  OAI21_X1   g23253(.A1(new_n23430_), .A2(new_n23550_), .B(new_n23548_), .ZN(new_n23551_));
  INV_X1     g23254(.I(new_n23532_), .ZN(new_n23552_));
  AOI21_X1   g23255(.A1(new_n23552_), .A2(new_n23538_), .B(new_n23535_), .ZN(new_n23553_));
  OAI22_X1   g23256(.A1(new_n6644_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n6647_), .ZN(new_n23554_));
  OAI21_X1   g23257(.A1(new_n13367_), .A2(new_n7284_), .B(new_n23554_), .ZN(new_n23555_));
  AOI21_X1   g23258(.A1(new_n23555_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n23556_));
  XOR2_X1    g23259(.A1(new_n14213_), .A2(new_n23556_), .Z(new_n23557_));
  INV_X1     g23260(.I(new_n23557_), .ZN(new_n23558_));
  AOI22_X1   g23261(.A1(new_n8631_), .A2(\b[55] ), .B1(\b[56] ), .B2(new_n9382_), .ZN(new_n23559_));
  AOI21_X1   g23262(.A1(\b[54] ), .A2(new_n9731_), .B(new_n23559_), .ZN(new_n23560_));
  OAI21_X1   g23263(.A1(new_n23560_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n23561_));
  XOR2_X1    g23264(.A1(new_n11748_), .A2(new_n23561_), .Z(new_n23562_));
  INV_X1     g23265(.I(new_n23489_), .ZN(new_n23563_));
  AOI21_X1   g23266(.A1(new_n23563_), .A2(new_n23492_), .B(new_n23488_), .ZN(new_n23564_));
  AOI22_X1   g23267(.A1(new_n11415_), .A2(new_n10858_), .B1(\b[51] ), .B2(new_n10145_), .ZN(new_n23565_));
  OAI21_X1   g23268(.A1(new_n23565_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23566_));
  XNOR2_X1   g23269(.A1(new_n10476_), .A2(new_n23566_), .ZN(new_n23567_));
  OAI22_X1   g23270(.A1(new_n10979_), .A2(new_n9296_), .B1(new_n8563_), .B2(new_n11401_), .ZN(new_n23568_));
  AOI21_X1   g23271(.A1(new_n23568_), .A2(new_n10973_), .B(new_n10964_), .ZN(new_n23569_));
  XNOR2_X1   g23272(.A1(new_n9299_), .A2(new_n23569_), .ZN(new_n23570_));
  INV_X1     g23273(.I(new_n23444_), .ZN(new_n23571_));
  NOR2_X1    g23274(.A1(new_n23466_), .A2(new_n23571_), .ZN(new_n23572_));
  NOR2_X1    g23275(.A1(new_n23572_), .A2(new_n23467_), .ZN(new_n23573_));
  NAND2_X1   g23276(.A1(new_n23450_), .A2(new_n23461_), .ZN(new_n23574_));
  NAND2_X1   g23277(.A1(new_n23574_), .A2(new_n23462_), .ZN(new_n23575_));
  NOR2_X1    g23278(.A1(new_n13476_), .A2(new_n5921_), .ZN(new_n23576_));
  XOR2_X1    g23279(.A1(new_n14736_), .A2(new_n5921_), .Z(new_n23577_));
  NAND2_X1   g23280(.A1(new_n23577_), .A2(\b[41] ), .ZN(new_n23578_));
  XOR2_X1    g23281(.A1(new_n23578_), .A2(new_n23576_), .Z(new_n23579_));
  NOR2_X1    g23282(.A1(new_n23457_), .A2(new_n23579_), .ZN(new_n23580_));
  INV_X1     g23283(.I(new_n23579_), .ZN(new_n23581_));
  NOR2_X1    g23284(.A1(new_n23581_), .A2(new_n23456_), .ZN(new_n23582_));
  NOR2_X1    g23285(.A1(new_n23580_), .A2(new_n23582_), .ZN(new_n23583_));
  INV_X1     g23286(.I(new_n23583_), .ZN(new_n23584_));
  XOR2_X1    g23287(.A1(new_n23456_), .A2(new_n23579_), .Z(new_n23585_));
  NOR2_X1    g23288(.A1(new_n23575_), .A2(new_n23585_), .ZN(new_n23586_));
  AOI21_X1   g23289(.A1(new_n23575_), .A2(new_n23584_), .B(new_n23586_), .ZN(new_n23587_));
  AOI22_X1   g23290(.A1(new_n13078_), .A2(\b[45] ), .B1(new_n8557_), .B2(new_n12218_), .ZN(new_n23588_));
  OAI21_X1   g23291(.A1(new_n23588_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23589_));
  XNOR2_X1   g23292(.A1(new_n8217_), .A2(new_n23589_), .ZN(new_n23590_));
  OAI22_X1   g23293(.A1(new_n13880_), .A2(new_n7199_), .B1(new_n6538_), .B2(new_n13885_), .ZN(new_n23591_));
  AOI21_X1   g23294(.A1(new_n23591_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23592_));
  XNOR2_X1   g23295(.A1(new_n7202_), .A2(new_n23592_), .ZN(new_n23593_));
  XNOR2_X1   g23296(.A1(new_n23590_), .A2(new_n23593_), .ZN(new_n23594_));
  NOR2_X1    g23297(.A1(new_n23594_), .A2(new_n23587_), .ZN(new_n23595_));
  INV_X1     g23298(.I(new_n23587_), .ZN(new_n23596_));
  NOR2_X1    g23299(.A1(new_n23590_), .A2(new_n23593_), .ZN(new_n23597_));
  INV_X1     g23300(.I(new_n23597_), .ZN(new_n23598_));
  NAND2_X1   g23301(.A1(new_n23590_), .A2(new_n23593_), .ZN(new_n23599_));
  AOI21_X1   g23302(.A1(new_n23598_), .A2(new_n23599_), .B(new_n23596_), .ZN(new_n23600_));
  NOR2_X1    g23303(.A1(new_n23595_), .A2(new_n23600_), .ZN(new_n23601_));
  XOR2_X1    g23304(.A1(new_n23601_), .A2(new_n23573_), .Z(new_n23602_));
  NOR2_X1    g23305(.A1(new_n23602_), .A2(new_n23570_), .ZN(new_n23603_));
  INV_X1     g23306(.I(new_n23570_), .ZN(new_n23604_));
  INV_X1     g23307(.I(new_n23573_), .ZN(new_n23605_));
  NOR2_X1    g23308(.A1(new_n23605_), .A2(new_n23601_), .ZN(new_n23606_));
  INV_X1     g23309(.I(new_n23606_), .ZN(new_n23607_));
  NAND2_X1   g23310(.A1(new_n23605_), .A2(new_n23601_), .ZN(new_n23608_));
  AOI21_X1   g23311(.A1(new_n23607_), .A2(new_n23608_), .B(new_n23604_), .ZN(new_n23609_));
  NOR2_X1    g23312(.A1(new_n23603_), .A2(new_n23609_), .ZN(new_n23610_));
  NOR2_X1    g23313(.A1(new_n23480_), .A2(new_n23471_), .ZN(new_n23611_));
  NOR2_X1    g23314(.A1(new_n23611_), .A2(new_n23478_), .ZN(new_n23612_));
  XOR2_X1    g23315(.A1(new_n23610_), .A2(new_n23612_), .Z(new_n23613_));
  NOR2_X1    g23316(.A1(new_n23613_), .A2(new_n23567_), .ZN(new_n23614_));
  INV_X1     g23317(.I(new_n23567_), .ZN(new_n23615_));
  INV_X1     g23318(.I(new_n23610_), .ZN(new_n23616_));
  NOR2_X1    g23319(.A1(new_n23616_), .A2(new_n23612_), .ZN(new_n23617_));
  INV_X1     g23320(.I(new_n23617_), .ZN(new_n23618_));
  NAND2_X1   g23321(.A1(new_n23616_), .A2(new_n23612_), .ZN(new_n23619_));
  AOI21_X1   g23322(.A1(new_n23618_), .A2(new_n23619_), .B(new_n23615_), .ZN(new_n23620_));
  NOR2_X1    g23323(.A1(new_n23620_), .A2(new_n23614_), .ZN(new_n23621_));
  XOR2_X1    g23324(.A1(new_n23621_), .A2(new_n23564_), .Z(new_n23622_));
  INV_X1     g23325(.I(new_n23564_), .ZN(new_n23623_));
  NOR2_X1    g23326(.A1(new_n23621_), .A2(new_n23623_), .ZN(new_n23624_));
  NAND2_X1   g23327(.A1(new_n23621_), .A2(new_n23623_), .ZN(new_n23625_));
  INV_X1     g23328(.I(new_n23625_), .ZN(new_n23626_));
  OAI21_X1   g23329(.A1(new_n23626_), .A2(new_n23624_), .B(new_n23562_), .ZN(new_n23627_));
  OAI21_X1   g23330(.A1(new_n23562_), .A2(new_n23622_), .B(new_n23627_), .ZN(new_n23628_));
  OAI22_X1   g23331(.A1(new_n7619_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n8309_), .ZN(new_n23629_));
  OAI21_X1   g23332(.A1(new_n12536_), .A2(new_n7947_), .B(new_n23629_), .ZN(new_n23630_));
  AOI21_X1   g23333(.A1(new_n23630_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23631_));
  XOR2_X1    g23334(.A1(new_n12969_), .A2(new_n23631_), .Z(new_n23632_));
  NOR2_X1    g23335(.A1(new_n23504_), .A2(new_n23502_), .ZN(new_n23633_));
  NOR2_X1    g23336(.A1(new_n23633_), .A2(new_n23501_), .ZN(new_n23634_));
  XOR2_X1    g23337(.A1(new_n23634_), .A2(new_n23632_), .Z(new_n23635_));
  NOR2_X1    g23338(.A1(new_n23634_), .A2(new_n23632_), .ZN(new_n23636_));
  INV_X1     g23339(.I(new_n23636_), .ZN(new_n23637_));
  NAND2_X1   g23340(.A1(new_n23634_), .A2(new_n23632_), .ZN(new_n23638_));
  AOI21_X1   g23341(.A1(new_n23637_), .A2(new_n23638_), .B(new_n23628_), .ZN(new_n23639_));
  AOI21_X1   g23342(.A1(new_n23628_), .A2(new_n23635_), .B(new_n23639_), .ZN(new_n23640_));
  AOI21_X1   g23343(.A1(new_n23515_), .A2(new_n23513_), .B(new_n23511_), .ZN(new_n23641_));
  NOR2_X1    g23344(.A1(new_n23640_), .A2(new_n23641_), .ZN(new_n23642_));
  NAND2_X1   g23345(.A1(new_n23640_), .A2(new_n23641_), .ZN(new_n23643_));
  INV_X1     g23346(.I(new_n23643_), .ZN(new_n23644_));
  OAI21_X1   g23347(.A1(new_n23644_), .A2(new_n23642_), .B(new_n23558_), .ZN(new_n23645_));
  XNOR2_X1   g23348(.A1(new_n23640_), .A2(new_n23641_), .ZN(new_n23646_));
  OAI21_X1   g23349(.A1(new_n23558_), .A2(new_n23646_), .B(new_n23645_), .ZN(new_n23647_));
  OAI21_X1   g23350(.A1(new_n5993_), .A2(new_n5997_), .B(new_n16487_), .ZN(new_n23648_));
  NAND2_X1   g23351(.A1(new_n23526_), .A2(new_n23529_), .ZN(new_n23649_));
  NAND2_X1   g23352(.A1(new_n23649_), .A2(new_n23528_), .ZN(new_n23650_));
  XNOR2_X1   g23353(.A1(new_n23650_), .A2(new_n23648_), .ZN(new_n23651_));
  XOR2_X1    g23354(.A1(new_n23651_), .A2(new_n23647_), .Z(new_n23652_));
  NOR2_X1    g23355(.A1(new_n23652_), .A2(\a[41] ), .ZN(new_n23653_));
  NAND2_X1   g23356(.A1(new_n23652_), .A2(\a[41] ), .ZN(new_n23654_));
  INV_X1     g23357(.I(new_n23654_), .ZN(new_n23655_));
  NOR2_X1    g23358(.A1(new_n23655_), .A2(new_n23653_), .ZN(new_n23656_));
  XOR2_X1    g23359(.A1(new_n23656_), .A2(new_n23553_), .Z(new_n23657_));
  NAND2_X1   g23360(.A1(new_n23551_), .A2(new_n23657_), .ZN(new_n23658_));
  INV_X1     g23361(.I(new_n23429_), .ZN(new_n23659_));
  AOI21_X1   g23362(.A1(new_n23175_), .A2(new_n23172_), .B(new_n23659_), .ZN(new_n23660_));
  AOI21_X1   g23363(.A1(new_n23660_), .A2(new_n23549_), .B(new_n23547_), .ZN(new_n23661_));
  INV_X1     g23364(.I(new_n23553_), .ZN(new_n23662_));
  INV_X1     g23365(.I(new_n23656_), .ZN(new_n23663_));
  NAND2_X1   g23366(.A1(new_n23663_), .A2(new_n23662_), .ZN(new_n23664_));
  NAND2_X1   g23367(.A1(new_n23656_), .A2(new_n23553_), .ZN(new_n23665_));
  NAND2_X1   g23368(.A1(new_n23664_), .A2(new_n23665_), .ZN(new_n23666_));
  NAND2_X1   g23369(.A1(new_n23661_), .A2(new_n23666_), .ZN(new_n23667_));
  NAND2_X1   g23370(.A1(new_n23667_), .A2(new_n23658_), .ZN(\f[104] ));
  OAI22_X1   g23371(.A1(new_n6644_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n6647_), .ZN(new_n23669_));
  OAI21_X1   g23372(.A1(new_n13785_), .A2(new_n7284_), .B(new_n23669_), .ZN(new_n23670_));
  AOI21_X1   g23373(.A1(new_n23670_), .A2(new_n6632_), .B(new_n6644_), .ZN(new_n23671_));
  XNOR2_X1   g23374(.A1(new_n14599_), .A2(new_n23671_), .ZN(new_n23672_));
  NOR2_X1    g23375(.A1(new_n23644_), .A2(new_n23557_), .ZN(new_n23673_));
  NOR2_X1    g23376(.A1(new_n23673_), .A2(new_n23642_), .ZN(new_n23674_));
  OAI21_X1   g23377(.A1(new_n23562_), .A2(new_n23624_), .B(new_n23625_), .ZN(new_n23675_));
  OAI22_X1   g23378(.A1(new_n8644_), .A2(new_n11744_), .B1(new_n12536_), .B2(new_n9388_), .ZN(new_n23676_));
  OAI21_X1   g23379(.A1(new_n11738_), .A2(new_n10154_), .B(new_n23676_), .ZN(new_n23677_));
  AOI21_X1   g23380(.A1(new_n23677_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n23678_));
  XNOR2_X1   g23381(.A1(new_n12128_), .A2(new_n23678_), .ZN(new_n23679_));
  AOI21_X1   g23382(.A1(new_n23615_), .A2(new_n23619_), .B(new_n23617_), .ZN(new_n23680_));
  OAI21_X1   g23383(.A1(new_n23570_), .A2(new_n23606_), .B(new_n23608_), .ZN(new_n23681_));
  AOI22_X1   g23384(.A1(new_n10969_), .A2(new_n10027_), .B1(new_n11394_), .B2(\b[49] ), .ZN(new_n23682_));
  OAI21_X1   g23385(.A1(new_n23682_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n23683_));
  XOR2_X1    g23386(.A1(new_n9642_), .A2(new_n23683_), .Z(new_n23684_));
  INV_X1     g23387(.I(new_n23684_), .ZN(new_n23685_));
  INV_X1     g23388(.I(new_n23582_), .ZN(new_n23686_));
  AOI21_X1   g23389(.A1(new_n23575_), .A2(new_n23686_), .B(new_n23580_), .ZN(new_n23687_));
  OAI22_X1   g23390(.A1(new_n13880_), .A2(new_n7865_), .B1(new_n6847_), .B2(new_n13885_), .ZN(new_n23688_));
  AOI21_X1   g23391(.A1(new_n23688_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23689_));
  XOR2_X1    g23392(.A1(new_n7516_), .A2(new_n23689_), .Z(new_n23690_));
  NOR2_X1    g23393(.A1(new_n13476_), .A2(new_n6229_), .ZN(new_n23691_));
  XOR2_X1    g23394(.A1(new_n14736_), .A2(new_n6229_), .Z(new_n23692_));
  NAND2_X1   g23395(.A1(new_n23692_), .A2(\b[42] ), .ZN(new_n23693_));
  XOR2_X1    g23396(.A1(new_n23693_), .A2(new_n23691_), .Z(new_n23694_));
  XOR2_X1    g23397(.A1(new_n23694_), .A2(\a[41] ), .Z(new_n23695_));
  NOR2_X1    g23398(.A1(new_n23695_), .A2(new_n23456_), .ZN(new_n23696_));
  NOR2_X1    g23399(.A1(new_n23694_), .A2(new_n5681_), .ZN(new_n23697_));
  INV_X1     g23400(.I(new_n23697_), .ZN(new_n23698_));
  NAND2_X1   g23401(.A1(new_n23694_), .A2(new_n5681_), .ZN(new_n23699_));
  AOI21_X1   g23402(.A1(new_n23698_), .A2(new_n23699_), .B(new_n23457_), .ZN(new_n23700_));
  NOR2_X1    g23403(.A1(new_n23696_), .A2(new_n23700_), .ZN(new_n23701_));
  XOR2_X1    g23404(.A1(new_n23690_), .A2(new_n23701_), .Z(new_n23702_));
  NOR2_X1    g23405(.A1(new_n23702_), .A2(new_n23687_), .ZN(new_n23703_));
  INV_X1     g23406(.I(new_n23687_), .ZN(new_n23704_));
  INV_X1     g23407(.I(new_n23690_), .ZN(new_n23705_));
  NOR2_X1    g23408(.A1(new_n23705_), .A2(new_n23701_), .ZN(new_n23706_));
  INV_X1     g23409(.I(new_n23706_), .ZN(new_n23707_));
  NAND2_X1   g23410(.A1(new_n23705_), .A2(new_n23701_), .ZN(new_n23708_));
  AOI21_X1   g23411(.A1(new_n23707_), .A2(new_n23708_), .B(new_n23704_), .ZN(new_n23709_));
  AOI22_X1   g23412(.A1(new_n13078_), .A2(\b[46] ), .B1(new_n8565_), .B2(new_n12218_), .ZN(new_n23710_));
  OAI21_X1   g23413(.A1(new_n23710_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23711_));
  XNOR2_X1   g23414(.A1(new_n8568_), .A2(new_n23711_), .ZN(new_n23712_));
  NAND2_X1   g23415(.A1(new_n23596_), .A2(new_n23599_), .ZN(new_n23713_));
  NAND2_X1   g23416(.A1(new_n23713_), .A2(new_n23598_), .ZN(new_n23714_));
  INV_X1     g23417(.I(new_n23714_), .ZN(new_n23715_));
  NOR2_X1    g23418(.A1(new_n23715_), .A2(new_n23712_), .ZN(new_n23716_));
  INV_X1     g23419(.I(new_n23712_), .ZN(new_n23717_));
  NOR2_X1    g23420(.A1(new_n23717_), .A2(new_n23714_), .ZN(new_n23718_));
  OAI22_X1   g23421(.A1(new_n23718_), .A2(new_n23716_), .B1(new_n23703_), .B2(new_n23709_), .ZN(new_n23719_));
  NOR2_X1    g23422(.A1(new_n23709_), .A2(new_n23703_), .ZN(new_n23720_));
  XNOR2_X1   g23423(.A1(new_n23712_), .A2(new_n23714_), .ZN(new_n23721_));
  NAND2_X1   g23424(.A1(new_n23721_), .A2(new_n23720_), .ZN(new_n23722_));
  AOI21_X1   g23425(.A1(new_n23722_), .A2(new_n23719_), .B(new_n23685_), .ZN(new_n23723_));
  INV_X1     g23426(.I(new_n23723_), .ZN(new_n23724_));
  NAND2_X1   g23427(.A1(new_n23722_), .A2(new_n23719_), .ZN(new_n23725_));
  NOR2_X1    g23428(.A1(new_n23725_), .A2(new_n23684_), .ZN(new_n23726_));
  INV_X1     g23429(.I(new_n23726_), .ZN(new_n23727_));
  NAND2_X1   g23430(.A1(new_n23727_), .A2(new_n23724_), .ZN(new_n23728_));
  XOR2_X1    g23431(.A1(new_n23725_), .A2(new_n23685_), .Z(new_n23729_));
  NOR2_X1    g23432(.A1(new_n23729_), .A2(new_n23681_), .ZN(new_n23730_));
  AOI21_X1   g23433(.A1(new_n23681_), .A2(new_n23728_), .B(new_n23730_), .ZN(new_n23731_));
  INV_X1     g23434(.I(new_n10863_), .ZN(new_n23732_));
  AOI22_X1   g23435(.A1(new_n11415_), .A2(new_n23732_), .B1(\b[52] ), .B2(new_n10145_), .ZN(new_n23733_));
  OAI21_X1   g23436(.A1(new_n23733_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23734_));
  XOR2_X1    g23437(.A1(new_n10866_), .A2(new_n23734_), .Z(new_n23735_));
  XNOR2_X1   g23438(.A1(new_n23731_), .A2(new_n23735_), .ZN(new_n23736_));
  NOR2_X1    g23439(.A1(new_n23736_), .A2(new_n23680_), .ZN(new_n23737_));
  INV_X1     g23440(.I(new_n23680_), .ZN(new_n23738_));
  NOR2_X1    g23441(.A1(new_n23731_), .A2(new_n23735_), .ZN(new_n23739_));
  INV_X1     g23442(.I(new_n23739_), .ZN(new_n23740_));
  NAND2_X1   g23443(.A1(new_n23731_), .A2(new_n23735_), .ZN(new_n23741_));
  AOI21_X1   g23444(.A1(new_n23740_), .A2(new_n23741_), .B(new_n23738_), .ZN(new_n23742_));
  NOR2_X1    g23445(.A1(new_n23737_), .A2(new_n23742_), .ZN(new_n23743_));
  XOR2_X1    g23446(.A1(new_n23743_), .A2(new_n23679_), .Z(new_n23744_));
  INV_X1     g23447(.I(new_n23744_), .ZN(new_n23745_));
  INV_X1     g23448(.I(new_n23679_), .ZN(new_n23746_));
  NOR2_X1    g23449(.A1(new_n23743_), .A2(new_n23746_), .ZN(new_n23747_));
  INV_X1     g23450(.I(new_n23747_), .ZN(new_n23748_));
  NAND2_X1   g23451(.A1(new_n23743_), .A2(new_n23746_), .ZN(new_n23749_));
  AOI21_X1   g23452(.A1(new_n23748_), .A2(new_n23749_), .B(new_n23675_), .ZN(new_n23750_));
  AOI21_X1   g23453(.A1(new_n23745_), .A2(new_n23675_), .B(new_n23750_), .ZN(new_n23751_));
  OAI22_X1   g23454(.A1(new_n7619_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n8309_), .ZN(new_n23752_));
  OAI21_X1   g23455(.A1(new_n12542_), .A2(new_n7947_), .B(new_n23752_), .ZN(new_n23753_));
  AOI21_X1   g23456(.A1(new_n23753_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23754_));
  XNOR2_X1   g23457(.A1(new_n13371_), .A2(new_n23754_), .ZN(new_n23755_));
  INV_X1     g23458(.I(new_n23628_), .ZN(new_n23756_));
  AOI21_X1   g23459(.A1(new_n23756_), .A2(new_n23638_), .B(new_n23636_), .ZN(new_n23757_));
  NOR2_X1    g23460(.A1(new_n23757_), .A2(new_n23755_), .ZN(new_n23758_));
  INV_X1     g23461(.I(new_n23758_), .ZN(new_n23759_));
  NAND2_X1   g23462(.A1(new_n23757_), .A2(new_n23755_), .ZN(new_n23760_));
  AOI21_X1   g23463(.A1(new_n23759_), .A2(new_n23760_), .B(new_n23751_), .ZN(new_n23761_));
  XOR2_X1    g23464(.A1(new_n23757_), .A2(new_n23755_), .Z(new_n23762_));
  AOI21_X1   g23465(.A1(new_n23751_), .A2(new_n23762_), .B(new_n23761_), .ZN(new_n23763_));
  XOR2_X1    g23466(.A1(new_n23763_), .A2(new_n23674_), .Z(new_n23764_));
  NOR2_X1    g23467(.A1(new_n23764_), .A2(new_n23672_), .ZN(new_n23765_));
  INV_X1     g23468(.I(new_n23674_), .ZN(new_n23766_));
  NOR2_X1    g23469(.A1(new_n23766_), .A2(new_n23763_), .ZN(new_n23767_));
  INV_X1     g23470(.I(new_n23767_), .ZN(new_n23768_));
  NAND2_X1   g23471(.A1(new_n23766_), .A2(new_n23763_), .ZN(new_n23769_));
  NAND2_X1   g23472(.A1(new_n23768_), .A2(new_n23769_), .ZN(new_n23770_));
  AOI21_X1   g23473(.A1(new_n23672_), .A2(new_n23770_), .B(new_n23765_), .ZN(new_n23771_));
  NAND2_X1   g23474(.A1(new_n23647_), .A2(new_n23650_), .ZN(new_n23772_));
  XOR2_X1    g23475(.A1(new_n23648_), .A2(\a[41] ), .Z(new_n23773_));
  OAI21_X1   g23476(.A1(new_n23647_), .A2(new_n23650_), .B(new_n23773_), .ZN(new_n23774_));
  NAND2_X1   g23477(.A1(new_n23774_), .A2(new_n23772_), .ZN(new_n23775_));
  INV_X1     g23478(.I(new_n23775_), .ZN(new_n23776_));
  XOR2_X1    g23479(.A1(new_n23771_), .A2(new_n23776_), .Z(new_n23777_));
  INV_X1     g23480(.I(new_n23777_), .ZN(new_n23778_));
  NAND2_X1   g23481(.A1(new_n23657_), .A2(new_n23778_), .ZN(new_n23779_));
  XOR2_X1    g23482(.A1(new_n23779_), .A2(new_n23664_), .Z(new_n23780_));
  XOR2_X1    g23483(.A1(new_n23551_), .A2(new_n23780_), .Z(\f[105] ));
  NOR2_X1    g23484(.A1(new_n23771_), .A2(new_n23775_), .ZN(new_n23782_));
  NOR2_X1    g23485(.A1(new_n23778_), .A2(new_n23663_), .ZN(new_n23783_));
  AOI21_X1   g23486(.A1(new_n23778_), .A2(new_n23663_), .B(new_n23662_), .ZN(new_n23784_));
  NOR2_X1    g23487(.A1(new_n23784_), .A2(new_n23783_), .ZN(new_n23785_));
  NAND2_X1   g23488(.A1(new_n23551_), .A2(new_n23785_), .ZN(new_n23786_));
  NOR2_X1    g23489(.A1(new_n7284_), .A2(new_n6647_), .ZN(new_n23787_));
  NAND2_X1   g23490(.A1(new_n16148_), .A2(new_n6632_), .ZN(new_n23788_));
  OAI21_X1   g23491(.A1(new_n23787_), .A2(new_n23788_), .B(new_n6631_), .ZN(new_n23789_));
  XNOR2_X1   g23492(.A1(new_n14978_), .A2(new_n23789_), .ZN(new_n23790_));
  AOI21_X1   g23493(.A1(new_n23751_), .A2(new_n23760_), .B(new_n23758_), .ZN(new_n23791_));
  OAI22_X1   g23494(.A1(new_n7619_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n8309_), .ZN(new_n23792_));
  OAI21_X1   g23495(.A1(new_n12970_), .A2(new_n7947_), .B(new_n23792_), .ZN(new_n23793_));
  AOI21_X1   g23496(.A1(new_n23793_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23794_));
  XOR2_X1    g23497(.A1(new_n13784_), .A2(new_n23794_), .Z(new_n23795_));
  INV_X1     g23498(.I(new_n23795_), .ZN(new_n23796_));
  INV_X1     g23499(.I(new_n23749_), .ZN(new_n23797_));
  AOI21_X1   g23500(.A1(new_n23675_), .A2(new_n23748_), .B(new_n23797_), .ZN(new_n23798_));
  INV_X1     g23501(.I(new_n23798_), .ZN(new_n23799_));
  AOI22_X1   g23502(.A1(new_n8631_), .A2(\b[57] ), .B1(\b[58] ), .B2(new_n9382_), .ZN(new_n23800_));
  AOI21_X1   g23503(.A1(\b[56] ), .A2(new_n9731_), .B(new_n23800_), .ZN(new_n23801_));
  OAI21_X1   g23504(.A1(new_n23801_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n23802_));
  XOR2_X1    g23505(.A1(new_n12546_), .A2(new_n23802_), .Z(new_n23803_));
  NAND2_X1   g23506(.A1(new_n23741_), .A2(new_n23738_), .ZN(new_n23804_));
  NAND2_X1   g23507(.A1(new_n23804_), .A2(new_n23740_), .ZN(new_n23805_));
  OAI22_X1   g23508(.A1(new_n10979_), .A2(new_n10032_), .B1(new_n9295_), .B2(new_n11401_), .ZN(new_n23806_));
  AOI21_X1   g23509(.A1(new_n23806_), .A2(new_n10973_), .B(new_n10964_), .ZN(new_n23807_));
  XNOR2_X1   g23510(.A1(new_n10035_), .A2(new_n23807_), .ZN(new_n23808_));
  OAI21_X1   g23511(.A1(new_n23687_), .A2(new_n23706_), .B(new_n23708_), .ZN(new_n23809_));
  INV_X1     g23512(.I(new_n23809_), .ZN(new_n23810_));
  OAI22_X1   g23513(.A1(new_n13880_), .A2(new_n7871_), .B1(new_n7198_), .B2(new_n13885_), .ZN(new_n23811_));
  AOI21_X1   g23514(.A1(new_n23811_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23812_));
  XNOR2_X1   g23515(.A1(new_n7874_), .A2(new_n23812_), .ZN(new_n23813_));
  NAND2_X1   g23516(.A1(new_n23699_), .A2(new_n23457_), .ZN(new_n23814_));
  NAND2_X1   g23517(.A1(new_n23814_), .A2(new_n23698_), .ZN(new_n23815_));
  NOR2_X1    g23518(.A1(new_n13476_), .A2(new_n6538_), .ZN(new_n23816_));
  XOR2_X1    g23519(.A1(new_n14736_), .A2(new_n6538_), .Z(new_n23817_));
  NAND2_X1   g23520(.A1(new_n23817_), .A2(\b[43] ), .ZN(new_n23818_));
  XOR2_X1    g23521(.A1(new_n23818_), .A2(new_n23816_), .Z(new_n23819_));
  INV_X1     g23522(.I(new_n23819_), .ZN(new_n23820_));
  XOR2_X1    g23523(.A1(new_n23815_), .A2(new_n23820_), .Z(new_n23821_));
  NOR2_X1    g23524(.A1(new_n23813_), .A2(new_n23821_), .ZN(new_n23822_));
  INV_X1     g23525(.I(new_n23813_), .ZN(new_n23823_));
  NOR2_X1    g23526(.A1(new_n23815_), .A2(new_n23819_), .ZN(new_n23824_));
  INV_X1     g23527(.I(new_n23824_), .ZN(new_n23825_));
  NAND2_X1   g23528(.A1(new_n23815_), .A2(new_n23819_), .ZN(new_n23826_));
  AOI21_X1   g23529(.A1(new_n23825_), .A2(new_n23826_), .B(new_n23823_), .ZN(new_n23827_));
  NOR2_X1    g23530(.A1(new_n23827_), .A2(new_n23822_), .ZN(new_n23828_));
  INV_X1     g23531(.I(new_n23828_), .ZN(new_n23829_));
  AOI22_X1   g23532(.A1(new_n13078_), .A2(\b[47] ), .B1(new_n9291_), .B2(new_n12218_), .ZN(new_n23830_));
  OAI21_X1   g23533(.A1(new_n23830_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23831_));
  XNOR2_X1   g23534(.A1(new_n8952_), .A2(new_n23831_), .ZN(new_n23832_));
  NOR2_X1    g23535(.A1(new_n23829_), .A2(new_n23832_), .ZN(new_n23833_));
  INV_X1     g23536(.I(new_n23832_), .ZN(new_n23834_));
  NOR2_X1    g23537(.A1(new_n23828_), .A2(new_n23834_), .ZN(new_n23835_));
  NOR2_X1    g23538(.A1(new_n23833_), .A2(new_n23835_), .ZN(new_n23836_));
  NOR2_X1    g23539(.A1(new_n23836_), .A2(new_n23810_), .ZN(new_n23837_));
  XOR2_X1    g23540(.A1(new_n23828_), .A2(new_n23832_), .Z(new_n23838_));
  NOR2_X1    g23541(.A1(new_n23838_), .A2(new_n23809_), .ZN(new_n23839_));
  NOR2_X1    g23542(.A1(new_n23837_), .A2(new_n23839_), .ZN(new_n23840_));
  INV_X1     g23543(.I(new_n23716_), .ZN(new_n23841_));
  OAI21_X1   g23544(.A1(new_n23717_), .A2(new_n23714_), .B(new_n23720_), .ZN(new_n23842_));
  NAND2_X1   g23545(.A1(new_n23841_), .A2(new_n23842_), .ZN(new_n23843_));
  INV_X1     g23546(.I(new_n23843_), .ZN(new_n23844_));
  NOR2_X1    g23547(.A1(new_n23840_), .A2(new_n23844_), .ZN(new_n23845_));
  NOR3_X1    g23548(.A1(new_n23837_), .A2(new_n23839_), .A3(new_n23843_), .ZN(new_n23846_));
  NOR2_X1    g23549(.A1(new_n23845_), .A2(new_n23846_), .ZN(new_n23847_));
  NOR2_X1    g23550(.A1(new_n23847_), .A2(new_n23808_), .ZN(new_n23848_));
  INV_X1     g23551(.I(new_n23808_), .ZN(new_n23849_));
  XOR2_X1    g23552(.A1(new_n23840_), .A2(new_n23843_), .Z(new_n23850_));
  NOR2_X1    g23553(.A1(new_n23850_), .A2(new_n23849_), .ZN(new_n23851_));
  NOR2_X1    g23554(.A1(new_n23851_), .A2(new_n23848_), .ZN(new_n23852_));
  NAND2_X1   g23555(.A1(new_n23724_), .A2(new_n23681_), .ZN(new_n23853_));
  NAND2_X1   g23556(.A1(new_n23853_), .A2(new_n23727_), .ZN(new_n23854_));
  INV_X1     g23557(.I(new_n23854_), .ZN(new_n23855_));
  AOI22_X1   g23558(.A1(new_n11415_), .A2(new_n11740_), .B1(\b[53] ), .B2(new_n10145_), .ZN(new_n23856_));
  OAI21_X1   g23559(.A1(new_n23856_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23857_));
  XNOR2_X1   g23560(.A1(new_n11298_), .A2(new_n23857_), .ZN(new_n23858_));
  NOR2_X1    g23561(.A1(new_n23855_), .A2(new_n23858_), .ZN(new_n23859_));
  INV_X1     g23562(.I(new_n23858_), .ZN(new_n23860_));
  NOR2_X1    g23563(.A1(new_n23854_), .A2(new_n23860_), .ZN(new_n23861_));
  NOR2_X1    g23564(.A1(new_n23859_), .A2(new_n23861_), .ZN(new_n23862_));
  NOR2_X1    g23565(.A1(new_n23862_), .A2(new_n23852_), .ZN(new_n23863_));
  INV_X1     g23566(.I(new_n23852_), .ZN(new_n23864_));
  XOR2_X1    g23567(.A1(new_n23854_), .A2(new_n23858_), .Z(new_n23865_));
  NOR2_X1    g23568(.A1(new_n23864_), .A2(new_n23865_), .ZN(new_n23866_));
  NOR2_X1    g23569(.A1(new_n23863_), .A2(new_n23866_), .ZN(new_n23867_));
  XOR2_X1    g23570(.A1(new_n23805_), .A2(new_n23867_), .Z(new_n23868_));
  NOR2_X1    g23571(.A1(new_n23868_), .A2(new_n23803_), .ZN(new_n23869_));
  INV_X1     g23572(.I(new_n23803_), .ZN(new_n23870_));
  INV_X1     g23573(.I(new_n23805_), .ZN(new_n23871_));
  NOR2_X1    g23574(.A1(new_n23871_), .A2(new_n23867_), .ZN(new_n23872_));
  INV_X1     g23575(.I(new_n23872_), .ZN(new_n23873_));
  NAND2_X1   g23576(.A1(new_n23871_), .A2(new_n23867_), .ZN(new_n23874_));
  AOI21_X1   g23577(.A1(new_n23873_), .A2(new_n23874_), .B(new_n23870_), .ZN(new_n23875_));
  NOR2_X1    g23578(.A1(new_n23875_), .A2(new_n23869_), .ZN(new_n23876_));
  NOR2_X1    g23579(.A1(new_n23799_), .A2(new_n23876_), .ZN(new_n23877_));
  NOR3_X1    g23580(.A1(new_n23798_), .A2(new_n23869_), .A3(new_n23875_), .ZN(new_n23878_));
  OAI21_X1   g23581(.A1(new_n23877_), .A2(new_n23878_), .B(new_n23796_), .ZN(new_n23879_));
  XOR2_X1    g23582(.A1(new_n23798_), .A2(new_n23876_), .Z(new_n23880_));
  OAI21_X1   g23583(.A1(new_n23796_), .A2(new_n23880_), .B(new_n23879_), .ZN(new_n23881_));
  INV_X1     g23584(.I(new_n23881_), .ZN(new_n23882_));
  NOR2_X1    g23585(.A1(new_n23882_), .A2(new_n23791_), .ZN(new_n23883_));
  INV_X1     g23586(.I(new_n23883_), .ZN(new_n23884_));
  NAND2_X1   g23587(.A1(new_n23882_), .A2(new_n23791_), .ZN(new_n23885_));
  AOI21_X1   g23588(.A1(new_n23884_), .A2(new_n23885_), .B(new_n23790_), .ZN(new_n23886_));
  INV_X1     g23589(.I(new_n23790_), .ZN(new_n23887_));
  XOR2_X1    g23590(.A1(new_n23881_), .A2(new_n23791_), .Z(new_n23888_));
  NOR2_X1    g23591(.A1(new_n23888_), .A2(new_n23887_), .ZN(new_n23889_));
  NOR2_X1    g23592(.A1(new_n23886_), .A2(new_n23889_), .ZN(new_n23890_));
  INV_X1     g23593(.I(new_n23890_), .ZN(new_n23891_));
  OAI21_X1   g23594(.A1(new_n23672_), .A2(new_n23767_), .B(new_n23769_), .ZN(new_n23892_));
  NAND2_X1   g23595(.A1(new_n23891_), .A2(new_n23892_), .ZN(new_n23893_));
  XOR2_X1    g23596(.A1(new_n23786_), .A2(new_n23893_), .Z(new_n23894_));
  XOR2_X1    g23597(.A1(new_n23894_), .A2(new_n23782_), .Z(\f[106] ));
  INV_X1     g23598(.I(new_n23782_), .ZN(new_n23896_));
  NOR2_X1    g23599(.A1(new_n23896_), .A2(new_n23890_), .ZN(new_n23897_));
  INV_X1     g23600(.I(new_n23897_), .ZN(new_n23898_));
  OAI21_X1   g23601(.A1(new_n23782_), .A2(new_n23891_), .B(new_n23892_), .ZN(new_n23899_));
  INV_X1     g23602(.I(new_n23899_), .ZN(new_n23900_));
  NAND3_X1   g23603(.A1(new_n23551_), .A2(new_n23785_), .A3(new_n23900_), .ZN(new_n23901_));
  NAND2_X1   g23604(.A1(new_n23901_), .A2(new_n23898_), .ZN(new_n23902_));
  AOI21_X1   g23605(.A1(new_n23887_), .A2(new_n23885_), .B(new_n23883_), .ZN(new_n23903_));
  OAI22_X1   g23606(.A1(new_n7619_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n8309_), .ZN(new_n23904_));
  OAI21_X1   g23607(.A1(new_n13367_), .A2(new_n7947_), .B(new_n23904_), .ZN(new_n23905_));
  AOI21_X1   g23608(.A1(new_n23905_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n23906_));
  XOR2_X1    g23609(.A1(new_n14213_), .A2(new_n23906_), .Z(new_n23907_));
  INV_X1     g23610(.I(new_n11745_), .ZN(new_n23908_));
  AOI22_X1   g23611(.A1(new_n11415_), .A2(new_n23908_), .B1(\b[54] ), .B2(new_n10145_), .ZN(new_n23909_));
  OAI21_X1   g23612(.A1(new_n23909_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n23910_));
  XOR2_X1    g23613(.A1(new_n11748_), .A2(new_n23910_), .Z(new_n23911_));
  INV_X1     g23614(.I(new_n23911_), .ZN(new_n23912_));
  INV_X1     g23615(.I(new_n23846_), .ZN(new_n23913_));
  AOI21_X1   g23616(.A1(new_n23913_), .A2(new_n23849_), .B(new_n23845_), .ZN(new_n23914_));
  INV_X1     g23617(.I(new_n23914_), .ZN(new_n23915_));
  AOI22_X1   g23618(.A1(new_n10969_), .A2(new_n10858_), .B1(new_n11394_), .B2(\b[51] ), .ZN(new_n23916_));
  OAI21_X1   g23619(.A1(new_n23916_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n23917_));
  XNOR2_X1   g23620(.A1(new_n10476_), .A2(new_n23917_), .ZN(new_n23918_));
  AOI22_X1   g23621(.A1(new_n13078_), .A2(\b[48] ), .B1(new_n23193_), .B2(new_n12218_), .ZN(new_n23919_));
  OAI21_X1   g23622(.A1(new_n23919_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n23920_));
  XOR2_X1    g23623(.A1(new_n9299_), .A2(new_n23920_), .Z(new_n23921_));
  OAI21_X1   g23624(.A1(new_n23813_), .A2(new_n23824_), .B(new_n23826_), .ZN(new_n23922_));
  OAI22_X1   g23625(.A1(new_n13880_), .A2(new_n8556_), .B1(new_n7864_), .B2(new_n13885_), .ZN(new_n23923_));
  AOI21_X1   g23626(.A1(new_n23923_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n23924_));
  XOR2_X1    g23627(.A1(new_n8217_), .A2(new_n23924_), .Z(new_n23925_));
  NOR2_X1    g23628(.A1(new_n13476_), .A2(new_n6847_), .ZN(new_n23926_));
  XOR2_X1    g23629(.A1(new_n14736_), .A2(new_n6847_), .Z(new_n23927_));
  NAND2_X1   g23630(.A1(new_n23927_), .A2(\b[44] ), .ZN(new_n23928_));
  XOR2_X1    g23631(.A1(new_n23928_), .A2(new_n23926_), .Z(new_n23929_));
  XOR2_X1    g23632(.A1(new_n23819_), .A2(new_n23929_), .Z(new_n23930_));
  NOR2_X1    g23633(.A1(new_n23820_), .A2(new_n23929_), .ZN(new_n23931_));
  NAND2_X1   g23634(.A1(new_n23820_), .A2(new_n23929_), .ZN(new_n23932_));
  INV_X1     g23635(.I(new_n23932_), .ZN(new_n23933_));
  OAI21_X1   g23636(.A1(new_n23931_), .A2(new_n23933_), .B(new_n23925_), .ZN(new_n23934_));
  OAI21_X1   g23637(.A1(new_n23925_), .A2(new_n23930_), .B(new_n23934_), .ZN(new_n23935_));
  XOR2_X1    g23638(.A1(new_n23935_), .A2(new_n23922_), .Z(new_n23936_));
  NOR2_X1    g23639(.A1(new_n23936_), .A2(new_n23921_), .ZN(new_n23937_));
  INV_X1     g23640(.I(new_n23921_), .ZN(new_n23938_));
  INV_X1     g23641(.I(new_n23922_), .ZN(new_n23939_));
  NAND2_X1   g23642(.A1(new_n23935_), .A2(new_n23939_), .ZN(new_n23940_));
  NOR2_X1    g23643(.A1(new_n23935_), .A2(new_n23939_), .ZN(new_n23941_));
  INV_X1     g23644(.I(new_n23941_), .ZN(new_n23942_));
  AOI21_X1   g23645(.A1(new_n23940_), .A2(new_n23942_), .B(new_n23938_), .ZN(new_n23943_));
  NOR2_X1    g23646(.A1(new_n23943_), .A2(new_n23937_), .ZN(new_n23944_));
  NOR2_X1    g23647(.A1(new_n23835_), .A2(new_n23810_), .ZN(new_n23945_));
  NOR2_X1    g23648(.A1(new_n23945_), .A2(new_n23833_), .ZN(new_n23946_));
  XOR2_X1    g23649(.A1(new_n23944_), .A2(new_n23946_), .Z(new_n23947_));
  NOR2_X1    g23650(.A1(new_n23947_), .A2(new_n23918_), .ZN(new_n23948_));
  INV_X1     g23651(.I(new_n23918_), .ZN(new_n23949_));
  INV_X1     g23652(.I(new_n23944_), .ZN(new_n23950_));
  NOR2_X1    g23653(.A1(new_n23950_), .A2(new_n23946_), .ZN(new_n23951_));
  INV_X1     g23654(.I(new_n23951_), .ZN(new_n23952_));
  NAND2_X1   g23655(.A1(new_n23950_), .A2(new_n23946_), .ZN(new_n23953_));
  AOI21_X1   g23656(.A1(new_n23952_), .A2(new_n23953_), .B(new_n23949_), .ZN(new_n23954_));
  NOR2_X1    g23657(.A1(new_n23954_), .A2(new_n23948_), .ZN(new_n23955_));
  XOR2_X1    g23658(.A1(new_n23955_), .A2(new_n23915_), .Z(new_n23956_));
  NAND2_X1   g23659(.A1(new_n23956_), .A2(new_n23912_), .ZN(new_n23957_));
  NOR2_X1    g23660(.A1(new_n23955_), .A2(new_n23915_), .ZN(new_n23958_));
  NAND2_X1   g23661(.A1(new_n23955_), .A2(new_n23915_), .ZN(new_n23959_));
  INV_X1     g23662(.I(new_n23959_), .ZN(new_n23960_));
  OAI21_X1   g23663(.A1(new_n23960_), .A2(new_n23958_), .B(new_n23911_), .ZN(new_n23961_));
  NAND2_X1   g23664(.A1(new_n23957_), .A2(new_n23961_), .ZN(new_n23962_));
  OAI22_X1   g23665(.A1(new_n8644_), .A2(new_n12542_), .B1(new_n12970_), .B2(new_n9388_), .ZN(new_n23963_));
  OAI21_X1   g23666(.A1(new_n12536_), .A2(new_n10154_), .B(new_n23963_), .ZN(new_n23964_));
  AOI21_X1   g23667(.A1(new_n23964_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n23965_));
  XOR2_X1    g23668(.A1(new_n12969_), .A2(new_n23965_), .Z(new_n23966_));
  NOR2_X1    g23669(.A1(new_n23852_), .A2(new_n23861_), .ZN(new_n23967_));
  NOR2_X1    g23670(.A1(new_n23967_), .A2(new_n23859_), .ZN(new_n23968_));
  XOR2_X1    g23671(.A1(new_n23968_), .A2(new_n23966_), .Z(new_n23969_));
  NOR2_X1    g23672(.A1(new_n23968_), .A2(new_n23966_), .ZN(new_n23970_));
  INV_X1     g23673(.I(new_n23970_), .ZN(new_n23971_));
  NAND2_X1   g23674(.A1(new_n23968_), .A2(new_n23966_), .ZN(new_n23972_));
  AOI21_X1   g23675(.A1(new_n23971_), .A2(new_n23972_), .B(new_n23962_), .ZN(new_n23973_));
  AOI21_X1   g23676(.A1(new_n23962_), .A2(new_n23969_), .B(new_n23973_), .ZN(new_n23974_));
  AOI21_X1   g23677(.A1(new_n23870_), .A2(new_n23874_), .B(new_n23872_), .ZN(new_n23975_));
  NOR2_X1    g23678(.A1(new_n23974_), .A2(new_n23975_), .ZN(new_n23976_));
  INV_X1     g23679(.I(new_n23976_), .ZN(new_n23977_));
  NAND2_X1   g23680(.A1(new_n23974_), .A2(new_n23975_), .ZN(new_n23978_));
  AOI21_X1   g23681(.A1(new_n23977_), .A2(new_n23978_), .B(new_n23907_), .ZN(new_n23979_));
  XOR2_X1    g23682(.A1(new_n23974_), .A2(new_n23975_), .Z(new_n23980_));
  AOI21_X1   g23683(.A1(new_n23907_), .A2(new_n23980_), .B(new_n23979_), .ZN(new_n23981_));
  OAI21_X1   g23684(.A1(new_n6644_), .A2(new_n7284_), .B(new_n16487_), .ZN(new_n23982_));
  NOR2_X1    g23685(.A1(new_n23877_), .A2(new_n23795_), .ZN(new_n23983_));
  NOR2_X1    g23686(.A1(new_n23983_), .A2(new_n23878_), .ZN(new_n23984_));
  XNOR2_X1   g23687(.A1(new_n23984_), .A2(new_n23982_), .ZN(new_n23985_));
  XOR2_X1    g23688(.A1(new_n23985_), .A2(new_n23981_), .Z(new_n23986_));
  NOR2_X1    g23689(.A1(new_n23986_), .A2(\a[44] ), .ZN(new_n23987_));
  NAND2_X1   g23690(.A1(new_n23986_), .A2(\a[44] ), .ZN(new_n23988_));
  INV_X1     g23691(.I(new_n23988_), .ZN(new_n23989_));
  NOR2_X1    g23692(.A1(new_n23989_), .A2(new_n23987_), .ZN(new_n23990_));
  XOR2_X1    g23693(.A1(new_n23990_), .A2(new_n23903_), .Z(new_n23991_));
  NAND2_X1   g23694(.A1(new_n23902_), .A2(new_n23991_), .ZN(new_n23992_));
  XOR2_X1    g23695(.A1(new_n23990_), .A2(new_n23903_), .Z(new_n23993_));
  OAI21_X1   g23696(.A1(new_n23902_), .A2(new_n23993_), .B(new_n23992_), .ZN(\f[107] ));
  INV_X1     g23697(.I(new_n23903_), .ZN(new_n23995_));
  INV_X1     g23698(.I(new_n23990_), .ZN(new_n23996_));
  NAND2_X1   g23699(.A1(new_n23996_), .A2(new_n23995_), .ZN(new_n23997_));
  OAI22_X1   g23700(.A1(new_n7619_), .A2(new_n14208_), .B1(new_n14592_), .B2(new_n8309_), .ZN(new_n23998_));
  OAI21_X1   g23701(.A1(new_n13785_), .A2(new_n7947_), .B(new_n23998_), .ZN(new_n23999_));
  AOI21_X1   g23702(.A1(new_n23999_), .A2(new_n7608_), .B(new_n7619_), .ZN(new_n24000_));
  XNOR2_X1   g23703(.A1(new_n14599_), .A2(new_n24000_), .ZN(new_n24001_));
  INV_X1     g23704(.I(new_n23907_), .ZN(new_n24002_));
  NAND2_X1   g23705(.A1(new_n23978_), .A2(new_n24002_), .ZN(new_n24003_));
  NAND2_X1   g23706(.A1(new_n24003_), .A2(new_n23977_), .ZN(new_n24004_));
  INV_X1     g23707(.I(new_n23962_), .ZN(new_n24005_));
  AOI21_X1   g23708(.A1(new_n24005_), .A2(new_n23972_), .B(new_n23970_), .ZN(new_n24006_));
  OAI22_X1   g23709(.A1(new_n8644_), .A2(new_n12970_), .B1(new_n13367_), .B2(new_n9388_), .ZN(new_n24007_));
  OAI21_X1   g23710(.A1(new_n12542_), .A2(new_n10154_), .B(new_n24007_), .ZN(new_n24008_));
  AOI21_X1   g23711(.A1(new_n24008_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n24009_));
  XNOR2_X1   g23712(.A1(new_n13371_), .A2(new_n24009_), .ZN(new_n24010_));
  OAI21_X1   g23713(.A1(new_n23911_), .A2(new_n23958_), .B(new_n23959_), .ZN(new_n24011_));
  INV_X1     g23714(.I(new_n24011_), .ZN(new_n24012_));
  AOI22_X1   g23715(.A1(new_n11415_), .A2(new_n12538_), .B1(\b[55] ), .B2(new_n10145_), .ZN(new_n24013_));
  OAI21_X1   g23716(.A1(new_n24013_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24014_));
  XOR2_X1    g23717(.A1(new_n12128_), .A2(new_n24014_), .Z(new_n24015_));
  AOI21_X1   g23718(.A1(new_n23949_), .A2(new_n23953_), .B(new_n23951_), .ZN(new_n24016_));
  AOI22_X1   g23719(.A1(new_n10969_), .A2(new_n23732_), .B1(new_n11394_), .B2(\b[52] ), .ZN(new_n24017_));
  OAI21_X1   g23720(.A1(new_n24017_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24018_));
  XOR2_X1    g23721(.A1(new_n10866_), .A2(new_n24018_), .Z(new_n24019_));
  INV_X1     g23722(.I(new_n24019_), .ZN(new_n24020_));
  AOI21_X1   g23723(.A1(new_n23938_), .A2(new_n23940_), .B(new_n23941_), .ZN(new_n24021_));
  INV_X1     g23724(.I(new_n24021_), .ZN(new_n24022_));
  INV_X1     g23725(.I(new_n23925_), .ZN(new_n24023_));
  AOI21_X1   g23726(.A1(new_n24023_), .A2(new_n23932_), .B(new_n23931_), .ZN(new_n24024_));
  OAI22_X1   g23727(.A1(new_n13880_), .A2(new_n8564_), .B1(new_n7870_), .B2(new_n13885_), .ZN(new_n24025_));
  AOI21_X1   g23728(.A1(new_n24025_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24026_));
  XOR2_X1    g23729(.A1(new_n8568_), .A2(new_n24026_), .Z(new_n24027_));
  NOR2_X1    g23730(.A1(new_n13476_), .A2(new_n7198_), .ZN(new_n24028_));
  XOR2_X1    g23731(.A1(new_n14736_), .A2(new_n7198_), .Z(new_n24029_));
  NAND2_X1   g23732(.A1(new_n24029_), .A2(\b[45] ), .ZN(new_n24030_));
  XOR2_X1    g23733(.A1(new_n24030_), .A2(new_n24028_), .Z(new_n24031_));
  NOR2_X1    g23734(.A1(new_n24031_), .A2(new_n6632_), .ZN(new_n24032_));
  INV_X1     g23735(.I(new_n24032_), .ZN(new_n24033_));
  NAND2_X1   g23736(.A1(new_n24031_), .A2(new_n6632_), .ZN(new_n24034_));
  AOI21_X1   g23737(.A1(new_n24033_), .A2(new_n24034_), .B(new_n23819_), .ZN(new_n24035_));
  XOR2_X1    g23738(.A1(new_n24031_), .A2(\a[44] ), .Z(new_n24036_));
  NOR2_X1    g23739(.A1(new_n24036_), .A2(new_n23820_), .ZN(new_n24037_));
  NOR2_X1    g23740(.A1(new_n24037_), .A2(new_n24035_), .ZN(new_n24038_));
  NOR2_X1    g23741(.A1(new_n24027_), .A2(new_n24038_), .ZN(new_n24039_));
  AND2_X2    g23742(.A1(new_n24027_), .A2(new_n24038_), .Z(new_n24040_));
  NOR2_X1    g23743(.A1(new_n24040_), .A2(new_n24039_), .ZN(new_n24041_));
  NOR2_X1    g23744(.A1(new_n24041_), .A2(new_n24024_), .ZN(new_n24042_));
  INV_X1     g23745(.I(new_n24024_), .ZN(new_n24043_));
  XNOR2_X1   g23746(.A1(new_n24027_), .A2(new_n24038_), .ZN(new_n24044_));
  NOR2_X1    g23747(.A1(new_n24044_), .A2(new_n24043_), .ZN(new_n24045_));
  NOR2_X1    g23748(.A1(new_n24042_), .A2(new_n24045_), .ZN(new_n24046_));
  AOI22_X1   g23749(.A1(new_n13078_), .A2(\b[49] ), .B1(new_n10027_), .B2(new_n12218_), .ZN(new_n24047_));
  OAI21_X1   g23750(.A1(new_n24047_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24048_));
  XOR2_X1    g23751(.A1(new_n9642_), .A2(new_n24048_), .Z(new_n24049_));
  XOR2_X1    g23752(.A1(new_n24046_), .A2(new_n24049_), .Z(new_n24050_));
  NAND2_X1   g23753(.A1(new_n24050_), .A2(new_n24022_), .ZN(new_n24051_));
  NOR2_X1    g23754(.A1(new_n24046_), .A2(new_n24049_), .ZN(new_n24052_));
  NAND2_X1   g23755(.A1(new_n24046_), .A2(new_n24049_), .ZN(new_n24053_));
  INV_X1     g23756(.I(new_n24053_), .ZN(new_n24054_));
  OAI21_X1   g23757(.A1(new_n24054_), .A2(new_n24052_), .B(new_n24021_), .ZN(new_n24055_));
  NAND2_X1   g23758(.A1(new_n24051_), .A2(new_n24055_), .ZN(new_n24056_));
  XOR2_X1    g23759(.A1(new_n24056_), .A2(new_n24020_), .Z(new_n24057_));
  NOR2_X1    g23760(.A1(new_n24057_), .A2(new_n24016_), .ZN(new_n24058_));
  INV_X1     g23761(.I(new_n24016_), .ZN(new_n24059_));
  AOI21_X1   g23762(.A1(new_n24051_), .A2(new_n24055_), .B(new_n24020_), .ZN(new_n24060_));
  NOR2_X1    g23763(.A1(new_n24056_), .A2(new_n24019_), .ZN(new_n24061_));
  NOR2_X1    g23764(.A1(new_n24061_), .A2(new_n24060_), .ZN(new_n24062_));
  NOR2_X1    g23765(.A1(new_n24062_), .A2(new_n24059_), .ZN(new_n24063_));
  NOR2_X1    g23766(.A1(new_n24058_), .A2(new_n24063_), .ZN(new_n24064_));
  XOR2_X1    g23767(.A1(new_n24064_), .A2(new_n24015_), .Z(new_n24065_));
  NOR2_X1    g23768(.A1(new_n24065_), .A2(new_n24012_), .ZN(new_n24066_));
  INV_X1     g23769(.I(new_n24015_), .ZN(new_n24067_));
  NOR2_X1    g23770(.A1(new_n24064_), .A2(new_n24067_), .ZN(new_n24068_));
  INV_X1     g23771(.I(new_n24068_), .ZN(new_n24069_));
  NAND2_X1   g23772(.A1(new_n24064_), .A2(new_n24067_), .ZN(new_n24070_));
  AOI21_X1   g23773(.A1(new_n24069_), .A2(new_n24070_), .B(new_n24011_), .ZN(new_n24071_));
  NOR2_X1    g23774(.A1(new_n24066_), .A2(new_n24071_), .ZN(new_n24072_));
  XOR2_X1    g23775(.A1(new_n24072_), .A2(new_n24010_), .Z(new_n24073_));
  NOR2_X1    g23776(.A1(new_n24073_), .A2(new_n24006_), .ZN(new_n24074_));
  INV_X1     g23777(.I(new_n24010_), .ZN(new_n24075_));
  NOR2_X1    g23778(.A1(new_n24072_), .A2(new_n24075_), .ZN(new_n24076_));
  INV_X1     g23779(.I(new_n24076_), .ZN(new_n24077_));
  NAND2_X1   g23780(.A1(new_n24072_), .A2(new_n24075_), .ZN(new_n24078_));
  NAND2_X1   g23781(.A1(new_n24077_), .A2(new_n24078_), .ZN(new_n24079_));
  AOI21_X1   g23782(.A1(new_n24006_), .A2(new_n24079_), .B(new_n24074_), .ZN(new_n24080_));
  XNOR2_X1   g23783(.A1(new_n24080_), .A2(new_n24004_), .ZN(new_n24081_));
  NOR2_X1    g23784(.A1(new_n24081_), .A2(new_n24001_), .ZN(new_n24082_));
  NOR2_X1    g23785(.A1(new_n24080_), .A2(new_n24004_), .ZN(new_n24083_));
  INV_X1     g23786(.I(new_n24083_), .ZN(new_n24084_));
  NAND2_X1   g23787(.A1(new_n24080_), .A2(new_n24004_), .ZN(new_n24085_));
  NAND2_X1   g23788(.A1(new_n24084_), .A2(new_n24085_), .ZN(new_n24086_));
  AOI21_X1   g23789(.A1(new_n24001_), .A2(new_n24086_), .B(new_n24082_), .ZN(new_n24087_));
  NOR2_X1    g23790(.A1(new_n23984_), .A2(new_n23981_), .ZN(new_n24088_));
  XOR2_X1    g23791(.A1(new_n23982_), .A2(new_n6632_), .Z(new_n24089_));
  AOI21_X1   g23792(.A1(new_n23984_), .A2(new_n23981_), .B(new_n24089_), .ZN(new_n24090_));
  NOR2_X1    g23793(.A1(new_n24090_), .A2(new_n24088_), .ZN(new_n24091_));
  XOR2_X1    g23794(.A1(new_n24087_), .A2(new_n24091_), .Z(new_n24092_));
  INV_X1     g23795(.I(new_n24092_), .ZN(new_n24093_));
  NAND2_X1   g23796(.A1(new_n23991_), .A2(new_n24093_), .ZN(new_n24094_));
  XOR2_X1    g23797(.A1(new_n24094_), .A2(new_n23997_), .Z(new_n24095_));
  XOR2_X1    g23798(.A1(new_n23902_), .A2(new_n24095_), .Z(\f[108] ));
  NOR3_X1    g23799(.A1(new_n24087_), .A2(new_n24088_), .A3(new_n24090_), .ZN(new_n24097_));
  INV_X1     g23800(.I(new_n24097_), .ZN(new_n24098_));
  NOR2_X1    g23801(.A1(new_n24093_), .A2(new_n23996_), .ZN(new_n24099_));
  AOI21_X1   g23802(.A1(new_n24093_), .A2(new_n23996_), .B(new_n23995_), .ZN(new_n24100_));
  NOR2_X1    g23803(.A1(new_n24100_), .A2(new_n24099_), .ZN(new_n24101_));
  INV_X1     g23804(.I(new_n24101_), .ZN(new_n24102_));
  AOI21_X1   g23805(.A1(new_n23901_), .A2(new_n23898_), .B(new_n24102_), .ZN(new_n24103_));
  NOR2_X1    g23806(.A1(new_n7947_), .A2(new_n8309_), .ZN(new_n24104_));
  NAND2_X1   g23807(.A1(new_n16148_), .A2(new_n7608_), .ZN(new_n24105_));
  OAI21_X1   g23808(.A1(new_n24104_), .A2(new_n24105_), .B(new_n7607_), .ZN(new_n24106_));
  XNOR2_X1   g23809(.A1(new_n14978_), .A2(new_n24106_), .ZN(new_n24107_));
  OAI21_X1   g23810(.A1(new_n24006_), .A2(new_n24076_), .B(new_n24078_), .ZN(new_n24108_));
  INV_X1     g23811(.I(new_n24108_), .ZN(new_n24109_));
  OAI22_X1   g23812(.A1(new_n8644_), .A2(new_n13367_), .B1(new_n13785_), .B2(new_n9388_), .ZN(new_n24110_));
  OAI21_X1   g23813(.A1(new_n12970_), .A2(new_n10154_), .B(new_n24110_), .ZN(new_n24111_));
  AOI21_X1   g23814(.A1(new_n24111_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n24112_));
  XOR2_X1    g23815(.A1(new_n13784_), .A2(new_n24112_), .Z(new_n24113_));
  OAI21_X1   g23816(.A1(new_n24012_), .A2(new_n24068_), .B(new_n24070_), .ZN(new_n24114_));
  INV_X1     g23817(.I(new_n12543_), .ZN(new_n24115_));
  AOI22_X1   g23818(.A1(new_n11415_), .A2(new_n24115_), .B1(\b[56] ), .B2(new_n10145_), .ZN(new_n24116_));
  OAI21_X1   g23819(.A1(new_n24116_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24117_));
  XOR2_X1    g23820(.A1(new_n12546_), .A2(new_n24117_), .Z(new_n24118_));
  NOR2_X1    g23821(.A1(new_n24060_), .A2(new_n24016_), .ZN(new_n24119_));
  NOR2_X1    g23822(.A1(new_n24119_), .A2(new_n24061_), .ZN(new_n24120_));
  AOI21_X1   g23823(.A1(new_n24022_), .A2(new_n24053_), .B(new_n24052_), .ZN(new_n24121_));
  AOI22_X1   g23824(.A1(new_n13078_), .A2(\b[50] ), .B1(new_n23440_), .B2(new_n12218_), .ZN(new_n24122_));
  OAI21_X1   g23825(.A1(new_n24122_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24123_));
  XOR2_X1    g23826(.A1(new_n10035_), .A2(new_n24123_), .Z(new_n24124_));
  NOR2_X1    g23827(.A1(new_n24040_), .A2(new_n24024_), .ZN(new_n24125_));
  NOR2_X1    g23828(.A1(new_n24125_), .A2(new_n24039_), .ZN(new_n24126_));
  OAI22_X1   g23829(.A1(new_n13880_), .A2(new_n9290_), .B1(new_n8218_), .B2(new_n13885_), .ZN(new_n24127_));
  AOI21_X1   g23830(.A1(new_n24127_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24128_));
  XOR2_X1    g23831(.A1(new_n8952_), .A2(new_n24128_), .Z(new_n24129_));
  NAND2_X1   g23832(.A1(new_n24034_), .A2(new_n23820_), .ZN(new_n24130_));
  NAND2_X1   g23833(.A1(new_n24130_), .A2(new_n24033_), .ZN(new_n24131_));
  NOR2_X1    g23834(.A1(new_n13476_), .A2(new_n7864_), .ZN(new_n24132_));
  XOR2_X1    g23835(.A1(new_n14736_), .A2(new_n7864_), .Z(new_n24133_));
  NAND2_X1   g23836(.A1(new_n24133_), .A2(\b[46] ), .ZN(new_n24134_));
  XOR2_X1    g23837(.A1(new_n24134_), .A2(new_n24132_), .Z(new_n24135_));
  INV_X1     g23838(.I(new_n24135_), .ZN(new_n24136_));
  XOR2_X1    g23839(.A1(new_n24131_), .A2(new_n24136_), .Z(new_n24137_));
  OR2_X2     g23840(.A1(new_n24129_), .A2(new_n24137_), .Z(new_n24138_));
  NOR2_X1    g23841(.A1(new_n24131_), .A2(new_n24135_), .ZN(new_n24139_));
  NAND2_X1   g23842(.A1(new_n24131_), .A2(new_n24135_), .ZN(new_n24140_));
  INV_X1     g23843(.I(new_n24140_), .ZN(new_n24141_));
  OAI21_X1   g23844(.A1(new_n24139_), .A2(new_n24141_), .B(new_n24129_), .ZN(new_n24142_));
  NAND2_X1   g23845(.A1(new_n24138_), .A2(new_n24142_), .ZN(new_n24143_));
  XNOR2_X1   g23846(.A1(new_n24126_), .A2(new_n24143_), .ZN(new_n24144_));
  NAND2_X1   g23847(.A1(new_n24126_), .A2(new_n24143_), .ZN(new_n24145_));
  NOR2_X1    g23848(.A1(new_n24126_), .A2(new_n24143_), .ZN(new_n24146_));
  INV_X1     g23849(.I(new_n24146_), .ZN(new_n24147_));
  NAND2_X1   g23850(.A1(new_n24147_), .A2(new_n24145_), .ZN(new_n24148_));
  NAND2_X1   g23851(.A1(new_n24148_), .A2(new_n24124_), .ZN(new_n24149_));
  OAI21_X1   g23852(.A1(new_n24124_), .A2(new_n24144_), .B(new_n24149_), .ZN(new_n24150_));
  AOI22_X1   g23853(.A1(new_n10969_), .A2(new_n11740_), .B1(new_n11394_), .B2(\b[53] ), .ZN(new_n24151_));
  OAI21_X1   g23854(.A1(new_n24151_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24152_));
  XNOR2_X1   g23855(.A1(new_n11298_), .A2(new_n24152_), .ZN(new_n24153_));
  NOR2_X1    g23856(.A1(new_n24150_), .A2(new_n24153_), .ZN(new_n24154_));
  INV_X1     g23857(.I(new_n24154_), .ZN(new_n24155_));
  NAND2_X1   g23858(.A1(new_n24150_), .A2(new_n24153_), .ZN(new_n24156_));
  AOI21_X1   g23859(.A1(new_n24155_), .A2(new_n24156_), .B(new_n24121_), .ZN(new_n24157_));
  INV_X1     g23860(.I(new_n24121_), .ZN(new_n24158_));
  XNOR2_X1   g23861(.A1(new_n24150_), .A2(new_n24153_), .ZN(new_n24159_));
  NOR2_X1    g23862(.A1(new_n24159_), .A2(new_n24158_), .ZN(new_n24160_));
  NOR2_X1    g23863(.A1(new_n24160_), .A2(new_n24157_), .ZN(new_n24161_));
  XNOR2_X1   g23864(.A1(new_n24161_), .A2(new_n24120_), .ZN(new_n24162_));
  NOR2_X1    g23865(.A1(new_n24162_), .A2(new_n24118_), .ZN(new_n24163_));
  INV_X1     g23866(.I(new_n24118_), .ZN(new_n24164_));
  NOR2_X1    g23867(.A1(new_n24161_), .A2(new_n24120_), .ZN(new_n24165_));
  INV_X1     g23868(.I(new_n24165_), .ZN(new_n24166_));
  NAND2_X1   g23869(.A1(new_n24161_), .A2(new_n24120_), .ZN(new_n24167_));
  AOI21_X1   g23870(.A1(new_n24166_), .A2(new_n24167_), .B(new_n24164_), .ZN(new_n24168_));
  NOR2_X1    g23871(.A1(new_n24163_), .A2(new_n24168_), .ZN(new_n24169_));
  NOR2_X1    g23872(.A1(new_n24169_), .A2(new_n24114_), .ZN(new_n24170_));
  INV_X1     g23873(.I(new_n24114_), .ZN(new_n24171_));
  INV_X1     g23874(.I(new_n24169_), .ZN(new_n24172_));
  NOR2_X1    g23875(.A1(new_n24172_), .A2(new_n24171_), .ZN(new_n24173_));
  NOR2_X1    g23876(.A1(new_n24173_), .A2(new_n24170_), .ZN(new_n24174_));
  NOR2_X1    g23877(.A1(new_n24174_), .A2(new_n24113_), .ZN(new_n24175_));
  INV_X1     g23878(.I(new_n24113_), .ZN(new_n24176_));
  XOR2_X1    g23879(.A1(new_n24169_), .A2(new_n24171_), .Z(new_n24177_));
  NOR2_X1    g23880(.A1(new_n24177_), .A2(new_n24176_), .ZN(new_n24178_));
  NOR2_X1    g23881(.A1(new_n24175_), .A2(new_n24178_), .ZN(new_n24179_));
  NOR2_X1    g23882(.A1(new_n24179_), .A2(new_n24109_), .ZN(new_n24180_));
  NOR3_X1    g23883(.A1(new_n24175_), .A2(new_n24108_), .A3(new_n24178_), .ZN(new_n24181_));
  NOR2_X1    g23884(.A1(new_n24180_), .A2(new_n24181_), .ZN(new_n24182_));
  NOR2_X1    g23885(.A1(new_n24182_), .A2(new_n24107_), .ZN(new_n24183_));
  INV_X1     g23886(.I(new_n24107_), .ZN(new_n24184_));
  XOR2_X1    g23887(.A1(new_n24179_), .A2(new_n24108_), .Z(new_n24185_));
  NOR2_X1    g23888(.A1(new_n24185_), .A2(new_n24184_), .ZN(new_n24186_));
  NOR2_X1    g23889(.A1(new_n24186_), .A2(new_n24183_), .ZN(new_n24187_));
  INV_X1     g23890(.I(new_n24187_), .ZN(new_n24188_));
  OAI21_X1   g23891(.A1(new_n24001_), .A2(new_n24083_), .B(new_n24085_), .ZN(new_n24189_));
  NAND2_X1   g23892(.A1(new_n24188_), .A2(new_n24189_), .ZN(new_n24190_));
  XOR2_X1    g23893(.A1(new_n24103_), .A2(new_n24190_), .Z(new_n24191_));
  XOR2_X1    g23894(.A1(new_n24191_), .A2(new_n24098_), .Z(\f[109] ));
  INV_X1     g23895(.I(new_n23785_), .ZN(new_n24193_));
  NOR3_X1    g23896(.A1(new_n23661_), .A2(new_n24193_), .A3(new_n23899_), .ZN(new_n24194_));
  OAI21_X1   g23897(.A1(new_n24194_), .A2(new_n23897_), .B(new_n24101_), .ZN(new_n24195_));
  NOR2_X1    g23898(.A1(new_n24098_), .A2(new_n24187_), .ZN(new_n24196_));
  INV_X1     g23899(.I(new_n24196_), .ZN(new_n24197_));
  OAI21_X1   g23900(.A1(new_n24097_), .A2(new_n24188_), .B(new_n24189_), .ZN(new_n24198_));
  OAI21_X1   g23901(.A1(new_n24195_), .A2(new_n24198_), .B(new_n24197_), .ZN(new_n24199_));
  OAI21_X1   g23902(.A1(new_n7619_), .A2(new_n7947_), .B(new_n16487_), .ZN(new_n24200_));
  OAI22_X1   g23903(.A1(new_n8644_), .A2(new_n13785_), .B1(new_n14208_), .B2(new_n9388_), .ZN(new_n24201_));
  OAI21_X1   g23904(.A1(new_n13367_), .A2(new_n10154_), .B(new_n24201_), .ZN(new_n24202_));
  AOI21_X1   g23905(.A1(new_n24202_), .A2(new_n8624_), .B(new_n8644_), .ZN(new_n24203_));
  XOR2_X1    g23906(.A1(new_n14213_), .A2(new_n24203_), .Z(new_n24204_));
  AOI22_X1   g23907(.A1(new_n10969_), .A2(new_n23908_), .B1(new_n11394_), .B2(\b[54] ), .ZN(new_n24205_));
  OAI21_X1   g23908(.A1(new_n24205_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24206_));
  XOR2_X1    g23909(.A1(new_n11748_), .A2(new_n24206_), .Z(new_n24207_));
  INV_X1     g23910(.I(new_n24124_), .ZN(new_n24208_));
  AOI21_X1   g23911(.A1(new_n24208_), .A2(new_n24145_), .B(new_n24146_), .ZN(new_n24209_));
  AOI22_X1   g23912(.A1(new_n13078_), .A2(\b[51] ), .B1(new_n10858_), .B2(new_n12218_), .ZN(new_n24210_));
  OAI21_X1   g23913(.A1(new_n24210_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24211_));
  XNOR2_X1   g23914(.A1(new_n10476_), .A2(new_n24211_), .ZN(new_n24212_));
  OAI21_X1   g23915(.A1(new_n24129_), .A2(new_n24139_), .B(new_n24140_), .ZN(new_n24213_));
  NOR2_X1    g23916(.A1(new_n13476_), .A2(new_n7870_), .ZN(new_n24214_));
  XOR2_X1    g23917(.A1(new_n14736_), .A2(new_n7870_), .Z(new_n24215_));
  NAND2_X1   g23918(.A1(new_n24215_), .A2(\b[47] ), .ZN(new_n24216_));
  XOR2_X1    g23919(.A1(new_n24216_), .A2(new_n24214_), .Z(new_n24217_));
  NOR2_X1    g23920(.A1(new_n24136_), .A2(new_n24217_), .ZN(new_n24218_));
  INV_X1     g23921(.I(new_n24217_), .ZN(new_n24219_));
  NOR2_X1    g23922(.A1(new_n24219_), .A2(new_n24135_), .ZN(new_n24220_));
  OAI21_X1   g23923(.A1(new_n24218_), .A2(new_n24220_), .B(new_n24213_), .ZN(new_n24221_));
  XOR2_X1    g23924(.A1(new_n24135_), .A2(new_n24217_), .Z(new_n24222_));
  OR2_X2     g23925(.A1(new_n24213_), .A2(new_n24222_), .Z(new_n24223_));
  NAND2_X1   g23926(.A1(new_n24223_), .A2(new_n24221_), .ZN(new_n24224_));
  OAI22_X1   g23927(.A1(new_n13880_), .A2(new_n9296_), .B1(new_n8563_), .B2(new_n13885_), .ZN(new_n24225_));
  AOI21_X1   g23928(.A1(new_n24225_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24226_));
  XNOR2_X1   g23929(.A1(new_n9299_), .A2(new_n24226_), .ZN(new_n24227_));
  XOR2_X1    g23930(.A1(new_n24224_), .A2(new_n24227_), .Z(new_n24228_));
  NOR2_X1    g23931(.A1(new_n24228_), .A2(new_n24212_), .ZN(new_n24229_));
  INV_X1     g23932(.I(new_n24212_), .ZN(new_n24230_));
  INV_X1     g23933(.I(new_n24224_), .ZN(new_n24231_));
  NOR2_X1    g23934(.A1(new_n24231_), .A2(new_n24227_), .ZN(new_n24232_));
  INV_X1     g23935(.I(new_n24232_), .ZN(new_n24233_));
  NAND2_X1   g23936(.A1(new_n24231_), .A2(new_n24227_), .ZN(new_n24234_));
  AOI21_X1   g23937(.A1(new_n24233_), .A2(new_n24234_), .B(new_n24230_), .ZN(new_n24235_));
  NOR2_X1    g23938(.A1(new_n24235_), .A2(new_n24229_), .ZN(new_n24236_));
  XOR2_X1    g23939(.A1(new_n24236_), .A2(new_n24209_), .Z(new_n24237_));
  NOR2_X1    g23940(.A1(new_n24237_), .A2(new_n24207_), .ZN(new_n24238_));
  INV_X1     g23941(.I(new_n24209_), .ZN(new_n24239_));
  NOR2_X1    g23942(.A1(new_n24236_), .A2(new_n24239_), .ZN(new_n24240_));
  INV_X1     g23943(.I(new_n24240_), .ZN(new_n24241_));
  NAND2_X1   g23944(.A1(new_n24236_), .A2(new_n24239_), .ZN(new_n24242_));
  NAND2_X1   g23945(.A1(new_n24241_), .A2(new_n24242_), .ZN(new_n24243_));
  AOI21_X1   g23946(.A1(new_n24207_), .A2(new_n24243_), .B(new_n24238_), .ZN(new_n24244_));
  AOI22_X1   g23947(.A1(new_n11415_), .A2(new_n13363_), .B1(\b[57] ), .B2(new_n10145_), .ZN(new_n24245_));
  OAI21_X1   g23948(.A1(new_n24245_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24246_));
  XNOR2_X1   g23949(.A1(new_n12969_), .A2(new_n24246_), .ZN(new_n24247_));
  AOI21_X1   g23950(.A1(new_n24158_), .A2(new_n24156_), .B(new_n24154_), .ZN(new_n24248_));
  XNOR2_X1   g23951(.A1(new_n24248_), .A2(new_n24247_), .ZN(new_n24249_));
  NOR2_X1    g23952(.A1(new_n24249_), .A2(new_n24244_), .ZN(new_n24250_));
  NOR2_X1    g23953(.A1(new_n24248_), .A2(new_n24247_), .ZN(new_n24251_));
  INV_X1     g23954(.I(new_n24251_), .ZN(new_n24252_));
  NAND2_X1   g23955(.A1(new_n24248_), .A2(new_n24247_), .ZN(new_n24253_));
  NAND2_X1   g23956(.A1(new_n24252_), .A2(new_n24253_), .ZN(new_n24254_));
  AOI21_X1   g23957(.A1(new_n24244_), .A2(new_n24254_), .B(new_n24250_), .ZN(new_n24255_));
  AOI21_X1   g23958(.A1(new_n24164_), .A2(new_n24167_), .B(new_n24165_), .ZN(new_n24256_));
  NOR2_X1    g23959(.A1(new_n24255_), .A2(new_n24256_), .ZN(new_n24257_));
  INV_X1     g23960(.I(new_n24257_), .ZN(new_n24258_));
  NAND2_X1   g23961(.A1(new_n24255_), .A2(new_n24256_), .ZN(new_n24259_));
  AOI21_X1   g23962(.A1(new_n24258_), .A2(new_n24259_), .B(new_n24204_), .ZN(new_n24260_));
  INV_X1     g23963(.I(new_n24204_), .ZN(new_n24261_));
  XNOR2_X1   g23964(.A1(new_n24255_), .A2(new_n24256_), .ZN(new_n24262_));
  NOR2_X1    g23965(.A1(new_n24262_), .A2(new_n24261_), .ZN(new_n24263_));
  NOR2_X1    g23966(.A1(new_n24263_), .A2(new_n24260_), .ZN(new_n24264_));
  INV_X1     g23967(.I(new_n24170_), .ZN(new_n24265_));
  AOI21_X1   g23968(.A1(new_n24176_), .A2(new_n24265_), .B(new_n24173_), .ZN(new_n24266_));
  XNOR2_X1   g23969(.A1(new_n24266_), .A2(new_n24264_), .ZN(new_n24267_));
  XOR2_X1    g23970(.A1(new_n24267_), .A2(new_n24200_), .Z(new_n24268_));
  OR2_X2     g23971(.A1(new_n24268_), .A2(\a[47] ), .Z(new_n24269_));
  NAND2_X1   g23972(.A1(new_n24268_), .A2(\a[47] ), .ZN(new_n24270_));
  NAND2_X1   g23973(.A1(new_n24269_), .A2(new_n24270_), .ZN(new_n24271_));
  INV_X1     g23974(.I(new_n24181_), .ZN(new_n24272_));
  AOI21_X1   g23975(.A1(new_n24272_), .A2(new_n24184_), .B(new_n24180_), .ZN(new_n24273_));
  INV_X1     g23976(.I(new_n24273_), .ZN(new_n24274_));
  XOR2_X1    g23977(.A1(new_n24271_), .A2(new_n24274_), .Z(new_n24275_));
  NAND2_X1   g23978(.A1(new_n24199_), .A2(new_n24275_), .ZN(new_n24276_));
  INV_X1     g23979(.I(new_n24198_), .ZN(new_n24277_));
  AOI21_X1   g23980(.A1(new_n24103_), .A2(new_n24277_), .B(new_n24196_), .ZN(new_n24278_));
  NAND2_X1   g23981(.A1(new_n24271_), .A2(new_n24274_), .ZN(new_n24279_));
  INV_X1     g23982(.I(new_n24271_), .ZN(new_n24280_));
  NAND2_X1   g23983(.A1(new_n24280_), .A2(new_n24273_), .ZN(new_n24281_));
  NAND2_X1   g23984(.A1(new_n24281_), .A2(new_n24279_), .ZN(new_n24282_));
  NAND2_X1   g23985(.A1(new_n24278_), .A2(new_n24282_), .ZN(new_n24283_));
  NAND2_X1   g23986(.A1(new_n24276_), .A2(new_n24283_), .ZN(\f[110] ));
  AOI22_X1   g23987(.A1(new_n8631_), .A2(\b[62] ), .B1(\b[63] ), .B2(new_n9382_), .ZN(new_n24285_));
  AOI21_X1   g23988(.A1(\b[61] ), .A2(new_n9731_), .B(new_n24285_), .ZN(new_n24286_));
  OAI21_X1   g23989(.A1(new_n24286_), .A2(\a[50] ), .B(new_n8631_), .ZN(new_n24287_));
  XOR2_X1    g23990(.A1(new_n14599_), .A2(new_n24287_), .Z(new_n24288_));
  INV_X1     g23991(.I(new_n24288_), .ZN(new_n24289_));
  NAND2_X1   g23992(.A1(new_n24259_), .A2(new_n24261_), .ZN(new_n24290_));
  NAND2_X1   g23993(.A1(new_n24290_), .A2(new_n24258_), .ZN(new_n24291_));
  AOI21_X1   g23994(.A1(new_n24244_), .A2(new_n24253_), .B(new_n24251_), .ZN(new_n24292_));
  INV_X1     g23995(.I(new_n24292_), .ZN(new_n24293_));
  INV_X1     g23996(.I(new_n13368_), .ZN(new_n24294_));
  AOI22_X1   g23997(.A1(new_n11415_), .A2(new_n24294_), .B1(\b[58] ), .B2(new_n10145_), .ZN(new_n24295_));
  OAI21_X1   g23998(.A1(new_n24295_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24296_));
  XOR2_X1    g23999(.A1(new_n13371_), .A2(new_n24296_), .Z(new_n24297_));
  OAI21_X1   g24000(.A1(new_n24207_), .A2(new_n24240_), .B(new_n24242_), .ZN(new_n24298_));
  AOI22_X1   g24001(.A1(new_n10969_), .A2(new_n12538_), .B1(new_n11394_), .B2(\b[55] ), .ZN(new_n24299_));
  OAI21_X1   g24002(.A1(new_n24299_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24300_));
  XOR2_X1    g24003(.A1(new_n12128_), .A2(new_n24300_), .Z(new_n24301_));
  INV_X1     g24004(.I(new_n24301_), .ZN(new_n24302_));
  AOI21_X1   g24005(.A1(new_n24230_), .A2(new_n24234_), .B(new_n24232_), .ZN(new_n24303_));
  INV_X1     g24006(.I(new_n24218_), .ZN(new_n24304_));
  AOI21_X1   g24007(.A1(new_n24213_), .A2(new_n24304_), .B(new_n24220_), .ZN(new_n24305_));
  OAI22_X1   g24008(.A1(new_n13880_), .A2(new_n10026_), .B1(new_n8948_), .B2(new_n13885_), .ZN(new_n24306_));
  AOI21_X1   g24009(.A1(new_n24306_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24307_));
  XNOR2_X1   g24010(.A1(new_n9642_), .A2(new_n24307_), .ZN(new_n24308_));
  INV_X1     g24011(.I(new_n24308_), .ZN(new_n24309_));
  NOR2_X1    g24012(.A1(new_n13476_), .A2(new_n8218_), .ZN(new_n24310_));
  XOR2_X1    g24013(.A1(new_n14736_), .A2(new_n8218_), .Z(new_n24311_));
  NAND2_X1   g24014(.A1(new_n24311_), .A2(\b[48] ), .ZN(new_n24312_));
  XOR2_X1    g24015(.A1(new_n24312_), .A2(new_n24310_), .Z(new_n24313_));
  XOR2_X1    g24016(.A1(new_n24313_), .A2(\a[47] ), .Z(new_n24314_));
  NOR2_X1    g24017(.A1(new_n24314_), .A2(new_n24217_), .ZN(new_n24315_));
  NOR2_X1    g24018(.A1(new_n24313_), .A2(new_n7608_), .ZN(new_n24316_));
  INV_X1     g24019(.I(new_n24316_), .ZN(new_n24317_));
  NAND2_X1   g24020(.A1(new_n24313_), .A2(new_n7608_), .ZN(new_n24318_));
  AOI21_X1   g24021(.A1(new_n24317_), .A2(new_n24318_), .B(new_n24219_), .ZN(new_n24319_));
  NOR2_X1    g24022(.A1(new_n24315_), .A2(new_n24319_), .ZN(new_n24320_));
  NOR2_X1    g24023(.A1(new_n24309_), .A2(new_n24320_), .ZN(new_n24321_));
  INV_X1     g24024(.I(new_n24321_), .ZN(new_n24322_));
  NAND2_X1   g24025(.A1(new_n24309_), .A2(new_n24320_), .ZN(new_n24323_));
  AOI21_X1   g24026(.A1(new_n24322_), .A2(new_n24323_), .B(new_n24305_), .ZN(new_n24324_));
  XOR2_X1    g24027(.A1(new_n24308_), .A2(new_n24320_), .Z(new_n24325_));
  INV_X1     g24028(.I(new_n24325_), .ZN(new_n24326_));
  AOI21_X1   g24029(.A1(new_n24305_), .A2(new_n24326_), .B(new_n24324_), .ZN(new_n24327_));
  AOI22_X1   g24030(.A1(new_n13078_), .A2(\b[52] ), .B1(new_n23732_), .B2(new_n12218_), .ZN(new_n24328_));
  OAI21_X1   g24031(.A1(new_n24328_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24329_));
  XOR2_X1    g24032(.A1(new_n10866_), .A2(new_n24329_), .Z(new_n24330_));
  XNOR2_X1   g24033(.A1(new_n24327_), .A2(new_n24330_), .ZN(new_n24331_));
  NOR2_X1    g24034(.A1(new_n24331_), .A2(new_n24303_), .ZN(new_n24332_));
  INV_X1     g24035(.I(new_n24303_), .ZN(new_n24333_));
  NOR2_X1    g24036(.A1(new_n24327_), .A2(new_n24330_), .ZN(new_n24334_));
  INV_X1     g24037(.I(new_n24334_), .ZN(new_n24335_));
  NAND2_X1   g24038(.A1(new_n24327_), .A2(new_n24330_), .ZN(new_n24336_));
  AOI21_X1   g24039(.A1(new_n24335_), .A2(new_n24336_), .B(new_n24333_), .ZN(new_n24337_));
  NOR2_X1    g24040(.A1(new_n24332_), .A2(new_n24337_), .ZN(new_n24338_));
  XOR2_X1    g24041(.A1(new_n24338_), .A2(new_n24302_), .Z(new_n24339_));
  NAND2_X1   g24042(.A1(new_n24339_), .A2(new_n24298_), .ZN(new_n24340_));
  INV_X1     g24043(.I(new_n24298_), .ZN(new_n24341_));
  NOR2_X1    g24044(.A1(new_n24338_), .A2(new_n24302_), .ZN(new_n24342_));
  NAND2_X1   g24045(.A1(new_n24338_), .A2(new_n24302_), .ZN(new_n24343_));
  INV_X1     g24046(.I(new_n24343_), .ZN(new_n24344_));
  OAI21_X1   g24047(.A1(new_n24344_), .A2(new_n24342_), .B(new_n24341_), .ZN(new_n24345_));
  NAND2_X1   g24048(.A1(new_n24340_), .A2(new_n24345_), .ZN(new_n24346_));
  XOR2_X1    g24049(.A1(new_n24346_), .A2(new_n24297_), .Z(new_n24347_));
  NAND2_X1   g24050(.A1(new_n24347_), .A2(new_n24293_), .ZN(new_n24348_));
  AND2_X2    g24051(.A1(new_n24346_), .A2(new_n24297_), .Z(new_n24349_));
  NOR2_X1    g24052(.A1(new_n24346_), .A2(new_n24297_), .ZN(new_n24350_));
  OAI21_X1   g24053(.A1(new_n24349_), .A2(new_n24350_), .B(new_n24292_), .ZN(new_n24351_));
  NAND2_X1   g24054(.A1(new_n24348_), .A2(new_n24351_), .ZN(new_n24352_));
  XNOR2_X1   g24055(.A1(new_n24352_), .A2(new_n24291_), .ZN(new_n24353_));
  INV_X1     g24056(.I(new_n24352_), .ZN(new_n24354_));
  NOR2_X1    g24057(.A1(new_n24354_), .A2(new_n24291_), .ZN(new_n24355_));
  INV_X1     g24058(.I(new_n24355_), .ZN(new_n24356_));
  NAND2_X1   g24059(.A1(new_n24354_), .A2(new_n24291_), .ZN(new_n24357_));
  AOI21_X1   g24060(.A1(new_n24356_), .A2(new_n24357_), .B(new_n24289_), .ZN(new_n24358_));
  AOI21_X1   g24061(.A1(new_n24289_), .A2(new_n24353_), .B(new_n24358_), .ZN(new_n24359_));
  INV_X1     g24062(.I(new_n24264_), .ZN(new_n24360_));
  INV_X1     g24063(.I(new_n24266_), .ZN(new_n24361_));
  XOR2_X1    g24064(.A1(new_n24200_), .A2(\a[47] ), .Z(new_n24362_));
  OAI21_X1   g24065(.A1(new_n24361_), .A2(new_n24360_), .B(new_n24362_), .ZN(new_n24363_));
  OAI21_X1   g24066(.A1(new_n24264_), .A2(new_n24266_), .B(new_n24363_), .ZN(new_n24364_));
  XOR2_X1    g24067(.A1(new_n24359_), .A2(new_n24364_), .Z(new_n24365_));
  NAND2_X1   g24068(.A1(new_n24275_), .A2(new_n24365_), .ZN(new_n24366_));
  XNOR2_X1   g24069(.A1(new_n24366_), .A2(new_n24279_), .ZN(new_n24367_));
  XOR2_X1    g24070(.A1(new_n24278_), .A2(new_n24367_), .Z(\f[111] ));
  NOR2_X1    g24071(.A1(new_n24359_), .A2(new_n24364_), .ZN(new_n24369_));
  NOR2_X1    g24072(.A1(new_n24365_), .A2(new_n24274_), .ZN(new_n24370_));
  NAND2_X1   g24073(.A1(new_n24365_), .A2(new_n24274_), .ZN(new_n24371_));
  AOI21_X1   g24074(.A1(new_n24280_), .A2(new_n24371_), .B(new_n24370_), .ZN(new_n24372_));
  NAND2_X1   g24075(.A1(new_n24199_), .A2(new_n24372_), .ZN(new_n24373_));
  NOR2_X1    g24076(.A1(new_n10154_), .A2(new_n9388_), .ZN(new_n24374_));
  NAND2_X1   g24077(.A1(new_n16148_), .A2(new_n8624_), .ZN(new_n24375_));
  OAI21_X1   g24078(.A1(new_n24374_), .A2(new_n24375_), .B(new_n8631_), .ZN(new_n24376_));
  XNOR2_X1   g24079(.A1(new_n14978_), .A2(new_n24376_), .ZN(new_n24377_));
  NOR2_X1    g24080(.A1(new_n24349_), .A2(new_n24292_), .ZN(new_n24378_));
  AOI22_X1   g24081(.A1(new_n11415_), .A2(new_n14202_), .B1(\b[59] ), .B2(new_n10145_), .ZN(new_n24379_));
  OAI21_X1   g24082(.A1(new_n24379_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24380_));
  XNOR2_X1   g24083(.A1(new_n13784_), .A2(new_n24380_), .ZN(new_n24381_));
  OAI21_X1   g24084(.A1(new_n24341_), .A2(new_n24342_), .B(new_n24343_), .ZN(new_n24382_));
  AOI22_X1   g24085(.A1(new_n10969_), .A2(new_n24115_), .B1(new_n11394_), .B2(\b[56] ), .ZN(new_n24383_));
  OAI21_X1   g24086(.A1(new_n24383_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24384_));
  XOR2_X1    g24087(.A1(new_n12546_), .A2(new_n24384_), .Z(new_n24385_));
  NAND2_X1   g24088(.A1(new_n24336_), .A2(new_n24333_), .ZN(new_n24386_));
  NAND2_X1   g24089(.A1(new_n24386_), .A2(new_n24335_), .ZN(new_n24387_));
  AOI22_X1   g24090(.A1(new_n13078_), .A2(\b[53] ), .B1(new_n11740_), .B2(new_n12218_), .ZN(new_n24388_));
  OAI21_X1   g24091(.A1(new_n24388_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24389_));
  XNOR2_X1   g24092(.A1(new_n11298_), .A2(new_n24389_), .ZN(new_n24390_));
  OAI21_X1   g24093(.A1(new_n24305_), .A2(new_n24321_), .B(new_n24323_), .ZN(new_n24391_));
  OAI22_X1   g24094(.A1(new_n13880_), .A2(new_n10032_), .B1(new_n9295_), .B2(new_n13885_), .ZN(new_n24392_));
  AOI21_X1   g24095(.A1(new_n24392_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24393_));
  XNOR2_X1   g24096(.A1(new_n10035_), .A2(new_n24393_), .ZN(new_n24394_));
  NAND2_X1   g24097(.A1(new_n24318_), .A2(new_n24219_), .ZN(new_n24395_));
  NAND2_X1   g24098(.A1(new_n24395_), .A2(new_n24317_), .ZN(new_n24396_));
  NOR2_X1    g24099(.A1(new_n13476_), .A2(new_n8563_), .ZN(new_n24397_));
  XOR2_X1    g24100(.A1(new_n14736_), .A2(new_n8563_), .Z(new_n24398_));
  NAND2_X1   g24101(.A1(new_n24398_), .A2(\b[49] ), .ZN(new_n24399_));
  XOR2_X1    g24102(.A1(new_n24399_), .A2(new_n24397_), .Z(new_n24400_));
  INV_X1     g24103(.I(new_n24400_), .ZN(new_n24401_));
  XOR2_X1    g24104(.A1(new_n24396_), .A2(new_n24401_), .Z(new_n24402_));
  NOR2_X1    g24105(.A1(new_n24394_), .A2(new_n24402_), .ZN(new_n24403_));
  NOR2_X1    g24106(.A1(new_n24396_), .A2(new_n24400_), .ZN(new_n24404_));
  INV_X1     g24107(.I(new_n24404_), .ZN(new_n24405_));
  NAND2_X1   g24108(.A1(new_n24396_), .A2(new_n24400_), .ZN(new_n24406_));
  NAND2_X1   g24109(.A1(new_n24405_), .A2(new_n24406_), .ZN(new_n24407_));
  AOI21_X1   g24110(.A1(new_n24394_), .A2(new_n24407_), .B(new_n24403_), .ZN(new_n24408_));
  XNOR2_X1   g24111(.A1(new_n24408_), .A2(new_n24391_), .ZN(new_n24409_));
  NOR2_X1    g24112(.A1(new_n24409_), .A2(new_n24390_), .ZN(new_n24410_));
  NOR2_X1    g24113(.A1(new_n24408_), .A2(new_n24391_), .ZN(new_n24411_));
  INV_X1     g24114(.I(new_n24411_), .ZN(new_n24412_));
  NAND2_X1   g24115(.A1(new_n24408_), .A2(new_n24391_), .ZN(new_n24413_));
  NAND2_X1   g24116(.A1(new_n24412_), .A2(new_n24413_), .ZN(new_n24414_));
  AOI21_X1   g24117(.A1(new_n24390_), .A2(new_n24414_), .B(new_n24410_), .ZN(new_n24415_));
  XNOR2_X1   g24118(.A1(new_n24415_), .A2(new_n24387_), .ZN(new_n24416_));
  NOR2_X1    g24119(.A1(new_n24416_), .A2(new_n24385_), .ZN(new_n24417_));
  NOR2_X1    g24120(.A1(new_n24415_), .A2(new_n24387_), .ZN(new_n24418_));
  INV_X1     g24121(.I(new_n24418_), .ZN(new_n24419_));
  NAND2_X1   g24122(.A1(new_n24415_), .A2(new_n24387_), .ZN(new_n24420_));
  NAND2_X1   g24123(.A1(new_n24419_), .A2(new_n24420_), .ZN(new_n24421_));
  AOI21_X1   g24124(.A1(new_n24385_), .A2(new_n24421_), .B(new_n24417_), .ZN(new_n24422_));
  XNOR2_X1   g24125(.A1(new_n24422_), .A2(new_n24382_), .ZN(new_n24423_));
  NOR2_X1    g24126(.A1(new_n24423_), .A2(new_n24381_), .ZN(new_n24424_));
  INV_X1     g24127(.I(new_n24381_), .ZN(new_n24425_));
  NOR2_X1    g24128(.A1(new_n24422_), .A2(new_n24382_), .ZN(new_n24426_));
  INV_X1     g24129(.I(new_n24426_), .ZN(new_n24427_));
  NAND2_X1   g24130(.A1(new_n24422_), .A2(new_n24382_), .ZN(new_n24428_));
  AOI21_X1   g24131(.A1(new_n24427_), .A2(new_n24428_), .B(new_n24425_), .ZN(new_n24429_));
  NOR2_X1    g24132(.A1(new_n24424_), .A2(new_n24429_), .ZN(new_n24430_));
  NOR3_X1    g24133(.A1(new_n24430_), .A2(new_n24350_), .A3(new_n24378_), .ZN(new_n24431_));
  NOR2_X1    g24134(.A1(new_n24378_), .A2(new_n24350_), .ZN(new_n24432_));
  INV_X1     g24135(.I(new_n24430_), .ZN(new_n24433_));
  NOR2_X1    g24136(.A1(new_n24433_), .A2(new_n24432_), .ZN(new_n24434_));
  NOR2_X1    g24137(.A1(new_n24434_), .A2(new_n24431_), .ZN(new_n24435_));
  NOR2_X1    g24138(.A1(new_n24435_), .A2(new_n24377_), .ZN(new_n24436_));
  INV_X1     g24139(.I(new_n24377_), .ZN(new_n24437_));
  XOR2_X1    g24140(.A1(new_n24430_), .A2(new_n24432_), .Z(new_n24438_));
  NOR2_X1    g24141(.A1(new_n24438_), .A2(new_n24437_), .ZN(new_n24439_));
  NOR2_X1    g24142(.A1(new_n24436_), .A2(new_n24439_), .ZN(new_n24440_));
  INV_X1     g24143(.I(new_n24440_), .ZN(new_n24441_));
  OAI21_X1   g24144(.A1(new_n24288_), .A2(new_n24355_), .B(new_n24357_), .ZN(new_n24442_));
  NAND2_X1   g24145(.A1(new_n24441_), .A2(new_n24442_), .ZN(new_n24443_));
  XOR2_X1    g24146(.A1(new_n24373_), .A2(new_n24443_), .Z(new_n24444_));
  XOR2_X1    g24147(.A1(new_n24444_), .A2(new_n24369_), .Z(\f[112] ));
  INV_X1     g24148(.I(new_n24369_), .ZN(new_n24446_));
  NOR2_X1    g24149(.A1(new_n24446_), .A2(new_n24440_), .ZN(new_n24447_));
  INV_X1     g24150(.I(new_n24447_), .ZN(new_n24448_));
  OAI21_X1   g24151(.A1(new_n24441_), .A2(new_n24369_), .B(new_n24442_), .ZN(new_n24449_));
  INV_X1     g24152(.I(new_n24449_), .ZN(new_n24450_));
  NAND3_X1   g24153(.A1(new_n24199_), .A2(new_n24372_), .A3(new_n24450_), .ZN(new_n24451_));
  NAND2_X1   g24154(.A1(new_n24451_), .A2(new_n24448_), .ZN(new_n24452_));
  OAI21_X1   g24155(.A1(new_n8644_), .A2(new_n10154_), .B(new_n16487_), .ZN(new_n24453_));
  AOI22_X1   g24156(.A1(new_n11415_), .A2(new_n14590_), .B1(\b[60] ), .B2(new_n10145_), .ZN(new_n24454_));
  OAI21_X1   g24157(.A1(new_n24454_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24455_));
  XNOR2_X1   g24158(.A1(new_n14213_), .A2(new_n24455_), .ZN(new_n24456_));
  AOI22_X1   g24159(.A1(new_n13078_), .A2(\b[54] ), .B1(new_n23908_), .B2(new_n12218_), .ZN(new_n24457_));
  OAI21_X1   g24160(.A1(new_n24457_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24458_));
  XOR2_X1    g24161(.A1(new_n11748_), .A2(new_n24458_), .Z(new_n24459_));
  INV_X1     g24162(.I(new_n24459_), .ZN(new_n24460_));
  OAI22_X1   g24163(.A1(new_n13880_), .A2(new_n10857_), .B1(new_n10025_), .B2(new_n13885_), .ZN(new_n24461_));
  AOI21_X1   g24164(.A1(new_n24461_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24462_));
  XOR2_X1    g24165(.A1(new_n10476_), .A2(new_n24462_), .Z(new_n24463_));
  INV_X1     g24166(.I(new_n24463_), .ZN(new_n24464_));
  NOR2_X1    g24167(.A1(new_n13476_), .A2(new_n8948_), .ZN(new_n24465_));
  XOR2_X1    g24168(.A1(new_n14736_), .A2(new_n8948_), .Z(new_n24466_));
  NAND2_X1   g24169(.A1(new_n24466_), .A2(\b[50] ), .ZN(new_n24467_));
  XOR2_X1    g24170(.A1(new_n24467_), .A2(new_n24465_), .Z(new_n24468_));
  NOR2_X1    g24171(.A1(new_n24401_), .A2(new_n24468_), .ZN(new_n24469_));
  INV_X1     g24172(.I(new_n24468_), .ZN(new_n24470_));
  NOR2_X1    g24173(.A1(new_n24470_), .A2(new_n24400_), .ZN(new_n24471_));
  OAI21_X1   g24174(.A1(new_n24469_), .A2(new_n24471_), .B(new_n24464_), .ZN(new_n24472_));
  XNOR2_X1   g24175(.A1(new_n24400_), .A2(new_n24468_), .ZN(new_n24473_));
  NAND2_X1   g24176(.A1(new_n24463_), .A2(new_n24473_), .ZN(new_n24474_));
  NAND2_X1   g24177(.A1(new_n24472_), .A2(new_n24474_), .ZN(new_n24475_));
  OR2_X2     g24178(.A1(new_n24394_), .A2(new_n24404_), .Z(new_n24476_));
  NAND2_X1   g24179(.A1(new_n24476_), .A2(new_n24406_), .ZN(new_n24477_));
  XNOR2_X1   g24180(.A1(new_n24477_), .A2(new_n24475_), .ZN(new_n24478_));
  INV_X1     g24181(.I(new_n24478_), .ZN(new_n24479_));
  AOI22_X1   g24182(.A1(new_n24406_), .A2(new_n24476_), .B1(new_n24472_), .B2(new_n24474_), .ZN(new_n24480_));
  NOR2_X1    g24183(.A1(new_n24477_), .A2(new_n24475_), .ZN(new_n24481_));
  NOR2_X1    g24184(.A1(new_n24481_), .A2(new_n24480_), .ZN(new_n24482_));
  NOR2_X1    g24185(.A1(new_n24460_), .A2(new_n24482_), .ZN(new_n24483_));
  AOI21_X1   g24186(.A1(new_n24479_), .A2(new_n24460_), .B(new_n24483_), .ZN(new_n24484_));
  AOI22_X1   g24187(.A1(new_n10969_), .A2(new_n13363_), .B1(new_n11394_), .B2(\b[57] ), .ZN(new_n24485_));
  OAI21_X1   g24188(.A1(new_n24485_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24486_));
  XNOR2_X1   g24189(.A1(new_n12969_), .A2(new_n24486_), .ZN(new_n24487_));
  OAI21_X1   g24190(.A1(new_n24390_), .A2(new_n24411_), .B(new_n24413_), .ZN(new_n24488_));
  XOR2_X1    g24191(.A1(new_n24487_), .A2(new_n24488_), .Z(new_n24489_));
  NOR2_X1    g24192(.A1(new_n24489_), .A2(new_n24484_), .ZN(new_n24490_));
  INV_X1     g24193(.I(new_n24484_), .ZN(new_n24491_));
  INV_X1     g24194(.I(new_n24488_), .ZN(new_n24492_));
  NOR2_X1    g24195(.A1(new_n24487_), .A2(new_n24492_), .ZN(new_n24493_));
  INV_X1     g24196(.I(new_n24493_), .ZN(new_n24494_));
  NAND2_X1   g24197(.A1(new_n24487_), .A2(new_n24492_), .ZN(new_n24495_));
  AOI21_X1   g24198(.A1(new_n24494_), .A2(new_n24495_), .B(new_n24491_), .ZN(new_n24496_));
  NOR2_X1    g24199(.A1(new_n24496_), .A2(new_n24490_), .ZN(new_n24497_));
  OAI21_X1   g24200(.A1(new_n24385_), .A2(new_n24418_), .B(new_n24420_), .ZN(new_n24498_));
  INV_X1     g24201(.I(new_n24498_), .ZN(new_n24499_));
  NOR2_X1    g24202(.A1(new_n24497_), .A2(new_n24499_), .ZN(new_n24500_));
  NOR3_X1    g24203(.A1(new_n24498_), .A2(new_n24496_), .A3(new_n24490_), .ZN(new_n24501_));
  NOR2_X1    g24204(.A1(new_n24500_), .A2(new_n24501_), .ZN(new_n24502_));
  NOR2_X1    g24205(.A1(new_n24502_), .A2(new_n24456_), .ZN(new_n24503_));
  INV_X1     g24206(.I(new_n24456_), .ZN(new_n24504_));
  XOR2_X1    g24207(.A1(new_n24497_), .A2(new_n24498_), .Z(new_n24505_));
  NOR2_X1    g24208(.A1(new_n24505_), .A2(new_n24504_), .ZN(new_n24506_));
  NOR2_X1    g24209(.A1(new_n24506_), .A2(new_n24503_), .ZN(new_n24507_));
  OAI21_X1   g24210(.A1(new_n24381_), .A2(new_n24426_), .B(new_n24428_), .ZN(new_n24508_));
  XOR2_X1    g24211(.A1(new_n24507_), .A2(new_n24508_), .Z(new_n24509_));
  XOR2_X1    g24212(.A1(new_n24509_), .A2(new_n24453_), .Z(new_n24510_));
  NOR2_X1    g24213(.A1(new_n24510_), .A2(\a[50] ), .ZN(new_n24511_));
  NAND2_X1   g24214(.A1(new_n24510_), .A2(\a[50] ), .ZN(new_n24512_));
  INV_X1     g24215(.I(new_n24512_), .ZN(new_n24513_));
  NOR2_X1    g24216(.A1(new_n24513_), .A2(new_n24511_), .ZN(new_n24514_));
  INV_X1     g24217(.I(new_n24431_), .ZN(new_n24515_));
  AOI21_X1   g24218(.A1(new_n24515_), .A2(new_n24437_), .B(new_n24434_), .ZN(new_n24516_));
  XOR2_X1    g24219(.A1(new_n24514_), .A2(new_n24516_), .Z(new_n24517_));
  NAND2_X1   g24220(.A1(new_n24452_), .A2(new_n24517_), .ZN(new_n24518_));
  XOR2_X1    g24221(.A1(new_n24514_), .A2(new_n24516_), .Z(new_n24519_));
  OAI21_X1   g24222(.A1(new_n24452_), .A2(new_n24519_), .B(new_n24518_), .ZN(\f[113] ));
  NOR2_X1    g24223(.A1(new_n24514_), .A2(new_n24516_), .ZN(new_n24521_));
  AOI22_X1   g24224(.A1(new_n11415_), .A2(new_n16148_), .B1(\b[61] ), .B2(new_n10145_), .ZN(new_n24522_));
  OAI21_X1   g24225(.A1(new_n24522_), .A2(\a[53] ), .B(new_n9712_), .ZN(new_n24523_));
  XOR2_X1    g24226(.A1(new_n14599_), .A2(new_n24523_), .Z(new_n24524_));
  INV_X1     g24227(.I(new_n24501_), .ZN(new_n24525_));
  AOI21_X1   g24228(.A1(new_n24525_), .A2(new_n24504_), .B(new_n24500_), .ZN(new_n24526_));
  AOI21_X1   g24229(.A1(new_n24484_), .A2(new_n24495_), .B(new_n24493_), .ZN(new_n24527_));
  AOI22_X1   g24230(.A1(new_n10969_), .A2(new_n24294_), .B1(new_n11394_), .B2(\b[58] ), .ZN(new_n24528_));
  OAI21_X1   g24231(.A1(new_n24528_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24529_));
  XOR2_X1    g24232(.A1(new_n13371_), .A2(new_n24529_), .Z(new_n24530_));
  INV_X1     g24233(.I(new_n24530_), .ZN(new_n24531_));
  NOR2_X1    g24234(.A1(new_n24459_), .A2(new_n24481_), .ZN(new_n24532_));
  AOI22_X1   g24235(.A1(new_n13078_), .A2(\b[55] ), .B1(new_n12218_), .B2(new_n12538_), .ZN(new_n24533_));
  OAI21_X1   g24236(.A1(new_n24533_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24534_));
  XOR2_X1    g24237(.A1(new_n12128_), .A2(new_n24534_), .Z(new_n24535_));
  INV_X1     g24238(.I(new_n24535_), .ZN(new_n24536_));
  OAI22_X1   g24239(.A1(new_n13880_), .A2(new_n10863_), .B1(new_n10031_), .B2(new_n13885_), .ZN(new_n24537_));
  AOI21_X1   g24240(.A1(new_n24537_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24538_));
  XNOR2_X1   g24241(.A1(new_n10866_), .A2(new_n24538_), .ZN(new_n24539_));
  NOR2_X1    g24242(.A1(new_n24463_), .A2(new_n24471_), .ZN(new_n24540_));
  NOR2_X1    g24243(.A1(new_n24540_), .A2(new_n24469_), .ZN(new_n24541_));
  NOR2_X1    g24244(.A1(new_n13476_), .A2(new_n9295_), .ZN(new_n24542_));
  XOR2_X1    g24245(.A1(new_n14736_), .A2(new_n9295_), .Z(new_n24543_));
  NAND2_X1   g24246(.A1(new_n24543_), .A2(\b[51] ), .ZN(new_n24544_));
  XOR2_X1    g24247(.A1(new_n24544_), .A2(new_n24542_), .Z(new_n24545_));
  XOR2_X1    g24248(.A1(new_n24545_), .A2(\a[50] ), .Z(new_n24546_));
  NOR2_X1    g24249(.A1(new_n24546_), .A2(new_n24400_), .ZN(new_n24547_));
  NOR2_X1    g24250(.A1(new_n24545_), .A2(new_n8624_), .ZN(new_n24548_));
  INV_X1     g24251(.I(new_n24548_), .ZN(new_n24549_));
  NAND2_X1   g24252(.A1(new_n24545_), .A2(new_n8624_), .ZN(new_n24550_));
  AOI21_X1   g24253(.A1(new_n24549_), .A2(new_n24550_), .B(new_n24401_), .ZN(new_n24551_));
  NOR2_X1    g24254(.A1(new_n24547_), .A2(new_n24551_), .ZN(new_n24552_));
  XOR2_X1    g24255(.A1(new_n24541_), .A2(new_n24552_), .Z(new_n24553_));
  NOR2_X1    g24256(.A1(new_n24553_), .A2(new_n24539_), .ZN(new_n24554_));
  INV_X1     g24257(.I(new_n24539_), .ZN(new_n24555_));
  OAI21_X1   g24258(.A1(new_n24547_), .A2(new_n24551_), .B(new_n24541_), .ZN(new_n24556_));
  OAI21_X1   g24259(.A1(new_n24540_), .A2(new_n24469_), .B(new_n24552_), .ZN(new_n24557_));
  AOI21_X1   g24260(.A1(new_n24556_), .A2(new_n24557_), .B(new_n24555_), .ZN(new_n24558_));
  NOR2_X1    g24261(.A1(new_n24554_), .A2(new_n24558_), .ZN(new_n24559_));
  XOR2_X1    g24262(.A1(new_n24559_), .A2(new_n24536_), .Z(new_n24560_));
  OAI21_X1   g24263(.A1(new_n24480_), .A2(new_n24532_), .B(new_n24560_), .ZN(new_n24561_));
  NOR2_X1    g24264(.A1(new_n24532_), .A2(new_n24480_), .ZN(new_n24562_));
  NOR2_X1    g24265(.A1(new_n24559_), .A2(new_n24536_), .ZN(new_n24563_));
  NAND2_X1   g24266(.A1(new_n24559_), .A2(new_n24536_), .ZN(new_n24564_));
  INV_X1     g24267(.I(new_n24564_), .ZN(new_n24565_));
  OAI21_X1   g24268(.A1(new_n24565_), .A2(new_n24563_), .B(new_n24562_), .ZN(new_n24566_));
  NAND2_X1   g24269(.A1(new_n24561_), .A2(new_n24566_), .ZN(new_n24567_));
  XOR2_X1    g24270(.A1(new_n24567_), .A2(new_n24531_), .Z(new_n24568_));
  NOR2_X1    g24271(.A1(new_n24568_), .A2(new_n24527_), .ZN(new_n24569_));
  INV_X1     g24272(.I(new_n24527_), .ZN(new_n24570_));
  AOI21_X1   g24273(.A1(new_n24561_), .A2(new_n24566_), .B(new_n24531_), .ZN(new_n24571_));
  NOR2_X1    g24274(.A1(new_n24567_), .A2(new_n24530_), .ZN(new_n24572_));
  NOR2_X1    g24275(.A1(new_n24572_), .A2(new_n24571_), .ZN(new_n24573_));
  NOR2_X1    g24276(.A1(new_n24573_), .A2(new_n24570_), .ZN(new_n24574_));
  NOR2_X1    g24277(.A1(new_n24569_), .A2(new_n24574_), .ZN(new_n24575_));
  XOR2_X1    g24278(.A1(new_n24575_), .A2(new_n24526_), .Z(new_n24576_));
  NOR2_X1    g24279(.A1(new_n24576_), .A2(new_n24524_), .ZN(new_n24577_));
  INV_X1     g24280(.I(new_n24526_), .ZN(new_n24578_));
  NOR2_X1    g24281(.A1(new_n24575_), .A2(new_n24578_), .ZN(new_n24579_));
  INV_X1     g24282(.I(new_n24579_), .ZN(new_n24580_));
  NAND2_X1   g24283(.A1(new_n24575_), .A2(new_n24578_), .ZN(new_n24581_));
  NAND2_X1   g24284(.A1(new_n24580_), .A2(new_n24581_), .ZN(new_n24582_));
  AOI21_X1   g24285(.A1(new_n24524_), .A2(new_n24582_), .B(new_n24577_), .ZN(new_n24583_));
  INV_X1     g24286(.I(new_n24508_), .ZN(new_n24584_));
  NOR2_X1    g24287(.A1(new_n24584_), .A2(new_n24507_), .ZN(new_n24585_));
  XOR2_X1    g24288(.A1(new_n24453_), .A2(new_n8624_), .Z(new_n24586_));
  AOI21_X1   g24289(.A1(new_n24584_), .A2(new_n24507_), .B(new_n24586_), .ZN(new_n24587_));
  NOR2_X1    g24290(.A1(new_n24587_), .A2(new_n24585_), .ZN(new_n24588_));
  INV_X1     g24291(.I(new_n24588_), .ZN(new_n24589_));
  XOR2_X1    g24292(.A1(new_n24583_), .A2(new_n24589_), .Z(new_n24590_));
  NAND2_X1   g24293(.A1(new_n24517_), .A2(new_n24590_), .ZN(new_n24591_));
  XNOR2_X1   g24294(.A1(new_n24591_), .A2(new_n24521_), .ZN(new_n24592_));
  XOR2_X1    g24295(.A1(new_n24452_), .A2(new_n24592_), .Z(\f[114] ));
  NOR2_X1    g24296(.A1(new_n24583_), .A2(new_n24589_), .ZN(new_n24594_));
  INV_X1     g24297(.I(new_n24372_), .ZN(new_n24595_));
  NOR3_X1    g24298(.A1(new_n24278_), .A2(new_n24595_), .A3(new_n24449_), .ZN(new_n24596_));
  INV_X1     g24299(.I(new_n24516_), .ZN(new_n24597_));
  NOR2_X1    g24300(.A1(new_n24590_), .A2(new_n24597_), .ZN(new_n24598_));
  NAND2_X1   g24301(.A1(new_n24590_), .A2(new_n24597_), .ZN(new_n24599_));
  AOI21_X1   g24302(.A1(new_n24514_), .A2(new_n24599_), .B(new_n24598_), .ZN(new_n24600_));
  OAI21_X1   g24303(.A1(new_n24596_), .A2(new_n24447_), .B(new_n24600_), .ZN(new_n24601_));
  NAND2_X1   g24304(.A1(new_n10145_), .A2(new_n9715_), .ZN(new_n24602_));
  NOR2_X1    g24305(.A1(new_n14596_), .A2(\a[53] ), .ZN(new_n24603_));
  AOI21_X1   g24306(.A1(new_n24602_), .A2(new_n24603_), .B(new_n9713_), .ZN(new_n24604_));
  XOR2_X1    g24307(.A1(new_n14978_), .A2(new_n24604_), .Z(new_n24605_));
  INV_X1     g24308(.I(new_n24571_), .ZN(new_n24606_));
  AOI21_X1   g24309(.A1(new_n24606_), .A2(new_n24570_), .B(new_n24572_), .ZN(new_n24607_));
  INV_X1     g24310(.I(new_n24607_), .ZN(new_n24608_));
  AOI22_X1   g24311(.A1(new_n10969_), .A2(new_n14202_), .B1(new_n11394_), .B2(\b[59] ), .ZN(new_n24609_));
  OAI21_X1   g24312(.A1(new_n24609_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24610_));
  XNOR2_X1   g24313(.A1(new_n13784_), .A2(new_n24610_), .ZN(new_n24611_));
  OAI21_X1   g24314(.A1(new_n24562_), .A2(new_n24563_), .B(new_n24564_), .ZN(new_n24612_));
  AOI22_X1   g24315(.A1(new_n13078_), .A2(\b[56] ), .B1(new_n12218_), .B2(new_n24115_), .ZN(new_n24613_));
  OAI21_X1   g24316(.A1(new_n24613_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24614_));
  XOR2_X1    g24317(.A1(new_n12546_), .A2(new_n24614_), .Z(new_n24615_));
  NAND2_X1   g24318(.A1(new_n24555_), .A2(new_n24556_), .ZN(new_n24616_));
  NAND2_X1   g24319(.A1(new_n24616_), .A2(new_n24557_), .ZN(new_n24617_));
  OAI22_X1   g24320(.A1(new_n13880_), .A2(new_n11739_), .B1(new_n10477_), .B2(new_n13885_), .ZN(new_n24618_));
  AOI21_X1   g24321(.A1(new_n24618_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24619_));
  XOR2_X1    g24322(.A1(new_n11298_), .A2(new_n24619_), .Z(new_n24620_));
  NAND2_X1   g24323(.A1(new_n24550_), .A2(new_n24401_), .ZN(new_n24621_));
  NAND2_X1   g24324(.A1(new_n24621_), .A2(new_n24549_), .ZN(new_n24622_));
  NOR2_X1    g24325(.A1(new_n13476_), .A2(new_n10025_), .ZN(new_n24623_));
  XOR2_X1    g24326(.A1(new_n14736_), .A2(new_n10025_), .Z(new_n24624_));
  NAND2_X1   g24327(.A1(new_n24624_), .A2(\b[52] ), .ZN(new_n24625_));
  XOR2_X1    g24328(.A1(new_n24625_), .A2(new_n24623_), .Z(new_n24626_));
  INV_X1     g24329(.I(new_n24626_), .ZN(new_n24627_));
  XOR2_X1    g24330(.A1(new_n24622_), .A2(new_n24627_), .Z(new_n24628_));
  NOR2_X1    g24331(.A1(new_n24622_), .A2(new_n24626_), .ZN(new_n24629_));
  NAND2_X1   g24332(.A1(new_n24622_), .A2(new_n24626_), .ZN(new_n24630_));
  INV_X1     g24333(.I(new_n24630_), .ZN(new_n24631_));
  OAI21_X1   g24334(.A1(new_n24629_), .A2(new_n24631_), .B(new_n24620_), .ZN(new_n24632_));
  OAI21_X1   g24335(.A1(new_n24620_), .A2(new_n24628_), .B(new_n24632_), .ZN(new_n24633_));
  XOR2_X1    g24336(.A1(new_n24617_), .A2(new_n24633_), .Z(new_n24634_));
  NOR2_X1    g24337(.A1(new_n24634_), .A2(new_n24615_), .ZN(new_n24635_));
  INV_X1     g24338(.I(new_n24615_), .ZN(new_n24636_));
  INV_X1     g24339(.I(new_n24617_), .ZN(new_n24637_));
  NAND2_X1   g24340(.A1(new_n24637_), .A2(new_n24633_), .ZN(new_n24638_));
  NOR2_X1    g24341(.A1(new_n24637_), .A2(new_n24633_), .ZN(new_n24639_));
  INV_X1     g24342(.I(new_n24639_), .ZN(new_n24640_));
  AOI21_X1   g24343(.A1(new_n24640_), .A2(new_n24638_), .B(new_n24636_), .ZN(new_n24641_));
  NOR2_X1    g24344(.A1(new_n24641_), .A2(new_n24635_), .ZN(new_n24642_));
  XNOR2_X1   g24345(.A1(new_n24642_), .A2(new_n24612_), .ZN(new_n24643_));
  NOR2_X1    g24346(.A1(new_n24643_), .A2(new_n24611_), .ZN(new_n24644_));
  INV_X1     g24347(.I(new_n24611_), .ZN(new_n24645_));
  NOR2_X1    g24348(.A1(new_n24642_), .A2(new_n24612_), .ZN(new_n24646_));
  INV_X1     g24349(.I(new_n24646_), .ZN(new_n24647_));
  NAND2_X1   g24350(.A1(new_n24642_), .A2(new_n24612_), .ZN(new_n24648_));
  AOI21_X1   g24351(.A1(new_n24647_), .A2(new_n24648_), .B(new_n24645_), .ZN(new_n24649_));
  NOR2_X1    g24352(.A1(new_n24644_), .A2(new_n24649_), .ZN(new_n24650_));
  NOR2_X1    g24353(.A1(new_n24650_), .A2(new_n24608_), .ZN(new_n24651_));
  INV_X1     g24354(.I(new_n24650_), .ZN(new_n24652_));
  NOR2_X1    g24355(.A1(new_n24652_), .A2(new_n24607_), .ZN(new_n24653_));
  NOR2_X1    g24356(.A1(new_n24653_), .A2(new_n24651_), .ZN(new_n24654_));
  NOR2_X1    g24357(.A1(new_n24654_), .A2(new_n24605_), .ZN(new_n24655_));
  INV_X1     g24358(.I(new_n24605_), .ZN(new_n24656_));
  XOR2_X1    g24359(.A1(new_n24650_), .A2(new_n24607_), .Z(new_n24657_));
  NOR2_X1    g24360(.A1(new_n24657_), .A2(new_n24656_), .ZN(new_n24658_));
  NOR2_X1    g24361(.A1(new_n24655_), .A2(new_n24658_), .ZN(new_n24659_));
  INV_X1     g24362(.I(new_n24659_), .ZN(new_n24660_));
  OAI21_X1   g24363(.A1(new_n24524_), .A2(new_n24579_), .B(new_n24581_), .ZN(new_n24661_));
  NAND2_X1   g24364(.A1(new_n24660_), .A2(new_n24661_), .ZN(new_n24662_));
  XOR2_X1    g24365(.A1(new_n24601_), .A2(new_n24662_), .Z(new_n24663_));
  XOR2_X1    g24366(.A1(new_n24663_), .A2(new_n24594_), .Z(\f[115] ));
  INV_X1     g24367(.I(new_n24594_), .ZN(new_n24665_));
  NOR2_X1    g24368(.A1(new_n24665_), .A2(new_n24659_), .ZN(new_n24666_));
  INV_X1     g24369(.I(new_n24666_), .ZN(new_n24667_));
  OAI21_X1   g24370(.A1(new_n24594_), .A2(new_n24660_), .B(new_n24661_), .ZN(new_n24668_));
  OAI21_X1   g24371(.A1(new_n24601_), .A2(new_n24668_), .B(new_n24667_), .ZN(new_n24669_));
  OAI21_X1   g24372(.A1(new_n9713_), .A2(new_n10137_), .B(new_n16487_), .ZN(new_n24670_));
  AOI22_X1   g24373(.A1(new_n10969_), .A2(new_n14590_), .B1(new_n11394_), .B2(\b[60] ), .ZN(new_n24671_));
  OAI21_X1   g24374(.A1(new_n24671_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24672_));
  XNOR2_X1   g24375(.A1(new_n14213_), .A2(new_n24672_), .ZN(new_n24673_));
  AOI21_X1   g24376(.A1(new_n24636_), .A2(new_n24638_), .B(new_n24639_), .ZN(new_n24674_));
  INV_X1     g24377(.I(new_n24674_), .ZN(new_n24675_));
  OAI21_X1   g24378(.A1(new_n24620_), .A2(new_n24629_), .B(new_n24630_), .ZN(new_n24676_));
  NOR2_X1    g24379(.A1(new_n13476_), .A2(new_n10031_), .ZN(new_n24677_));
  XOR2_X1    g24380(.A1(new_n14736_), .A2(new_n10031_), .Z(new_n24678_));
  NAND2_X1   g24381(.A1(new_n24678_), .A2(\b[53] ), .ZN(new_n24679_));
  XOR2_X1    g24382(.A1(new_n24679_), .A2(new_n24677_), .Z(new_n24680_));
  NOR2_X1    g24383(.A1(new_n24627_), .A2(new_n24680_), .ZN(new_n24681_));
  INV_X1     g24384(.I(new_n24680_), .ZN(new_n24682_));
  NOR2_X1    g24385(.A1(new_n24682_), .A2(new_n24626_), .ZN(new_n24683_));
  NOR2_X1    g24386(.A1(new_n24681_), .A2(new_n24683_), .ZN(new_n24684_));
  INV_X1     g24387(.I(new_n24684_), .ZN(new_n24685_));
  XOR2_X1    g24388(.A1(new_n24626_), .A2(new_n24680_), .Z(new_n24686_));
  NOR2_X1    g24389(.A1(new_n24676_), .A2(new_n24686_), .ZN(new_n24687_));
  AOI21_X1   g24390(.A1(new_n24676_), .A2(new_n24685_), .B(new_n24687_), .ZN(new_n24688_));
  AOI22_X1   g24391(.A1(new_n13078_), .A2(\b[57] ), .B1(new_n12218_), .B2(new_n13363_), .ZN(new_n24689_));
  OAI21_X1   g24392(.A1(new_n24689_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24690_));
  XNOR2_X1   g24393(.A1(new_n12969_), .A2(new_n24690_), .ZN(new_n24691_));
  OAI22_X1   g24394(.A1(new_n13880_), .A2(new_n11745_), .B1(new_n10862_), .B2(new_n13885_), .ZN(new_n24692_));
  AOI21_X1   g24395(.A1(new_n24692_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24693_));
  XNOR2_X1   g24396(.A1(new_n11748_), .A2(new_n24693_), .ZN(new_n24694_));
  XNOR2_X1   g24397(.A1(new_n24691_), .A2(new_n24694_), .ZN(new_n24695_));
  NOR2_X1    g24398(.A1(new_n24695_), .A2(new_n24688_), .ZN(new_n24696_));
  INV_X1     g24399(.I(new_n24688_), .ZN(new_n24697_));
  NOR2_X1    g24400(.A1(new_n24691_), .A2(new_n24694_), .ZN(new_n24698_));
  INV_X1     g24401(.I(new_n24698_), .ZN(new_n24699_));
  NAND2_X1   g24402(.A1(new_n24691_), .A2(new_n24694_), .ZN(new_n24700_));
  AOI21_X1   g24403(.A1(new_n24699_), .A2(new_n24700_), .B(new_n24697_), .ZN(new_n24701_));
  NOR2_X1    g24404(.A1(new_n24696_), .A2(new_n24701_), .ZN(new_n24702_));
  NOR2_X1    g24405(.A1(new_n24702_), .A2(new_n24675_), .ZN(new_n24703_));
  INV_X1     g24406(.I(new_n24702_), .ZN(new_n24704_));
  NOR2_X1    g24407(.A1(new_n24704_), .A2(new_n24674_), .ZN(new_n24705_));
  NOR2_X1    g24408(.A1(new_n24705_), .A2(new_n24703_), .ZN(new_n24706_));
  NOR2_X1    g24409(.A1(new_n24706_), .A2(new_n24673_), .ZN(new_n24707_));
  INV_X1     g24410(.I(new_n24673_), .ZN(new_n24708_));
  XOR2_X1    g24411(.A1(new_n24702_), .A2(new_n24674_), .Z(new_n24709_));
  NOR2_X1    g24412(.A1(new_n24709_), .A2(new_n24708_), .ZN(new_n24710_));
  NOR2_X1    g24413(.A1(new_n24707_), .A2(new_n24710_), .ZN(new_n24711_));
  OAI21_X1   g24414(.A1(new_n24611_), .A2(new_n24646_), .B(new_n24648_), .ZN(new_n24712_));
  XOR2_X1    g24415(.A1(new_n24711_), .A2(new_n24712_), .Z(new_n24713_));
  XOR2_X1    g24416(.A1(new_n24713_), .A2(new_n24670_), .Z(new_n24714_));
  NOR2_X1    g24417(.A1(new_n24714_), .A2(\a[53] ), .ZN(new_n24715_));
  NAND2_X1   g24418(.A1(new_n24714_), .A2(\a[53] ), .ZN(new_n24716_));
  INV_X1     g24419(.I(new_n24716_), .ZN(new_n24717_));
  NOR2_X1    g24420(.A1(new_n24717_), .A2(new_n24715_), .ZN(new_n24718_));
  INV_X1     g24421(.I(new_n24651_), .ZN(new_n24719_));
  AOI21_X1   g24422(.A1(new_n24719_), .A2(new_n24656_), .B(new_n24653_), .ZN(new_n24720_));
  XOR2_X1    g24423(.A1(new_n24718_), .A2(new_n24720_), .Z(new_n24721_));
  NAND2_X1   g24424(.A1(new_n24669_), .A2(new_n24721_), .ZN(new_n24722_));
  INV_X1     g24425(.I(new_n24600_), .ZN(new_n24723_));
  AOI21_X1   g24426(.A1(new_n24451_), .A2(new_n24448_), .B(new_n24723_), .ZN(new_n24724_));
  INV_X1     g24427(.I(new_n24668_), .ZN(new_n24725_));
  AOI21_X1   g24428(.A1(new_n24724_), .A2(new_n24725_), .B(new_n24666_), .ZN(new_n24726_));
  INV_X1     g24429(.I(new_n24718_), .ZN(new_n24727_));
  INV_X1     g24430(.I(new_n24720_), .ZN(new_n24728_));
  NAND2_X1   g24431(.A1(new_n24727_), .A2(new_n24728_), .ZN(new_n24729_));
  NAND2_X1   g24432(.A1(new_n24718_), .A2(new_n24720_), .ZN(new_n24730_));
  NAND2_X1   g24433(.A1(new_n24729_), .A2(new_n24730_), .ZN(new_n24731_));
  NAND2_X1   g24434(.A1(new_n24726_), .A2(new_n24731_), .ZN(new_n24732_));
  NAND2_X1   g24435(.A1(new_n24732_), .A2(new_n24722_), .ZN(\f[116] ));
  INV_X1     g24436(.I(new_n24712_), .ZN(new_n24734_));
  NOR2_X1    g24437(.A1(new_n24711_), .A2(new_n24734_), .ZN(new_n24735_));
  XOR2_X1    g24438(.A1(new_n24670_), .A2(new_n9718_), .Z(new_n24736_));
  AOI21_X1   g24439(.A1(new_n24711_), .A2(new_n24734_), .B(new_n24736_), .ZN(new_n24737_));
  NOR2_X1    g24440(.A1(new_n24737_), .A2(new_n24735_), .ZN(new_n24738_));
  INV_X1     g24441(.I(new_n24703_), .ZN(new_n24739_));
  AOI21_X1   g24442(.A1(new_n24708_), .A2(new_n24739_), .B(new_n24705_), .ZN(new_n24740_));
  AOI22_X1   g24443(.A1(new_n10969_), .A2(new_n16148_), .B1(new_n11394_), .B2(\b[61] ), .ZN(new_n24741_));
  OAI21_X1   g24444(.A1(new_n24741_), .A2(\a[56] ), .B(new_n10975_), .ZN(new_n24742_));
  XOR2_X1    g24445(.A1(new_n14599_), .A2(new_n24742_), .Z(new_n24743_));
  AOI21_X1   g24446(.A1(new_n24697_), .A2(new_n24700_), .B(new_n24698_), .ZN(new_n24744_));
  INV_X1     g24447(.I(new_n24744_), .ZN(new_n24745_));
  AOI22_X1   g24448(.A1(new_n13078_), .A2(\b[58] ), .B1(new_n12218_), .B2(new_n24294_), .ZN(new_n24746_));
  OAI21_X1   g24449(.A1(new_n24746_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24747_));
  NOR2_X1    g24450(.A1(new_n13371_), .A2(new_n24747_), .ZN(new_n24748_));
  NAND2_X1   g24451(.A1(new_n13371_), .A2(new_n24747_), .ZN(new_n24749_));
  INV_X1     g24452(.I(new_n24749_), .ZN(new_n24750_));
  INV_X1     g24453(.I(new_n24681_), .ZN(new_n24751_));
  AOI21_X1   g24454(.A1(new_n24676_), .A2(new_n24751_), .B(new_n24683_), .ZN(new_n24752_));
  OAI22_X1   g24455(.A1(new_n13880_), .A2(new_n12537_), .B1(new_n11738_), .B2(new_n13885_), .ZN(new_n24753_));
  AOI21_X1   g24456(.A1(new_n24753_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24754_));
  XNOR2_X1   g24457(.A1(new_n12128_), .A2(new_n24754_), .ZN(new_n24755_));
  NOR2_X1    g24458(.A1(new_n13476_), .A2(new_n10477_), .ZN(new_n24756_));
  XOR2_X1    g24459(.A1(new_n14736_), .A2(new_n10477_), .Z(new_n24757_));
  NAND2_X1   g24460(.A1(new_n24757_), .A2(\b[54] ), .ZN(new_n24758_));
  XOR2_X1    g24461(.A1(new_n24758_), .A2(new_n24756_), .Z(new_n24759_));
  XOR2_X1    g24462(.A1(new_n24759_), .A2(\a[53] ), .Z(new_n24760_));
  NOR2_X1    g24463(.A1(new_n24760_), .A2(new_n24680_), .ZN(new_n24761_));
  NOR2_X1    g24464(.A1(new_n24759_), .A2(new_n9718_), .ZN(new_n24762_));
  INV_X1     g24465(.I(new_n24762_), .ZN(new_n24763_));
  NAND2_X1   g24466(.A1(new_n24759_), .A2(new_n9718_), .ZN(new_n24764_));
  AOI21_X1   g24467(.A1(new_n24763_), .A2(new_n24764_), .B(new_n24682_), .ZN(new_n24765_));
  NOR2_X1    g24468(.A1(new_n24761_), .A2(new_n24765_), .ZN(new_n24766_));
  XOR2_X1    g24469(.A1(new_n24755_), .A2(new_n24766_), .Z(new_n24767_));
  NOR2_X1    g24470(.A1(new_n24767_), .A2(new_n24752_), .ZN(new_n24768_));
  INV_X1     g24471(.I(new_n24752_), .ZN(new_n24769_));
  INV_X1     g24472(.I(new_n24755_), .ZN(new_n24770_));
  NOR2_X1    g24473(.A1(new_n24770_), .A2(new_n24766_), .ZN(new_n24771_));
  INV_X1     g24474(.I(new_n24771_), .ZN(new_n24772_));
  NAND2_X1   g24475(.A1(new_n24770_), .A2(new_n24766_), .ZN(new_n24773_));
  AOI21_X1   g24476(.A1(new_n24772_), .A2(new_n24773_), .B(new_n24769_), .ZN(new_n24774_));
  NOR2_X1    g24477(.A1(new_n24774_), .A2(new_n24768_), .ZN(new_n24775_));
  NOR3_X1    g24478(.A1(new_n24775_), .A2(new_n24748_), .A3(new_n24750_), .ZN(new_n24776_));
  NOR2_X1    g24479(.A1(new_n24750_), .A2(new_n24748_), .ZN(new_n24777_));
  NOR3_X1    g24480(.A1(new_n24777_), .A2(new_n24768_), .A3(new_n24774_), .ZN(new_n24778_));
  OAI21_X1   g24481(.A1(new_n24776_), .A2(new_n24778_), .B(new_n24745_), .ZN(new_n24779_));
  XOR2_X1    g24482(.A1(new_n24775_), .A2(new_n24777_), .Z(new_n24780_));
  OAI21_X1   g24483(.A1(new_n24780_), .A2(new_n24745_), .B(new_n24779_), .ZN(new_n24781_));
  INV_X1     g24484(.I(new_n24781_), .ZN(new_n24782_));
  NOR2_X1    g24485(.A1(new_n24782_), .A2(new_n24743_), .ZN(new_n24783_));
  INV_X1     g24486(.I(new_n24783_), .ZN(new_n24784_));
  NAND2_X1   g24487(.A1(new_n24782_), .A2(new_n24743_), .ZN(new_n24785_));
  AOI21_X1   g24488(.A1(new_n24784_), .A2(new_n24785_), .B(new_n24740_), .ZN(new_n24786_));
  XNOR2_X1   g24489(.A1(new_n24781_), .A2(new_n24743_), .ZN(new_n24787_));
  AOI21_X1   g24490(.A1(new_n24740_), .A2(new_n24787_), .B(new_n24786_), .ZN(new_n24788_));
  XNOR2_X1   g24491(.A1(new_n24788_), .A2(new_n24738_), .ZN(new_n24789_));
  INV_X1     g24492(.I(new_n24789_), .ZN(new_n24790_));
  NAND2_X1   g24493(.A1(new_n24721_), .A2(new_n24790_), .ZN(new_n24791_));
  XOR2_X1    g24494(.A1(new_n24791_), .A2(new_n24729_), .Z(new_n24792_));
  XOR2_X1    g24495(.A1(new_n24669_), .A2(new_n24792_), .Z(\f[117] ));
  NAND2_X1   g24496(.A1(new_n24788_), .A2(new_n24738_), .ZN(new_n24794_));
  NOR2_X1    g24497(.A1(new_n24790_), .A2(new_n24728_), .ZN(new_n24795_));
  AOI21_X1   g24498(.A1(new_n24728_), .A2(new_n24790_), .B(new_n24727_), .ZN(new_n24796_));
  NOR2_X1    g24499(.A1(new_n24796_), .A2(new_n24795_), .ZN(new_n24797_));
  NAND2_X1   g24500(.A1(new_n24669_), .A2(new_n24797_), .ZN(new_n24798_));
  NAND2_X1   g24501(.A1(new_n11394_), .A2(new_n10967_), .ZN(new_n24799_));
  NOR2_X1    g24502(.A1(new_n14596_), .A2(\a[56] ), .ZN(new_n24800_));
  AOI21_X1   g24503(.A1(new_n24799_), .A2(new_n24800_), .B(new_n10964_), .ZN(new_n24801_));
  XOR2_X1    g24504(.A1(new_n14978_), .A2(new_n24801_), .Z(new_n24802_));
  NOR2_X1    g24505(.A1(new_n24776_), .A2(new_n24744_), .ZN(new_n24803_));
  NOR2_X1    g24506(.A1(new_n24803_), .A2(new_n24778_), .ZN(new_n24804_));
  AOI22_X1   g24507(.A1(new_n13078_), .A2(\b[59] ), .B1(new_n12218_), .B2(new_n14202_), .ZN(new_n24805_));
  OAI21_X1   g24508(.A1(new_n24805_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24806_));
  XNOR2_X1   g24509(.A1(new_n13784_), .A2(new_n24806_), .ZN(new_n24807_));
  OAI21_X1   g24510(.A1(new_n24752_), .A2(new_n24771_), .B(new_n24773_), .ZN(new_n24808_));
  OAI22_X1   g24511(.A1(new_n13880_), .A2(new_n12543_), .B1(new_n11744_), .B2(new_n13885_), .ZN(new_n24809_));
  AOI21_X1   g24512(.A1(new_n24809_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24810_));
  XNOR2_X1   g24513(.A1(new_n12546_), .A2(new_n24810_), .ZN(new_n24811_));
  NAND2_X1   g24514(.A1(new_n24764_), .A2(new_n24682_), .ZN(new_n24812_));
  NAND2_X1   g24515(.A1(new_n24812_), .A2(new_n24763_), .ZN(new_n24813_));
  NOR2_X1    g24516(.A1(new_n13476_), .A2(new_n10862_), .ZN(new_n24814_));
  XOR2_X1    g24517(.A1(new_n14736_), .A2(new_n10862_), .Z(new_n24815_));
  NAND2_X1   g24518(.A1(new_n24815_), .A2(\b[55] ), .ZN(new_n24816_));
  XOR2_X1    g24519(.A1(new_n24816_), .A2(new_n24814_), .Z(new_n24817_));
  INV_X1     g24520(.I(new_n24817_), .ZN(new_n24818_));
  XOR2_X1    g24521(.A1(new_n24813_), .A2(new_n24818_), .Z(new_n24819_));
  NOR2_X1    g24522(.A1(new_n24811_), .A2(new_n24819_), .ZN(new_n24820_));
  NOR2_X1    g24523(.A1(new_n24813_), .A2(new_n24817_), .ZN(new_n24821_));
  INV_X1     g24524(.I(new_n24821_), .ZN(new_n24822_));
  NAND2_X1   g24525(.A1(new_n24813_), .A2(new_n24817_), .ZN(new_n24823_));
  NAND2_X1   g24526(.A1(new_n24822_), .A2(new_n24823_), .ZN(new_n24824_));
  AOI21_X1   g24527(.A1(new_n24811_), .A2(new_n24824_), .B(new_n24820_), .ZN(new_n24825_));
  XNOR2_X1   g24528(.A1(new_n24825_), .A2(new_n24808_), .ZN(new_n24826_));
  NOR2_X1    g24529(.A1(new_n24825_), .A2(new_n24808_), .ZN(new_n24827_));
  AND2_X2    g24530(.A1(new_n24825_), .A2(new_n24808_), .Z(new_n24828_));
  OAI21_X1   g24531(.A1(new_n24828_), .A2(new_n24827_), .B(new_n24807_), .ZN(new_n24829_));
  OAI21_X1   g24532(.A1(new_n24807_), .A2(new_n24826_), .B(new_n24829_), .ZN(new_n24830_));
  NAND2_X1   g24533(.A1(new_n24830_), .A2(new_n24804_), .ZN(new_n24831_));
  NOR2_X1    g24534(.A1(new_n24830_), .A2(new_n24804_), .ZN(new_n24832_));
  INV_X1     g24535(.I(new_n24832_), .ZN(new_n24833_));
  AOI21_X1   g24536(.A1(new_n24833_), .A2(new_n24831_), .B(new_n24802_), .ZN(new_n24834_));
  INV_X1     g24537(.I(new_n24802_), .ZN(new_n24835_));
  XNOR2_X1   g24538(.A1(new_n24830_), .A2(new_n24804_), .ZN(new_n24836_));
  NOR2_X1    g24539(.A1(new_n24836_), .A2(new_n24835_), .ZN(new_n24837_));
  NOR2_X1    g24540(.A1(new_n24837_), .A2(new_n24834_), .ZN(new_n24838_));
  INV_X1     g24541(.I(new_n24740_), .ZN(new_n24839_));
  AOI21_X1   g24542(.A1(new_n24839_), .A2(new_n24785_), .B(new_n24783_), .ZN(new_n24840_));
  NOR2_X1    g24543(.A1(new_n24838_), .A2(new_n24840_), .ZN(new_n24841_));
  XOR2_X1    g24544(.A1(new_n24798_), .A2(new_n24841_), .Z(new_n24842_));
  XOR2_X1    g24545(.A1(new_n24842_), .A2(new_n24794_), .Z(\f[118] ));
  NOR2_X1    g24546(.A1(new_n24794_), .A2(new_n24838_), .ZN(new_n24844_));
  INV_X1     g24547(.I(new_n24797_), .ZN(new_n24845_));
  AOI21_X1   g24548(.A1(new_n24794_), .A2(new_n24838_), .B(new_n24840_), .ZN(new_n24846_));
  INV_X1     g24549(.I(new_n24846_), .ZN(new_n24847_));
  NOR3_X1    g24550(.A1(new_n24726_), .A2(new_n24845_), .A3(new_n24847_), .ZN(new_n24848_));
  NOR2_X1    g24551(.A1(new_n24848_), .A2(new_n24844_), .ZN(new_n24849_));
  OAI21_X1   g24552(.A1(new_n10964_), .A2(new_n11401_), .B(new_n16487_), .ZN(new_n24850_));
  AOI22_X1   g24553(.A1(new_n13078_), .A2(\b[60] ), .B1(new_n12218_), .B2(new_n14590_), .ZN(new_n24851_));
  OAI21_X1   g24554(.A1(new_n24851_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24852_));
  XNOR2_X1   g24555(.A1(new_n14213_), .A2(new_n24852_), .ZN(new_n24853_));
  OAI22_X1   g24556(.A1(new_n13880_), .A2(new_n13362_), .B1(new_n12536_), .B2(new_n13885_), .ZN(new_n24854_));
  AOI21_X1   g24557(.A1(new_n24854_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24855_));
  XOR2_X1    g24558(.A1(new_n12969_), .A2(new_n24855_), .Z(new_n24856_));
  INV_X1     g24559(.I(new_n24856_), .ZN(new_n24857_));
  NOR2_X1    g24560(.A1(new_n13476_), .A2(new_n11738_), .ZN(new_n24858_));
  XOR2_X1    g24561(.A1(new_n14736_), .A2(new_n11738_), .Z(new_n24859_));
  NAND2_X1   g24562(.A1(new_n24859_), .A2(\b[56] ), .ZN(new_n24860_));
  XOR2_X1    g24563(.A1(new_n24860_), .A2(new_n24858_), .Z(new_n24861_));
  NOR2_X1    g24564(.A1(new_n24818_), .A2(new_n24861_), .ZN(new_n24862_));
  INV_X1     g24565(.I(new_n24861_), .ZN(new_n24863_));
  NOR2_X1    g24566(.A1(new_n24863_), .A2(new_n24817_), .ZN(new_n24864_));
  OAI21_X1   g24567(.A1(new_n24862_), .A2(new_n24864_), .B(new_n24857_), .ZN(new_n24865_));
  XNOR2_X1   g24568(.A1(new_n24817_), .A2(new_n24861_), .ZN(new_n24866_));
  NAND2_X1   g24569(.A1(new_n24856_), .A2(new_n24866_), .ZN(new_n24867_));
  OR2_X2     g24570(.A1(new_n24811_), .A2(new_n24821_), .Z(new_n24868_));
  AOI22_X1   g24571(.A1(new_n24823_), .A2(new_n24868_), .B1(new_n24865_), .B2(new_n24867_), .ZN(new_n24869_));
  NAND2_X1   g24572(.A1(new_n24865_), .A2(new_n24867_), .ZN(new_n24870_));
  NAND2_X1   g24573(.A1(new_n24868_), .A2(new_n24823_), .ZN(new_n24871_));
  NOR2_X1    g24574(.A1(new_n24871_), .A2(new_n24870_), .ZN(new_n24872_));
  NOR2_X1    g24575(.A1(new_n24872_), .A2(new_n24869_), .ZN(new_n24873_));
  NOR2_X1    g24576(.A1(new_n24873_), .A2(new_n24853_), .ZN(new_n24874_));
  XOR2_X1    g24577(.A1(new_n24871_), .A2(new_n24870_), .Z(new_n24875_));
  AOI21_X1   g24578(.A1(new_n24853_), .A2(new_n24875_), .B(new_n24874_), .ZN(new_n24876_));
  NOR2_X1    g24579(.A1(new_n24827_), .A2(new_n24807_), .ZN(new_n24877_));
  NOR2_X1    g24580(.A1(new_n24877_), .A2(new_n24828_), .ZN(new_n24878_));
  XNOR2_X1   g24581(.A1(new_n24876_), .A2(new_n24878_), .ZN(new_n24879_));
  XOR2_X1    g24582(.A1(new_n24879_), .A2(new_n24850_), .Z(new_n24880_));
  NOR2_X1    g24583(.A1(new_n24880_), .A2(\a[56] ), .ZN(new_n24881_));
  NAND2_X1   g24584(.A1(new_n24880_), .A2(\a[56] ), .ZN(new_n24882_));
  INV_X1     g24585(.I(new_n24882_), .ZN(new_n24883_));
  NOR2_X1    g24586(.A1(new_n24883_), .A2(new_n24881_), .ZN(new_n24884_));
  AOI21_X1   g24587(.A1(new_n24835_), .A2(new_n24831_), .B(new_n24832_), .ZN(new_n24885_));
  XOR2_X1    g24588(.A1(new_n24884_), .A2(new_n24885_), .Z(new_n24886_));
  INV_X1     g24589(.I(new_n24884_), .ZN(new_n24887_));
  INV_X1     g24590(.I(new_n24885_), .ZN(new_n24888_));
  NAND2_X1   g24591(.A1(new_n24887_), .A2(new_n24888_), .ZN(new_n24889_));
  NAND2_X1   g24592(.A1(new_n24884_), .A2(new_n24885_), .ZN(new_n24890_));
  NAND2_X1   g24593(.A1(new_n24889_), .A2(new_n24890_), .ZN(new_n24891_));
  MUX2_X1    g24594(.I0(new_n24886_), .I1(new_n24891_), .S(new_n24849_), .Z(\f[119] ));
  INV_X1     g24595(.I(new_n24869_), .ZN(new_n24893_));
  OAI21_X1   g24596(.A1(new_n24853_), .A2(new_n24872_), .B(new_n24893_), .ZN(new_n24894_));
  INV_X1     g24597(.I(new_n24894_), .ZN(new_n24895_));
  AOI22_X1   g24598(.A1(new_n13078_), .A2(\b[61] ), .B1(new_n12218_), .B2(new_n16148_), .ZN(new_n24896_));
  OAI21_X1   g24599(.A1(new_n24896_), .A2(\a[59] ), .B(new_n12214_), .ZN(new_n24897_));
  NOR2_X1    g24600(.A1(new_n14599_), .A2(new_n24897_), .ZN(new_n24898_));
  NAND2_X1   g24601(.A1(new_n14599_), .A2(new_n24897_), .ZN(new_n24899_));
  INV_X1     g24602(.I(new_n24899_), .ZN(new_n24900_));
  NOR2_X1    g24603(.A1(new_n24900_), .A2(new_n24898_), .ZN(new_n24901_));
  INV_X1     g24604(.I(new_n24901_), .ZN(new_n24902_));
  NOR2_X1    g24605(.A1(new_n24856_), .A2(new_n24864_), .ZN(new_n24903_));
  NOR2_X1    g24606(.A1(new_n24903_), .A2(new_n24862_), .ZN(new_n24904_));
  OAI22_X1   g24607(.A1(new_n13880_), .A2(new_n13368_), .B1(new_n12542_), .B2(new_n13885_), .ZN(new_n24905_));
  AOI21_X1   g24608(.A1(new_n24905_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24906_));
  XNOR2_X1   g24609(.A1(new_n13371_), .A2(new_n24906_), .ZN(new_n24907_));
  NOR2_X1    g24610(.A1(new_n13476_), .A2(new_n11744_), .ZN(new_n24908_));
  XOR2_X1    g24611(.A1(new_n14736_), .A2(new_n11744_), .Z(new_n24909_));
  NAND2_X1   g24612(.A1(new_n24909_), .A2(\b[57] ), .ZN(new_n24910_));
  XOR2_X1    g24613(.A1(new_n24910_), .A2(new_n24908_), .Z(new_n24911_));
  NOR2_X1    g24614(.A1(new_n24911_), .A2(new_n10973_), .ZN(new_n24912_));
  INV_X1     g24615(.I(new_n24912_), .ZN(new_n24913_));
  NAND2_X1   g24616(.A1(new_n24911_), .A2(new_n10973_), .ZN(new_n24914_));
  AOI21_X1   g24617(.A1(new_n24913_), .A2(new_n24914_), .B(new_n24817_), .ZN(new_n24915_));
  XOR2_X1    g24618(.A1(new_n24911_), .A2(\a[56] ), .Z(new_n24916_));
  NOR2_X1    g24619(.A1(new_n24916_), .A2(new_n24818_), .ZN(new_n24917_));
  NOR2_X1    g24620(.A1(new_n24917_), .A2(new_n24915_), .ZN(new_n24918_));
  XNOR2_X1   g24621(.A1(new_n24907_), .A2(new_n24918_), .ZN(new_n24919_));
  NOR2_X1    g24622(.A1(new_n24919_), .A2(new_n24904_), .ZN(new_n24920_));
  INV_X1     g24623(.I(new_n24904_), .ZN(new_n24921_));
  NOR2_X1    g24624(.A1(new_n24907_), .A2(new_n24918_), .ZN(new_n24922_));
  INV_X1     g24625(.I(new_n24922_), .ZN(new_n24923_));
  NAND2_X1   g24626(.A1(new_n24907_), .A2(new_n24918_), .ZN(new_n24924_));
  AOI21_X1   g24627(.A1(new_n24923_), .A2(new_n24924_), .B(new_n24921_), .ZN(new_n24925_));
  NOR2_X1    g24628(.A1(new_n24920_), .A2(new_n24925_), .ZN(new_n24926_));
  NOR2_X1    g24629(.A1(new_n24902_), .A2(new_n24926_), .ZN(new_n24927_));
  INV_X1     g24630(.I(new_n24927_), .ZN(new_n24928_));
  NAND2_X1   g24631(.A1(new_n24902_), .A2(new_n24926_), .ZN(new_n24929_));
  AOI21_X1   g24632(.A1(new_n24928_), .A2(new_n24929_), .B(new_n24895_), .ZN(new_n24930_));
  XNOR2_X1   g24633(.A1(new_n24926_), .A2(new_n24901_), .ZN(new_n24931_));
  AOI21_X1   g24634(.A1(new_n24895_), .A2(new_n24931_), .B(new_n24930_), .ZN(new_n24932_));
  NOR2_X1    g24635(.A1(new_n24876_), .A2(new_n24878_), .ZN(new_n24933_));
  NAND2_X1   g24636(.A1(new_n24876_), .A2(new_n24878_), .ZN(new_n24934_));
  XOR2_X1    g24637(.A1(new_n24850_), .A2(\a[56] ), .Z(new_n24935_));
  AOI21_X1   g24638(.A1(new_n24934_), .A2(new_n24935_), .B(new_n24933_), .ZN(new_n24936_));
  XNOR2_X1   g24639(.A1(new_n24932_), .A2(new_n24936_), .ZN(new_n24937_));
  INV_X1     g24640(.I(new_n24937_), .ZN(new_n24938_));
  NAND2_X1   g24641(.A1(new_n24886_), .A2(new_n24938_), .ZN(new_n24939_));
  XNOR2_X1   g24642(.A1(new_n24939_), .A2(new_n24889_), .ZN(new_n24940_));
  XOR2_X1    g24643(.A1(new_n24849_), .A2(new_n24940_), .Z(\f[120] ));
  NAND2_X1   g24644(.A1(new_n24932_), .A2(new_n24936_), .ZN(new_n24942_));
  INV_X1     g24645(.I(new_n24844_), .ZN(new_n24943_));
  NAND3_X1   g24646(.A1(new_n24669_), .A2(new_n24797_), .A3(new_n24846_), .ZN(new_n24944_));
  NOR2_X1    g24647(.A1(new_n24938_), .A2(new_n24888_), .ZN(new_n24945_));
  AOI21_X1   g24648(.A1(new_n24888_), .A2(new_n24938_), .B(new_n24887_), .ZN(new_n24946_));
  NOR2_X1    g24649(.A1(new_n24946_), .A2(new_n24945_), .ZN(new_n24947_));
  INV_X1     g24650(.I(new_n24947_), .ZN(new_n24948_));
  AOI21_X1   g24651(.A1(new_n24944_), .A2(new_n24943_), .B(new_n24948_), .ZN(new_n24949_));
  NAND2_X1   g24652(.A1(new_n13078_), .A2(new_n12216_), .ZN(new_n24950_));
  NOR2_X1    g24653(.A1(new_n14596_), .A2(\a[59] ), .ZN(new_n24951_));
  AOI21_X1   g24654(.A1(new_n24950_), .A2(new_n24951_), .B(new_n12643_), .ZN(new_n24952_));
  XOR2_X1    g24655(.A1(new_n14978_), .A2(new_n24952_), .Z(new_n24953_));
  INV_X1     g24656(.I(new_n24953_), .ZN(new_n24954_));
  NAND2_X1   g24657(.A1(new_n24924_), .A2(new_n24921_), .ZN(new_n24955_));
  NAND2_X1   g24658(.A1(new_n24955_), .A2(new_n24923_), .ZN(new_n24956_));
  OAI22_X1   g24659(.A1(new_n13880_), .A2(new_n14201_), .B1(new_n12970_), .B2(new_n13885_), .ZN(new_n24957_));
  AOI21_X1   g24660(.A1(new_n24957_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n24958_));
  XOR2_X1    g24661(.A1(new_n13784_), .A2(new_n24958_), .Z(new_n24959_));
  NAND2_X1   g24662(.A1(new_n24914_), .A2(new_n24818_), .ZN(new_n24960_));
  NAND2_X1   g24663(.A1(new_n24960_), .A2(new_n24913_), .ZN(new_n24961_));
  NOR2_X1    g24664(.A1(new_n13476_), .A2(new_n12536_), .ZN(new_n24962_));
  XOR2_X1    g24665(.A1(new_n14736_), .A2(new_n12536_), .Z(new_n24963_));
  NAND2_X1   g24666(.A1(new_n24963_), .A2(\b[58] ), .ZN(new_n24964_));
  XOR2_X1    g24667(.A1(new_n24964_), .A2(new_n24962_), .Z(new_n24965_));
  INV_X1     g24668(.I(new_n24965_), .ZN(new_n24966_));
  XOR2_X1    g24669(.A1(new_n24961_), .A2(new_n24966_), .Z(new_n24967_));
  OR2_X2     g24670(.A1(new_n24959_), .A2(new_n24967_), .Z(new_n24968_));
  NOR2_X1    g24671(.A1(new_n24961_), .A2(new_n24965_), .ZN(new_n24969_));
  NAND2_X1   g24672(.A1(new_n24961_), .A2(new_n24965_), .ZN(new_n24970_));
  INV_X1     g24673(.I(new_n24970_), .ZN(new_n24971_));
  OAI21_X1   g24674(.A1(new_n24969_), .A2(new_n24971_), .B(new_n24959_), .ZN(new_n24972_));
  AOI21_X1   g24675(.A1(new_n24968_), .A2(new_n24972_), .B(new_n24956_), .ZN(new_n24973_));
  NAND2_X1   g24676(.A1(new_n24968_), .A2(new_n24972_), .ZN(new_n24974_));
  AOI21_X1   g24677(.A1(new_n24923_), .A2(new_n24955_), .B(new_n24974_), .ZN(new_n24975_));
  OAI21_X1   g24678(.A1(new_n24973_), .A2(new_n24975_), .B(new_n24954_), .ZN(new_n24976_));
  XNOR2_X1   g24679(.A1(new_n24956_), .A2(new_n24974_), .ZN(new_n24977_));
  NAND2_X1   g24680(.A1(new_n24977_), .A2(new_n24953_), .ZN(new_n24978_));
  NAND2_X1   g24681(.A1(new_n24978_), .A2(new_n24976_), .ZN(new_n24979_));
  OAI21_X1   g24682(.A1(new_n24895_), .A2(new_n24927_), .B(new_n24929_), .ZN(new_n24980_));
  NAND2_X1   g24683(.A1(new_n24979_), .A2(new_n24980_), .ZN(new_n24981_));
  XOR2_X1    g24684(.A1(new_n24949_), .A2(new_n24981_), .Z(new_n24982_));
  XOR2_X1    g24685(.A1(new_n24982_), .A2(new_n24942_), .Z(\f[121] ));
  INV_X1     g24686(.I(new_n24979_), .ZN(new_n24984_));
  NOR2_X1    g24687(.A1(new_n24942_), .A2(new_n24984_), .ZN(new_n24985_));
  NAND2_X1   g24688(.A1(new_n24942_), .A2(new_n24984_), .ZN(new_n24986_));
  AND2_X2    g24689(.A1(new_n24986_), .A2(new_n24980_), .Z(new_n24987_));
  AOI21_X1   g24690(.A1(new_n24949_), .A2(new_n24987_), .B(new_n24985_), .ZN(new_n24988_));
  NOR2_X1    g24691(.A1(new_n24973_), .A2(new_n24953_), .ZN(new_n24989_));
  NOR2_X1    g24692(.A1(new_n24989_), .A2(new_n24975_), .ZN(new_n24990_));
  OAI21_X1   g24693(.A1(new_n12643_), .A2(new_n12637_), .B(new_n16487_), .ZN(new_n24991_));
  OAI21_X1   g24694(.A1(new_n24959_), .A2(new_n24969_), .B(new_n24970_), .ZN(new_n24992_));
  NOR2_X1    g24695(.A1(new_n13476_), .A2(new_n12542_), .ZN(new_n24993_));
  XOR2_X1    g24696(.A1(new_n14736_), .A2(new_n12542_), .Z(new_n24994_));
  NAND2_X1   g24697(.A1(new_n24994_), .A2(\b[59] ), .ZN(new_n24995_));
  XOR2_X1    g24698(.A1(new_n24995_), .A2(new_n24993_), .Z(new_n24996_));
  NOR2_X1    g24699(.A1(new_n24966_), .A2(new_n24996_), .ZN(new_n24997_));
  INV_X1     g24700(.I(new_n24996_), .ZN(new_n24998_));
  NOR2_X1    g24701(.A1(new_n24998_), .A2(new_n24965_), .ZN(new_n24999_));
  OAI21_X1   g24702(.A1(new_n24997_), .A2(new_n24999_), .B(new_n24992_), .ZN(new_n25000_));
  INV_X1     g24703(.I(new_n24992_), .ZN(new_n25001_));
  XNOR2_X1   g24704(.A1(new_n24965_), .A2(new_n24996_), .ZN(new_n25002_));
  NAND2_X1   g24705(.A1(new_n25001_), .A2(new_n25002_), .ZN(new_n25003_));
  NAND2_X1   g24706(.A1(new_n25003_), .A2(new_n25000_), .ZN(new_n25004_));
  OAI22_X1   g24707(.A1(new_n13880_), .A2(new_n14209_), .B1(new_n13367_), .B2(new_n13885_), .ZN(new_n25005_));
  AOI21_X1   g24708(.A1(new_n25005_), .A2(new_n13476_), .B(new_n13879_), .ZN(new_n25006_));
  XOR2_X1    g24709(.A1(new_n14213_), .A2(new_n25006_), .Z(new_n25007_));
  XOR2_X1    g24710(.A1(new_n25004_), .A2(new_n25007_), .Z(new_n25008_));
  XOR2_X1    g24711(.A1(new_n25008_), .A2(new_n24991_), .Z(new_n25009_));
  XOR2_X1    g24712(.A1(new_n25009_), .A2(\a[59] ), .Z(new_n25010_));
  NOR2_X1    g24713(.A1(new_n25010_), .A2(new_n24990_), .ZN(new_n25011_));
  NAND2_X1   g24714(.A1(new_n25010_), .A2(new_n24990_), .ZN(new_n25012_));
  INV_X1     g24715(.I(new_n25012_), .ZN(new_n25013_));
  NOR2_X1    g24716(.A1(new_n25013_), .A2(new_n25011_), .ZN(new_n25014_));
  XOR2_X1    g24717(.A1(new_n24988_), .A2(new_n25014_), .Z(\f[122] ));
  INV_X1     g24718(.I(new_n25004_), .ZN(new_n25016_));
  NOR2_X1    g24719(.A1(new_n25016_), .A2(new_n25007_), .ZN(new_n25017_));
  NAND2_X1   g24720(.A1(new_n25016_), .A2(new_n25007_), .ZN(new_n25018_));
  XOR2_X1    g24721(.A1(new_n24991_), .A2(\a[59] ), .Z(new_n25019_));
  AOI21_X1   g24722(.A1(new_n25019_), .A2(new_n25018_), .B(new_n25017_), .ZN(new_n25020_));
  NOR2_X1    g24723(.A1(new_n25001_), .A2(new_n24997_), .ZN(new_n25021_));
  NOR2_X1    g24724(.A1(new_n25021_), .A2(new_n24999_), .ZN(new_n25022_));
  AOI22_X1   g24725(.A1(new_n13472_), .A2(new_n16148_), .B1(\b[61] ), .B2(new_n13884_), .ZN(new_n25023_));
  OAI21_X1   g24726(.A1(new_n25023_), .A2(\a[62] ), .B(new_n13466_), .ZN(new_n25024_));
  XOR2_X1    g24727(.A1(new_n14599_), .A2(new_n25024_), .Z(new_n25025_));
  NOR2_X1    g24728(.A1(new_n13476_), .A2(new_n12970_), .ZN(new_n25026_));
  XOR2_X1    g24729(.A1(new_n14736_), .A2(new_n12970_), .Z(new_n25027_));
  NAND2_X1   g24730(.A1(new_n25027_), .A2(\b[60] ), .ZN(new_n25028_));
  XOR2_X1    g24731(.A1(new_n25028_), .A2(new_n25026_), .Z(new_n25029_));
  XOR2_X1    g24732(.A1(new_n25029_), .A2(\a[59] ), .Z(new_n25030_));
  NOR2_X1    g24733(.A1(new_n25030_), .A2(new_n24996_), .ZN(new_n25031_));
  NOR2_X1    g24734(.A1(new_n25029_), .A2(new_n12222_), .ZN(new_n25032_));
  INV_X1     g24735(.I(new_n25032_), .ZN(new_n25033_));
  NAND2_X1   g24736(.A1(new_n25029_), .A2(new_n12222_), .ZN(new_n25034_));
  AOI21_X1   g24737(.A1(new_n25033_), .A2(new_n25034_), .B(new_n24998_), .ZN(new_n25035_));
  NOR2_X1    g24738(.A1(new_n25031_), .A2(new_n25035_), .ZN(new_n25036_));
  XOR2_X1    g24739(.A1(new_n25025_), .A2(new_n25036_), .Z(new_n25037_));
  INV_X1     g24740(.I(new_n25036_), .ZN(new_n25038_));
  AND2_X2    g24741(.A1(new_n25025_), .A2(new_n25038_), .Z(new_n25039_));
  NOR2_X1    g24742(.A1(new_n25025_), .A2(new_n25038_), .ZN(new_n25040_));
  OAI21_X1   g24743(.A1(new_n25039_), .A2(new_n25040_), .B(new_n25022_), .ZN(new_n25041_));
  OAI21_X1   g24744(.A1(new_n25022_), .A2(new_n25037_), .B(new_n25041_), .ZN(new_n25042_));
  NAND2_X1   g24745(.A1(new_n25042_), .A2(new_n25020_), .ZN(new_n25043_));
  INV_X1     g24746(.I(new_n25043_), .ZN(new_n25044_));
  NOR2_X1    g24747(.A1(new_n25042_), .A2(new_n25020_), .ZN(new_n25045_));
  NOR2_X1    g24748(.A1(new_n25044_), .A2(new_n25045_), .ZN(new_n25046_));
  AOI21_X1   g24749(.A1(new_n25012_), .A2(new_n25046_), .B(new_n25014_), .ZN(new_n25047_));
  XNOR2_X1   g24750(.A1(new_n24988_), .A2(new_n25047_), .ZN(\f[123] ));
  OAI21_X1   g24751(.A1(new_n24848_), .A2(new_n24844_), .B(new_n24947_), .ZN(new_n25049_));
  INV_X1     g24752(.I(new_n24985_), .ZN(new_n25050_));
  INV_X1     g24753(.I(new_n24987_), .ZN(new_n25051_));
  OAI21_X1   g24754(.A1(new_n25049_), .A2(new_n25051_), .B(new_n25050_), .ZN(new_n25052_));
  NOR2_X1    g24755(.A1(new_n25013_), .A2(new_n25011_), .ZN(new_n25053_));
  INV_X1     g24756(.I(new_n25053_), .ZN(new_n25054_));
  INV_X1     g24757(.I(new_n25040_), .ZN(new_n25055_));
  OAI21_X1   g24758(.A1(new_n25022_), .A2(new_n25039_), .B(new_n25055_), .ZN(new_n25056_));
  NAND2_X1   g24759(.A1(new_n13884_), .A2(new_n13469_), .ZN(new_n25057_));
  NOR2_X1    g24760(.A1(new_n14596_), .A2(\a[62] ), .ZN(new_n25058_));
  AOI21_X1   g24761(.A1(new_n25057_), .A2(new_n25058_), .B(new_n13879_), .ZN(new_n25059_));
  XOR2_X1    g24762(.A1(new_n14978_), .A2(new_n25059_), .Z(new_n25060_));
  NAND2_X1   g24763(.A1(new_n25034_), .A2(new_n24998_), .ZN(new_n25061_));
  NAND2_X1   g24764(.A1(new_n25061_), .A2(new_n25033_), .ZN(new_n25062_));
  NOR2_X1    g24765(.A1(new_n13476_), .A2(new_n13367_), .ZN(new_n25063_));
  XOR2_X1    g24766(.A1(new_n14736_), .A2(new_n13367_), .Z(new_n25064_));
  NAND2_X1   g24767(.A1(new_n25064_), .A2(\b[61] ), .ZN(new_n25065_));
  XOR2_X1    g24768(.A1(new_n25065_), .A2(new_n25063_), .Z(new_n25066_));
  INV_X1     g24769(.I(new_n25066_), .ZN(new_n25067_));
  XOR2_X1    g24770(.A1(new_n25062_), .A2(new_n25067_), .Z(new_n25068_));
  NOR2_X1    g24771(.A1(new_n25062_), .A2(new_n25066_), .ZN(new_n25069_));
  NAND2_X1   g24772(.A1(new_n25062_), .A2(new_n25066_), .ZN(new_n25070_));
  INV_X1     g24773(.I(new_n25070_), .ZN(new_n25071_));
  OAI21_X1   g24774(.A1(new_n25069_), .A2(new_n25071_), .B(new_n25060_), .ZN(new_n25072_));
  OAI21_X1   g24775(.A1(new_n25060_), .A2(new_n25068_), .B(new_n25072_), .ZN(new_n25073_));
  NAND2_X1   g24776(.A1(new_n25056_), .A2(new_n25073_), .ZN(new_n25074_));
  AOI21_X1   g24777(.A1(new_n25052_), .A2(new_n25054_), .B(new_n25074_), .ZN(new_n25075_));
  INV_X1     g24778(.I(new_n25074_), .ZN(new_n25076_));
  NOR3_X1    g24779(.A1(new_n24988_), .A2(new_n25053_), .A3(new_n25076_), .ZN(new_n25077_));
  OAI21_X1   g24780(.A1(new_n25075_), .A2(new_n25077_), .B(new_n25043_), .ZN(new_n25078_));
  OR3_X2     g24781(.A1(new_n25075_), .A2(new_n25043_), .A3(new_n25077_), .Z(new_n25079_));
  NAND2_X1   g24782(.A1(new_n25079_), .A2(new_n25078_), .ZN(\f[124] ));
  OAI21_X1   g24783(.A1(new_n25056_), .A2(new_n25073_), .B(new_n25044_), .ZN(new_n25081_));
  NOR3_X1    g24784(.A1(new_n24988_), .A2(new_n25053_), .A3(new_n25081_), .ZN(new_n25082_));
  OAI21_X1   g24785(.A1(new_n25060_), .A2(new_n25069_), .B(new_n25070_), .ZN(new_n25083_));
  AOI21_X1   g24786(.A1(new_n13466_), .A2(new_n13884_), .B(new_n16486_), .ZN(new_n25084_));
  NOR2_X1    g24787(.A1(new_n13476_), .A2(new_n13785_), .ZN(new_n25085_));
  XOR2_X1    g24788(.A1(new_n14736_), .A2(new_n13785_), .Z(new_n25086_));
  NAND2_X1   g24789(.A1(new_n25086_), .A2(\b[62] ), .ZN(new_n25087_));
  XOR2_X1    g24790(.A1(new_n25087_), .A2(new_n25085_), .Z(new_n25088_));
  INV_X1     g24791(.I(new_n25088_), .ZN(new_n25089_));
  XOR2_X1    g24792(.A1(new_n25084_), .A2(new_n25089_), .Z(new_n25090_));
  XOR2_X1    g24793(.A1(new_n25090_), .A2(new_n25067_), .Z(new_n25091_));
  XOR2_X1    g24794(.A1(new_n25091_), .A2(\a[62] ), .Z(new_n25092_));
  XOR2_X1    g24795(.A1(new_n25092_), .A2(new_n25083_), .Z(new_n25093_));
  OAI21_X1   g24796(.A1(new_n25082_), .A2(new_n25076_), .B(new_n25093_), .ZN(new_n25094_));
  INV_X1     g24797(.I(new_n25081_), .ZN(new_n25095_));
  NAND3_X1   g24798(.A1(new_n25052_), .A2(new_n25054_), .A3(new_n25095_), .ZN(new_n25096_));
  NOR2_X1    g24799(.A1(new_n25092_), .A2(new_n25083_), .ZN(new_n25097_));
  INV_X1     g24800(.I(new_n25097_), .ZN(new_n25098_));
  NAND2_X1   g24801(.A1(new_n25092_), .A2(new_n25083_), .ZN(new_n25099_));
  NAND2_X1   g24802(.A1(new_n25098_), .A2(new_n25099_), .ZN(new_n25100_));
  NAND3_X1   g24803(.A1(new_n25096_), .A2(new_n25074_), .A3(new_n25100_), .ZN(new_n25101_));
  NAND2_X1   g24804(.A1(new_n25101_), .A2(new_n25094_), .ZN(\f[125] ));
  INV_X1     g24805(.I(new_n25099_), .ZN(new_n25103_));
  AOI21_X1   g24806(.A1(new_n25096_), .A2(new_n25074_), .B(new_n25097_), .ZN(new_n25104_));
  AND2_X2    g24807(.A1(new_n25084_), .A2(\a[62] ), .Z(new_n25105_));
  NOR2_X1    g24808(.A1(new_n25084_), .A2(\a[62] ), .ZN(new_n25106_));
  OAI22_X1   g24809(.A1(new_n25105_), .A2(new_n25106_), .B1(new_n25067_), .B2(new_n25089_), .ZN(new_n25107_));
  OAI21_X1   g24810(.A1(new_n25066_), .A2(new_n25088_), .B(new_n25107_), .ZN(new_n25108_));
  NOR2_X1    g24811(.A1(new_n13476_), .A2(new_n14208_), .ZN(new_n25109_));
  XOR2_X1    g24812(.A1(new_n14736_), .A2(new_n14208_), .Z(new_n25110_));
  NAND2_X1   g24813(.A1(new_n25110_), .A2(\b[63] ), .ZN(new_n25111_));
  XOR2_X1    g24814(.A1(new_n25111_), .A2(new_n25109_), .Z(new_n25112_));
  XOR2_X1    g24815(.A1(new_n25112_), .A2(\a[62] ), .Z(new_n25113_));
  NOR2_X1    g24816(.A1(new_n25113_), .A2(new_n25066_), .ZN(new_n25114_));
  NOR2_X1    g24817(.A1(new_n25112_), .A2(new_n13476_), .ZN(new_n25115_));
  INV_X1     g24818(.I(new_n25115_), .ZN(new_n25116_));
  NAND2_X1   g24819(.A1(new_n25112_), .A2(new_n13476_), .ZN(new_n25117_));
  AOI21_X1   g24820(.A1(new_n25116_), .A2(new_n25117_), .B(new_n25067_), .ZN(new_n25118_));
  NOR2_X1    g24821(.A1(new_n25114_), .A2(new_n25118_), .ZN(new_n25119_));
  XOR2_X1    g24822(.A1(new_n25108_), .A2(new_n25119_), .Z(new_n25120_));
  OAI21_X1   g24823(.A1(new_n25104_), .A2(new_n25103_), .B(new_n25120_), .ZN(new_n25121_));
  OAI21_X1   g24824(.A1(new_n25082_), .A2(new_n25076_), .B(new_n25098_), .ZN(new_n25122_));
  XNOR2_X1   g24825(.A1(new_n25108_), .A2(new_n25119_), .ZN(new_n25123_));
  NAND3_X1   g24826(.A1(new_n25122_), .A2(new_n25099_), .A3(new_n25123_), .ZN(new_n25124_));
  NAND2_X1   g24827(.A1(new_n25121_), .A2(new_n25124_), .ZN(\f[126] ));
  OAI21_X1   g24828(.A1(new_n25114_), .A2(new_n25118_), .B(new_n25108_), .ZN(new_n25126_));
  NOR3_X1    g24829(.A1(new_n25113_), .A2(new_n14592_), .A3(new_n14736_), .ZN(new_n25127_));
  XOR2_X1    g24830(.A1(new_n25127_), .A2(new_n25116_), .Z(new_n25128_));
  XOR2_X1    g24831(.A1(new_n25128_), .A2(new_n25066_), .Z(new_n25129_));
  NAND2_X1   g24832(.A1(new_n25123_), .A2(new_n25129_), .ZN(new_n25130_));
  XNOR2_X1   g24833(.A1(new_n25130_), .A2(new_n25126_), .ZN(new_n25131_));
  INV_X1     g24834(.I(new_n25131_), .ZN(new_n25132_));
  NAND3_X1   g24835(.A1(new_n25122_), .A2(new_n25099_), .A3(new_n25132_), .ZN(new_n25133_));
  OAI21_X1   g24836(.A1(new_n25104_), .A2(new_n25103_), .B(new_n25131_), .ZN(new_n25134_));
  NAND2_X1   g24837(.A1(new_n25134_), .A2(new_n25133_), .ZN(\f[127] ));
endmodule


