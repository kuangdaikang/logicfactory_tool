// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:57 2022

module ti  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43,
    v44, v45, v46,
    \v47.0 , \v47.1 , \v47.2 , \v47.3 , \v47.4 , \v47.5 , \v47.6 , \v47.7 ,
    \v47.8 , \v47.9 , \v47.10 , \v47.11 , \v47.12 , \v47.13 , \v47.14 ,
    \v47.15 , \v47.16 , \v47.17 , \v47.18 , \v47.19 , \v47.20 , \v47.21 ,
    \v47.22 , \v47.23 , \v47.24 , \v47.25 , \v47.26 , \v47.27 , \v47.28 ,
    \v47.29 , \v47.30 , \v47.31 , \v47.32 , \v47.33 , \v47.34 , \v47.35 ,
    \v47.36 , \v47.37 , \v47.38 , \v47.39 , \v47.40 , \v47.41 , \v47.42 ,
    \v47.43 , \v47.44 , \v47.45 , \v47.46 , \v47.47 , \v47.48 , \v47.49 ,
    \v47.50 , \v47.51 , \v47.52 , \v47.53 , \v47.54 , \v47.55 , \v47.56 ,
    \v47.57 , \v47.58 , \v47.59 , \v47.60 , \v47.61 , \v47.62 , \v47.63 ,
    \v47.64 , \v47.65 , \v47.66 , \v47.67 , \v47.68 , \v47.69 , \v47.70 ,
    \v47.71   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42,
    v43, v44, v45, v46;
  output \v47.0 , \v47.1 , \v47.2 , \v47.3 , \v47.4 , \v47.5 , \v47.6 ,
    \v47.7 , \v47.8 , \v47.9 , \v47.10 , \v47.11 , \v47.12 , \v47.13 ,
    \v47.14 , \v47.15 , \v47.16 , \v47.17 , \v47.18 , \v47.19 , \v47.20 ,
    \v47.21 , \v47.22 , \v47.23 , \v47.24 , \v47.25 , \v47.26 , \v47.27 ,
    \v47.28 , \v47.29 , \v47.30 , \v47.31 , \v47.32 , \v47.33 , \v47.34 ,
    \v47.35 , \v47.36 , \v47.37 , \v47.38 , \v47.39 , \v47.40 , \v47.41 ,
    \v47.42 , \v47.43 , \v47.44 , \v47.45 , \v47.46 , \v47.47 , \v47.48 ,
    \v47.49 , \v47.50 , \v47.51 , \v47.52 , \v47.53 , \v47.54 , \v47.55 ,
    \v47.56 , \v47.57 , \v47.58 , \v47.59 , \v47.60 , \v47.61 , \v47.62 ,
    \v47.63 , \v47.64 , \v47.65 , \v47.66 , \v47.67 , \v47.68 , \v47.69 ,
    \v47.70 , \v47.71 ;
  wire new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1158_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_;
  assign new_n121_ = v21 & v22;
  assign new_n122_ = v11 & ~v22;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = ~v5 & ~v6;
  assign new_n125_ = ~v3 & ~v41;
  assign new_n126_ = v1 & new_n125_;
  assign new_n127_ = ~new_n124_ & ~new_n126_;
  assign new_n128_ = ~v3 & new_n127_;
  assign new_n129_ = ~new_n123_ & ~new_n128_;
  assign new_n130_ = ~v46 & new_n129_;
  assign new_n131_ = v20 & new_n121_;
  assign new_n132_ = v20 & ~new_n131_;
  assign new_n133_ = v18 & v19;
  assign new_n134_ = v39 & v40;
  assign new_n135_ = ~new_n133_ & ~new_n134_;
  assign new_n136_ = ~new_n132_ & ~new_n135_;
  assign new_n137_ = v46 & new_n136_;
  assign new_n138_ = ~new_n130_ & ~new_n137_;
  assign new_n139_ = v43 & ~new_n138_;
  assign new_n140_ = v19 & ~v40;
  assign new_n141_ = ~v40 & ~new_n140_;
  assign new_n142_ = v46 & ~new_n141_;
  assign new_n143_ = ~v43 & new_n142_;
  assign new_n144_ = ~v39 & new_n143_;
  assign new_n145_ = v13 & new_n144_;
  assign new_n146_ = v11 & new_n145_;
  assign new_n147_ = ~new_n139_ & ~new_n146_;
  assign new_n148_ = v42 & ~new_n147_;
  assign new_n149_ = ~new_n121_ & ~new_n133_;
  assign new_n150_ = v19 & ~new_n121_;
  assign new_n151_ = v18 & new_n150_;
  assign new_n152_ = ~new_n149_ & ~new_n151_;
  assign new_n153_ = ~v43 & ~new_n152_;
  assign new_n154_ = ~v43 & ~new_n153_;
  assign new_n155_ = v46 & ~new_n154_;
  assign new_n156_ = ~v42 & new_n155_;
  assign new_n157_ = ~new_n148_ & ~new_n156_;
  assign new_n158_ = ~v45 & ~new_n157_;
  assign new_n159_ = v45 & ~v46;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~v44 & ~new_n160_;
  assign new_n162_ = ~v19 & new_n134_;
  assign new_n163_ = ~v19 & ~new_n162_;
  assign new_n164_ = v46 & ~new_n163_;
  assign new_n165_ = v46 & ~new_n164_;
  assign new_n166_ = ~v43 & ~new_n165_;
  assign new_n167_ = ~v42 & new_n164_;
  assign new_n168_ = v42 & ~v46;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = v43 & ~new_n169_;
  assign new_n171_ = ~new_n166_ & ~new_n170_;
  assign new_n172_ = v45 & ~new_n171_;
  assign new_n173_ = ~v45 & ~v46;
  assign new_n174_ = ~v42 & new_n173_;
  assign new_n175_ = ~new_n172_ & ~new_n174_;
  assign new_n176_ = v44 & ~new_n175_;
  assign new_n177_ = ~new_n161_ & ~new_n176_;
  assign new_n178_ = v35 & ~new_n177_;
  assign new_n179_ = ~v42 & v43;
  assign new_n180_ = ~v35 & new_n179_;
  assign new_n181_ = v44 & new_n159_;
  assign new_n182_ = new_n180_ & new_n181_;
  assign \v47.0  = new_n178_ | new_n182_;
  assign new_n184_ = ~v20 & v21;
  assign new_n185_ = v22 & ~v36;
  assign new_n186_ = new_n184_ & new_n185_;
  assign new_n187_ = v22 & ~new_n186_;
  assign new_n188_ = v41 & ~new_n124_;
  assign new_n189_ = v1 & ~new_n188_;
  assign new_n190_ = ~new_n187_ & ~new_n189_;
  assign new_n191_ = ~v3 & new_n190_;
  assign new_n192_ = ~new_n129_ & ~new_n191_;
  assign new_n193_ = ~v46 & ~new_n192_;
  assign new_n194_ = ~v36 & new_n135_;
  assign new_n195_ = ~v20 & new_n194_;
  assign new_n196_ = ~new_n136_ & ~new_n195_;
  assign new_n197_ = v46 & ~new_n196_;
  assign new_n198_ = ~new_n193_ & ~new_n197_;
  assign new_n199_ = v43 & ~new_n198_;
  assign new_n200_ = v11 & v13;
  assign new_n201_ = v13 & ~new_n200_;
  assign new_n202_ = ~new_n141_ & ~new_n201_;
  assign new_n203_ = ~v19 & ~v40;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = v46 & ~new_n204_;
  assign new_n206_ = ~v43 & new_n205_;
  assign new_n207_ = ~v39 & new_n206_;
  assign new_n208_ = ~new_n199_ & ~new_n207_;
  assign new_n209_ = v42 & ~new_n208_;
  assign new_n210_ = ~v20 & ~v36;
  assign new_n211_ = v22 & ~new_n210_;
  assign new_n212_ = ~v43 & ~new_n211_;
  assign new_n213_ = ~v43 & ~new_n212_;
  assign new_n214_ = v46 & ~new_n213_;
  assign new_n215_ = v43 & ~v46;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = ~v42 & ~new_n216_;
  assign new_n218_ = ~new_n209_ & ~new_n217_;
  assign new_n219_ = ~v44 & ~new_n218_;
  assign new_n220_ = v44 & ~v46;
  assign new_n221_ = ~new_n219_ & ~new_n220_;
  assign new_n222_ = ~v45 & ~new_n221_;
  assign new_n223_ = ~v42 & ~v44;
  assign new_n224_ = ~v42 & ~new_n223_;
  assign new_n225_ = ~v46 & ~new_n224_;
  assign new_n226_ = v44 & new_n164_;
  assign new_n227_ = ~v42 & new_n226_;
  assign new_n228_ = ~new_n225_ & ~new_n227_;
  assign new_n229_ = ~v43 & ~new_n228_;
  assign new_n230_ = ~v44 & v46;
  assign new_n231_ = ~new_n220_ & ~new_n230_;
  assign new_n232_ = v43 & ~new_n231_;
  assign new_n233_ = v42 & new_n232_;
  assign new_n234_ = ~new_n229_ & ~new_n233_;
  assign new_n235_ = v45 & ~new_n234_;
  assign new_n236_ = ~new_n222_ & ~new_n235_;
  assign \v47.1  = v35 & ~new_n236_;
  assign new_n238_ = v22 & ~new_n121_;
  assign new_n239_ = ~new_n189_ & ~new_n238_;
  assign new_n240_ = ~v3 & new_n239_;
  assign new_n241_ = ~new_n129_ & ~new_n240_;
  assign new_n242_ = ~v46 & ~new_n241_;
  assign new_n243_ = ~v20 & ~new_n135_;
  assign new_n244_ = ~new_n135_ & ~new_n243_;
  assign new_n245_ = v46 & ~new_n244_;
  assign new_n246_ = ~new_n242_ & ~new_n245_;
  assign new_n247_ = v43 & ~new_n246_;
  assign new_n248_ = ~v13 & ~new_n141_;
  assign new_n249_ = ~new_n203_ & ~new_n248_;
  assign new_n250_ = v46 & ~new_n249_;
  assign new_n251_ = ~v43 & new_n250_;
  assign new_n252_ = ~v39 & new_n251_;
  assign new_n253_ = ~new_n247_ & ~new_n252_;
  assign new_n254_ = v42 & ~new_n253_;
  assign new_n255_ = ~v21 & ~new_n133_;
  assign new_n256_ = ~v13 & v18;
  assign new_n257_ = v19 & ~v22;
  assign new_n258_ = new_n256_ & new_n257_;
  assign new_n259_ = ~new_n131_ & ~new_n258_;
  assign new_n260_ = ~new_n255_ & new_n259_;
  assign new_n261_ = v20 & new_n260_;
  assign new_n262_ = ~v43 & ~new_n261_;
  assign new_n263_ = ~v43 & ~new_n262_;
  assign new_n264_ = v46 & ~new_n263_;
  assign new_n265_ = ~new_n215_ & ~new_n264_;
  assign new_n266_ = ~v42 & ~new_n265_;
  assign new_n267_ = ~new_n254_ & ~new_n266_;
  assign new_n268_ = ~v45 & ~new_n267_;
  assign new_n269_ = ~v19 & new_n179_;
  assign new_n270_ = v43 & ~new_n269_;
  assign new_n271_ = ~v46 & ~new_n270_;
  assign new_n272_ = v43 & v46;
  assign new_n273_ = v42 & new_n272_;
  assign new_n274_ = ~new_n271_ & ~new_n273_;
  assign new_n275_ = v45 & ~new_n274_;
  assign new_n276_ = ~new_n268_ & ~new_n275_;
  assign new_n277_ = ~v44 & ~new_n276_;
  assign new_n278_ = v42 & v45;
  assign new_n279_ = v45 & ~new_n278_;
  assign new_n280_ = v43 & ~new_n279_;
  assign new_n281_ = v42 & ~v43;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = ~v46 & ~new_n282_;
  assign new_n284_ = ~new_n179_ & ~new_n281_;
  assign new_n285_ = ~new_n163_ & ~new_n284_;
  assign new_n286_ = v46 & new_n285_;
  assign new_n287_ = v45 & new_n286_;
  assign new_n288_ = ~new_n283_ & ~new_n287_;
  assign new_n289_ = v44 & ~new_n288_;
  assign new_n290_ = ~new_n277_ & ~new_n289_;
  assign \v47.2  = v35 & ~new_n290_;
  assign new_n292_ = ~v19 & ~v39;
  assign new_n293_ = v40 & v46;
  assign new_n294_ = new_n292_ & new_n293_;
  assign new_n295_ = v46 & ~new_n294_;
  assign new_n296_ = ~v42 & ~new_n295_;
  assign new_n297_ = ~v19 & v40;
  assign new_n298_ = ~v19 & ~new_n297_;
  assign new_n299_ = v46 & ~new_n298_;
  assign new_n300_ = v42 & new_n299_;
  assign new_n301_ = ~new_n296_ & ~new_n300_;
  assign new_n302_ = v45 & ~new_n301_;
  assign new_n303_ = ~new_n174_ & ~new_n302_;
  assign new_n304_ = v44 & ~new_n303_;
  assign new_n305_ = ~new_n140_ & ~new_n297_;
  assign new_n306_ = v13 & ~new_n305_;
  assign new_n307_ = ~v11 & new_n306_;
  assign new_n308_ = ~new_n203_ & ~new_n307_;
  assign new_n309_ = v42 & ~new_n308_;
  assign new_n310_ = ~v39 & new_n309_;
  assign new_n311_ = ~v21 & ~v42;
  assign new_n312_ = new_n133_ & new_n311_;
  assign new_n313_ = ~new_n310_ & ~new_n312_;
  assign new_n314_ = v46 & ~new_n313_;
  assign new_n315_ = ~v45 & new_n314_;
  assign new_n316_ = ~v44 & new_n315_;
  assign new_n317_ = ~new_n304_ & ~new_n316_;
  assign new_n318_ = ~v43 & ~new_n317_;
  assign new_n319_ = ~v4 & new_n124_;
  assign new_n320_ = v3 & v41;
  assign new_n321_ = ~new_n319_ & ~new_n320_;
  assign new_n322_ = ~v46 & ~new_n321_;
  assign new_n323_ = ~v22 & new_n322_;
  assign new_n324_ = ~v11 & new_n323_;
  assign new_n325_ = v46 & ~new_n135_;
  assign new_n326_ = v22 & new_n325_;
  assign new_n327_ = v21 & new_n326_;
  assign new_n328_ = v20 & new_n327_;
  assign new_n329_ = ~new_n324_ & ~new_n328_;
  assign new_n330_ = ~v45 & ~new_n329_;
  assign new_n331_ = ~new_n159_ & ~new_n330_;
  assign new_n332_ = v42 & ~new_n331_;
  assign new_n333_ = v19 & v45;
  assign new_n334_ = v45 & ~new_n333_;
  assign new_n335_ = ~v46 & ~new_n334_;
  assign new_n336_ = ~v42 & new_n335_;
  assign new_n337_ = ~new_n332_ & ~new_n336_;
  assign new_n338_ = ~v44 & ~new_n337_;
  assign new_n339_ = v45 & new_n164_;
  assign new_n340_ = ~v42 & new_n339_;
  assign new_n341_ = v42 & new_n173_;
  assign new_n342_ = ~new_n340_ & ~new_n341_;
  assign new_n343_ = v44 & ~new_n342_;
  assign new_n344_ = ~new_n338_ & ~new_n343_;
  assign new_n345_ = v43 & ~new_n344_;
  assign new_n346_ = ~new_n318_ & ~new_n345_;
  assign \v47.3  = v35 & ~new_n346_;
  assign new_n348_ = ~v44 & v45;
  assign new_n349_ = new_n281_ & new_n348_;
  assign new_n350_ = v12 & ~v42;
  assign new_n351_ = v44 & ~v45;
  assign new_n352_ = v43 & new_n351_;
  assign new_n353_ = new_n350_ & new_n352_;
  assign new_n354_ = ~new_n349_ & ~new_n353_;
  assign new_n355_ = v43 & v45;
  assign new_n356_ = v43 & ~new_n355_;
  assign new_n357_ = v44 & ~new_n356_;
  assign new_n358_ = v4 & ~v11;
  assign new_n359_ = ~v11 & ~new_n358_;
  assign new_n360_ = ~v6 & ~new_n359_;
  assign new_n361_ = ~v5 & new_n360_;
  assign new_n362_ = ~v3 & ~new_n126_;
  assign new_n363_ = v11 & ~new_n362_;
  assign new_n364_ = ~v3 & ~new_n189_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = ~new_n361_ & new_n365_;
  assign new_n367_ = ~v22 & ~new_n366_;
  assign new_n368_ = v11 & ~new_n121_;
  assign new_n369_ = ~v3 & ~new_n368_;
  assign new_n370_ = v1 & new_n369_;
  assign new_n371_ = v3 & ~v11;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign new_n373_ = ~v41 & ~new_n372_;
  assign new_n374_ = ~v3 & ~new_n124_;
  assign new_n375_ = v22 & ~new_n374_;
  assign new_n376_ = v21 & new_n375_;
  assign new_n377_ = ~new_n373_ & ~new_n376_;
  assign new_n378_ = ~new_n367_ & new_n377_;
  assign new_n379_ = ~v45 & ~new_n378_;
  assign new_n380_ = ~v18 & v45;
  assign new_n381_ = ~new_n379_ & ~new_n380_;
  assign new_n382_ = ~v44 & ~new_n381_;
  assign new_n383_ = v43 & new_n382_;
  assign new_n384_ = ~new_n357_ & ~new_n383_;
  assign new_n385_ = v42 & ~new_n384_;
  assign new_n386_ = ~v12 & v44;
  assign new_n387_ = v44 & ~new_n386_;
  assign new_n388_ = ~v45 & ~new_n387_;
  assign new_n389_ = v43 & new_n388_;
  assign new_n390_ = ~v43 & new_n348_;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = ~v42 & ~new_n391_;
  assign new_n393_ = ~new_n385_ & ~new_n392_;
  assign new_n394_ = new_n354_ & new_n393_;
  assign new_n395_ = ~v46 & ~new_n394_;
  assign new_n396_ = ~new_n202_ & ~new_n307_;
  assign new_n397_ = v42 & ~new_n396_;
  assign new_n398_ = ~v39 & new_n397_;
  assign new_n399_ = v13 & v18;
  assign new_n400_ = new_n257_ & new_n399_;
  assign new_n401_ = ~new_n255_ & ~new_n400_;
  assign new_n402_ = ~v42 & ~new_n401_;
  assign new_n403_ = ~new_n398_ & ~new_n402_;
  assign new_n404_ = ~v45 & ~new_n403_;
  assign new_n405_ = ~v44 & new_n404_;
  assign new_n406_ = v40 & ~v42;
  assign new_n407_ = new_n292_ & new_n406_;
  assign new_n408_ = new_n163_ & ~new_n407_;
  assign new_n409_ = v45 & ~new_n408_;
  assign new_n410_ = v44 & new_n409_;
  assign new_n411_ = ~new_n405_ & ~new_n410_;
  assign new_n412_ = ~v43 & ~new_n411_;
  assign new_n413_ = ~v45 & ~new_n135_;
  assign new_n414_ = ~v44 & new_n413_;
  assign new_n415_ = v42 & new_n414_;
  assign new_n416_ = v22 & new_n415_;
  assign new_n417_ = v21 & new_n416_;
  assign new_n418_ = v20 & new_n417_;
  assign new_n419_ = ~v39 & v40;
  assign new_n420_ = ~v19 & new_n419_;
  assign new_n421_ = v44 & v45;
  assign new_n422_ = ~v42 & new_n421_;
  assign new_n423_ = new_n420_ & new_n422_;
  assign new_n424_ = ~new_n418_ & ~new_n423_;
  assign new_n425_ = v43 & ~new_n424_;
  assign new_n426_ = ~new_n412_ & ~new_n425_;
  assign new_n427_ = v46 & ~new_n426_;
  assign new_n428_ = ~new_n395_ & ~new_n427_;
  assign \v47.4  = v35 & ~new_n428_;
  assign new_n430_ = v8 & ~v33;
  assign new_n431_ = v7 & new_n430_;
  assign new_n432_ = v8 & ~new_n431_;
  assign new_n433_ = v6 & ~new_n432_;
  assign new_n434_ = ~v7 & ~v8;
  assign new_n435_ = v8 & ~v32;
  assign new_n436_ = v7 & new_n435_;
  assign new_n437_ = ~new_n434_ & ~new_n436_;
  assign new_n438_ = ~v6 & ~new_n437_;
  assign new_n439_ = ~new_n433_ & ~new_n438_;
  assign new_n440_ = ~v30 & ~new_n439_;
  assign new_n441_ = ~v8 & ~v32;
  assign new_n442_ = ~v6 & new_n441_;
  assign new_n443_ = v6 & ~v33;
  assign new_n444_ = ~new_n442_ & ~new_n443_;
  assign new_n445_ = ~v7 & ~new_n444_;
  assign new_n446_ = ~new_n440_ & ~new_n445_;
  assign new_n447_ = v4 & ~new_n446_;
  assign new_n448_ = v8 & ~new_n436_;
  assign new_n449_ = v6 & ~new_n448_;
  assign new_n450_ = ~new_n431_ & ~new_n434_;
  assign new_n451_ = ~v6 & ~new_n450_;
  assign new_n452_ = ~new_n449_ & ~new_n451_;
  assign new_n453_ = ~v29 & ~new_n452_;
  assign new_n454_ = v6 & ~v32;
  assign new_n455_ = ~v8 & ~v33;
  assign new_n456_ = ~v6 & new_n455_;
  assign new_n457_ = ~new_n454_ & ~new_n456_;
  assign new_n458_ = ~v7 & ~new_n457_;
  assign new_n459_ = ~new_n453_ & ~new_n458_;
  assign new_n460_ = ~v4 & ~new_n459_;
  assign new_n461_ = ~new_n447_ & ~new_n460_;
  assign new_n462_ = v5 & ~new_n461_;
  assign new_n463_ = v7 & v8;
  assign new_n464_ = ~v32 & ~v33;
  assign new_n465_ = new_n463_ & new_n464_;
  assign new_n466_ = v8 & ~new_n465_;
  assign new_n467_ = ~v30 & ~new_n466_;
  assign new_n468_ = v4 & new_n467_;
  assign new_n469_ = v32 & v33;
  assign new_n470_ = v8 & ~new_n469_;
  assign new_n471_ = v7 & new_n470_;
  assign new_n472_ = v8 & ~new_n471_;
  assign new_n473_ = ~v4 & ~new_n472_;
  assign new_n474_ = ~new_n468_ & ~new_n473_;
  assign new_n475_ = ~v29 & ~new_n474_;
  assign new_n476_ = v8 & ~v30;
  assign new_n477_ = v7 & new_n476_;
  assign new_n478_ = v7 & ~new_n477_;
  assign new_n479_ = ~new_n469_ & ~new_n478_;
  assign new_n480_ = ~v8 & ~v30;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = ~v4 & ~new_n481_;
  assign new_n483_ = v4 & ~v7;
  assign new_n484_ = new_n464_ & new_n483_;
  assign new_n485_ = ~new_n482_ & ~new_n484_;
  assign new_n486_ = ~new_n475_ & new_n485_;
  assign new_n487_ = v6 & ~new_n486_;
  assign new_n488_ = ~v5 & new_n487_;
  assign new_n489_ = ~new_n462_ & ~new_n488_;
  assign new_n490_ = v46 & ~new_n489_;
  assign new_n491_ = ~v45 & new_n490_;
  assign new_n492_ = ~v44 & new_n491_;
  assign \v47.5  = v35 & new_n492_;
  assign new_n494_ = v41 & new_n374_;
  assign new_n495_ = ~new_n123_ & ~new_n494_;
  assign new_n496_ = ~v22 & v41;
  assign new_n497_ = v41 & ~new_n496_;
  assign new_n498_ = v3 & ~new_n497_;
  assign new_n499_ = ~v18 & v19;
  assign new_n500_ = v19 & ~new_n499_;
  assign new_n501_ = ~new_n124_ & new_n500_;
  assign new_n502_ = ~v22 & ~new_n501_;
  assign new_n503_ = ~new_n126_ & ~new_n502_;
  assign new_n504_ = ~new_n498_ & new_n503_;
  assign new_n505_ = ~v11 & ~new_n504_;
  assign new_n506_ = v7 & ~v8;
  assign new_n507_ = ~v4 & ~v6;
  assign new_n508_ = ~v4 & ~new_n507_;
  assign new_n509_ = ~new_n506_ & ~new_n508_;
  assign new_n510_ = ~v7 & v8;
  assign new_n511_ = v41 & ~new_n238_;
  assign new_n512_ = ~v3 & new_n511_;
  assign new_n513_ = new_n510_ & ~new_n512_;
  assign new_n514_ = ~new_n509_ & new_n513_;
  assign new_n515_ = v5 & ~new_n514_;
  assign new_n516_ = v4 & v5;
  assign new_n517_ = ~new_n506_ & ~new_n516_;
  assign new_n518_ = ~v5 & ~new_n510_;
  assign new_n519_ = ~new_n512_ & ~new_n518_;
  assign new_n520_ = ~new_n517_ & new_n519_;
  assign new_n521_ = v6 & ~new_n520_;
  assign new_n522_ = ~v3 & ~new_n238_;
  assign new_n523_ = ~v1 & new_n522_;
  assign new_n524_ = ~new_n521_ & ~new_n523_;
  assign new_n525_ = ~new_n515_ & new_n524_;
  assign new_n526_ = ~new_n505_ & new_n525_;
  assign new_n527_ = ~new_n495_ & new_n526_;
  assign new_n528_ = ~v46 & ~new_n527_;
  assign new_n529_ = v18 & new_n203_;
  assign new_n530_ = ~v40 & ~new_n529_;
  assign new_n531_ = v46 & ~new_n530_;
  assign new_n532_ = ~v39 & new_n531_;
  assign new_n533_ = ~new_n528_ & ~new_n532_;
  assign new_n534_ = v43 & ~new_n533_;
  assign new_n535_ = v42 & new_n534_;
  assign new_n536_ = ~v22 & ~new_n133_;
  assign new_n537_ = ~new_n121_ & ~new_n536_;
  assign new_n538_ = v46 & ~new_n537_;
  assign new_n539_ = ~v43 & new_n538_;
  assign new_n540_ = ~v42 & new_n539_;
  assign new_n541_ = ~new_n535_ & ~new_n540_;
  assign new_n542_ = ~v45 & ~new_n541_;
  assign new_n543_ = ~v40 & v42;
  assign new_n544_ = v45 & v46;
  assign new_n545_ = v43 & new_n544_;
  assign new_n546_ = new_n543_ & new_n545_;
  assign new_n547_ = ~new_n542_ & ~new_n546_;
  assign new_n548_ = ~v44 & ~new_n547_;
  assign new_n549_ = v42 & v43;
  assign new_n550_ = v44 & new_n173_;
  assign new_n551_ = new_n549_ & new_n550_;
  assign new_n552_ = ~new_n548_ & ~new_n551_;
  assign \v47.6  = v35 & ~new_n552_;
  assign new_n554_ = ~v18 & ~v19;
  assign new_n555_ = ~v40 & v46;
  assign new_n556_ = ~v39 & new_n555_;
  assign new_n557_ = new_n554_ & new_n556_;
  assign new_n558_ = ~new_n528_ & ~new_n557_;
  assign new_n559_ = v43 & ~new_n558_;
  assign new_n560_ = ~v43 & v46;
  assign new_n561_ = ~new_n559_ & ~new_n560_;
  assign new_n562_ = v42 & ~new_n561_;
  assign new_n563_ = ~new_n540_ & ~new_n562_;
  assign new_n564_ = ~v45 & ~new_n563_;
  assign new_n565_ = ~v39 & v42;
  assign new_n566_ = new_n545_ & new_n565_;
  assign new_n567_ = ~new_n564_ & ~new_n566_;
  assign new_n568_ = ~v44 & ~new_n567_;
  assign new_n569_ = ~new_n551_ & ~new_n568_;
  assign \v47.7  = v35 & ~new_n569_;
  assign new_n571_ = v13 & ~v39;
  assign new_n572_ = ~v40 & new_n560_;
  assign new_n573_ = new_n571_ & new_n572_;
  assign new_n574_ = ~v18 & ~v22;
  assign new_n575_ = new_n215_ & new_n574_;
  assign new_n576_ = ~new_n573_ & ~new_n575_;
  assign new_n577_ = v19 & ~new_n576_;
  assign new_n578_ = ~v11 & new_n577_;
  assign new_n579_ = v38 & new_n272_;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = ~v45 & ~new_n580_;
  assign new_n582_ = ~v38 & v43;
  assign new_n583_ = new_n544_ & new_n582_;
  assign new_n584_ = ~new_n581_ & ~new_n583_;
  assign new_n585_ = ~v44 & ~new_n584_;
  assign new_n586_ = v43 & v44;
  assign new_n587_ = new_n173_ & new_n586_;
  assign new_n588_ = ~new_n585_ & ~new_n587_;
  assign new_n589_ = v42 & ~new_n588_;
  assign new_n590_ = v44 & new_n544_;
  assign new_n591_ = new_n420_ & new_n590_;
  assign new_n592_ = ~new_n589_ & ~new_n591_;
  assign \v47.8  = v35 & ~new_n592_;
  assign new_n594_ = v37 & ~v38;
  assign new_n595_ = v37 & ~new_n594_;
  assign new_n596_ = v46 & ~new_n595_;
  assign new_n597_ = v43 & new_n596_;
  assign new_n598_ = ~new_n578_ & ~new_n597_;
  assign new_n599_ = ~v45 & ~new_n598_;
  assign new_n600_ = ~v37 & v43;
  assign new_n601_ = new_n544_ & new_n600_;
  assign new_n602_ = ~new_n599_ & ~new_n601_;
  assign new_n603_ = ~v44 & ~new_n602_;
  assign new_n604_ = ~new_n587_ & ~new_n603_;
  assign new_n605_ = v42 & ~new_n604_;
  assign new_n606_ = ~new_n591_ & ~new_n605_;
  assign \v47.9  = v35 & ~new_n606_;
  assign new_n608_ = v43 & ~v44;
  assign new_n609_ = v43 & ~new_n608_;
  assign new_n610_ = ~v42 & ~new_n609_;
  assign new_n611_ = v42 & new_n608_;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = v45 & ~new_n612_;
  assign new_n614_ = v3 & new_n188_;
  assign new_n615_ = ~new_n319_ & ~new_n614_;
  assign new_n616_ = ~new_n123_ & ~new_n615_;
  assign new_n617_ = ~v22 & ~new_n500_;
  assign new_n618_ = ~v11 & new_n617_;
  assign new_n619_ = v22 & ~new_n189_;
  assign new_n620_ = v21 & new_n619_;
  assign new_n621_ = ~v3 & new_n620_;
  assign new_n622_ = ~new_n618_ & ~new_n621_;
  assign new_n623_ = ~new_n616_ & new_n622_;
  assign new_n624_ = ~v44 & ~new_n623_;
  assign new_n625_ = ~v44 & ~new_n624_;
  assign new_n626_ = v42 & ~new_n625_;
  assign new_n627_ = ~v42 & v44;
  assign new_n628_ = ~v12 & new_n627_;
  assign new_n629_ = ~new_n626_ & ~new_n628_;
  assign new_n630_ = ~v45 & ~new_n629_;
  assign new_n631_ = v43 & new_n630_;
  assign new_n632_ = ~new_n613_ & ~new_n631_;
  assign new_n633_ = ~v46 & ~new_n632_;
  assign new_n634_ = ~v43 & ~new_n308_;
  assign new_n635_ = ~v39 & new_n634_;
  assign new_n636_ = ~v37 & v38;
  assign new_n637_ = ~v37 & ~new_n636_;
  assign new_n638_ = v43 & ~new_n637_;
  assign new_n639_ = ~new_n635_ & ~new_n638_;
  assign new_n640_ = v42 & ~new_n639_;
  assign new_n641_ = ~v10 & ~v22;
  assign new_n642_ = ~new_n121_ & ~new_n641_;
  assign new_n643_ = ~v43 & ~new_n642_;
  assign new_n644_ = ~v42 & new_n643_;
  assign new_n645_ = ~new_n640_ & ~new_n644_;
  assign new_n646_ = ~v45 & ~new_n645_;
  assign new_n647_ = ~v44 & new_n646_;
  assign new_n648_ = v40 & new_n421_;
  assign new_n649_ = new_n292_ & new_n648_;
  assign new_n650_ = ~new_n647_ & ~new_n649_;
  assign new_n651_ = v46 & ~new_n650_;
  assign new_n652_ = ~new_n633_ & ~new_n651_;
  assign \v47.10  = v35 & ~new_n652_;
  assign new_n654_ = v37 & v43;
  assign new_n655_ = ~new_n635_ & ~new_n654_;
  assign new_n656_ = v46 & ~new_n655_;
  assign new_n657_ = ~v46 & ~new_n622_;
  assign new_n658_ = v43 & new_n657_;
  assign new_n659_ = ~new_n656_ & ~new_n658_;
  assign new_n660_ = v42 & ~new_n659_;
  assign new_n661_ = ~v42 & new_n560_;
  assign new_n662_ = new_n121_ & new_n661_;
  assign new_n663_ = ~new_n660_ & ~new_n662_;
  assign new_n664_ = ~v45 & ~new_n663_;
  assign new_n665_ = v43 & new_n159_;
  assign new_n666_ = ~v42 & new_n665_;
  assign new_n667_ = ~new_n664_ & ~new_n666_;
  assign new_n668_ = ~v44 & ~new_n667_;
  assign new_n669_ = v40 & new_n544_;
  assign new_n670_ = new_n292_ & new_n669_;
  assign new_n671_ = new_n173_ & new_n549_;
  assign new_n672_ = ~new_n670_ & ~new_n671_;
  assign new_n673_ = v44 & ~new_n672_;
  assign new_n674_ = ~new_n668_ & ~new_n673_;
  assign \v47.12  = v35 & ~new_n674_;
  assign new_n676_ = ~v11 & ~v18;
  assign new_n677_ = new_n257_ & new_n676_;
  assign new_n678_ = ~new_n621_ & ~new_n677_;
  assign new_n679_ = ~v45 & ~new_n678_;
  assign new_n680_ = ~v45 & ~new_n679_;
  assign new_n681_ = ~v46 & ~new_n680_;
  assign new_n682_ = ~v45 & v46;
  assign new_n683_ = v38 & new_n682_;
  assign new_n684_ = ~new_n681_ & ~new_n683_;
  assign new_n685_ = v43 & ~new_n684_;
  assign new_n686_ = ~v11 & v13;
  assign new_n687_ = v19 & ~v39;
  assign new_n688_ = new_n686_ & new_n687_;
  assign new_n689_ = ~v40 & ~v43;
  assign new_n690_ = new_n682_ & new_n689_;
  assign new_n691_ = new_n688_ & new_n690_;
  assign new_n692_ = ~new_n685_ & ~new_n691_;
  assign new_n693_ = v42 & ~new_n692_;
  assign new_n694_ = v46 & ~new_n642_;
  assign new_n695_ = ~v45 & new_n694_;
  assign new_n696_ = ~v43 & new_n695_;
  assign new_n697_ = ~v42 & new_n696_;
  assign new_n698_ = ~new_n693_ & ~new_n697_;
  assign new_n699_ = ~v44 & ~new_n698_;
  assign new_n700_ = ~new_n673_ & ~new_n699_;
  assign \v47.13  = v35 & ~new_n700_;
  assign new_n702_ = v46 & ~new_n305_;
  assign new_n703_ = ~v43 & new_n702_;
  assign new_n704_ = ~v39 & new_n703_;
  assign new_n705_ = v13 & new_n704_;
  assign new_n706_ = ~v46 & ~new_n500_;
  assign new_n707_ = v43 & new_n706_;
  assign new_n708_ = ~v22 & new_n707_;
  assign new_n709_ = ~new_n705_ & ~new_n708_;
  assign new_n710_ = ~v11 & ~new_n709_;
  assign new_n711_ = v38 & v43;
  assign new_n712_ = ~v37 & new_n711_;
  assign new_n713_ = new_n292_ & new_n689_;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = v46 & ~new_n714_;
  assign new_n716_ = ~v46 & ~new_n189_;
  assign new_n717_ = v43 & new_n716_;
  assign new_n718_ = v22 & new_n717_;
  assign new_n719_ = v21 & new_n718_;
  assign new_n720_ = ~v3 & new_n719_;
  assign new_n721_ = ~new_n715_ & ~new_n720_;
  assign new_n722_ = ~new_n710_ & new_n721_;
  assign new_n723_ = v42 & ~new_n722_;
  assign new_n724_ = ~v43 & new_n694_;
  assign new_n725_ = ~v42 & new_n724_;
  assign new_n726_ = ~new_n723_ & ~new_n725_;
  assign new_n727_ = ~v45 & ~new_n726_;
  assign new_n728_ = ~new_n666_ & ~new_n727_;
  assign new_n729_ = ~v44 & ~new_n728_;
  assign new_n730_ = ~new_n673_ & ~new_n729_;
  assign \v47.14  = v35 & ~new_n730_;
  assign new_n732_ = ~v11 & ~v19;
  assign new_n733_ = v42 & ~v45;
  assign new_n734_ = ~v22 & new_n733_;
  assign new_n735_ = new_n732_ & new_n734_;
  assign new_n736_ = ~v45 & ~new_n735_;
  assign new_n737_ = ~v46 & ~new_n736_;
  assign new_n738_ = ~new_n594_ & ~new_n636_;
  assign new_n739_ = v46 & ~new_n738_;
  assign new_n740_ = ~v45 & new_n739_;
  assign new_n741_ = v42 & new_n740_;
  assign new_n742_ = ~new_n737_ & ~new_n741_;
  assign new_n743_ = v43 & ~new_n742_;
  assign new_n744_ = v13 & v40;
  assign new_n745_ = ~v11 & new_n744_;
  assign new_n746_ = v40 & ~new_n745_;
  assign new_n747_ = v42 & ~new_n746_;
  assign new_n748_ = ~v39 & new_n747_;
  assign new_n749_ = ~v19 & new_n748_;
  assign new_n750_ = ~v22 & ~v42;
  assign new_n751_ = ~v10 & new_n750_;
  assign new_n752_ = ~new_n749_ & ~new_n751_;
  assign new_n753_ = v46 & ~new_n752_;
  assign new_n754_ = ~v45 & new_n753_;
  assign new_n755_ = ~v43 & new_n754_;
  assign new_n756_ = ~new_n743_ & ~new_n755_;
  assign new_n757_ = ~v44 & ~new_n756_;
  assign \v47.15  = v35 & new_n757_;
  assign new_n759_ = ~v45 & ~new_n622_;
  assign new_n760_ = ~v45 & ~new_n759_;
  assign new_n761_ = ~v46 & ~new_n760_;
  assign new_n762_ = new_n594_ & new_n682_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = v43 & ~new_n763_;
  assign new_n765_ = v46 & ~new_n308_;
  assign new_n766_ = ~v45 & new_n765_;
  assign new_n767_ = ~v43 & new_n766_;
  assign new_n768_ = ~v39 & new_n767_;
  assign new_n769_ = ~new_n764_ & ~new_n768_;
  assign new_n770_ = v42 & ~new_n769_;
  assign new_n771_ = ~new_n697_ & ~new_n770_;
  assign new_n772_ = ~v44 & ~new_n771_;
  assign new_n773_ = ~new_n673_ & ~new_n772_;
  assign \v47.16  = v35 & ~new_n773_;
  assign new_n775_ = v46 & ~new_n639_;
  assign new_n776_ = ~new_n658_ & ~new_n775_;
  assign new_n777_ = v42 & ~new_n776_;
  assign new_n778_ = ~new_n725_ & ~new_n777_;
  assign new_n779_ = ~v44 & ~new_n778_;
  assign new_n780_ = new_n220_ & new_n549_;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = ~v45 & ~new_n781_;
  assign new_n783_ = ~new_n591_ & ~new_n782_;
  assign \v47.17  = v35 & ~new_n783_;
  assign new_n785_ = ~v44 & new_n616_;
  assign new_n786_ = v42 & new_n785_;
  assign new_n787_ = ~new_n628_ & ~new_n786_;
  assign new_n788_ = ~v45 & ~new_n787_;
  assign new_n789_ = v43 & new_n788_;
  assign new_n790_ = ~new_n613_ & ~new_n789_;
  assign new_n791_ = ~v46 & ~new_n790_;
  assign \v47.18  = v35 & new_n791_;
  assign new_n793_ = v35 & new_n641_;
  assign new_n794_ = ~v42 & new_n793_;
  assign new_n795_ = ~v43 & new_n794_;
  assign new_n796_ = ~v44 & new_n795_;
  assign new_n797_ = ~v45 & new_n796_;
  assign \v47.19  = v46 & new_n797_;
  assign new_n799_ = v26 & v27;
  assign new_n800_ = v28 & new_n421_;
  assign new_n801_ = new_n799_ & new_n800_;
  assign new_n802_ = v24 & v25;
  assign new_n803_ = v23 & new_n802_;
  assign new_n804_ = ~v44 & ~v45;
  assign new_n805_ = new_n281_ & new_n804_;
  assign new_n806_ = new_n803_ & new_n805_;
  assign new_n807_ = ~new_n801_ & ~new_n806_;
  assign new_n808_ = v46 & ~new_n807_;
  assign \v47.20  = v35 & new_n808_;
  assign new_n810_ = ~v26 & v27;
  assign new_n811_ = new_n800_ & new_n810_;
  assign new_n812_ = ~v23 & new_n802_;
  assign new_n813_ = new_n805_ & new_n812_;
  assign new_n814_ = ~new_n811_ & ~new_n813_;
  assign new_n815_ = v46 & ~new_n814_;
  assign \v47.21  = v35 & new_n815_;
  assign new_n817_ = v26 & ~v27;
  assign new_n818_ = new_n800_ & new_n817_;
  assign new_n819_ = ~v24 & v25;
  assign new_n820_ = v23 & new_n819_;
  assign new_n821_ = new_n805_ & new_n820_;
  assign new_n822_ = ~new_n818_ & ~new_n821_;
  assign new_n823_ = v46 & ~new_n822_;
  assign \v47.22  = v35 & new_n823_;
  assign new_n825_ = ~v26 & ~v27;
  assign new_n826_ = new_n800_ & new_n825_;
  assign new_n827_ = ~v23 & new_n819_;
  assign new_n828_ = new_n805_ & new_n827_;
  assign new_n829_ = ~new_n826_ & ~new_n828_;
  assign new_n830_ = v46 & ~new_n829_;
  assign \v47.23  = v35 & new_n830_;
  assign new_n832_ = v23 & v24;
  assign new_n833_ = v25 & new_n421_;
  assign new_n834_ = new_n832_ & new_n833_;
  assign new_n835_ = v27 & v28;
  assign new_n836_ = v26 & new_n835_;
  assign new_n837_ = new_n805_ & new_n836_;
  assign new_n838_ = ~new_n834_ & ~new_n837_;
  assign new_n839_ = v46 & ~new_n838_;
  assign \v47.24  = v35 & new_n839_;
  assign new_n841_ = ~v23 & v24;
  assign new_n842_ = new_n833_ & new_n841_;
  assign new_n843_ = ~v26 & new_n835_;
  assign new_n844_ = new_n805_ & new_n843_;
  assign new_n845_ = ~new_n842_ & ~new_n844_;
  assign new_n846_ = v46 & ~new_n845_;
  assign \v47.25  = v35 & new_n846_;
  assign new_n848_ = v23 & ~v24;
  assign new_n849_ = new_n833_ & new_n848_;
  assign new_n850_ = ~v27 & v28;
  assign new_n851_ = v26 & new_n850_;
  assign new_n852_ = new_n805_ & new_n851_;
  assign new_n853_ = ~new_n849_ & ~new_n852_;
  assign new_n854_ = v46 & ~new_n853_;
  assign \v47.26  = v35 & new_n854_;
  assign new_n856_ = ~v23 & ~v24;
  assign new_n857_ = new_n833_ & new_n856_;
  assign new_n858_ = ~v26 & new_n850_;
  assign new_n859_ = new_n805_ & new_n858_;
  assign new_n860_ = ~new_n857_ & ~new_n859_;
  assign new_n861_ = v46 & ~new_n860_;
  assign \v47.27  = v35 & new_n861_;
  assign new_n863_ = v4 & new_n124_;
  assign new_n864_ = v41 & ~new_n863_;
  assign new_n865_ = ~new_n123_ & ~new_n864_;
  assign new_n866_ = ~v46 & new_n865_;
  assign new_n867_ = v43 & new_n866_;
  assign new_n868_ = ~v9 & new_n867_;
  assign new_n869_ = ~v28 & new_n560_;
  assign new_n870_ = ~v27 & new_n869_;
  assign new_n871_ = ~new_n868_ & ~new_n870_;
  assign new_n872_ = ~v45 & ~new_n871_;
  assign new_n873_ = ~v9 & ~v43;
  assign new_n874_ = new_n159_ & new_n873_;
  assign new_n875_ = ~new_n872_ & ~new_n874_;
  assign new_n876_ = ~v44 & ~new_n875_;
  assign new_n877_ = ~v43 & new_n181_;
  assign new_n878_ = v17 & new_n877_;
  assign new_n879_ = ~new_n876_ & ~new_n878_;
  assign new_n880_ = v42 & ~new_n879_;
  assign new_n881_ = ~v25 & new_n544_;
  assign new_n882_ = ~v24 & new_n881_;
  assign new_n883_ = ~v9 & new_n350_;
  assign new_n884_ = v43 & new_n173_;
  assign new_n885_ = new_n883_ & new_n884_;
  assign new_n886_ = ~new_n882_ & ~new_n885_;
  assign new_n887_ = v44 & ~new_n886_;
  assign new_n888_ = ~new_n880_ & ~new_n887_;
  assign \v47.28  = v35 & ~new_n888_;
  assign new_n890_ = ~v43 & v44;
  assign new_n891_ = v5 & new_n890_;
  assign new_n892_ = v15 & new_n608_;
  assign new_n893_ = ~new_n891_ & ~new_n892_;
  assign new_n894_ = ~v42 & ~new_n893_;
  assign new_n895_ = v12 & new_n611_;
  assign new_n896_ = ~new_n894_ & ~new_n895_;
  assign new_n897_ = ~v46 & ~new_n896_;
  assign new_n898_ = v44 & v46;
  assign new_n899_ = ~v28 & new_n898_;
  assign new_n900_ = ~v27 & new_n899_;
  assign new_n901_ = ~new_n897_ & ~new_n900_;
  assign new_n902_ = v45 & ~new_n901_;
  assign new_n903_ = ~v44 & new_n682_;
  assign new_n904_ = ~v43 & new_n903_;
  assign new_n905_ = v42 & new_n904_;
  assign new_n906_ = ~v25 & new_n905_;
  assign new_n907_ = ~v24 & new_n906_;
  assign new_n908_ = ~new_n902_ & ~new_n907_;
  assign \v47.29  = v35 & ~new_n908_;
  assign new_n910_ = ~v24 & ~v25;
  assign new_n911_ = v23 & new_n910_;
  assign new_n912_ = ~v43 & new_n682_;
  assign new_n913_ = new_n911_ & new_n912_;
  assign new_n914_ = v11 & v12;
  assign new_n915_ = new_n665_ & new_n914_;
  assign new_n916_ = ~new_n913_ & ~new_n915_;
  assign new_n917_ = v42 & ~new_n916_;
  assign new_n918_ = v15 & ~v42;
  assign new_n919_ = v14 & new_n918_;
  assign new_n920_ = new_n665_ & new_n919_;
  assign new_n921_ = ~new_n917_ & ~new_n920_;
  assign new_n922_ = ~v44 & ~new_n921_;
  assign new_n923_ = ~v28 & v46;
  assign new_n924_ = new_n817_ & new_n923_;
  assign new_n925_ = ~v43 & ~v46;
  assign new_n926_ = ~v42 & new_n925_;
  assign new_n927_ = new_n516_ & new_n926_;
  assign new_n928_ = ~new_n924_ & ~new_n927_;
  assign new_n929_ = v45 & ~new_n928_;
  assign new_n930_ = v44 & new_n929_;
  assign new_n931_ = ~new_n922_ & ~new_n930_;
  assign \v47.30  = v35 & ~new_n931_;
  assign new_n933_ = ~v45 & new_n865_;
  assign new_n934_ = v43 & new_n933_;
  assign new_n935_ = ~v43 & v45;
  assign new_n936_ = ~new_n934_ & ~new_n935_;
  assign new_n937_ = ~v46 & ~new_n936_;
  assign new_n938_ = ~v9 & new_n937_;
  assign new_n939_ = ~v27 & ~v28;
  assign new_n940_ = v26 & new_n939_;
  assign new_n941_ = new_n912_ & new_n940_;
  assign new_n942_ = ~new_n938_ & ~new_n941_;
  assign new_n943_ = ~v44 & ~new_n942_;
  assign new_n944_ = v17 & ~v43;
  assign new_n945_ = v16 & new_n944_;
  assign new_n946_ = new_n181_ & new_n945_;
  assign new_n947_ = ~new_n943_ & ~new_n946_;
  assign new_n948_ = v42 & ~new_n947_;
  assign new_n949_ = new_n848_ & new_n881_;
  assign new_n950_ = ~new_n885_ & ~new_n949_;
  assign new_n951_ = v44 & ~new_n950_;
  assign new_n952_ = ~new_n948_ & ~new_n951_;
  assign \v47.31  = v35 & ~new_n952_;
  assign new_n954_ = ~v35 & ~v42;
  assign new_n955_ = v43 & new_n954_;
  assign new_n956_ = v44 & new_n955_;
  assign new_n957_ = v45 & new_n956_;
  assign \v47.32  = ~v46 & new_n957_;
  assign new_n959_ = v9 & new_n865_;
  assign new_n960_ = ~v5 & v6;
  assign new_n961_ = ~v4 & v5;
  assign new_n962_ = ~new_n960_ & ~new_n961_;
  assign new_n963_ = ~new_n510_ & ~new_n962_;
  assign new_n964_ = ~new_n959_ & ~new_n963_;
  assign new_n965_ = ~v45 & ~new_n964_;
  assign new_n966_ = ~v44 & new_n965_;
  assign new_n967_ = ~new_n421_ & ~new_n966_;
  assign new_n968_ = v43 & ~new_n967_;
  assign new_n969_ = ~v17 & v44;
  assign new_n970_ = v16 & new_n969_;
  assign new_n971_ = v9 & ~v44;
  assign new_n972_ = ~new_n970_ & ~new_n971_;
  assign new_n973_ = v45 & ~new_n972_;
  assign new_n974_ = ~v43 & new_n973_;
  assign new_n975_ = ~new_n968_ & ~new_n974_;
  assign new_n976_ = v42 & ~new_n975_;
  assign new_n977_ = v9 & new_n350_;
  assign new_n978_ = new_n352_ & new_n977_;
  assign new_n979_ = ~new_n976_ & ~new_n978_;
  assign new_n980_ = ~v46 & ~new_n979_;
  assign \v47.33  = v35 & new_n980_;
  assign new_n982_ = ~v29 & new_n421_;
  assign new_n983_ = ~v4 & new_n960_;
  assign new_n984_ = v6 & ~v29;
  assign new_n985_ = ~v5 & new_n984_;
  assign new_n986_ = ~v5 & ~new_n985_;
  assign new_n987_ = v4 & ~new_n986_;
  assign new_n988_ = ~new_n983_ & ~new_n987_;
  assign new_n989_ = ~new_n510_ & ~new_n988_;
  assign new_n990_ = ~v29 & new_n865_;
  assign new_n991_ = v9 & new_n990_;
  assign new_n992_ = ~new_n989_ & ~new_n991_;
  assign new_n993_ = ~v45 & ~new_n992_;
  assign new_n994_ = ~v44 & new_n993_;
  assign new_n995_ = ~new_n982_ & ~new_n994_;
  assign new_n996_ = v43 & ~new_n995_;
  assign new_n997_ = ~v29 & new_n974_;
  assign new_n998_ = ~new_n996_ & ~new_n997_;
  assign new_n999_ = v42 & ~new_n998_;
  assign new_n1000_ = v12 & ~v29;
  assign new_n1001_ = v9 & new_n1000_;
  assign new_n1002_ = new_n179_ & new_n351_;
  assign new_n1003_ = new_n1001_ & new_n1002_;
  assign new_n1004_ = ~new_n999_ & ~new_n1003_;
  assign new_n1005_ = ~v46 & ~new_n1004_;
  assign \v47.34  = v35 & new_n1005_;
  assign new_n1007_ = ~v44 & ~new_n936_;
  assign new_n1008_ = v42 & new_n1007_;
  assign new_n1009_ = ~new_n353_ & ~new_n1008_;
  assign new_n1010_ = v9 & ~new_n1009_;
  assign new_n1011_ = ~v17 & v42;
  assign new_n1012_ = v16 & new_n1011_;
  assign new_n1013_ = ~v43 & new_n421_;
  assign new_n1014_ = new_n1012_ & new_n1013_;
  assign new_n1015_ = ~new_n1010_ & ~new_n1014_;
  assign new_n1016_ = ~v46 & ~new_n1015_;
  assign new_n1017_ = v35 & new_n1016_;
  assign new_n1018_ = ~v30 & new_n1017_;
  assign \v47.35  = ~v29 & new_n1018_;
  assign new_n1020_ = v24 & ~v25;
  assign new_n1021_ = ~v23 & new_n1020_;
  assign new_n1022_ = new_n912_ & new_n1021_;
  assign new_n1023_ = v11 & ~v12;
  assign new_n1024_ = new_n665_ & new_n1023_;
  assign new_n1025_ = ~new_n1022_ & ~new_n1024_;
  assign new_n1026_ = v42 & ~new_n1025_;
  assign new_n1027_ = ~v15 & ~v42;
  assign new_n1028_ = v14 & new_n1027_;
  assign new_n1029_ = new_n665_ & new_n1028_;
  assign new_n1030_ = ~new_n1026_ & ~new_n1029_;
  assign new_n1031_ = ~v44 & ~new_n1030_;
  assign new_n1032_ = new_n810_ & new_n923_;
  assign new_n1033_ = v4 & ~v5;
  assign new_n1034_ = new_n926_ & new_n1033_;
  assign new_n1035_ = ~new_n1032_ & ~new_n1034_;
  assign new_n1036_ = v45 & ~new_n1035_;
  assign new_n1037_ = v44 & new_n1036_;
  assign new_n1038_ = ~new_n1031_ & ~new_n1037_;
  assign new_n1039_ = v35 & ~new_n1038_;
  assign \v47.36  = new_n182_ | new_n1039_;
  assign new_n1041_ = ~v45 & new_n866_;
  assign new_n1042_ = v9 & new_n1041_;
  assign new_n1043_ = ~v26 & v46;
  assign new_n1044_ = v24 & new_n1043_;
  assign new_n1045_ = ~new_n1042_ & ~new_n1044_;
  assign new_n1046_ = v43 & ~new_n1045_;
  assign new_n1047_ = ~v28 & new_n682_;
  assign new_n1048_ = new_n810_ & new_n1047_;
  assign new_n1049_ = v9 & new_n159_;
  assign new_n1050_ = ~new_n1048_ & ~new_n1049_;
  assign new_n1051_ = ~v43 & ~new_n1050_;
  assign new_n1052_ = ~new_n1046_ & ~new_n1051_;
  assign new_n1053_ = ~v44 & ~new_n1052_;
  assign new_n1054_ = ~v17 & ~v43;
  assign new_n1055_ = v16 & new_n1054_;
  assign new_n1056_ = new_n181_ & new_n1055_;
  assign new_n1057_ = ~new_n1053_ & ~new_n1056_;
  assign new_n1058_ = v42 & ~new_n1057_;
  assign new_n1059_ = new_n841_ & new_n881_;
  assign new_n1060_ = new_n884_ & new_n977_;
  assign new_n1061_ = ~new_n1059_ & ~new_n1060_;
  assign new_n1062_ = v44 & ~new_n1061_;
  assign new_n1063_ = ~new_n1058_ & ~new_n1062_;
  assign \v47.37  = v35 & ~new_n1063_;
  assign new_n1065_ = v43 & new_n230_;
  assign new_n1066_ = v42 & new_n1065_;
  assign new_n1067_ = v35 & new_n1066_;
  assign new_n1068_ = ~v26 & new_n1067_;
  assign \v47.38  = ~v24 & new_n1068_;
  assign new_n1070_ = ~new_n802_ & ~new_n910_;
  assign new_n1071_ = v46 & ~new_n1070_;
  assign new_n1072_ = ~v26 & new_n1071_;
  assign new_n1073_ = ~new_n1042_ & ~new_n1072_;
  assign new_n1074_ = v43 & ~new_n1073_;
  assign new_n1075_ = ~new_n1051_ & ~new_n1074_;
  assign new_n1076_ = ~v44 & ~new_n1075_;
  assign new_n1077_ = ~new_n1056_ & ~new_n1076_;
  assign new_n1078_ = v42 & ~new_n1077_;
  assign new_n1079_ = ~new_n1062_ & ~new_n1078_;
  assign \v47.39  = v35 & ~new_n1079_;
  assign new_n1081_ = ~new_n819_ & ~new_n1020_;
  assign new_n1082_ = v46 & ~new_n1081_;
  assign new_n1083_ = ~v44 & new_n1082_;
  assign new_n1084_ = v43 & new_n1083_;
  assign new_n1085_ = v42 & new_n1084_;
  assign new_n1086_ = v35 & new_n1085_;
  assign \v47.40  = ~v26 & new_n1086_;
  assign new_n1088_ = ~new_n1042_ & ~new_n1043_;
  assign new_n1089_ = v43 & ~new_n1088_;
  assign new_n1090_ = ~new_n1051_ & ~new_n1089_;
  assign new_n1091_ = ~v44 & ~new_n1090_;
  assign new_n1092_ = ~new_n1056_ & ~new_n1091_;
  assign new_n1093_ = v42 & ~new_n1092_;
  assign new_n1094_ = ~new_n1062_ & ~new_n1093_;
  assign \v47.41  = v35 & ~new_n1094_;
  assign new_n1096_ = v6 & ~new_n516_;
  assign new_n1097_ = v5 & ~v6;
  assign new_n1098_ = v4 & new_n1097_;
  assign new_n1099_ = ~new_n1096_ & ~new_n1098_;
  assign new_n1100_ = ~new_n506_ & ~new_n1099_;
  assign new_n1101_ = ~v46 & new_n1100_;
  assign new_n1102_ = ~v45 & new_n1101_;
  assign new_n1103_ = ~v44 & new_n1102_;
  assign new_n1104_ = v43 & new_n1103_;
  assign new_n1105_ = v42 & new_n1104_;
  assign \v47.42  = v35 & new_n1105_;
  assign new_n1107_ = ~v4 & ~v5;
  assign new_n1108_ = ~v5 & ~v32;
  assign new_n1109_ = ~v5 & ~new_n1108_;
  assign new_n1110_ = v4 & ~new_n1109_;
  assign new_n1111_ = ~new_n1107_ & ~new_n1110_;
  assign new_n1112_ = v6 & ~new_n1111_;
  assign new_n1113_ = ~v4 & new_n1097_;
  assign new_n1114_ = ~new_n1112_ & ~new_n1113_;
  assign new_n1115_ = ~new_n506_ & ~new_n1114_;
  assign new_n1116_ = ~v46 & new_n1115_;
  assign new_n1117_ = ~v45 & new_n1116_;
  assign new_n1118_ = ~v44 & new_n1117_;
  assign new_n1119_ = v43 & new_n1118_;
  assign new_n1120_ = v42 & new_n1119_;
  assign \v47.43  = v35 & new_n1120_;
  assign new_n1122_ = v23 & new_n1020_;
  assign new_n1123_ = new_n912_ & new_n1122_;
  assign new_n1124_ = ~v11 & ~v12;
  assign new_n1125_ = new_n665_ & new_n1124_;
  assign new_n1126_ = ~new_n1123_ & ~new_n1125_;
  assign new_n1127_ = v42 & ~new_n1126_;
  assign new_n1128_ = ~v14 & new_n1027_;
  assign new_n1129_ = new_n665_ & new_n1128_;
  assign new_n1130_ = ~new_n1127_ & ~new_n1129_;
  assign new_n1131_ = ~v44 & ~new_n1130_;
  assign new_n1132_ = new_n799_ & new_n923_;
  assign new_n1133_ = new_n926_ & new_n1107_;
  assign new_n1134_ = ~new_n1132_ & ~new_n1133_;
  assign new_n1135_ = v45 & ~new_n1134_;
  assign new_n1136_ = v44 & new_n1135_;
  assign new_n1137_ = ~new_n1131_ & ~new_n1136_;
  assign \v47.45  = v35 & ~new_n1137_;
  assign new_n1139_ = v26 & v42;
  assign new_n1140_ = new_n608_ & new_n1139_;
  assign new_n1141_ = v23 & new_n421_;
  assign new_n1142_ = ~new_n1140_ & ~new_n1141_;
  assign new_n1143_ = ~v25 & ~new_n1142_;
  assign new_n1144_ = v25 & v26;
  assign new_n1145_ = new_n611_ & new_n1144_;
  assign new_n1146_ = ~new_n1143_ & ~new_n1145_;
  assign new_n1147_ = v24 & ~new_n1146_;
  assign new_n1148_ = v27 & ~v28;
  assign new_n1149_ = v26 & new_n1148_;
  assign new_n1150_ = new_n805_ & new_n1149_;
  assign new_n1151_ = ~new_n1147_ & ~new_n1150_;
  assign new_n1152_ = v46 & ~new_n1151_;
  assign new_n1153_ = ~v16 & new_n1011_;
  assign new_n1154_ = new_n159_ & new_n890_;
  assign new_n1155_ = new_n1153_ & new_n1154_;
  assign new_n1156_ = ~new_n1152_ & ~new_n1155_;
  assign \v47.46  = v35 & ~new_n1156_;
  assign new_n1158_ = v26 & new_n1067_;
  assign \v47.47  = ~v24 & new_n1158_;
  assign new_n1160_ = v23 & ~v25;
  assign new_n1161_ = new_n421_ & new_n1160_;
  assign new_n1162_ = ~new_n1145_ & ~new_n1161_;
  assign new_n1163_ = v24 & ~new_n1162_;
  assign new_n1164_ = ~v25 & v43;
  assign new_n1165_ = ~v24 & new_n1164_;
  assign new_n1166_ = ~v43 & ~v45;
  assign new_n1167_ = new_n1148_ & new_n1166_;
  assign new_n1168_ = ~new_n1165_ & ~new_n1167_;
  assign new_n1169_ = ~v44 & ~new_n1168_;
  assign new_n1170_ = v42 & new_n1169_;
  assign new_n1171_ = v26 & new_n1170_;
  assign new_n1172_ = ~new_n1163_ & ~new_n1171_;
  assign new_n1173_ = v46 & ~new_n1172_;
  assign new_n1174_ = ~new_n1155_ & ~new_n1173_;
  assign \v47.48  = v35 & ~new_n1174_;
  assign \v47.49  = v26 & new_n1086_;
  assign new_n1177_ = ~v43 & ~new_n1167_;
  assign new_n1178_ = v46 & ~new_n1177_;
  assign new_n1179_ = ~v44 & new_n1178_;
  assign new_n1180_ = v26 & new_n1179_;
  assign new_n1181_ = ~v16 & new_n1054_;
  assign new_n1182_ = new_n181_ & new_n1181_;
  assign new_n1183_ = ~new_n1180_ & ~new_n1182_;
  assign new_n1184_ = v42 & ~new_n1183_;
  assign new_n1185_ = new_n590_ & new_n1122_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign \v47.50  = v35 & ~new_n1186_;
  assign new_n1188_ = ~v45 & new_n130_;
  assign new_n1189_ = ~v46 & ~new_n1188_;
  assign new_n1190_ = v43 & ~new_n1189_;
  assign new_n1191_ = ~v43 & new_n159_;
  assign new_n1192_ = ~new_n1190_ & ~new_n1191_;
  assign new_n1193_ = ~v44 & ~new_n1192_;
  assign new_n1194_ = ~new_n877_ & ~new_n1193_;
  assign new_n1195_ = v42 & ~new_n1194_;
  assign new_n1196_ = v43 & new_n220_;
  assign new_n1197_ = ~v43 & new_n230_;
  assign new_n1198_ = new_n641_ & new_n1197_;
  assign new_n1199_ = ~new_n1196_ & ~new_n1198_;
  assign new_n1200_ = ~v45 & ~new_n1199_;
  assign new_n1201_ = ~v43 & ~v44;
  assign new_n1202_ = new_n159_ & new_n1201_;
  assign new_n1203_ = ~new_n1200_ & ~new_n1202_;
  assign new_n1204_ = ~v42 & ~new_n1203_;
  assign new_n1205_ = ~new_n1195_ & ~new_n1204_;
  assign new_n1206_ = v35 & ~new_n1205_;
  assign \v47.51  = new_n182_ | new_n1206_;
  assign new_n1208_ = ~v40 & ~new_n203_;
  assign new_n1209_ = ~v39 & ~new_n1208_;
  assign new_n1210_ = ~v38 & ~new_n594_;
  assign new_n1211_ = v37 & new_n1210_;
  assign new_n1212_ = ~new_n1209_ & new_n1211_;
  assign new_n1213_ = ~new_n135_ & new_n1212_;
  assign new_n1214_ = ~v28 & new_n1213_;
  assign new_n1215_ = ~new_n136_ & new_n1214_;
  assign new_n1216_ = v46 & ~new_n1215_;
  assign new_n1217_ = ~new_n130_ & ~new_n1216_;
  assign new_n1218_ = v43 & ~new_n1217_;
  assign new_n1219_ = v42 & new_n1218_;
  assign new_n1220_ = v13 & ~v22;
  assign new_n1221_ = v21 & ~new_n1220_;
  assign new_n1222_ = v19 & ~new_n1221_;
  assign new_n1223_ = v18 & new_n1222_;
  assign new_n1224_ = ~new_n131_ & ~new_n641_;
  assign new_n1225_ = v20 & new_n1224_;
  assign new_n1226_ = ~new_n1223_ & new_n1225_;
  assign new_n1227_ = v46 & ~new_n1226_;
  assign new_n1228_ = ~v43 & new_n1227_;
  assign new_n1229_ = ~v42 & new_n1228_;
  assign new_n1230_ = ~new_n1219_ & ~new_n1229_;
  assign new_n1231_ = ~v45 & ~new_n1230_;
  assign new_n1232_ = ~new_n1191_ & ~new_n1231_;
  assign new_n1233_ = ~v44 & ~new_n1232_;
  assign new_n1234_ = v43 & ~v45;
  assign new_n1235_ = ~v42 & new_n1234_;
  assign new_n1236_ = v42 & new_n935_;
  assign new_n1237_ = ~new_n1235_ & ~new_n1236_;
  assign new_n1238_ = ~v46 & ~new_n1237_;
  assign new_n1239_ = v44 & new_n1238_;
  assign new_n1240_ = ~new_n1233_ & ~new_n1239_;
  assign new_n1241_ = v35 & ~new_n1240_;
  assign \v47.52  = new_n182_ | new_n1241_;
  assign new_n1243_ = ~v45 & new_n129_;
  assign new_n1244_ = v43 & new_n1243_;
  assign new_n1245_ = ~new_n935_ & ~new_n1244_;
  assign new_n1246_ = ~v44 & ~new_n1245_;
  assign new_n1247_ = ~new_n1013_ & ~new_n1246_;
  assign new_n1248_ = v42 & ~new_n1247_;
  assign new_n1249_ = ~new_n352_ & ~new_n390_;
  assign new_n1250_ = ~v42 & ~new_n1249_;
  assign new_n1251_ = ~new_n1248_ & ~new_n1250_;
  assign new_n1252_ = v35 & ~new_n1251_;
  assign new_n1253_ = v43 & new_n421_;
  assign new_n1254_ = new_n954_ & new_n1253_;
  assign new_n1255_ = ~new_n1252_ & ~new_n1254_;
  assign \v47.54  = ~v46 & ~new_n1255_;
  assign new_n1257_ = v35 & v42;
  assign new_n1258_ = ~v43 & new_n1257_;
  assign new_n1259_ = v44 & new_n1258_;
  assign new_n1260_ = ~v45 & new_n1259_;
  assign \v47.55  = ~v46 & new_n1260_;
  assign new_n1262_ = v35 & ~v42;
  assign new_n1263_ = ~v43 & new_n1262_;
  assign new_n1264_ = v44 & new_n1263_;
  assign new_n1265_ = ~v45 & new_n1264_;
  assign \v47.56  = ~v46 & new_n1265_;
  assign \v47.58  = ~v28 & new_n1067_;
  assign \v47.59  = v28 & new_n1067_;
  assign new_n1269_ = v35 & new_n939_;
  assign new_n1270_ = v42 & new_n1269_;
  assign new_n1271_ = v43 & new_n1270_;
  assign new_n1272_ = ~v44 & new_n1271_;
  assign \v47.60  = v46 & new_n1272_;
  assign new_n1274_ = ~v42 & new_n230_;
  assign new_n1275_ = new_n641_ & new_n1274_;
  assign new_n1276_ = v42 & new_n220_;
  assign new_n1277_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1278_ = ~v45 & ~new_n1277_;
  assign new_n1279_ = ~v43 & new_n1278_;
  assign \v47.62  = v35 & new_n1279_;
  assign new_n1281_ = ~v28 & v42;
  assign new_n1282_ = v27 & new_n1281_;
  assign new_n1283_ = new_n1065_ & new_n1282_;
  assign new_n1284_ = ~v42 & ~v43;
  assign new_n1285_ = new_n550_ & new_n1284_;
  assign new_n1286_ = ~new_n1283_ & ~new_n1285_;
  assign \v47.63  = v35 & ~new_n1286_;
  assign new_n1288_ = v28 & new_n1065_;
  assign new_n1289_ = ~v43 & new_n220_;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_;
  assign new_n1291_ = ~v45 & ~new_n1290_;
  assign new_n1292_ = v42 & new_n1291_;
  assign \v47.64  = v35 & new_n1292_;
  assign new_n1294_ = ~v20 & v28;
  assign new_n1295_ = v35 & new_n1294_;
  assign new_n1296_ = v42 & new_n1295_;
  assign new_n1297_ = v43 & new_n1296_;
  assign new_n1298_ = ~v44 & new_n1297_;
  assign new_n1299_ = ~v45 & new_n1298_;
  assign \v47.65  = v46 & new_n1299_;
  assign new_n1301_ = v20 & v28;
  assign new_n1302_ = new_n1065_ & new_n1301_;
  assign new_n1303_ = ~new_n1289_ & ~new_n1302_;
  assign new_n1304_ = ~v45 & ~new_n1303_;
  assign new_n1305_ = v42 & new_n1304_;
  assign \v47.66  = v35 & new_n1305_;
  assign new_n1307_ = v35 & new_n835_;
  assign new_n1308_ = v42 & new_n1307_;
  assign new_n1309_ = v43 & new_n1308_;
  assign new_n1310_ = ~v44 & new_n1309_;
  assign new_n1311_ = ~v45 & new_n1310_;
  assign \v47.68  = v46 & new_n1311_;
  assign new_n1313_ = v35 & new_n850_;
  assign new_n1314_ = v42 & new_n1313_;
  assign new_n1315_ = v43 & new_n1314_;
  assign new_n1316_ = ~v44 & new_n1315_;
  assign new_n1317_ = ~v45 & new_n1316_;
  assign \v47.69  = v46 & new_n1317_;
  assign new_n1319_ = ~v46 & ~new_n1251_;
  assign new_n1320_ = new_n682_ & new_n1201_;
  assign new_n1321_ = new_n751_ & new_n1320_;
  assign new_n1322_ = ~new_n1319_ & ~new_n1321_;
  assign new_n1323_ = v35 & ~new_n1322_;
  assign \v47.70  = new_n182_ | new_n1323_;
  assign \v47.11  = 1'b0;
  assign \v47.44  = 1'b0;
  assign \v47.53  = 1'b0;
  assign \v47.61  = 1'b0;
  assign \v47.67  = 1'b0;
  assign \v47.57  = \v47.55 ;
  assign \v47.71  = \v47.54 ;
endmodule


