// Benchmark "bar" written by ABC on Tue Sep  5 17:54:35 2023

module bar ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1044_, new_n1045_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1279_,
    new_n1280_, new_n1281_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1349_, new_n1350_, new_n1351_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1497_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1517_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1539_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1591_, new_n1592_, new_n1593_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1621_, new_n1622_, new_n1623_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1721_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1755_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1776_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1799_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1822_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1910_, new_n1911_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1979_, new_n1980_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1994_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2019_,
    new_n2021_, new_n2023_, new_n2025_, new_n2028_, new_n2029_, new_n2032_,
    new_n2035_, new_n2036_, new_n2039_, new_n2042_, new_n2044_, new_n2047_,
    new_n2050_, new_n2053_, new_n2056_, new_n2058_, new_n2060_, new_n2062_,
    new_n2064_, new_n2065_, new_n2068_, new_n2069_, new_n2071_, new_n2072_,
    new_n2075_, new_n2076_, new_n2079_, new_n2081_, new_n2083_, new_n2086_,
    new_n2089_, new_n2092_, new_n2095_, new_n2097_, new_n2100_, new_n2102_,
    new_n2104_, new_n2106_, new_n2108_, new_n2111_, new_n2114_, new_n2117_,
    new_n2120_, new_n2122_;
  INV_X1     g0000(.I(\shift[6] ), .ZN(new_n264_));
  INV_X1     g0001(.I(\shift[5] ), .ZN(new_n265_));
  NOR2_X1    g0002(.A1(\shift[2] ), .A2(\shift[3] ), .ZN(new_n266_));
  INV_X1     g0003(.I(new_n266_), .ZN(new_n267_));
  NAND3_X1   g0004(.A1(new_n267_), .A2(\shift[4] ), .A3(new_n265_), .ZN(new_n268_));
  NAND2_X1   g0005(.A1(new_n268_), .A2(new_n264_), .ZN(new_n269_));
  INV_X1     g0006(.I(\shift[4] ), .ZN(new_n270_));
  NOR2_X1    g0007(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1     g0008(.I(new_n271_), .ZN(new_n272_));
  NAND2_X1   g0009(.A1(new_n266_), .A2(new_n270_), .ZN(new_n273_));
  NAND3_X1   g0010(.A1(new_n272_), .A2(new_n265_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1     g0011(.I(\shift[2] ), .ZN(new_n275_));
  INV_X1     g0012(.I(\shift[3] ), .ZN(new_n276_));
  NOR2_X1    g0013(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1    g0014(.A1(\shift[2] ), .A2(\shift[3] ), .ZN(new_n278_));
  INV_X1     g0015(.I(\shift[0] ), .ZN(new_n279_));
  OAI21_X1   g0016(.A1(\a[40] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n280_));
  NOR3_X1    g0017(.A1(new_n279_), .A2(\a[37] ), .A3(\shift[1] ), .ZN(new_n281_));
  XOR2_X1    g0018(.A1(new_n280_), .A2(new_n281_), .Z(new_n282_));
  XNOR2_X1   g0019(.A1(\shift[0] ), .A2(\shift[1] ), .ZN(new_n283_));
  INV_X1     g0020(.I(\shift[1] ), .ZN(new_n284_));
  NOR2_X1    g0021(.A1(new_n284_), .A2(\a[38] ), .ZN(new_n285_));
  NOR2_X1    g0022(.A1(\a[39] ), .A2(\shift[1] ), .ZN(new_n286_));
  NOR4_X1    g0023(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  NOR2_X1    g0024(.A1(\shift[4] ), .A2(\shift[5] ), .ZN(new_n288_));
  NOR2_X1    g0025(.A1(new_n274_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1   g0026(.A1(new_n289_), .A2(new_n264_), .B(new_n269_), .ZN(\result[0] ));
  INV_X1     g0027(.I(new_n277_), .ZN(new_n291_));
  NOR2_X1    g0028(.A1(\a[101] ), .A2(\shift[1] ), .ZN(new_n292_));
  NOR3_X1    g0029(.A1(new_n279_), .A2(\a[98] ), .A3(\shift[1] ), .ZN(new_n293_));
  INV_X1     g0030(.I(new_n293_), .ZN(new_n294_));
  NOR2_X1    g0031(.A1(new_n292_), .A2(\shift[0] ), .ZN(new_n295_));
  INV_X1     g0032(.I(\a[98] ), .ZN(new_n296_));
  NAND3_X1   g0033(.A1(new_n296_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n297_));
  NAND2_X1   g0034(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1   g0035(.A1(new_n298_), .A2(new_n294_), .ZN(new_n299_));
  NOR2_X1    g0036(.A1(new_n284_), .A2(\a[99] ), .ZN(new_n300_));
  NOR2_X1    g0037(.A1(\a[100] ), .A2(\shift[1] ), .ZN(new_n301_));
  NOR3_X1    g0038(.A1(new_n283_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1   g0039(.A1(new_n299_), .A2(new_n302_), .B(new_n291_), .ZN(new_n303_));
  NOR2_X1    g0040(.A1(\a[113] ), .A2(\shift[1] ), .ZN(new_n304_));
  NOR3_X1    g0041(.A1(new_n279_), .A2(\a[110] ), .A3(\shift[1] ), .ZN(new_n305_));
  NOR3_X1    g0042(.A1(new_n279_), .A2(\a[110] ), .A3(\shift[1] ), .ZN(new_n306_));
  NOR3_X1    g0043(.A1(new_n306_), .A2(\shift[0] ), .A3(new_n304_), .ZN(new_n307_));
  NOR2_X1    g0044(.A1(new_n307_), .A2(new_n305_), .ZN(new_n308_));
  XOR2_X1    g0045(.A1(\shift[0] ), .A2(\shift[1] ), .Z(new_n309_));
  NOR2_X1    g0046(.A1(new_n284_), .A2(\a[111] ), .ZN(new_n310_));
  NOR2_X1    g0047(.A1(\a[112] ), .A2(\shift[1] ), .ZN(new_n311_));
  NOR2_X1    g0048(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1   g0049(.A1(new_n312_), .A2(new_n309_), .ZN(new_n313_));
  OAI21_X1   g0050(.A1(new_n308_), .A2(new_n313_), .B(new_n278_), .ZN(new_n314_));
  INV_X1     g0051(.I(new_n278_), .ZN(new_n315_));
  NOR2_X1    g0052(.A1(\a[105] ), .A2(\shift[1] ), .ZN(new_n316_));
  NOR3_X1    g0053(.A1(new_n279_), .A2(\a[102] ), .A3(\shift[1] ), .ZN(new_n317_));
  NOR3_X1    g0054(.A1(new_n279_), .A2(\a[102] ), .A3(\shift[1] ), .ZN(new_n318_));
  NOR3_X1    g0055(.A1(new_n318_), .A2(\shift[0] ), .A3(new_n316_), .ZN(new_n319_));
  NOR2_X1    g0056(.A1(new_n319_), .A2(new_n317_), .ZN(new_n320_));
  INV_X1     g0057(.I(\a[103] ), .ZN(new_n321_));
  NOR2_X1    g0058(.A1(\a[104] ), .A2(\shift[1] ), .ZN(new_n322_));
  AOI21_X1   g0059(.A1(new_n321_), .A2(\shift[1] ), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1   g0060(.A1(new_n309_), .A2(new_n323_), .ZN(new_n324_));
  NOR3_X1    g0061(.A1(new_n320_), .A2(new_n315_), .A3(new_n324_), .ZN(new_n325_));
  NOR2_X1    g0062(.A1(\a[109] ), .A2(\shift[1] ), .ZN(new_n326_));
  NOR3_X1    g0063(.A1(new_n279_), .A2(\a[106] ), .A3(\shift[1] ), .ZN(new_n327_));
  NOR3_X1    g0064(.A1(new_n279_), .A2(\a[106] ), .A3(\shift[1] ), .ZN(new_n328_));
  NOR3_X1    g0065(.A1(new_n328_), .A2(\shift[0] ), .A3(new_n326_), .ZN(new_n329_));
  NOR2_X1    g0066(.A1(new_n329_), .A2(new_n327_), .ZN(new_n330_));
  NOR2_X1    g0067(.A1(new_n284_), .A2(\a[107] ), .ZN(new_n331_));
  NOR2_X1    g0068(.A1(\a[108] ), .A2(\shift[1] ), .ZN(new_n332_));
  NOR2_X1    g0069(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1   g0070(.A1(new_n333_), .A2(new_n309_), .ZN(new_n334_));
  NOR3_X1    g0071(.A1(new_n330_), .A2(new_n315_), .A3(new_n334_), .ZN(new_n335_));
  NOR4_X1    g0072(.A1(new_n303_), .A2(new_n325_), .A3(new_n335_), .A4(new_n314_), .ZN(new_n336_));
  NOR2_X1    g0073(.A1(new_n336_), .A2(new_n270_), .ZN(new_n337_));
  NOR2_X1    g0074(.A1(\a[117] ), .A2(\shift[1] ), .ZN(new_n338_));
  NOR3_X1    g0075(.A1(new_n279_), .A2(\a[114] ), .A3(\shift[1] ), .ZN(new_n339_));
  NOR3_X1    g0076(.A1(new_n279_), .A2(\a[114] ), .A3(\shift[1] ), .ZN(new_n340_));
  NOR3_X1    g0077(.A1(new_n340_), .A2(\shift[0] ), .A3(new_n338_), .ZN(new_n341_));
  NOR2_X1    g0078(.A1(new_n341_), .A2(new_n339_), .ZN(new_n342_));
  NOR2_X1    g0079(.A1(new_n284_), .A2(\a[115] ), .ZN(new_n343_));
  NOR2_X1    g0080(.A1(\a[116] ), .A2(\shift[1] ), .ZN(new_n344_));
  NOR2_X1    g0081(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1   g0082(.A1(new_n345_), .A2(new_n309_), .ZN(new_n346_));
  OAI21_X1   g0083(.A1(new_n342_), .A2(new_n346_), .B(new_n277_), .ZN(new_n347_));
  INV_X1     g0084(.I(\a[0] ), .ZN(new_n348_));
  NAND2_X1   g0085(.A1(new_n348_), .A2(\shift[0] ), .ZN(new_n349_));
  OR2_X2     g0086(.A1(\a[127] ), .A2(\shift[0] ), .Z(new_n350_));
  NAND2_X1   g0087(.A1(new_n350_), .A2(new_n349_), .ZN(new_n351_));
  INV_X1     g0088(.I(\a[1] ), .ZN(new_n352_));
  NAND2_X1   g0089(.A1(\a[126] ), .A2(\shift[1] ), .ZN(new_n353_));
  NAND3_X1   g0090(.A1(new_n353_), .A2(new_n352_), .A3(\shift[0] ), .ZN(new_n354_));
  INV_X1     g0091(.I(new_n354_), .ZN(new_n355_));
  AOI21_X1   g0092(.A1(new_n352_), .A2(\shift[0] ), .B(new_n353_), .ZN(new_n356_));
  NOR4_X1    g0093(.A1(new_n355_), .A2(new_n351_), .A3(new_n283_), .A4(new_n356_), .ZN(new_n357_));
  NOR2_X1    g0094(.A1(new_n357_), .A2(new_n315_), .ZN(new_n358_));
  NOR2_X1    g0095(.A1(\a[121] ), .A2(\shift[1] ), .ZN(new_n359_));
  NOR2_X1    g0096(.A1(new_n359_), .A2(\shift[0] ), .ZN(new_n360_));
  NOR3_X1    g0097(.A1(new_n279_), .A2(\a[118] ), .A3(\shift[1] ), .ZN(new_n361_));
  XOR2_X1    g0098(.A1(new_n360_), .A2(new_n361_), .Z(new_n362_));
  NOR2_X1    g0099(.A1(new_n284_), .A2(\a[119] ), .ZN(new_n363_));
  NOR2_X1    g0100(.A1(\a[120] ), .A2(\shift[1] ), .ZN(new_n364_));
  NOR3_X1    g0101(.A1(new_n283_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1   g0102(.A1(new_n362_), .A2(new_n365_), .A3(new_n278_), .ZN(new_n366_));
  NOR2_X1    g0103(.A1(\a[125] ), .A2(\shift[1] ), .ZN(new_n367_));
  NOR3_X1    g0104(.A1(new_n279_), .A2(\a[122] ), .A3(\shift[1] ), .ZN(new_n368_));
  INV_X1     g0105(.I(new_n368_), .ZN(new_n369_));
  NOR2_X1    g0106(.A1(new_n367_), .A2(\shift[0] ), .ZN(new_n370_));
  INV_X1     g0107(.I(\a[122] ), .ZN(new_n371_));
  NAND3_X1   g0108(.A1(new_n371_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n372_));
  NAND2_X1   g0109(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1   g0110(.A1(new_n373_), .A2(new_n369_), .ZN(new_n374_));
  INV_X1     g0111(.I(\a[123] ), .ZN(new_n375_));
  NOR2_X1    g0112(.A1(\a[124] ), .A2(\shift[1] ), .ZN(new_n376_));
  AOI21_X1   g0113(.A1(new_n375_), .A2(\shift[1] ), .B(new_n376_), .ZN(new_n377_));
  NAND4_X1   g0114(.A1(new_n374_), .A2(new_n278_), .A3(new_n309_), .A4(new_n377_), .ZN(new_n378_));
  NAND4_X1   g0115(.A1(new_n366_), .A2(new_n358_), .A3(new_n378_), .A4(new_n347_), .ZN(new_n379_));
  OAI21_X1   g0116(.A1(new_n379_), .A2(new_n270_), .B(new_n265_), .ZN(new_n380_));
  NOR2_X1    g0117(.A1(new_n380_), .A2(new_n337_), .ZN(new_n381_));
  NOR2_X1    g0118(.A1(\a[85] ), .A2(\shift[1] ), .ZN(new_n382_));
  NOR3_X1    g0119(.A1(new_n279_), .A2(\a[82] ), .A3(\shift[1] ), .ZN(new_n383_));
  INV_X1     g0120(.I(new_n383_), .ZN(new_n384_));
  NOR2_X1    g0121(.A1(new_n382_), .A2(\shift[0] ), .ZN(new_n385_));
  INV_X1     g0122(.I(\a[82] ), .ZN(new_n386_));
  NAND3_X1   g0123(.A1(new_n386_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n387_));
  NAND2_X1   g0124(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1   g0125(.A1(new_n388_), .A2(new_n384_), .ZN(new_n389_));
  NOR2_X1    g0126(.A1(new_n284_), .A2(\a[83] ), .ZN(new_n390_));
  NOR2_X1    g0127(.A1(\a[84] ), .A2(\shift[1] ), .ZN(new_n391_));
  NOR3_X1    g0128(.A1(new_n283_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1   g0129(.A1(new_n389_), .A2(new_n392_), .B(new_n291_), .ZN(new_n393_));
  NOR2_X1    g0130(.A1(\a[97] ), .A2(\shift[1] ), .ZN(new_n394_));
  NOR3_X1    g0131(.A1(new_n279_), .A2(\a[94] ), .A3(\shift[1] ), .ZN(new_n395_));
  NOR3_X1    g0132(.A1(new_n279_), .A2(\a[94] ), .A3(\shift[1] ), .ZN(new_n396_));
  NOR3_X1    g0133(.A1(new_n396_), .A2(\shift[0] ), .A3(new_n394_), .ZN(new_n397_));
  NOR2_X1    g0134(.A1(new_n397_), .A2(new_n395_), .ZN(new_n398_));
  NOR2_X1    g0135(.A1(new_n284_), .A2(\a[95] ), .ZN(new_n399_));
  NOR2_X1    g0136(.A1(\a[96] ), .A2(\shift[1] ), .ZN(new_n400_));
  NOR2_X1    g0137(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1   g0138(.A1(new_n401_), .A2(new_n309_), .ZN(new_n402_));
  OAI21_X1   g0139(.A1(new_n398_), .A2(new_n402_), .B(new_n278_), .ZN(new_n403_));
  NOR2_X1    g0140(.A1(new_n393_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1    g0141(.A1(\a[89] ), .A2(\shift[1] ), .ZN(new_n405_));
  NOR3_X1    g0142(.A1(new_n279_), .A2(\a[86] ), .A3(\shift[1] ), .ZN(new_n406_));
  INV_X1     g0143(.I(new_n406_), .ZN(new_n407_));
  NOR2_X1    g0144(.A1(new_n405_), .A2(\shift[0] ), .ZN(new_n408_));
  INV_X1     g0145(.I(\a[86] ), .ZN(new_n409_));
  NAND3_X1   g0146(.A1(new_n409_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n410_));
  NAND2_X1   g0147(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1   g0148(.A1(new_n411_), .A2(new_n407_), .ZN(new_n412_));
  NOR2_X1    g0149(.A1(new_n284_), .A2(\a[87] ), .ZN(new_n413_));
  NOR2_X1    g0150(.A1(\a[88] ), .A2(\shift[1] ), .ZN(new_n414_));
  NOR3_X1    g0151(.A1(new_n283_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1   g0152(.A1(new_n412_), .A2(new_n415_), .A3(new_n278_), .ZN(new_n416_));
  NOR2_X1    g0153(.A1(\a[93] ), .A2(\shift[1] ), .ZN(new_n417_));
  NOR3_X1    g0154(.A1(new_n279_), .A2(\a[90] ), .A3(\shift[1] ), .ZN(new_n418_));
  INV_X1     g0155(.I(new_n418_), .ZN(new_n419_));
  NOR2_X1    g0156(.A1(new_n417_), .A2(\shift[0] ), .ZN(new_n420_));
  INV_X1     g0157(.I(\a[90] ), .ZN(new_n421_));
  NAND3_X1   g0158(.A1(new_n421_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n422_));
  NAND2_X1   g0159(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1   g0160(.A1(new_n423_), .A2(new_n419_), .ZN(new_n424_));
  NOR2_X1    g0161(.A1(new_n284_), .A2(\a[91] ), .ZN(new_n425_));
  NOR2_X1    g0162(.A1(\a[92] ), .A2(\shift[1] ), .ZN(new_n426_));
  NOR3_X1    g0163(.A1(new_n283_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1   g0164(.A1(new_n424_), .A2(new_n427_), .A3(new_n278_), .ZN(new_n428_));
  NAND4_X1   g0165(.A1(new_n404_), .A2(new_n270_), .A3(new_n416_), .A4(new_n428_), .ZN(new_n429_));
  NOR2_X1    g0166(.A1(\a[69] ), .A2(\shift[1] ), .ZN(new_n430_));
  NOR3_X1    g0167(.A1(new_n279_), .A2(\a[66] ), .A3(\shift[1] ), .ZN(new_n431_));
  NOR3_X1    g0168(.A1(new_n279_), .A2(\a[66] ), .A3(\shift[1] ), .ZN(new_n432_));
  NOR3_X1    g0169(.A1(new_n432_), .A2(\shift[0] ), .A3(new_n430_), .ZN(new_n433_));
  NOR2_X1    g0170(.A1(new_n433_), .A2(new_n431_), .ZN(new_n434_));
  NOR2_X1    g0171(.A1(new_n284_), .A2(\a[67] ), .ZN(new_n435_));
  NOR2_X1    g0172(.A1(\a[68] ), .A2(\shift[1] ), .ZN(new_n436_));
  NOR2_X1    g0173(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1   g0174(.A1(new_n437_), .A2(new_n309_), .ZN(new_n438_));
  OAI21_X1   g0175(.A1(new_n434_), .A2(new_n438_), .B(new_n277_), .ZN(new_n439_));
  NOR2_X1    g0176(.A1(new_n315_), .A2(new_n270_), .ZN(new_n440_));
  INV_X1     g0177(.I(new_n440_), .ZN(new_n441_));
  NOR2_X1    g0178(.A1(\a[81] ), .A2(\shift[1] ), .ZN(new_n442_));
  NOR3_X1    g0179(.A1(new_n279_), .A2(\a[78] ), .A3(\shift[1] ), .ZN(new_n443_));
  NOR3_X1    g0180(.A1(new_n279_), .A2(\a[78] ), .A3(\shift[1] ), .ZN(new_n444_));
  NOR3_X1    g0181(.A1(new_n444_), .A2(\shift[0] ), .A3(new_n442_), .ZN(new_n445_));
  NOR2_X1    g0182(.A1(new_n445_), .A2(new_n443_), .ZN(new_n446_));
  NOR2_X1    g0183(.A1(new_n284_), .A2(\a[79] ), .ZN(new_n447_));
  NOR2_X1    g0184(.A1(\a[80] ), .A2(\shift[1] ), .ZN(new_n448_));
  NOR2_X1    g0185(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1   g0186(.A1(new_n449_), .A2(new_n309_), .ZN(new_n450_));
  NOR2_X1    g0187(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1    g0188(.A1(new_n451_), .A2(new_n441_), .ZN(new_n452_));
  NOR2_X1    g0189(.A1(\a[73] ), .A2(\shift[1] ), .ZN(new_n453_));
  NOR2_X1    g0190(.A1(new_n453_), .A2(\shift[0] ), .ZN(new_n454_));
  NOR3_X1    g0191(.A1(new_n279_), .A2(\a[70] ), .A3(\shift[1] ), .ZN(new_n455_));
  XOR2_X1    g0192(.A1(new_n454_), .A2(new_n455_), .Z(new_n456_));
  INV_X1     g0193(.I(\a[71] ), .ZN(new_n457_));
  NOR2_X1    g0194(.A1(\a[72] ), .A2(\shift[1] ), .ZN(new_n458_));
  AOI21_X1   g0195(.A1(new_n457_), .A2(\shift[1] ), .B(new_n458_), .ZN(new_n459_));
  AND2_X2    g0196(.A1(new_n309_), .A2(new_n459_), .Z(new_n460_));
  NAND3_X1   g0197(.A1(new_n456_), .A2(new_n460_), .A3(new_n278_), .ZN(new_n461_));
  NOR2_X1    g0198(.A1(\a[77] ), .A2(\shift[1] ), .ZN(new_n462_));
  NOR3_X1    g0199(.A1(new_n279_), .A2(\a[74] ), .A3(\shift[1] ), .ZN(new_n463_));
  INV_X1     g0200(.I(new_n463_), .ZN(new_n464_));
  NOR2_X1    g0201(.A1(new_n462_), .A2(\shift[0] ), .ZN(new_n465_));
  INV_X1     g0202(.I(\a[74] ), .ZN(new_n466_));
  NAND3_X1   g0203(.A1(new_n466_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n467_));
  NAND2_X1   g0204(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1   g0205(.A1(new_n468_), .A2(new_n464_), .ZN(new_n469_));
  NOR2_X1    g0206(.A1(new_n284_), .A2(\a[75] ), .ZN(new_n470_));
  NOR2_X1    g0207(.A1(\a[76] ), .A2(\shift[1] ), .ZN(new_n471_));
  NOR2_X1    g0208(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1   g0209(.A1(new_n469_), .A2(new_n278_), .A3(new_n309_), .A4(new_n472_), .ZN(new_n473_));
  NAND4_X1   g0210(.A1(new_n452_), .A2(new_n439_), .A3(new_n461_), .A4(new_n473_), .ZN(new_n474_));
  NAND3_X1   g0211(.A1(new_n429_), .A2(new_n474_), .A3(new_n265_), .ZN(new_n475_));
  OAI21_X1   g0212(.A1(new_n381_), .A2(new_n475_), .B(new_n264_), .ZN(new_n476_));
  NOR2_X1    g0213(.A1(\a[53] ), .A2(\shift[1] ), .ZN(new_n477_));
  NOR3_X1    g0214(.A1(new_n279_), .A2(\a[50] ), .A3(\shift[1] ), .ZN(new_n478_));
  INV_X1     g0215(.I(new_n478_), .ZN(new_n479_));
  NOR2_X1    g0216(.A1(new_n477_), .A2(\shift[0] ), .ZN(new_n480_));
  INV_X1     g0217(.I(\a[50] ), .ZN(new_n481_));
  NAND3_X1   g0218(.A1(new_n481_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n482_));
  NAND2_X1   g0219(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1   g0220(.A1(new_n483_), .A2(new_n479_), .ZN(new_n484_));
  NOR2_X1    g0221(.A1(new_n284_), .A2(\a[51] ), .ZN(new_n485_));
  NOR2_X1    g0222(.A1(\a[52] ), .A2(\shift[1] ), .ZN(new_n486_));
  NOR3_X1    g0223(.A1(new_n283_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1   g0224(.A1(new_n484_), .A2(new_n487_), .B(new_n291_), .ZN(new_n488_));
  NOR2_X1    g0225(.A1(\a[65] ), .A2(\shift[1] ), .ZN(new_n489_));
  NOR3_X1    g0226(.A1(new_n279_), .A2(\a[62] ), .A3(\shift[1] ), .ZN(new_n490_));
  NOR3_X1    g0227(.A1(new_n279_), .A2(\a[62] ), .A3(\shift[1] ), .ZN(new_n491_));
  NOR3_X1    g0228(.A1(new_n491_), .A2(\shift[0] ), .A3(new_n489_), .ZN(new_n492_));
  NOR2_X1    g0229(.A1(new_n492_), .A2(new_n490_), .ZN(new_n493_));
  INV_X1     g0230(.I(\a[63] ), .ZN(new_n494_));
  NOR2_X1    g0231(.A1(\a[64] ), .A2(\shift[1] ), .ZN(new_n495_));
  AOI21_X1   g0232(.A1(new_n494_), .A2(\shift[1] ), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1   g0233(.A1(new_n309_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1   g0234(.A1(new_n493_), .A2(new_n497_), .B(new_n278_), .ZN(new_n498_));
  NOR2_X1    g0235(.A1(\a[57] ), .A2(\shift[1] ), .ZN(new_n499_));
  NOR3_X1    g0236(.A1(new_n279_), .A2(\a[54] ), .A3(\shift[1] ), .ZN(new_n500_));
  NOR3_X1    g0237(.A1(new_n279_), .A2(\a[54] ), .A3(\shift[1] ), .ZN(new_n501_));
  NOR3_X1    g0238(.A1(new_n501_), .A2(\shift[0] ), .A3(new_n499_), .ZN(new_n502_));
  NOR2_X1    g0239(.A1(new_n502_), .A2(new_n500_), .ZN(new_n503_));
  NOR2_X1    g0240(.A1(new_n284_), .A2(\a[55] ), .ZN(new_n504_));
  NOR2_X1    g0241(.A1(\a[56] ), .A2(\shift[1] ), .ZN(new_n505_));
  NOR2_X1    g0242(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1   g0243(.A1(new_n506_), .A2(new_n309_), .ZN(new_n507_));
  NOR3_X1    g0244(.A1(new_n503_), .A2(new_n315_), .A3(new_n507_), .ZN(new_n508_));
  NOR2_X1    g0245(.A1(\a[61] ), .A2(\shift[1] ), .ZN(new_n509_));
  NOR3_X1    g0246(.A1(new_n279_), .A2(\a[58] ), .A3(\shift[1] ), .ZN(new_n510_));
  NOR3_X1    g0247(.A1(new_n279_), .A2(\a[58] ), .A3(\shift[1] ), .ZN(new_n511_));
  NOR3_X1    g0248(.A1(new_n511_), .A2(\shift[0] ), .A3(new_n509_), .ZN(new_n512_));
  NOR2_X1    g0249(.A1(new_n512_), .A2(new_n510_), .ZN(new_n513_));
  NOR2_X1    g0250(.A1(new_n284_), .A2(\a[59] ), .ZN(new_n514_));
  NOR2_X1    g0251(.A1(\a[60] ), .A2(\shift[1] ), .ZN(new_n515_));
  NOR2_X1    g0252(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1   g0253(.A1(new_n516_), .A2(new_n309_), .ZN(new_n517_));
  NOR3_X1    g0254(.A1(new_n513_), .A2(new_n315_), .A3(new_n517_), .ZN(new_n518_));
  NOR4_X1    g0255(.A1(new_n488_), .A2(new_n508_), .A3(new_n518_), .A4(new_n498_), .ZN(new_n519_));
  AOI21_X1   g0256(.A1(new_n519_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n520_));
  NOR3_X1    g0257(.A1(new_n279_), .A2(\a[50] ), .A3(\shift[1] ), .ZN(new_n521_));
  NOR3_X1    g0258(.A1(new_n521_), .A2(\shift[0] ), .A3(new_n477_), .ZN(new_n522_));
  NOR2_X1    g0259(.A1(new_n522_), .A2(new_n478_), .ZN(new_n523_));
  NOR2_X1    g0260(.A1(new_n485_), .A2(new_n486_), .ZN(new_n524_));
  NAND2_X1   g0261(.A1(new_n524_), .A2(new_n309_), .ZN(new_n525_));
  OAI21_X1   g0262(.A1(new_n523_), .A2(new_n525_), .B(new_n277_), .ZN(new_n526_));
  INV_X1     g0263(.I(new_n490_), .ZN(new_n527_));
  NOR2_X1    g0264(.A1(new_n489_), .A2(\shift[0] ), .ZN(new_n528_));
  INV_X1     g0265(.I(\a[62] ), .ZN(new_n529_));
  NAND3_X1   g0266(.A1(new_n529_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n530_));
  NAND2_X1   g0267(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1   g0268(.A1(new_n531_), .A2(new_n527_), .ZN(new_n532_));
  AND2_X2    g0269(.A1(new_n309_), .A2(new_n496_), .Z(new_n533_));
  NAND2_X1   g0270(.A1(new_n533_), .A2(new_n532_), .ZN(new_n534_));
  NAND3_X1   g0271(.A1(new_n534_), .A2(new_n526_), .A3(new_n278_), .ZN(new_n535_));
  INV_X1     g0272(.I(new_n500_), .ZN(new_n536_));
  NOR2_X1    g0273(.A1(new_n499_), .A2(\shift[0] ), .ZN(new_n537_));
  INV_X1     g0274(.I(\a[54] ), .ZN(new_n538_));
  NAND3_X1   g0275(.A1(new_n538_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n539_));
  NAND2_X1   g0276(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1   g0277(.A1(new_n540_), .A2(new_n536_), .ZN(new_n541_));
  NOR3_X1    g0278(.A1(new_n283_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n542_));
  NAND2_X1   g0279(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1     g0280(.I(new_n510_), .ZN(new_n544_));
  NOR2_X1    g0281(.A1(new_n509_), .A2(\shift[0] ), .ZN(new_n545_));
  INV_X1     g0282(.I(\a[58] ), .ZN(new_n546_));
  NAND3_X1   g0283(.A1(new_n546_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n547_));
  NAND2_X1   g0284(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1   g0285(.A1(new_n548_), .A2(new_n544_), .ZN(new_n549_));
  NOR3_X1    g0286(.A1(new_n283_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n550_));
  NAND2_X1   g0287(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1   g0288(.A1(new_n543_), .A2(new_n551_), .B(new_n315_), .ZN(new_n552_));
  NOR4_X1    g0289(.A1(new_n535_), .A2(new_n552_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n553_));
  NOR2_X1    g0290(.A1(new_n520_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1     g0291(.I(\a[2] ), .ZN(new_n555_));
  NOR2_X1    g0292(.A1(\a[5] ), .A2(\shift[1] ), .ZN(new_n556_));
  NAND3_X1   g0293(.A1(new_n555_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n557_));
  INV_X1     g0294(.I(new_n557_), .ZN(new_n558_));
  NOR3_X1    g0295(.A1(new_n279_), .A2(\a[2] ), .A3(\shift[1] ), .ZN(new_n559_));
  NOR3_X1    g0296(.A1(new_n559_), .A2(\shift[0] ), .A3(new_n556_), .ZN(new_n560_));
  NOR2_X1    g0297(.A1(new_n560_), .A2(new_n558_), .ZN(new_n561_));
  NOR2_X1    g0298(.A1(new_n284_), .A2(\a[3] ), .ZN(new_n562_));
  NOR2_X1    g0299(.A1(\a[4] ), .A2(\shift[1] ), .ZN(new_n563_));
  NOR2_X1    g0300(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1   g0301(.A1(new_n564_), .A2(new_n309_), .ZN(new_n565_));
  OAI21_X1   g0302(.A1(new_n561_), .A2(new_n565_), .B(new_n277_), .ZN(new_n566_));
  NOR2_X1    g0303(.A1(\a[17] ), .A2(\shift[1] ), .ZN(new_n567_));
  NOR3_X1    g0304(.A1(new_n279_), .A2(\a[14] ), .A3(\shift[1] ), .ZN(new_n568_));
  INV_X1     g0305(.I(new_n568_), .ZN(new_n569_));
  NOR2_X1    g0306(.A1(new_n567_), .A2(\shift[0] ), .ZN(new_n570_));
  INV_X1     g0307(.I(\a[14] ), .ZN(new_n571_));
  NAND3_X1   g0308(.A1(new_n571_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n572_));
  NAND2_X1   g0309(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1   g0310(.A1(new_n573_), .A2(new_n569_), .ZN(new_n574_));
  NOR2_X1    g0311(.A1(new_n284_), .A2(\a[15] ), .ZN(new_n575_));
  NOR2_X1    g0312(.A1(\a[16] ), .A2(\shift[1] ), .ZN(new_n576_));
  NOR3_X1    g0313(.A1(new_n283_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1   g0314(.A1(new_n574_), .A2(new_n577_), .B(new_n315_), .ZN(new_n578_));
  NAND2_X1   g0315(.A1(new_n578_), .A2(new_n566_), .ZN(new_n579_));
  NOR2_X1    g0316(.A1(\a[9] ), .A2(\shift[1] ), .ZN(new_n580_));
  NOR3_X1    g0317(.A1(new_n279_), .A2(\a[6] ), .A3(\shift[1] ), .ZN(new_n581_));
  INV_X1     g0318(.I(new_n581_), .ZN(new_n582_));
  NOR2_X1    g0319(.A1(new_n580_), .A2(\shift[0] ), .ZN(new_n583_));
  INV_X1     g0320(.I(\a[6] ), .ZN(new_n584_));
  NAND3_X1   g0321(.A1(new_n584_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n585_));
  NAND2_X1   g0322(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1   g0323(.A1(new_n586_), .A2(new_n582_), .ZN(new_n587_));
  NOR2_X1    g0324(.A1(new_n284_), .A2(\a[7] ), .ZN(new_n588_));
  NOR2_X1    g0325(.A1(\a[8] ), .A2(\shift[1] ), .ZN(new_n589_));
  NOR3_X1    g0326(.A1(new_n283_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND3_X1   g0327(.A1(new_n587_), .A2(new_n590_), .A3(new_n278_), .ZN(new_n591_));
  NOR2_X1    g0328(.A1(\a[13] ), .A2(\shift[1] ), .ZN(new_n592_));
  NOR3_X1    g0329(.A1(new_n279_), .A2(\a[10] ), .A3(\shift[1] ), .ZN(new_n593_));
  INV_X1     g0330(.I(new_n593_), .ZN(new_n594_));
  NOR2_X1    g0331(.A1(new_n592_), .A2(\shift[0] ), .ZN(new_n595_));
  INV_X1     g0332(.I(\a[10] ), .ZN(new_n596_));
  NAND3_X1   g0333(.A1(new_n596_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n597_));
  NAND2_X1   g0334(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1   g0335(.A1(new_n598_), .A2(new_n594_), .ZN(new_n599_));
  NOR2_X1    g0336(.A1(new_n284_), .A2(\a[11] ), .ZN(new_n600_));
  NOR2_X1    g0337(.A1(\a[12] ), .A2(\shift[1] ), .ZN(new_n601_));
  NOR3_X1    g0338(.A1(new_n283_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1   g0339(.A1(new_n599_), .A2(new_n602_), .A3(new_n278_), .ZN(new_n603_));
  NAND2_X1   g0340(.A1(new_n591_), .A2(new_n603_), .ZN(new_n604_));
  NOR4_X1    g0341(.A1(new_n579_), .A2(new_n604_), .A3(new_n270_), .A4(\shift[5] ), .ZN(new_n605_));
  NOR2_X1    g0342(.A1(new_n556_), .A2(\shift[0] ), .ZN(new_n606_));
  NAND3_X1   g0343(.A1(new_n555_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n607_));
  NAND2_X1   g0344(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1   g0345(.A1(new_n608_), .A2(new_n557_), .ZN(new_n609_));
  NOR3_X1    g0346(.A1(new_n283_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n610_));
  AOI21_X1   g0347(.A1(new_n609_), .A2(new_n610_), .B(new_n291_), .ZN(new_n611_));
  NOR3_X1    g0348(.A1(new_n279_), .A2(\a[14] ), .A3(\shift[1] ), .ZN(new_n612_));
  NOR3_X1    g0349(.A1(new_n612_), .A2(\shift[0] ), .A3(new_n567_), .ZN(new_n613_));
  NOR2_X1    g0350(.A1(new_n613_), .A2(new_n568_), .ZN(new_n614_));
  NOR2_X1    g0351(.A1(new_n575_), .A2(new_n576_), .ZN(new_n615_));
  NAND2_X1   g0352(.A1(new_n615_), .A2(new_n309_), .ZN(new_n616_));
  OAI21_X1   g0353(.A1(new_n614_), .A2(new_n616_), .B(new_n278_), .ZN(new_n617_));
  NOR3_X1    g0354(.A1(new_n279_), .A2(\a[6] ), .A3(\shift[1] ), .ZN(new_n618_));
  NOR3_X1    g0355(.A1(new_n618_), .A2(\shift[0] ), .A3(new_n580_), .ZN(new_n619_));
  NOR2_X1    g0356(.A1(new_n619_), .A2(new_n581_), .ZN(new_n620_));
  NOR2_X1    g0357(.A1(new_n588_), .A2(new_n589_), .ZN(new_n621_));
  NAND2_X1   g0358(.A1(new_n621_), .A2(new_n309_), .ZN(new_n622_));
  NOR3_X1    g0359(.A1(new_n620_), .A2(new_n315_), .A3(new_n622_), .ZN(new_n623_));
  NOR3_X1    g0360(.A1(new_n279_), .A2(\a[10] ), .A3(\shift[1] ), .ZN(new_n624_));
  NOR3_X1    g0361(.A1(new_n624_), .A2(\shift[0] ), .A3(new_n592_), .ZN(new_n625_));
  NOR2_X1    g0362(.A1(new_n625_), .A2(new_n593_), .ZN(new_n626_));
  NOR2_X1    g0363(.A1(new_n600_), .A2(new_n601_), .ZN(new_n627_));
  NAND2_X1   g0364(.A1(new_n627_), .A2(new_n309_), .ZN(new_n628_));
  NOR3_X1    g0365(.A1(new_n626_), .A2(new_n315_), .A3(new_n628_), .ZN(new_n629_));
  NOR4_X1    g0366(.A1(new_n611_), .A2(new_n623_), .A3(new_n629_), .A4(new_n617_), .ZN(new_n630_));
  AOI21_X1   g0367(.A1(new_n630_), .A2(\shift[4] ), .B(new_n265_), .ZN(new_n631_));
  NOR2_X1    g0368(.A1(new_n631_), .A2(new_n605_), .ZN(new_n632_));
  NOR2_X1    g0369(.A1(\a[21] ), .A2(\shift[1] ), .ZN(new_n633_));
  NOR2_X1    g0370(.A1(new_n633_), .A2(\shift[0] ), .ZN(new_n634_));
  NOR3_X1    g0371(.A1(new_n279_), .A2(\a[18] ), .A3(\shift[1] ), .ZN(new_n635_));
  XOR2_X1    g0372(.A1(new_n634_), .A2(new_n635_), .Z(new_n636_));
  INV_X1     g0373(.I(\a[19] ), .ZN(new_n637_));
  NOR2_X1    g0374(.A1(\a[20] ), .A2(\shift[1] ), .ZN(new_n638_));
  AOI21_X1   g0375(.A1(new_n637_), .A2(\shift[1] ), .B(new_n638_), .ZN(new_n639_));
  AND2_X2    g0376(.A1(new_n309_), .A2(new_n639_), .Z(new_n640_));
  AOI21_X1   g0377(.A1(new_n636_), .A2(new_n640_), .B(new_n291_), .ZN(new_n641_));
  NOR2_X1    g0378(.A1(\a[33] ), .A2(\shift[1] ), .ZN(new_n642_));
  NOR2_X1    g0379(.A1(new_n642_), .A2(\shift[0] ), .ZN(new_n643_));
  INV_X1     g0380(.I(\a[30] ), .ZN(new_n644_));
  NAND3_X1   g0381(.A1(new_n644_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n645_));
  NOR2_X1    g0382(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1   g0383(.A1(\a[33] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n647_));
  NOR3_X1    g0384(.A1(new_n279_), .A2(\a[30] ), .A3(\shift[1] ), .ZN(new_n648_));
  NOR2_X1    g0385(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1    g0386(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1    g0387(.A1(new_n284_), .A2(\a[31] ), .ZN(new_n651_));
  NOR2_X1    g0388(.A1(\a[32] ), .A2(\shift[1] ), .ZN(new_n652_));
  NOR2_X1    g0389(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1   g0390(.A1(new_n653_), .A2(new_n309_), .ZN(new_n654_));
  OAI21_X1   g0391(.A1(new_n650_), .A2(new_n654_), .B(new_n278_), .ZN(new_n655_));
  NOR2_X1    g0392(.A1(\a[25] ), .A2(\shift[1] ), .ZN(new_n656_));
  NOR3_X1    g0393(.A1(new_n279_), .A2(\a[22] ), .A3(\shift[1] ), .ZN(new_n657_));
  NOR3_X1    g0394(.A1(new_n279_), .A2(\a[22] ), .A3(\shift[1] ), .ZN(new_n658_));
  NOR3_X1    g0395(.A1(new_n658_), .A2(\shift[0] ), .A3(new_n656_), .ZN(new_n659_));
  NOR2_X1    g0396(.A1(new_n659_), .A2(new_n657_), .ZN(new_n660_));
  INV_X1     g0397(.I(\a[23] ), .ZN(new_n661_));
  NAND2_X1   g0398(.A1(new_n661_), .A2(\shift[1] ), .ZN(new_n662_));
  OR2_X2     g0399(.A1(\a[24] ), .A2(\shift[1] ), .Z(new_n663_));
  NAND3_X1   g0400(.A1(new_n309_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NOR3_X1    g0401(.A1(new_n660_), .A2(new_n315_), .A3(new_n664_), .ZN(new_n665_));
  NOR2_X1    g0402(.A1(\a[29] ), .A2(\shift[1] ), .ZN(new_n666_));
  NOR3_X1    g0403(.A1(new_n279_), .A2(\a[26] ), .A3(\shift[1] ), .ZN(new_n667_));
  NOR3_X1    g0404(.A1(new_n279_), .A2(\a[26] ), .A3(\shift[1] ), .ZN(new_n668_));
  NOR3_X1    g0405(.A1(new_n668_), .A2(\shift[0] ), .A3(new_n666_), .ZN(new_n669_));
  NOR2_X1    g0406(.A1(new_n669_), .A2(new_n667_), .ZN(new_n670_));
  NOR2_X1    g0407(.A1(new_n284_), .A2(\a[27] ), .ZN(new_n671_));
  NOR2_X1    g0408(.A1(\a[28] ), .A2(\shift[1] ), .ZN(new_n672_));
  NOR2_X1    g0409(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1   g0410(.A1(new_n673_), .A2(new_n309_), .ZN(new_n674_));
  NOR3_X1    g0411(.A1(new_n670_), .A2(new_n315_), .A3(new_n674_), .ZN(new_n675_));
  OR4_X2     g0412(.A1(new_n641_), .A2(new_n655_), .A3(new_n665_), .A4(new_n675_), .Z(new_n676_));
  NOR2_X1    g0413(.A1(new_n265_), .A2(\shift[4] ), .ZN(new_n677_));
  NOR2_X1    g0414(.A1(new_n270_), .A2(\shift[5] ), .ZN(new_n678_));
  NOR2_X1    g0415(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1     g0416(.I(new_n679_), .ZN(new_n680_));
  NOR2_X1    g0417(.A1(\a[37] ), .A2(\shift[1] ), .ZN(new_n681_));
  NOR3_X1    g0418(.A1(new_n279_), .A2(\a[34] ), .A3(\shift[1] ), .ZN(new_n682_));
  INV_X1     g0419(.I(new_n682_), .ZN(new_n683_));
  NOR2_X1    g0420(.A1(new_n681_), .A2(\shift[0] ), .ZN(new_n684_));
  INV_X1     g0421(.I(\a[34] ), .ZN(new_n685_));
  NAND3_X1   g0422(.A1(new_n685_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n686_));
  NAND2_X1   g0423(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1   g0424(.A1(new_n687_), .A2(new_n683_), .ZN(new_n688_));
  NOR2_X1    g0425(.A1(new_n284_), .A2(\a[35] ), .ZN(new_n689_));
  NOR2_X1    g0426(.A1(\a[36] ), .A2(\shift[1] ), .ZN(new_n690_));
  NOR3_X1    g0427(.A1(new_n283_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1   g0428(.A1(new_n688_), .A2(new_n691_), .B(new_n291_), .ZN(new_n692_));
  NOR2_X1    g0429(.A1(\a[49] ), .A2(\shift[1] ), .ZN(new_n693_));
  NOR3_X1    g0430(.A1(new_n279_), .A2(\a[46] ), .A3(\shift[1] ), .ZN(new_n694_));
  NOR3_X1    g0431(.A1(new_n279_), .A2(\a[46] ), .A3(\shift[1] ), .ZN(new_n695_));
  NOR3_X1    g0432(.A1(new_n695_), .A2(\shift[0] ), .A3(new_n693_), .ZN(new_n696_));
  NOR2_X1    g0433(.A1(new_n696_), .A2(new_n694_), .ZN(new_n697_));
  NOR2_X1    g0434(.A1(new_n284_), .A2(\a[47] ), .ZN(new_n698_));
  NOR2_X1    g0435(.A1(\a[48] ), .A2(\shift[1] ), .ZN(new_n699_));
  NOR2_X1    g0436(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1   g0437(.A1(new_n700_), .A2(new_n309_), .ZN(new_n701_));
  OAI21_X1   g0438(.A1(new_n697_), .A2(new_n701_), .B(new_n440_), .ZN(new_n702_));
  NOR2_X1    g0439(.A1(new_n692_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1    g0440(.A1(new_n703_), .A2(new_n680_), .ZN(new_n704_));
  OAI21_X1   g0441(.A1(new_n676_), .A2(\shift[4] ), .B(new_n704_), .ZN(new_n705_));
  AOI21_X1   g0442(.A1(new_n554_), .A2(new_n632_), .B(new_n705_), .ZN(new_n706_));
  OAI21_X1   g0443(.A1(new_n706_), .A2(new_n264_), .B(new_n476_), .ZN(\result[1] ));
  NAND2_X1   g0444(.A1(new_n270_), .A2(new_n265_), .ZN(new_n708_));
  NOR2_X1    g0445(.A1(new_n441_), .A2(new_n277_), .ZN(new_n709_));
  INV_X1     g0446(.I(new_n709_), .ZN(new_n710_));
  NAND4_X1   g0447(.A1(new_n710_), .A2(new_n265_), .A3(new_n708_), .A4(new_n273_), .ZN(new_n711_));
  NAND2_X1   g0448(.A1(new_n711_), .A2(new_n264_), .ZN(new_n712_));
  XOR2_X1    g0449(.A1(new_n273_), .A2(\shift[5] ), .Z(new_n713_));
  NOR2_X1    g0450(.A1(new_n272_), .A2(\shift[5] ), .ZN(new_n714_));
  NOR2_X1    g0451(.A1(new_n271_), .A2(new_n265_), .ZN(new_n715_));
  NOR3_X1    g0452(.A1(new_n714_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1   g0453(.A1(new_n710_), .A2(new_n273_), .A3(new_n679_), .ZN(new_n717_));
  NOR2_X1    g0454(.A1(new_n717_), .A2(new_n716_), .ZN(new_n718_));
  OAI21_X1   g0455(.A1(new_n718_), .A2(new_n264_), .B(new_n712_), .ZN(\result[2] ));
  NAND2_X1   g0456(.A1(new_n344_), .A2(\shift[0] ), .ZN(new_n721_));
  OAI21_X1   g0457(.A1(\a[119] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n722_));
  NAND2_X1   g0458(.A1(new_n722_), .A2(new_n721_), .ZN(new_n723_));
  INV_X1     g0459(.I(\a[117] ), .ZN(new_n724_));
  NAND2_X1   g0460(.A1(new_n724_), .A2(\shift[1] ), .ZN(new_n725_));
  OR2_X2     g0461(.A1(\a[118] ), .A2(\shift[1] ), .Z(new_n726_));
  NAND3_X1   g0462(.A1(new_n309_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1     g0463(.I(new_n727_), .ZN(new_n728_));
  AOI21_X1   g0464(.A1(new_n728_), .A2(new_n723_), .B(new_n291_), .ZN(new_n729_));
  OAI21_X1   g0465(.A1(\a[3] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n730_));
  NOR3_X1    g0466(.A1(new_n279_), .A2(\a[0] ), .A3(\shift[1] ), .ZN(new_n731_));
  XOR2_X1    g0467(.A1(new_n730_), .A2(new_n731_), .Z(new_n732_));
  NAND2_X1   g0468(.A1(new_n352_), .A2(\shift[1] ), .ZN(new_n733_));
  NAND2_X1   g0469(.A1(new_n555_), .A2(new_n284_), .ZN(new_n734_));
  NAND3_X1   g0470(.A1(new_n309_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NOR2_X1    g0471(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1   g0472(.A1(new_n364_), .A2(\shift[0] ), .ZN(new_n738_));
  OAI21_X1   g0473(.A1(\a[123] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n739_));
  NAND2_X1   g0474(.A1(new_n739_), .A2(new_n738_), .ZN(new_n740_));
  INV_X1     g0475(.I(\a[121] ), .ZN(new_n741_));
  NAND2_X1   g0476(.A1(new_n741_), .A2(\shift[1] ), .ZN(new_n742_));
  NAND2_X1   g0477(.A1(new_n371_), .A2(new_n284_), .ZN(new_n743_));
  AND2_X2    g0478(.A1(new_n743_), .A2(new_n742_), .Z(new_n744_));
  NAND4_X1   g0479(.A1(new_n744_), .A2(new_n278_), .A3(new_n740_), .A4(new_n309_), .ZN(new_n745_));
  NAND2_X1   g0480(.A1(new_n376_), .A2(\shift[0] ), .ZN(new_n747_));
  OAI21_X1   g0481(.A1(\a[127] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n748_));
  NAND2_X1   g0482(.A1(new_n748_), .A2(new_n747_), .ZN(new_n749_));
  NOR2_X1    g0483(.A1(new_n284_), .A2(\a[125] ), .ZN(new_n750_));
  NOR2_X1    g0484(.A1(\a[126] ), .A2(\shift[1] ), .ZN(new_n751_));
  NOR2_X1    g0485(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1   g0486(.A1(new_n749_), .A2(new_n278_), .A3(new_n309_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1   g0487(.A1(new_n745_), .A2(new_n753_), .ZN(new_n754_));
  NOR4_X1    g0488(.A1(new_n754_), .A2(new_n729_), .A3(new_n736_), .A4(new_n315_), .ZN(new_n755_));
  AOI21_X1   g0489(.A1(new_n755_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n756_));
  INV_X1     g0490(.I(new_n723_), .ZN(new_n757_));
  OAI21_X1   g0491(.A1(new_n757_), .A2(new_n727_), .B(new_n277_), .ZN(new_n758_));
  NOR2_X1    g0492(.A1(\a[3] ), .A2(\shift[1] ), .ZN(new_n759_));
  NOR2_X1    g0493(.A1(new_n759_), .A2(\shift[0] ), .ZN(new_n760_));
  XOR2_X1    g0494(.A1(new_n760_), .A2(new_n731_), .Z(new_n761_));
  NAND2_X1   g0495(.A1(new_n734_), .A2(new_n733_), .ZN(new_n762_));
  NOR2_X1    g0496(.A1(new_n762_), .A2(new_n283_), .ZN(new_n763_));
  AOI21_X1   g0497(.A1(new_n761_), .A2(new_n763_), .B(new_n315_), .ZN(new_n764_));
  NAND4_X1   g0498(.A1(new_n764_), .A2(new_n758_), .A3(new_n745_), .A4(new_n753_), .ZN(new_n765_));
  NOR3_X1    g0499(.A1(new_n765_), .A2(\shift[4] ), .A3(new_n265_), .ZN(new_n766_));
  NOR2_X1    g0500(.A1(new_n756_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1   g0501(.A1(new_n436_), .A2(\shift[0] ), .ZN(new_n769_));
  OAI21_X1   g0502(.A1(\a[71] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n770_));
  NAND2_X1   g0503(.A1(new_n770_), .A2(new_n769_), .ZN(new_n771_));
  INV_X1     g0504(.I(new_n771_), .ZN(new_n772_));
  INV_X1     g0505(.I(\a[69] ), .ZN(new_n773_));
  NAND2_X1   g0506(.A1(new_n773_), .A2(\shift[1] ), .ZN(new_n774_));
  OR2_X2     g0507(.A1(\a[70] ), .A2(\shift[1] ), .Z(new_n775_));
  NAND3_X1   g0508(.A1(new_n309_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1   g0509(.A1(new_n772_), .A2(new_n776_), .B(new_n277_), .ZN(new_n777_));
  NAND2_X1   g0510(.A1(new_n448_), .A2(\shift[0] ), .ZN(new_n779_));
  OAI21_X1   g0511(.A1(\a[83] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n780_));
  NAND2_X1   g0512(.A1(new_n780_), .A2(new_n779_), .ZN(new_n781_));
  INV_X1     g0513(.I(\a[81] ), .ZN(new_n782_));
  NAND2_X1   g0514(.A1(new_n782_), .A2(\shift[1] ), .ZN(new_n783_));
  OAI21_X1   g0515(.A1(\a[82] ), .A2(\shift[1] ), .B(new_n783_), .ZN(new_n784_));
  NOR2_X1    g0516(.A1(new_n784_), .A2(new_n283_), .ZN(new_n785_));
  NAND2_X1   g0517(.A1(new_n785_), .A2(new_n781_), .ZN(new_n786_));
  NAND3_X1   g0518(.A1(new_n777_), .A2(new_n786_), .A3(new_n278_), .ZN(new_n787_));
  NAND2_X1   g0519(.A1(new_n458_), .A2(\shift[0] ), .ZN(new_n789_));
  OAI21_X1   g0520(.A1(\a[75] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n790_));
  NAND2_X1   g0521(.A1(new_n790_), .A2(new_n789_), .ZN(new_n791_));
  INV_X1     g0522(.I(\a[73] ), .ZN(new_n792_));
  NAND2_X1   g0523(.A1(new_n792_), .A2(\shift[1] ), .ZN(new_n793_));
  NAND2_X1   g0524(.A1(new_n466_), .A2(new_n284_), .ZN(new_n794_));
  NAND3_X1   g0525(.A1(new_n309_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1     g0526(.I(new_n795_), .ZN(new_n796_));
  NAND3_X1   g0527(.A1(new_n796_), .A2(new_n791_), .A3(new_n278_), .ZN(new_n797_));
  NAND2_X1   g0528(.A1(new_n471_), .A2(\shift[0] ), .ZN(new_n799_));
  OAI21_X1   g0529(.A1(\a[79] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n800_));
  NAND2_X1   g0530(.A1(new_n800_), .A2(new_n799_), .ZN(new_n801_));
  INV_X1     g0531(.I(\a[77] ), .ZN(new_n802_));
  NAND2_X1   g0532(.A1(new_n802_), .A2(\shift[1] ), .ZN(new_n803_));
  OAI21_X1   g0533(.A1(\a[78] ), .A2(\shift[1] ), .B(new_n803_), .ZN(new_n804_));
  NOR2_X1    g0534(.A1(new_n804_), .A2(new_n283_), .ZN(new_n805_));
  NAND3_X1   g0535(.A1(new_n805_), .A2(new_n278_), .A3(new_n801_), .ZN(new_n806_));
  NAND2_X1   g0536(.A1(new_n797_), .A2(new_n806_), .ZN(new_n807_));
  NOR4_X1    g0537(.A1(new_n807_), .A2(new_n787_), .A3(new_n270_), .A4(\shift[5] ), .ZN(new_n808_));
  INV_X1     g0538(.I(new_n776_), .ZN(new_n809_));
  AOI21_X1   g0539(.A1(new_n809_), .A2(new_n771_), .B(new_n291_), .ZN(new_n810_));
  INV_X1     g0540(.I(new_n781_), .ZN(new_n811_));
  NAND2_X1   g0541(.A1(new_n386_), .A2(new_n284_), .ZN(new_n812_));
  NAND3_X1   g0542(.A1(new_n309_), .A2(new_n783_), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1   g0543(.A1(new_n811_), .A2(new_n813_), .B(new_n278_), .ZN(new_n814_));
  INV_X1     g0544(.I(new_n791_), .ZN(new_n815_));
  NOR3_X1    g0545(.A1(new_n815_), .A2(new_n795_), .A3(new_n315_), .ZN(new_n816_));
  INV_X1     g0546(.I(new_n801_), .ZN(new_n817_));
  INV_X1     g0547(.I(\a[78] ), .ZN(new_n818_));
  NAND2_X1   g0548(.A1(new_n818_), .A2(new_n284_), .ZN(new_n819_));
  NAND3_X1   g0549(.A1(new_n309_), .A2(new_n803_), .A3(new_n819_), .ZN(new_n820_));
  NOR3_X1    g0550(.A1(new_n817_), .A2(new_n820_), .A3(new_n315_), .ZN(new_n821_));
  NOR4_X1    g0551(.A1(new_n810_), .A2(new_n814_), .A3(new_n816_), .A4(new_n821_), .ZN(new_n822_));
  AOI21_X1   g0552(.A1(new_n822_), .A2(\shift[4] ), .B(new_n265_), .ZN(new_n823_));
  NOR2_X1    g0553(.A1(new_n823_), .A2(new_n808_), .ZN(new_n824_));
  INV_X1     g0554(.I(\a[87] ), .ZN(new_n825_));
  NOR3_X1    g0555(.A1(new_n279_), .A2(\a[84] ), .A3(\shift[1] ), .ZN(new_n828_));
  AOI21_X1   g0556(.A1(new_n825_), .A2(new_n284_), .B(\shift[0] ), .ZN(new_n829_));
  NOR2_X1    g0557(.A1(new_n829_), .A2(new_n828_), .ZN(new_n830_));
  INV_X1     g0558(.I(\a[85] ), .ZN(new_n831_));
  NAND2_X1   g0559(.A1(new_n831_), .A2(\shift[1] ), .ZN(new_n832_));
  OAI21_X1   g0560(.A1(\a[86] ), .A2(\shift[1] ), .B(new_n832_), .ZN(new_n833_));
  NOR3_X1    g0561(.A1(new_n833_), .A2(new_n830_), .A3(new_n283_), .ZN(new_n834_));
  NOR2_X1    g0562(.A1(new_n834_), .A2(new_n291_), .ZN(new_n835_));
  NAND2_X1   g0563(.A1(new_n400_), .A2(\shift[0] ), .ZN(new_n837_));
  OAI21_X1   g0564(.A1(\a[99] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n838_));
  AND2_X2    g0565(.A1(new_n838_), .A2(new_n837_), .Z(new_n839_));
  MUX2_X1    g0566(.I0(\a[98] ), .I1(\a[97] ), .S(\shift[1] ), .Z(new_n840_));
  NAND2_X1   g0567(.A1(new_n309_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1   g0568(.A1(new_n839_), .A2(new_n841_), .B(new_n278_), .ZN(new_n842_));
  NAND2_X1   g0569(.A1(new_n414_), .A2(\shift[0] ), .ZN(new_n844_));
  OAI21_X1   g0570(.A1(\a[91] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n845_));
  NAND2_X1   g0571(.A1(new_n845_), .A2(new_n844_), .ZN(new_n846_));
  MUX2_X1    g0572(.I0(\a[90] ), .I1(\a[89] ), .S(\shift[1] ), .Z(new_n847_));
  NAND4_X1   g0573(.A1(new_n846_), .A2(new_n278_), .A3(new_n309_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1   g0574(.A1(new_n426_), .A2(\shift[0] ), .ZN(new_n850_));
  OAI21_X1   g0575(.A1(\a[95] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n851_));
  NAND2_X1   g0576(.A1(new_n851_), .A2(new_n850_), .ZN(new_n852_));
  MUX2_X1    g0577(.I0(\a[94] ), .I1(\a[93] ), .S(\shift[1] ), .Z(new_n853_));
  NAND4_X1   g0578(.A1(new_n852_), .A2(new_n278_), .A3(new_n309_), .A4(new_n853_), .ZN(new_n854_));
  NAND2_X1   g0579(.A1(new_n848_), .A2(new_n854_), .ZN(new_n855_));
  NOR3_X1    g0580(.A1(new_n855_), .A2(new_n835_), .A3(new_n842_), .ZN(new_n856_));
  NAND2_X1   g0581(.A1(new_n856_), .A2(new_n270_), .ZN(new_n857_));
  NAND2_X1   g0582(.A1(new_n301_), .A2(\shift[0] ), .ZN(new_n859_));
  OAI21_X1   g0583(.A1(\a[103] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n860_));
  AND2_X2    g0584(.A1(new_n860_), .A2(new_n859_), .Z(new_n861_));
  INV_X1     g0585(.I(\a[101] ), .ZN(new_n862_));
  NOR2_X1    g0586(.A1(\a[102] ), .A2(\shift[1] ), .ZN(new_n863_));
  AOI21_X1   g0587(.A1(new_n862_), .A2(\shift[1] ), .B(new_n863_), .ZN(new_n864_));
  NAND2_X1   g0588(.A1(new_n309_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1   g0589(.A1(new_n861_), .A2(new_n865_), .B(new_n277_), .ZN(new_n866_));
  NAND2_X1   g0590(.A1(new_n311_), .A2(\shift[0] ), .ZN(new_n868_));
  OAI21_X1   g0591(.A1(\a[115] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n869_));
  NAND2_X1   g0592(.A1(new_n869_), .A2(new_n868_), .ZN(new_n870_));
  INV_X1     g0593(.I(\a[113] ), .ZN(new_n871_));
  NAND2_X1   g0594(.A1(new_n871_), .A2(\shift[1] ), .ZN(new_n872_));
  INV_X1     g0595(.I(\a[114] ), .ZN(new_n873_));
  NAND2_X1   g0596(.A1(new_n873_), .A2(new_n284_), .ZN(new_n874_));
  NAND4_X1   g0597(.A1(new_n870_), .A2(new_n309_), .A3(new_n872_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1   g0598(.A1(new_n875_), .A2(new_n278_), .ZN(new_n876_));
  INV_X1     g0599(.I(new_n876_), .ZN(new_n877_));
  NAND2_X1   g0600(.A1(new_n322_), .A2(\shift[0] ), .ZN(new_n879_));
  OAI21_X1   g0601(.A1(\a[107] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n880_));
  AND2_X2    g0602(.A1(new_n880_), .A2(new_n879_), .Z(new_n881_));
  INV_X1     g0603(.I(\a[105] ), .ZN(new_n882_));
  NOR2_X1    g0604(.A1(\a[106] ), .A2(\shift[1] ), .ZN(new_n883_));
  AOI21_X1   g0605(.A1(new_n882_), .A2(\shift[1] ), .B(new_n883_), .ZN(new_n884_));
  NAND2_X1   g0606(.A1(new_n309_), .A2(new_n884_), .ZN(new_n885_));
  NOR3_X1    g0607(.A1(new_n881_), .A2(new_n885_), .A3(new_n315_), .ZN(new_n886_));
  NAND2_X1   g0608(.A1(new_n332_), .A2(\shift[0] ), .ZN(new_n888_));
  OAI21_X1   g0609(.A1(\a[111] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n889_));
  AND2_X2    g0610(.A1(new_n889_), .A2(new_n888_), .Z(new_n890_));
  INV_X1     g0611(.I(\a[109] ), .ZN(new_n891_));
  NAND2_X1   g0612(.A1(new_n891_), .A2(\shift[1] ), .ZN(new_n892_));
  INV_X1     g0613(.I(\a[110] ), .ZN(new_n893_));
  NAND2_X1   g0614(.A1(new_n893_), .A2(new_n284_), .ZN(new_n894_));
  NAND3_X1   g0615(.A1(new_n309_), .A2(new_n892_), .A3(new_n894_), .ZN(new_n895_));
  NOR3_X1    g0616(.A1(new_n890_), .A2(new_n895_), .A3(new_n315_), .ZN(new_n896_));
  NOR2_X1    g0617(.A1(new_n886_), .A2(new_n896_), .ZN(new_n897_));
  NAND4_X1   g0618(.A1(new_n877_), .A2(new_n897_), .A3(\shift[4] ), .A4(new_n866_), .ZN(new_n898_));
  NAND3_X1   g0619(.A1(new_n857_), .A2(new_n898_), .A3(new_n679_), .ZN(new_n899_));
  AOI21_X1   g0620(.A1(new_n767_), .A2(new_n824_), .B(new_n899_), .ZN(new_n900_));
  OAI21_X1   g0621(.A1(\a[43] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n901_));
  NOR3_X1    g0622(.A1(new_n279_), .A2(\a[40] ), .A3(\shift[1] ), .ZN(new_n902_));
  XOR2_X1    g0623(.A1(new_n901_), .A2(new_n902_), .Z(new_n903_));
  INV_X1     g0624(.I(\a[41] ), .ZN(new_n904_));
  NAND2_X1   g0625(.A1(new_n904_), .A2(\shift[1] ), .ZN(new_n905_));
  OR2_X2     g0626(.A1(\a[42] ), .A2(\shift[1] ), .Z(new_n906_));
  NAND3_X1   g0627(.A1(new_n309_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  NOR3_X1    g0628(.A1(new_n903_), .A2(new_n315_), .A3(new_n907_), .ZN(new_n908_));
  NOR3_X1    g0629(.A1(new_n279_), .A2(\a[36] ), .A3(\shift[1] ), .ZN(new_n909_));
  NOR2_X1    g0630(.A1(new_n286_), .A2(\shift[0] ), .ZN(new_n910_));
  NOR2_X1    g0631(.A1(new_n910_), .A2(new_n909_), .ZN(new_n911_));
  NOR2_X1    g0632(.A1(new_n284_), .A2(\a[37] ), .ZN(new_n912_));
  NOR2_X1    g0633(.A1(\a[38] ), .A2(\shift[1] ), .ZN(new_n913_));
  NOR4_X1    g0634(.A1(new_n911_), .A2(new_n283_), .A3(new_n912_), .A4(new_n913_), .ZN(new_n914_));
  NOR2_X1    g0635(.A1(new_n914_), .A2(new_n291_), .ZN(new_n915_));
  NAND2_X1   g0636(.A1(new_n699_), .A2(\shift[0] ), .ZN(new_n917_));
  OAI21_X1   g0637(.A1(\a[51] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n918_));
  NAND2_X1   g0638(.A1(new_n918_), .A2(new_n917_), .ZN(new_n919_));
  INV_X1     g0639(.I(new_n919_), .ZN(new_n920_));
  NOR2_X1    g0640(.A1(new_n284_), .A2(\a[49] ), .ZN(new_n921_));
  NOR2_X1    g0641(.A1(\a[50] ), .A2(\shift[1] ), .ZN(new_n922_));
  NOR2_X1    g0642(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1   g0643(.A1(new_n923_), .A2(new_n309_), .ZN(new_n924_));
  OAI21_X1   g0644(.A1(new_n920_), .A2(new_n924_), .B(new_n278_), .ZN(new_n925_));
  NOR3_X1    g0645(.A1(new_n908_), .A2(new_n915_), .A3(new_n925_), .ZN(new_n926_));
  NOR2_X1    g0646(.A1(new_n926_), .A2(new_n270_), .ZN(new_n927_));
  NAND2_X1   g0647(.A1(new_n486_), .A2(\shift[0] ), .ZN(new_n929_));
  OAI21_X1   g0648(.A1(\a[55] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n930_));
  NAND2_X1   g0649(.A1(new_n930_), .A2(new_n929_), .ZN(new_n931_));
  INV_X1     g0650(.I(new_n931_), .ZN(new_n932_));
  INV_X1     g0651(.I(\a[53] ), .ZN(new_n933_));
  NOR2_X1    g0652(.A1(\a[54] ), .A2(\shift[1] ), .ZN(new_n934_));
  AOI21_X1   g0653(.A1(new_n933_), .A2(\shift[1] ), .B(new_n934_), .ZN(new_n935_));
  NAND2_X1   g0654(.A1(new_n309_), .A2(new_n935_), .ZN(new_n936_));
  OAI21_X1   g0655(.A1(new_n932_), .A2(new_n936_), .B(new_n277_), .ZN(new_n937_));
  NAND2_X1   g0656(.A1(new_n495_), .A2(\shift[0] ), .ZN(new_n939_));
  OAI21_X1   g0657(.A1(\a[67] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n940_));
  NAND2_X1   g0658(.A1(new_n940_), .A2(new_n939_), .ZN(new_n941_));
  MUX2_X1    g0659(.I0(\a[66] ), .I1(\a[65] ), .S(\shift[1] ), .Z(new_n942_));
  NAND3_X1   g0660(.A1(new_n941_), .A2(new_n309_), .A3(new_n942_), .ZN(new_n943_));
  NAND3_X1   g0661(.A1(new_n937_), .A2(new_n943_), .A3(new_n278_), .ZN(new_n944_));
  NAND2_X1   g0662(.A1(new_n505_), .A2(\shift[0] ), .ZN(new_n946_));
  OAI21_X1   g0663(.A1(\a[59] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n947_));
  NAND2_X1   g0664(.A1(new_n947_), .A2(new_n946_), .ZN(new_n948_));
  MUX2_X1    g0665(.I0(\a[58] ), .I1(\a[57] ), .S(\shift[1] ), .Z(new_n949_));
  NAND4_X1   g0666(.A1(new_n948_), .A2(new_n278_), .A3(new_n309_), .A4(new_n949_), .ZN(new_n950_));
  NAND2_X1   g0667(.A1(new_n515_), .A2(\shift[0] ), .ZN(new_n952_));
  OAI21_X1   g0668(.A1(\a[63] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n953_));
  NAND2_X1   g0669(.A1(new_n953_), .A2(new_n952_), .ZN(new_n954_));
  INV_X1     g0670(.I(\a[61] ), .ZN(new_n955_));
  NAND2_X1   g0671(.A1(new_n955_), .A2(\shift[1] ), .ZN(new_n956_));
  NAND2_X1   g0672(.A1(new_n529_), .A2(new_n284_), .ZN(new_n957_));
  NAND2_X1   g0673(.A1(new_n957_), .A2(new_n956_), .ZN(new_n958_));
  NOR2_X1    g0674(.A1(new_n958_), .A2(new_n283_), .ZN(new_n959_));
  NAND2_X1   g0675(.A1(new_n959_), .A2(new_n954_), .ZN(new_n960_));
  OAI21_X1   g0676(.A1(new_n960_), .A2(new_n315_), .B(new_n950_), .ZN(new_n961_));
  NOR3_X1    g0677(.A1(new_n944_), .A2(new_n270_), .A3(new_n961_), .ZN(new_n962_));
  NOR3_X1    g0678(.A1(new_n927_), .A2(new_n962_), .A3(\shift[5] ), .ZN(new_n963_));
  NAND2_X1   g0679(.A1(new_n638_), .A2(\shift[0] ), .ZN(new_n965_));
  OAI21_X1   g0680(.A1(\a[23] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n966_));
  NAND2_X1   g0681(.A1(new_n966_), .A2(new_n965_), .ZN(new_n967_));
  INV_X1     g0682(.I(\a[21] ), .ZN(new_n968_));
  NAND2_X1   g0683(.A1(new_n968_), .A2(\shift[1] ), .ZN(new_n969_));
  OR2_X2     g0684(.A1(\a[22] ), .A2(\shift[1] ), .Z(new_n970_));
  NAND2_X1   g0685(.A1(new_n970_), .A2(new_n969_), .ZN(new_n971_));
  NOR2_X1    g0686(.A1(new_n971_), .A2(new_n283_), .ZN(new_n972_));
  AOI21_X1   g0687(.A1(new_n972_), .A2(new_n967_), .B(new_n291_), .ZN(new_n973_));
  NAND2_X1   g0688(.A1(new_n652_), .A2(\shift[0] ), .ZN(new_n975_));
  OAI21_X1   g0689(.A1(\a[35] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n976_));
  NAND2_X1   g0690(.A1(new_n976_), .A2(new_n975_), .ZN(new_n977_));
  NOR2_X1    g0691(.A1(new_n284_), .A2(\a[33] ), .ZN(new_n978_));
  NOR2_X1    g0692(.A1(\a[34] ), .A2(\shift[1] ), .ZN(new_n979_));
  NOR2_X1    g0693(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  NAND3_X1   g0694(.A1(new_n977_), .A2(new_n309_), .A3(new_n980_), .ZN(new_n981_));
  NAND2_X1   g0695(.A1(new_n981_), .A2(new_n278_), .ZN(new_n982_));
  NOR2_X1    g0696(.A1(\a[27] ), .A2(\shift[1] ), .ZN(new_n983_));
  MUX2_X1    g0697(.I0(new_n983_), .I1(new_n663_), .S(\shift[0] ), .Z(new_n984_));
  INV_X1     g0698(.I(\a[25] ), .ZN(new_n985_));
  NAND2_X1   g0699(.A1(new_n985_), .A2(\shift[1] ), .ZN(new_n986_));
  OR2_X2     g0700(.A1(\a[26] ), .A2(\shift[1] ), .Z(new_n987_));
  NAND3_X1   g0701(.A1(new_n309_), .A2(new_n986_), .A3(new_n987_), .ZN(new_n988_));
  NOR3_X1    g0702(.A1(new_n988_), .A2(new_n984_), .A3(new_n315_), .ZN(new_n989_));
  NAND2_X1   g0703(.A1(new_n672_), .A2(\shift[0] ), .ZN(new_n991_));
  OAI21_X1   g0704(.A1(\a[31] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n992_));
  NAND2_X1   g0705(.A1(new_n992_), .A2(new_n991_), .ZN(new_n993_));
  INV_X1     g0706(.I(new_n993_), .ZN(new_n994_));
  NOR2_X1    g0707(.A1(new_n284_), .A2(\a[29] ), .ZN(new_n995_));
  NOR2_X1    g0708(.A1(\a[30] ), .A2(\shift[1] ), .ZN(new_n996_));
  NOR2_X1    g0709(.A1(new_n995_), .A2(new_n996_), .ZN(new_n997_));
  NAND2_X1   g0710(.A1(new_n997_), .A2(new_n309_), .ZN(new_n998_));
  NOR3_X1    g0711(.A1(new_n994_), .A2(new_n998_), .A3(new_n315_), .ZN(new_n999_));
  NOR4_X1    g0712(.A1(new_n982_), .A2(new_n999_), .A3(new_n973_), .A4(new_n989_), .ZN(new_n1000_));
  NAND2_X1   g0713(.A1(new_n1000_), .A2(new_n270_), .ZN(new_n1001_));
  NAND2_X1   g0714(.A1(new_n563_), .A2(\shift[0] ), .ZN(new_n1003_));
  OAI21_X1   g0715(.A1(\a[7] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n1004_));
  NAND2_X1   g0716(.A1(new_n1004_), .A2(new_n1003_), .ZN(new_n1005_));
  INV_X1     g0717(.I(\a[5] ), .ZN(new_n1006_));
  NAND2_X1   g0718(.A1(new_n1006_), .A2(\shift[1] ), .ZN(new_n1007_));
  OAI21_X1   g0719(.A1(\a[6] ), .A2(\shift[1] ), .B(new_n1007_), .ZN(new_n1008_));
  NOR2_X1    g0720(.A1(new_n1008_), .A2(new_n283_), .ZN(new_n1009_));
  AOI21_X1   g0721(.A1(new_n1009_), .A2(new_n1005_), .B(new_n291_), .ZN(new_n1010_));
  NAND2_X1   g0722(.A1(new_n576_), .A2(\shift[0] ), .ZN(new_n1012_));
  OAI21_X1   g0723(.A1(\a[19] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n1013_));
  NAND2_X1   g0724(.A1(new_n1013_), .A2(new_n1012_), .ZN(new_n1014_));
  INV_X1     g0725(.I(new_n1014_), .ZN(new_n1015_));
  INV_X1     g0726(.I(\a[17] ), .ZN(new_n1016_));
  NAND2_X1   g0727(.A1(new_n1016_), .A2(\shift[1] ), .ZN(new_n1017_));
  OR2_X2     g0728(.A1(\a[18] ), .A2(\shift[1] ), .Z(new_n1018_));
  NAND3_X1   g0729(.A1(new_n309_), .A2(new_n1017_), .A3(new_n1018_), .ZN(new_n1019_));
  OAI21_X1   g0730(.A1(new_n1015_), .A2(new_n1019_), .B(new_n278_), .ZN(new_n1020_));
  NAND2_X1   g0731(.A1(new_n589_), .A2(\shift[0] ), .ZN(new_n1022_));
  OAI21_X1   g0732(.A1(\a[11] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n1023_));
  AND2_X2    g0733(.A1(new_n1023_), .A2(new_n1022_), .Z(new_n1024_));
  INV_X1     g0734(.I(\a[9] ), .ZN(new_n1025_));
  NAND2_X1   g0735(.A1(new_n1025_), .A2(\shift[1] ), .ZN(new_n1026_));
  NAND2_X1   g0736(.A1(new_n596_), .A2(new_n284_), .ZN(new_n1027_));
  NAND3_X1   g0737(.A1(new_n309_), .A2(new_n1026_), .A3(new_n1027_), .ZN(new_n1028_));
  NOR3_X1    g0738(.A1(new_n1024_), .A2(new_n1028_), .A3(new_n315_), .ZN(new_n1029_));
  NAND2_X1   g0739(.A1(new_n601_), .A2(\shift[0] ), .ZN(new_n1031_));
  OAI21_X1   g0740(.A1(\a[15] ), .A2(\shift[1] ), .B(new_n279_), .ZN(new_n1032_));
  AND2_X2    g0741(.A1(new_n1032_), .A2(new_n1031_), .Z(new_n1033_));
  INV_X1     g0742(.I(\a[13] ), .ZN(new_n1034_));
  NAND2_X1   g0743(.A1(new_n1034_), .A2(\shift[1] ), .ZN(new_n1035_));
  NAND2_X1   g0744(.A1(new_n571_), .A2(new_n284_), .ZN(new_n1036_));
  NAND3_X1   g0745(.A1(new_n309_), .A2(new_n1035_), .A3(new_n1036_), .ZN(new_n1037_));
  NOR3_X1    g0746(.A1(new_n1033_), .A2(new_n1037_), .A3(new_n315_), .ZN(new_n1038_));
  NOR4_X1    g0747(.A1(new_n1010_), .A2(new_n1020_), .A3(new_n1029_), .A4(new_n1038_), .ZN(new_n1039_));
  AOI21_X1   g0748(.A1(new_n1039_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1040_));
  NAND2_X1   g0749(.A1(new_n1040_), .A2(new_n1001_), .ZN(new_n1041_));
  OAI21_X1   g0750(.A1(new_n963_), .A2(new_n1041_), .B(\shift[6] ), .ZN(new_n1042_));
  OAI21_X1   g0751(.A1(new_n900_), .A2(\shift[6] ), .B(new_n1042_), .ZN(\result[3] ));
  NOR2_X1    g0752(.A1(\shift[2] ), .A2(\shift[3] ), .ZN(new_n1044_));
  NOR4_X1    g0753(.A1(new_n267_), .A2(new_n270_), .A3(\shift[5] ), .A4(new_n1044_), .ZN(new_n1045_));
  OAI21_X1   g0754(.A1(new_n264_), .A2(new_n1045_), .B(new_n269_), .ZN(\result[4] ));
  OAI21_X1   g0755(.A1(new_n342_), .A2(new_n346_), .B(new_n278_), .ZN(new_n1047_));
  AOI21_X1   g0756(.A1(new_n882_), .A2(new_n284_), .B(\shift[0] ), .ZN(new_n1048_));
  XOR2_X1    g0757(.A1(new_n1048_), .A2(new_n318_), .Z(new_n1049_));
  AND2_X2    g0758(.A1(new_n309_), .A2(new_n323_), .Z(new_n1050_));
  AOI21_X1   g0759(.A1(new_n1049_), .A2(new_n1050_), .B(new_n291_), .ZN(new_n1051_));
  NOR3_X1    g0760(.A1(new_n308_), .A2(new_n315_), .A3(new_n313_), .ZN(new_n1052_));
  NOR4_X1    g0761(.A1(new_n1051_), .A2(new_n335_), .A3(new_n1047_), .A4(new_n1052_), .ZN(new_n1053_));
  NOR2_X1    g0762(.A1(new_n1053_), .A2(new_n270_), .ZN(new_n1054_));
  NAND2_X1   g0763(.A1(new_n357_), .A2(new_n278_), .ZN(new_n1055_));
  AOI21_X1   g0764(.A1(new_n609_), .A2(new_n610_), .B(new_n315_), .ZN(new_n1056_));
  NOR3_X1    g0765(.A1(new_n279_), .A2(\a[118] ), .A3(\shift[1] ), .ZN(new_n1057_));
  NOR3_X1    g0766(.A1(new_n361_), .A2(\shift[0] ), .A3(new_n359_), .ZN(new_n1058_));
  NOR2_X1    g0767(.A1(new_n1058_), .A2(new_n1057_), .ZN(new_n1059_));
  NOR2_X1    g0768(.A1(new_n363_), .A2(new_n364_), .ZN(new_n1060_));
  NAND2_X1   g0769(.A1(new_n1060_), .A2(new_n309_), .ZN(new_n1061_));
  OAI21_X1   g0770(.A1(new_n1059_), .A2(new_n1061_), .B(new_n277_), .ZN(new_n1062_));
  NAND4_X1   g0771(.A1(new_n1055_), .A2(new_n378_), .A3(new_n1056_), .A4(new_n1062_), .ZN(new_n1063_));
  OAI21_X1   g0772(.A1(new_n1063_), .A2(new_n270_), .B(new_n265_), .ZN(new_n1064_));
  NOR2_X1    g0773(.A1(new_n1064_), .A2(new_n1054_), .ZN(new_n1065_));
  NOR3_X1    g0774(.A1(new_n279_), .A2(\a[90] ), .A3(\shift[1] ), .ZN(new_n1066_));
  NOR3_X1    g0775(.A1(new_n1066_), .A2(\shift[0] ), .A3(new_n417_), .ZN(new_n1067_));
  NOR2_X1    g0776(.A1(new_n1067_), .A2(new_n418_), .ZN(new_n1068_));
  NOR2_X1    g0777(.A1(new_n425_), .A2(new_n426_), .ZN(new_n1069_));
  NAND2_X1   g0778(.A1(new_n1069_), .A2(new_n309_), .ZN(new_n1070_));
  NOR3_X1    g0779(.A1(new_n1068_), .A2(new_n315_), .A3(new_n1070_), .ZN(new_n1071_));
  NOR3_X1    g0780(.A1(new_n279_), .A2(\a[98] ), .A3(\shift[1] ), .ZN(new_n1072_));
  NOR3_X1    g0781(.A1(new_n1072_), .A2(\shift[0] ), .A3(new_n292_), .ZN(new_n1073_));
  NOR2_X1    g0782(.A1(new_n1073_), .A2(new_n293_), .ZN(new_n1074_));
  NOR2_X1    g0783(.A1(new_n300_), .A2(new_n301_), .ZN(new_n1075_));
  NAND2_X1   g0784(.A1(new_n1075_), .A2(new_n309_), .ZN(new_n1076_));
  OAI21_X1   g0785(.A1(new_n1074_), .A2(new_n1076_), .B(new_n278_), .ZN(new_n1077_));
  AOI21_X1   g0786(.A1(new_n412_), .A2(new_n415_), .B(new_n291_), .ZN(new_n1078_));
  NOR3_X1    g0787(.A1(new_n398_), .A2(new_n315_), .A3(new_n402_), .ZN(new_n1079_));
  NOR4_X1    g0788(.A1(new_n1071_), .A2(new_n1078_), .A3(new_n1079_), .A4(new_n1077_), .ZN(new_n1080_));
  NAND2_X1   g0789(.A1(new_n1080_), .A2(new_n270_), .ZN(new_n1081_));
  NOR3_X1    g0790(.A1(new_n279_), .A2(\a[82] ), .A3(\shift[1] ), .ZN(new_n1082_));
  NOR3_X1    g0791(.A1(new_n1082_), .A2(\shift[0] ), .A3(new_n382_), .ZN(new_n1083_));
  NOR2_X1    g0792(.A1(new_n1083_), .A2(new_n383_), .ZN(new_n1084_));
  NOR2_X1    g0793(.A1(new_n390_), .A2(new_n391_), .ZN(new_n1085_));
  NAND2_X1   g0794(.A1(new_n1085_), .A2(new_n309_), .ZN(new_n1086_));
  NOR2_X1    g0795(.A1(new_n1084_), .A2(new_n1086_), .ZN(new_n1087_));
  NOR3_X1    g0796(.A1(new_n279_), .A2(\a[74] ), .A3(\shift[1] ), .ZN(new_n1088_));
  NOR3_X1    g0797(.A1(new_n1088_), .A2(\shift[0] ), .A3(new_n462_), .ZN(new_n1089_));
  NOR2_X1    g0798(.A1(new_n1089_), .A2(new_n463_), .ZN(new_n1090_));
  NAND2_X1   g0799(.A1(new_n472_), .A2(new_n309_), .ZN(new_n1091_));
  NOR2_X1    g0800(.A1(new_n1090_), .A2(new_n1091_), .ZN(new_n1092_));
  NOR3_X1    g0801(.A1(new_n1087_), .A2(new_n1092_), .A3(new_n315_), .ZN(new_n1093_));
  NAND2_X1   g0802(.A1(new_n456_), .A2(new_n460_), .ZN(new_n1094_));
  AOI22_X1   g0803(.A1(new_n1094_), .A2(new_n277_), .B1(new_n278_), .B2(new_n451_), .ZN(new_n1095_));
  NAND3_X1   g0804(.A1(new_n1095_), .A2(\shift[4] ), .A3(new_n1093_), .ZN(new_n1096_));
  NAND3_X1   g0805(.A1(new_n1096_), .A2(new_n1081_), .A3(new_n265_), .ZN(new_n1097_));
  OAI21_X1   g0806(.A1(new_n1065_), .A2(new_n1097_), .B(new_n264_), .ZN(new_n1098_));
  NOR2_X1    g0807(.A1(new_n523_), .A2(new_n525_), .ZN(new_n1099_));
  NOR3_X1    g0808(.A1(new_n697_), .A2(new_n315_), .A3(new_n701_), .ZN(new_n1100_));
  NOR3_X1    g0809(.A1(new_n1100_), .A2(new_n1099_), .A3(new_n267_), .ZN(new_n1101_));
  OAI21_X1   g0810(.A1(new_n434_), .A2(new_n438_), .B(new_n278_), .ZN(new_n1102_));
  AOI21_X1   g0811(.A1(new_n541_), .A2(new_n542_), .B(new_n291_), .ZN(new_n1103_));
  NOR3_X1    g0812(.A1(new_n493_), .A2(new_n315_), .A3(new_n497_), .ZN(new_n1104_));
  NOR4_X1    g0813(.A1(new_n518_), .A2(new_n1103_), .A3(new_n1104_), .A4(new_n1102_), .ZN(new_n1105_));
  AOI21_X1   g0814(.A1(new_n1105_), .A2(new_n270_), .B(new_n1101_), .ZN(new_n1106_));
  OR3_X2     g0815(.A1(new_n1100_), .A2(new_n267_), .A3(new_n1099_), .Z(new_n1107_));
  NOR3_X1    g0816(.A1(new_n1107_), .A2(new_n1105_), .A3(\shift[4] ), .ZN(new_n1108_));
  NOR3_X1    g0817(.A1(new_n1108_), .A2(new_n1106_), .A3(\shift[5] ), .ZN(new_n1109_));
  NOR3_X1    g0818(.A1(new_n283_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n1110_));
  OAI21_X1   g0819(.A1(new_n667_), .A2(new_n669_), .B(new_n1110_), .ZN(new_n1111_));
  NAND2_X1   g0820(.A1(new_n688_), .A2(new_n691_), .ZN(new_n1112_));
  NAND3_X1   g0821(.A1(new_n1111_), .A2(new_n1112_), .A3(new_n278_), .ZN(new_n1113_));
  NOR2_X1    g0822(.A1(new_n656_), .A2(\shift[0] ), .ZN(new_n1114_));
  XOR2_X1    g0823(.A1(new_n1114_), .A2(new_n658_), .Z(new_n1115_));
  NAND2_X1   g0824(.A1(new_n663_), .A2(new_n662_), .ZN(new_n1116_));
  NOR2_X1    g0825(.A1(new_n1116_), .A2(new_n283_), .ZN(new_n1117_));
  AOI21_X1   g0826(.A1(new_n1115_), .A2(new_n1117_), .B(new_n291_), .ZN(new_n1118_));
  NOR3_X1    g0827(.A1(new_n650_), .A2(new_n315_), .A3(new_n654_), .ZN(new_n1119_));
  NOR3_X1    g0828(.A1(new_n1113_), .A2(new_n1118_), .A3(new_n1119_), .ZN(new_n1120_));
  NOR3_X1    g0829(.A1(new_n279_), .A2(\a[18] ), .A3(\shift[1] ), .ZN(new_n1121_));
  NOR3_X1    g0830(.A1(new_n635_), .A2(\shift[0] ), .A3(new_n633_), .ZN(new_n1122_));
  NOR2_X1    g0831(.A1(new_n1122_), .A2(new_n1121_), .ZN(new_n1123_));
  NAND2_X1   g0832(.A1(new_n309_), .A2(new_n639_), .ZN(new_n1124_));
  OAI21_X1   g0833(.A1(new_n1123_), .A2(new_n1124_), .B(new_n278_), .ZN(new_n1125_));
  AOI21_X1   g0834(.A1(new_n587_), .A2(new_n590_), .B(new_n291_), .ZN(new_n1126_));
  NOR3_X1    g0835(.A1(new_n614_), .A2(new_n315_), .A3(new_n616_), .ZN(new_n1127_));
  NOR4_X1    g0836(.A1(new_n629_), .A2(new_n1126_), .A3(new_n1127_), .A4(new_n1125_), .ZN(new_n1128_));
  NAND4_X1   g0837(.A1(new_n1120_), .A2(\shift[4] ), .A3(new_n265_), .A4(new_n1128_), .ZN(new_n1129_));
  OAI21_X1   g0838(.A1(new_n1109_), .A2(new_n1129_), .B(\shift[6] ), .ZN(new_n1130_));
  NAND2_X1   g0839(.A1(new_n1130_), .A2(new_n1098_), .ZN(\result[5] ));
  INV_X1     g0840(.I(new_n714_), .ZN(new_n1132_));
  NOR2_X1    g0841(.A1(new_n267_), .A2(\shift[5] ), .ZN(new_n1133_));
  INV_X1     g0842(.I(new_n1133_), .ZN(new_n1134_));
  OAI21_X1   g0843(.A1(new_n270_), .A2(new_n266_), .B(new_n1134_), .ZN(new_n1135_));
  OAI21_X1   g0844(.A1(new_n1132_), .A2(new_n1135_), .B(\shift[6] ), .ZN(new_n1136_));
  NAND2_X1   g0845(.A1(new_n1136_), .A2(new_n269_), .ZN(\result[6] ));
  OAI21_X1   g0846(.A1(new_n757_), .A2(new_n727_), .B(new_n278_), .ZN(new_n1138_));
  NAND2_X1   g0847(.A1(new_n880_), .A2(new_n879_), .ZN(new_n1139_));
  INV_X1     g0848(.I(new_n885_), .ZN(new_n1140_));
  AOI21_X1   g0849(.A1(new_n1140_), .A2(new_n1139_), .B(new_n291_), .ZN(new_n1141_));
  NOR2_X1    g0850(.A1(new_n875_), .A2(new_n315_), .ZN(new_n1142_));
  NOR4_X1    g0851(.A1(new_n1141_), .A2(new_n1142_), .A3(new_n896_), .A4(new_n1138_), .ZN(new_n1143_));
  NOR2_X1    g0852(.A1(new_n1143_), .A2(new_n270_), .ZN(new_n1144_));
  NAND2_X1   g0853(.A1(new_n1009_), .A2(new_n1005_), .ZN(new_n1145_));
  NAND3_X1   g0854(.A1(new_n1145_), .A2(new_n278_), .A3(new_n753_), .ZN(new_n1146_));
  INV_X1     g0855(.I(new_n740_), .ZN(new_n1147_));
  NAND3_X1   g0856(.A1(new_n309_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n1148_));
  OAI21_X1   g0857(.A1(new_n1147_), .A2(new_n1148_), .B(new_n277_), .ZN(new_n1149_));
  INV_X1     g0858(.I(new_n1149_), .ZN(new_n1150_));
  NOR3_X1    g0859(.A1(new_n732_), .A2(new_n315_), .A3(new_n735_), .ZN(new_n1151_));
  NOR4_X1    g0860(.A1(new_n1146_), .A2(new_n1150_), .A3(new_n270_), .A4(new_n1151_), .ZN(new_n1152_));
  NOR3_X1    g0861(.A1(new_n1144_), .A2(new_n1152_), .A3(\shift[5] ), .ZN(new_n1153_));
  INV_X1     g0862(.I(new_n854_), .ZN(new_n1154_));
  OAI21_X1   g0863(.A1(new_n861_), .A2(new_n865_), .B(new_n278_), .ZN(new_n1155_));
  NAND2_X1   g0864(.A1(new_n309_), .A2(new_n847_), .ZN(new_n1156_));
  INV_X1     g0865(.I(new_n1156_), .ZN(new_n1157_));
  AOI21_X1   g0866(.A1(new_n1157_), .A2(new_n846_), .B(new_n291_), .ZN(new_n1158_));
  NAND2_X1   g0867(.A1(new_n838_), .A2(new_n837_), .ZN(new_n1159_));
  NAND4_X1   g0868(.A1(new_n1159_), .A2(new_n278_), .A3(new_n309_), .A4(new_n840_), .ZN(new_n1160_));
  INV_X1     g0869(.I(new_n1160_), .ZN(new_n1161_));
  NOR4_X1    g0870(.A1(new_n1158_), .A2(new_n1154_), .A3(new_n1161_), .A4(new_n1155_), .ZN(new_n1162_));
  NAND2_X1   g0871(.A1(new_n1162_), .A2(new_n270_), .ZN(new_n1163_));
  NOR3_X1    g0872(.A1(new_n821_), .A2(new_n315_), .A3(new_n834_), .ZN(new_n1164_));
  OAI21_X1   g0873(.A1(new_n815_), .A2(new_n795_), .B(new_n277_), .ZN(new_n1165_));
  NAND3_X1   g0874(.A1(new_n785_), .A2(new_n278_), .A3(new_n781_), .ZN(new_n1166_));
  NAND4_X1   g0875(.A1(new_n1164_), .A2(\shift[4] ), .A3(new_n1165_), .A4(new_n1166_), .ZN(new_n1167_));
  NAND3_X1   g0876(.A1(new_n1163_), .A2(new_n1167_), .A3(new_n265_), .ZN(new_n1168_));
  OAI21_X1   g0877(.A1(new_n1153_), .A2(new_n1168_), .B(new_n264_), .ZN(new_n1169_));
  NAND4_X1   g0878(.A1(new_n919_), .A2(new_n278_), .A3(new_n309_), .A4(new_n923_), .ZN(new_n1170_));
  OAI21_X1   g0879(.A1(new_n903_), .A2(new_n907_), .B(new_n277_), .ZN(new_n1171_));
  INV_X1     g0880(.I(new_n935_), .ZN(new_n1172_));
  NOR2_X1    g0881(.A1(new_n1172_), .A2(new_n283_), .ZN(new_n1173_));
  AOI21_X1   g0882(.A1(new_n1173_), .A2(new_n931_), .B(new_n315_), .ZN(new_n1174_));
  NAND3_X1   g0883(.A1(new_n1171_), .A2(new_n1174_), .A3(new_n1170_), .ZN(new_n1175_));
  AND2_X2    g0884(.A1(new_n953_), .A2(new_n952_), .Z(new_n1176_));
  NAND3_X1   g0885(.A1(new_n309_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n1177_));
  NOR3_X1    g0886(.A1(new_n1176_), .A2(new_n1177_), .A3(new_n315_), .ZN(new_n1178_));
  OAI21_X1   g0887(.A1(new_n772_), .A2(new_n776_), .B(new_n278_), .ZN(new_n1179_));
  AND2_X2    g0888(.A1(new_n947_), .A2(new_n946_), .Z(new_n1180_));
  NAND2_X1   g0889(.A1(new_n309_), .A2(new_n949_), .ZN(new_n1181_));
  NOR2_X1    g0890(.A1(new_n1180_), .A2(new_n1181_), .ZN(new_n1182_));
  NOR2_X1    g0891(.A1(new_n1182_), .A2(new_n291_), .ZN(new_n1183_));
  NOR2_X1    g0892(.A1(new_n943_), .A2(new_n315_), .ZN(new_n1184_));
  NOR4_X1    g0893(.A1(new_n1183_), .A2(new_n1178_), .A3(new_n1179_), .A4(new_n1184_), .ZN(new_n1185_));
  INV_X1     g0894(.I(new_n1185_), .ZN(new_n1186_));
  OAI21_X1   g0895(.A1(new_n1186_), .A2(\shift[4] ), .B(new_n1175_), .ZN(new_n1187_));
  NOR3_X1    g0896(.A1(new_n1185_), .A2(new_n1175_), .A3(\shift[4] ), .ZN(new_n1188_));
  NOR2_X1    g0897(.A1(new_n1188_), .A2(\shift[5] ), .ZN(new_n1189_));
  INV_X1     g0898(.I(new_n967_), .ZN(new_n1190_));
  NAND3_X1   g0899(.A1(new_n309_), .A2(new_n969_), .A3(new_n970_), .ZN(new_n1191_));
  OAI21_X1   g0900(.A1(new_n1190_), .A2(new_n1191_), .B(new_n278_), .ZN(new_n1192_));
  NOR2_X1    g0901(.A1(new_n1024_), .A2(new_n1028_), .ZN(new_n1193_));
  NOR2_X1    g0902(.A1(new_n1193_), .A2(new_n291_), .ZN(new_n1194_));
  NOR3_X1    g0903(.A1(new_n1015_), .A2(new_n1019_), .A3(new_n315_), .ZN(new_n1195_));
  NOR4_X1    g0904(.A1(new_n1194_), .A2(new_n1038_), .A3(new_n1192_), .A4(new_n1195_), .ZN(new_n1196_));
  INV_X1     g0905(.I(new_n911_), .ZN(new_n1197_));
  NOR2_X1    g0906(.A1(new_n912_), .A2(new_n913_), .ZN(new_n1198_));
  NAND3_X1   g0907(.A1(new_n1197_), .A2(new_n309_), .A3(new_n1198_), .ZN(new_n1199_));
  NAND3_X1   g0908(.A1(new_n993_), .A2(new_n309_), .A3(new_n997_), .ZN(new_n1200_));
  NAND3_X1   g0909(.A1(new_n1199_), .A2(new_n1200_), .A3(new_n278_), .ZN(new_n1201_));
  NOR2_X1    g0910(.A1(new_n988_), .A2(new_n984_), .ZN(new_n1202_));
  NOR2_X1    g0911(.A1(new_n1202_), .A2(new_n291_), .ZN(new_n1203_));
  AND4_X2    g0912(.A1(new_n278_), .A2(new_n977_), .A3(new_n309_), .A4(new_n980_), .Z(new_n1204_));
  NOR3_X1    g0913(.A1(new_n1201_), .A2(new_n1203_), .A3(new_n1204_), .ZN(new_n1205_));
  NAND4_X1   g0914(.A1(new_n1205_), .A2(new_n1196_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1206_));
  AOI21_X1   g0915(.A1(new_n1189_), .A2(new_n1187_), .B(new_n1206_), .ZN(new_n1207_));
  OAI21_X1   g0916(.A1(new_n1207_), .A2(new_n264_), .B(new_n1169_), .ZN(\result[7] ));
  NAND4_X1   g0917(.A1(new_n267_), .A2(\shift[4] ), .A3(new_n265_), .A4(new_n264_), .ZN(\result[8] ));
  OAI21_X1   g0918(.A1(new_n1059_), .A2(new_n1061_), .B(new_n278_), .ZN(new_n1210_));
  NOR2_X1    g0919(.A1(new_n326_), .A2(\shift[0] ), .ZN(new_n1211_));
  XOR2_X1    g0920(.A1(new_n1211_), .A2(new_n328_), .Z(new_n1212_));
  INV_X1     g0921(.I(new_n334_), .ZN(new_n1213_));
  AOI21_X1   g0922(.A1(new_n1212_), .A2(new_n1213_), .B(new_n291_), .ZN(new_n1214_));
  NOR3_X1    g0923(.A1(new_n342_), .A2(new_n315_), .A3(new_n346_), .ZN(new_n1215_));
  NOR4_X1    g0924(.A1(new_n1214_), .A2(new_n1052_), .A3(new_n1210_), .A4(new_n1215_), .ZN(new_n1216_));
  NOR2_X1    g0925(.A1(new_n1216_), .A2(new_n270_), .ZN(new_n1217_));
  NOR2_X1    g0926(.A1(new_n620_), .A2(new_n622_), .ZN(new_n1218_));
  NOR3_X1    g0927(.A1(new_n1218_), .A2(new_n315_), .A3(new_n357_), .ZN(new_n1219_));
  NOR3_X1    g0928(.A1(new_n279_), .A2(\a[122] ), .A3(\shift[1] ), .ZN(new_n1220_));
  NOR3_X1    g0929(.A1(new_n1220_), .A2(\shift[0] ), .A3(new_n367_), .ZN(new_n1221_));
  NOR2_X1    g0930(.A1(new_n1221_), .A2(new_n368_), .ZN(new_n1222_));
  NAND2_X1   g0931(.A1(new_n309_), .A2(new_n377_), .ZN(new_n1223_));
  OAI21_X1   g0932(.A1(new_n1222_), .A2(new_n1223_), .B(new_n277_), .ZN(new_n1224_));
  NAND3_X1   g0933(.A1(new_n609_), .A2(new_n610_), .A3(new_n278_), .ZN(new_n1225_));
  NAND4_X1   g0934(.A1(new_n1219_), .A2(\shift[4] ), .A3(new_n1224_), .A4(new_n1225_), .ZN(new_n1226_));
  NAND2_X1   g0935(.A1(new_n1226_), .A2(new_n265_), .ZN(new_n1227_));
  NOR2_X1    g0936(.A1(new_n1227_), .A2(new_n1217_), .ZN(new_n1228_));
  OAI21_X1   g0937(.A1(new_n320_), .A2(new_n324_), .B(new_n278_), .ZN(new_n1229_));
  AOI21_X1   g0938(.A1(new_n424_), .A2(new_n427_), .B(new_n291_), .ZN(new_n1230_));
  NOR3_X1    g0939(.A1(new_n1074_), .A2(new_n315_), .A3(new_n1076_), .ZN(new_n1231_));
  NOR4_X1    g0940(.A1(new_n1079_), .A2(new_n1230_), .A3(new_n1231_), .A4(new_n1229_), .ZN(new_n1232_));
  NAND2_X1   g0941(.A1(new_n1232_), .A2(new_n270_), .ZN(new_n1233_));
  NOR3_X1    g0942(.A1(new_n279_), .A2(\a[86] ), .A3(\shift[1] ), .ZN(new_n1234_));
  NOR3_X1    g0943(.A1(new_n1234_), .A2(\shift[0] ), .A3(new_n405_), .ZN(new_n1235_));
  NOR2_X1    g0944(.A1(new_n1235_), .A2(new_n406_), .ZN(new_n1236_));
  NOR2_X1    g0945(.A1(new_n413_), .A2(new_n414_), .ZN(new_n1237_));
  NAND2_X1   g0946(.A1(new_n1237_), .A2(new_n309_), .ZN(new_n1238_));
  NOR2_X1    g0947(.A1(new_n1236_), .A2(new_n1238_), .ZN(new_n1239_));
  NOR3_X1    g0948(.A1(new_n451_), .A2(new_n1239_), .A3(new_n315_), .ZN(new_n1240_));
  OAI21_X1   g0949(.A1(new_n1090_), .A2(new_n1091_), .B(new_n277_), .ZN(new_n1241_));
  NAND3_X1   g0950(.A1(new_n389_), .A2(new_n392_), .A3(new_n278_), .ZN(new_n1242_));
  NAND4_X1   g0951(.A1(new_n1240_), .A2(\shift[4] ), .A3(new_n1241_), .A4(new_n1242_), .ZN(new_n1243_));
  NAND3_X1   g0952(.A1(new_n1233_), .A2(new_n1243_), .A3(new_n265_), .ZN(new_n1244_));
  OAI21_X1   g0953(.A1(new_n1228_), .A2(new_n1244_), .B(new_n264_), .ZN(new_n1245_));
  NOR2_X1    g0954(.A1(new_n503_), .A2(new_n507_), .ZN(new_n1246_));
  NOR3_X1    g0955(.A1(new_n523_), .A2(new_n315_), .A3(new_n525_), .ZN(new_n1247_));
  NOR4_X1    g0956(.A1(new_n1100_), .A2(new_n1247_), .A3(new_n1246_), .A4(new_n267_), .ZN(new_n1248_));
  NOR3_X1    g0957(.A1(new_n279_), .A2(\a[70] ), .A3(\shift[1] ), .ZN(new_n1249_));
  NOR3_X1    g0958(.A1(new_n455_), .A2(\shift[0] ), .A3(new_n453_), .ZN(new_n1250_));
  NOR2_X1    g0959(.A1(new_n1250_), .A2(new_n1249_), .ZN(new_n1251_));
  NAND2_X1   g0960(.A1(new_n309_), .A2(new_n459_), .ZN(new_n1252_));
  OAI21_X1   g0961(.A1(new_n1251_), .A2(new_n1252_), .B(new_n278_), .ZN(new_n1253_));
  AOI21_X1   g0962(.A1(new_n549_), .A2(new_n550_), .B(new_n291_), .ZN(new_n1254_));
  NOR3_X1    g0963(.A1(new_n434_), .A2(new_n315_), .A3(new_n438_), .ZN(new_n1255_));
  NOR4_X1    g0964(.A1(new_n1104_), .A2(new_n1254_), .A3(new_n1255_), .A4(new_n1253_), .ZN(new_n1256_));
  AOI21_X1   g0965(.A1(new_n1256_), .A2(new_n270_), .B(new_n1248_), .ZN(new_n1257_));
  NOR2_X1    g0966(.A1(new_n693_), .A2(\shift[0] ), .ZN(new_n1258_));
  XOR2_X1    g0967(.A1(new_n1258_), .A2(new_n695_), .Z(new_n1259_));
  NOR3_X1    g0968(.A1(new_n283_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n1260_));
  NAND3_X1   g0969(.A1(new_n1259_), .A2(new_n1260_), .A3(new_n278_), .ZN(new_n1261_));
  NAND3_X1   g0970(.A1(new_n484_), .A2(new_n487_), .A3(new_n278_), .ZN(new_n1262_));
  NAND4_X1   g0971(.A1(new_n1261_), .A2(new_n266_), .A3(new_n543_), .A4(new_n1262_), .ZN(new_n1263_));
  NOR3_X1    g0972(.A1(new_n1256_), .A2(new_n1263_), .A3(\shift[4] ), .ZN(new_n1264_));
  NOR3_X1    g0973(.A1(new_n1264_), .A2(new_n1257_), .A3(\shift[5] ), .ZN(new_n1265_));
  OAI21_X1   g0974(.A1(new_n660_), .A2(new_n664_), .B(new_n278_), .ZN(new_n1266_));
  AOI21_X1   g0975(.A1(new_n599_), .A2(new_n602_), .B(new_n291_), .ZN(new_n1267_));
  NOR3_X1    g0976(.A1(new_n1123_), .A2(new_n315_), .A3(new_n1124_), .ZN(new_n1268_));
  NOR4_X1    g0977(.A1(new_n1127_), .A2(new_n1267_), .A3(new_n1268_), .A4(new_n1266_), .ZN(new_n1269_));
  OAI21_X1   g0978(.A1(new_n650_), .A2(new_n654_), .B(new_n278_), .ZN(new_n1270_));
  OAI21_X1   g0979(.A1(new_n670_), .A2(new_n674_), .B(new_n277_), .ZN(new_n1271_));
  INV_X1     g0980(.I(new_n1271_), .ZN(new_n1272_));
  NAND3_X1   g0981(.A1(new_n688_), .A2(new_n691_), .A3(new_n278_), .ZN(new_n1273_));
  INV_X1     g0982(.I(new_n1273_), .ZN(new_n1274_));
  NOR3_X1    g0983(.A1(new_n1272_), .A2(new_n1274_), .A3(new_n1270_), .ZN(new_n1275_));
  NAND4_X1   g0984(.A1(new_n1275_), .A2(\shift[4] ), .A3(new_n1269_), .A4(new_n265_), .ZN(new_n1276_));
  OAI21_X1   g0985(.A1(new_n1265_), .A2(new_n1276_), .B(\shift[6] ), .ZN(new_n1277_));
  NAND2_X1   g0986(.A1(new_n1277_), .A2(new_n1245_), .ZN(\result[9] ));
  NOR2_X1    g0987(.A1(new_n710_), .A2(\shift[5] ), .ZN(new_n1279_));
  INV_X1     g0988(.I(new_n1279_), .ZN(new_n1280_));
  NOR2_X1    g0989(.A1(new_n1280_), .A2(new_n1135_), .ZN(new_n1281_));
  OAI21_X1   g0990(.A1(new_n1281_), .A2(new_n264_), .B(new_n269_), .ZN(\result[10] ));
  OAI21_X1   g0991(.A1(new_n1147_), .A2(new_n1148_), .B(new_n278_), .ZN(new_n1283_));
  NAND2_X1   g0992(.A1(new_n889_), .A2(new_n888_), .ZN(new_n1284_));
  NAND2_X1   g0993(.A1(new_n894_), .A2(new_n892_), .ZN(new_n1285_));
  NOR2_X1    g0994(.A1(new_n1285_), .A2(new_n283_), .ZN(new_n1286_));
  AOI21_X1   g0995(.A1(new_n1286_), .A2(new_n1284_), .B(new_n291_), .ZN(new_n1287_));
  NOR3_X1    g0996(.A1(new_n757_), .A2(new_n727_), .A3(new_n315_), .ZN(new_n1288_));
  NOR4_X1    g0997(.A1(new_n1142_), .A2(new_n1283_), .A3(new_n1288_), .A4(new_n1287_), .ZN(new_n1289_));
  NOR2_X1    g0998(.A1(new_n1289_), .A2(new_n270_), .ZN(new_n1290_));
  NAND3_X1   g0999(.A1(new_n761_), .A2(new_n278_), .A3(new_n763_), .ZN(new_n1291_));
  NAND2_X1   g1000(.A1(new_n1023_), .A2(new_n1022_), .ZN(new_n1292_));
  OAI21_X1   g1001(.A1(\a[10] ), .A2(\shift[1] ), .B(new_n1026_), .ZN(new_n1293_));
  NOR2_X1    g1002(.A1(new_n1293_), .A2(new_n283_), .ZN(new_n1294_));
  AOI21_X1   g1003(.A1(new_n1294_), .A2(new_n1292_), .B(new_n315_), .ZN(new_n1295_));
  NAND3_X1   g1004(.A1(new_n749_), .A2(new_n309_), .A3(new_n752_), .ZN(new_n1296_));
  NAND2_X1   g1005(.A1(new_n1296_), .A2(new_n277_), .ZN(new_n1297_));
  NAND3_X1   g1006(.A1(new_n1009_), .A2(new_n278_), .A3(new_n1005_), .ZN(new_n1298_));
  NAND4_X1   g1007(.A1(new_n1291_), .A2(new_n1295_), .A3(new_n1297_), .A4(new_n1298_), .ZN(new_n1299_));
  OAI21_X1   g1008(.A1(new_n1299_), .A2(new_n270_), .B(new_n265_), .ZN(new_n1300_));
  NOR2_X1    g1009(.A1(new_n1300_), .A2(new_n1290_), .ZN(new_n1301_));
  OAI21_X1   g1010(.A1(new_n881_), .A2(new_n885_), .B(new_n278_), .ZN(new_n1302_));
  AND2_X2    g1011(.A1(new_n309_), .A2(new_n853_), .Z(new_n1303_));
  AOI21_X1   g1012(.A1(new_n1303_), .A2(new_n852_), .B(new_n291_), .ZN(new_n1304_));
  NOR3_X1    g1013(.A1(new_n861_), .A2(new_n865_), .A3(new_n315_), .ZN(new_n1305_));
  NOR4_X1    g1014(.A1(new_n1304_), .A2(new_n1161_), .A3(new_n1302_), .A4(new_n1305_), .ZN(new_n1306_));
  NAND2_X1   g1015(.A1(new_n1306_), .A2(new_n270_), .ZN(new_n1307_));
  NOR3_X1    g1016(.A1(new_n811_), .A2(new_n813_), .A3(new_n315_), .ZN(new_n1308_));
  NAND3_X1   g1017(.A1(new_n846_), .A2(new_n309_), .A3(new_n847_), .ZN(new_n1309_));
  NAND2_X1   g1018(.A1(new_n1309_), .A2(new_n278_), .ZN(new_n1310_));
  AOI21_X1   g1019(.A1(new_n805_), .A2(new_n801_), .B(new_n291_), .ZN(new_n1311_));
  NOR4_X1    g1020(.A1(new_n833_), .A2(new_n830_), .A3(new_n315_), .A4(new_n283_), .ZN(new_n1312_));
  NOR4_X1    g1021(.A1(new_n1310_), .A2(new_n1311_), .A3(new_n1308_), .A4(new_n1312_), .ZN(new_n1313_));
  AOI21_X1   g1022(.A1(new_n1313_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1314_));
  NAND2_X1   g1023(.A1(new_n1314_), .A2(new_n1307_), .ZN(new_n1315_));
  OAI21_X1   g1024(.A1(new_n1301_), .A2(new_n1315_), .B(new_n264_), .ZN(new_n1316_));
  NAND3_X1   g1025(.A1(new_n1173_), .A2(new_n278_), .A3(new_n931_), .ZN(new_n1317_));
  NOR2_X1    g1026(.A1(new_n1182_), .A2(new_n267_), .ZN(new_n1318_));
  NAND3_X1   g1027(.A1(new_n1318_), .A2(new_n1170_), .A3(new_n1317_), .ZN(new_n1319_));
  OAI21_X1   g1028(.A1(new_n815_), .A2(new_n795_), .B(new_n278_), .ZN(new_n1320_));
  NOR2_X1    g1029(.A1(new_n1176_), .A2(new_n1177_), .ZN(new_n1321_));
  NOR2_X1    g1030(.A1(new_n1321_), .A2(new_n291_), .ZN(new_n1322_));
  NOR3_X1    g1031(.A1(new_n772_), .A2(new_n776_), .A3(new_n315_), .ZN(new_n1323_));
  NOR4_X1    g1032(.A1(new_n1322_), .A2(new_n1184_), .A3(new_n1320_), .A4(new_n1323_), .ZN(new_n1324_));
  INV_X1     g1033(.I(new_n1324_), .ZN(new_n1325_));
  OAI21_X1   g1034(.A1(new_n1325_), .A2(\shift[4] ), .B(new_n1319_), .ZN(new_n1326_));
  NOR3_X1    g1035(.A1(new_n1324_), .A2(new_n1319_), .A3(\shift[4] ), .ZN(new_n1327_));
  NOR2_X1    g1036(.A1(new_n1327_), .A2(\shift[5] ), .ZN(new_n1328_));
  OR2_X2     g1037(.A1(new_n988_), .A2(new_n984_), .Z(new_n1329_));
  NAND2_X1   g1038(.A1(new_n1018_), .A2(new_n1017_), .ZN(new_n1330_));
  NOR2_X1    g1039(.A1(new_n1330_), .A2(new_n283_), .ZN(new_n1331_));
  NAND2_X1   g1040(.A1(new_n1331_), .A2(new_n1014_), .ZN(new_n1332_));
  NAND3_X1   g1041(.A1(new_n1329_), .A2(new_n278_), .A3(new_n1332_), .ZN(new_n1333_));
  NAND2_X1   g1042(.A1(new_n1032_), .A2(new_n1031_), .ZN(new_n1334_));
  NAND2_X1   g1043(.A1(new_n1036_), .A2(new_n1035_), .ZN(new_n1335_));
  NOR2_X1    g1044(.A1(new_n1335_), .A2(new_n283_), .ZN(new_n1336_));
  AOI21_X1   g1045(.A1(new_n1336_), .A2(new_n1334_), .B(new_n291_), .ZN(new_n1337_));
  NOR3_X1    g1046(.A1(new_n1190_), .A2(new_n1191_), .A3(new_n315_), .ZN(new_n1338_));
  OR2_X2     g1047(.A1(new_n1338_), .A2(new_n1337_), .Z(new_n1339_));
  OAI21_X1   g1048(.A1(new_n1339_), .A2(new_n1333_), .B(\shift[4] ), .ZN(new_n1340_));
  OAI21_X1   g1049(.A1(new_n903_), .A2(new_n907_), .B(new_n440_), .ZN(new_n1341_));
  NAND2_X1   g1050(.A1(new_n1200_), .A2(new_n277_), .ZN(new_n1342_));
  NAND2_X1   g1051(.A1(new_n914_), .A2(new_n278_), .ZN(new_n1343_));
  NAND2_X1   g1052(.A1(new_n1343_), .A2(new_n1342_), .ZN(new_n1344_));
  NOR4_X1    g1053(.A1(new_n1344_), .A2(\shift[5] ), .A3(new_n1204_), .A4(new_n1341_), .ZN(new_n1345_));
  NAND2_X1   g1054(.A1(new_n1340_), .A2(new_n1345_), .ZN(new_n1346_));
  AOI21_X1   g1055(.A1(new_n1328_), .A2(new_n1326_), .B(new_n1346_), .ZN(new_n1347_));
  OAI21_X1   g1056(.A1(new_n1347_), .A2(new_n264_), .B(new_n1316_), .ZN(\result[11] ));
  AOI21_X1   g1057(.A1(new_n287_), .A2(new_n278_), .B(new_n710_), .ZN(new_n1349_));
  INV_X1     g1058(.I(new_n1349_), .ZN(new_n1350_));
  NOR3_X1    g1059(.A1(new_n1350_), .A2(\shift[5] ), .A3(new_n1135_), .ZN(new_n1351_));
  OAI21_X1   g1060(.A1(new_n1351_), .A2(new_n264_), .B(new_n269_), .ZN(\result[12] ));
  NOR3_X1    g1061(.A1(new_n1059_), .A2(new_n315_), .A3(new_n1061_), .ZN(new_n1353_));
  OAI21_X1   g1062(.A1(new_n1222_), .A2(new_n1223_), .B(new_n278_), .ZN(new_n1354_));
  INV_X1     g1063(.I(new_n305_), .ZN(new_n1355_));
  NOR2_X1    g1064(.A1(new_n304_), .A2(\shift[0] ), .ZN(new_n1356_));
  NAND3_X1   g1065(.A1(new_n893_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n1357_));
  NAND2_X1   g1066(.A1(new_n1356_), .A2(new_n1357_), .ZN(new_n1358_));
  NAND2_X1   g1067(.A1(new_n1358_), .A2(new_n1355_), .ZN(new_n1359_));
  INV_X1     g1068(.I(new_n313_), .ZN(new_n1360_));
  AOI21_X1   g1069(.A1(new_n1360_), .A2(new_n1359_), .B(new_n291_), .ZN(new_n1361_));
  NOR4_X1    g1070(.A1(new_n1361_), .A2(new_n1353_), .A3(new_n1215_), .A4(new_n1354_), .ZN(new_n1362_));
  NOR2_X1    g1071(.A1(new_n1362_), .A2(new_n270_), .ZN(new_n1363_));
  NAND3_X1   g1072(.A1(new_n309_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n1364_));
  NAND2_X1   g1073(.A1(new_n352_), .A2(\shift[0] ), .ZN(new_n1365_));
  NAND3_X1   g1074(.A1(new_n1365_), .A2(\a[126] ), .A3(\shift[1] ), .ZN(new_n1366_));
  NAND2_X1   g1075(.A1(new_n1366_), .A2(new_n354_), .ZN(new_n1367_));
  OAI21_X1   g1076(.A1(new_n1367_), .A2(new_n1364_), .B(new_n277_), .ZN(new_n1368_));
  AOI21_X1   g1077(.A1(new_n599_), .A2(new_n602_), .B(new_n315_), .ZN(new_n1369_));
  NAND4_X1   g1078(.A1(new_n591_), .A2(new_n1369_), .A3(new_n1225_), .A4(new_n1368_), .ZN(new_n1370_));
  OAI21_X1   g1079(.A1(new_n1370_), .A2(new_n270_), .B(new_n265_), .ZN(new_n1371_));
  NOR2_X1    g1080(.A1(new_n1363_), .A2(new_n1371_), .ZN(new_n1372_));
  NAND3_X1   g1081(.A1(new_n299_), .A2(new_n302_), .A3(new_n278_), .ZN(new_n1373_));
  OAI21_X1   g1082(.A1(new_n330_), .A2(new_n334_), .B(new_n278_), .ZN(new_n1374_));
  NOR2_X1    g1083(.A1(new_n325_), .A2(new_n1374_), .ZN(new_n1375_));
  OAI21_X1   g1084(.A1(new_n398_), .A2(new_n402_), .B(new_n277_), .ZN(new_n1376_));
  NAND4_X1   g1085(.A1(new_n1375_), .A2(new_n270_), .A3(new_n1373_), .A4(new_n1376_), .ZN(new_n1377_));
  NOR3_X1    g1086(.A1(new_n1236_), .A2(new_n315_), .A3(new_n1238_), .ZN(new_n1378_));
  OAI21_X1   g1087(.A1(new_n1068_), .A2(new_n1070_), .B(new_n278_), .ZN(new_n1379_));
  NOR2_X1    g1088(.A1(new_n1378_), .A2(new_n1379_), .ZN(new_n1380_));
  OAI21_X1   g1089(.A1(new_n446_), .A2(new_n450_), .B(new_n277_), .ZN(new_n1381_));
  NAND4_X1   g1090(.A1(new_n1380_), .A2(\shift[4] ), .A3(new_n1242_), .A4(new_n1381_), .ZN(new_n1382_));
  NAND3_X1   g1091(.A1(new_n1377_), .A2(new_n1382_), .A3(new_n265_), .ZN(new_n1383_));
  OAI21_X1   g1092(.A1(new_n1372_), .A2(new_n1383_), .B(new_n264_), .ZN(new_n1384_));
  NAND3_X1   g1093(.A1(new_n541_), .A2(new_n542_), .A3(new_n278_), .ZN(new_n1385_));
  AOI21_X1   g1094(.A1(new_n549_), .A2(new_n550_), .B(new_n315_), .ZN(new_n1386_));
  OAI21_X1   g1095(.A1(new_n697_), .A2(new_n701_), .B(new_n277_), .ZN(new_n1387_));
  NAND4_X1   g1096(.A1(new_n1385_), .A2(new_n1386_), .A3(new_n1387_), .A4(new_n1262_), .ZN(new_n1388_));
  NOR3_X1    g1097(.A1(new_n1251_), .A2(new_n315_), .A3(new_n1252_), .ZN(new_n1389_));
  OAI21_X1   g1098(.A1(new_n1090_), .A2(new_n1091_), .B(new_n278_), .ZN(new_n1390_));
  AOI21_X1   g1099(.A1(new_n533_), .A2(new_n532_), .B(new_n291_), .ZN(new_n1391_));
  NOR4_X1    g1100(.A1(new_n1391_), .A2(new_n1389_), .A3(new_n1255_), .A4(new_n1390_), .ZN(new_n1392_));
  INV_X1     g1101(.I(new_n1392_), .ZN(new_n1393_));
  OAI21_X1   g1102(.A1(new_n1393_), .A2(\shift[4] ), .B(new_n1388_), .ZN(new_n1394_));
  NOR3_X1    g1103(.A1(new_n1392_), .A2(new_n1388_), .A3(\shift[4] ), .ZN(new_n1395_));
  NOR2_X1    g1104(.A1(new_n1395_), .A2(\shift[5] ), .ZN(new_n1396_));
  OAI21_X1   g1105(.A1(new_n670_), .A2(new_n674_), .B(new_n278_), .ZN(new_n1397_));
  AOI21_X1   g1106(.A1(new_n574_), .A2(new_n577_), .B(new_n291_), .ZN(new_n1398_));
  NOR4_X1    g1107(.A1(new_n665_), .A2(new_n1268_), .A3(new_n1398_), .A4(new_n1397_), .ZN(new_n1399_));
  OAI21_X1   g1108(.A1(new_n650_), .A2(new_n654_), .B(new_n277_), .ZN(new_n1400_));
  NAND4_X1   g1109(.A1(new_n1400_), .A2(new_n1273_), .A3(new_n265_), .A4(new_n440_), .ZN(new_n1401_));
  INV_X1     g1110(.I(new_n1401_), .ZN(new_n1402_));
  OAI21_X1   g1111(.A1(new_n270_), .A2(new_n1399_), .B(new_n1402_), .ZN(new_n1403_));
  AOI21_X1   g1112(.A1(new_n1396_), .A2(new_n1394_), .B(new_n1403_), .ZN(new_n1404_));
  OAI21_X1   g1113(.A1(new_n1404_), .A2(new_n264_), .B(new_n1384_), .ZN(\result[13] ));
  NOR3_X1    g1114(.A1(new_n1147_), .A2(new_n1148_), .A3(new_n315_), .ZN(new_n1406_));
  NAND2_X1   g1115(.A1(new_n1296_), .A2(new_n278_), .ZN(new_n1407_));
  AND3_X2    g1116(.A1(new_n309_), .A2(new_n872_), .A3(new_n874_), .Z(new_n1408_));
  AOI21_X1   g1117(.A1(new_n1408_), .A2(new_n870_), .B(new_n291_), .ZN(new_n1409_));
  NOR4_X1    g1118(.A1(new_n1409_), .A2(new_n1406_), .A3(new_n1407_), .A4(new_n1288_), .ZN(new_n1410_));
  NOR2_X1    g1119(.A1(new_n1410_), .A2(new_n270_), .ZN(new_n1411_));
  INV_X1     g1120(.I(new_n1005_), .ZN(new_n1412_));
  NAND2_X1   g1121(.A1(new_n584_), .A2(new_n284_), .ZN(new_n1413_));
  NAND3_X1   g1122(.A1(new_n309_), .A2(new_n1007_), .A3(new_n1413_), .ZN(new_n1414_));
  NOR3_X1    g1123(.A1(new_n1412_), .A2(new_n1414_), .A3(new_n315_), .ZN(new_n1415_));
  NAND2_X1   g1124(.A1(new_n1294_), .A2(new_n1292_), .ZN(new_n1416_));
  NAND2_X1   g1125(.A1(new_n1336_), .A2(new_n1334_), .ZN(new_n1417_));
  NAND3_X1   g1126(.A1(new_n1416_), .A2(new_n1417_), .A3(new_n278_), .ZN(new_n1418_));
  AOI21_X1   g1127(.A1(new_n761_), .A2(new_n763_), .B(new_n291_), .ZN(new_n1419_));
  NOR4_X1    g1128(.A1(new_n1418_), .A2(new_n270_), .A3(new_n1415_), .A4(new_n1419_), .ZN(new_n1420_));
  NOR3_X1    g1129(.A1(new_n1411_), .A2(new_n1420_), .A3(\shift[5] ), .ZN(new_n1421_));
  NAND2_X1   g1130(.A1(new_n860_), .A2(new_n859_), .ZN(new_n1422_));
  INV_X1     g1131(.I(new_n864_), .ZN(new_n1423_));
  NOR2_X1    g1132(.A1(new_n1423_), .A2(new_n283_), .ZN(new_n1424_));
  NAND3_X1   g1133(.A1(new_n1424_), .A2(new_n278_), .A3(new_n1422_), .ZN(new_n1425_));
  OAI21_X1   g1134(.A1(new_n890_), .A2(new_n895_), .B(new_n278_), .ZN(new_n1426_));
  NOR2_X1    g1135(.A1(new_n1426_), .A2(new_n886_), .ZN(new_n1427_));
  OAI21_X1   g1136(.A1(new_n839_), .A2(new_n841_), .B(new_n277_), .ZN(new_n1428_));
  NAND4_X1   g1137(.A1(new_n1427_), .A2(new_n270_), .A3(new_n1425_), .A4(new_n1428_), .ZN(new_n1429_));
  NAND3_X1   g1138(.A1(new_n852_), .A2(new_n309_), .A3(new_n853_), .ZN(new_n1430_));
  NAND3_X1   g1139(.A1(new_n1309_), .A2(new_n1430_), .A3(new_n278_), .ZN(new_n1431_));
  AOI21_X1   g1140(.A1(new_n785_), .A2(new_n781_), .B(new_n291_), .ZN(new_n1432_));
  NOR3_X1    g1141(.A1(new_n1431_), .A2(new_n1432_), .A3(new_n1312_), .ZN(new_n1433_));
  NAND2_X1   g1142(.A1(new_n1433_), .A2(\shift[4] ), .ZN(new_n1434_));
  NAND3_X1   g1143(.A1(new_n1434_), .A2(new_n1429_), .A3(new_n265_), .ZN(new_n1435_));
  OAI21_X1   g1144(.A1(new_n1421_), .A2(new_n1435_), .B(new_n264_), .ZN(new_n1436_));
  AOI21_X1   g1145(.A1(new_n959_), .A2(new_n954_), .B(new_n315_), .ZN(new_n1437_));
  OAI21_X1   g1146(.A1(new_n920_), .A2(new_n924_), .B(new_n277_), .ZN(new_n1438_));
  NAND4_X1   g1147(.A1(new_n1317_), .A2(new_n950_), .A3(new_n1438_), .A4(new_n1437_), .ZN(new_n1439_));
  OAI21_X1   g1148(.A1(new_n817_), .A2(new_n820_), .B(new_n278_), .ZN(new_n1440_));
  AND2_X2    g1149(.A1(new_n309_), .A2(new_n942_), .Z(new_n1441_));
  AOI21_X1   g1150(.A1(new_n1441_), .A2(new_n941_), .B(new_n291_), .ZN(new_n1442_));
  NOR4_X1    g1151(.A1(new_n1442_), .A2(new_n816_), .A3(new_n1323_), .A4(new_n1440_), .ZN(new_n1443_));
  INV_X1     g1152(.I(new_n1443_), .ZN(new_n1444_));
  OAI21_X1   g1153(.A1(new_n1444_), .A2(\shift[4] ), .B(new_n1439_), .ZN(new_n1445_));
  NOR3_X1    g1154(.A1(new_n1443_), .A2(new_n1439_), .A3(\shift[4] ), .ZN(new_n1446_));
  NOR2_X1    g1155(.A1(new_n1446_), .A2(\shift[5] ), .ZN(new_n1447_));
  NAND3_X1   g1156(.A1(new_n1329_), .A2(new_n278_), .A3(new_n1200_), .ZN(new_n1448_));
  AOI21_X1   g1157(.A1(new_n1331_), .A2(new_n1014_), .B(new_n291_), .ZN(new_n1449_));
  OR2_X2     g1158(.A1(new_n1338_), .A2(new_n1449_), .Z(new_n1450_));
  OAI21_X1   g1159(.A1(new_n1450_), .A2(new_n1448_), .B(\shift[4] ), .ZN(new_n1451_));
  NAND2_X1   g1160(.A1(new_n981_), .A2(new_n277_), .ZN(new_n1452_));
  NAND2_X1   g1161(.A1(new_n1343_), .A2(new_n1452_), .ZN(new_n1453_));
  NOR4_X1    g1162(.A1(new_n1453_), .A2(\shift[5] ), .A3(new_n441_), .A4(new_n908_), .ZN(new_n1454_));
  NAND2_X1   g1163(.A1(new_n1451_), .A2(new_n1454_), .ZN(new_n1455_));
  AOI21_X1   g1164(.A1(new_n1447_), .A2(new_n1445_), .B(new_n1455_), .ZN(new_n1456_));
  OAI21_X1   g1165(.A1(new_n1456_), .A2(new_n264_), .B(new_n1436_), .ZN(\result[15] ));
  NAND4_X1   g1166(.A1(new_n272_), .A2(new_n273_), .A3(new_n267_), .A4(new_n265_), .ZN(new_n1458_));
  NAND2_X1   g1167(.A1(new_n1458_), .A2(new_n264_), .ZN(new_n1459_));
  NOR4_X1    g1168(.A1(new_n287_), .A2(\shift[4] ), .A3(new_n277_), .A4(new_n315_), .ZN(new_n1460_));
  NOR4_X1    g1169(.A1(new_n1460_), .A2(new_n709_), .A3(new_n680_), .A4(new_n716_), .ZN(new_n1461_));
  OAI21_X1   g1170(.A1(new_n1461_), .A2(new_n264_), .B(new_n1459_), .ZN(\result[16] ));
  NAND4_X1   g1171(.A1(new_n566_), .A2(new_n578_), .A3(new_n591_), .A4(new_n603_), .ZN(new_n1463_));
  OAI21_X1   g1172(.A1(\shift[4] ), .A2(new_n1463_), .B(new_n379_), .ZN(new_n1464_));
  NOR3_X1    g1173(.A1(new_n630_), .A2(new_n379_), .A3(\shift[4] ), .ZN(new_n1465_));
  NOR2_X1    g1174(.A1(new_n1465_), .A2(\shift[5] ), .ZN(new_n1466_));
  NAND2_X1   g1175(.A1(new_n336_), .A2(new_n270_), .ZN(new_n1467_));
  NOR4_X1    g1176(.A1(new_n393_), .A2(new_n1378_), .A3(new_n1071_), .A4(new_n403_), .ZN(new_n1468_));
  AOI21_X1   g1177(.A1(new_n1468_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1469_));
  NAND2_X1   g1178(.A1(new_n1469_), .A2(new_n1467_), .ZN(new_n1470_));
  AOI21_X1   g1179(.A1(new_n1466_), .A2(new_n1464_), .B(new_n1470_), .ZN(new_n1471_));
  INV_X1     g1180(.I(new_n443_), .ZN(new_n1472_));
  NOR2_X1    g1181(.A1(new_n442_), .A2(\shift[0] ), .ZN(new_n1473_));
  NAND3_X1   g1182(.A1(new_n818_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n1474_));
  NAND2_X1   g1183(.A1(new_n1473_), .A2(new_n1474_), .ZN(new_n1475_));
  NAND2_X1   g1184(.A1(new_n1475_), .A2(new_n1472_), .ZN(new_n1476_));
  NOR3_X1    g1185(.A1(new_n283_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n1477_));
  NAND2_X1   g1186(.A1(new_n1476_), .A2(new_n1477_), .ZN(new_n1478_));
  NAND3_X1   g1187(.A1(new_n439_), .A2(new_n1478_), .A3(new_n440_), .ZN(new_n1479_));
  NAND2_X1   g1188(.A1(new_n461_), .A2(new_n473_), .ZN(new_n1480_));
  NOR2_X1    g1189(.A1(new_n1480_), .A2(new_n1479_), .ZN(new_n1481_));
  NOR2_X1    g1190(.A1(new_n519_), .A2(new_n270_), .ZN(new_n1482_));
  NOR3_X1    g1191(.A1(new_n1482_), .A2(\shift[5] ), .A3(new_n1481_), .ZN(new_n1483_));
  NOR4_X1    g1192(.A1(new_n641_), .A2(new_n655_), .A3(new_n665_), .A4(new_n675_), .ZN(new_n1484_));
  NOR3_X1    g1193(.A1(new_n279_), .A2(\a[34] ), .A3(\shift[1] ), .ZN(new_n1485_));
  NOR3_X1    g1194(.A1(new_n1485_), .A2(\shift[0] ), .A3(new_n681_), .ZN(new_n1486_));
  NOR2_X1    g1195(.A1(new_n1486_), .A2(new_n682_), .ZN(new_n1487_));
  NOR2_X1    g1196(.A1(new_n689_), .A2(new_n690_), .ZN(new_n1488_));
  NAND2_X1   g1197(.A1(new_n1488_), .A2(new_n309_), .ZN(new_n1489_));
  OAI21_X1   g1198(.A1(new_n1487_), .A2(new_n1489_), .B(new_n277_), .ZN(new_n1490_));
  NAND2_X1   g1199(.A1(new_n1259_), .A2(new_n1260_), .ZN(new_n1491_));
  NAND4_X1   g1200(.A1(new_n1491_), .A2(new_n1490_), .A3(new_n265_), .A4(new_n440_), .ZN(new_n1492_));
  INV_X1     g1201(.I(new_n1492_), .ZN(new_n1493_));
  OAI21_X1   g1202(.A1(new_n1484_), .A2(new_n270_), .B(new_n1493_), .ZN(new_n1494_));
  OAI21_X1   g1203(.A1(new_n1483_), .A2(new_n1494_), .B(\shift[6] ), .ZN(new_n1495_));
  OAI21_X1   g1204(.A1(new_n1471_), .A2(\shift[6] ), .B(new_n1495_), .ZN(\result[17] ));
  NOR4_X1    g1205(.A1(new_n270_), .A2(\shift[2] ), .A3(\shift[3] ), .A4(\shift[5] ), .ZN(new_n1497_));
  OAI21_X1   g1206(.A1(new_n264_), .A2(new_n1497_), .B(new_n1459_), .ZN(\result[18] ));
  INV_X1     g1207(.I(new_n1039_), .ZN(new_n1499_));
  OAI21_X1   g1208(.A1(new_n1499_), .A2(\shift[4] ), .B(new_n765_), .ZN(new_n1500_));
  NOR3_X1    g1209(.A1(new_n765_), .A2(new_n1039_), .A3(\shift[4] ), .ZN(new_n1501_));
  NOR2_X1    g1210(.A1(new_n1501_), .A2(\shift[5] ), .ZN(new_n1502_));
  INV_X1     g1211(.I(new_n866_), .ZN(new_n1503_));
  NOR4_X1    g1212(.A1(new_n1503_), .A2(new_n876_), .A3(new_n886_), .A4(new_n896_), .ZN(new_n1504_));
  NAND4_X1   g1213(.A1(new_n1504_), .A2(\shift[4] ), .A3(new_n856_), .A4(new_n265_), .ZN(new_n1505_));
  AOI21_X1   g1214(.A1(new_n1502_), .A2(new_n1500_), .B(new_n1505_), .ZN(new_n1506_));
  NOR3_X1    g1215(.A1(new_n807_), .A2(new_n787_), .A3(new_n270_), .ZN(new_n1507_));
  AOI21_X1   g1216(.A1(new_n1173_), .A2(new_n931_), .B(new_n291_), .ZN(new_n1508_));
  NAND2_X1   g1217(.A1(new_n943_), .A2(new_n278_), .ZN(new_n1509_));
  INV_X1     g1218(.I(new_n950_), .ZN(new_n1510_));
  NOR4_X1    g1219(.A1(new_n1508_), .A2(new_n1509_), .A3(new_n1510_), .A4(new_n1178_), .ZN(new_n1511_));
  NOR2_X1    g1220(.A1(new_n1511_), .A2(new_n270_), .ZN(new_n1512_));
  NOR3_X1    g1221(.A1(new_n1512_), .A2(new_n1507_), .A3(\shift[5] ), .ZN(new_n1513_));
  NAND4_X1   g1222(.A1(new_n926_), .A2(new_n1000_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1514_));
  OAI21_X1   g1223(.A1(new_n1513_), .A2(new_n1514_), .B(\shift[6] ), .ZN(new_n1515_));
  OAI21_X1   g1224(.A1(new_n1506_), .A2(\shift[6] ), .B(new_n1515_), .ZN(\result[19] ));
  NOR3_X1    g1225(.A1(new_n267_), .A2(\shift[4] ), .A3(new_n265_), .ZN(new_n1517_));
  OAI21_X1   g1226(.A1(new_n264_), .A2(new_n1517_), .B(new_n1459_), .ZN(\result[20] ));
  INV_X1     g1227(.I(new_n1128_), .ZN(new_n1519_));
  OAI21_X1   g1228(.A1(new_n1519_), .A2(\shift[4] ), .B(new_n1063_), .ZN(new_n1520_));
  NOR3_X1    g1229(.A1(new_n1128_), .A2(new_n1063_), .A3(\shift[4] ), .ZN(new_n1521_));
  NOR2_X1    g1230(.A1(new_n1521_), .A2(\shift[5] ), .ZN(new_n1522_));
  NAND2_X1   g1231(.A1(new_n1053_), .A2(new_n270_), .ZN(new_n1523_));
  NOR2_X1    g1232(.A1(new_n1071_), .A2(new_n1077_), .ZN(new_n1524_));
  NOR2_X1    g1233(.A1(new_n1078_), .A2(new_n1079_), .ZN(new_n1525_));
  NAND3_X1   g1234(.A1(new_n1525_), .A2(new_n1524_), .A3(\shift[4] ), .ZN(new_n1526_));
  NAND3_X1   g1235(.A1(new_n1523_), .A2(new_n1526_), .A3(new_n265_), .ZN(new_n1527_));
  AOI21_X1   g1236(.A1(new_n1522_), .A2(new_n1520_), .B(new_n1527_), .ZN(new_n1528_));
  AOI21_X1   g1237(.A1(new_n389_), .A2(new_n392_), .B(new_n315_), .ZN(new_n1529_));
  OAI21_X1   g1238(.A1(new_n1251_), .A2(new_n1252_), .B(new_n277_), .ZN(new_n1530_));
  NAND3_X1   g1239(.A1(new_n1476_), .A2(new_n1477_), .A3(new_n278_), .ZN(new_n1531_));
  NAND4_X1   g1240(.A1(new_n473_), .A2(new_n1529_), .A3(new_n1530_), .A4(new_n1531_), .ZN(new_n1532_));
  NOR2_X1    g1241(.A1(new_n1532_), .A2(new_n265_), .ZN(new_n1533_));
  OAI21_X1   g1242(.A1(new_n1101_), .A2(new_n265_), .B(new_n270_), .ZN(new_n1534_));
  NOR2_X1    g1243(.A1(new_n1533_), .A2(new_n1534_), .ZN(new_n1535_));
  NAND4_X1   g1244(.A1(new_n1120_), .A2(new_n270_), .A3(\shift[5] ), .A4(new_n1105_), .ZN(new_n1536_));
  OAI21_X1   g1245(.A1(new_n1535_), .A2(new_n1536_), .B(\shift[6] ), .ZN(new_n1537_));
  OAI21_X1   g1246(.A1(new_n1528_), .A2(\shift[6] ), .B(new_n1537_), .ZN(\result[21] ));
  NOR3_X1    g1247(.A1(new_n267_), .A2(\shift[4] ), .A3(new_n265_), .ZN(new_n1539_));
  OAI21_X1   g1248(.A1(new_n264_), .A2(new_n1539_), .B(new_n1459_), .ZN(\result[22] ));
  NAND2_X1   g1249(.A1(new_n270_), .A2(new_n265_), .ZN(new_n1541_));
  NAND2_X1   g1250(.A1(\shift[4] ), .A2(\shift[5] ), .ZN(new_n1542_));
  NOR3_X1    g1251(.A1(new_n680_), .A2(new_n1541_), .A3(new_n1542_), .ZN(new_n1543_));
  NAND3_X1   g1252(.A1(new_n1196_), .A2(new_n1162_), .A3(new_n1543_), .ZN(new_n1544_));
  INV_X1     g1253(.I(new_n1143_), .ZN(new_n1545_));
  INV_X1     g1254(.I(new_n1296_), .ZN(new_n1546_));
  NOR2_X1    g1255(.A1(new_n1412_), .A2(new_n1414_), .ZN(new_n1547_));
  NOR3_X1    g1256(.A1(new_n1546_), .A2(new_n1547_), .A3(new_n315_), .ZN(new_n1548_));
  NAND4_X1   g1257(.A1(new_n1548_), .A2(\shift[4] ), .A3(new_n1149_), .A4(new_n1291_), .ZN(new_n1549_));
  OAI21_X1   g1258(.A1(new_n1545_), .A2(\shift[4] ), .B(new_n1549_), .ZN(new_n1550_));
  OAI21_X1   g1259(.A1(new_n1550_), .A2(new_n1544_), .B(new_n264_), .ZN(new_n1551_));
  NOR2_X1    g1260(.A1(new_n834_), .A2(new_n315_), .ZN(new_n1552_));
  NAND4_X1   g1261(.A1(new_n1552_), .A2(new_n806_), .A3(new_n1166_), .A4(new_n1165_), .ZN(new_n1553_));
  OAI21_X1   g1262(.A1(new_n1553_), .A2(\shift[4] ), .B(new_n265_), .ZN(new_n1554_));
  NAND2_X1   g1263(.A1(new_n1205_), .A2(\shift[4] ), .ZN(new_n1555_));
  NOR2_X1    g1264(.A1(new_n1553_), .A2(\shift[4] ), .ZN(new_n1556_));
  OAI21_X1   g1265(.A1(new_n1555_), .A2(new_n1556_), .B(\shift[5] ), .ZN(new_n1557_));
  NOR2_X1    g1266(.A1(new_n1179_), .A2(new_n1178_), .ZN(new_n1558_));
  INV_X1     g1267(.I(new_n1183_), .ZN(new_n1559_));
  INV_X1     g1268(.I(new_n1184_), .ZN(new_n1560_));
  NAND4_X1   g1269(.A1(new_n1559_), .A2(new_n265_), .A3(new_n1558_), .A4(new_n1560_), .ZN(new_n1561_));
  NAND4_X1   g1270(.A1(new_n1171_), .A2(\shift[5] ), .A3(new_n1174_), .A4(new_n1170_), .ZN(new_n1562_));
  NAND3_X1   g1271(.A1(new_n1561_), .A2(new_n1562_), .A3(new_n679_), .ZN(new_n1563_));
  AOI21_X1   g1272(.A1(new_n1557_), .A2(new_n1554_), .B(new_n1563_), .ZN(new_n1564_));
  OAI21_X1   g1273(.A1(new_n1564_), .A2(new_n264_), .B(new_n1551_), .ZN(\result[23] ));
  NAND4_X1   g1274(.A1(new_n1543_), .A2(new_n266_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n1566_));
  NAND2_X1   g1275(.A1(new_n1566_), .A2(new_n264_), .ZN(new_n1567_));
  NOR3_X1    g1276(.A1(new_n287_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n1568_));
  OR2_X2     g1277(.A1(new_n1568_), .A2(new_n265_), .Z(new_n1569_));
  AOI21_X1   g1278(.A1(new_n1568_), .A2(new_n265_), .B(new_n713_), .ZN(new_n1570_));
  NAND2_X1   g1279(.A1(new_n266_), .A2(\shift[5] ), .ZN(new_n1571_));
  NAND3_X1   g1280(.A1(new_n1134_), .A2(new_n679_), .A3(new_n1571_), .ZN(new_n1572_));
  AOI21_X1   g1281(.A1(new_n1569_), .A2(new_n1570_), .B(new_n1572_), .ZN(new_n1573_));
  OAI21_X1   g1282(.A1(new_n1573_), .A2(new_n264_), .B(new_n1567_), .ZN(\result[24] ));
  NAND3_X1   g1283(.A1(new_n1232_), .A2(new_n1269_), .A3(new_n1543_), .ZN(new_n1575_));
  INV_X1     g1284(.I(new_n1216_), .ZN(new_n1576_));
  OAI21_X1   g1285(.A1(new_n1576_), .A2(\shift[4] ), .B(new_n1226_), .ZN(new_n1577_));
  OAI21_X1   g1286(.A1(new_n1577_), .A2(new_n1575_), .B(new_n264_), .ZN(new_n1578_));
  AOI21_X1   g1287(.A1(new_n412_), .A2(new_n415_), .B(new_n315_), .ZN(new_n1579_));
  NAND4_X1   g1288(.A1(new_n1531_), .A2(new_n1579_), .A3(new_n1241_), .A4(new_n1242_), .ZN(new_n1580_));
  OAI21_X1   g1289(.A1(new_n1580_), .A2(\shift[4] ), .B(new_n265_), .ZN(new_n1581_));
  INV_X1     g1290(.I(new_n1270_), .ZN(new_n1582_));
  NAND4_X1   g1291(.A1(new_n1582_), .A2(\shift[4] ), .A3(new_n1271_), .A4(new_n1273_), .ZN(new_n1583_));
  NOR2_X1    g1292(.A1(new_n1580_), .A2(\shift[4] ), .ZN(new_n1584_));
  OAI21_X1   g1293(.A1(new_n1584_), .A2(new_n1583_), .B(\shift[5] ), .ZN(new_n1585_));
  NAND2_X1   g1294(.A1(new_n1256_), .A2(new_n265_), .ZN(new_n1586_));
  AOI21_X1   g1295(.A1(new_n1248_), .A2(\shift[5] ), .B(new_n680_), .ZN(new_n1587_));
  NAND2_X1   g1296(.A1(new_n1586_), .A2(new_n1587_), .ZN(new_n1588_));
  AOI21_X1   g1297(.A1(new_n1581_), .A2(new_n1585_), .B(new_n1588_), .ZN(new_n1589_));
  OAI21_X1   g1298(.A1(new_n1589_), .A2(new_n264_), .B(new_n1578_), .ZN(\result[25] ));
  NOR2_X1    g1299(.A1(new_n709_), .A2(new_n265_), .ZN(new_n1591_));
  NOR3_X1    g1300(.A1(new_n1279_), .A2(new_n713_), .A3(new_n1591_), .ZN(new_n1592_));
  OAI21_X1   g1301(.A1(new_n1592_), .A2(new_n1572_), .B(\shift[6] ), .ZN(new_n1593_));
  NAND2_X1   g1302(.A1(new_n1593_), .A2(new_n1459_), .ZN(\result[26] ));
  NOR3_X1    g1303(.A1(new_n736_), .A2(new_n315_), .A3(new_n1193_), .ZN(new_n1595_));
  AOI21_X1   g1304(.A1(new_n277_), .A2(new_n1296_), .B(new_n1415_), .ZN(new_n1596_));
  OAI21_X1   g1305(.A1(new_n988_), .A2(new_n984_), .B(new_n278_), .ZN(new_n1597_));
  NOR4_X1    g1306(.A1(new_n1195_), .A2(new_n1338_), .A3(new_n1597_), .A4(new_n1337_), .ZN(new_n1598_));
  AOI22_X1   g1307(.A1(new_n1595_), .A2(new_n1596_), .B1(new_n1598_), .B2(new_n270_), .ZN(new_n1599_));
  NOR3_X1    g1308(.A1(new_n1299_), .A2(new_n1598_), .A3(\shift[4] ), .ZN(new_n1600_));
  NOR3_X1    g1309(.A1(new_n1599_), .A2(new_n1600_), .A3(\shift[5] ), .ZN(new_n1601_));
  INV_X1     g1310(.I(new_n1289_), .ZN(new_n1602_));
  AOI21_X1   g1311(.A1(new_n1306_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1603_));
  OAI21_X1   g1312(.A1(\shift[4] ), .A2(new_n1602_), .B(new_n1603_), .ZN(new_n1604_));
  OAI21_X1   g1313(.A1(new_n1601_), .A2(new_n1604_), .B(new_n264_), .ZN(new_n1605_));
  NAND3_X1   g1314(.A1(new_n786_), .A2(new_n278_), .A3(new_n1309_), .ZN(new_n1606_));
  OAI21_X1   g1315(.A1(new_n817_), .A2(new_n820_), .B(new_n277_), .ZN(new_n1607_));
  INV_X1     g1316(.I(new_n1312_), .ZN(new_n1608_));
  NAND2_X1   g1317(.A1(new_n1608_), .A2(new_n1607_), .ZN(new_n1609_));
  NOR4_X1    g1318(.A1(new_n1609_), .A2(new_n1606_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1610_));
  AOI21_X1   g1319(.A1(new_n1313_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n1611_));
  NOR2_X1    g1320(.A1(new_n1341_), .A2(new_n1204_), .ZN(new_n1612_));
  AOI22_X1   g1321(.A1(new_n914_), .A2(new_n278_), .B1(new_n1200_), .B2(new_n277_), .ZN(new_n1613_));
  AOI21_X1   g1322(.A1(new_n1612_), .A2(new_n1613_), .B(new_n265_), .ZN(new_n1614_));
  NOR4_X1    g1323(.A1(new_n1611_), .A2(new_n1614_), .A3(new_n1345_), .A4(new_n1610_), .ZN(new_n1615_));
  NAND2_X1   g1324(.A1(new_n1324_), .A2(new_n265_), .ZN(new_n1616_));
  NAND4_X1   g1325(.A1(new_n1318_), .A2(\shift[5] ), .A3(new_n1317_), .A4(new_n1170_), .ZN(new_n1617_));
  NAND3_X1   g1326(.A1(new_n1616_), .A2(new_n679_), .A3(new_n1617_), .ZN(new_n1618_));
  OAI21_X1   g1327(.A1(new_n1615_), .A2(new_n1618_), .B(\shift[6] ), .ZN(new_n1619_));
  NAND2_X1   g1328(.A1(new_n1605_), .A2(new_n1619_), .ZN(\result[27] ));
  NAND2_X1   g1329(.A1(new_n1350_), .A2(\shift[5] ), .ZN(new_n1621_));
  AOI21_X1   g1330(.A1(new_n1349_), .A2(new_n265_), .B(new_n713_), .ZN(new_n1622_));
  AOI21_X1   g1331(.A1(new_n1621_), .A2(new_n1622_), .B(new_n1572_), .ZN(new_n1623_));
  OAI21_X1   g1332(.A1(new_n1623_), .A2(new_n264_), .B(new_n1459_), .ZN(\result[28] ));
  NOR2_X1    g1333(.A1(new_n357_), .A2(new_n291_), .ZN(new_n1625_));
  OAI21_X1   g1334(.A1(new_n626_), .A2(new_n628_), .B(new_n278_), .ZN(new_n1626_));
  NOR2_X1    g1335(.A1(new_n1625_), .A2(new_n1626_), .ZN(new_n1627_));
  NOR2_X1    g1336(.A1(new_n561_), .A2(new_n565_), .ZN(new_n1628_));
  OAI21_X1   g1337(.A1(new_n1628_), .A2(new_n1218_), .B(new_n278_), .ZN(new_n1629_));
  AOI22_X1   g1338(.A1(new_n1399_), .A2(new_n270_), .B1(new_n1627_), .B2(new_n1629_), .ZN(new_n1630_));
  NOR3_X1    g1339(.A1(new_n1399_), .A2(new_n1370_), .A3(\shift[4] ), .ZN(new_n1631_));
  NOR3_X1    g1340(.A1(new_n1630_), .A2(new_n1631_), .A3(\shift[5] ), .ZN(new_n1632_));
  NAND2_X1   g1341(.A1(new_n1362_), .A2(new_n270_), .ZN(new_n1633_));
  INV_X1     g1342(.I(new_n395_), .ZN(new_n1634_));
  NOR2_X1    g1343(.A1(new_n394_), .A2(\shift[0] ), .ZN(new_n1635_));
  INV_X1     g1344(.I(\a[94] ), .ZN(new_n1636_));
  NAND3_X1   g1345(.A1(new_n1636_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n1637_));
  NAND2_X1   g1346(.A1(new_n1635_), .A2(new_n1637_), .ZN(new_n1638_));
  NAND2_X1   g1347(.A1(new_n1638_), .A2(new_n1634_), .ZN(new_n1639_));
  NOR3_X1    g1348(.A1(new_n283_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n1640_));
  AOI21_X1   g1349(.A1(new_n1639_), .A2(new_n1640_), .B(new_n291_), .ZN(new_n1641_));
  NOR4_X1    g1350(.A1(new_n325_), .A2(new_n1641_), .A3(new_n1231_), .A4(new_n1374_), .ZN(new_n1642_));
  AOI21_X1   g1351(.A1(new_n1642_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1643_));
  NAND2_X1   g1352(.A1(new_n1643_), .A2(new_n1633_), .ZN(new_n1644_));
  OAI21_X1   g1353(.A1(new_n1632_), .A2(new_n1644_), .B(new_n264_), .ZN(new_n1645_));
  AOI21_X1   g1354(.A1(new_n424_), .A2(new_n427_), .B(new_n315_), .ZN(new_n1646_));
  NAND2_X1   g1355(.A1(new_n1646_), .A2(new_n416_), .ZN(new_n1647_));
  NAND2_X1   g1356(.A1(new_n1381_), .A2(new_n1242_), .ZN(new_n1648_));
  NOR4_X1    g1357(.A1(new_n1647_), .A2(new_n1648_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1649_));
  NOR3_X1    g1358(.A1(new_n1084_), .A2(new_n315_), .A3(new_n1086_), .ZN(new_n1650_));
  AOI21_X1   g1359(.A1(new_n1476_), .A2(new_n1477_), .B(new_n291_), .ZN(new_n1651_));
  NOR4_X1    g1360(.A1(new_n1378_), .A2(new_n1650_), .A3(new_n1651_), .A4(new_n1379_), .ZN(new_n1652_));
  AOI21_X1   g1361(.A1(new_n1652_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n1653_));
  XOR2_X1    g1362(.A1(new_n643_), .A2(new_n648_), .Z(new_n1654_));
  INV_X1     g1363(.I(new_n654_), .ZN(new_n1655_));
  AOI21_X1   g1364(.A1(new_n1654_), .A2(new_n1655_), .B(new_n291_), .ZN(new_n1656_));
  NAND2_X1   g1365(.A1(new_n1273_), .A2(new_n440_), .ZN(new_n1657_));
  OAI21_X1   g1366(.A1(new_n1657_), .A2(new_n1656_), .B(\shift[5] ), .ZN(new_n1658_));
  NAND2_X1   g1367(.A1(new_n1658_), .A2(new_n1401_), .ZN(new_n1659_));
  NOR3_X1    g1368(.A1(new_n1659_), .A2(new_n1653_), .A3(new_n1649_), .ZN(new_n1660_));
  NAND2_X1   g1369(.A1(new_n1392_), .A2(new_n265_), .ZN(new_n1661_));
  NOR2_X1    g1370(.A1(new_n513_), .A2(new_n517_), .ZN(new_n1662_));
  NOR3_X1    g1371(.A1(new_n1662_), .A2(new_n1246_), .A3(new_n315_), .ZN(new_n1663_));
  AOI21_X1   g1372(.A1(new_n1491_), .A2(new_n277_), .B(new_n1247_), .ZN(new_n1664_));
  NAND3_X1   g1373(.A1(new_n1664_), .A2(\shift[5] ), .A3(new_n1663_), .ZN(new_n1665_));
  NAND3_X1   g1374(.A1(new_n1661_), .A2(new_n1665_), .A3(new_n679_), .ZN(new_n1666_));
  OAI21_X1   g1375(.A1(new_n1660_), .A2(new_n1666_), .B(\shift[6] ), .ZN(new_n1667_));
  NAND2_X1   g1376(.A1(new_n1645_), .A2(new_n1667_), .ZN(\result[29] ));
  NOR2_X1    g1377(.A1(new_n1033_), .A2(new_n1037_), .ZN(new_n1669_));
  NOR3_X1    g1378(.A1(new_n1193_), .A2(new_n1669_), .A3(new_n315_), .ZN(new_n1670_));
  NOR2_X1    g1379(.A1(new_n1419_), .A2(new_n1415_), .ZN(new_n1671_));
  NAND2_X1   g1380(.A1(new_n1200_), .A2(new_n278_), .ZN(new_n1672_));
  NOR4_X1    g1381(.A1(new_n1672_), .A2(new_n1338_), .A3(new_n1449_), .A4(new_n989_), .ZN(new_n1673_));
  AOI22_X1   g1382(.A1(new_n1673_), .A2(new_n270_), .B1(new_n1671_), .B2(new_n1670_), .ZN(new_n1674_));
  OAI21_X1   g1383(.A1(new_n736_), .A2(new_n291_), .B(new_n1298_), .ZN(new_n1675_));
  NOR4_X1    g1384(.A1(new_n1673_), .A2(new_n1675_), .A3(\shift[4] ), .A4(new_n1418_), .ZN(new_n1676_));
  NOR3_X1    g1385(.A1(new_n1674_), .A2(new_n1676_), .A3(\shift[5] ), .ZN(new_n1677_));
  NAND2_X1   g1386(.A1(new_n1410_), .A2(new_n270_), .ZN(new_n1678_));
  INV_X1     g1387(.I(new_n1428_), .ZN(new_n1679_));
  NOR4_X1    g1388(.A1(new_n1679_), .A2(new_n886_), .A3(new_n1305_), .A4(new_n1426_), .ZN(new_n1680_));
  NAND2_X1   g1389(.A1(new_n1680_), .A2(\shift[4] ), .ZN(new_n1681_));
  NAND3_X1   g1390(.A1(new_n1681_), .A2(new_n1678_), .A3(new_n265_), .ZN(new_n1682_));
  OAI21_X1   g1391(.A1(new_n1677_), .A2(new_n1682_), .B(new_n264_), .ZN(new_n1683_));
  OAI21_X1   g1392(.A1(new_n811_), .A2(new_n813_), .B(new_n277_), .ZN(new_n1684_));
  NAND2_X1   g1393(.A1(new_n1608_), .A2(new_n1684_), .ZN(new_n1685_));
  NOR4_X1    g1394(.A1(new_n1685_), .A2(\shift[4] ), .A3(new_n265_), .A4(new_n1431_), .ZN(new_n1686_));
  AOI21_X1   g1395(.A1(new_n1433_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n1687_));
  NOR2_X1    g1396(.A1(new_n908_), .A2(new_n441_), .ZN(new_n1688_));
  AOI22_X1   g1397(.A1(new_n914_), .A2(new_n278_), .B1(new_n981_), .B2(new_n277_), .ZN(new_n1689_));
  AOI21_X1   g1398(.A1(new_n1688_), .A2(new_n1689_), .B(new_n265_), .ZN(new_n1690_));
  NOR4_X1    g1399(.A1(new_n1687_), .A2(new_n1690_), .A3(new_n1454_), .A4(new_n1686_), .ZN(new_n1691_));
  NAND2_X1   g1400(.A1(new_n1443_), .A2(new_n265_), .ZN(new_n1692_));
  NOR3_X1    g1401(.A1(new_n1321_), .A2(new_n1182_), .A3(new_n315_), .ZN(new_n1693_));
  NAND4_X1   g1402(.A1(new_n1693_), .A2(\shift[5] ), .A3(new_n1317_), .A4(new_n1438_), .ZN(new_n1694_));
  NAND3_X1   g1403(.A1(new_n1692_), .A2(new_n679_), .A3(new_n1694_), .ZN(new_n1695_));
  OAI21_X1   g1404(.A1(new_n1691_), .A2(new_n1695_), .B(\shift[6] ), .ZN(new_n1696_));
  NAND2_X1   g1405(.A1(new_n1683_), .A2(new_n1696_), .ZN(\result[31] ));
  OAI21_X1   g1406(.A1(new_n1132_), .A2(new_n1135_), .B(new_n264_), .ZN(new_n1698_));
  NAND2_X1   g1407(.A1(new_n287_), .A2(new_n278_), .ZN(new_n1699_));
  AOI21_X1   g1408(.A1(new_n1699_), .A2(new_n266_), .B(new_n270_), .ZN(new_n1700_));
  NOR3_X1    g1409(.A1(new_n1700_), .A2(new_n1133_), .A3(new_n1280_), .ZN(new_n1701_));
  OAI21_X1   g1410(.A1(new_n1701_), .A2(new_n264_), .B(new_n1698_), .ZN(\result[32] ));
  AOI21_X1   g1411(.A1(new_n1484_), .A2(new_n270_), .B(new_n630_), .ZN(new_n1703_));
  NOR3_X1    g1412(.A1(new_n1484_), .A2(new_n1463_), .A3(\shift[4] ), .ZN(new_n1704_));
  NOR3_X1    g1413(.A1(new_n1703_), .A2(new_n1704_), .A3(\shift[5] ), .ZN(new_n1705_));
  INV_X1     g1414(.I(new_n379_), .ZN(new_n1706_));
  NAND4_X1   g1415(.A1(new_n1706_), .A2(\shift[4] ), .A3(new_n265_), .A4(new_n336_), .ZN(new_n1707_));
  OAI21_X1   g1416(.A1(new_n1705_), .A2(new_n1707_), .B(new_n264_), .ZN(new_n1708_));
  OAI21_X1   g1417(.A1(new_n1084_), .A2(new_n1086_), .B(new_n277_), .ZN(new_n1709_));
  AOI21_X1   g1418(.A1(new_n1639_), .A2(new_n1640_), .B(new_n315_), .ZN(new_n1710_));
  NAND4_X1   g1419(.A1(new_n1709_), .A2(new_n1710_), .A3(new_n416_), .A4(new_n428_), .ZN(new_n1711_));
  NOR3_X1    g1420(.A1(new_n1711_), .A2(\shift[4] ), .A3(new_n265_), .ZN(new_n1712_));
  AOI21_X1   g1421(.A1(new_n1468_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n1713_));
  OAI21_X1   g1422(.A1(new_n692_), .A2(new_n702_), .B(\shift[5] ), .ZN(new_n1714_));
  NAND2_X1   g1423(.A1(new_n1492_), .A2(new_n1714_), .ZN(new_n1715_));
  NOR3_X1    g1424(.A1(new_n1713_), .A2(new_n1712_), .A3(new_n1715_), .ZN(new_n1716_));
  NAND2_X1   g1425(.A1(new_n519_), .A2(new_n270_), .ZN(new_n1717_));
  NAND3_X1   g1426(.A1(new_n1717_), .A2(new_n474_), .A3(new_n679_), .ZN(new_n1718_));
  OAI21_X1   g1427(.A1(new_n1716_), .A2(new_n1718_), .B(\shift[6] ), .ZN(new_n1719_));
  NAND2_X1   g1428(.A1(new_n1708_), .A2(new_n1719_), .ZN(\result[33] ));
  NOR2_X1    g1429(.A1(new_n1592_), .A2(new_n717_), .ZN(new_n1721_));
  OAI21_X1   g1430(.A1(new_n1721_), .A2(new_n264_), .B(new_n1698_), .ZN(\result[34] ));
  NAND3_X1   g1431(.A1(new_n1504_), .A2(new_n1000_), .A3(new_n1543_), .ZN(new_n1723_));
  NOR2_X1    g1432(.A1(new_n765_), .A2(new_n265_), .ZN(new_n1724_));
  NOR2_X1    g1433(.A1(new_n1499_), .A2(\shift[5] ), .ZN(new_n1725_));
  NOR3_X1    g1434(.A1(new_n1725_), .A2(new_n1723_), .A3(new_n1724_), .ZN(new_n1726_));
  NOR2_X1    g1435(.A1(new_n1511_), .A2(new_n265_), .ZN(new_n1727_));
  NOR4_X1    g1436(.A1(new_n855_), .A2(new_n265_), .A3(new_n835_), .A4(new_n842_), .ZN(new_n1728_));
  NOR3_X1    g1437(.A1(new_n1727_), .A2(\shift[4] ), .A3(new_n1728_), .ZN(new_n1729_));
  NAND4_X1   g1438(.A1(new_n822_), .A2(new_n926_), .A3(new_n270_), .A4(\shift[5] ), .ZN(new_n1730_));
  OAI21_X1   g1439(.A1(new_n1729_), .A2(new_n1730_), .B(\shift[6] ), .ZN(new_n1731_));
  OAI21_X1   g1440(.A1(\shift[6] ), .A2(new_n1726_), .B(new_n1731_), .ZN(\result[35] ));
  NAND3_X1   g1441(.A1(new_n266_), .A2(\shift[4] ), .A3(new_n265_), .ZN(new_n1733_));
  NAND2_X1   g1442(.A1(new_n1733_), .A2(new_n264_), .ZN(new_n1734_));
  INV_X1     g1443(.I(new_n273_), .ZN(new_n1735_));
  INV_X1     g1444(.I(new_n1044_), .ZN(new_n1736_));
  NOR2_X1    g1445(.A1(new_n1736_), .A2(new_n270_), .ZN(new_n1737_));
  NOR4_X1    g1446(.A1(new_n1737_), .A2(new_n1735_), .A3(\shift[5] ), .A4(new_n266_), .ZN(new_n1738_));
  OAI21_X1   g1447(.A1(new_n1738_), .A2(new_n264_), .B(new_n1734_), .ZN(\result[36] ));
  NOR4_X1    g1448(.A1(new_n1113_), .A2(new_n270_), .A3(new_n1118_), .A4(new_n1119_), .ZN(new_n1740_));
  OAI21_X1   g1449(.A1(new_n1128_), .A2(new_n270_), .B(new_n265_), .ZN(new_n1741_));
  NOR2_X1    g1450(.A1(new_n1741_), .A2(new_n1740_), .ZN(new_n1742_));
  AND4_X2    g1451(.A1(new_n378_), .A2(new_n1055_), .A3(new_n1056_), .A4(new_n1062_), .Z(new_n1743_));
  NAND4_X1   g1452(.A1(new_n1743_), .A2(\shift[4] ), .A3(new_n1053_), .A4(new_n265_), .ZN(new_n1744_));
  OAI21_X1   g1453(.A1(new_n1742_), .A2(new_n1744_), .B(new_n264_), .ZN(new_n1745_));
  INV_X1     g1454(.I(new_n1080_), .ZN(new_n1746_));
  OAI21_X1   g1455(.A1(new_n1746_), .A2(\shift[4] ), .B(new_n1532_), .ZN(new_n1747_));
  NOR3_X1    g1456(.A1(new_n1080_), .A2(new_n1532_), .A3(\shift[4] ), .ZN(new_n1748_));
  NOR2_X1    g1457(.A1(new_n1748_), .A2(\shift[5] ), .ZN(new_n1749_));
  NAND2_X1   g1458(.A1(new_n1105_), .A2(new_n270_), .ZN(new_n1750_));
  AOI21_X1   g1459(.A1(new_n1101_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1751_));
  NAND2_X1   g1460(.A1(new_n1750_), .A2(new_n1751_), .ZN(new_n1752_));
  AOI21_X1   g1461(.A1(new_n1749_), .A2(new_n1747_), .B(new_n1752_), .ZN(new_n1753_));
  OAI21_X1   g1462(.A1(new_n1753_), .A2(new_n264_), .B(new_n1745_), .ZN(\result[37] ));
  NAND2_X1   g1463(.A1(new_n1458_), .A2(\shift[6] ), .ZN(new_n1755_));
  NAND2_X1   g1464(.A1(new_n1755_), .A2(new_n1734_), .ZN(\result[38] ));
  NOR2_X1    g1465(.A1(new_n1192_), .A2(new_n1038_), .ZN(new_n1757_));
  NOR2_X1    g1466(.A1(new_n1194_), .A2(new_n1195_), .ZN(new_n1758_));
  AOI21_X1   g1467(.A1(new_n1758_), .A2(new_n1757_), .B(new_n270_), .ZN(new_n1759_));
  NOR4_X1    g1468(.A1(new_n1201_), .A2(new_n1203_), .A3(new_n270_), .A4(new_n1204_), .ZN(new_n1760_));
  NOR3_X1    g1469(.A1(new_n1759_), .A2(new_n1760_), .A3(\shift[5] ), .ZN(new_n1761_));
  NOR3_X1    g1470(.A1(new_n1146_), .A2(new_n1150_), .A3(new_n1151_), .ZN(new_n1762_));
  NAND4_X1   g1471(.A1(new_n1762_), .A2(new_n1143_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1763_));
  OAI21_X1   g1472(.A1(new_n1761_), .A2(new_n1763_), .B(new_n264_), .ZN(new_n1764_));
  AOI21_X1   g1473(.A1(new_n1424_), .A2(new_n1422_), .B(new_n315_), .ZN(new_n1765_));
  NAND2_X1   g1474(.A1(new_n1309_), .A2(new_n277_), .ZN(new_n1766_));
  NAND4_X1   g1475(.A1(new_n1765_), .A2(new_n1766_), .A3(new_n854_), .A4(new_n1160_), .ZN(new_n1767_));
  OAI21_X1   g1476(.A1(\shift[4] ), .A2(new_n1767_), .B(new_n1553_), .ZN(new_n1768_));
  NOR3_X1    g1477(.A1(new_n1162_), .A2(new_n1553_), .A3(\shift[4] ), .ZN(new_n1769_));
  NOR2_X1    g1478(.A1(new_n1769_), .A2(\shift[5] ), .ZN(new_n1770_));
  NAND4_X1   g1479(.A1(new_n1559_), .A2(new_n270_), .A3(new_n1558_), .A4(new_n1560_), .ZN(new_n1771_));
  NAND4_X1   g1480(.A1(new_n1171_), .A2(\shift[4] ), .A3(new_n1174_), .A4(new_n1170_), .ZN(new_n1772_));
  NAND3_X1   g1481(.A1(new_n1771_), .A2(new_n1772_), .A3(new_n265_), .ZN(new_n1773_));
  AOI21_X1   g1482(.A1(new_n1770_), .A2(new_n1768_), .B(new_n1773_), .ZN(new_n1774_));
  OAI21_X1   g1483(.A1(new_n1774_), .A2(new_n264_), .B(new_n1764_), .ZN(\result[39] ));
  NOR4_X1    g1484(.A1(new_n287_), .A2(new_n270_), .A3(\shift[5] ), .A4(new_n267_), .ZN(new_n1776_));
  OAI21_X1   g1485(.A1(new_n1776_), .A2(\shift[6] ), .B(new_n1755_), .ZN(\result[40] ));
  NOR4_X1    g1486(.A1(new_n1272_), .A2(new_n1274_), .A3(new_n270_), .A4(new_n1270_), .ZN(new_n1778_));
  OAI21_X1   g1487(.A1(new_n1269_), .A2(new_n270_), .B(new_n265_), .ZN(new_n1779_));
  NOR2_X1    g1488(.A1(new_n1779_), .A2(new_n1778_), .ZN(new_n1780_));
  NAND2_X1   g1489(.A1(new_n587_), .A2(new_n590_), .ZN(new_n1781_));
  NAND3_X1   g1490(.A1(new_n1055_), .A2(new_n1781_), .A3(new_n278_), .ZN(new_n1782_));
  NAND2_X1   g1491(.A1(new_n1224_), .A2(new_n1225_), .ZN(new_n1783_));
  NOR2_X1    g1492(.A1(new_n1783_), .A2(new_n1782_), .ZN(new_n1784_));
  NAND4_X1   g1493(.A1(new_n1784_), .A2(\shift[4] ), .A3(new_n1216_), .A4(new_n265_), .ZN(new_n1785_));
  OAI21_X1   g1494(.A1(new_n1780_), .A2(new_n1785_), .B(new_n264_), .ZN(new_n1786_));
  NAND3_X1   g1495(.A1(new_n1639_), .A2(new_n1640_), .A3(new_n278_), .ZN(new_n1787_));
  AOI21_X1   g1496(.A1(new_n1049_), .A2(new_n1050_), .B(new_n315_), .ZN(new_n1788_));
  OAI21_X1   g1497(.A1(new_n1068_), .A2(new_n1070_), .B(new_n277_), .ZN(new_n1789_));
  NAND4_X1   g1498(.A1(new_n1788_), .A2(new_n1787_), .A3(new_n1789_), .A4(new_n1373_), .ZN(new_n1790_));
  OAI21_X1   g1499(.A1(\shift[4] ), .A2(new_n1790_), .B(new_n1580_), .ZN(new_n1791_));
  NOR3_X1    g1500(.A1(new_n1232_), .A2(new_n1580_), .A3(\shift[4] ), .ZN(new_n1792_));
  NOR2_X1    g1501(.A1(new_n1792_), .A2(\shift[5] ), .ZN(new_n1793_));
  NAND2_X1   g1502(.A1(new_n1256_), .A2(new_n270_), .ZN(new_n1794_));
  AOI21_X1   g1503(.A1(new_n1248_), .A2(\shift[4] ), .B(\shift[5] ), .ZN(new_n1795_));
  NAND2_X1   g1504(.A1(new_n1794_), .A2(new_n1795_), .ZN(new_n1796_));
  AOI21_X1   g1505(.A1(new_n1793_), .A2(new_n1791_), .B(new_n1796_), .ZN(new_n1797_));
  OAI21_X1   g1506(.A1(new_n1797_), .A2(new_n264_), .B(new_n1786_), .ZN(\result[41] ));
  NOR4_X1    g1507(.A1(new_n270_), .A2(\shift[2] ), .A3(\shift[3] ), .A4(\shift[5] ), .ZN(new_n1799_));
  OAI21_X1   g1508(.A1(\shift[6] ), .A2(new_n1799_), .B(new_n1755_), .ZN(\result[42] ));
  NOR2_X1    g1509(.A1(new_n1598_), .A2(new_n270_), .ZN(new_n1801_));
  NOR3_X1    g1510(.A1(new_n1344_), .A2(new_n1204_), .A3(new_n1341_), .ZN(new_n1802_));
  NOR3_X1    g1511(.A1(new_n1801_), .A2(new_n1802_), .A3(\shift[5] ), .ZN(new_n1803_));
  AND4_X2    g1512(.A1(new_n1291_), .A2(new_n1295_), .A3(new_n1297_), .A4(new_n1298_), .Z(new_n1804_));
  NAND4_X1   g1513(.A1(new_n1804_), .A2(new_n1289_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1805_));
  OAI21_X1   g1514(.A1(new_n1805_), .A2(new_n1803_), .B(new_n264_), .ZN(new_n1806_));
  AOI21_X1   g1515(.A1(new_n1140_), .A2(new_n1139_), .B(new_n315_), .ZN(new_n1807_));
  NAND2_X1   g1516(.A1(new_n1430_), .A2(new_n277_), .ZN(new_n1808_));
  NAND4_X1   g1517(.A1(new_n1807_), .A2(new_n1425_), .A3(new_n1808_), .A4(new_n1160_), .ZN(new_n1809_));
  AOI21_X1   g1518(.A1(new_n1157_), .A2(new_n846_), .B(new_n315_), .ZN(new_n1810_));
  NAND4_X1   g1519(.A1(new_n1810_), .A2(new_n1608_), .A3(new_n1166_), .A4(new_n1607_), .ZN(new_n1811_));
  OAI21_X1   g1520(.A1(new_n1809_), .A2(\shift[4] ), .B(new_n1811_), .ZN(new_n1812_));
  NOR3_X1    g1521(.A1(new_n1811_), .A2(new_n1306_), .A3(\shift[4] ), .ZN(new_n1813_));
  NOR2_X1    g1522(.A1(new_n1813_), .A2(\shift[5] ), .ZN(new_n1814_));
  NOR2_X1    g1523(.A1(new_n1184_), .A2(new_n1320_), .ZN(new_n1815_));
  NOR2_X1    g1524(.A1(new_n1322_), .A2(new_n1323_), .ZN(new_n1816_));
  NAND3_X1   g1525(.A1(new_n1816_), .A2(new_n270_), .A3(new_n1815_), .ZN(new_n1817_));
  NAND4_X1   g1526(.A1(new_n1318_), .A2(\shift[4] ), .A3(new_n1317_), .A4(new_n1170_), .ZN(new_n1818_));
  NAND3_X1   g1527(.A1(new_n1817_), .A2(new_n265_), .A3(new_n1818_), .ZN(new_n1819_));
  AOI21_X1   g1528(.A1(new_n1814_), .A2(new_n1812_), .B(new_n1819_), .ZN(new_n1820_));
  OAI21_X1   g1529(.A1(new_n1820_), .A2(new_n264_), .B(new_n1806_), .ZN(\result[43] ));
  NOR4_X1    g1530(.A1(new_n1350_), .A2(new_n270_), .A3(\shift[5] ), .A4(new_n267_), .ZN(new_n1822_));
  OAI21_X1   g1531(.A1(new_n1822_), .A2(\shift[6] ), .B(new_n1755_), .ZN(\result[44] ));
  NOR2_X1    g1532(.A1(new_n1399_), .A2(new_n270_), .ZN(new_n1824_));
  NAND3_X1   g1533(.A1(new_n1400_), .A2(new_n1273_), .A3(new_n440_), .ZN(new_n1825_));
  NAND2_X1   g1534(.A1(new_n1825_), .A2(new_n265_), .ZN(new_n1826_));
  NOR2_X1    g1535(.A1(new_n1824_), .A2(new_n1826_), .ZN(new_n1827_));
  INV_X1     g1536(.I(new_n1370_), .ZN(new_n1828_));
  NAND4_X1   g1537(.A1(new_n1828_), .A2(\shift[4] ), .A3(new_n1362_), .A4(new_n265_), .ZN(new_n1829_));
  OAI21_X1   g1538(.A1(new_n1827_), .A2(new_n1829_), .B(new_n264_), .ZN(new_n1830_));
  NAND3_X1   g1539(.A1(new_n1049_), .A2(new_n1050_), .A3(new_n278_), .ZN(new_n1831_));
  AOI21_X1   g1540(.A1(new_n1212_), .A2(new_n1213_), .B(new_n315_), .ZN(new_n1832_));
  NAND4_X1   g1541(.A1(new_n1832_), .A2(new_n1831_), .A3(new_n1373_), .A4(new_n1376_), .ZN(new_n1833_));
  NAND4_X1   g1542(.A1(new_n416_), .A2(new_n1646_), .A3(new_n1381_), .A4(new_n1242_), .ZN(new_n1834_));
  OAI21_X1   g1543(.A1(new_n1833_), .A2(\shift[4] ), .B(new_n1834_), .ZN(new_n1835_));
  NOR3_X1    g1544(.A1(new_n1642_), .A2(new_n1834_), .A3(\shift[4] ), .ZN(new_n1836_));
  NOR2_X1    g1545(.A1(new_n1836_), .A2(\shift[5] ), .ZN(new_n1837_));
  NAND2_X1   g1546(.A1(new_n1392_), .A2(new_n270_), .ZN(new_n1838_));
  NAND3_X1   g1547(.A1(new_n1664_), .A2(\shift[4] ), .A3(new_n1663_), .ZN(new_n1839_));
  NAND3_X1   g1548(.A1(new_n1838_), .A2(new_n1839_), .A3(new_n265_), .ZN(new_n1840_));
  AOI21_X1   g1549(.A1(new_n1837_), .A2(new_n1835_), .B(new_n1840_), .ZN(new_n1841_));
  OAI21_X1   g1550(.A1(new_n1841_), .A2(new_n264_), .B(new_n1830_), .ZN(\result[45] ));
  NOR2_X1    g1551(.A1(new_n1673_), .A2(new_n270_), .ZN(new_n1843_));
  NOR3_X1    g1552(.A1(new_n1453_), .A2(new_n441_), .A3(new_n908_), .ZN(new_n1844_));
  NOR3_X1    g1553(.A1(new_n1843_), .A2(new_n1844_), .A3(\shift[5] ), .ZN(new_n1845_));
  NOR3_X1    g1554(.A1(new_n1418_), .A2(new_n1415_), .A3(new_n1419_), .ZN(new_n1846_));
  NAND4_X1   g1555(.A1(new_n1846_), .A2(\shift[4] ), .A3(new_n1410_), .A4(new_n265_), .ZN(new_n1847_));
  OAI21_X1   g1556(.A1(new_n1845_), .A2(new_n1847_), .B(new_n264_), .ZN(new_n1848_));
  NAND3_X1   g1557(.A1(new_n1140_), .A2(new_n278_), .A3(new_n1139_), .ZN(new_n1849_));
  AOI21_X1   g1558(.A1(new_n1286_), .A2(new_n1284_), .B(new_n315_), .ZN(new_n1850_));
  NAND4_X1   g1559(.A1(new_n1849_), .A2(new_n1425_), .A3(new_n1850_), .A4(new_n1428_), .ZN(new_n1851_));
  AOI21_X1   g1560(.A1(new_n1303_), .A2(new_n852_), .B(new_n315_), .ZN(new_n1852_));
  NAND4_X1   g1561(.A1(new_n1852_), .A2(new_n1608_), .A3(new_n1684_), .A4(new_n848_), .ZN(new_n1853_));
  OAI21_X1   g1562(.A1(new_n1851_), .A2(\shift[4] ), .B(new_n1853_), .ZN(new_n1854_));
  NOR3_X1    g1563(.A1(new_n1680_), .A2(\shift[4] ), .A3(new_n1853_), .ZN(new_n1855_));
  NOR2_X1    g1564(.A1(new_n1855_), .A2(\shift[5] ), .ZN(new_n1856_));
  NAND2_X1   g1565(.A1(new_n1443_), .A2(new_n270_), .ZN(new_n1857_));
  NAND4_X1   g1566(.A1(new_n1693_), .A2(\shift[4] ), .A3(new_n1317_), .A4(new_n1438_), .ZN(new_n1858_));
  NAND3_X1   g1567(.A1(new_n1857_), .A2(new_n1858_), .A3(new_n265_), .ZN(new_n1859_));
  AOI21_X1   g1568(.A1(new_n1856_), .A2(new_n1854_), .B(new_n1859_), .ZN(new_n1860_));
  OAI21_X1   g1569(.A1(new_n1860_), .A2(new_n264_), .B(new_n1848_), .ZN(\result[47] ));
  NOR2_X1    g1570(.A1(\shift[2] ), .A2(\shift[3] ), .ZN(new_n1862_));
  NOR3_X1    g1571(.A1(new_n1699_), .A2(\shift[4] ), .A3(new_n267_), .ZN(new_n1863_));
  NOR2_X1    g1572(.A1(new_n1863_), .A2(\shift[5] ), .ZN(new_n1864_));
  AOI21_X1   g1573(.A1(new_n1864_), .A2(new_n1862_), .B(new_n274_), .ZN(new_n1865_));
  OAI21_X1   g1574(.A1(new_n1865_), .A2(\shift[6] ), .B(new_n1593_), .ZN(\result[48] ));
  OAI21_X1   g1575(.A1(new_n692_), .A2(new_n702_), .B(new_n265_), .ZN(new_n1867_));
  AOI21_X1   g1576(.A1(new_n676_), .A2(\shift[4] ), .B(new_n1867_), .ZN(new_n1868_));
  NOR3_X1    g1577(.A1(new_n1222_), .A2(new_n315_), .A3(new_n1223_), .ZN(new_n1869_));
  NOR2_X1    g1578(.A1(new_n1353_), .A2(new_n1869_), .ZN(new_n1870_));
  NAND4_X1   g1579(.A1(new_n1870_), .A2(\shift[4] ), .A3(new_n347_), .A4(new_n358_), .ZN(new_n1871_));
  NAND2_X1   g1580(.A1(new_n630_), .A2(new_n270_), .ZN(new_n1872_));
  NAND3_X1   g1581(.A1(new_n1872_), .A2(new_n1871_), .A3(new_n265_), .ZN(new_n1873_));
  OAI21_X1   g1582(.A1(new_n1873_), .A2(new_n1868_), .B(new_n264_), .ZN(new_n1874_));
  INV_X1     g1583(.I(new_n336_), .ZN(new_n1875_));
  OAI21_X1   g1584(.A1(new_n1875_), .A2(\shift[4] ), .B(new_n1711_), .ZN(new_n1876_));
  NOR3_X1    g1585(.A1(new_n336_), .A2(new_n1711_), .A3(\shift[4] ), .ZN(new_n1877_));
  NOR2_X1    g1586(.A1(new_n1877_), .A2(\shift[5] ), .ZN(new_n1878_));
  OAI21_X1   g1587(.A1(new_n535_), .A2(new_n552_), .B(\shift[4] ), .ZN(new_n1879_));
  NAND3_X1   g1588(.A1(new_n1879_), .A2(new_n1481_), .A3(new_n265_), .ZN(new_n1880_));
  AOI21_X1   g1589(.A1(new_n1878_), .A2(new_n1876_), .B(new_n1880_), .ZN(new_n1881_));
  OAI21_X1   g1590(.A1(new_n1881_), .A2(new_n264_), .B(new_n1874_), .ZN(\result[49] ));
  NOR2_X1    g1591(.A1(\shift[4] ), .A2(\shift[5] ), .ZN(new_n1883_));
  NOR2_X1    g1592(.A1(new_n274_), .A2(new_n1883_), .ZN(new_n1884_));
  NAND4_X1   g1593(.A1(new_n709_), .A2(new_n270_), .A3(new_n265_), .A4(new_n267_), .ZN(new_n1885_));
  NAND2_X1   g1594(.A1(new_n1885_), .A2(\shift[6] ), .ZN(new_n1886_));
  OAI21_X1   g1595(.A1(new_n1884_), .A2(\shift[6] ), .B(new_n1886_), .ZN(\result[50] ));
  NOR4_X1    g1596(.A1(new_n908_), .A2(new_n270_), .A3(new_n915_), .A4(new_n925_), .ZN(new_n1888_));
  OAI21_X1   g1597(.A1(new_n1000_), .A2(new_n270_), .B(new_n265_), .ZN(new_n1889_));
  NOR2_X1    g1598(.A1(new_n1889_), .A2(new_n1888_), .ZN(new_n1890_));
  NAND2_X1   g1599(.A1(new_n1039_), .A2(new_n270_), .ZN(new_n1891_));
  INV_X1     g1600(.I(new_n753_), .ZN(new_n1892_));
  NOR2_X1    g1601(.A1(new_n1892_), .A2(new_n1406_), .ZN(new_n1893_));
  NAND4_X1   g1602(.A1(new_n1893_), .A2(\shift[4] ), .A3(new_n758_), .A4(new_n764_), .ZN(new_n1894_));
  NAND3_X1   g1603(.A1(new_n1891_), .A2(new_n1894_), .A3(new_n265_), .ZN(new_n1895_));
  OAI21_X1   g1604(.A1(new_n1890_), .A2(new_n1895_), .B(new_n264_), .ZN(new_n1896_));
  AOI21_X1   g1605(.A1(new_n1504_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n1897_));
  NAND3_X1   g1606(.A1(new_n866_), .A2(new_n278_), .A3(new_n875_), .ZN(new_n1898_));
  OR2_X2     g1607(.A1(new_n886_), .A2(new_n896_), .Z(new_n1899_));
  NOR4_X1    g1608(.A1(new_n1899_), .A2(new_n1898_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1900_));
  NOR2_X1    g1609(.A1(new_n1897_), .A2(new_n1900_), .ZN(new_n1901_));
  NOR4_X1    g1610(.A1(new_n944_), .A2(new_n270_), .A3(new_n961_), .A4(\shift[5] ), .ZN(new_n1902_));
  AOI21_X1   g1611(.A1(new_n1511_), .A2(\shift[4] ), .B(new_n265_), .ZN(new_n1903_));
  NOR2_X1    g1612(.A1(new_n1903_), .A2(new_n1902_), .ZN(new_n1904_));
  NAND2_X1   g1613(.A1(new_n822_), .A2(new_n270_), .ZN(new_n1905_));
  AOI21_X1   g1614(.A1(new_n856_), .A2(\shift[4] ), .B(new_n680_), .ZN(new_n1906_));
  NAND2_X1   g1615(.A1(new_n1906_), .A2(new_n1905_), .ZN(new_n1907_));
  AOI21_X1   g1616(.A1(new_n1901_), .A2(new_n1904_), .B(new_n1907_), .ZN(new_n1908_));
  OAI21_X1   g1617(.A1(new_n1908_), .A2(new_n264_), .B(new_n1896_), .ZN(\result[51] ));
  NOR2_X1    g1618(.A1(new_n1566_), .A2(new_n1736_), .ZN(new_n1910_));
  OAI21_X1   g1619(.A1(new_n716_), .A2(new_n1572_), .B(\shift[6] ), .ZN(new_n1911_));
  OAI21_X1   g1620(.A1(new_n1910_), .A2(\shift[6] ), .B(new_n1911_), .ZN(\result[52] ));
  NOR2_X1    g1621(.A1(new_n1519_), .A2(\shift[4] ), .ZN(new_n1913_));
  NOR2_X1    g1622(.A1(new_n670_), .A2(new_n674_), .ZN(new_n1914_));
  NOR2_X1    g1623(.A1(new_n1487_), .A2(new_n1489_), .ZN(new_n1915_));
  NOR3_X1    g1624(.A1(new_n1914_), .A2(new_n1915_), .A3(new_n315_), .ZN(new_n1916_));
  NOR2_X1    g1625(.A1(new_n1118_), .A2(new_n1119_), .ZN(new_n1917_));
  NAND3_X1   g1626(.A1(new_n1917_), .A2(\shift[4] ), .A3(new_n1916_), .ZN(new_n1918_));
  NAND4_X1   g1627(.A1(new_n1918_), .A2(new_n1743_), .A3(new_n1101_), .A4(new_n1543_), .ZN(new_n1919_));
  OAI21_X1   g1628(.A1(new_n1919_), .A2(new_n1913_), .B(new_n264_), .ZN(new_n1920_));
  AOI21_X1   g1629(.A1(new_n1053_), .A2(new_n270_), .B(\shift[5] ), .ZN(new_n1921_));
  NAND2_X1   g1630(.A1(new_n1212_), .A2(new_n1213_), .ZN(new_n1922_));
  INV_X1     g1631(.I(new_n339_), .ZN(new_n1923_));
  NOR2_X1    g1632(.A1(new_n338_), .A2(\shift[0] ), .ZN(new_n1924_));
  NAND3_X1   g1633(.A1(new_n873_), .A2(new_n284_), .A3(\shift[0] ), .ZN(new_n1925_));
  NAND2_X1   g1634(.A1(new_n1924_), .A2(new_n1925_), .ZN(new_n1926_));
  NAND2_X1   g1635(.A1(new_n1926_), .A2(new_n1923_), .ZN(new_n1927_));
  NAND3_X1   g1636(.A1(new_n1927_), .A2(new_n309_), .A3(new_n345_), .ZN(new_n1928_));
  NAND3_X1   g1637(.A1(new_n1922_), .A2(new_n1928_), .A3(new_n278_), .ZN(new_n1929_));
  NAND2_X1   g1638(.A1(new_n1360_), .A2(new_n1359_), .ZN(new_n1930_));
  NOR2_X1    g1639(.A1(new_n320_), .A2(new_n324_), .ZN(new_n1931_));
  OAI22_X1   g1640(.A1(new_n1930_), .A2(new_n315_), .B1(new_n1931_), .B2(new_n291_), .ZN(new_n1932_));
  NOR4_X1    g1641(.A1(new_n1932_), .A2(new_n1929_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1933_));
  NOR2_X1    g1642(.A1(new_n1933_), .A2(new_n1921_), .ZN(new_n1934_));
  NOR3_X1    g1643(.A1(new_n283_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n1935_));
  OAI21_X1   g1644(.A1(new_n431_), .A2(new_n433_), .B(new_n1935_), .ZN(new_n1936_));
  NAND3_X1   g1645(.A1(new_n1936_), .A2(new_n551_), .A3(new_n278_), .ZN(new_n1937_));
  OAI22_X1   g1646(.A1(new_n534_), .A2(new_n315_), .B1(new_n1246_), .B2(new_n291_), .ZN(new_n1938_));
  NOR4_X1    g1647(.A1(new_n1938_), .A2(new_n270_), .A3(new_n1937_), .A4(\shift[5] ), .ZN(new_n1939_));
  AOI21_X1   g1648(.A1(new_n1105_), .A2(\shift[4] ), .B(new_n265_), .ZN(new_n1940_));
  NOR2_X1    g1649(.A1(new_n1940_), .A2(new_n1939_), .ZN(new_n1941_));
  NAND3_X1   g1650(.A1(new_n1095_), .A2(\shift[5] ), .A3(new_n1093_), .ZN(new_n1942_));
  NAND3_X1   g1651(.A1(new_n1525_), .A2(new_n1524_), .A3(new_n265_), .ZN(new_n1943_));
  NAND3_X1   g1652(.A1(new_n1942_), .A2(new_n1943_), .A3(new_n679_), .ZN(new_n1944_));
  AOI21_X1   g1653(.A1(new_n1934_), .A2(new_n1941_), .B(new_n1944_), .ZN(new_n1945_));
  OAI21_X1   g1654(.A1(new_n1945_), .A2(new_n264_), .B(new_n1920_), .ZN(\result[53] ));
  NAND2_X1   g1655(.A1(new_n1567_), .A2(new_n1911_), .ZN(\result[54] ));
  AOI21_X1   g1656(.A1(new_n1758_), .A2(new_n1757_), .B(new_n265_), .ZN(new_n1948_));
  NAND2_X1   g1657(.A1(new_n1562_), .A2(new_n270_), .ZN(new_n1949_));
  NOR2_X1    g1658(.A1(new_n1949_), .A2(new_n1948_), .ZN(new_n1950_));
  NOR3_X1    g1659(.A1(new_n999_), .A2(new_n315_), .A3(new_n914_), .ZN(new_n1951_));
  AOI21_X1   g1660(.A1(new_n1329_), .A2(new_n277_), .B(new_n1204_), .ZN(new_n1952_));
  NAND3_X1   g1661(.A1(new_n1952_), .A2(new_n265_), .A3(new_n1951_), .ZN(new_n1953_));
  NAND4_X1   g1662(.A1(new_n1548_), .A2(\shift[5] ), .A3(new_n1149_), .A4(new_n1291_), .ZN(new_n1954_));
  NAND3_X1   g1663(.A1(new_n1953_), .A2(new_n1954_), .A3(new_n270_), .ZN(new_n1955_));
  OAI21_X1   g1664(.A1(new_n1950_), .A2(new_n1955_), .B(new_n264_), .ZN(new_n1956_));
  OAI21_X1   g1665(.A1(new_n1545_), .A2(\shift[4] ), .B(new_n1767_), .ZN(new_n1957_));
  NOR3_X1    g1666(.A1(new_n1143_), .A2(new_n1767_), .A3(\shift[4] ), .ZN(new_n1958_));
  NOR2_X1    g1667(.A1(new_n1958_), .A2(\shift[5] ), .ZN(new_n1959_));
  INV_X1     g1668(.I(new_n1553_), .ZN(new_n1960_));
  NAND4_X1   g1669(.A1(new_n1960_), .A2(new_n1185_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n1961_));
  AOI21_X1   g1670(.A1(new_n1959_), .A2(new_n1957_), .B(new_n1961_), .ZN(new_n1962_));
  OAI21_X1   g1671(.A1(new_n1962_), .A2(new_n264_), .B(new_n1956_), .ZN(\result[55] ));
  NAND4_X1   g1672(.A1(new_n267_), .A2(new_n270_), .A3(\shift[5] ), .A4(new_n264_), .ZN(\result[56] ));
  NOR2_X1    g1673(.A1(new_n1269_), .A2(new_n265_), .ZN(new_n1965_));
  OAI21_X1   g1674(.A1(new_n1263_), .A2(new_n265_), .B(new_n270_), .ZN(new_n1966_));
  NOR2_X1    g1675(.A1(new_n1966_), .A2(new_n1965_), .ZN(new_n1967_));
  NAND4_X1   g1676(.A1(new_n1582_), .A2(new_n265_), .A3(new_n1271_), .A4(new_n1273_), .ZN(new_n1968_));
  NAND4_X1   g1677(.A1(new_n1219_), .A2(\shift[5] ), .A3(new_n1224_), .A4(new_n1225_), .ZN(new_n1969_));
  NAND3_X1   g1678(.A1(new_n1968_), .A2(new_n1969_), .A3(new_n270_), .ZN(new_n1970_));
  OAI21_X1   g1679(.A1(new_n1967_), .A2(new_n1970_), .B(new_n264_), .ZN(new_n1971_));
  OAI21_X1   g1680(.A1(new_n1576_), .A2(\shift[4] ), .B(new_n1790_), .ZN(new_n1972_));
  NOR3_X1    g1681(.A1(new_n1216_), .A2(new_n1790_), .A3(\shift[4] ), .ZN(new_n1973_));
  NOR2_X1    g1682(.A1(new_n1973_), .A2(\shift[5] ), .ZN(new_n1974_));
  INV_X1     g1683(.I(new_n1580_), .ZN(new_n1975_));
  NAND4_X1   g1684(.A1(new_n1975_), .A2(\shift[4] ), .A3(new_n265_), .A4(new_n1256_), .ZN(new_n1976_));
  AOI21_X1   g1685(.A1(new_n1974_), .A2(new_n1972_), .B(new_n1976_), .ZN(new_n1977_));
  OAI21_X1   g1686(.A1(new_n1977_), .A2(new_n264_), .B(new_n1971_), .ZN(\result[57] ));
  NAND2_X1   g1687(.A1(new_n1543_), .A2(new_n266_), .ZN(new_n1979_));
  NOR3_X1    g1688(.A1(new_n1979_), .A2(new_n1735_), .A3(new_n709_), .ZN(new_n1980_));
  OAI21_X1   g1689(.A1(new_n1980_), .A2(\shift[6] ), .B(new_n1136_), .ZN(\result[58] ));
  NOR3_X1    g1690(.A1(new_n1339_), .A2(new_n1333_), .A3(\shift[4] ), .ZN(new_n1982_));
  NAND3_X1   g1691(.A1(new_n948_), .A2(new_n309_), .A3(new_n949_), .ZN(new_n1983_));
  AND4_X2    g1692(.A1(new_n266_), .A2(new_n1317_), .A3(new_n1983_), .A4(new_n1170_), .Z(new_n1984_));
  NAND2_X1   g1693(.A1(new_n1612_), .A2(new_n1613_), .ZN(new_n1985_));
  NAND4_X1   g1694(.A1(new_n1985_), .A2(new_n1804_), .A3(new_n1984_), .A4(new_n1543_), .ZN(new_n1986_));
  OAI21_X1   g1695(.A1(new_n1986_), .A2(new_n1982_), .B(new_n264_), .ZN(new_n1987_));
  OAI21_X1   g1696(.A1(new_n1602_), .A2(\shift[4] ), .B(new_n1809_), .ZN(new_n1988_));
  NOR3_X1    g1697(.A1(new_n1809_), .A2(new_n1289_), .A3(\shift[4] ), .ZN(new_n1989_));
  NOR2_X1    g1698(.A1(new_n1989_), .A2(\shift[5] ), .ZN(new_n1990_));
  NAND4_X1   g1699(.A1(new_n1324_), .A2(\shift[4] ), .A3(new_n1313_), .A4(new_n265_), .ZN(new_n1991_));
  AOI21_X1   g1700(.A1(new_n1990_), .A2(new_n1988_), .B(new_n1991_), .ZN(new_n1992_));
  OAI21_X1   g1701(.A1(new_n1992_), .A2(new_n264_), .B(new_n1987_), .ZN(\result[59] ));
  NOR3_X1    g1702(.A1(new_n1349_), .A2(new_n1735_), .A3(new_n1979_), .ZN(new_n1994_));
  OAI21_X1   g1703(.A1(new_n1994_), .A2(\shift[6] ), .B(new_n1136_), .ZN(\result[60] ));
  AND2_X2    g1704(.A1(new_n1399_), .A2(new_n270_), .Z(new_n1996_));
  INV_X1     g1705(.I(new_n1388_), .ZN(new_n1997_));
  NAND4_X1   g1706(.A1(new_n1997_), .A2(new_n1828_), .A3(new_n1825_), .A4(new_n1543_), .ZN(new_n1998_));
  OAI21_X1   g1707(.A1(new_n1998_), .A2(new_n1996_), .B(new_n264_), .ZN(new_n1999_));
  INV_X1     g1708(.I(new_n1362_), .ZN(new_n2000_));
  OAI21_X1   g1709(.A1(new_n2000_), .A2(\shift[4] ), .B(new_n1833_), .ZN(new_n2001_));
  NOR3_X1    g1710(.A1(new_n1833_), .A2(new_n1362_), .A3(\shift[4] ), .ZN(new_n2002_));
  NOR2_X1    g1711(.A1(new_n2002_), .A2(\shift[5] ), .ZN(new_n2003_));
  NAND4_X1   g1712(.A1(new_n1392_), .A2(new_n1652_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n2004_));
  AOI21_X1   g1713(.A1(new_n2003_), .A2(new_n2001_), .B(new_n2004_), .ZN(new_n2005_));
  OAI21_X1   g1714(.A1(new_n2005_), .A2(new_n264_), .B(new_n1999_), .ZN(\result[61] ));
  NOR3_X1    g1715(.A1(new_n1450_), .A2(new_n1448_), .A3(\shift[4] ), .ZN(new_n2007_));
  INV_X1     g1716(.I(new_n1439_), .ZN(new_n2008_));
  NAND2_X1   g1717(.A1(new_n1688_), .A2(new_n1689_), .ZN(new_n2009_));
  NAND4_X1   g1718(.A1(new_n2009_), .A2(new_n2008_), .A3(new_n1846_), .A4(new_n1543_), .ZN(new_n2010_));
  OAI21_X1   g1719(.A1(new_n2010_), .A2(new_n2007_), .B(new_n264_), .ZN(new_n2011_));
  INV_X1     g1720(.I(new_n1410_), .ZN(new_n2012_));
  OAI21_X1   g1721(.A1(new_n2012_), .A2(\shift[4] ), .B(new_n1851_), .ZN(new_n2013_));
  NOR3_X1    g1722(.A1(new_n1410_), .A2(new_n1851_), .A3(\shift[4] ), .ZN(new_n2014_));
  NOR2_X1    g1723(.A1(new_n2014_), .A2(\shift[5] ), .ZN(new_n2015_));
  NAND4_X1   g1724(.A1(new_n1443_), .A2(new_n1433_), .A3(\shift[4] ), .A4(new_n265_), .ZN(new_n2016_));
  AOI21_X1   g1725(.A1(new_n2015_), .A2(new_n2013_), .B(new_n2016_), .ZN(new_n2017_));
  OAI21_X1   g1726(.A1(new_n2017_), .A2(new_n264_), .B(new_n2011_), .ZN(\result[63] ));
  NAND2_X1   g1727(.A1(new_n268_), .A2(\shift[6] ), .ZN(new_n2019_));
  OAI21_X1   g1728(.A1(new_n289_), .A2(\shift[6] ), .B(new_n2019_), .ZN(\result[64] ));
  OAI21_X1   g1729(.A1(new_n381_), .A2(new_n475_), .B(\shift[6] ), .ZN(new_n2021_));
  OAI21_X1   g1730(.A1(new_n706_), .A2(\shift[6] ), .B(new_n2021_), .ZN(\result[65] ));
  NAND2_X1   g1731(.A1(new_n711_), .A2(\shift[6] ), .ZN(new_n2023_));
  OAI21_X1   g1732(.A1(new_n718_), .A2(\shift[6] ), .B(new_n2023_), .ZN(\result[66] ));
  OAI21_X1   g1733(.A1(new_n963_), .A2(new_n1041_), .B(new_n264_), .ZN(new_n2025_));
  OAI21_X1   g1734(.A1(new_n900_), .A2(new_n264_), .B(new_n2025_), .ZN(\result[67] ));
  OAI21_X1   g1735(.A1(\shift[6] ), .A2(new_n1045_), .B(new_n2019_), .ZN(\result[68] ));
  OAI21_X1   g1736(.A1(new_n1109_), .A2(new_n1129_), .B(new_n264_), .ZN(new_n2028_));
  OAI21_X1   g1737(.A1(new_n1065_), .A2(new_n1097_), .B(\shift[6] ), .ZN(new_n2029_));
  NAND2_X1   g1738(.A1(new_n2028_), .A2(new_n2029_), .ZN(\result[69] ));
  NAND2_X1   g1739(.A1(new_n1698_), .A2(new_n2019_), .ZN(\result[70] ));
  OAI21_X1   g1740(.A1(new_n1153_), .A2(new_n1168_), .B(\shift[6] ), .ZN(new_n2032_));
  OAI21_X1   g1741(.A1(new_n1207_), .A2(\shift[6] ), .B(new_n2032_), .ZN(\result[71] ));
  NAND4_X1   g1742(.A1(new_n267_), .A2(\shift[4] ), .A3(new_n265_), .A4(\shift[6] ), .ZN(\result[72] ));
  OAI21_X1   g1743(.A1(new_n1265_), .A2(new_n1276_), .B(new_n264_), .ZN(new_n2035_));
  OAI21_X1   g1744(.A1(new_n1228_), .A2(new_n1244_), .B(\shift[6] ), .ZN(new_n2036_));
  NAND2_X1   g1745(.A1(new_n2035_), .A2(new_n2036_), .ZN(\result[73] ));
  OAI21_X1   g1746(.A1(new_n1281_), .A2(\shift[6] ), .B(new_n2019_), .ZN(\result[74] ));
  OAI21_X1   g1747(.A1(new_n1301_), .A2(new_n1315_), .B(\shift[6] ), .ZN(new_n2039_));
  OAI21_X1   g1748(.A1(new_n1347_), .A2(\shift[6] ), .B(new_n2039_), .ZN(\result[75] ));
  OAI21_X1   g1749(.A1(new_n1351_), .A2(\shift[6] ), .B(new_n2019_), .ZN(\result[76] ));
  OAI21_X1   g1750(.A1(new_n1372_), .A2(new_n1383_), .B(\shift[6] ), .ZN(new_n2042_));
  OAI21_X1   g1751(.A1(new_n1404_), .A2(\shift[6] ), .B(new_n2042_), .ZN(\result[77] ));
  OAI21_X1   g1752(.A1(new_n1421_), .A2(new_n1435_), .B(\shift[6] ), .ZN(new_n2044_));
  OAI21_X1   g1753(.A1(new_n1456_), .A2(\shift[6] ), .B(new_n2044_), .ZN(\result[79] ));
  OAI21_X1   g1754(.A1(new_n1461_), .A2(\shift[6] ), .B(new_n1755_), .ZN(\result[80] ));
  OAI21_X1   g1755(.A1(new_n1483_), .A2(new_n1494_), .B(new_n264_), .ZN(new_n2047_));
  OAI21_X1   g1756(.A1(new_n1471_), .A2(new_n264_), .B(new_n2047_), .ZN(\result[81] ));
  OAI21_X1   g1757(.A1(\shift[6] ), .A2(new_n1497_), .B(new_n1755_), .ZN(\result[82] ));
  OAI21_X1   g1758(.A1(new_n1513_), .A2(new_n1514_), .B(new_n264_), .ZN(new_n2050_));
  OAI21_X1   g1759(.A1(new_n1506_), .A2(new_n264_), .B(new_n2050_), .ZN(\result[83] ));
  OAI21_X1   g1760(.A1(\shift[6] ), .A2(new_n1517_), .B(new_n1755_), .ZN(\result[84] ));
  OAI21_X1   g1761(.A1(new_n1535_), .A2(new_n1536_), .B(new_n264_), .ZN(new_n2053_));
  OAI21_X1   g1762(.A1(new_n1528_), .A2(new_n264_), .B(new_n2053_), .ZN(\result[85] ));
  OAI21_X1   g1763(.A1(\shift[6] ), .A2(new_n1539_), .B(new_n1755_), .ZN(\result[86] ));
  OAI21_X1   g1764(.A1(new_n1550_), .A2(new_n1544_), .B(\shift[6] ), .ZN(new_n2056_));
  OAI21_X1   g1765(.A1(new_n1564_), .A2(\shift[6] ), .B(new_n2056_), .ZN(\result[87] ));
  NAND2_X1   g1766(.A1(new_n1566_), .A2(\shift[6] ), .ZN(new_n2058_));
  OAI21_X1   g1767(.A1(new_n1573_), .A2(\shift[6] ), .B(new_n2058_), .ZN(\result[88] ));
  OAI21_X1   g1768(.A1(new_n1577_), .A2(new_n1575_), .B(\shift[6] ), .ZN(new_n2060_));
  OAI21_X1   g1769(.A1(new_n1589_), .A2(\shift[6] ), .B(new_n2060_), .ZN(\result[89] ));
  OAI21_X1   g1770(.A1(new_n1592_), .A2(new_n1572_), .B(new_n264_), .ZN(new_n2062_));
  NAND2_X1   g1771(.A1(new_n2062_), .A2(new_n1755_), .ZN(\result[90] ));
  OAI21_X1   g1772(.A1(new_n1615_), .A2(new_n1618_), .B(new_n264_), .ZN(new_n2064_));
  OAI21_X1   g1773(.A1(new_n1601_), .A2(new_n1604_), .B(\shift[6] ), .ZN(new_n2065_));
  NAND2_X1   g1774(.A1(new_n2065_), .A2(new_n2064_), .ZN(\result[91] ));
  OAI21_X1   g1775(.A1(new_n1623_), .A2(\shift[6] ), .B(new_n1755_), .ZN(\result[92] ));
  OAI21_X1   g1776(.A1(new_n1660_), .A2(new_n1666_), .B(new_n264_), .ZN(new_n2068_));
  OAI21_X1   g1777(.A1(new_n1632_), .A2(new_n1644_), .B(\shift[6] ), .ZN(new_n2069_));
  NAND2_X1   g1778(.A1(new_n2069_), .A2(new_n2068_), .ZN(\result[93] ));
  OAI21_X1   g1779(.A1(new_n1691_), .A2(new_n1695_), .B(new_n264_), .ZN(new_n2071_));
  OAI21_X1   g1780(.A1(new_n1677_), .A2(new_n1682_), .B(\shift[6] ), .ZN(new_n2072_));
  NAND2_X1   g1781(.A1(new_n2072_), .A2(new_n2071_), .ZN(\result[95] ));
  OAI21_X1   g1782(.A1(new_n1701_), .A2(\shift[6] ), .B(new_n1136_), .ZN(\result[96] ));
  OAI21_X1   g1783(.A1(new_n1716_), .A2(new_n1718_), .B(new_n264_), .ZN(new_n2075_));
  OAI21_X1   g1784(.A1(new_n1705_), .A2(new_n1707_), .B(\shift[6] ), .ZN(new_n2076_));
  NAND2_X1   g1785(.A1(new_n2076_), .A2(new_n2075_), .ZN(\result[97] ));
  OAI21_X1   g1786(.A1(new_n1721_), .A2(\shift[6] ), .B(new_n1136_), .ZN(\result[98] ));
  OAI21_X1   g1787(.A1(new_n1729_), .A2(new_n1730_), .B(new_n264_), .ZN(new_n2079_));
  OAI21_X1   g1788(.A1(new_n264_), .A2(new_n1726_), .B(new_n2079_), .ZN(\result[99] ));
  NAND2_X1   g1789(.A1(new_n1733_), .A2(\shift[6] ), .ZN(new_n2081_));
  OAI21_X1   g1790(.A1(new_n1738_), .A2(\shift[6] ), .B(new_n2081_), .ZN(\result[100] ));
  OAI21_X1   g1791(.A1(new_n1742_), .A2(new_n1744_), .B(\shift[6] ), .ZN(new_n2083_));
  OAI21_X1   g1792(.A1(new_n1753_), .A2(\shift[6] ), .B(new_n2083_), .ZN(\result[101] ));
  NAND2_X1   g1793(.A1(new_n1459_), .A2(new_n2081_), .ZN(\result[102] ));
  OAI21_X1   g1794(.A1(new_n1761_), .A2(new_n1763_), .B(\shift[6] ), .ZN(new_n2086_));
  OAI21_X1   g1795(.A1(new_n1774_), .A2(\shift[6] ), .B(new_n2086_), .ZN(\result[103] ));
  OAI21_X1   g1796(.A1(new_n1776_), .A2(new_n264_), .B(new_n1459_), .ZN(\result[104] ));
  OAI21_X1   g1797(.A1(new_n1780_), .A2(new_n1785_), .B(\shift[6] ), .ZN(new_n2089_));
  OAI21_X1   g1798(.A1(new_n1797_), .A2(\shift[6] ), .B(new_n2089_), .ZN(\result[105] ));
  OAI21_X1   g1799(.A1(new_n264_), .A2(new_n1799_), .B(new_n1459_), .ZN(\result[106] ));
  OAI21_X1   g1800(.A1(new_n1805_), .A2(new_n1803_), .B(\shift[6] ), .ZN(new_n2092_));
  OAI21_X1   g1801(.A1(new_n1820_), .A2(\shift[6] ), .B(new_n2092_), .ZN(\result[107] ));
  OAI21_X1   g1802(.A1(new_n1822_), .A2(new_n264_), .B(new_n1459_), .ZN(\result[108] ));
  OAI21_X1   g1803(.A1(new_n1827_), .A2(new_n1829_), .B(\shift[6] ), .ZN(new_n2095_));
  OAI21_X1   g1804(.A1(new_n1841_), .A2(\shift[6] ), .B(new_n2095_), .ZN(\result[109] ));
  OAI21_X1   g1805(.A1(new_n1845_), .A2(new_n1847_), .B(\shift[6] ), .ZN(new_n2097_));
  OAI21_X1   g1806(.A1(new_n1860_), .A2(\shift[6] ), .B(new_n2097_), .ZN(\result[111] ));
  OAI21_X1   g1807(.A1(new_n1865_), .A2(new_n264_), .B(new_n2062_), .ZN(\result[112] ));
  OAI21_X1   g1808(.A1(new_n1873_), .A2(new_n1868_), .B(\shift[6] ), .ZN(new_n2100_));
  OAI21_X1   g1809(.A1(new_n1881_), .A2(\shift[6] ), .B(new_n2100_), .ZN(\result[113] ));
  NAND2_X1   g1810(.A1(new_n1885_), .A2(new_n264_), .ZN(new_n2102_));
  OAI21_X1   g1811(.A1(new_n1884_), .A2(new_n264_), .B(new_n2102_), .ZN(\result[114] ));
  OAI21_X1   g1812(.A1(new_n1890_), .A2(new_n1895_), .B(\shift[6] ), .ZN(new_n2104_));
  OAI21_X1   g1813(.A1(new_n1908_), .A2(\shift[6] ), .B(new_n2104_), .ZN(\result[115] ));
  OAI21_X1   g1814(.A1(new_n716_), .A2(new_n1572_), .B(new_n264_), .ZN(new_n2106_));
  OAI21_X1   g1815(.A1(new_n1910_), .A2(new_n264_), .B(new_n2106_), .ZN(\result[116] ));
  OAI21_X1   g1816(.A1(new_n1919_), .A2(new_n1913_), .B(\shift[6] ), .ZN(new_n2108_));
  OAI21_X1   g1817(.A1(new_n1945_), .A2(\shift[6] ), .B(new_n2108_), .ZN(\result[117] ));
  NAND2_X1   g1818(.A1(new_n2058_), .A2(new_n2106_), .ZN(\result[118] ));
  OAI21_X1   g1819(.A1(new_n1950_), .A2(new_n1955_), .B(\shift[6] ), .ZN(new_n2111_));
  OAI21_X1   g1820(.A1(new_n1962_), .A2(\shift[6] ), .B(new_n2111_), .ZN(\result[119] ));
  NAND4_X1   g1821(.A1(new_n267_), .A2(new_n270_), .A3(\shift[5] ), .A4(\shift[6] ), .ZN(\result[120] ));
  OAI21_X1   g1822(.A1(new_n1967_), .A2(new_n1970_), .B(\shift[6] ), .ZN(new_n2114_));
  OAI21_X1   g1823(.A1(new_n1977_), .A2(\shift[6] ), .B(new_n2114_), .ZN(\result[121] ));
  OAI21_X1   g1824(.A1(new_n1980_), .A2(new_n264_), .B(new_n1698_), .ZN(\result[122] ));
  OAI21_X1   g1825(.A1(new_n1986_), .A2(new_n1982_), .B(\shift[6] ), .ZN(new_n2117_));
  OAI21_X1   g1826(.A1(new_n1992_), .A2(\shift[6] ), .B(new_n2117_), .ZN(\result[123] ));
  OAI21_X1   g1827(.A1(new_n1994_), .A2(new_n264_), .B(new_n1698_), .ZN(\result[124] ));
  OAI21_X1   g1828(.A1(new_n1998_), .A2(new_n1996_), .B(\shift[6] ), .ZN(new_n2120_));
  OAI21_X1   g1829(.A1(new_n2005_), .A2(\shift[6] ), .B(new_n2120_), .ZN(\result[125] ));
  OAI21_X1   g1830(.A1(new_n2010_), .A2(new_n2007_), .B(\shift[6] ), .ZN(new_n2122_));
  OAI21_X1   g1831(.A1(new_n2017_), .A2(\shift[6] ), .B(new_n2122_), .ZN(\result[127] ));
  OAI21_X1   g1832(.A1(new_n1281_), .A2(new_n264_), .B(new_n269_), .ZN(\result[14] ));
  NAND2_X1   g1833(.A1(new_n1593_), .A2(new_n1459_), .ZN(\result[30] ));
  OAI21_X1   g1834(.A1(\shift[6] ), .A2(new_n1799_), .B(new_n1755_), .ZN(\result[46] ));
  OAI21_X1   g1835(.A1(new_n1980_), .A2(\shift[6] ), .B(new_n1136_), .ZN(\result[62] ));
  OAI21_X1   g1836(.A1(new_n1281_), .A2(\shift[6] ), .B(new_n2019_), .ZN(\result[78] ));
  NAND2_X1   g1837(.A1(new_n2062_), .A2(new_n1755_), .ZN(\result[94] ));
  OAI21_X1   g1838(.A1(new_n264_), .A2(new_n1799_), .B(new_n1459_), .ZN(\result[110] ));
  OAI21_X1   g1839(.A1(new_n1980_), .A2(new_n264_), .B(new_n1698_), .ZN(\result[126] ));
endmodule


