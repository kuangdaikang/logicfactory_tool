// Benchmark "source.pla" written by ABC on Fri Feb 25 15:13:09 2022

module opa  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16,
    \v17.0 , \v17.1 , \v17.2 , \v17.3 , \v17.4 , \v17.5 , \v17.6 , \v17.7 ,
    \v17.8 , \v17.9 , \v17.10 , \v17.11 , \v17.12 , \v17.13 , \v17.14 ,
    \v17.15 , \v17.16 , \v17.17 , \v17.18 , \v17.19 , \v17.20 , \v17.21 ,
    \v17.22 , \v17.23 , \v17.24 , \v17.25 , \v17.26 , \v17.27 , \v17.28 ,
    \v17.29 , \v17.30 , \v17.31 , \v17.32 , \v17.33 , \v17.34 , \v17.35 ,
    \v17.36 , \v17.37 , \v17.38 , \v17.39 , \v17.40 , \v17.41 , \v17.42 ,
    \v17.43 , \v17.44 , \v17.45 , \v17.46 , \v17.47 , \v17.48 , \v17.49 ,
    \v17.50 , \v17.51 , \v17.52 , \v17.53 , \v17.54 , \v17.55 , \v17.56 ,
    \v17.57 , \v17.58 , \v17.59 , \v17.60 , \v17.61 , \v17.62 , \v17.63 ,
    \v17.64 , \v17.65 , \v17.66 , \v17.67 , \v17.68   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16;
  output \v17.0 , \v17.1 , \v17.2 , \v17.3 , \v17.4 , \v17.5 , \v17.6 ,
    \v17.7 , \v17.8 , \v17.9 , \v17.10 , \v17.11 , \v17.12 , \v17.13 ,
    \v17.14 , \v17.15 , \v17.16 , \v17.17 , \v17.18 , \v17.19 , \v17.20 ,
    \v17.21 , \v17.22 , \v17.23 , \v17.24 , \v17.25 , \v17.26 , \v17.27 ,
    \v17.28 , \v17.29 , \v17.30 , \v17.31 , \v17.32 , \v17.33 , \v17.34 ,
    \v17.35 , \v17.36 , \v17.37 , \v17.38 , \v17.39 , \v17.40 , \v17.41 ,
    \v17.42 , \v17.43 , \v17.44 , \v17.45 , \v17.46 , \v17.47 , \v17.48 ,
    \v17.49 , \v17.50 , \v17.51 , \v17.52 , \v17.53 , \v17.54 , \v17.55 ,
    \v17.56 , \v17.57 , \v17.58 , \v17.59 , \v17.60 , \v17.61 , \v17.62 ,
    \v17.63 , \v17.64 , \v17.65 , \v17.66 , \v17.67 , \v17.68 ;
  wire new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n198_, new_n199_,
    new_n201_, new_n202_, new_n203_, new_n205_, new_n206_, new_n207_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_;
  assign new_n88_ = v2 & ~v4;
  assign new_n89_ = v4 & v6;
  assign new_n90_ = ~v2 & new_n89_;
  assign new_n91_ = ~new_n88_ & ~new_n90_;
  assign new_n92_ = v5 & ~new_n91_;
  assign new_n93_ = ~v3 & new_n92_;
  assign new_n94_ = v5 & ~v6;
  assign new_n95_ = v2 & ~new_n94_;
  assign new_n96_ = ~v5 & v6;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = ~v4 & ~new_n97_;
  assign new_n99_ = v3 & new_n98_;
  assign new_n100_ = ~new_n93_ & ~new_n99_;
  assign new_n101_ = v1 & ~new_n100_;
  assign new_n102_ = v6 & ~v13;
  assign new_n103_ = v2 & new_n102_;
  assign new_n104_ = ~v4 & ~new_n103_;
  assign new_n105_ = ~v1 & ~new_n104_;
  assign new_n106_ = v4 & ~v6;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = v5 & ~new_n107_;
  assign new_n109_ = ~v1 & ~v4;
  assign new_n110_ = ~v5 & ~v6;
  assign new_n111_ = new_n109_ & new_n110_;
  assign new_n112_ = ~new_n108_ & ~new_n111_;
  assign new_n113_ = v3 & ~new_n112_;
  assign new_n114_ = ~new_n101_ & ~new_n113_;
  assign \v17.0  = ~v0 & ~new_n114_;
  assign new_n116_ = ~v1 & ~new_n110_;
  assign new_n117_ = ~v4 & ~v6;
  assign new_n118_ = ~v3 & ~new_n117_;
  assign new_n119_ = ~new_n116_ & ~new_n118_;
  assign new_n120_ = ~v2 & ~new_n119_;
  assign new_n121_ = ~v3 & ~v4;
  assign new_n122_ = ~v1 & ~new_n121_;
  assign new_n123_ = v1 & v2;
  assign new_n124_ = ~v3 & ~new_n123_;
  assign new_n125_ = ~new_n89_ & ~new_n124_;
  assign new_n126_ = ~v7 & ~v9;
  assign new_n127_ = ~v16 & ~new_n126_;
  assign new_n128_ = ~v15 & new_n127_;
  assign new_n129_ = ~v14 & new_n128_;
  assign new_n130_ = ~v12 & new_n129_;
  assign new_n131_ = ~v8 & new_n130_;
  assign new_n132_ = v3 & new_n131_;
  assign new_n133_ = v5 & ~new_n132_;
  assign new_n134_ = v2 & ~new_n133_;
  assign new_n135_ = v1 & ~v5;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = ~new_n125_ & new_n136_;
  assign new_n138_ = ~new_n122_ & new_n137_;
  assign new_n139_ = ~new_n120_ & new_n138_;
  assign \v17.1  = ~v0 & ~new_n139_;
  assign new_n141_ = v6 & new_n131_;
  assign new_n142_ = v4 & new_n141_;
  assign new_n143_ = v2 & new_n142_;
  assign new_n144_ = ~v2 & new_n117_;
  assign new_n145_ = ~new_n143_ & ~new_n144_;
  assign new_n146_ = v1 & ~new_n145_;
  assign new_n147_ = ~v1 & v13;
  assign new_n148_ = v6 & ~new_n147_;
  assign new_n149_ = v2 & new_n148_;
  assign new_n150_ = v5 & ~new_n149_;
  assign new_n151_ = ~v4 & new_n150_;
  assign new_n152_ = ~new_n146_ & ~new_n151_;
  assign new_n153_ = v3 & ~new_n152_;
  assign new_n154_ = ~v1 & v6;
  assign new_n155_ = v3 & ~new_n154_;
  assign new_n156_ = v2 & ~new_n155_;
  assign new_n157_ = v1 & ~v3;
  assign new_n158_ = ~v4 & ~new_n157_;
  assign new_n159_ = ~new_n156_ & new_n158_;
  assign new_n160_ = ~v5 & ~new_n159_;
  assign new_n161_ = v1 & v6;
  assign new_n162_ = v4 & ~new_n161_;
  assign new_n163_ = ~v4 & v6;
  assign new_n164_ = ~new_n116_ & ~new_n163_;
  assign new_n165_ = ~v2 & ~new_n164_;
  assign new_n166_ = ~new_n162_ & ~new_n165_;
  assign new_n167_ = ~v3 & ~new_n166_;
  assign new_n168_ = ~v4 & ~new_n110_;
  assign new_n169_ = ~v2 & new_n168_;
  assign new_n170_ = ~v1 & new_n169_;
  assign new_n171_ = ~new_n167_ & ~new_n170_;
  assign new_n172_ = ~new_n160_ & new_n171_;
  assign new_n173_ = ~new_n153_ & new_n172_;
  assign \v17.2  = ~v0 & ~new_n173_;
  assign new_n175_ = ~v0 & ~v1;
  assign new_n176_ = v2 & new_n175_;
  assign new_n177_ = v3 & new_n176_;
  assign new_n178_ = v4 & new_n177_;
  assign new_n179_ = v5 & new_n178_;
  assign \v17.3  = ~v6 & new_n179_;
  assign new_n181_ = ~v2 & new_n175_;
  assign new_n182_ = v3 & new_n181_;
  assign new_n183_ = v4 & new_n182_;
  assign new_n184_ = v5 & new_n183_;
  assign \v17.4  = ~v6 & new_n184_;
  assign new_n186_ = ~v0 & v1;
  assign new_n187_ = ~v2 & new_n186_;
  assign new_n188_ = v3 & new_n187_;
  assign new_n189_ = v4 & new_n188_;
  assign new_n190_ = ~v5 & new_n189_;
  assign \v17.5  = v6 & new_n190_;
  assign \v17.6  = ~v6 & new_n190_;
  assign new_n193_ = v2 & new_n186_;
  assign new_n194_ = v3 & new_n193_;
  assign new_n195_ = ~v4 & new_n194_;
  assign new_n196_ = v5 & new_n195_;
  assign \v17.7  = ~v6 & new_n196_;
  assign new_n198_ = ~v4 & new_n177_;
  assign new_n199_ = v5 & new_n198_;
  assign \v17.8  = v6 & new_n199_;
  assign new_n201_ = ~v3 & new_n187_;
  assign new_n202_ = ~v4 & new_n201_;
  assign new_n203_ = v5 & new_n202_;
  assign \v17.9  = v6 & new_n203_;
  assign new_n205_ = ~v3 & new_n193_;
  assign new_n206_ = ~v4 & new_n205_;
  assign new_n207_ = ~v5 & new_n206_;
  assign \v17.10  = ~v6 & new_n207_;
  assign new_n209_ = v4 & new_n194_;
  assign new_n210_ = v5 & new_n209_;
  assign new_n211_ = v6 & new_n210_;
  assign new_n212_ = v7 & new_n211_;
  assign new_n213_ = v8 & new_n212_;
  assign new_n214_ = ~v9 & new_n213_;
  assign new_n215_ = ~v12 & new_n214_;
  assign new_n216_ = ~v14 & new_n215_;
  assign new_n217_ = ~v15 & new_n216_;
  assign \v17.11  = ~v16 & new_n217_;
  assign new_n219_ = ~v7 & new_n211_;
  assign new_n220_ = v8 & new_n219_;
  assign new_n221_ = ~v9 & new_n220_;
  assign new_n222_ = ~v12 & new_n221_;
  assign new_n223_ = ~v14 & new_n222_;
  assign new_n224_ = ~v15 & new_n223_;
  assign \v17.12  = ~v16 & new_n224_;
  assign new_n226_ = ~v8 & new_n219_;
  assign new_n227_ = ~v9 & new_n226_;
  assign new_n228_ = ~v12 & new_n227_;
  assign new_n229_ = ~v14 & new_n228_;
  assign new_n230_ = ~v15 & new_n229_;
  assign \v17.13  = ~v16 & new_n230_;
  assign new_n232_ = ~v1 & ~v6;
  assign new_n233_ = v2 & ~new_n232_;
  assign new_n234_ = v5 & ~new_n233_;
  assign new_n235_ = v2 & v5;
  assign new_n236_ = v6 & ~new_n235_;
  assign new_n237_ = ~v1 & new_n236_;
  assign new_n238_ = ~v2 & ~v6;
  assign new_n239_ = v1 & new_n238_;
  assign new_n240_ = ~new_n237_ & ~new_n239_;
  assign new_n241_ = ~new_n234_ & new_n240_;
  assign new_n242_ = ~v4 & ~new_n241_;
  assign new_n243_ = v3 & new_n242_;
  assign \v17.14  = ~v0 & new_n243_;
  assign new_n245_ = ~v2 & ~new_n110_;
  assign new_n246_ = ~v1 & new_n245_;
  assign new_n247_ = v2 & ~new_n89_;
  assign new_n248_ = v5 & ~new_n163_;
  assign new_n249_ = ~new_n247_ & new_n248_;
  assign new_n250_ = v1 & ~new_n249_;
  assign new_n251_ = v2 & ~v5;
  assign new_n252_ = ~new_n106_ & ~new_n251_;
  assign new_n253_ = ~new_n250_ & new_n252_;
  assign new_n254_ = ~new_n246_ & new_n253_;
  assign new_n255_ = ~v3 & ~new_n254_;
  assign new_n256_ = v4 & new_n131_;
  assign new_n257_ = v3 & new_n256_;
  assign new_n258_ = ~new_n135_ & ~new_n257_;
  assign new_n259_ = v2 & ~new_n258_;
  assign new_n260_ = ~v1 & v4;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = ~new_n255_ & new_n261_;
  assign new_n263_ = ~v10 & ~new_n262_;
  assign new_n264_ = v3 & ~v6;
  assign new_n265_ = ~new_n121_ & ~new_n264_;
  assign new_n266_ = v5 & ~new_n265_;
  assign new_n267_ = v1 & new_n266_;
  assign new_n268_ = ~v8 & v9;
  assign new_n269_ = v7 & new_n268_;
  assign new_n270_ = ~v12 & ~v14;
  assign new_n271_ = ~v15 & ~v16;
  assign new_n272_ = new_n270_ & new_n271_;
  assign new_n273_ = new_n269_ & new_n272_;
  assign new_n274_ = v6 & ~new_n273_;
  assign new_n275_ = v5 & new_n274_;
  assign new_n276_ = v4 & ~new_n275_;
  assign new_n277_ = v3 & new_n276_;
  assign new_n278_ = ~new_n267_ & ~new_n277_;
  assign new_n279_ = v2 & ~new_n278_;
  assign new_n280_ = ~new_n94_ & ~new_n96_;
  assign new_n281_ = v1 & new_n280_;
  assign new_n282_ = v4 & ~new_n281_;
  assign new_n283_ = v3 & new_n282_;
  assign new_n284_ = ~new_n279_ & ~new_n283_;
  assign new_n285_ = ~new_n263_ & new_n284_;
  assign \v17.15  = ~v0 & ~new_n285_;
  assign new_n287_ = ~v7 & v9;
  assign new_n288_ = v7 & ~v9;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign new_n290_ = ~v16 & ~new_n289_;
  assign new_n291_ = ~v15 & new_n290_;
  assign new_n292_ = ~v14 & new_n291_;
  assign new_n293_ = ~v12 & new_n292_;
  assign new_n294_ = ~v8 & new_n293_;
  assign new_n295_ = v6 & new_n294_;
  assign new_n296_ = v5 & new_n295_;
  assign new_n297_ = v4 & new_n296_;
  assign new_n298_ = v3 & new_n297_;
  assign new_n299_ = ~v4 & ~v5;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = v2 & ~new_n300_;
  assign new_n302_ = ~v3 & ~v5;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = v1 & ~new_n303_;
  assign new_n305_ = ~new_n165_ & ~new_n251_;
  assign new_n306_ = ~new_n162_ & new_n305_;
  assign new_n307_ = ~v3 & ~new_n306_;
  assign new_n308_ = ~new_n304_ & ~new_n307_;
  assign new_n309_ = v10 & ~new_n308_;
  assign \v17.16  = ~v0 & new_n309_;
  assign new_n311_ = ~v2 & v6;
  assign new_n312_ = ~v4 & ~new_n311_;
  assign new_n313_ = ~v1 & ~new_n312_;
  assign new_n314_ = v1 & new_n251_;
  assign new_n315_ = ~v4 & ~new_n314_;
  assign new_n316_ = ~v6 & ~new_n315_;
  assign new_n317_ = ~v2 & new_n163_;
  assign new_n318_ = ~new_n316_ & ~new_n317_;
  assign new_n319_ = ~new_n313_ & new_n318_;
  assign new_n320_ = ~v3 & ~new_n319_;
  assign new_n321_ = v4 & ~v5;
  assign new_n322_ = ~v2 & v3;
  assign new_n323_ = new_n117_ & new_n322_;
  assign new_n324_ = ~new_n321_ & ~new_n323_;
  assign new_n325_ = v1 & ~new_n324_;
  assign new_n326_ = ~v4 & v5;
  assign new_n327_ = v3 & new_n326_;
  assign new_n328_ = ~new_n321_ & ~new_n327_;
  assign new_n329_ = ~v6 & ~new_n328_;
  assign new_n330_ = v5 & ~new_n123_;
  assign new_n331_ = ~v4 & new_n330_;
  assign new_n332_ = v3 & new_n331_;
  assign new_n333_ = ~new_n329_ & ~new_n332_;
  assign new_n334_ = ~new_n325_ & new_n333_;
  assign new_n335_ = ~new_n320_ & new_n334_;
  assign \v17.17  = ~v0 & ~new_n335_;
  assign new_n337_ = ~v3 & v4;
  assign new_n338_ = ~v2 & new_n337_;
  assign new_n339_ = v3 & ~v4;
  assign new_n340_ = v2 & new_n339_;
  assign new_n341_ = ~new_n338_ & ~new_n340_;
  assign new_n342_ = v5 & ~new_n341_;
  assign new_n343_ = v1 & new_n342_;
  assign new_n344_ = new_n299_ & new_n322_;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = v6 & ~new_n345_;
  assign new_n347_ = ~v1 & v3;
  assign new_n348_ = new_n299_ & new_n347_;
  assign new_n349_ = ~new_n346_ & ~new_n348_;
  assign \v17.18  = ~v0 & ~new_n349_;
  assign new_n351_ = v2 & new_n299_;
  assign new_n352_ = ~v2 & v4;
  assign new_n353_ = new_n94_ & new_n352_;
  assign new_n354_ = ~new_n351_ & ~new_n353_;
  assign new_n355_ = v1 & ~new_n354_;
  assign new_n356_ = ~v1 & ~v2;
  assign new_n357_ = v5 & v6;
  assign new_n358_ = v4 & new_n357_;
  assign new_n359_ = new_n356_ & new_n358_;
  assign new_n360_ = ~new_n355_ & ~new_n359_;
  assign new_n361_ = v3 & ~new_n360_;
  assign \v17.19  = ~v0 & new_n361_;
  assign new_n363_ = v2 & v3;
  assign new_n364_ = v4 & v5;
  assign new_n365_ = new_n363_ & new_n364_;
  assign new_n366_ = ~v2 & ~v3;
  assign new_n367_ = new_n299_ & new_n366_;
  assign new_n368_ = ~new_n365_ & ~new_n367_;
  assign new_n369_ = ~v6 & ~new_n368_;
  assign new_n370_ = v1 & new_n369_;
  assign new_n371_ = ~v2 & v5;
  assign new_n372_ = v6 & ~new_n371_;
  assign new_n373_ = v4 & new_n372_;
  assign new_n374_ = v3 & new_n373_;
  assign new_n375_ = ~v1 & new_n374_;
  assign new_n376_ = ~new_n370_ & ~new_n375_;
  assign \v17.20  = ~v0 & ~new_n376_;
  assign new_n378_ = v5 & new_n131_;
  assign new_n379_ = v4 & new_n378_;
  assign new_n380_ = v3 & new_n379_;
  assign new_n381_ = v1 & new_n380_;
  assign new_n382_ = ~v3 & new_n299_;
  assign new_n383_ = ~new_n381_ & ~new_n382_;
  assign new_n384_ = v6 & ~new_n383_;
  assign new_n385_ = ~v1 & ~v3;
  assign new_n386_ = new_n299_ & new_n385_;
  assign new_n387_ = ~new_n384_ & ~new_n386_;
  assign new_n388_ = v2 & ~new_n387_;
  assign new_n389_ = ~v1 & new_n366_;
  assign new_n390_ = ~v4 & new_n94_;
  assign new_n391_ = new_n389_ & new_n390_;
  assign new_n392_ = ~new_n388_ & ~new_n391_;
  assign \v17.21  = ~v0 & ~new_n392_;
  assign new_n394_ = ~v1 & new_n321_;
  assign new_n395_ = v1 & ~v4;
  assign new_n396_ = new_n94_ & new_n395_;
  assign new_n397_ = ~new_n394_ & ~new_n396_;
  assign new_n398_ = v2 & ~new_n397_;
  assign new_n399_ = ~v6 & ~v11;
  assign new_n400_ = ~v5 & ~new_n399_;
  assign new_n401_ = v4 & new_n400_;
  assign new_n402_ = v1 & new_n401_;
  assign new_n403_ = ~new_n398_ & ~new_n402_;
  assign new_n404_ = v3 & ~new_n403_;
  assign \v17.22  = ~v0 & new_n404_;
  assign new_n406_ = v2 & ~new_n161_;
  assign new_n407_ = v1 & new_n311_;
  assign new_n408_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = ~v5 & ~new_n408_;
  assign new_n410_ = v4 & new_n409_;
  assign new_n411_ = v3 & new_n410_;
  assign \v17.23  = ~v0 & new_n411_;
  assign new_n413_ = v4 & new_n96_;
  assign new_n414_ = ~new_n390_ & ~new_n413_;
  assign new_n415_ = v3 & ~new_n414_;
  assign new_n416_ = v2 & new_n415_;
  assign new_n417_ = v1 & new_n416_;
  assign \v17.24  = ~v0 & new_n417_;
  assign new_n419_ = v1 & new_n143_;
  assign new_n420_ = ~v1 & ~new_n102_;
  assign new_n421_ = v2 & ~new_n420_;
  assign new_n422_ = ~v4 & ~new_n421_;
  assign new_n423_ = ~new_n419_ & ~new_n422_;
  assign new_n424_ = v3 & ~new_n423_;
  assign new_n425_ = v3 & v4;
  assign new_n426_ = ~v2 & ~new_n425_;
  assign new_n427_ = ~v1 & new_n426_;
  assign new_n428_ = ~new_n424_ & ~new_n427_;
  assign new_n429_ = v5 & ~new_n428_;
  assign new_n430_ = v5 & ~new_n339_;
  assign new_n431_ = ~v6 & ~new_n430_;
  assign new_n432_ = v1 & new_n431_;
  assign new_n433_ = ~v1 & ~new_n425_;
  assign new_n434_ = ~new_n121_ & ~new_n433_;
  assign new_n435_ = v6 & ~new_n434_;
  assign new_n436_ = ~new_n394_ & ~new_n435_;
  assign new_n437_ = ~new_n432_ & new_n436_;
  assign new_n438_ = ~v2 & ~new_n437_;
  assign new_n439_ = ~v4 & new_n96_;
  assign new_n440_ = ~new_n337_ & ~new_n439_;
  assign new_n441_ = ~v1 & ~new_n440_;
  assign new_n442_ = ~v5 & ~new_n356_;
  assign new_n443_ = ~new_n106_ & ~new_n442_;
  assign new_n444_ = ~v3 & ~new_n443_;
  assign new_n445_ = ~new_n441_ & ~new_n444_;
  assign new_n446_ = ~new_n438_ & new_n445_;
  assign new_n447_ = ~new_n429_ & new_n446_;
  assign \v17.25  = ~v0 & ~new_n447_;
  assign new_n449_ = v5 & new_n102_;
  assign new_n450_ = ~v4 & ~new_n449_;
  assign new_n451_ = v2 & ~new_n450_;
  assign new_n452_ = ~v4 & new_n110_;
  assign new_n453_ = ~new_n364_ & ~new_n452_;
  assign new_n454_ = ~new_n451_ & new_n453_;
  assign new_n455_ = ~v1 & ~new_n454_;
  assign new_n456_ = v2 & ~new_n364_;
  assign new_n457_ = ~new_n96_ & ~new_n456_;
  assign new_n458_ = v1 & ~new_n457_;
  assign new_n459_ = v2 & new_n110_;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~new_n455_ & new_n460_;
  assign new_n462_ = v3 & ~new_n461_;
  assign new_n463_ = new_n89_ & new_n366_;
  assign new_n464_ = ~new_n88_ & ~new_n463_;
  assign new_n465_ = v5 & ~new_n464_;
  assign new_n466_ = v1 & new_n465_;
  assign new_n467_ = ~new_n462_ & ~new_n466_;
  assign \v17.26  = ~v0 & ~new_n467_;
  assign new_n469_ = ~v2 & ~new_n121_;
  assign new_n470_ = v2 & ~v3;
  assign new_n471_ = ~new_n364_ & ~new_n470_;
  assign new_n472_ = ~new_n469_ & new_n471_;
  assign new_n473_ = ~v6 & ~new_n472_;
  assign new_n474_ = v3 & ~new_n96_;
  assign new_n475_ = ~v4 & ~new_n474_;
  assign new_n476_ = ~new_n380_ & ~new_n475_;
  assign new_n477_ = v2 & ~new_n476_;
  assign new_n478_ = ~v3 & ~new_n248_;
  assign new_n479_ = ~new_n477_ & ~new_n478_;
  assign new_n480_ = ~new_n473_ & new_n479_;
  assign new_n481_ = v1 & ~new_n480_;
  assign new_n482_ = ~v4 & ~new_n371_;
  assign new_n483_ = ~v3 & ~new_n482_;
  assign new_n484_ = ~v6 & ~new_n321_;
  assign new_n485_ = ~new_n326_ & new_n484_;
  assign new_n486_ = ~v2 & ~new_n485_;
  assign new_n487_ = ~new_n168_ & ~new_n357_;
  assign new_n488_ = v3 & ~new_n487_;
  assign new_n489_ = ~new_n486_ & ~new_n488_;
  assign new_n490_ = ~new_n483_ & new_n489_;
  assign new_n491_ = ~v1 & ~new_n490_;
  assign new_n492_ = v2 & new_n302_;
  assign new_n493_ = new_n322_ & new_n326_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = ~new_n491_ & new_n494_;
  assign new_n496_ = ~new_n481_ & new_n495_;
  assign \v17.27  = ~v0 & ~new_n496_;
  assign new_n498_ = v2 & new_n379_;
  assign new_n499_ = ~new_n163_ & ~new_n238_;
  assign new_n500_ = ~new_n498_ & new_n499_;
  assign new_n501_ = v1 & ~new_n500_;
  assign new_n502_ = ~v1 & ~v5;
  assign new_n503_ = v4 & ~new_n502_;
  assign new_n504_ = ~v2 & ~new_n503_;
  assign new_n505_ = ~v4 & ~new_n102_;
  assign new_n506_ = ~v1 & new_n505_;
  assign new_n507_ = ~new_n504_ & ~new_n506_;
  assign new_n508_ = ~new_n501_ & new_n507_;
  assign new_n509_ = v3 & ~new_n508_;
  assign new_n510_ = v2 & v4;
  assign new_n511_ = new_n94_ & new_n510_;
  assign new_n512_ = ~new_n302_ & ~new_n511_;
  assign new_n513_ = v1 & ~new_n512_;
  assign new_n514_ = v3 & ~new_n109_;
  assign new_n515_ = ~v5 & ~new_n514_;
  assign new_n516_ = v2 & new_n515_;
  assign new_n517_ = ~v3 & v5;
  assign new_n518_ = ~v6 & ~new_n517_;
  assign new_n519_ = ~v2 & ~new_n518_;
  assign new_n520_ = v3 & ~new_n357_;
  assign new_n521_ = v4 & ~new_n520_;
  assign new_n522_ = ~new_n519_ & ~new_n521_;
  assign new_n523_ = ~v1 & ~new_n522_;
  assign new_n524_ = ~v2 & ~new_n117_;
  assign new_n525_ = ~new_n106_ & ~new_n524_;
  assign new_n526_ = ~v3 & ~new_n525_;
  assign new_n527_ = ~new_n523_ & ~new_n526_;
  assign new_n528_ = ~new_n516_ & new_n527_;
  assign new_n529_ = ~new_n513_ & new_n528_;
  assign new_n530_ = ~new_n509_ & new_n529_;
  assign \v17.28  = ~v0 & ~new_n530_;
  assign new_n532_ = new_n88_ & new_n94_;
  assign new_n533_ = ~new_n413_ & ~new_n532_;
  assign new_n534_ = v1 & ~new_n533_;
  assign new_n535_ = v2 & new_n321_;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = v3 & ~new_n536_;
  assign \v17.29  = ~v0 & new_n537_;
  assign new_n539_ = v1 & new_n88_;
  assign new_n540_ = ~new_n389_ & ~new_n539_;
  assign new_n541_ = v6 & ~new_n540_;
  assign new_n542_ = v3 & ~v5;
  assign new_n543_ = ~new_n517_ & ~new_n542_;
  assign new_n544_ = ~v4 & ~new_n543_;
  assign new_n545_ = v1 & new_n544_;
  assign new_n546_ = v3 & v5;
  assign new_n547_ = ~new_n302_ & ~new_n546_;
  assign new_n548_ = ~v1 & ~new_n547_;
  assign new_n549_ = v5 & ~v8;
  assign new_n550_ = new_n425_ & new_n549_;
  assign new_n551_ = v9 & ~v12;
  assign new_n552_ = ~v14 & new_n271_;
  assign new_n553_ = new_n551_ & new_n552_;
  assign new_n554_ = new_n550_ & new_n553_;
  assign new_n555_ = ~new_n548_ & ~new_n554_;
  assign new_n556_ = ~new_n545_ & new_n555_;
  assign new_n557_ = v2 & ~new_n556_;
  assign new_n558_ = ~v2 & new_n517_;
  assign new_n559_ = ~v4 & ~new_n558_;
  assign new_n560_ = ~v1 & ~new_n559_;
  assign new_n561_ = ~v4 & ~new_n135_;
  assign new_n562_ = ~v3 & ~new_n561_;
  assign new_n563_ = ~new_n321_ & ~new_n562_;
  assign new_n564_ = ~v2 & ~new_n563_;
  assign new_n565_ = v6 & ~new_n302_;
  assign new_n566_ = v4 & ~new_n565_;
  assign new_n567_ = ~new_n564_ & ~new_n566_;
  assign new_n568_ = ~new_n560_ & new_n567_;
  assign new_n569_ = ~new_n557_ & new_n568_;
  assign new_n570_ = ~new_n541_ & new_n569_;
  assign \v17.30  = ~v0 & ~new_n570_;
  assign new_n572_ = ~v5 & ~new_n161_;
  assign new_n573_ = ~v4 & new_n572_;
  assign new_n574_ = ~v2 & new_n573_;
  assign new_n575_ = v1 & new_n510_;
  assign new_n576_ = v6 & v7;
  assign new_n577_ = v5 & new_n576_;
  assign new_n578_ = new_n575_ & new_n577_;
  assign new_n579_ = ~v9 & ~v12;
  assign new_n580_ = ~v8 & new_n579_;
  assign new_n581_ = new_n552_ & new_n580_;
  assign new_n582_ = new_n578_ & new_n581_;
  assign new_n583_ = ~new_n574_ & ~new_n582_;
  assign new_n584_ = v3 & ~new_n583_;
  assign \v17.31  = ~v0 & new_n584_;
  assign new_n586_ = ~v3 & ~new_n235_;
  assign new_n587_ = v8 & v9;
  assign new_n588_ = v7 & ~new_n587_;
  assign new_n589_ = ~new_n268_ & ~new_n588_;
  assign new_n590_ = ~v16 & ~new_n589_;
  assign new_n591_ = ~v15 & new_n590_;
  assign new_n592_ = ~v14 & new_n591_;
  assign new_n593_ = ~v12 & new_n592_;
  assign new_n594_ = v5 & new_n593_;
  assign new_n595_ = v3 & new_n594_;
  assign new_n596_ = v2 & new_n595_;
  assign new_n597_ = new_n161_ & ~new_n596_;
  assign new_n598_ = ~new_n586_ & new_n597_;
  assign new_n599_ = v4 & ~new_n598_;
  assign new_n600_ = ~v1 & v2;
  assign new_n601_ = new_n546_ & new_n600_;
  assign new_n602_ = ~v2 & ~v5;
  assign new_n603_ = v1 & new_n602_;
  assign new_n604_ = ~new_n601_ & ~new_n603_;
  assign new_n605_ = ~v6 & ~new_n604_;
  assign new_n606_ = ~v1 & new_n302_;
  assign new_n607_ = v1 & v3;
  assign new_n608_ = ~v4 & new_n357_;
  assign new_n609_ = new_n607_ & new_n608_;
  assign new_n610_ = ~new_n606_ & ~new_n609_;
  assign new_n611_ = v2 & ~new_n610_;
  assign new_n612_ = v2 & ~v6;
  assign new_n613_ = ~v5 & ~new_n612_;
  assign new_n614_ = v1 & new_n613_;
  assign new_n615_ = ~v1 & v5;
  assign new_n616_ = ~v6 & ~new_n615_;
  assign new_n617_ = ~v2 & ~new_n616_;
  assign new_n618_ = ~new_n614_ & ~new_n617_;
  assign new_n619_ = ~v3 & ~new_n618_;
  assign new_n620_ = new_n356_ & new_n542_;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = ~new_n611_ & new_n621_;
  assign new_n623_ = ~new_n605_ & new_n622_;
  assign new_n624_ = ~new_n599_ & new_n623_;
  assign \v17.32  = ~v0 & ~new_n624_;
  assign new_n626_ = v6 & ~v7;
  assign new_n627_ = v4 & new_n626_;
  assign new_n628_ = new_n607_ & new_n627_;
  assign new_n629_ = new_n552_ & new_n579_;
  assign new_n630_ = new_n628_ & new_n629_;
  assign new_n631_ = ~new_n121_ & ~new_n630_;
  assign new_n632_ = v5 & ~new_n631_;
  assign new_n633_ = v2 & new_n632_;
  assign \v17.33  = ~v0 & new_n633_;
  assign new_n635_ = v4 & v12;
  assign new_n636_ = v1 & new_n635_;
  assign new_n637_ = ~new_n502_ & ~new_n636_;
  assign new_n638_ = ~v2 & ~new_n637_;
  assign new_n639_ = ~v5 & v12;
  assign new_n640_ = v2 & new_n639_;
  assign new_n641_ = ~new_n638_ & ~new_n640_;
  assign new_n642_ = ~v3 & ~new_n641_;
  assign new_n643_ = ~v4 & v12;
  assign new_n644_ = v4 & ~v7;
  assign new_n645_ = new_n268_ & new_n644_;
  assign new_n646_ = new_n272_ & new_n645_;
  assign new_n647_ = ~new_n643_ & ~new_n646_;
  assign new_n648_ = v5 & ~new_n647_;
  assign new_n649_ = v3 & new_n648_;
  assign new_n650_ = v2 & new_n649_;
  assign new_n651_ = v1 & new_n650_;
  assign new_n652_ = ~new_n642_ & ~new_n651_;
  assign new_n653_ = v6 & ~new_n652_;
  assign new_n654_ = ~v2 & ~v4;
  assign new_n655_ = new_n94_ & new_n654_;
  assign new_n656_ = ~new_n251_ & ~new_n655_;
  assign new_n657_ = v12 & ~new_n656_;
  assign new_n658_ = ~v1 & new_n657_;
  assign new_n659_ = ~new_n321_ & ~new_n658_;
  assign new_n660_ = ~v3 & ~new_n659_;
  assign new_n661_ = ~new_n653_ & ~new_n660_;
  assign \v17.34  = ~v0 & ~new_n661_;
  assign new_n663_ = ~v7 & new_n268_;
  assign new_n664_ = new_n272_ & new_n663_;
  assign new_n665_ = v4 & ~new_n664_;
  assign new_n666_ = v5 & ~new_n665_;
  assign new_n667_ = v3 & new_n666_;
  assign new_n668_ = v1 & new_n667_;
  assign new_n669_ = ~new_n302_ & ~new_n668_;
  assign new_n670_ = v6 & ~new_n669_;
  assign new_n671_ = ~new_n606_ & ~new_n670_;
  assign new_n672_ = v2 & ~new_n671_;
  assign new_n673_ = ~v2 & new_n94_;
  assign new_n674_ = ~v4 & ~new_n673_;
  assign new_n675_ = ~v1 & ~new_n674_;
  assign new_n676_ = v2 & new_n357_;
  assign new_n677_ = v4 & ~new_n676_;
  assign new_n678_ = ~new_n675_ & ~new_n677_;
  assign new_n679_ = ~v3 & ~new_n678_;
  assign new_n680_ = ~new_n672_ & ~new_n679_;
  assign \v17.35  = ~v0 & ~new_n680_;
  assign new_n682_ = v4 & ~new_n357_;
  assign new_n683_ = ~v3 & new_n682_;
  assign new_n684_ = v1 & new_n683_;
  assign \v17.36  = ~v0 & new_n684_;
  assign new_n686_ = ~v7 & ~v8;
  assign new_n687_ = v5 & new_n686_;
  assign new_n688_ = new_n363_ & new_n687_;
  assign new_n689_ = new_n553_ & new_n688_;
  assign new_n690_ = ~new_n302_ & ~new_n689_;
  assign new_n691_ = v6 & ~new_n690_;
  assign new_n692_ = v1 & new_n691_;
  assign new_n693_ = ~v3 & ~v6;
  assign new_n694_ = ~v1 & new_n693_;
  assign new_n695_ = ~new_n692_ & ~new_n694_;
  assign new_n696_ = v4 & ~new_n695_;
  assign \v17.37  = ~v0 & new_n696_;
  assign new_n698_ = ~v4 & ~new_n245_;
  assign new_n699_ = ~v1 & ~new_n698_;
  assign new_n700_ = ~new_n677_ & ~new_n699_;
  assign new_n701_ = ~v3 & ~new_n700_;
  assign new_n702_ = ~new_n672_ & ~new_n701_;
  assign \v17.38  = ~v0 & ~new_n702_;
  assign new_n704_ = ~new_n313_ & ~new_n682_;
  assign new_n705_ = ~v3 & ~new_n704_;
  assign new_n706_ = v1 & new_n363_;
  assign new_n707_ = new_n358_ & new_n706_;
  assign new_n708_ = new_n664_ & new_n707_;
  assign new_n709_ = ~new_n705_ & ~new_n708_;
  assign \v17.39  = ~v0 & ~new_n709_;
  assign new_n711_ = ~v3 & new_n117_;
  assign new_n712_ = v8 & new_n579_;
  assign new_n713_ = new_n552_ & new_n712_;
  assign new_n714_ = new_n628_ & new_n713_;
  assign new_n715_ = ~new_n711_ & ~new_n714_;
  assign new_n716_ = v5 & ~new_n715_;
  assign new_n717_ = v2 & new_n716_;
  assign \v17.40  = ~v0 & new_n717_;
  assign new_n719_ = ~new_n121_ & ~new_n714_;
  assign new_n720_ = v5 & ~new_n719_;
  assign new_n721_ = v2 & new_n720_;
  assign \v17.41  = ~v0 & new_n721_;
  assign new_n723_ = v1 & ~v6;
  assign new_n724_ = ~v5 & ~new_n723_;
  assign new_n725_ = ~v4 & new_n724_;
  assign new_n726_ = v2 & new_n725_;
  assign new_n727_ = ~v1 & ~new_n88_;
  assign new_n728_ = v2 & v6;
  assign new_n729_ = v4 & ~new_n728_;
  assign new_n730_ = ~new_n727_ & ~new_n729_;
  assign new_n731_ = v5 & ~new_n730_;
  assign new_n732_ = ~new_n726_ & ~new_n731_;
  assign new_n733_ = ~v3 & ~new_n732_;
  assign new_n734_ = new_n608_ & new_n706_;
  assign new_n735_ = ~new_n733_ & ~new_n734_;
  assign \v17.42  = ~v0 & ~new_n735_;
  assign new_n737_ = ~v0 & v2;
  assign new_n738_ = ~v3 & new_n737_;
  assign new_n739_ = ~v4 & new_n738_;
  assign \v17.43  = v5 & new_n739_;
  assign new_n741_ = ~v5 & ~new_n88_;
  assign new_n742_ = ~v1 & ~new_n741_;
  assign new_n743_ = ~new_n94_ & ~new_n168_;
  assign new_n744_ = v2 & ~new_n743_;
  assign new_n745_ = ~v2 & new_n364_;
  assign new_n746_ = ~new_n744_ & ~new_n745_;
  assign new_n747_ = ~new_n742_ & new_n746_;
  assign new_n748_ = ~v3 & ~new_n747_;
  assign new_n749_ = new_n123_ & new_n608_;
  assign new_n750_ = ~new_n748_ & ~new_n749_;
  assign \v17.44  = ~v0 & ~new_n750_;
  assign \v17.45  = v5 & new_n206_;
  assign new_n753_ = ~v3 & ~new_n89_;
  assign new_n754_ = ~v1 & new_n753_;
  assign new_n755_ = ~new_n714_ & ~new_n754_;
  assign new_n756_ = v2 & ~new_n755_;
  assign new_n757_ = ~v3 & new_n106_;
  assign new_n758_ = ~new_n756_ & ~new_n757_;
  assign new_n759_ = v5 & ~new_n758_;
  assign \v17.46  = ~v0 & new_n759_;
  assign new_n761_ = ~v7 & v8;
  assign new_n762_ = v5 & new_n761_;
  assign new_n763_ = new_n425_ & new_n762_;
  assign new_n764_ = new_n629_ & new_n763_;
  assign new_n765_ = ~new_n121_ & ~new_n764_;
  assign new_n766_ = v6 & ~new_n765_;
  assign new_n767_ = v1 & new_n766_;
  assign new_n768_ = v1 & v4;
  assign new_n769_ = v5 & ~new_n768_;
  assign new_n770_ = ~v1 & ~new_n163_;
  assign new_n771_ = ~new_n682_ & ~new_n770_;
  assign new_n772_ = ~new_n769_ & new_n771_;
  assign new_n773_ = ~v3 & ~new_n772_;
  assign new_n774_ = ~new_n767_ & ~new_n773_;
  assign new_n775_ = v2 & ~new_n774_;
  assign \v17.47  = ~v0 & new_n775_;
  assign new_n777_ = v2 & new_n94_;
  assign new_n778_ = ~v4 & ~new_n777_;
  assign new_n779_ = ~v1 & ~new_n778_;
  assign new_n780_ = ~v4 & ~new_n723_;
  assign new_n781_ = ~v5 & ~new_n780_;
  assign new_n782_ = ~v2 & new_n781_;
  assign new_n783_ = ~v8 & ~v9;
  assign new_n784_ = ~new_n588_ & ~new_n783_;
  assign new_n785_ = ~v16 & ~new_n784_;
  assign new_n786_ = ~v15 & new_n785_;
  assign new_n787_ = ~v14 & new_n786_;
  assign new_n788_ = ~v12 & new_n787_;
  assign new_n789_ = v5 & new_n788_;
  assign new_n790_ = v2 & new_n789_;
  assign new_n791_ = v6 & ~new_n790_;
  assign new_n792_ = v4 & ~new_n791_;
  assign new_n793_ = ~new_n782_ & ~new_n792_;
  assign new_n794_ = ~new_n779_ & new_n793_;
  assign new_n795_ = v3 & ~new_n794_;
  assign new_n796_ = ~v4 & ~new_n94_;
  assign new_n797_ = ~v3 & new_n796_;
  assign new_n798_ = ~v2 & new_n797_;
  assign new_n799_ = v1 & new_n798_;
  assign new_n800_ = ~new_n795_ & ~new_n799_;
  assign \v17.48  = ~v0 & ~new_n800_;
  assign new_n802_ = v7 & ~v8;
  assign new_n803_ = new_n235_ & new_n802_;
  assign new_n804_ = new_n553_ & new_n803_;
  assign new_n805_ = v6 & ~new_n804_;
  assign new_n806_ = v1 & new_n805_;
  assign new_n807_ = v4 & ~new_n806_;
  assign new_n808_ = v3 & new_n807_;
  assign \v17.49  = ~v0 & new_n808_;
  assign new_n810_ = new_n123_ & new_n577_;
  assign new_n811_ = ~v8 & new_n551_;
  assign new_n812_ = new_n552_ & new_n811_;
  assign new_n813_ = new_n810_ & new_n812_;
  assign new_n814_ = ~new_n572_ & ~new_n813_;
  assign new_n815_ = v4 & ~new_n814_;
  assign new_n816_ = v3 & new_n815_;
  assign \v17.50  = ~v0 & new_n816_;
  assign new_n818_ = v6 & ~new_n356_;
  assign new_n819_ = ~v5 & ~new_n818_;
  assign new_n820_ = ~new_n813_ & ~new_n819_;
  assign new_n821_ = v4 & ~new_n820_;
  assign new_n822_ = v3 & new_n821_;
  assign \v17.51  = ~v0 & new_n822_;
  assign new_n824_ = v5 & ~new_n273_;
  assign new_n825_ = v2 & ~new_n824_;
  assign new_n826_ = new_n161_ & ~new_n825_;
  assign new_n827_ = v4 & ~new_n826_;
  assign new_n828_ = v3 & new_n827_;
  assign \v17.52  = ~v0 & new_n828_;
  assign new_n830_ = ~v4 & new_n182_;
  assign \v17.53  = ~v5 & new_n830_;
  assign new_n832_ = v1 & v5;
  assign new_n833_ = ~v2 & ~new_n832_;
  assign new_n834_ = ~v1 & ~new_n94_;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = ~v4 & ~new_n835_;
  assign new_n837_ = ~new_n582_ & ~new_n836_;
  assign new_n838_ = v3 & ~new_n837_;
  assign \v17.54  = ~v0 & new_n838_;
  assign new_n840_ = new_n510_ & new_n577_;
  assign new_n841_ = new_n581_ & new_n840_;
  assign new_n842_ = ~new_n654_ & ~new_n841_;
  assign new_n843_ = v1 & ~new_n842_;
  assign new_n844_ = v5 & ~new_n728_;
  assign new_n845_ = ~v4 & ~new_n844_;
  assign new_n846_ = ~v1 & new_n845_;
  assign new_n847_ = ~new_n843_ & ~new_n846_;
  assign new_n848_ = v3 & ~new_n847_;
  assign \v17.55  = ~v0 & new_n848_;
  assign new_n850_ = v5 & ~new_n311_;
  assign new_n851_ = ~v1 & ~new_n850_;
  assign new_n852_ = ~new_n110_ & ~new_n357_;
  assign new_n853_ = ~v2 & ~new_n852_;
  assign new_n854_ = ~new_n851_ & ~new_n853_;
  assign new_n855_ = ~v4 & ~new_n854_;
  assign new_n856_ = ~new_n582_ & ~new_n855_;
  assign new_n857_ = v3 & ~new_n856_;
  assign \v17.56  = ~v0 & new_n857_;
  assign new_n859_ = v2 & ~new_n502_;
  assign new_n860_ = v12 & ~new_n859_;
  assign new_n861_ = ~v4 & new_n860_;
  assign new_n862_ = v3 & new_n861_;
  assign \v17.57  = ~v0 & new_n862_;
  assign \v17.58  = ~v5 & new_n195_;
  assign new_n865_ = ~new_n251_ & ~new_n371_;
  assign new_n866_ = ~v6 & ~new_n865_;
  assign new_n867_ = ~v3 & new_n866_;
  assign new_n868_ = ~v1 & new_n867_;
  assign new_n869_ = v3 & new_n357_;
  assign new_n870_ = new_n123_ & new_n869_;
  assign new_n871_ = ~new_n868_ & ~new_n870_;
  assign new_n872_ = ~v4 & ~new_n871_;
  assign \v17.59  = ~v0 & new_n872_;
  assign new_n874_ = v1 & ~v2;
  assign new_n875_ = new_n364_ & new_n874_;
  assign new_n876_ = ~new_n351_ & ~new_n875_;
  assign new_n877_ = v6 & ~new_n876_;
  assign new_n878_ = ~v3 & new_n877_;
  assign \v17.60  = ~v0 & new_n878_;
  assign \v17.61  = 1'b0;
  assign \v17.62  = 1'b0;
  assign \v17.63  = 1'b0;
  assign \v17.64  = 1'b0;
  assign \v17.65  = 1'b0;
  assign \v17.66  = 1'b0;
  assign \v17.67  = 1'b0;
  assign \v17.68  = 1'b0;
endmodule


