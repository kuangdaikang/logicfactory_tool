// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:34 2022

module pope  ( 
    v0, v1, v2, v3, v4, v5,
    \v6.0 , \v6.1 , \v6.2 , \v6.3 , \v6.4 , \v6.5 , \v6.6 , \v6.7 , \v6.8 ,
    \v6.9 , \v6.10 , \v6.11 , \v6.12 , \v6.13 , \v6.14 , \v6.15 , \v6.16 ,
    \v6.17 , \v6.18 , \v6.19 , \v6.20 , \v6.21 , \v6.22 , \v6.23 , \v6.24 ,
    \v6.25 , \v6.26 , \v6.27 , \v6.28 , \v6.29 , \v6.30 , \v6.31 , \v6.32 ,
    \v6.33 , \v6.34 , \v6.35 , \v6.36 , \v6.37 , \v6.38 , \v6.39 , \v6.40 ,
    \v6.41 , \v6.42 , \v6.43 , \v6.44 , \v6.45 , \v6.46 , \v6.47   );
  input  v0, v1, v2, v3, v4, v5;
  output \v6.0 , \v6.1 , \v6.2 , \v6.3 , \v6.4 , \v6.5 , \v6.6 , \v6.7 ,
    \v6.8 , \v6.9 , \v6.10 , \v6.11 , \v6.12 , \v6.13 , \v6.14 , \v6.15 ,
    \v6.16 , \v6.17 , \v6.18 , \v6.19 , \v6.20 , \v6.21 , \v6.22 , \v6.23 ,
    \v6.24 , \v6.25 , \v6.26 , \v6.27 , \v6.28 , \v6.29 , \v6.30 , \v6.31 ,
    \v6.32 , \v6.33 , \v6.34 , \v6.35 , \v6.36 , \v6.37 , \v6.38 , \v6.39 ,
    \v6.40 , \v6.41 , \v6.42 , \v6.43 , \v6.44 , \v6.45 , \v6.46 , \v6.47 ;
  wire new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_,
    new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_,
    new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n318_, new_n319_,
    new_n320_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n525_, new_n526_,
    new_n528_, new_n529_, new_n530_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n541_,
    new_n543_, new_n544_, new_n545_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n685_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_;
  assign new_n56_ = ~v3 & v4;
  assign new_n57_ = v3 & ~v4;
  assign new_n58_ = ~new_n56_ & ~new_n57_;
  assign new_n59_ = v1 & v2;
  assign new_n60_ = ~v1 & ~v2;
  assign new_n61_ = ~new_n59_ & ~new_n60_;
  assign new_n62_ = ~v1 & v2;
  assign new_n63_ = v1 & ~v2;
  assign new_n64_ = ~new_n62_ & ~new_n63_;
  assign new_n65_ = ~v0 & ~v5;
  assign new_n66_ = ~v0 & ~new_n65_;
  assign new_n67_ = ~new_n64_ & ~new_n66_;
  assign new_n68_ = new_n61_ & ~new_n67_;
  assign new_n69_ = ~new_n58_ & ~new_n68_;
  assign new_n70_ = v3 & v4;
  assign new_n71_ = ~v3 & ~v4;
  assign new_n72_ = ~new_n70_ & ~new_n71_;
  assign new_n73_ = ~v5 & ~new_n64_;
  assign new_n74_ = ~v0 & ~v1;
  assign new_n75_ = v2 & v5;
  assign new_n76_ = new_n74_ & new_n75_;
  assign new_n77_ = ~new_n73_ & ~new_n76_;
  assign new_n78_ = new_n61_ & new_n77_;
  assign new_n79_ = ~new_n72_ & ~new_n78_;
  assign new_n80_ = ~v2 & v4;
  assign new_n81_ = v1 & new_n80_;
  assign new_n82_ = v2 & ~v4;
  assign new_n83_ = ~v1 & new_n82_;
  assign new_n84_ = ~new_n81_ & ~new_n83_;
  assign new_n85_ = v5 & ~new_n84_;
  assign new_n86_ = v3 & new_n85_;
  assign new_n87_ = ~v0 & new_n86_;
  assign new_n88_ = ~new_n79_ & ~new_n87_;
  assign \v6.0  = new_n69_ | ~new_n88_;
  assign new_n90_ = v0 & new_n70_;
  assign new_n91_ = ~v0 & new_n71_;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign new_n93_ = ~v2 & ~new_n92_;
  assign new_n94_ = v0 & new_n71_;
  assign new_n95_ = ~v4 & ~new_n94_;
  assign new_n96_ = v2 & ~new_n95_;
  assign new_n97_ = ~new_n93_ & ~new_n96_;
  assign new_n98_ = new_n58_ & ~new_n94_;
  assign new_n99_ = ~v2 & ~new_n98_;
  assign new_n100_ = v0 & v2;
  assign new_n101_ = new_n57_ & new_n100_;
  assign new_n102_ = ~new_n99_ & ~new_n101_;
  assign new_n103_ = v5 & ~new_n102_;
  assign new_n104_ = new_n97_ & ~new_n103_;
  assign new_n105_ = ~v0 & v1;
  assign new_n106_ = new_n75_ & new_n105_;
  assign new_n107_ = v0 & ~v1;
  assign new_n108_ = ~v2 & ~v5;
  assign new_n109_ = new_n107_ & new_n108_;
  assign new_n110_ = ~new_n106_ & ~new_n109_;
  assign new_n111_ = v3 & ~v5;
  assign new_n112_ = ~v2 & new_n111_;
  assign new_n113_ = new_n105_ & new_n112_;
  assign new_n114_ = new_n110_ & ~new_n113_;
  assign new_n115_ = ~v4 & ~new_n114_;
  assign new_n116_ = v3 & v5;
  assign new_n117_ = ~v1 & new_n116_;
  assign new_n118_ = ~v3 & ~v5;
  assign new_n119_ = v1 & new_n118_;
  assign new_n120_ = ~new_n117_ & ~new_n119_;
  assign new_n121_ = ~v0 & ~new_n120_;
  assign new_n122_ = v0 & v1;
  assign new_n123_ = new_n118_ & new_n122_;
  assign new_n124_ = ~new_n121_ & ~new_n123_;
  assign new_n125_ = v4 & ~new_n124_;
  assign new_n126_ = ~v2 & new_n125_;
  assign new_n127_ = ~new_n115_ & ~new_n126_;
  assign \v6.1  = ~new_n104_ | ~new_n127_;
  assign new_n129_ = ~v2 & v3;
  assign new_n130_ = ~v1 & new_n129_;
  assign new_n131_ = v2 & ~v3;
  assign new_n132_ = v1 & new_n131_;
  assign new_n133_ = ~new_n130_ & ~new_n132_;
  assign new_n134_ = ~v0 & ~v4;
  assign new_n135_ = ~v0 & ~new_n134_;
  assign new_n136_ = ~new_n133_ & ~new_n135_;
  assign new_n137_ = ~new_n74_ & ~new_n122_;
  assign new_n138_ = v2 & v3;
  assign new_n139_ = ~v2 & ~v3;
  assign new_n140_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = ~new_n137_ & ~new_n140_;
  assign new_n142_ = v1 & v3;
  assign new_n143_ = ~v1 & ~v3;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = ~v0 & ~new_n144_;
  assign new_n146_ = ~v1 & v3;
  assign new_n147_ = v0 & new_n146_;
  assign new_n148_ = ~new_n145_ & ~new_n147_;
  assign new_n149_ = v2 & ~new_n148_;
  assign new_n150_ = ~new_n141_ & ~new_n149_;
  assign new_n151_ = ~v4 & ~new_n150_;
  assign new_n152_ = ~v1 & ~new_n60_;
  assign new_n153_ = v3 & ~new_n152_;
  assign new_n154_ = ~v1 & new_n139_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = v4 & ~new_n155_;
  assign new_n157_ = ~v0 & new_n156_;
  assign new_n158_ = ~new_n151_ & ~new_n157_;
  assign new_n159_ = ~new_n136_ & new_n158_;
  assign new_n160_ = v1 & ~new_n58_;
  assign new_n161_ = v0 & new_n143_;
  assign new_n162_ = ~new_n160_ & ~new_n161_;
  assign new_n163_ = ~v5 & ~new_n162_;
  assign new_n164_ = v4 & v5;
  assign new_n165_ = v3 & new_n164_;
  assign new_n166_ = new_n122_ & new_n165_;
  assign new_n167_ = ~new_n163_ & ~new_n166_;
  assign new_n168_ = ~v2 & ~new_n167_;
  assign new_n169_ = ~v3 & v5;
  assign new_n170_ = ~new_n111_ & ~new_n169_;
  assign new_n171_ = ~v1 & ~new_n170_;
  assign new_n172_ = v1 & new_n116_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_ = v4 & ~new_n173_;
  assign new_n175_ = ~v4 & v5;
  assign new_n176_ = new_n143_ & new_n175_;
  assign new_n177_ = ~new_n174_ & ~new_n176_;
  assign new_n178_ = v0 & ~new_n177_;
  assign new_n179_ = new_n74_ & new_n165_;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = v2 & ~new_n180_;
  assign new_n182_ = ~new_n168_ & ~new_n181_;
  assign \v6.2  = ~new_n159_ | ~new_n182_;
  assign new_n184_ = ~new_n116_ & ~new_n118_;
  assign new_n185_ = v0 & ~new_n61_;
  assign new_n186_ = ~new_n74_ & ~new_n185_;
  assign new_n187_ = ~new_n184_ & ~new_n186_;
  assign new_n188_ = ~v0 & ~new_n61_;
  assign new_n189_ = v0 & new_n60_;
  assign new_n190_ = ~new_n188_ & ~new_n189_;
  assign new_n191_ = ~new_n170_ & ~new_n190_;
  assign new_n192_ = ~v0 & v3;
  assign new_n193_ = v0 & ~v3;
  assign new_n194_ = ~new_n192_ & ~new_n193_;
  assign new_n195_ = v2 & ~new_n194_;
  assign new_n196_ = v0 & ~v2;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = v5 & ~new_n197_;
  assign new_n199_ = ~v0 & new_n108_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = v1 & ~new_n200_;
  assign new_n202_ = v2 & new_n111_;
  assign new_n203_ = new_n107_ & new_n202_;
  assign new_n204_ = ~new_n201_ & ~new_n203_;
  assign new_n205_ = ~new_n191_ & new_n204_;
  assign new_n206_ = ~new_n187_ & new_n205_;
  assign new_n207_ = ~v1 & new_n75_;
  assign new_n208_ = v1 & new_n108_;
  assign new_n209_ = ~new_n207_ & ~new_n208_;
  assign new_n210_ = ~new_n58_ & ~new_n209_;
  assign new_n211_ = ~v1 & new_n56_;
  assign new_n212_ = v1 & new_n57_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~v5 & ~new_n213_;
  assign new_n215_ = v2 & new_n214_;
  assign new_n216_ = ~new_n210_ & ~new_n215_;
  assign new_n217_ = v0 & ~new_n216_;
  assign new_n218_ = new_n129_ & new_n164_;
  assign new_n219_ = ~v4 & ~v5;
  assign new_n220_ = new_n131_ & new_n219_;
  assign new_n221_ = ~new_n218_ & ~new_n220_;
  assign new_n222_ = v1 & ~new_n221_;
  assign new_n223_ = ~v4 & ~new_n170_;
  assign new_n224_ = v2 & new_n223_;
  assign new_n225_ = ~v1 & new_n224_;
  assign new_n226_ = ~new_n222_ & ~new_n225_;
  assign new_n227_ = ~v0 & ~new_n226_;
  assign new_n228_ = ~new_n217_ & ~new_n227_;
  assign \v6.3  = ~new_n206_ | ~new_n228_;
  assign new_n230_ = v2 & new_n175_;
  assign new_n231_ = v4 & ~v5;
  assign new_n232_ = ~v2 & new_n231_;
  assign new_n233_ = ~new_n230_ & ~new_n232_;
  assign new_n234_ = v1 & ~v3;
  assign new_n235_ = ~v0 & new_n234_;
  assign new_n236_ = ~v0 & ~new_n235_;
  assign new_n237_ = ~new_n233_ & ~new_n236_;
  assign new_n238_ = new_n56_ & new_n59_;
  assign new_n239_ = new_n57_ & new_n60_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = v0 & ~new_n240_;
  assign new_n242_ = v1 & new_n138_;
  assign new_n243_ = ~new_n60_ & ~new_n242_;
  assign new_n244_ = ~v0 & ~new_n243_;
  assign new_n245_ = ~new_n241_ & ~new_n244_;
  assign new_n246_ = ~new_n164_ & ~new_n219_;
  assign new_n247_ = v3 & ~new_n246_;
  assign new_n248_ = ~v3 & new_n219_;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = ~new_n137_ & ~new_n249_;
  assign new_n251_ = ~v3 & new_n164_;
  assign new_n252_ = ~new_n111_ & ~new_n251_;
  assign new_n253_ = ~v1 & ~new_n252_;
  assign new_n254_ = v0 & new_n253_;
  assign new_n255_ = ~new_n250_ & ~new_n254_;
  assign new_n256_ = v2 & ~new_n255_;
  assign new_n257_ = ~v1 & ~new_n143_;
  assign new_n258_ = ~v5 & ~new_n257_;
  assign new_n259_ = ~v4 & new_n258_;
  assign new_n260_ = new_n146_ & new_n164_;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = v0 & ~new_n261_;
  assign new_n263_ = v3 & new_n219_;
  assign new_n264_ = new_n105_ & new_n263_;
  assign new_n265_ = ~new_n262_ & ~new_n264_;
  assign new_n266_ = ~v2 & ~new_n265_;
  assign new_n267_ = ~new_n256_ & ~new_n266_;
  assign new_n268_ = new_n245_ & new_n267_;
  assign \v6.4  = new_n237_ | ~new_n268_;
  assign new_n270_ = ~new_n146_ & ~new_n234_;
  assign new_n271_ = v0 & ~new_n270_;
  assign new_n272_ = ~v0 & new_n142_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = v2 & ~new_n273_;
  assign new_n275_ = new_n107_ & new_n129_;
  assign new_n276_ = ~new_n274_ & ~new_n275_;
  assign new_n277_ = ~new_n141_ & new_n276_;
  assign new_n278_ = ~v4 & ~new_n277_;
  assign new_n279_ = ~v0 & ~new_n192_;
  assign new_n280_ = v2 & ~new_n279_;
  assign new_n281_ = ~v0 & new_n129_;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = v1 & ~new_n282_;
  assign new_n284_ = ~new_n129_ & ~new_n131_;
  assign new_n285_ = ~v1 & ~new_n284_;
  assign new_n286_ = v0 & new_n285_;
  assign new_n287_ = ~new_n283_ & ~new_n286_;
  assign new_n288_ = v4 & ~new_n287_;
  assign new_n289_ = ~new_n278_ & ~new_n288_;
  assign new_n290_ = v0 & ~new_n184_;
  assign new_n291_ = ~v0 & new_n118_;
  assign new_n292_ = ~new_n290_ & ~new_n291_;
  assign new_n293_ = v4 & ~new_n292_;
  assign new_n294_ = ~v0 & new_n219_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = v1 & ~new_n295_;
  assign new_n297_ = ~v3 & ~new_n56_;
  assign new_n298_ = v5 & ~new_n297_;
  assign new_n299_ = ~v0 & new_n298_;
  assign new_n300_ = new_n193_ & new_n219_;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = ~v1 & ~new_n301_;
  assign new_n303_ = ~new_n296_ & ~new_n302_;
  assign new_n304_ = ~v2 & ~new_n303_;
  assign new_n305_ = ~new_n175_ & ~new_n231_;
  assign new_n306_ = v1 & ~new_n305_;
  assign new_n307_ = ~v1 & new_n175_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = ~v3 & ~new_n308_;
  assign new_n310_ = ~new_n260_ & ~new_n309_;
  assign new_n311_ = ~v0 & ~new_n310_;
  assign new_n312_ = v3 & new_n231_;
  assign new_n313_ = new_n107_ & new_n312_;
  assign new_n314_ = ~new_n311_ & ~new_n313_;
  assign new_n315_ = v2 & ~new_n314_;
  assign new_n316_ = ~new_n304_ & ~new_n315_;
  assign \v6.5  = ~new_n289_ | ~new_n316_;
  assign new_n318_ = ~v2 & new_n122_;
  assign new_n319_ = v3 & new_n318_;
  assign new_n320_ = v4 & new_n319_;
  assign \v6.6  = v5 & new_n320_;
  assign new_n322_ = ~v0 & new_n82_;
  assign new_n323_ = ~new_n196_ & ~new_n322_;
  assign new_n324_ = ~v1 & v4;
  assign new_n325_ = v1 & ~v4;
  assign new_n326_ = ~new_n324_ & ~new_n325_;
  assign new_n327_ = ~v2 & ~new_n326_;
  assign new_n328_ = ~v0 & new_n327_;
  assign new_n329_ = v2 & v4;
  assign new_n330_ = new_n107_ & new_n329_;
  assign new_n331_ = ~new_n328_ & ~new_n330_;
  assign new_n332_ = new_n323_ & new_n331_;
  assign new_n333_ = ~new_n170_ & ~new_n332_;
  assign new_n334_ = v1 & v4;
  assign new_n335_ = ~v0 & new_n334_;
  assign new_n336_ = ~v1 & ~v4;
  assign new_n337_ = v0 & new_n336_;
  assign new_n338_ = ~new_n335_ & ~new_n337_;
  assign new_n339_ = new_n184_ & ~new_n202_;
  assign new_n340_ = ~new_n338_ & ~new_n339_;
  assign new_n341_ = v0 & new_n59_;
  assign new_n342_ = ~v0 & new_n60_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = ~new_n184_ & ~new_n343_;
  assign new_n345_ = v5 & ~new_n284_;
  assign new_n346_ = v1 & new_n345_;
  assign new_n347_ = v0 & new_n346_;
  assign new_n348_ = ~new_n344_ & ~new_n347_;
  assign new_n349_ = v0 & new_n324_;
  assign new_n350_ = ~v0 & new_n325_;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign new_n352_ = ~new_n184_ & ~new_n351_;
  assign new_n353_ = ~new_n334_ & ~new_n336_;
  assign new_n354_ = v5 & ~new_n353_;
  assign new_n355_ = ~v0 & new_n354_;
  assign new_n356_ = new_n122_ & new_n231_;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_ = ~v3 & ~new_n357_;
  assign new_n359_ = ~new_n352_ & ~new_n358_;
  assign new_n360_ = ~v2 & ~new_n359_;
  assign new_n361_ = ~new_n212_ & ~new_n324_;
  assign new_n362_ = v5 & ~new_n361_;
  assign new_n363_ = new_n143_ & new_n219_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = v2 & ~new_n364_;
  assign new_n366_ = ~v0 & new_n365_;
  assign new_n367_ = ~new_n360_ & ~new_n366_;
  assign new_n368_ = new_n348_ & new_n367_;
  assign new_n369_ = ~new_n340_ & new_n368_;
  assign \v6.7  = new_n333_ | ~new_n369_;
  assign new_n371_ = ~v0 & ~new_n105_;
  assign new_n372_ = v2 & ~new_n371_;
  assign new_n373_ = ~new_n342_ & ~new_n372_;
  assign new_n374_ = v5 & ~new_n373_;
  assign new_n375_ = v2 & ~v5;
  assign new_n376_ = new_n122_ & new_n375_;
  assign new_n377_ = ~new_n374_ & ~new_n376_;
  assign new_n378_ = ~v0 & new_n75_;
  assign new_n379_ = ~new_n196_ & ~new_n378_;
  assign new_n380_ = ~v1 & ~new_n379_;
  assign new_n381_ = new_n105_ & new_n108_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = v3 & ~new_n382_;
  assign new_n384_ = ~v2 & new_n118_;
  assign new_n385_ = new_n122_ & new_n384_;
  assign new_n386_ = ~new_n383_ & ~new_n385_;
  assign new_n387_ = new_n377_ & new_n386_;
  assign new_n388_ = ~v2 & ~v4;
  assign new_n389_ = ~new_n329_ & ~new_n388_;
  assign new_n390_ = ~v0 & ~new_n389_;
  assign new_n391_ = v0 & new_n329_;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = new_n71_ & new_n196_;
  assign new_n394_ = new_n392_ & ~new_n393_;
  assign new_n395_ = ~v1 & ~new_n394_;
  assign new_n396_ = v2 & ~new_n72_;
  assign new_n397_ = ~v2 & new_n56_;
  assign new_n398_ = ~new_n396_ & ~new_n397_;
  assign new_n399_ = v1 & ~new_n398_;
  assign new_n400_ = ~v0 & new_n399_;
  assign new_n401_ = ~new_n395_ & ~new_n400_;
  assign new_n402_ = ~v5 & ~new_n401_;
  assign \v6.8  = ~new_n387_ | new_n402_;
  assign new_n404_ = ~v0 & ~new_n284_;
  assign new_n405_ = new_n140_ & ~new_n404_;
  assign new_n406_ = ~v1 & ~new_n405_;
  assign new_n407_ = v0 & new_n138_;
  assign new_n408_ = ~new_n404_ & ~new_n407_;
  assign new_n409_ = v1 & ~new_n408_;
  assign new_n410_ = ~new_n406_ & ~new_n409_;
  assign new_n411_ = ~v1 & ~new_n62_;
  assign new_n412_ = ~v3 & ~new_n411_;
  assign new_n413_ = ~new_n130_ & ~new_n412_;
  assign new_n414_ = v0 & ~new_n413_;
  assign new_n415_ = new_n105_ & new_n138_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = v5 & ~new_n416_;
  assign new_n418_ = new_n410_ & ~new_n417_;
  assign new_n419_ = v2 & new_n57_;
  assign new_n420_ = ~new_n397_ & ~new_n419_;
  assign new_n421_ = ~v0 & ~new_n420_;
  assign new_n422_ = v2 & new_n56_;
  assign new_n423_ = ~new_n388_ & ~new_n422_;
  assign new_n424_ = v0 & ~new_n423_;
  assign new_n425_ = ~new_n421_ & ~new_n424_;
  assign new_n426_ = v1 & ~new_n425_;
  assign new_n427_ = new_n107_ & new_n422_;
  assign new_n428_ = ~new_n426_ & ~new_n427_;
  assign new_n429_ = ~v5 & ~new_n428_;
  assign \v6.9  = ~new_n418_ | new_n429_;
  assign new_n431_ = v1 & ~new_n389_;
  assign new_n432_ = ~new_n83_ & ~new_n431_;
  assign new_n433_ = ~v5 & ~new_n432_;
  assign new_n434_ = ~new_n207_ & ~new_n433_;
  assign new_n435_ = ~v3 & ~new_n434_;
  assign new_n436_ = new_n62_ & new_n312_;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = v0 & ~new_n437_;
  assign new_n439_ = v4 & ~new_n164_;
  assign new_n440_ = v3 & ~new_n439_;
  assign new_n441_ = v2 & new_n440_;
  assign new_n442_ = ~v1 & new_n441_;
  assign new_n443_ = ~v0 & new_n442_;
  assign \v6.10  = new_n438_ | new_n443_;
  assign new_n445_ = ~v2 & v5;
  assign new_n446_ = v0 & new_n445_;
  assign new_n447_ = ~v0 & v2;
  assign new_n448_ = new_n219_ & new_n447_;
  assign new_n449_ = ~new_n446_ & ~new_n448_;
  assign new_n450_ = ~v3 & ~new_n449_;
  assign \v6.11  = v1 & new_n450_;
  assign new_n452_ = ~v0 & ~v2;
  assign new_n453_ = new_n70_ & new_n452_;
  assign new_n454_ = new_n71_ & new_n100_;
  assign new_n455_ = ~new_n453_ & ~new_n454_;
  assign new_n456_ = ~v1 & v5;
  assign new_n457_ = ~v1 & ~new_n456_;
  assign new_n458_ = ~new_n455_ & ~new_n457_;
  assign new_n459_ = v0 & new_n129_;
  assign new_n460_ = new_n140_ & ~new_n459_;
  assign new_n461_ = v5 & ~new_n460_;
  assign new_n462_ = ~new_n199_ & ~new_n461_;
  assign new_n463_ = v4 & ~new_n170_;
  assign new_n464_ = v2 & new_n463_;
  assign new_n465_ = new_n139_ & new_n219_;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign new_n467_ = v0 & ~new_n466_;
  assign new_n468_ = v3 & new_n175_;
  assign new_n469_ = new_n452_ & new_n468_;
  assign new_n470_ = ~new_n467_ & ~new_n469_;
  assign new_n471_ = new_n462_ & new_n470_;
  assign new_n472_ = ~v1 & ~new_n471_;
  assign new_n473_ = v0 & v3;
  assign new_n474_ = v0 & ~new_n473_;
  assign new_n475_ = v0 & new_n56_;
  assign new_n476_ = new_n474_ & ~new_n475_;
  assign new_n477_ = v2 & ~new_n476_;
  assign new_n478_ = new_n57_ & new_n452_;
  assign new_n479_ = ~new_n477_ & ~new_n478_;
  assign new_n480_ = v5 & ~new_n479_;
  assign new_n481_ = v1 & new_n480_;
  assign new_n482_ = ~new_n472_ & ~new_n481_;
  assign \v6.12  = new_n458_ | ~new_n482_;
  assign new_n484_ = v0 & v5;
  assign new_n485_ = v0 & ~new_n484_;
  assign new_n486_ = ~new_n284_ & ~new_n485_;
  assign new_n487_ = new_n140_ & ~new_n486_;
  assign new_n488_ = ~new_n326_ & ~new_n487_;
  assign new_n489_ = ~v0 & ~new_n447_;
  assign new_n490_ = ~v0 & new_n139_;
  assign new_n491_ = new_n489_ & ~new_n490_;
  assign new_n492_ = new_n116_ & new_n452_;
  assign new_n493_ = new_n491_ & ~new_n492_;
  assign new_n494_ = ~new_n353_ & ~new_n493_;
  assign new_n495_ = new_n56_ & new_n62_;
  assign new_n496_ = new_n57_ & new_n63_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = ~v5 & ~new_n497_;
  assign new_n499_ = v0 & new_n498_;
  assign new_n500_ = ~new_n494_ & ~new_n499_;
  assign \v6.13  = new_n488_ | ~new_n500_;
  assign new_n502_ = v1 & new_n75_;
  assign new_n503_ = ~new_n60_ & ~new_n502_;
  assign new_n504_ = new_n105_ & new_n445_;
  assign new_n505_ = new_n503_ & ~new_n504_;
  assign new_n506_ = v5 & ~new_n64_;
  assign new_n507_ = v0 & new_n506_;
  assign new_n508_ = new_n105_ & new_n375_;
  assign new_n509_ = ~new_n507_ & ~new_n508_;
  assign new_n510_ = v3 & ~new_n509_;
  assign new_n511_ = ~v3 & ~new_n209_;
  assign new_n512_ = ~v0 & new_n511_;
  assign new_n513_ = ~new_n510_ & ~new_n512_;
  assign new_n514_ = new_n505_ & new_n513_;
  assign new_n515_ = ~new_n80_ & ~new_n82_;
  assign new_n516_ = v1 & ~new_n515_;
  assign new_n517_ = new_n57_ & new_n62_;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign new_n519_ = v0 & ~new_n518_;
  assign new_n520_ = ~v2 & new_n70_;
  assign new_n521_ = new_n105_ & new_n520_;
  assign new_n522_ = ~new_n519_ & ~new_n521_;
  assign new_n523_ = ~v5 & ~new_n522_;
  assign \v6.14  = ~new_n514_ | new_n523_;
  assign new_n525_ = v2 & new_n169_;
  assign new_n526_ = ~v1 & new_n525_;
  assign \v6.15  = v0 & new_n526_;
  assign new_n528_ = v2 & new_n122_;
  assign new_n529_ = v3 & new_n528_;
  assign new_n530_ = v4 & new_n529_;
  assign \v6.16  = ~v5 & new_n530_;
  assign new_n532_ = new_n60_ & new_n70_;
  assign new_n533_ = new_n59_ & new_n71_;
  assign new_n534_ = ~new_n532_ & ~new_n533_;
  assign new_n535_ = v0 & ~new_n534_;
  assign new_n536_ = v3 & ~new_n353_;
  assign new_n537_ = ~v2 & new_n536_;
  assign new_n538_ = ~v0 & new_n537_;
  assign new_n539_ = ~new_n535_ & ~new_n538_;
  assign \v6.17  = ~v5 & ~new_n539_;
  assign new_n541_ = ~v5 & ~new_n534_;
  assign \v6.18  = v0 & new_n541_;
  assign new_n543_ = ~v2 & new_n107_;
  assign new_n544_ = v3 & new_n543_;
  assign new_n545_ = v4 & new_n544_;
  assign \v6.19  = ~v5 & new_n545_;
  assign new_n547_ = ~v0 & v4;
  assign new_n548_ = v0 & ~v4;
  assign new_n549_ = ~new_n547_ & ~new_n548_;
  assign new_n550_ = ~v0 & new_n57_;
  assign new_n551_ = new_n549_ & ~new_n550_;
  assign new_n552_ = ~new_n61_ & ~new_n551_;
  assign new_n553_ = v0 & new_n62_;
  assign new_n554_ = ~v0 & new_n63_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = v0 & new_n431_;
  assign new_n557_ = new_n74_ & new_n82_;
  assign new_n558_ = ~new_n556_ & ~new_n557_;
  assign new_n559_ = new_n555_ & new_n558_;
  assign new_n560_ = v3 & ~new_n559_;
  assign new_n561_ = ~v1 & ~new_n392_;
  assign new_n562_ = v0 & new_n334_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = ~v3 & ~new_n563_;
  assign new_n565_ = ~new_n560_ & ~new_n564_;
  assign new_n566_ = ~new_n552_ & new_n565_;
  assign new_n567_ = ~v5 & ~new_n72_;
  assign new_n568_ = v1 & new_n567_;
  assign new_n569_ = ~v1 & new_n164_;
  assign new_n570_ = ~new_n568_ & ~new_n569_;
  assign new_n571_ = ~v2 & ~new_n570_;
  assign new_n572_ = ~v3 & new_n175_;
  assign new_n573_ = new_n62_ & new_n572_;
  assign new_n574_ = ~new_n571_ & ~new_n573_;
  assign new_n575_ = v0 & ~new_n574_;
  assign new_n576_ = ~new_n75_ & ~new_n108_;
  assign new_n577_ = v1 & ~new_n576_;
  assign new_n578_ = ~v1 & new_n375_;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign new_n580_ = ~v4 & ~new_n579_;
  assign new_n581_ = ~v3 & new_n580_;
  assign new_n582_ = new_n62_ & new_n165_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = ~v0 & ~new_n583_;
  assign new_n585_ = ~new_n575_ & ~new_n584_;
  assign \v6.20  = ~new_n566_ | ~new_n585_;
  assign new_n587_ = ~new_n196_ & ~new_n447_;
  assign new_n588_ = ~new_n100_ & ~new_n452_;
  assign new_n589_ = v3 & ~new_n588_;
  assign new_n590_ = new_n587_ & ~new_n589_;
  assign new_n591_ = ~new_n353_ & ~new_n590_;
  assign new_n592_ = ~new_n100_ & ~new_n281_;
  assign new_n593_ = ~new_n326_ & ~new_n592_;
  assign new_n594_ = ~new_n475_ & ~new_n550_;
  assign new_n595_ = v2 & ~new_n594_;
  assign new_n596_ = v1 & new_n595_;
  assign new_n597_ = ~v0 & new_n154_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~new_n593_ & new_n598_;
  assign new_n600_ = ~new_n591_ & new_n599_;
  assign new_n601_ = v1 & new_n219_;
  assign new_n602_ = ~new_n569_ & ~new_n601_;
  assign new_n603_ = ~v2 & ~new_n602_;
  assign new_n604_ = ~new_n573_ & ~new_n603_;
  assign new_n605_ = v0 & ~new_n604_;
  assign new_n606_ = ~v4 & ~new_n576_;
  assign new_n607_ = v1 & new_n606_;
  assign new_n608_ = new_n62_ & new_n231_;
  assign new_n609_ = ~new_n607_ & ~new_n608_;
  assign new_n610_ = ~v3 & ~new_n609_;
  assign new_n611_ = ~new_n582_ & ~new_n610_;
  assign new_n612_ = ~v0 & ~new_n611_;
  assign new_n613_ = ~new_n605_ & ~new_n612_;
  assign \v6.21  = ~new_n600_ | ~new_n613_;
  assign new_n615_ = v0 & ~new_n353_;
  assign new_n616_ = ~new_n74_ & ~new_n615_;
  assign new_n617_ = v2 & ~new_n616_;
  assign new_n618_ = new_n122_ & new_n388_;
  assign new_n619_ = ~new_n617_ & ~new_n618_;
  assign new_n620_ = ~v5 & ~new_n619_;
  assign new_n621_ = v0 & ~new_n107_;
  assign new_n622_ = v5 & ~new_n621_;
  assign new_n623_ = v4 & new_n622_;
  assign new_n624_ = ~v2 & new_n623_;
  assign new_n625_ = ~new_n620_ & ~new_n624_;
  assign new_n626_ = v5 & ~new_n58_;
  assign new_n627_ = ~v0 & ~v3;
  assign new_n628_ = new_n231_ & new_n627_;
  assign new_n629_ = ~new_n626_ & ~new_n628_;
  assign new_n630_ = v2 & ~new_n629_;
  assign new_n631_ = v0 & new_n164_;
  assign new_n632_ = ~new_n65_ & ~new_n631_;
  assign new_n633_ = v3 & ~new_n632_;
  assign new_n634_ = ~v2 & new_n633_;
  assign new_n635_ = ~new_n630_ & ~new_n634_;
  assign new_n636_ = v1 & ~new_n635_;
  assign new_n637_ = ~v0 & ~new_n233_;
  assign new_n638_ = new_n100_ & new_n175_;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign new_n640_ = v3 & ~new_n639_;
  assign new_n641_ = v0 & new_n422_;
  assign new_n642_ = ~new_n640_ & ~new_n641_;
  assign new_n643_ = ~v1 & ~new_n642_;
  assign new_n644_ = ~new_n636_ & ~new_n643_;
  assign \v6.22  = ~new_n625_ | ~new_n644_;
  assign new_n646_ = ~new_n184_ & ~new_n389_;
  assign new_n647_ = ~new_n312_ & ~new_n572_;
  assign new_n648_ = ~v2 & ~new_n647_;
  assign new_n649_ = ~v0 & new_n648_;
  assign new_n650_ = new_n100_ & new_n572_;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = ~new_n646_ & new_n651_;
  assign new_n653_ = v1 & new_n129_;
  assign new_n654_ = ~new_n62_ & ~new_n653_;
  assign new_n655_ = ~v4 & ~new_n654_;
  assign new_n656_ = v4 & ~new_n137_;
  assign new_n657_ = v3 & new_n656_;
  assign new_n658_ = v2 & new_n657_;
  assign new_n659_ = ~new_n655_ & ~new_n658_;
  assign new_n660_ = ~v5 & ~new_n659_;
  assign new_n661_ = ~v0 & new_n59_;
  assign new_n662_ = ~new_n189_ & ~new_n661_;
  assign new_n663_ = v5 & ~new_n662_;
  assign new_n664_ = ~v4 & new_n663_;
  assign new_n665_ = ~v3 & new_n664_;
  assign new_n666_ = ~new_n660_ & ~new_n665_;
  assign \v6.23  = ~new_n652_ | ~new_n666_;
  assign new_n668_ = ~new_n342_ & new_n371_;
  assign new_n669_ = new_n74_ & new_n138_;
  assign new_n670_ = new_n668_ & ~new_n669_;
  assign new_n671_ = new_n74_ & new_n422_;
  assign \v6.25  = ~new_n670_ | new_n671_;
  assign new_n673_ = ~v0 & ~new_n74_;
  assign new_n674_ = ~new_n661_ & new_n673_;
  assign new_n675_ = new_n105_ & new_n139_;
  assign new_n676_ = new_n674_ & ~new_n675_;
  assign \v6.26  = new_n521_ | ~new_n676_;
  assign new_n678_ = ~v4 & new_n544_;
  assign \v6.27  = ~v5 & new_n678_;
  assign new_n680_ = ~v0 & new_n62_;
  assign new_n681_ = new_n572_ & new_n680_;
  assign \v6.28  = \v6.25  | new_n681_;
  assign new_n683_ = new_n468_ & new_n554_;
  assign \v6.29  = \v6.26  | new_n683_;
  assign new_n685_ = new_n105_ & new_n129_;
  assign \v6.31  = ~new_n674_ | new_n685_;
  assign new_n687_ = ~v2 & ~new_n58_;
  assign \v6.32  = v1 & new_n687_;
  assign new_n689_ = ~new_n371_ & ~new_n389_;
  assign new_n690_ = ~v2 & ~new_n353_;
  assign new_n691_ = ~v0 & new_n690_;
  assign new_n692_ = new_n82_ & new_n122_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = ~new_n689_ & new_n693_;
  assign new_n695_ = new_n56_ & new_n447_;
  assign new_n696_ = new_n420_ & ~new_n695_;
  assign new_n697_ = ~v1 & ~new_n696_;
  assign new_n698_ = new_n122_ & new_n397_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign \v6.33  = ~new_n694_ | ~new_n699_;
  assign new_n701_ = v1 & ~new_n59_;
  assign new_n702_ = ~new_n58_ & ~new_n701_;
  assign \v6.34  = ~new_n72_ | new_n702_;
  assign new_n704_ = v2 & new_n70_;
  assign new_n705_ = ~v2 & new_n71_;
  assign \v6.35  = new_n704_ | new_n705_;
  assign new_n707_ = v1 & new_n82_;
  assign \v6.36  = new_n687_ | new_n707_;
  assign new_n709_ = ~new_n185_ & ~new_n452_;
  assign new_n710_ = new_n122_ & new_n129_;
  assign new_n711_ = new_n709_ & ~new_n710_;
  assign new_n712_ = ~v4 & ~new_n711_;
  assign new_n713_ = ~new_n140_ & ~new_n371_;
  assign new_n714_ = new_n74_ & new_n139_;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = v4 & ~new_n715_;
  assign \v6.37  = new_n712_ | new_n716_;
  assign new_n718_ = ~new_n196_ & ~new_n680_;
  assign new_n719_ = v4 & ~new_n718_;
  assign \v6.38  = v3 & new_n719_;
  assign new_n721_ = v2 & ~new_n673_;
  assign new_n722_ = ~new_n342_ & ~new_n721_;
  assign new_n723_ = ~new_n105_ & ~new_n107_;
  assign new_n724_ = ~v3 & ~new_n723_;
  assign new_n725_ = ~v2 & new_n724_;
  assign new_n726_ = new_n722_ & ~new_n725_;
  assign new_n727_ = ~v2 & ~new_n273_;
  assign new_n728_ = new_n105_ & new_n131_;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = ~v4 & ~new_n729_;
  assign new_n731_ = new_n105_ & new_n704_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign \v6.39  = ~new_n726_ | ~new_n732_;
  assign new_n734_ = v3 & ~new_n389_;
  assign new_n735_ = ~new_n139_ & ~new_n734_;
  assign new_n736_ = ~new_n82_ & ~new_n520_;
  assign new_n737_ = v1 & ~new_n736_;
  assign new_n738_ = new_n735_ & ~new_n737_;
  assign new_n739_ = new_n70_ & new_n196_;
  assign new_n740_ = ~new_n322_ & ~new_n739_;
  assign new_n741_ = ~v1 & ~new_n740_;
  assign new_n742_ = new_n105_ & new_n422_;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign \v6.40  = ~new_n738_ | ~new_n743_;
  assign new_n745_ = ~new_n554_ & new_n673_;
  assign new_n746_ = ~new_n58_ & ~new_n745_;
  assign \v6.41  = ~new_n72_ | new_n746_;
  assign \v6.42  = ~v0 & new_n707_;
  assign new_n749_ = v3 & ~new_n515_;
  assign new_n750_ = ~new_n131_ & ~new_n749_;
  assign new_n751_ = v1 & ~new_n750_;
  assign new_n752_ = ~v0 & new_n751_;
  assign \v6.43  = new_n427_ | new_n752_;
  assign new_n754_ = ~new_n342_ & new_n587_;
  assign new_n755_ = new_n122_ & new_n138_;
  assign new_n756_ = new_n754_ & ~new_n755_;
  assign new_n757_ = ~new_n100_ & ~new_n554_;
  assign new_n758_ = ~v4 & ~new_n757_;
  assign new_n759_ = ~v3 & new_n758_;
  assign new_n760_ = new_n107_ & new_n704_;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign \v6.45  = ~new_n756_ | ~new_n761_;
  assign new_n763_ = ~new_n140_ & ~new_n673_;
  assign new_n764_ = new_n284_ & ~new_n490_;
  assign new_n765_ = v1 & ~new_n764_;
  assign new_n766_ = ~new_n275_ & ~new_n765_;
  assign new_n767_ = ~new_n763_ & new_n766_;
  assign new_n768_ = ~v4 & ~new_n284_;
  assign new_n769_ = ~v1 & new_n768_;
  assign new_n770_ = new_n59_ & new_n70_;
  assign new_n771_ = ~new_n769_ & ~new_n770_;
  assign new_n772_ = ~v0 & ~new_n771_;
  assign \v6.46  = ~new_n767_ | new_n772_;
  assign new_n774_ = new_n70_ & new_n107_;
  assign new_n775_ = new_n71_ & new_n105_;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign \v6.47  = ~v2 & ~new_n776_;
  assign \v6.24  = 1'b1;
  assign \v6.30  = 1'b0;
  assign \v6.44  = \v6.43 ;
endmodule


